magic
tech c035u
timestamp 1394208763
<< metal1 >>
rect 135 1573 191 1585
rect 205 1573 839 1585
rect 853 1573 1679 1585
rect 1693 1573 2495 1585
rect 2509 1573 3287 1585
rect 3301 1573 4103 1585
rect 4117 1573 4871 1585
rect 4885 1573 5663 1585
rect 85 1551 599 1561
rect 613 1551 1439 1561
rect 1453 1551 2375 1561
rect 2389 1551 3167 1561
rect 3181 1551 3887 1561
rect 3901 1551 4655 1561
rect 4669 1551 5543 1561
rect 61 1529 575 1539
rect 589 1529 1559 1539
rect 1573 1529 2279 1539
rect 2293 1529 3047 1539
rect 3061 1529 3983 1539
rect 3997 1529 4631 1539
rect 4645 1529 5423 1539
rect 37 1506 719 1516
rect 733 1506 1415 1516
rect 1429 1506 2255 1516
rect 2269 1506 3023 1516
rect 3037 1506 3863 1516
rect 3877 1506 4751 1516
rect 4765 1506 5399 1516
rect 493 1483 1199 1493
rect 1213 1483 2039 1493
rect 2053 1483 2927 1493
rect 2941 1483 3767 1493
rect 3781 1483 4439 1493
rect 4453 1483 5207 1493
rect 5221 1483 6143 1493
rect 469 1461 1175 1471
rect 1189 1461 2159 1471
rect 2173 1461 2831 1471
rect 2845 1461 3647 1471
rect 3661 1461 4535 1471
rect 4549 1461 5183 1471
rect 5197 1461 6023 1471
rect 445 1438 1319 1448
rect 1333 1438 2015 1448
rect 2029 1438 2807 1448
rect 2821 1438 3623 1448
rect 3637 1438 4415 1448
rect 4429 1438 5303 1448
rect 5317 1438 5999 1448
rect 349 1415 959 1425
rect 973 1415 1799 1425
rect 1813 1415 2711 1425
rect 2725 1415 3527 1425
rect 3541 1415 4223 1425
rect 4237 1415 4991 1425
rect 5005 1415 5903 1425
rect 325 1393 935 1403
rect 949 1393 1919 1403
rect 1933 1393 2615 1403
rect 2629 1393 3407 1403
rect 3421 1393 4319 1403
rect 4333 1393 4967 1403
rect 4981 1393 5783 1403
rect 301 1370 1079 1380
rect 1093 1370 1775 1380
rect 1789 1370 2591 1380
rect 2605 1370 3383 1380
rect 3397 1370 4199 1380
rect 4213 1370 5087 1380
rect 5101 1370 5759 1380
<< m2contact >>
rect 121 1573 135 1587
rect 191 1572 205 1586
rect 839 1572 853 1586
rect 1679 1572 1693 1586
rect 2495 1572 2509 1586
rect 3287 1572 3301 1586
rect 4103 1572 4117 1586
rect 4871 1572 4885 1586
rect 5663 1572 5677 1586
rect 71 1549 85 1563
rect 599 1549 613 1563
rect 1439 1549 1453 1563
rect 2375 1549 2389 1563
rect 3167 1549 3181 1563
rect 3887 1549 3901 1563
rect 4655 1549 4669 1563
rect 5543 1549 5557 1563
rect 47 1527 61 1541
rect 575 1527 589 1541
rect 1559 1527 1573 1541
rect 2279 1527 2293 1541
rect 3047 1527 3061 1541
rect 3983 1527 3997 1541
rect 4631 1527 4645 1541
rect 5423 1527 5437 1541
rect 23 1504 37 1518
rect 719 1504 733 1518
rect 1415 1504 1429 1518
rect 2255 1504 2269 1518
rect 3023 1504 3037 1518
rect 3863 1504 3877 1518
rect 4751 1504 4765 1518
rect 5399 1504 5413 1518
rect 479 1481 493 1495
rect 1199 1481 1213 1495
rect 2039 1481 2053 1495
rect 2927 1481 2941 1495
rect 3767 1481 3781 1495
rect 4439 1481 4453 1495
rect 5207 1481 5221 1495
rect 6143 1481 6157 1495
rect 455 1459 469 1473
rect 1175 1459 1189 1473
rect 2159 1459 2173 1473
rect 2831 1459 2845 1473
rect 3647 1459 3661 1473
rect 4535 1459 4549 1473
rect 5183 1459 5197 1473
rect 6023 1459 6037 1473
rect 431 1436 445 1450
rect 1319 1436 1333 1450
rect 2015 1436 2029 1450
rect 2807 1436 2821 1450
rect 3623 1436 3637 1450
rect 4415 1436 4429 1450
rect 5303 1436 5317 1450
rect 5999 1436 6013 1450
rect 335 1413 349 1427
rect 959 1413 973 1427
rect 1799 1413 1813 1427
rect 2711 1413 2725 1427
rect 3527 1413 3541 1427
rect 4223 1413 4237 1427
rect 4991 1413 5005 1427
rect 5903 1413 5917 1427
rect 311 1391 325 1405
rect 935 1391 949 1405
rect 1919 1391 1933 1405
rect 2615 1391 2629 1405
rect 3407 1391 3421 1405
rect 4319 1391 4333 1405
rect 4967 1391 4981 1405
rect 5783 1391 5797 1405
rect 287 1368 301 1382
rect 1079 1368 1093 1382
rect 1775 1368 1789 1382
rect 2591 1368 2605 1382
rect 3383 1368 3397 1382
rect 4199 1368 4213 1382
rect 5087 1368 5101 1382
rect 5759 1368 5773 1382
<< metal2 >>
rect 24 1518 36 1618
rect 48 1541 60 1618
rect 72 1563 84 1618
rect 122 1587 134 1618
rect 24 1339 36 1504
rect 48 1339 60 1527
rect 72 1339 84 1549
rect 192 1339 204 1572
rect 288 1382 300 1618
rect 312 1405 324 1618
rect 336 1427 348 1618
rect 432 1450 444 1618
rect 456 1473 468 1618
rect 480 1495 492 1618
rect 288 1339 300 1368
rect 312 1339 324 1391
rect 336 1339 348 1413
rect 432 1339 444 1436
rect 456 1339 468 1459
rect 480 1339 492 1481
rect 576 1339 588 1527
rect 600 1339 612 1549
rect 720 1339 732 1504
rect 840 1339 852 1572
rect 936 1339 948 1391
rect 960 1339 972 1413
rect 1080 1339 1092 1368
rect 1176 1339 1188 1459
rect 1200 1339 1212 1481
rect 1320 1339 1332 1436
rect 1416 1339 1428 1504
rect 1440 1339 1452 1549
rect 1560 1339 1572 1527
rect 1680 1339 1692 1572
rect 1776 1339 1788 1368
rect 1800 1339 1812 1413
rect 1920 1339 1932 1391
rect 2016 1339 2028 1436
rect 2040 1339 2052 1481
rect 2160 1339 2172 1459
rect 2256 1339 2268 1504
rect 2280 1339 2292 1527
rect 2376 1339 2388 1549
rect 2496 1339 2508 1572
rect 2592 1339 2604 1368
rect 2616 1339 2628 1391
rect 2712 1339 2724 1413
rect 2808 1339 2820 1436
rect 2832 1339 2844 1459
rect 2928 1339 2940 1481
rect 3024 1339 3036 1504
rect 3048 1339 3060 1527
rect 3168 1339 3180 1549
rect 3288 1339 3300 1572
rect 3384 1339 3396 1368
rect 3408 1339 3420 1391
rect 3528 1339 3540 1413
rect 3624 1339 3636 1436
rect 3648 1339 3660 1459
rect 3768 1339 3780 1481
rect 3864 1339 3876 1504
rect 3888 1339 3900 1549
rect 3984 1339 3996 1527
rect 4104 1339 4116 1572
rect 4200 1339 4212 1368
rect 4224 1339 4236 1413
rect 4320 1339 4332 1391
rect 4416 1339 4428 1436
rect 4440 1339 4452 1481
rect 4536 1339 4548 1459
rect 4632 1339 4644 1527
rect 4656 1339 4668 1549
rect 4752 1339 4764 1504
rect 4872 1339 4884 1572
rect 4968 1339 4980 1391
rect 4992 1339 5004 1413
rect 5088 1339 5100 1368
rect 5184 1339 5196 1459
rect 5208 1339 5220 1481
rect 5304 1339 5316 1436
rect 5400 1339 5412 1504
rect 5424 1339 5436 1527
rect 5544 1339 5556 1549
rect 5664 1339 5676 1572
rect 5760 1339 5772 1368
rect 5784 1339 5796 1391
rect 5904 1339 5916 1413
rect 6000 1339 6012 1436
rect 6024 1339 6036 1459
rect 6144 1339 6156 1481
rect 120 528 180 540
rect 240 383 252 540
rect 384 451 396 540
rect 528 473 540 540
rect 648 528 708 540
rect 768 528 828 540
rect 888 495 900 540
rect 1008 528 1068 540
rect 1128 517 1140 540
rect 1248 528 1308 540
rect 1128 505 1333 517
rect 888 483 1235 495
rect 528 461 1044 473
rect 384 439 828 451
rect 72 371 252 383
rect 72 0 84 371
rect 816 0 828 439
rect 1032 0 1044 461
rect 1223 0 1235 483
rect 1321 43 1333 505
rect 1368 70 1380 540
rect 1488 528 1548 540
rect 1608 528 1668 540
rect 1728 92 1740 541
rect 4080 540 4092 542
rect 4848 540 4860 542
rect 1848 528 1908 540
rect 1968 114 1980 540
rect 2088 528 2148 540
rect 2208 136 2220 540
rect 2304 528 2364 540
rect 2424 528 2484 540
rect 2544 158 2556 540
rect 2640 528 2700 540
rect 2760 180 2772 540
rect 2856 528 2916 540
rect 2976 202 2988 540
rect 3096 528 3156 540
rect 3216 528 3276 540
rect 3336 224 3348 540
rect 3456 528 3516 540
rect 3576 246 3588 540
rect 3696 528 3756 540
rect 3816 268 3828 540
rect 3912 528 3972 540
rect 4032 528 4092 540
rect 4152 290 4164 540
rect 4248 528 4308 540
rect 4368 312 4380 540
rect 4464 528 4524 540
rect 4584 334 4596 540
rect 4680 528 4740 540
rect 4800 528 4860 540
rect 4920 356 4932 540
rect 5016 528 5076 540
rect 5136 378 5148 540
rect 5232 528 5292 540
rect 5352 400 5364 540
rect 5472 528 5532 540
rect 5592 528 5652 540
rect 5712 422 5724 540
rect 5832 528 5892 540
rect 5952 444 5964 540
rect 6072 528 6132 540
rect 6192 466 6204 540
rect 6192 454 9108 466
rect 5952 432 8892 444
rect 5712 410 8148 422
rect 5352 388 7956 400
rect 5136 366 7740 378
rect 4920 344 6996 356
rect 4584 322 6804 334
rect 4368 300 6588 312
rect 4152 278 5844 290
rect 3816 256 5652 268
rect 3576 234 5436 246
rect 3336 212 4692 224
rect 2976 190 4501 202
rect 2760 168 4284 180
rect 2543 146 3540 158
rect 2208 124 3348 136
rect 1968 102 3132 114
rect 1728 80 2388 92
rect 1368 58 2196 70
rect 1321 31 1980 43
rect 1968 0 1980 31
rect 2184 0 2196 58
rect 2376 0 2388 80
rect 3120 0 3132 102
rect 3336 0 3348 124
rect 3528 0 3540 146
rect 4272 0 4284 168
rect 4489 0 4501 190
rect 4680 0 4692 212
rect 5424 0 5436 234
rect 5640 0 5652 256
rect 5832 0 5844 278
rect 6576 0 6588 300
rect 6792 0 6804 322
rect 6984 0 6996 344
rect 7728 0 7740 366
rect 7944 0 7956 388
rect 8136 0 8148 410
rect 8880 0 8892 432
rect 9096 0 9108 454
use nor3 nor3_2
timestamp 1386235396
transform 1 0 0 0 1 540
box 0 0 144 799
use and2 and2_10
timestamp 1386234845
transform 1 0 144 0 1 540
box 0 0 120 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 264 0 1 540
box 0 0 144 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 408 0 1 540
box 0 0 144 799
use nor2 nor2_12
timestamp 1386235306
transform 1 0 552 0 1 540
box 0 0 120 799
use and2 and2_11
timestamp 1386234845
transform 1 0 672 0 1 540
box 0 0 120 799
use and2 and2_12
timestamp 1386234845
transform 1 0 792 0 1 540
box 0 0 120 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 912 0 1 540
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 1032 0 1 540
box 0 0 120 799
use nor2 nor2_6
timestamp 1386235306
transform 1 0 1152 0 1 540
box 0 0 120 799
use and2 and2_5
timestamp 1386234845
transform 1 0 1272 0 1 540
box 0 0 120 799
use nor2 nor2_13
timestamp 1386235306
transform 1 0 1392 0 1 540
box 0 0 120 799
use and2 and2_13
timestamp 1386234845
transform 1 0 1512 0 1 540
box 0 0 120 799
use and2 and2_14
timestamp 1386234845
transform 1 0 1632 0 1 540
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 1752 0 1 540
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 1872 0 1 540
box 0 0 120 799
use nor2 nor2_7
timestamp 1386235306
transform 1 0 1992 0 1 540
box 0 0 120 799
use and2 and2_6
timestamp 1386234845
transform 1 0 2112 0 1 540
box 0 0 120 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 2232 0 1 540
box 0 0 96 799
use nor2 nor2_14
timestamp 1386235306
transform 1 0 2328 0 1 540
box 0 0 120 799
use and2 and2_15
timestamp 1386234845
transform 1 0 2448 0 1 540
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 2568 0 1 540
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 2664 0 1 540
box 0 0 120 799
use nand2 nand2_3
timestamp 1386234792
transform 1 0 2784 0 1 540
box 0 0 96 799
use nor2 nor2_8
timestamp 1386235306
transform 1 0 2880 0 1 540
box 0 0 120 799
use nor2 nor2_15
timestamp 1386235306
transform 1 0 3000 0 1 540
box 0 0 120 799
use and2 and2_16
timestamp 1386234845
transform 1 0 3120 0 1 540
box 0 0 120 799
use and2 and2_17
timestamp 1386234845
transform 1 0 3240 0 1 540
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 3360 0 1 540
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 3480 0 1 540
box 0 0 120 799
use nor2 nor2_9
timestamp 1386235306
transform 1 0 3600 0 1 540
box 0 0 120 799
use and2 and2_7
timestamp 1386234845
transform 1 0 3720 0 1 540
box 0 0 120 799
use nand2 nand2_7
timestamp 1386234792
transform 1 0 3840 0 1 540
box 0 0 96 799
use nor2 nor2_16
timestamp 1386235306
transform 1 0 3936 0 1 540
box 0 0 120 799
use and2 and2_18
timestamp 1386234845
transform 1 0 4056 0 1 540
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 4176 0 1 540
box 0 0 96 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 4272 0 1 540
box 0 0 120 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 4392 0 1 540
box 0 0 96 799
use nor2 nor2_10
timestamp 1386235306
transform 1 0 4488 0 1 540
box 0 0 120 799
use nand2 nand2_8
timestamp 1386234792
transform 1 0 4608 0 1 540
box 0 0 96 799
use nor2 nor2_17
timestamp 1386235306
transform 1 0 4704 0 1 540
box 0 0 120 799
use and2 and2_19
timestamp 1386234845
transform 1 0 4824 0 1 540
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 4944 0 1 540
box 0 0 96 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 5040 0 1 540
box 0 0 120 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 5160 0 1 540
box 0 0 96 799
use nor2 nor2_11
timestamp 1386235306
transform 1 0 5256 0 1 540
box 0 0 120 799
use and2 and2_20
timestamp 1386234845
transform 1 0 5376 0 1 540
box 0 0 120 799
use and2 and2_21
timestamp 1386234845
transform 1 0 5496 0 1 540
box 0 0 120 799
use and2 and2_22
timestamp 1386234845
transform 1 0 5616 0 1 540
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 5736 0 1 540
box 0 0 120 799
use and2 and2_4
timestamp 1386234845
transform 1 0 5856 0 1 540
box 0 0 120 799
use and2 and2_8
timestamp 1386234845
transform 1 0 5976 0 1 540
box 0 0 120 799
use and2 and2_9
timestamp 1386234845
transform 1 0 6096 0 1 540
box 0 0 120 799
<< labels >>
rlabel metal2 72 0 84 0 1 Rw[0]
rlabel metal2 816 0 828 0 1 Rs1[0]
rlabel metal2 1032 0 1044 0 1 Rs2[0]
rlabel metal2 1223 0 1235 0 1 Rw[1]
rlabel metal2 1968 0 1980 0 1 Rs1[1]
rlabel metal2 2184 0 2196 0 1 Rs2[1]
rlabel metal2 2376 0 2388 0 1 Rw[2]
rlabel metal2 3120 0 3132 0 1 Rs1[2]
rlabel metal2 3336 0 3348 0 1 Rs2[2]
rlabel metal2 3528 0 3540 0 1 Rw[3]
rlabel metal2 4272 0 4284 0 1 Rs1[3]
rlabel metal2 4489 0 4501 0 1 Rs2[3]
rlabel metal2 4680 0 4692 0 1 Rw[4]
rlabel metal2 5424 0 5436 0 1 Rs1[4]
rlabel metal2 5640 0 5652 0 1 Rs2[4]
rlabel metal2 5832 0 5844 0 1 Rw[5]
rlabel metal2 6576 0 6588 0 1 Rs1[5]
rlabel metal2 6792 0 6804 0 1 Rs2[5]
rlabel metal2 6984 0 6996 0 1 Rw[6]
rlabel metal2 7728 0 7740 0 1 Rs1[6]
rlabel metal2 7944 0 7956 0 1 Rs2[6]
rlabel metal2 8136 0 8148 0 1 Rw[7]
rlabel metal2 8880 0 8892 0 1 Rs1[7]
rlabel metal2 9096 0 9108 0 1 Rs2[7]
rlabel metal2 24 1618 36 1618 5 RwIn[0]
rlabel metal2 48 1618 60 1618 5 RwIn[1]
rlabel metal2 72 1618 84 1618 5 RwIn[2]
rlabel metal2 122 1618 134 1618 5 We
rlabel metal2 288 1618 300 1618 5 Rs1In[0]
rlabel metal2 312 1618 324 1618 5 Rs1In[1]
rlabel metal2 336 1618 348 1618 5 Rs1In[2]
rlabel metal2 432 1618 444 1618 5 Rs2In[0]
rlabel metal2 456 1618 468 1618 5 Rs2In[1]
rlabel metal2 480 1618 492 1618 5 Rs2In[2]
<< end >>
