magic
tech c035u
timestamp 1394313755
<< metal1 >>
rect -40 15949 51 15959
rect -40 15842 28 15852
rect -40 15819 28 15829
rect -40 15781 28 15806
rect -40 15136 28 15161
rect -40 15113 28 15123
rect -40 15090 28 15100
rect -40 15067 28 15077
rect 9209 14984 9273 14994
rect -40 14949 51 14959
rect 8993 14962 9273 14972
rect -40 14842 28 14852
rect -40 14819 28 14829
rect -40 14781 28 14806
rect -40 14136 28 14161
rect -40 14113 28 14123
rect -40 14090 28 14100
rect -40 14067 28 14077
rect 9209 13984 9273 13994
rect -40 13949 51 13959
rect 8993 13962 9273 13972
rect -40 13842 28 13852
rect -40 13819 28 13829
rect -40 13781 28 13806
rect -40 13136 28 13161
rect -40 13113 28 13123
rect -40 13090 28 13100
rect -40 13067 28 13077
rect 9209 12984 9273 12994
rect -40 12949 51 12959
rect 8993 12962 9273 12972
rect -40 12842 28 12852
rect -40 12819 28 12829
rect -40 12781 28 12806
rect -40 12136 28 12161
rect -40 12113 28 12123
rect -40 12090 28 12100
rect -40 12067 28 12077
rect 9209 11984 9273 11994
rect -40 11949 51 11959
rect 8993 11962 9273 11972
rect -40 11842 28 11852
rect -40 11819 28 11829
rect -40 11781 28 11806
rect -40 11136 28 11161
rect -40 11113 28 11123
rect -40 11090 28 11100
rect -40 11067 28 11077
rect 9209 10984 9273 10994
rect -40 10949 51 10959
rect 8993 10962 9273 10972
rect -40 10842 28 10852
rect -40 10819 28 10829
rect -40 10781 28 10806
rect -40 10136 28 10161
rect -40 10113 28 10123
rect -40 10090 28 10100
rect -40 10067 28 10077
rect 9209 9984 9273 9994
rect -40 9949 51 9959
rect 8993 9962 9273 9972
rect -40 9842 28 9852
rect -40 9819 28 9829
rect -40 9781 28 9806
rect -40 9136 28 9161
rect -40 9113 28 9123
rect -40 9090 28 9100
rect -40 9067 28 9077
rect 9209 8984 9273 8994
rect -40 8949 51 8959
rect 8993 8962 9273 8972
rect -40 8842 28 8852
rect -40 8819 28 8829
rect -40 8781 28 8806
rect -40 8136 28 8161
rect -40 8113 28 8123
rect -40 8090 28 8100
rect -40 8067 28 8077
rect 9209 7984 9273 7994
rect -40 7949 51 7959
rect 8993 7962 9273 7972
rect -40 7842 28 7852
rect -40 7819 28 7829
rect -40 7781 28 7806
rect -40 7136 28 7161
rect -40 7113 28 7123
rect -40 7090 28 7100
rect -40 7067 28 7077
rect 9209 6984 9273 6994
rect -40 6949 51 6959
rect 8993 6962 9273 6972
rect -40 6842 28 6852
rect -40 6819 28 6829
rect -40 6781 28 6806
rect -40 6136 28 6161
rect -40 6113 28 6123
rect -40 6090 28 6100
rect -40 6067 28 6077
rect 9209 5984 9273 5994
rect -40 5949 51 5959
rect 8993 5962 9273 5972
rect -40 5842 28 5852
rect -40 5819 28 5829
rect -40 5781 28 5806
rect -40 5136 28 5161
rect -40 5113 28 5123
rect -40 5090 28 5100
rect -40 5067 28 5077
rect 9209 4984 9273 4994
rect -40 4949 51 4959
rect 8993 4962 9273 4972
rect -40 4842 28 4852
rect -40 4819 28 4829
rect -40 4781 28 4806
rect -40 4136 28 4161
rect -40 4113 28 4123
rect -40 4090 28 4100
rect -40 4067 28 4077
rect 9209 3984 9273 3994
rect -40 3949 51 3959
rect 8993 3962 9273 3972
rect -40 3842 28 3852
rect -40 3819 28 3829
rect -40 3781 28 3806
rect -40 3136 28 3161
rect -40 3113 28 3123
rect -40 3090 28 3100
rect -40 3067 28 3077
rect 9209 2984 9273 2994
rect -40 2949 51 2959
rect 8993 2962 9273 2972
rect -40 2842 28 2852
rect -40 2819 28 2829
rect -40 2781 28 2806
rect -40 2136 28 2161
rect -40 2113 28 2123
rect -40 2090 28 2100
rect -40 2067 28 2077
rect 9209 1984 9273 1994
rect -40 1949 51 1959
rect 8993 1962 9273 1972
rect -40 1842 28 1852
rect -40 1819 28 1829
rect -40 1781 28 1806
rect -40 1136 28 1161
rect -40 1113 28 1123
rect -40 1090 28 1100
rect -40 1067 28 1077
rect 9209 984 9273 994
rect -40 949 51 959
rect 8993 962 9273 972
rect -40 842 28 852
rect -40 819 28 829
rect -40 781 28 806
rect -40 136 28 161
rect -40 113 28 123
rect -40 90 28 100
rect -40 67 28 77
rect 9209 -16 9273 -6
rect 8993 -38 9273 -28
<< m2contact >>
rect 51 15947 65 15961
rect 9195 14982 9209 14996
rect 51 14947 65 14961
rect 8979 14960 8993 14974
rect 9195 13982 9209 13996
rect 51 13947 65 13961
rect 8979 13960 8993 13974
rect 9195 12982 9209 12996
rect 51 12947 65 12961
rect 8979 12960 8993 12974
rect 9195 11982 9209 11996
rect 51 11947 65 11961
rect 8979 11960 8993 11974
rect 9195 10982 9209 10996
rect 51 10947 65 10961
rect 8979 10960 8993 10974
rect 9195 9982 9209 9996
rect 51 9947 65 9961
rect 8979 9960 8993 9974
rect 9195 8982 9209 8996
rect 51 8947 65 8961
rect 8979 8960 8993 8974
rect 9195 7982 9209 7996
rect 51 7947 65 7961
rect 8979 7960 8993 7974
rect 9195 6982 9209 6996
rect 51 6947 65 6961
rect 8979 6960 8993 6974
rect 9195 5982 9209 5996
rect 51 5947 65 5961
rect 8979 5960 8993 5974
rect 9195 4982 9209 4996
rect 51 4947 65 4961
rect 8979 4960 8993 4974
rect 9195 3982 9209 3996
rect 51 3947 65 3961
rect 8979 3960 8993 3974
rect 9195 2982 9209 2996
rect 51 2947 65 2961
rect 8979 2960 8993 2974
rect 9195 1982 9209 1996
rect 51 1947 65 1961
rect 8979 1960 8993 1974
rect 9195 982 9209 996
rect 51 947 65 961
rect 8979 960 8993 974
rect 9195 -18 9209 -4
rect 8979 -40 8993 -26
<< metal2 >>
rect 52 17588 64 17601
rect 76 17588 88 17601
rect 100 17588 112 17601
rect 150 17588 162 17601
rect 316 17588 328 17601
rect 340 17588 352 17601
rect 364 17588 376 17601
rect 460 17588 472 17601
rect 484 17588 496 17601
rect 508 17588 520 17601
rect 52 15939 64 15947
rect 100 15939 112 15970
rect 844 15939 856 15970
rect 1060 15939 1072 15970
rect 1252 15939 1264 15970
rect 1996 15939 2008 15970
rect 2212 15939 2224 15970
rect 2404 15939 2416 15970
rect 3148 15939 3160 15970
rect 3364 15939 3376 15970
rect 3556 15939 3568 15970
rect 4300 15939 4312 15970
rect 4516 15939 4528 15970
rect 4708 15939 4720 15970
rect 5452 15939 5464 15970
rect 5668 15939 5680 15970
rect 5860 15939 5872 15970
rect 6604 15939 6616 15970
rect 6820 15939 6832 15970
rect 7012 15939 7024 15970
rect 7756 15939 7768 15970
rect 7972 15939 7984 15970
rect 8164 15939 8176 15970
rect 8908 15939 8920 15970
rect 9124 15939 9136 15970
rect 52 14939 64 14947
rect 100 14939 112 15000
rect 844 14939 856 15000
rect 1060 14939 1072 15000
rect 1252 14939 1264 15000
rect 1996 14939 2008 15000
rect 2212 14939 2224 15000
rect 2404 14939 2416 15000
rect 3148 14939 3160 15000
rect 3364 14939 3376 15000
rect 3556 14939 3568 15000
rect 4300 14939 4312 15000
rect 4516 14939 4528 15000
rect 4708 14939 4720 15000
rect 5452 14939 5464 15000
rect 5668 14939 5680 15000
rect 5860 14939 5872 15000
rect 6604 14939 6616 15000
rect 6820 14939 6832 15000
rect 7012 14939 7024 15000
rect 7756 14939 7768 15000
rect 7972 14939 7984 15000
rect 8164 14939 8176 15000
rect 8908 14939 8920 15000
rect 8980 14974 8992 15000
rect 9124 14939 9136 15000
rect 9196 14996 9208 15000
rect 52 13939 64 13947
rect 100 13939 112 14000
rect 844 13939 856 14000
rect 1060 13939 1072 14000
rect 1252 13939 1264 14000
rect 1996 13939 2008 14000
rect 2212 13939 2224 14000
rect 2404 13939 2416 14000
rect 3148 13939 3160 14000
rect 3364 13939 3376 14000
rect 3556 13939 3568 14000
rect 4300 13939 4312 14000
rect 4516 13939 4528 14000
rect 4708 13939 4720 14000
rect 5452 13939 5464 14000
rect 5668 13939 5680 14000
rect 5860 13939 5872 14000
rect 6604 13939 6616 14000
rect 6820 13939 6832 14000
rect 7012 13939 7024 14000
rect 7756 13939 7768 14000
rect 7972 13939 7984 14000
rect 8164 13939 8176 14000
rect 8908 13939 8920 14000
rect 8980 13974 8992 14000
rect 9124 13939 9136 14000
rect 9196 13996 9208 14000
rect 52 12939 64 12947
rect 100 12939 112 13000
rect 844 12939 856 13000
rect 1060 12939 1072 13000
rect 1252 12939 1264 13000
rect 1996 12939 2008 13000
rect 2212 12939 2224 13000
rect 2404 12939 2416 13000
rect 3148 12939 3160 13000
rect 3364 12939 3376 13000
rect 3556 12939 3568 13000
rect 4300 12939 4312 13000
rect 4516 12939 4528 13000
rect 4708 12939 4720 13000
rect 5452 12939 5464 13000
rect 5668 12939 5680 13000
rect 5860 12939 5872 13000
rect 6604 12939 6616 13000
rect 6820 12939 6832 13000
rect 7012 12939 7024 13000
rect 7756 12939 7768 13000
rect 7972 12939 7984 13000
rect 8164 12939 8176 13000
rect 8908 12939 8920 13000
rect 8980 12974 8992 13000
rect 9124 12939 9136 13000
rect 9196 12996 9208 13000
rect 52 11939 64 11947
rect 100 11939 112 12000
rect 844 11939 856 12000
rect 1060 11939 1072 12000
rect 1252 11939 1264 12000
rect 1996 11939 2008 12000
rect 2212 11939 2224 12000
rect 2404 11939 2416 12000
rect 3148 11939 3160 12000
rect 3364 11939 3376 12000
rect 3556 11939 3568 12000
rect 4300 11939 4312 12000
rect 4516 11939 4528 12000
rect 4708 11939 4720 12000
rect 5452 11939 5464 12000
rect 5668 11939 5680 12000
rect 5860 11939 5872 12000
rect 6604 11939 6616 12000
rect 6820 11939 6832 12000
rect 7012 11939 7024 12000
rect 7756 11939 7768 12000
rect 7972 11939 7984 12000
rect 8164 11939 8176 12000
rect 8908 11939 8920 12000
rect 8980 11974 8992 12000
rect 9124 11939 9136 12000
rect 9196 11996 9208 12000
rect 52 10939 64 10947
rect 100 10939 112 11000
rect 844 10939 856 11000
rect 1060 10939 1072 11000
rect 1252 10939 1264 11000
rect 1996 10939 2008 11000
rect 2212 10939 2224 11000
rect 2404 10939 2416 11000
rect 3148 10939 3160 11000
rect 3364 10939 3376 11000
rect 3556 10939 3568 11000
rect 4300 10939 4312 11000
rect 4516 10939 4528 11000
rect 4708 10939 4720 11000
rect 5452 10939 5464 11000
rect 5668 10939 5680 11000
rect 5860 10939 5872 11000
rect 6604 10939 6616 11000
rect 6820 10939 6832 11000
rect 7012 10939 7024 11000
rect 7756 10939 7768 11000
rect 7972 10939 7984 11000
rect 8164 10939 8176 11000
rect 8908 10939 8920 11000
rect 8980 10974 8992 11000
rect 9124 10939 9136 11000
rect 9196 10996 9208 11000
rect 52 9939 64 9947
rect 100 9939 112 10000
rect 844 9939 856 10000
rect 1060 9939 1072 10000
rect 1252 9939 1264 10000
rect 1996 9939 2008 10000
rect 2212 9939 2224 10000
rect 2404 9939 2416 10000
rect 3148 9939 3160 10000
rect 3364 9939 3376 10000
rect 3556 9939 3568 10000
rect 4300 9939 4312 10000
rect 4516 9939 4528 10000
rect 4708 9939 4720 10000
rect 5452 9939 5464 10000
rect 5668 9939 5680 10000
rect 5860 9939 5872 10000
rect 6604 9939 6616 10000
rect 6820 9939 6832 10000
rect 7012 9939 7024 10000
rect 7756 9939 7768 10000
rect 7972 9939 7984 10000
rect 8164 9939 8176 10000
rect 8908 9939 8920 10000
rect 8980 9974 8992 10000
rect 9124 9939 9136 10000
rect 9196 9996 9208 10000
rect 52 8939 64 8947
rect 100 8939 112 9000
rect 844 8939 856 9000
rect 1060 8939 1072 9000
rect 1252 8939 1264 9000
rect 1996 8939 2008 9000
rect 2212 8939 2224 9000
rect 2404 8939 2416 9000
rect 3148 8939 3160 9000
rect 3364 8939 3376 9000
rect 3556 8939 3568 9000
rect 4300 8939 4312 9000
rect 4516 8939 4528 9000
rect 4708 8939 4720 9000
rect 5452 8939 5464 9000
rect 5668 8939 5680 9000
rect 5860 8939 5872 9000
rect 6604 8939 6616 9000
rect 6820 8939 6832 9000
rect 7012 8939 7024 9000
rect 7756 8939 7768 9000
rect 7972 8939 7984 9000
rect 8164 8939 8176 9000
rect 8908 8939 8920 9000
rect 8980 8974 8992 9000
rect 9124 8939 9136 9000
rect 9196 8996 9208 9000
rect 52 7939 64 7947
rect 100 7939 112 8000
rect 844 7939 856 8000
rect 1060 7939 1072 8000
rect 1252 7939 1264 8000
rect 1996 7939 2008 8000
rect 2212 7939 2224 8000
rect 2404 7939 2416 8000
rect 3148 7939 3160 8000
rect 3364 7939 3376 8000
rect 3556 7939 3568 8000
rect 4300 7939 4312 8000
rect 4516 7939 4528 8000
rect 4708 7939 4720 8000
rect 5452 7939 5464 8000
rect 5668 7939 5680 8000
rect 5860 7939 5872 8000
rect 6604 7939 6616 8000
rect 6820 7939 6832 8000
rect 7012 7939 7024 8000
rect 7756 7939 7768 8000
rect 7972 7939 7984 8000
rect 8164 7939 8176 8000
rect 8908 7939 8920 8000
rect 8980 7974 8992 8000
rect 9124 7939 9136 8000
rect 9196 7996 9208 8000
rect 52 6939 64 6947
rect 100 6939 112 7000
rect 844 6939 856 7000
rect 1060 6939 1072 7000
rect 1252 6939 1264 7000
rect 1996 6939 2008 7000
rect 2212 6939 2224 7000
rect 2404 6939 2416 7000
rect 3148 6939 3160 7000
rect 3364 6939 3376 7000
rect 3556 6939 3568 7000
rect 4300 6939 4312 7000
rect 4516 6939 4528 7000
rect 4708 6939 4720 7000
rect 5452 6939 5464 7000
rect 5668 6939 5680 7000
rect 5860 6939 5872 7000
rect 6604 6939 6616 7000
rect 6820 6939 6832 7000
rect 7012 6939 7024 7000
rect 7756 6939 7768 7000
rect 7972 6939 7984 7000
rect 8164 6939 8176 7000
rect 8908 6939 8920 7000
rect 8980 6974 8992 7000
rect 9124 6939 9136 7000
rect 9196 6996 9208 7000
rect 52 5939 64 5947
rect 100 5939 112 6000
rect 844 5939 856 6000
rect 1060 5939 1072 6000
rect 1252 5939 1264 6000
rect 1996 5939 2008 6000
rect 2212 5939 2224 6000
rect 2404 5939 2416 6000
rect 3148 5939 3160 6000
rect 3364 5939 3376 6000
rect 3556 5939 3568 6000
rect 4300 5939 4312 6000
rect 4516 5939 4528 6000
rect 4708 5939 4720 6000
rect 5452 5939 5464 6000
rect 5668 5939 5680 6000
rect 5860 5939 5872 6000
rect 6604 5939 6616 6000
rect 6820 5939 6832 6000
rect 7012 5939 7024 6000
rect 7756 5939 7768 6000
rect 7972 5939 7984 6000
rect 8164 5939 8176 6000
rect 8908 5939 8920 6000
rect 8980 5974 8992 6000
rect 9124 5939 9136 6000
rect 9196 5996 9208 6000
rect 52 4939 64 4947
rect 100 4939 112 5000
rect 844 4939 856 5000
rect 1060 4939 1072 5000
rect 1252 4939 1264 5000
rect 1996 4939 2008 5000
rect 2212 4939 2224 5000
rect 2404 4939 2416 5000
rect 3148 4939 3160 5000
rect 3364 4939 3376 5000
rect 3556 4939 3568 5000
rect 4300 4939 4312 5000
rect 4516 4939 4528 5000
rect 4708 4939 4720 5000
rect 5452 4939 5464 5000
rect 5668 4939 5680 5000
rect 5860 4939 5872 5000
rect 6604 4939 6616 5000
rect 6820 4939 6832 5000
rect 7012 4939 7024 5000
rect 7756 4939 7768 5000
rect 7972 4939 7984 5000
rect 8164 4939 8176 5000
rect 8908 4939 8920 5000
rect 8980 4974 8992 5000
rect 9124 4939 9136 5000
rect 9196 4996 9208 5000
rect 52 3939 64 3947
rect 100 3939 112 4000
rect 844 3939 856 4000
rect 1060 3939 1072 4000
rect 1252 3939 1264 4000
rect 1996 3939 2008 4000
rect 2212 3939 2224 4000
rect 2404 3939 2416 4000
rect 3148 3939 3160 4000
rect 3364 3939 3376 4000
rect 3556 3939 3568 4000
rect 4300 3939 4312 4000
rect 4516 3939 4528 4000
rect 4708 3939 4720 4000
rect 5452 3939 5464 4000
rect 5668 3939 5680 4000
rect 5860 3939 5872 4000
rect 6604 3939 6616 4000
rect 6820 3939 6832 4000
rect 7012 3939 7024 4000
rect 7756 3939 7768 4000
rect 7972 3939 7984 4000
rect 8164 3939 8176 4000
rect 8908 3939 8920 4000
rect 8980 3974 8992 4000
rect 9124 3939 9136 4000
rect 9196 3996 9208 4000
rect 52 2939 64 2947
rect 100 2939 112 3000
rect 844 2939 856 3000
rect 1060 2939 1072 3000
rect 1252 2939 1264 3000
rect 1996 2939 2008 3000
rect 2212 2939 2224 3000
rect 2404 2939 2416 3000
rect 3148 2939 3160 3000
rect 3364 2939 3376 3000
rect 3556 2939 3568 3000
rect 4300 2939 4312 3000
rect 4516 2939 4528 3000
rect 4708 2939 4720 3000
rect 5452 2939 5464 3000
rect 5668 2939 5680 3000
rect 5860 2939 5872 3000
rect 6604 2939 6616 3000
rect 6820 2939 6832 3000
rect 7012 2939 7024 3000
rect 7756 2939 7768 3000
rect 7972 2939 7984 3000
rect 8164 2939 8176 3000
rect 8908 2939 8920 3000
rect 8980 2974 8992 3000
rect 9124 2939 9136 3000
rect 9196 2996 9208 3000
rect 52 1939 64 1947
rect 100 1939 112 2000
rect 844 1939 856 2000
rect 1060 1939 1072 2000
rect 1252 1939 1264 2000
rect 1996 1939 2008 2000
rect 2212 1939 2224 2000
rect 2404 1939 2416 2000
rect 3148 1939 3160 2000
rect 3364 1939 3376 2000
rect 3556 1939 3568 2000
rect 4300 1939 4312 2000
rect 4516 1939 4528 2000
rect 4708 1939 4720 2000
rect 5452 1939 5464 2000
rect 5668 1939 5680 2000
rect 5860 1939 5872 2000
rect 6604 1939 6616 2000
rect 6820 1939 6832 2000
rect 7012 1939 7024 2000
rect 7756 1939 7768 2000
rect 7972 1939 7984 2000
rect 8164 1939 8176 2000
rect 8908 1939 8920 2000
rect 8980 1974 8992 2000
rect 9124 1939 9136 2000
rect 9196 1996 9208 2000
rect 52 939 64 947
rect 100 939 112 1000
rect 844 939 856 1000
rect 1060 939 1072 1000
rect 1252 939 1264 1000
rect 1996 939 2008 1000
rect 2212 939 2224 1000
rect 2404 939 2416 1000
rect 3148 939 3160 1000
rect 3364 939 3376 1000
rect 3556 939 3568 1000
rect 4300 939 4312 1000
rect 4516 939 4528 1000
rect 4708 939 4720 1000
rect 5452 939 5464 1000
rect 5668 939 5680 1000
rect 5860 939 5872 1000
rect 6604 939 6616 1000
rect 6820 939 6832 1000
rect 7012 939 7024 1000
rect 7756 939 7768 1000
rect 7972 939 7984 1000
rect 8164 939 8176 1000
rect 8908 939 8920 1000
rect 8980 974 8992 1000
rect 9124 939 9136 1000
rect 9196 996 9208 1000
rect 100 -61 112 0
rect 844 -61 856 0
rect 1060 -61 1072 0
rect 1252 -61 1264 0
rect 1996 -61 2008 0
rect 2212 -61 2224 0
rect 2404 -61 2416 0
rect 3148 -61 3160 0
rect 3364 -61 3376 0
rect 3556 -61 3568 0
rect 4300 -61 4312 0
rect 4516 -61 4528 0
rect 4708 -61 4720 0
rect 5452 -61 5464 0
rect 5668 -61 5680 0
rect 5860 -61 5872 0
rect 6604 -61 6616 0
rect 6820 -61 6832 0
rect 7012 -61 7024 0
rect 7756 -61 7768 0
rect 7972 -61 7984 0
rect 8164 -61 8176 0
rect 8908 -61 8920 0
rect 8980 -26 8992 0
rect 9124 -61 9136 0
rect 9196 -4 9208 0
use regBlock_decoder  regBlock_decoder_0
timestamp 1394304361
transform 1 0 28 0 1 15970
box 0 0 9216 1618
use regBlock_slice  regBlock_slice_0
array 0 0 9313 0 15 1000
timestamp 1394295027
transform 1 0 28 0 1 0
box 0 0 9216 939
<< labels >>
rlabel metal1 9273 -16 9273 -6 7 Rd2[0]
rlabel metal1 9273 984 9273 994 7 Rd2[1]
rlabel metal1 9273 1984 9273 1994 7 Rd2[2]
rlabel metal1 9273 2984 9273 2994 7 Rd2[3]
rlabel metal1 9273 3984 9273 3994 7 Rd2[4]
rlabel metal1 9273 4984 9273 4994 7 Rd2[5]
rlabel metal1 9273 5984 9273 5994 7 Rd2[6]
rlabel metal1 9273 6984 9273 6994 7 Rd2[7]
rlabel metal1 9273 7984 9273 7994 7 Rd2[8]
rlabel metal1 9273 8984 9273 8994 7 Rd2[9]
rlabel metal1 9273 9984 9273 9994 7 Rd2[10]
rlabel metal1 9273 10984 9273 10994 7 Rd2[11]
rlabel metal1 9273 11984 9273 11994 7 Rd2[12]
rlabel metal1 9273 12984 9273 12994 7 Rd2[13]
rlabel metal1 9273 13984 9273 13994 7 Rd2[14]
rlabel metal1 9273 14984 9273 14994 7 Rd2[15]
rlabel metal1 9273 -38 9273 -28 7 Rd1[0]
rlabel metal1 9273 962 9273 972 7 Rd1[1]
rlabel metal1 9273 1962 9273 1972 7 Rd1[2]
rlabel metal1 9273 2962 9273 2972 7 Rd1[3]
rlabel metal1 9273 3962 9273 3972 7 Rd1[4]
rlabel metal1 9273 4962 9273 4972 7 Rd1[5]
rlabel metal1 9273 5962 9273 5972 7 Rd1[6]
rlabel metal1 9273 6962 9273 6972 7 Rd1[7]
rlabel metal1 9273 7962 9273 7972 7 Rd1[8]
rlabel metal1 9273 8962 9273 8972 7 Rd1[9]
rlabel metal1 9273 9962 9273 9972 7 Rd1[10]
rlabel metal1 9273 10962 9273 10972 7 Rd1[11]
rlabel metal1 9273 11962 9273 11972 7 Rd1[12]
rlabel metal1 9273 12962 9273 12972 7 Rd1[13]
rlabel metal1 9273 13962 9273 13972 7 Rd1[14]
rlabel metal1 9273 14962 9273 14972 7 Rd1[15]
rlabel metal1 -40 67 -40 77 3 nReset
rlabel metal1 -40 1067 -40 1077 3 nReset
rlabel metal1 -40 2067 -40 2077 3 nReset
rlabel metal1 -40 3067 -40 3077 3 nReset
rlabel metal1 -40 4067 -40 4077 3 nReset
rlabel metal1 -40 5067 -40 5077 3 nReset
rlabel metal1 -40 6067 -40 6077 3 nReset
rlabel metal1 -40 7067 -40 7077 3 nReset
rlabel metal1 -40 8067 -40 8077 3 nReset
rlabel metal1 -40 9067 -40 9077 3 nReset
rlabel metal1 -40 10067 -40 10077 3 nReset
rlabel metal1 -40 11067 -40 11077 3 nReset
rlabel metal1 -40 12067 -40 12077 3 nReset
rlabel metal1 -40 13067 -40 13077 3 nReset
rlabel metal1 -40 14067 -40 14077 3 nReset
rlabel metal1 -40 15067 -40 15077 3 nReset
rlabel metal1 -40 90 -40 100 3 Test
rlabel metal1 -40 1090 -40 1100 3 Test
rlabel metal1 -40 2090 -40 2100 3 Test
rlabel metal1 -40 3090 -40 3100 3 Test
rlabel metal1 -40 4090 -40 4100 3 Test
rlabel metal1 -40 5090 -40 5100 3 Test
rlabel metal1 -40 6090 -40 6100 3 Test
rlabel metal1 -40 7090 -40 7100 3 Test
rlabel metal1 -40 8090 -40 8100 3 Test
rlabel metal1 -40 9090 -40 9100 3 Test
rlabel metal1 -40 10090 -40 10100 3 Test
rlabel metal1 -40 11090 -40 11100 3 Test
rlabel metal1 -40 12090 -40 12100 3 Test
rlabel metal1 -40 13090 -40 13100 3 Test
rlabel metal1 -40 14090 -40 14100 3 Test
rlabel metal1 -40 15090 -40 15100 3 Test
rlabel metal1 -40 113 -40 123 3 Clock
rlabel metal1 -40 1113 -40 1123 3 Clock
rlabel metal1 -40 2113 -40 2123 3 Clock
rlabel metal1 -40 3113 -40 3123 3 Clock
rlabel metal1 -40 4113 -40 4123 3 Clock
rlabel metal1 -40 5113 -40 5123 3 Clock
rlabel metal1 -40 6113 -40 6123 3 Clock
rlabel metal1 -40 7113 -40 7123 3 Clock
rlabel metal1 -40 8113 -40 8123 3 Clock
rlabel metal1 -40 9113 -40 9123 3 Clock
rlabel metal1 -40 10113 -40 10123 3 Clock
rlabel metal1 -40 11113 -40 11123 3 Clock
rlabel metal1 -40 12113 -40 12123 3 Clock
rlabel metal1 -40 13113 -40 13123 3 Clock
rlabel metal1 -40 14113 -40 14123 3 Clock
rlabel metal1 -40 15113 -40 15123 3 Clock
rlabel metal1 -40 136 -40 161 3 GND!
rlabel metal1 -40 1136 -40 1161 3 GND!
rlabel metal1 -40 2136 -40 2161 3 GND!
rlabel metal1 -40 3136 -40 3161 3 GND!
rlabel metal1 -40 4136 -40 4161 3 GND!
rlabel metal1 -40 5136 -40 5161 3 GND!
rlabel metal1 -40 6136 -40 6161 3 GND!
rlabel metal1 -40 7136 -40 7161 3 GND!
rlabel metal1 -40 8136 -40 8161 3 GND!
rlabel metal1 -40 9136 -40 9161 3 GND!
rlabel metal1 -40 10136 -40 10161 3 GND!
rlabel metal1 -40 11136 -40 11161 3 GND!
rlabel metal1 -40 12136 -40 12161 3 GND!
rlabel metal1 -40 13136 -40 13161 3 GND!
rlabel metal1 -40 14136 -40 14161 3 GND!
rlabel metal1 -40 15136 -40 15161 3 GND!
rlabel metal1 -40 781 -40 806 3 Vdd!
rlabel metal1 -40 1781 -40 1806 3 Vdd!
rlabel metal1 -40 2781 -40 2806 3 Vdd!
rlabel metal1 -40 3781 -40 3806 3 Vdd!
rlabel metal1 -40 4781 -40 4806 3 Vdd!
rlabel metal1 -40 5781 -40 5806 3 Vdd!
rlabel metal1 -40 6781 -40 6806 3 Vdd!
rlabel metal1 -40 7781 -40 7806 3 Vdd!
rlabel metal1 -40 8781 -40 8806 3 Vdd!
rlabel metal1 -40 9781 -40 9806 3 Vdd!
rlabel metal1 -40 10781 -40 10806 3 Vdd!
rlabel metal1 -40 11781 -40 11806 3 Vdd!
rlabel metal1 -40 12781 -40 12806 3 Vdd!
rlabel metal1 -40 13781 -40 13806 3 Vdd!
rlabel metal1 -40 14781 -40 14806 3 Vdd!
rlabel metal1 -40 15781 -40 15806 3 Vdd!
rlabel metal1 -40 819 -40 829 3 SDI
rlabel metal1 -40 1819 -40 1829 3 SDI
rlabel metal1 -40 2819 -40 2829 3 SDI
rlabel metal1 -40 3819 -40 3829 3 SDI
rlabel metal1 -40 4819 -40 4829 3 SDI
rlabel metal1 -40 5819 -40 5829 3 SDI
rlabel metal1 -40 6819 -40 6829 3 SDI
rlabel metal1 -40 7819 -40 7829 3 SDI
rlabel metal1 -40 8819 -40 8829 3 SDI
rlabel metal1 -40 9819 -40 9829 3 SDI
rlabel metal1 -40 10819 -40 10829 3 SDI
rlabel metal1 -40 11819 -40 11829 3 SDI
rlabel metal1 -40 12819 -40 12829 3 SDI
rlabel metal1 -40 13819 -40 13829 3 SDI
rlabel metal1 -40 14819 -40 14829 3 SDI
rlabel metal1 -40 15819 -40 15829 3 SDI
rlabel metal1 -40 842 -40 852 3 ScanReturn
rlabel metal1 -40 1842 -40 1852 3 ScanReturn
rlabel metal1 -40 2842 -40 2852 3 ScanReturn
rlabel metal1 -40 3842 -40 3852 3 ScanReturn
rlabel metal1 -40 4842 -40 4852 3 ScanReturn
rlabel metal1 -40 5842 -40 5852 3 ScanReturn
rlabel metal1 -40 6842 -40 6852 3 ScanReturn
rlabel metal1 -40 7842 -40 7852 3 ScanReturn
rlabel metal1 -40 8842 -40 8852 3 ScanReturn
rlabel metal1 -40 9842 -40 9852 3 ScanReturn
rlabel metal1 -40 10842 -40 10852 3 ScanReturn
rlabel metal1 -40 11842 -40 11852 3 ScanReturn
rlabel metal1 -40 12842 -40 12852 3 ScanReturn
rlabel metal1 -40 13842 -40 13852 3 ScanReturn
rlabel metal1 -40 14842 -40 14852 3 ScanReturn
rlabel metal1 -40 15842 -40 15852 3 ScanReturn
rlabel metal1 -40 949 -40 959 3 WData[0]
rlabel metal1 -40 1949 -40 1959 3 WData[1]
rlabel metal1 -40 2949 -40 2959 3 WData[2]
rlabel metal1 -40 3949 -40 3959 3 WData[3]
rlabel metal1 -40 4949 -40 4959 3 WData[4]
rlabel metal1 -40 5949 -40 5959 3 WData[5]
rlabel metal1 -40 6949 -40 6959 3 WData[6]
rlabel metal1 -40 7949 -40 7959 3 WData[7]
rlabel metal1 -40 8949 -40 8959 3 WData[8]
rlabel metal1 -40 9949 -40 9959 3 WData[9]
rlabel metal1 -40 10949 -40 10959 3 WData[10]
rlabel metal1 -40 11949 -40 11959 3 WData[11]
rlabel metal1 -40 12949 -40 12959 3 WData[12]
rlabel metal1 -40 13949 -40 13959 3 WData[13]
rlabel metal1 -40 14949 -40 14959 3 WData[14]
rlabel metal1 -40 15949 -40 15959 3 WData[15]
rlabel metal2 316 17601 328 17601 5 Rs1[0]
rlabel metal2 340 17601 352 17601 5 Rs1[1]
rlabel metal2 364 17601 376 17601 5 Rs1[2]
rlabel metal2 460 17601 472 17601 5 Rs2[0]
rlabel metal2 484 17601 496 17601 5 Rs2[1]
rlabel metal2 508 17601 520 17601 5 Rs2[2]
rlabel metal2 52 17601 64 17601 5 Rw[0]
rlabel metal2 76 17601 88 17601 5 Rw[1]
rlabel metal2 100 17601 112 17601 5 Rw[2]
rlabel metal2 150 17601 162 17601 5 RegWe
<< end >>
