../../../Design/Implementation/verilog/behavioural/io_leds.sv