magic
tech c035u
timestamp 1394493540
<< nwell >>
rect 0 798 168 1196
<< pwell >>
rect 0 397 168 798
<< pohmic >>
rect 0 473 6 483
rect 162 473 168 483
<< nohmic >>
rect 0 1133 6 1143
rect 162 1133 168 1143
<< psubstratetap >>
rect 6 473 162 489
<< nsubstratetap >>
rect 6 1127 162 1143
<< metal1 >>
rect 3709 1464 4751 1474
rect 3589 1442 4655 1452
rect 3349 1420 4463 1430
rect 3109 1399 4271 1409
rect 2989 1377 4175 1387
rect 877 1355 1271 1365
rect 3829 1355 4079 1365
rect 4093 1355 4847 1365
rect 997 1333 1247 1343
rect 1333 1333 1488 1343
rect 1549 1333 1607 1343
rect 3469 1333 3983 1343
rect 3997 1333 4559 1343
rect 1093 1311 1128 1321
rect 1213 1311 1367 1321
rect 1453 1311 1583 1321
rect 1933 1311 1967 1321
rect 2197 1311 2471 1321
rect 3229 1311 3887 1321
rect 3901 1311 4367 1321
rect 4597 1311 6407 1321
rect 685 1289 839 1299
rect 853 1289 1031 1299
rect 1045 1289 3071 1299
rect 3085 1289 3311 1299
rect 3325 1289 3551 1299
rect 3565 1289 3791 1299
rect 3805 1289 4967 1299
rect 4981 1289 5303 1299
rect 565 1267 1511 1277
rect 1525 1267 3167 1277
rect 3181 1267 3287 1277
rect 3301 1267 3647 1277
rect 3661 1267 3767 1277
rect 3781 1267 4943 1277
rect 4957 1267 5183 1277
rect 5197 1267 5279 1277
rect 5293 1267 5927 1277
rect 5941 1267 6911 1277
rect 445 1245 815 1255
rect 829 1245 1151 1255
rect 1165 1245 1727 1255
rect 1741 1245 3383 1255
rect 3397 1245 3503 1255
rect 3517 1245 3623 1255
rect 3637 1245 3743 1255
rect 3757 1245 6887 1255
rect 7117 1245 7223 1255
rect 325 1223 959 1233
rect 973 1223 1391 1233
rect 1405 1223 2831 1233
rect 2845 1223 4919 1233
rect 5005 1223 5038 1233
rect 5365 1223 5423 1233
rect 5869 1223 6047 1233
rect 6109 1223 6143 1233
rect 6253 1223 6287 1233
rect 6301 1223 6503 1233
rect 6517 1223 6623 1233
rect 6637 1223 6743 1233
rect 6973 1223 7199 1233
rect 205 1201 1703 1211
rect 1717 1201 2711 1211
rect 2725 1201 2807 1211
rect 2821 1201 5063 1211
rect 5245 1201 5399 1211
rect 5485 1201 5519 1211
rect 5989 1201 6023 1211
rect 6037 1201 7247 1211
rect 7309 1201 7343 1211
rect 0 1179 168 1189
rect 0 1156 168 1166
rect 0 1127 6 1143
rect 162 1127 168 1143
rect 0 1118 168 1127
rect 0 489 168 498
rect 0 473 6 489
rect 162 473 168 489
rect 0 450 168 460
rect 0 427 168 437
rect 0 404 168 414
rect 253 382 791 392
rect 805 382 1415 392
rect 1429 382 5543 392
rect 5557 382 6167 392
rect 6181 382 7367 392
rect 373 360 2735 370
rect 2749 360 5159 370
rect 5173 360 6191 370
rect 6205 360 6863 370
rect 6877 360 7007 370
rect 7117 360 7151 370
rect 493 338 935 348
rect 949 338 1055 348
rect 1069 338 1751 348
rect 1765 338 2903 348
rect 2917 338 3023 348
rect 3037 338 3143 348
rect 3157 338 3263 348
rect 3277 338 5567 348
rect 5581 338 5783 348
rect 5797 338 5903 348
rect 5917 338 7031 348
rect 613 316 2927 326
rect 2941 316 3047 326
rect 3061 316 3407 326
rect 3421 316 3527 326
rect 4165 316 4247 326
rect 4261 316 4343 326
rect 4357 316 4439 326
rect 4453 316 4535 326
rect 4549 316 4631 326
rect 4645 316 4727 326
rect 4741 316 4823 326
rect 5150 316 5615 326
rect 6349 316 6383 326
rect 733 294 911 304
rect 925 294 2951 304
rect 2965 294 3191 304
rect 3205 294 3431 304
rect 3445 294 3671 304
rect 3685 294 5807 304
rect 5821 294 7055 304
rect 349 272 1655 282
rect 1669 272 1991 282
rect 2005 272 2351 282
rect 2869 271 3863 281
rect 3877 271 3959 281
rect 3973 271 4055 281
rect 5793 272 6455 282
rect 1813 250 1871 260
rect 2773 249 4151 259
rect 4353 250 4487 260
rect 5581 250 6575 260
rect 85 227 3911 237
rect 4021 227 5687 237
rect 5989 228 6695 238
rect 517 205 2087 215
rect 2245 205 4339 215
rect 4693 205 6863 215
rect 6877 205 6883 215
rect 685 183 2159 193
rect 2893 183 4775 193
rect 6349 183 6815 193
rect 709 161 2375 171
rect 3229 161 4871 171
rect 6709 161 7415 171
rect 781 139 2543 149
rect 3349 139 5663 149
rect 997 117 2591 127
rect 3397 117 4583 127
rect 1141 95 5111 105
rect 1477 73 4199 83
rect 5125 71 5779 81
rect 1837 51 4295 61
rect 2581 29 4391 39
rect 3565 7 4103 17
<< m2contact >>
rect 3695 1462 3709 1476
rect 4751 1462 4765 1476
rect 3575 1440 3589 1454
rect 4655 1440 4669 1454
rect 3335 1419 3349 1433
rect 4463 1418 4477 1432
rect 3095 1397 3109 1411
rect 4271 1396 4285 1410
rect 2975 1375 2989 1389
rect 4175 1375 4189 1389
rect 863 1353 877 1367
rect 1271 1353 1285 1367
rect 3815 1353 3829 1367
rect 4079 1353 4093 1367
rect 4847 1353 4861 1367
rect 983 1331 997 1345
rect 1247 1331 1261 1345
rect 1319 1331 1333 1345
rect 1488 1331 1502 1345
rect 1535 1331 1549 1345
rect 1607 1331 1621 1345
rect 3455 1331 3469 1345
rect 3983 1331 3997 1345
rect 4559 1331 4573 1345
rect 1079 1309 1093 1323
rect 1128 1309 1142 1323
rect 1199 1309 1213 1323
rect 1367 1309 1381 1323
rect 1439 1309 1453 1323
rect 1583 1309 1597 1323
rect 1919 1309 1933 1323
rect 1967 1309 1981 1323
rect 2183 1309 2197 1323
rect 2471 1309 2485 1323
rect 3215 1309 3229 1323
rect 3887 1309 3901 1323
rect 4367 1309 4381 1323
rect 4583 1309 4597 1323
rect 6407 1309 6421 1323
rect 671 1287 685 1301
rect 839 1287 853 1301
rect 1031 1287 1045 1301
rect 3071 1287 3085 1301
rect 3311 1287 3325 1301
rect 3551 1287 3565 1301
rect 3791 1287 3805 1301
rect 4967 1287 4981 1301
rect 5303 1287 5317 1301
rect 551 1265 565 1279
rect 1511 1265 1525 1279
rect 3167 1265 3181 1279
rect 3287 1265 3301 1279
rect 3647 1265 3661 1279
rect 3767 1265 3781 1279
rect 4943 1265 4957 1279
rect 5183 1265 5197 1279
rect 5279 1265 5293 1279
rect 5927 1265 5941 1279
rect 6911 1265 6925 1279
rect 431 1243 445 1257
rect 815 1243 829 1257
rect 1151 1243 1165 1257
rect 1727 1243 1741 1257
rect 3383 1243 3397 1257
rect 3503 1243 3517 1257
rect 3623 1243 3637 1257
rect 3743 1243 3757 1257
rect 6887 1243 6901 1257
rect 7103 1243 7117 1257
rect 7223 1243 7237 1257
rect 311 1221 325 1235
rect 959 1221 973 1235
rect 1391 1221 1405 1235
rect 2831 1221 2845 1235
rect 4919 1221 4933 1235
rect 4991 1221 5005 1235
rect 5038 1221 5052 1235
rect 5351 1221 5365 1235
rect 5423 1221 5437 1235
rect 5855 1221 5869 1235
rect 6047 1221 6061 1235
rect 6095 1221 6109 1235
rect 6143 1221 6157 1235
rect 6239 1221 6253 1235
rect 6287 1221 6301 1235
rect 6503 1221 6517 1235
rect 6623 1221 6637 1235
rect 6743 1221 6757 1235
rect 6959 1221 6973 1235
rect 7199 1221 7213 1235
rect 191 1199 205 1213
rect 1703 1199 1717 1213
rect 2711 1199 2725 1213
rect 2807 1199 2821 1213
rect 5063 1199 5077 1213
rect 5231 1199 5245 1213
rect 5399 1199 5413 1213
rect 5471 1199 5485 1213
rect 5519 1199 5533 1213
rect 5975 1199 5989 1213
rect 6023 1199 6037 1213
rect 7247 1199 7261 1213
rect 7295 1199 7309 1213
rect 7343 1199 7357 1213
rect 239 380 253 394
rect 791 380 805 394
rect 1415 380 1429 394
rect 5543 380 5557 394
rect 6167 380 6181 394
rect 7367 380 7381 394
rect 359 358 373 372
rect 2735 358 2749 372
rect 5159 358 5173 372
rect 6191 358 6205 372
rect 6863 358 6877 372
rect 7007 358 7021 372
rect 7103 358 7117 372
rect 7151 358 7165 372
rect 479 336 493 350
rect 935 336 949 350
rect 1055 336 1069 350
rect 1751 336 1765 350
rect 2903 336 2917 350
rect 3023 336 3037 350
rect 3143 336 3157 350
rect 3263 336 3277 350
rect 5567 336 5581 350
rect 5783 336 5797 350
rect 5903 336 5917 350
rect 7031 336 7045 350
rect 599 314 613 328
rect 2927 314 2941 328
rect 3047 314 3061 328
rect 3407 314 3421 328
rect 3527 314 3541 328
rect 4151 314 4165 328
rect 4247 314 4261 328
rect 4343 314 4357 328
rect 4439 314 4453 328
rect 4535 314 4549 328
rect 4631 314 4645 328
rect 4727 314 4741 328
rect 4823 314 4837 328
rect 5136 314 5150 328
rect 5615 314 5629 328
rect 6335 314 6349 328
rect 6383 314 6397 328
rect 719 292 733 306
rect 911 292 925 306
rect 2951 292 2965 306
rect 3191 292 3205 306
rect 3431 292 3445 306
rect 3671 292 3685 306
rect 5807 292 5821 306
rect 7055 291 7069 305
rect 335 270 349 284
rect 1655 270 1669 284
rect 1991 270 2005 284
rect 2351 270 2365 284
rect 2855 269 2869 283
rect 3863 269 3877 283
rect 3959 269 3973 283
rect 4055 269 4069 283
rect 5779 270 5793 284
rect 6455 270 6469 284
rect 1799 248 1813 262
rect 1871 248 1885 262
rect 2759 247 2773 261
rect 4151 247 4165 261
rect 4339 248 4353 262
rect 4487 248 4501 262
rect 5567 248 5581 262
rect 6575 248 6589 262
rect 71 225 85 239
rect 3911 225 3925 239
rect 4007 225 4021 239
rect 5687 225 5701 239
rect 5975 226 5989 240
rect 6695 226 6709 240
rect 503 203 517 217
rect 2087 203 2101 217
rect 2231 203 2245 217
rect 4339 203 4353 217
rect 4679 203 4693 217
rect 6863 203 6877 217
rect 671 181 685 195
rect 2159 181 2173 195
rect 2879 181 2893 195
rect 4775 181 4789 195
rect 6335 181 6349 195
rect 6815 181 6829 195
rect 695 159 709 173
rect 2375 159 2389 173
rect 3215 159 3229 173
rect 4871 159 4885 173
rect 6695 159 6709 173
rect 7415 159 7429 173
rect 767 137 781 151
rect 2543 137 2557 151
rect 3335 137 3349 151
rect 5663 137 5677 151
rect 983 115 997 129
rect 2591 115 2605 129
rect 3383 115 3397 129
rect 4583 115 4597 129
rect 1127 93 1141 107
rect 5111 93 5125 107
rect 1463 71 1477 85
rect 4199 71 4213 85
rect 5111 69 5125 83
rect 5779 69 5793 83
rect 1823 49 1837 63
rect 4295 49 4309 63
rect 2567 27 2581 41
rect 4391 27 4405 41
rect 3551 5 3565 19
rect 4103 5 4117 19
<< metal2 >>
rect 192 1213 204 1481
rect 312 1235 324 1481
rect 432 1257 444 1481
rect 552 1279 564 1481
rect 672 1301 684 1481
rect 192 1196 204 1199
rect 312 1196 324 1221
rect 432 1196 444 1243
rect 552 1196 564 1265
rect 672 1196 684 1287
rect 816 1196 828 1243
rect 840 1196 852 1287
rect 864 1196 876 1353
rect 960 1196 972 1221
rect 984 1196 996 1331
rect 1032 1196 1044 1287
rect 1080 1196 1092 1309
rect 1128 1196 1140 1309
rect 1152 1196 1164 1243
rect 1200 1196 1212 1309
rect 1248 1196 1260 1331
rect 1272 1196 1284 1353
rect 1320 1196 1332 1331
rect 1368 1196 1380 1309
rect 1392 1196 1404 1221
rect 1440 1196 1452 1309
rect 1488 1196 1500 1331
rect 1512 1196 1524 1265
rect 1536 1196 1548 1331
rect 1584 1196 1596 1309
rect 1608 1196 1620 1331
rect 1704 1196 1716 1199
rect 1728 1196 1740 1243
rect 1848 1196 1860 1481
rect 1920 1196 1932 1309
rect 1968 1196 1980 1309
rect 2184 1196 2196 1309
rect 2280 1196 2292 1481
rect 2472 1323 2484 1481
rect 2472 1196 2484 1309
rect 2544 1196 2556 1481
rect 2640 1196 2652 1481
rect 2712 1196 2724 1199
rect 2808 1196 2820 1199
rect 2832 1196 2844 1221
rect 2976 1196 2988 1375
rect 3072 1196 3084 1287
rect 3096 1196 3108 1397
rect 3168 1196 3180 1265
rect 3216 1196 3228 1309
rect 3288 1196 3300 1265
rect 3312 1196 3324 1287
rect 3336 1196 3348 1419
rect 3384 1196 3396 1243
rect 3456 1196 3468 1331
rect 3504 1196 3516 1243
rect 3552 1196 3564 1287
rect 3576 1196 3588 1440
rect 3624 1196 3636 1243
rect 3648 1196 3660 1265
rect 3696 1196 3708 1462
rect 3744 1196 3756 1243
rect 3768 1196 3780 1265
rect 3792 1196 3804 1287
rect 3816 1196 3828 1353
rect 3888 1196 3900 1309
rect 3984 1196 3996 1331
rect 4080 1196 4092 1353
rect 4176 1196 4188 1375
rect 4272 1196 4284 1396
rect 4368 1196 4380 1309
rect 4464 1196 4476 1418
rect 4560 1196 4572 1331
rect 4584 1196 4596 1309
rect 4656 1196 4668 1440
rect 4752 1196 4764 1462
rect 4848 1196 4860 1353
rect 4920 1196 4932 1221
rect 4944 1196 4956 1265
rect 4968 1196 4980 1287
rect 4992 1196 5004 1221
rect 5040 1196 5052 1221
rect 5064 1196 5076 1199
rect 5184 1196 5196 1265
rect 5232 1196 5244 1199
rect 5280 1196 5292 1265
rect 5304 1196 5316 1287
rect 5352 1196 5364 1221
rect 5400 1196 5412 1199
rect 5424 1196 5436 1221
rect 5472 1196 5484 1199
rect 5520 1196 5532 1199
rect 5856 1196 5868 1221
rect 5928 1196 5940 1265
rect 5976 1196 5988 1199
rect 6024 1196 6036 1199
rect 6048 1196 6060 1221
rect 6096 1196 6108 1221
rect 6144 1196 6156 1221
rect 6240 1196 6252 1221
rect 6288 1196 6300 1221
rect 6312 1196 6324 1481
rect 6408 1196 6420 1309
rect 6504 1196 6516 1221
rect 6528 1196 6540 1481
rect 6624 1196 6636 1221
rect 6648 1196 6660 1481
rect 6744 1196 6756 1221
rect 6768 1196 6780 1481
rect 6888 1196 6900 1243
rect 6912 1196 6924 1265
rect 6960 1196 6972 1221
rect 7104 1196 7116 1243
rect 7152 1196 7164 1481
rect 7200 1196 7212 1221
rect 7224 1196 7236 1243
rect 7248 1196 7260 1199
rect 7296 1196 7308 1199
rect 7344 1196 7356 1199
rect 240 394 252 397
rect 360 372 372 397
rect 480 350 492 397
rect 600 328 612 397
rect 720 306 732 397
rect 792 394 804 397
rect 912 306 924 397
rect 936 350 948 397
rect 1056 350 1068 397
rect 1416 394 1428 397
rect 1656 284 1668 397
rect 1752 350 1764 397
rect 72 -143 84 225
rect 336 -143 348 270
rect 1800 262 1812 397
rect 1872 262 1884 397
rect 1992 284 2004 397
rect 2088 217 2100 397
rect 504 -143 516 203
rect 2160 195 2172 397
rect 2352 284 2364 397
rect 672 -143 684 181
rect 696 -143 708 159
rect 768 -143 780 137
rect 984 -143 996 115
rect 1128 -143 1140 93
rect 1464 -143 1476 71
rect 1824 -143 1836 49
rect 2232 -143 2244 203
rect 2376 173 2388 397
rect 2544 151 2556 397
rect 2592 129 2604 397
rect 2736 372 2748 397
rect 2760 261 2772 397
rect 2856 283 2868 397
rect 2904 350 2916 397
rect 2928 328 2940 397
rect 2952 306 2964 397
rect 3024 350 3036 397
rect 3048 328 3060 397
rect 3144 350 3156 397
rect 3192 306 3204 397
rect 3264 350 3276 397
rect 3408 328 3420 397
rect 3432 306 3444 397
rect 3528 328 3540 397
rect 3672 306 3684 397
rect 3864 283 3876 397
rect 3912 239 3924 397
rect 3960 283 3972 397
rect 4008 239 4020 397
rect 4056 283 4068 397
rect 2568 -143 2580 27
rect 2880 -143 2892 181
rect 3216 -143 3228 159
rect 3336 -143 3348 137
rect 3384 -143 3396 115
rect 4104 19 4116 397
rect 4152 328 4164 397
rect 4152 261 4164 314
rect 4200 85 4212 397
rect 4248 328 4260 397
rect 4296 63 4308 397
rect 4344 328 4356 397
rect 4340 217 4352 248
rect 4392 41 4404 397
rect 4440 328 4452 397
rect 4488 262 4500 397
rect 4536 328 4548 397
rect 4584 129 4596 397
rect 4632 328 4644 397
rect 4680 217 4692 397
rect 4728 328 4740 397
rect 4776 195 4788 397
rect 4824 328 4836 397
rect 4872 173 4884 397
rect 5112 107 5124 397
rect 5160 372 5172 397
rect 5544 394 5556 397
rect 5568 350 5580 397
rect 5616 328 5628 397
rect 3552 -143 3564 5
rect 5112 -143 5124 69
rect 5137 -143 5149 314
rect 5568 -143 5580 248
rect 5664 151 5676 397
rect 5688 239 5700 397
rect 5736 -143 5748 397
rect 5784 350 5796 397
rect 5808 306 5820 397
rect 5904 350 5916 397
rect 6168 394 6180 397
rect 6192 372 6204 397
rect 6336 328 6348 397
rect 6384 328 6396 397
rect 6456 284 6468 397
rect 5780 83 5792 270
rect 6576 262 6588 397
rect 6696 240 6708 397
rect 5976 -143 5988 226
rect 6816 195 6828 397
rect 6864 372 6876 397
rect 7008 372 7020 397
rect 7032 350 7044 397
rect 7056 305 7068 397
rect 7152 372 7164 508
rect 7368 394 7380 397
rect 6336 -143 6348 181
rect 6696 -143 6708 159
rect 6864 -143 6876 203
rect 7104 -143 7116 358
rect 7416 173 7428 397
use inv  inv_0
timestamp 1386238110
transform 1 0 168 0 1 397
box 0 0 120 799
use inv  inv_1
timestamp 1386238110
transform 1 0 288 0 1 397
box 0 0 120 799
use inv  inv_2
timestamp 1386238110
transform 1 0 408 0 1 397
box 0 0 120 799
use inv  inv_3
timestamp 1386238110
transform 1 0 528 0 1 397
box 0 0 120 799
use inv  inv_4
timestamp 1386238110
transform 1 0 648 0 1 397
box 0 0 120 799
use nand3  nand3_0
timestamp 1386234893
transform 1 0 768 0 1 397
box 0 0 120 799
use nand3  nand3_1
timestamp 1386234893
transform 1 0 888 0 1 397
box 0 0 120 799
use nand2  nand2_0
timestamp 1386234792
transform 1 0 1008 0 1 397
box 0 0 96 799
use nor2  nor2_0
timestamp 1386235306
transform 1 0 1104 0 1 397
box 0 0 120 799
use nor2  nor2_1
timestamp 1386235306
transform 1 0 1224 0 1 397
box 0 0 120 799
use nand3  nand3_2
timestamp 1386234893
transform 1 0 1344 0 1 397
box 0 0 120 799
use nand2  nand2_1
timestamp 1386234792
transform 1 0 1464 0 1 397
box 0 0 96 799
use nor2  nor2_2
timestamp 1386235306
transform 1 0 1560 0 1 397
box 0 0 120 799
use nor3  nor3_0
timestamp 1386235396
transform 1 0 1680 0 1 397
box 0 0 144 799
use and2  and2_4
timestamp 1386234845
transform 1 0 1824 0 1 397
box 0 0 120 799
use xor2  xor2_3
timestamp 1386237344
transform 1 0 1944 0 1 397
box 0 0 192 799
use xor2  xor2_4
timestamp 1386237344
transform 1 0 2136 0 1 397
box 0 0 192 799
use xor2  xor2_5
timestamp 1386237344
transform 1 0 2328 0 1 397
box 0 0 192 799
use rowcrosser  rowcrosser_1
timestamp 1386086759
transform 1 0 2520 0 1 397
box 0 0 48 799
use inv  inv_6
timestamp 1386238110
transform 1 0 2568 0 1 397
box 0 0 120 799
use nand2  nand2_2
timestamp 1386234792
transform 1 0 2688 0 1 397
box 0 0 96 799
use nand2  nand2_3
timestamp 1386234792
transform 1 0 2784 0 1 397
box 0 0 96 799
use nand3  nand3_4
timestamp 1386234893
transform 1 0 2880 0 1 397
box 0 0 120 799
use nand3  nand3_5
timestamp 1386234893
transform 1 0 3000 0 1 397
box 0 0 120 799
use nand3  nand3_6
timestamp 1386234893
transform 1 0 3120 0 1 397
box 0 0 120 799
use nand3  nand3_7
timestamp 1386234893
transform 1 0 3240 0 1 397
box 0 0 120 799
use nand3  nand3_8
timestamp 1386234893
transform 1 0 3360 0 1 397
box 0 0 120 799
use nand3  nand3_9
timestamp 1386234893
transform 1 0 3480 0 1 397
box 0 0 120 799
use nand3  nand3_10
timestamp 1386234893
transform 1 0 3600 0 1 397
box 0 0 120 799
use nand3  nand3_11
timestamp 1386234893
transform 1 0 3720 0 1 397
box 0 0 120 799
use nand2  nand2_4
timestamp 1386234792
transform 1 0 3840 0 1 397
box 0 0 96 799
use nand2  nand2_5
timestamp 1386234792
transform 1 0 3936 0 1 397
box 0 0 96 799
use nand2  nand2_6
timestamp 1386234792
transform 1 0 4032 0 1 397
box 0 0 96 799
use nand2  nand2_7
timestamp 1386234792
transform 1 0 4128 0 1 397
box 0 0 96 799
use nand2  nand2_8
timestamp 1386234792
transform 1 0 4224 0 1 397
box 0 0 96 799
use nand2  nand2_9
timestamp 1386234792
transform 1 0 4320 0 1 397
box 0 0 96 799
use nand2  nand2_10
timestamp 1386234792
transform 1 0 4416 0 1 397
box 0 0 96 799
use nand2  nand2_11
timestamp 1386234792
transform 1 0 4512 0 1 397
box 0 0 96 799
use nand2  nand2_12
timestamp 1386234792
transform 1 0 4608 0 1 397
box 0 0 96 799
use nand2  nand2_13
timestamp 1386234792
transform 1 0 4704 0 1 397
box 0 0 96 799
use nand2  nand2_14
timestamp 1386234792
transform 1 0 4800 0 1 397
box 0 0 96 799
use nand3  nand3_3
timestamp 1386234893
transform 1 0 4896 0 1 397
box 0 0 120 799
use nor2  nor2_3
timestamp 1386235306
transform 1 0 5016 0 1 397
box 0 0 120 799
use nor2  nor2_4
timestamp 1386235306
transform 1 0 5136 0 1 397
box 0 0 120 799
use nor2  nor2_5
timestamp 1386235306
transform 1 0 5256 0 1 397
box 0 0 120 799
use nor2  nor2_6
timestamp 1386235306
transform 1 0 5376 0 1 397
box 0 0 120 799
use nor3  nor3_1
timestamp 1386235396
transform 1 0 5496 0 1 397
box 0 0 144 799
use and2  and2_3
timestamp 1386234845
transform 1 0 5640 0 1 397
box 0 0 120 799
use nor2  nor2_7
timestamp 1386235306
transform 1 0 5760 0 1 397
box 0 0 120 799
use nor2  nor2_8
timestamp 1386235306
transform 1 0 5880 0 1 397
box 0 0 120 799
use nor2  nor2_9
timestamp 1386235306
transform 1 0 6000 0 1 397
box 0 0 120 799
use nor3  nor3_2
timestamp 1386235396
transform 1 0 6120 0 1 397
box 0 0 144 799
use nand2  nand2_15
timestamp 1386234792
transform 1 0 6264 0 1 397
box 0 0 96 799
use nor2  nor2_10
timestamp 1386235306
transform 1 0 6360 0 1 397
box 0 0 120 799
use and2  and2_0
timestamp 1386234845
transform 1 0 6480 0 1 397
box 0 0 120 799
use and2  and2_1
timestamp 1386234845
transform 1 0 6600 0 1 397
box 0 0 120 799
use and2  and2_2
timestamp 1386234845
transform 1 0 6720 0 1 397
box 0 0 120 799
use nor3  nor3_3
timestamp 1386235396
transform 1 0 6840 0 1 397
box 0 0 144 799
use nor3  nor3_4
timestamp 1386235396
transform 1 0 6984 0 1 397
box 0 0 144 799
use rowcrosser  rowcrosser_0
timestamp 1386086759
transform 1 0 7128 0 1 397
box 0 0 48 799
use nor3  nor3_5
timestamp 1386235396
transform 1 0 7176 0 1 397
box 0 0 144 799
use nor2  nor2_11
timestamp 1386235306
transform 1 0 7320 0 1 397
box 0 0 120 799
<< labels >>
rlabel metal1 504 344 504 344 1 nC
rlabel metal1 747 297 747 297 1 nE
rlabel metal1 272 386 272 386 1 nA
rlabel metal1 378 364 378 364 1 nB
rlabel metal1 627 319 627 319 1 nD
rlabel metal2 192 1481 204 1481 5 OpCode[4]
rlabel metal2 312 1481 324 1481 5 OpCode[3]
rlabel metal2 432 1481 444 1481 5 OpCode[2]
rlabel metal2 552 1481 564 1481 5 OpCode[1]
rlabel metal2 672 1481 684 1481 5 OpCode[0]
rlabel metal2 2640 1481 2652 1481 5 Z
rlabel metal2 2544 1481 2556 1481 5 N
rlabel metal2 2280 1481 2292 1481 5 V
rlabel metal2 1848 1481 1860 1481 5 Cin
rlabel metal2 2472 1481 2484 1481 5 C
rlabel metal2 6768 1481 6780 1481 5 imm4[0]
rlabel metal2 6648 1481 6660 1481 5 imm4[1]
rlabel metal2 6528 1481 6540 1481 5 imm4[2]
rlabel metal2 6312 1481 6324 1481 5 imm4[3]
rlabel metal2 6245 1198 6245 1198 1 N
rlabel metal1 5502 231 5502 231 1 ShSign
rlabel metal1 0 1118 0 1143 3 Vdd!
rlabel metal1 0 473 0 498 3 GND!
rlabel metal2 7152 1481 7164 1481 5 OutEn
rlabel metal1 0 1156 0 1166 3 Scan
rlabel metal1 0 1179 0 1189 3 ScanReturn
rlabel metal1 0 404 0 414 3 nReset
rlabel metal1 0 427 0 437 3 Test
rlabel metal1 0 450 0 460 3 Clock
rlabel metal2 5736 -143 5748 -143 1 ShInBit
rlabel metal2 2880 -143 2892 -143 1 NAND
rlabel metal2 336 -143 348 -143 1 SUB
rlabel metal2 504 -143 516 -143 1 CIn_slice
rlabel metal2 672 -143 684 -143 1 LastCIn
rlabel metal2 696 -143 708 -143 1 COut
rlabel metal2 984 -143 996 -143 1 nZ
rlabel metal2 1128 -143 1140 -143 1 FAOut
rlabel metal2 1464 -143 1476 -143 1 AND
rlabel metal2 1824 -143 1836 -143 1 OR
rlabel metal2 2232 -143 2244 -143 1 XOR
rlabel metal2 2568 -143 2580 -143 1 NOT
rlabel metal2 3552 -143 3564 -143 1 ShL
rlabel metal2 5137 -143 5149 -143 1 ShR
rlabel metal2 6696 -143 6708 -143 1 ShOut
rlabel metal2 3336 -143 3348 -143 1 ASign
rlabel metal2 3384 -143 3396 -143 1 ShB
rlabel metal2 5112 -143 5124 -143 1 Sh8
rlabel metal2 5568 -143 5580 -143 1 Sh4
rlabel metal2 5976 -143 5988 -143 1 Sh2
rlabel metal2 6336 -143 6348 -143 1 Sh1
rlabel metal2 3216 -143 3228 -143 1 NOR
rlabel metal2 768 -143 780 -143 1 N
rlabel metal2 72 -143 84 -143 1 ZeroA
rlabel metal2 6864 -143 6876 -143 1 LLI
rlabel metal2 7104 -143 7116 -143 1 Outen
<< end >>
