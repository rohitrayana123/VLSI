magic
tech c035u
timestamp 1395342641
<< metal4 >>
rect 6166 49274 7726 50834
rect 10638 49274 12198 50834
rect 15110 49274 16670 50834
rect 19582 49274 21142 50834
rect 24054 49274 25614 50834
rect 28526 49274 30086 50834
rect 32998 49274 34558 50834
rect 37470 49274 39030 50834
rect 41942 49274 43502 50834
rect -544 42736 1016 44296
rect 48652 42736 50212 44296
rect -544 37576 1016 39136
rect 48652 37576 50212 39136
rect -544 32416 1016 33976
rect 48652 32416 50212 33976
rect -544 27256 1016 28816
rect 48652 27256 50212 28816
rect -544 22096 1016 23656
rect 48652 22096 50212 23656
rect -544 16936 1016 18496
rect 48652 16936 50212 18496
rect -544 11776 1016 13336
rect 48652 11776 50212 13336
rect -544 6616 1016 8176
rect 48652 6616 50212 8176
rect 6166 78 7726 1638
rect 10638 78 12198 1638
rect 15110 78 16670 1638
rect 19582 78 21142 1638
rect 24054 78 25614 1638
rect 28526 78 30086 1638
rect 32998 78 34558 1638
rect 37470 78 39030 1638
rect 41942 78 43502 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 -622 -1 0 50912
box 0 0 6450 6450
use fillpp_mt fillpp_mt_805
timestamp 1300117811
transform 0 -1 5914 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_804
timestamp 1300117811
transform 0 -1 6000 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_803
timestamp 1300117811
transform 0 -1 6086 1 0 44462
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 7806 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_802
timestamp 1300117811
transform 0 -1 7892 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_801
timestamp 1300117811
transform 0 -1 7978 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_800
timestamp 1300117811
transform 0 -1 8064 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_799
timestamp 1300117811
transform 0 -1 8150 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_798
timestamp 1300117811
transform 0 -1 8236 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_797
timestamp 1300117811
transform 0 -1 8322 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_796
timestamp 1300117811
transform 0 -1 8408 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_795
timestamp 1300117811
transform 0 -1 8494 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_794
timestamp 1300117811
transform 0 -1 8580 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_793
timestamp 1300117811
transform 0 -1 8666 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_792
timestamp 1300117811
transform 0 -1 8752 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_791
timestamp 1300117811
transform 0 -1 8838 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_790
timestamp 1300117811
transform 0 -1 8924 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_789
timestamp 1300117811
transform 0 -1 9010 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_788
timestamp 1300117811
transform 0 -1 9096 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform 0 -1 9182 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform 0 -1 9268 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform 0 -1 9354 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform 0 -1 9440 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform 0 -1 9526 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform 0 -1 9612 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform 0 -1 9698 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform 0 -1 9784 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform 0 -1 9870 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform 0 -1 9956 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform 0 -1 10042 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform 0 -1 10128 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform 0 -1 10214 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform 0 -1 10300 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform 0 -1 10386 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform 0 -1 10472 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform 0 -1 10558 1 0 44462
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 12278 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform 0 -1 12364 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform 0 -1 12450 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform 0 -1 12536 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform 0 -1 12622 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform 0 -1 12708 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform 0 -1 12794 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform 0 -1 12880 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform 0 -1 12966 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform 0 -1 13052 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform 0 -1 13138 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform 0 -1 13224 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform 0 -1 13310 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform 0 -1 13396 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform 0 -1 13482 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform 0 -1 13568 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform 0 -1 13654 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform 0 -1 13740 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform 0 -1 13826 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform 0 -1 13912 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform 0 -1 13998 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform 0 -1 14084 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform 0 -1 14170 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform 0 -1 14256 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform 0 -1 14342 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform 0 -1 14428 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform 0 -1 14514 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform 0 -1 14600 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform 0 -1 14686 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform 0 -1 14772 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform 0 -1 14858 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform 0 -1 14944 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform 0 -1 15030 1 0 44462
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 16750 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform 0 -1 16836 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform 0 -1 16922 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform 0 -1 17008 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform 0 -1 17094 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform 0 -1 17180 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform 0 -1 17266 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform 0 -1 17352 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform 0 -1 17438 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform 0 -1 17524 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform 0 -1 17610 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform 0 -1 17696 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform 0 -1 17782 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform 0 -1 17868 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform 0 -1 17954 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform 0 -1 18040 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform 0 -1 18126 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform 0 -1 18212 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform 0 -1 18298 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform 0 -1 18384 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform 0 -1 18470 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform 0 -1 18556 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform 0 -1 18642 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform 0 -1 18728 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform 0 -1 18814 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform 0 -1 18900 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform 0 -1 18986 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform 0 -1 19072 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform 0 -1 19158 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform 0 -1 19244 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform 0 -1 19330 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform 0 -1 19416 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform 0 -1 19502 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 21222 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform 0 -1 21308 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform 0 -1 21394 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform 0 -1 21480 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform 0 -1 21566 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform 0 -1 21652 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform 0 -1 21738 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform 0 -1 21824 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform 0 -1 21910 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform 0 -1 21996 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform 0 -1 22082 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform 0 -1 22168 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform 0 -1 22254 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform 0 -1 22340 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform 0 -1 22426 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform 0 -1 22512 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform 0 -1 22598 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform 0 -1 22684 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform 0 -1 22770 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform 0 -1 22856 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform 0 -1 22942 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform 0 -1 23028 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform 0 -1 23114 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform 0 -1 23200 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform 0 -1 23286 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform 0 -1 23372 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform 0 -1 23458 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform 0 -1 23544 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform 0 -1 23630 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform 0 -1 23716 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform 0 -1 23802 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform 0 -1 23888 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform 0 -1 23974 1 0 44462
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 25694 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform 0 -1 25780 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform 0 -1 25866 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform 0 -1 25952 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform 0 -1 26038 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform 0 -1 26124 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform 0 -1 26210 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform 0 -1 26296 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform 0 -1 26382 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform 0 -1 26468 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform 0 -1 26554 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform 0 -1 26640 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform 0 -1 26726 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform 0 -1 26812 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform 0 -1 26898 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform 0 -1 26984 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform 0 -1 27070 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform 0 -1 27156 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform 0 -1 27242 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform 0 -1 27328 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform 0 -1 27414 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform 0 -1 27500 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform 0 -1 27586 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform 0 -1 27672 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform 0 -1 27758 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform 0 -1 27844 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform 0 -1 27930 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform 0 -1 28016 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform 0 -1 28102 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform 0 -1 28188 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform 0 -1 28274 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform 0 -1 28360 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform 0 -1 28446 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 30166 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform 0 -1 30252 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform 0 -1 30338 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform 0 -1 30424 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform 0 -1 30510 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform 0 -1 30596 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform 0 -1 30682 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform 0 -1 30768 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform 0 -1 30854 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform 0 -1 30940 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform 0 -1 31026 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform 0 -1 31112 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform 0 -1 31198 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform 0 -1 31284 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform 0 -1 31370 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform 0 -1 31456 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform 0 -1 31542 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform 0 -1 31628 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform 0 -1 31714 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform 0 -1 31800 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform 0 -1 31886 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform 0 -1 31972 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform 0 -1 32058 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform 0 -1 32144 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform 0 -1 32230 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform 0 -1 32316 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform 0 -1 32402 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform 0 -1 32488 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform 0 -1 32574 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform 0 -1 32660 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform 0 -1 32746 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform 0 -1 32832 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform 0 -1 32918 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 34638 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform 0 -1 34724 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform 0 -1 34810 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform 0 -1 34896 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform 0 -1 34982 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform 0 -1 35068 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform 0 -1 35154 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform 0 -1 35240 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform 0 -1 35326 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform 0 -1 35412 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform 0 -1 35498 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform 0 -1 35584 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform 0 -1 35670 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform 0 -1 35756 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform 0 -1 35842 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform 0 -1 35928 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform 0 -1 36014 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform 0 -1 36100 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform 0 -1 36186 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform 0 -1 36272 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform 0 -1 36358 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform 0 -1 36444 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform 0 -1 36530 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform 0 -1 36616 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform 0 -1 36702 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform 0 -1 36788 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform 0 -1 36874 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform 0 -1 36960 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform 0 -1 37046 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform 0 -1 37132 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform 0 -1 37218 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform 0 -1 37304 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform 0 -1 37390 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 39110 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform 0 -1 39196 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform 0 -1 39282 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform 0 -1 39368 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform 0 -1 39454 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform 0 -1 39540 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform 0 -1 39626 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform 0 -1 39712 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform 0 -1 39798 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform 0 -1 39884 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform 0 -1 39970 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform 0 -1 40056 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform 0 -1 40142 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform 0 -1 40228 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform 0 -1 40314 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform 0 -1 40400 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 40486 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 40572 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 40658 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 40744 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 40830 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 40916 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 41002 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 41088 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 41174 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 41260 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 41346 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 41432 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 41518 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 41604 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 41690 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 41776 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 41862 1 0 44462
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 43582 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 43668 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 43754 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 43840 1 0 44462
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 50290 0 -1 50912
box 0 0 6450 6450
use fillpp_mt fillpp_mt_806
timestamp 1300117811
transform -1 0 5828 0 -1 44462
box 0 0 6450 86
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 5828 0 -1 44376
box 0 0 6450 1720
use fillpp_mt fillpp_mt_807
timestamp 1300117811
transform -1 0 5828 0 -1 42656
box 0 0 6450 86
use fillpp_mt fillpp_mt_808
timestamp 1300117811
transform -1 0 5828 0 -1 42570
box 0 0 6450 86
use fillpp_mt fillpp_mt_809
timestamp 1300117811
transform -1 0 5828 0 -1 42484
box 0 0 6450 86
use fillpp_mt fillpp_mt_810
timestamp 1300117811
transform -1 0 5828 0 -1 42398
box 0 0 6450 86
use fillpp_mt fillpp_mt_811
timestamp 1300117811
transform -1 0 5828 0 -1 42312
box 0 0 6450 86
use fillpp_mt fillpp_mt_812
timestamp 1300117811
transform -1 0 5828 0 -1 42226
box 0 0 6450 86
use fillpp_mt fillpp_mt_813
timestamp 1300117811
transform -1 0 5828 0 -1 42140
box 0 0 6450 86
use fillpp_mt fillpp_mt_814
timestamp 1300117811
transform -1 0 5828 0 -1 42054
box 0 0 6450 86
use fillpp_mt fillpp_mt_815
timestamp 1300117811
transform -1 0 5828 0 -1 41968
box 0 0 6450 86
use fillpp_mt fillpp_mt_816
timestamp 1300117811
transform -1 0 5828 0 -1 41882
box 0 0 6450 86
use fillpp_mt fillpp_mt_817
timestamp 1300117811
transform -1 0 5828 0 -1 41796
box 0 0 6450 86
use fillpp_mt fillpp_mt_818
timestamp 1300117811
transform -1 0 5828 0 -1 41710
box 0 0 6450 86
use fillpp_mt fillpp_mt_819
timestamp 1300117811
transform -1 0 5828 0 -1 41624
box 0 0 6450 86
use fillpp_mt fillpp_mt_820
timestamp 1300117811
transform -1 0 5828 0 -1 41538
box 0 0 6450 86
use fillpp_mt fillpp_mt_821
timestamp 1300117811
transform -1 0 5828 0 -1 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_822
timestamp 1300117811
transform -1 0 5828 0 -1 41366
box 0 0 6450 86
use fillpp_mt fillpp_mt_823
timestamp 1300117811
transform -1 0 5828 0 -1 41280
box 0 0 6450 86
use fillpp_mt fillpp_mt_824
timestamp 1300117811
transform -1 0 5828 0 -1 41194
box 0 0 6450 86
use fillpp_mt fillpp_mt_825
timestamp 1300117811
transform -1 0 5828 0 -1 41108
box 0 0 6450 86
use fillpp_mt fillpp_mt_826
timestamp 1300117811
transform -1 0 5828 0 -1 41022
box 0 0 6450 86
use fillpp_mt fillpp_mt_827
timestamp 1300117811
transform -1 0 5828 0 -1 40936
box 0 0 6450 86
use fillpp_mt fillpp_mt_828
timestamp 1300117811
transform -1 0 5828 0 -1 40850
box 0 0 6450 86
use fillpp_mt fillpp_mt_829
timestamp 1300117811
transform -1 0 5828 0 -1 40764
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 1 0 43840 0 1 44376
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 43840 0 1 42656
box 0 0 6450 1720
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 1 0 43840 0 1 42570
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 1 0 43840 0 1 42484
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 1 0 43840 0 1 42398
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 1 0 43840 0 1 42312
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 1 0 43840 0 1 42226
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 1 0 43840 0 1 42140
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 1 0 43840 0 1 42054
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 1 0 43840 0 1 41968
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 1 0 43840 0 1 41882
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 1 0 43840 0 1 41796
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 1 0 43840 0 1 41710
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 1 0 43840 0 1 41624
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 1 0 43840 0 1 41538
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 1 0 43840 0 1 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 1 0 43840 0 1 41366
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 1 0 43840 0 1 41280
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 1 0 43840 0 1 41194
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 1 0 43840 0 1 41108
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 1 0 43840 0 1 41022
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 1 0 43840 0 1 40936
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 1 0 43840 0 1 40850
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 1 0 43840 0 1 40764
box 0 0 6450 86
use fillpp_mt fillpp_mt_830
timestamp 1300117811
transform -1 0 5828 0 -1 40678
box 0 0 6450 86
use fillpp_mt fillpp_mt_831
timestamp 1300117811
transform -1 0 5828 0 -1 40592
box 0 0 6450 86
use fillpp_mt fillpp_mt_832
timestamp 1300117811
transform -1 0 5828 0 -1 40506
box 0 0 6450 86
use fillpp_mt fillpp_mt_833
timestamp 1300117811
transform -1 0 5828 0 -1 40420
box 0 0 6450 86
use fillpp_mt fillpp_mt_834
timestamp 1300117811
transform -1 0 5828 0 -1 40334
box 0 0 6450 86
use fillpp_mt fillpp_mt_835
timestamp 1300117811
transform -1 0 5828 0 -1 40248
box 0 0 6450 86
use fillpp_mt fillpp_mt_836
timestamp 1300117811
transform -1 0 5828 0 -1 40162
box 0 0 6450 86
use fillpp_mt fillpp_mt_837
timestamp 1300117811
transform -1 0 5828 0 -1 40076
box 0 0 6450 86
use fillpp_mt fillpp_mt_838
timestamp 1300117811
transform -1 0 5828 0 -1 39990
box 0 0 6450 86
use fillpp_mt fillpp_mt_839
timestamp 1300117811
transform -1 0 5828 0 -1 39904
box 0 0 6450 86
use fillpp_mt fillpp_mt_840
timestamp 1300117811
transform -1 0 5828 0 -1 39818
box 0 0 6450 86
use fillpp_mt fillpp_mt_841
timestamp 1300117811
transform -1 0 5828 0 -1 39732
box 0 0 6450 86
use fillpp_mt fillpp_mt_842
timestamp 1300117811
transform -1 0 5828 0 -1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_843
timestamp 1300117811
transform -1 0 5828 0 -1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_844
timestamp 1300117811
transform -1 0 5828 0 -1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_845
timestamp 1300117811
transform -1 0 5828 0 -1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_846
timestamp 1300117811
transform -1 0 5828 0 -1 39302
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 5828 0 -1 39216
box 0 0 6450 1720
use fillpp_mt fillpp_mt_847
timestamp 1300117811
transform -1 0 5828 0 -1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_848
timestamp 1300117811
transform -1 0 5828 0 -1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_849
timestamp 1300117811
transform -1 0 5828 0 -1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_850
timestamp 1300117811
transform -1 0 5828 0 -1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_851
timestamp 1300117811
transform -1 0 5828 0 -1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_852
timestamp 1300117811
transform -1 0 5828 0 -1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_853
timestamp 1300117811
transform -1 0 5828 0 -1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_854
timestamp 1300117811
transform -1 0 5828 0 -1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_855
timestamp 1300117811
transform -1 0 5828 0 -1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_856
timestamp 1300117811
transform -1 0 5828 0 -1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_857
timestamp 1300117811
transform -1 0 5828 0 -1 36636
box 0 0 6450 86
use fillpp_mt fillpp_mt_858
timestamp 1300117811
transform -1 0 5828 0 -1 36550
box 0 0 6450 86
use fillpp_mt fillpp_mt_859
timestamp 1300117811
transform -1 0 5828 0 -1 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_860
timestamp 1300117811
transform -1 0 5828 0 -1 36378
box 0 0 6450 86
use fillpp_mt fillpp_mt_861
timestamp 1300117811
transform -1 0 5828 0 -1 36292
box 0 0 6450 86
use fillpp_mt fillpp_mt_862
timestamp 1300117811
transform -1 0 5828 0 -1 36206
box 0 0 6450 86
use fillpp_mt fillpp_mt_863
timestamp 1300117811
transform -1 0 5828 0 -1 36120
box 0 0 6450 86
use fillpp_mt fillpp_mt_864
timestamp 1300117811
transform -1 0 5828 0 -1 36034
box 0 0 6450 86
use fillpp_mt fillpp_mt_865
timestamp 1300117811
transform -1 0 5828 0 -1 35948
box 0 0 6450 86
use fillpp_mt fillpp_mt_866
timestamp 1300117811
transform -1 0 5828 0 -1 35862
box 0 0 6450 86
use fillpp_mt fillpp_mt_867
timestamp 1300117811
transform -1 0 5828 0 -1 35776
box 0 0 6450 86
use fillpp_mt fillpp_mt_868
timestamp 1300117811
transform -1 0 5828 0 -1 35690
box 0 0 6450 86
use fillpp_mt fillpp_mt_869
timestamp 1300117811
transform -1 0 5828 0 -1 35604
box 0 0 6450 86
use fillpp_mt fillpp_mt_870
timestamp 1300117811
transform -1 0 5828 0 -1 35518
box 0 0 6450 86
use fillpp_mt fillpp_mt_871
timestamp 1300117811
transform -1 0 5828 0 -1 35432
box 0 0 6450 86
use fillpp_mt fillpp_mt_872
timestamp 1300117811
transform -1 0 5828 0 -1 35346
box 0 0 6450 86
use fillpp_mt fillpp_mt_873
timestamp 1300117811
transform -1 0 5828 0 -1 35260
box 0 0 6450 86
use fillpp_mt fillpp_mt_874
timestamp 1300117811
transform -1 0 5828 0 -1 35174
box 0 0 6450 86
use fillpp_mt fillpp_mt_875
timestamp 1300117811
transform -1 0 5828 0 -1 35088
box 0 0 6450 86
use fillpp_mt fillpp_mt_876
timestamp 1300117811
transform -1 0 5828 0 -1 35002
box 0 0 6450 86
use fillpp_mt fillpp_mt_877
timestamp 1300117811
transform -1 0 5828 0 -1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_878
timestamp 1300117811
transform -1 0 5828 0 -1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_879
timestamp 1300117811
transform -1 0 5828 0 -1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_880
timestamp 1300117811
transform -1 0 5828 0 -1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_881
timestamp 1300117811
transform -1 0 5828 0 -1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_882
timestamp 1300117811
transform -1 0 5828 0 -1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_883
timestamp 1300117811
transform -1 0 5828 0 -1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_884
timestamp 1300117811
transform -1 0 5828 0 -1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_885
timestamp 1300117811
transform -1 0 5828 0 -1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_886
timestamp 1300117811
transform -1 0 5828 0 -1 34142
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 5828 0 -1 34056
box 0 0 6450 1720
use control control_0
timestamp 1395324901
transform 1 0 12032 0 1 32499
box 0 0 28280 8252
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 1 0 43840 0 1 40678
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 1 0 43840 0 1 40592
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 1 0 43840 0 1 40506
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 1 0 43840 0 1 40420
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 1 0 43840 0 1 40334
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 1 0 43840 0 1 40248
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 1 0 43840 0 1 40162
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 1 0 43840 0 1 40076
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 1 0 43840 0 1 39990
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 1 0 43840 0 1 39904
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 1 0 43840 0 1 39818
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 1 0 43840 0 1 39732
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 1 0 43840 0 1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 1 0 43840 0 1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 1 0 43840 0 1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 1 0 43840 0 1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 1 0 43840 0 1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 1 0 43840 0 1 39216
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 43840 0 1 37496
box 0 0 6450 1720
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 1 0 43840 0 1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 1 0 43840 0 1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 1 0 43840 0 1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 1 0 43840 0 1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 1 0 43840 0 1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 1 0 43840 0 1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 1 0 43840 0 1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 1 0 43840 0 1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 1 0 43840 0 1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 1 0 43840 0 1 36636
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 1 0 43840 0 1 36550
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 1 0 43840 0 1 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 1 0 43840 0 1 36378
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 1 0 43840 0 1 36292
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 1 0 43840 0 1 36206
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 1 0 43840 0 1 36120
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 1 0 43840 0 1 36034
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 1 0 43840 0 1 35948
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 1 0 43840 0 1 35862
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 1 0 43840 0 1 35776
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 1 0 43840 0 1 35690
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 1 0 43840 0 1 35604
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 1 0 43840 0 1 35518
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 1 0 43840 0 1 35432
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 1 0 43840 0 1 35346
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 1 0 43840 0 1 35260
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 1 0 43840 0 1 35174
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 1 0 43840 0 1 35088
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 1 0 43840 0 1 35002
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 1 0 43840 0 1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 1 0 43840 0 1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 1 0 43840 0 1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 1 0 43840 0 1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 1 0 43840 0 1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 1 0 43840 0 1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 1 0 43840 0 1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 1 0 43840 0 1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 1 0 43840 0 1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 1 0 43840 0 1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 1 0 43840 0 1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_887
timestamp 1300117811
transform -1 0 5828 0 -1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_888
timestamp 1300117811
transform -1 0 5828 0 -1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_889
timestamp 1300117811
transform -1 0 5828 0 -1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_890
timestamp 1300117811
transform -1 0 5828 0 -1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_891
timestamp 1300117811
transform -1 0 5828 0 -1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_892
timestamp 1300117811
transform -1 0 5828 0 -1 31906
box 0 0 6450 86
use fillpp_mt fillpp_mt_893
timestamp 1300117811
transform -1 0 5828 0 -1 31820
box 0 0 6450 86
use fillpp_mt fillpp_mt_894
timestamp 1300117811
transform -1 0 5828 0 -1 31734
box 0 0 6450 86
use fillpp_mt fillpp_mt_895
timestamp 1300117811
transform -1 0 5828 0 -1 31648
box 0 0 6450 86
use fillpp_mt fillpp_mt_896
timestamp 1300117811
transform -1 0 5828 0 -1 31562
box 0 0 6450 86
use fillpp_mt fillpp_mt_897
timestamp 1300117811
transform -1 0 5828 0 -1 31476
box 0 0 6450 86
use fillpp_mt fillpp_mt_898
timestamp 1300117811
transform -1 0 5828 0 -1 31390
box 0 0 6450 86
use fillpp_mt fillpp_mt_899
timestamp 1300117811
transform -1 0 5828 0 -1 31304
box 0 0 6450 86
use fillpp_mt fillpp_mt_900
timestamp 1300117811
transform -1 0 5828 0 -1 31218
box 0 0 6450 86
use fillpp_mt fillpp_mt_901
timestamp 1300117811
transform -1 0 5828 0 -1 31132
box 0 0 6450 86
use fillpp_mt fillpp_mt_902
timestamp 1300117811
transform -1 0 5828 0 -1 31046
box 0 0 6450 86
use fillpp_mt fillpp_mt_903
timestamp 1300117811
transform -1 0 5828 0 -1 30960
box 0 0 6450 86
use fillpp_mt fillpp_mt_904
timestamp 1300117811
transform -1 0 5828 0 -1 30874
box 0 0 6450 86
use fillpp_mt fillpp_mt_905
timestamp 1300117811
transform -1 0 5828 0 -1 30788
box 0 0 6450 86
use fillpp_mt fillpp_mt_906
timestamp 1300117811
transform -1 0 5828 0 -1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_907
timestamp 1300117811
transform -1 0 5828 0 -1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_908
timestamp 1300117811
transform -1 0 5828 0 -1 30530
box 0 0 6450 86
use fillpp_mt fillpp_mt_909
timestamp 1300117811
transform -1 0 5828 0 -1 30444
box 0 0 6450 86
use fillpp_mt fillpp_mt_910
timestamp 1300117811
transform -1 0 5828 0 -1 30358
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 43840 0 1 32336
box 0 0 6450 1720
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 1 0 43840 0 1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 1 0 43840 0 1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 1 0 43840 0 1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 1 0 43840 0 1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 1 0 43840 0 1 31906
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 1 0 43840 0 1 31820
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 1 0 43840 0 1 31734
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 1 0 43840 0 1 31648
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 1 0 43840 0 1 31562
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 1 0 43840 0 1 31476
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 1 0 43840 0 1 31390
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 1 0 43840 0 1 31304
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 1 0 43840 0 1 31218
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 1 0 43840 0 1 31132
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 1 0 43840 0 1 31046
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 1 0 43840 0 1 30960
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 1 0 43840 0 1 30874
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 1 0 43840 0 1 30788
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 1 0 43840 0 1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 1 0 43840 0 1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 1 0 43840 0 1 30530
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 1 0 43840 0 1 30444
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 1 0 43840 0 1 30358
box 0 0 6450 86
use fillpp_mt fillpp_mt_911
timestamp 1300117811
transform -1 0 5828 0 -1 30272
box 0 0 6450 86
use fillpp_mt fillpp_mt_912
timestamp 1300117811
transform -1 0 5828 0 -1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_913
timestamp 1300117811
transform -1 0 5828 0 -1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_914
timestamp 1300117811
transform -1 0 5828 0 -1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_915
timestamp 1300117811
transform -1 0 5828 0 -1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_916
timestamp 1300117811
transform -1 0 5828 0 -1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_917
timestamp 1300117811
transform -1 0 5828 0 -1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_918
timestamp 1300117811
transform -1 0 5828 0 -1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_919
timestamp 1300117811
transform -1 0 5828 0 -1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_920
timestamp 1300117811
transform -1 0 5828 0 -1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_921
timestamp 1300117811
transform -1 0 5828 0 -1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_922
timestamp 1300117811
transform -1 0 5828 0 -1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_923
timestamp 1300117811
transform -1 0 5828 0 -1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_924
timestamp 1300117811
transform -1 0 5828 0 -1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_925
timestamp 1300117811
transform -1 0 5828 0 -1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_926
timestamp 1300117811
transform -1 0 5828 0 -1 28982
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 5828 0 -1 28896
box 0 0 6450 1720
use fillpp_mt fillpp_mt_927
timestamp 1300117811
transform -1 0 5828 0 -1 27176
box 0 0 6450 86
use fillpp_mt fillpp_mt_928
timestamp 1300117811
transform -1 0 5828 0 -1 27090
box 0 0 6450 86
use fillpp_mt fillpp_mt_929
timestamp 1300117811
transform -1 0 5828 0 -1 27004
box 0 0 6450 86
use fillpp_mt fillpp_mt_930
timestamp 1300117811
transform -1 0 5828 0 -1 26918
box 0 0 6450 86
use fillpp_mt fillpp_mt_931
timestamp 1300117811
transform -1 0 5828 0 -1 26832
box 0 0 6450 86
use fillpp_mt fillpp_mt_932
timestamp 1300117811
transform -1 0 5828 0 -1 26746
box 0 0 6450 86
use fillpp_mt fillpp_mt_933
timestamp 1300117811
transform -1 0 5828 0 -1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_934
timestamp 1300117811
transform -1 0 5828 0 -1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_935
timestamp 1300117811
transform -1 0 5828 0 -1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_936
timestamp 1300117811
transform -1 0 5828 0 -1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_937
timestamp 1300117811
transform -1 0 5828 0 -1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_938
timestamp 1300117811
transform -1 0 5828 0 -1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_939
timestamp 1300117811
transform -1 0 5828 0 -1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_940
timestamp 1300117811
transform -1 0 5828 0 -1 26058
box 0 0 6450 86
use fillpp_mt fillpp_mt_941
timestamp 1300117811
transform -1 0 5828 0 -1 25972
box 0 0 6450 86
use fillpp_mt fillpp_mt_942
timestamp 1300117811
transform -1 0 5828 0 -1 25886
box 0 0 6450 86
use fillpp_mt fillpp_mt_943
timestamp 1300117811
transform -1 0 5828 0 -1 25800
box 0 0 6450 86
use fillpp_mt fillpp_mt_944
timestamp 1300117811
transform -1 0 5828 0 -1 25714
box 0 0 6450 86
use fillpp_mt fillpp_mt_945
timestamp 1300117811
transform -1 0 5828 0 -1 25628
box 0 0 6450 86
use fillpp_mt fillpp_mt_946
timestamp 1300117811
transform -1 0 5828 0 -1 25542
box 0 0 6450 86
use fillpp_mt fillpp_mt_947
timestamp 1300117811
transform -1 0 5828 0 -1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_948
timestamp 1300117811
transform -1 0 5828 0 -1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_949
timestamp 1300117811
transform -1 0 5828 0 -1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_950
timestamp 1300117811
transform -1 0 5828 0 -1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_951
timestamp 1300117811
transform -1 0 5828 0 -1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_952
timestamp 1300117811
transform -1 0 5828 0 -1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_953
timestamp 1300117811
transform -1 0 5828 0 -1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_954
timestamp 1300117811
transform -1 0 5828 0 -1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_955
timestamp 1300117811
transform -1 0 5828 0 -1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_956
timestamp 1300117811
transform -1 0 5828 0 -1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_957
timestamp 1300117811
transform -1 0 5828 0 -1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_958
timestamp 1300117811
transform -1 0 5828 0 -1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_959
timestamp 1300117811
transform -1 0 5828 0 -1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_960
timestamp 1300117811
transform -1 0 5828 0 -1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_961
timestamp 1300117811
transform -1 0 5828 0 -1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_962
timestamp 1300117811
transform -1 0 5828 0 -1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_963
timestamp 1300117811
transform -1 0 5828 0 -1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_964
timestamp 1300117811
transform -1 0 5828 0 -1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_965
timestamp 1300117811
transform -1 0 5828 0 -1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_966
timestamp 1300117811
transform -1 0 5828 0 -1 23822
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 5828 0 -1 23736
box 0 0 6450 1720
use fillpp_mt fillpp_mt_967
timestamp 1300117811
transform -1 0 5828 0 -1 22016
box 0 0 6450 86
use fillpp_mt fillpp_mt_968
timestamp 1300117811
transform -1 0 5828 0 -1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_969
timestamp 1300117811
transform -1 0 5828 0 -1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_970
timestamp 1300117811
transform -1 0 5828 0 -1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_971
timestamp 1300117811
transform -1 0 5828 0 -1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_972
timestamp 1300117811
transform -1 0 5828 0 -1 21586
box 0 0 6450 86
use fillpp_mt fillpp_mt_973
timestamp 1300117811
transform -1 0 5828 0 -1 21500
box 0 0 6450 86
use fillpp_mt fillpp_mt_974
timestamp 1300117811
transform -1 0 5828 0 -1 21414
box 0 0 6450 86
use fillpp_mt fillpp_mt_975
timestamp 1300117811
transform -1 0 5828 0 -1 21328
box 0 0 6450 86
use fillpp_mt fillpp_mt_976
timestamp 1300117811
transform -1 0 5828 0 -1 21242
box 0 0 6450 86
use fillpp_mt fillpp_mt_977
timestamp 1300117811
transform -1 0 5828 0 -1 21156
box 0 0 6450 86
use fillpp_mt fillpp_mt_978
timestamp 1300117811
transform -1 0 5828 0 -1 21070
box 0 0 6450 86
use fillpp_mt fillpp_mt_979
timestamp 1300117811
transform -1 0 5828 0 -1 20984
box 0 0 6450 86
use fillpp_mt fillpp_mt_980
timestamp 1300117811
transform -1 0 5828 0 -1 20898
box 0 0 6450 86
use fillpp_mt fillpp_mt_981
timestamp 1300117811
transform -1 0 5828 0 -1 20812
box 0 0 6450 86
use fillpp_mt fillpp_mt_982
timestamp 1300117811
transform -1 0 5828 0 -1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_983
timestamp 1300117811
transform -1 0 5828 0 -1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_984
timestamp 1300117811
transform -1 0 5828 0 -1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_985
timestamp 1300117811
transform -1 0 5828 0 -1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_986
timestamp 1300117811
transform -1 0 5828 0 -1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_987
timestamp 1300117811
transform -1 0 5828 0 -1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_988
timestamp 1300117811
transform -1 0 5828 0 -1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_989
timestamp 1300117811
transform -1 0 5828 0 -1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_990
timestamp 1300117811
transform -1 0 5828 0 -1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_991
timestamp 1300117811
transform -1 0 5828 0 -1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_992
timestamp 1300117811
transform -1 0 5828 0 -1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_993
timestamp 1300117811
transform -1 0 5828 0 -1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_994
timestamp 1300117811
transform -1 0 5828 0 -1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_995
timestamp 1300117811
transform -1 0 5828 0 -1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_996
timestamp 1300117811
transform -1 0 5828 0 -1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_997
timestamp 1300117811
transform -1 0 5828 0 -1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_998
timestamp 1300117811
transform -1 0 5828 0 -1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_999
timestamp 1300117811
transform -1 0 5828 0 -1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_1000
timestamp 1300117811
transform -1 0 5828 0 -1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_1001
timestamp 1300117811
transform -1 0 5828 0 -1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_1002
timestamp 1300117811
transform -1 0 5828 0 -1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_1003
timestamp 1300117811
transform -1 0 5828 0 -1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_1004
timestamp 1300117811
transform -1 0 5828 0 -1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_1005
timestamp 1300117811
transform -1 0 5828 0 -1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_1006
timestamp 1300117811
transform -1 0 5828 0 -1 18662
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 5828 0 -1 18576
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1007
timestamp 1300117811
transform -1 0 5828 0 -1 16856
box 0 0 6450 86
use fillpp_mt fillpp_mt_1008
timestamp 1300117811
transform -1 0 5828 0 -1 16770
box 0 0 6450 86
use fillpp_mt fillpp_mt_1009
timestamp 1300117811
transform -1 0 5828 0 -1 16684
box 0 0 6450 86
use fillpp_mt fillpp_mt_1010
timestamp 1300117811
transform -1 0 5828 0 -1 16598
box 0 0 6450 86
use fillpp_mt fillpp_mt_1011
timestamp 1300117811
transform -1 0 5828 0 -1 16512
box 0 0 6450 86
use fillpp_mt fillpp_mt_1012
timestamp 1300117811
transform -1 0 5828 0 -1 16426
box 0 0 6450 86
use fillpp_mt fillpp_mt_1013
timestamp 1300117811
transform -1 0 5828 0 -1 16340
box 0 0 6450 86
use fillpp_mt fillpp_mt_1014
timestamp 1300117811
transform -1 0 5828 0 -1 16254
box 0 0 6450 86
use fillpp_mt fillpp_mt_1015
timestamp 1300117811
transform -1 0 5828 0 -1 16168
box 0 0 6450 86
use fillpp_mt fillpp_mt_1016
timestamp 1300117811
transform -1 0 5828 0 -1 16082
box 0 0 6450 86
use fillpp_mt fillpp_mt_1017
timestamp 1300117811
transform -1 0 5828 0 -1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_1018
timestamp 1300117811
transform -1 0 5828 0 -1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_1019
timestamp 1300117811
transform -1 0 5828 0 -1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_1020
timestamp 1300117811
transform -1 0 5828 0 -1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_1021
timestamp 1300117811
transform -1 0 5828 0 -1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_1022
timestamp 1300117811
transform -1 0 5828 0 -1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_1023
timestamp 1300117811
transform -1 0 5828 0 -1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_1024
timestamp 1300117811
transform -1 0 5828 0 -1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_1025
timestamp 1300117811
transform -1 0 5828 0 -1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_1026
timestamp 1300117811
transform -1 0 5828 0 -1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_1027
timestamp 1300117811
transform -1 0 5828 0 -1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_1028
timestamp 1300117811
transform -1 0 5828 0 -1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_1029
timestamp 1300117811
transform -1 0 5828 0 -1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_1030
timestamp 1300117811
transform -1 0 5828 0 -1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_1031
timestamp 1300117811
transform -1 0 5828 0 -1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_1032
timestamp 1300117811
transform -1 0 5828 0 -1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_1033
timestamp 1300117811
transform -1 0 5828 0 -1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_1034
timestamp 1300117811
transform -1 0 5828 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_1035
timestamp 1300117811
transform -1 0 5828 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_1036
timestamp 1300117811
transform -1 0 5828 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_1037
timestamp 1300117811
transform -1 0 5828 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_1038
timestamp 1300117811
transform -1 0 5828 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_1039
timestamp 1300117811
transform -1 0 5828 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_1040
timestamp 1300117811
transform -1 0 5828 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_1041
timestamp 1300117811
transform -1 0 5828 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_1042
timestamp 1300117811
transform -1 0 5828 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_1043
timestamp 1300117811
transform -1 0 5828 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_1044
timestamp 1300117811
transform -1 0 5828 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_1045
timestamp 1300117811
transform -1 0 5828 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_1046
timestamp 1300117811
transform -1 0 5828 0 -1 13502
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 5828 0 -1 13416
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1047
timestamp 1300117811
transform -1 0 5828 0 -1 11696
box 0 0 6450 86
use fillpp_mt fillpp_mt_1048
timestamp 1300117811
transform -1 0 5828 0 -1 11610
box 0 0 6450 86
use fillpp_mt fillpp_mt_1049
timestamp 1300117811
transform -1 0 5828 0 -1 11524
box 0 0 6450 86
use fillpp_mt fillpp_mt_1050
timestamp 1300117811
transform -1 0 5828 0 -1 11438
box 0 0 6450 86
use fillpp_mt fillpp_mt_1051
timestamp 1300117811
transform -1 0 5828 0 -1 11352
box 0 0 6450 86
use fillpp_mt fillpp_mt_1052
timestamp 1300117811
transform -1 0 5828 0 -1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_1053
timestamp 1300117811
transform -1 0 5828 0 -1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_1054
timestamp 1300117811
transform -1 0 5828 0 -1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_1055
timestamp 1300117811
transform -1 0 5828 0 -1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_1056
timestamp 1300117811
transform -1 0 5828 0 -1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_1057
timestamp 1300117811
transform -1 0 5828 0 -1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_1058
timestamp 1300117811
transform -1 0 5828 0 -1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_1059
timestamp 1300117811
transform -1 0 5828 0 -1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_1060
timestamp 1300117811
transform -1 0 5828 0 -1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_1061
timestamp 1300117811
transform -1 0 5828 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_1062
timestamp 1300117811
transform -1 0 5828 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_1063
timestamp 1300117811
transform -1 0 5828 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_1064
timestamp 1300117811
transform -1 0 5828 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_1065
timestamp 1300117811
transform -1 0 5828 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_1066
timestamp 1300117811
transform -1 0 5828 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_1067
timestamp 1300117811
transform -1 0 5828 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_1068
timestamp 1300117811
transform -1 0 5828 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_1069
timestamp 1300117811
transform -1 0 5828 0 -1 9804
box 0 0 6450 86
use datapath datapath_0
timestamp 1395340701
transform 1 0 12579 0 1 9710
box 414 43 25445 20615
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 1 0 43840 0 1 30272
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 1 0 43840 0 1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 1 0 43840 0 1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 1 0 43840 0 1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 1 0 43840 0 1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 1 0 43840 0 1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 1 0 43840 0 1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 1 0 43840 0 1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 1 0 43840 0 1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 1 0 43840 0 1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 1 0 43840 0 1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 1 0 43840 0 1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 1 0 43840 0 1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 1 0 43840 0 1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 1 0 43840 0 1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 1 0 43840 0 1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 1 0 43840 0 1 28896
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 43840 0 1 27176
box 0 0 6450 1720
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 1 0 43840 0 1 27090
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 1 0 43840 0 1 27004
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 1 0 43840 0 1 26918
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 1 0 43840 0 1 26832
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 1 0 43840 0 1 26746
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 1 0 43840 0 1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 1 0 43840 0 1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 1 0 43840 0 1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 1 0 43840 0 1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 1 0 43840 0 1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 1 0 43840 0 1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 1 0 43840 0 1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 1 0 43840 0 1 26058
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 1 0 43840 0 1 25972
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 1 0 43840 0 1 25886
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 1 0 43840 0 1 25800
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 1 0 43840 0 1 25714
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 1 0 43840 0 1 25628
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 1 0 43840 0 1 25542
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 1 0 43840 0 1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 1 0 43840 0 1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 1 0 43840 0 1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 1 0 43840 0 1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 1 0 43840 0 1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 1 0 43840 0 1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 1 0 43840 0 1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 1 0 43840 0 1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 1 0 43840 0 1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 1 0 43840 0 1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 43840 0 1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 43840 0 1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 43840 0 1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 43840 0 1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 43840 0 1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 43840 0 1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 43840 0 1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 43840 0 1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 43840 0 1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 43840 0 1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 43840 0 1 23736
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 43840 0 1 22016
box 0 0 6450 1720
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 43840 0 1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 43840 0 1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 43840 0 1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 43840 0 1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 43840 0 1 21586
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 43840 0 1 21500
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 43840 0 1 21414
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 43840 0 1 21328
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 43840 0 1 21242
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 43840 0 1 21156
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 43840 0 1 21070
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 43840 0 1 20984
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 43840 0 1 20898
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 43840 0 1 20812
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 43840 0 1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 43840 0 1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 43840 0 1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 43840 0 1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 43840 0 1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 43840 0 1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 43840 0 1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 43840 0 1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 43840 0 1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 43840 0 1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 43840 0 1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 43840 0 1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 43840 0 1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 43840 0 1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 43840 0 1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 43840 0 1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 43840 0 1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 43840 0 1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 43840 0 1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 43840 0 1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 43840 0 1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 43840 0 1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 43840 0 1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 43840 0 1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 43840 0 1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 43840 0 1 18576
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 43840 0 1 16856
box 0 0 6450 1720
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 43840 0 1 16770
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 43840 0 1 16684
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 43840 0 1 16598
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 43840 0 1 16512
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 43840 0 1 16426
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 43840 0 1 16340
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 43840 0 1 16254
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 43840 0 1 16168
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 43840 0 1 16082
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 43840 0 1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 43840 0 1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 43840 0 1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 43840 0 1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 43840 0 1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 43840 0 1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 43840 0 1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 43840 0 1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 43840 0 1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 43840 0 1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 43840 0 1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 43840 0 1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 43840 0 1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 43840 0 1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 43840 0 1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 43840 0 1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 43840 0 1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 43840 0 1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 43840 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 43840 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 43840 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 43840 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 43840 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 43840 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 43840 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 43840 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 43840 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 43840 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 43840 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 43840 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 43840 0 1 13416
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 43840 0 1 11696
box 0 0 6450 1720
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 43840 0 1 11610
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 43840 0 1 11524
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 43840 0 1 11438
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 43840 0 1 11352
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 43840 0 1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 43840 0 1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 43840 0 1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 43840 0 1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 43840 0 1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 43840 0 1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 43840 0 1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 43840 0 1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 43840 0 1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 43840 0 1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 43840 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 43840 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 43840 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 43840 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 43840 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 43840 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 43840 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 43840 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_1070
timestamp 1300117811
transform -1 0 5828 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_1071
timestamp 1300117811
transform -1 0 5828 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_1072
timestamp 1300117811
transform -1 0 5828 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_1073
timestamp 1300117811
transform -1 0 5828 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_1074
timestamp 1300117811
transform -1 0 5828 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_1075
timestamp 1300117811
transform -1 0 5828 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_1076
timestamp 1300117811
transform -1 0 5828 0 -1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_1077
timestamp 1300117811
transform -1 0 5828 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_1078
timestamp 1300117811
transform -1 0 5828 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_1079
timestamp 1300117811
transform -1 0 5828 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_1080
timestamp 1300117811
transform -1 0 5828 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_1081
timestamp 1300117811
transform -1 0 5828 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_1082
timestamp 1300117811
transform -1 0 5828 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_1083
timestamp 1300117811
transform -1 0 5828 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_1084
timestamp 1300117811
transform -1 0 5828 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_1085
timestamp 1300117811
transform -1 0 5828 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_1086
timestamp 1300117811
transform -1 0 5828 0 -1 8342
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 5828 0 -1 8256
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1087
timestamp 1300117811
transform -1 0 5828 0 -1 6536
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 43840 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 43840 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 43840 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 43840 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 43840 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 43840 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 43840 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 43840 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 43840 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 43840 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 43840 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 43840 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 43840 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 43840 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 43840 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 43840 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 43840 0 1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 43840 0 1 8256
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 43840 0 1 6536
box 0 0 6450 1720
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 43840 0 1 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 -622 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 5828 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 5914 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 6000 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6086 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 7806 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 7892 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 7978 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8064 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8150 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8236 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8322 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 8408 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 8494 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 8580 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 8666 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 8752 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 8838 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 8924 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9010 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9096 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9182 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9268 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9354 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 9440 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 9526 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 9612 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 9698 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 9784 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 9870 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 9956 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 10042 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 10128 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 10214 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 10300 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 10386 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 10472 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10558 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12278 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12364 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 12450 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 12536 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 12622 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 12708 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 12794 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 12880 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 12966 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 13052 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 13138 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 13224 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 13310 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 13396 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 13482 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 13568 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 13654 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 13740 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 13826 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 13912 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 13998 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 14084 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 14170 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 14256 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 14342 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 14428 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 14514 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 14600 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 14686 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 14772 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 14858 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 14944 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 15030 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 16750 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 16836 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 16922 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 17008 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 17094 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 17180 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 17266 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 17352 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 17438 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 17524 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 17610 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 17696 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 17782 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 17868 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 17954 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 18040 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 18126 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 18212 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 18298 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 18384 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 18470 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 18556 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 18642 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 18728 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 18814 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 18900 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 18986 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 19072 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 19158 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 19244 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 19330 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 19416 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 19502 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 21222 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 21308 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 21394 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 21480 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 21566 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 21652 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 21738 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 21824 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 21910 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 21996 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 22082 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 22168 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 22254 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 22340 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 22426 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 22512 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 22598 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 22684 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 22770 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 22856 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 22942 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 23028 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 23114 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 23200 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 23286 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 23372 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 23458 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 23544 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 23630 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 23716 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 23802 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 23888 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 23974 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 25694 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 25780 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 25866 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 25952 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 26038 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 26124 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 26210 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 26296 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 26382 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 26468 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 26554 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 26640 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 26726 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 26812 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 26898 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 26984 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 27070 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 27156 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 27242 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 27328 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 27414 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 27500 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 27586 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 27672 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 27758 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 27844 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 27930 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 28016 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 28102 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 28188 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 28274 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 28360 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 28446 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 30166 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 30252 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 30338 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 30424 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 30510 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 30596 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 30682 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 0 1 30768 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 0 1 30854 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 0 1 30940 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 0 1 31026 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 0 1 31112 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 0 1 31198 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 0 1 31284 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 0 1 31370 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 0 1 31456 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 0 1 31542 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 0 1 31628 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 0 1 31714 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 0 1 31800 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 0 1 31886 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 0 1 31972 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 0 1 32058 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 0 1 32144 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 0 1 32230 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 0 1 32316 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 0 1 32402 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 0 1 32488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 0 1 32574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 0 1 32660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 0 1 32746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 0 1 32832 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 32918 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 0 1 34638 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 0 1 34724 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 0 1 34810 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 0 1 34896 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 0 1 34982 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 0 1 35068 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 0 1 35154 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 0 1 35240 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 0 1 35326 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 0 1 35412 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 0 1 35498 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 0 1 35584 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 0 1 35670 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 0 1 35756 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 0 1 35842 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 0 1 35928 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 0 1 36014 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 0 1 36100 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 0 1 36186 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 0 1 36272 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 0 1 36358 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 0 1 36444 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 0 1 36530 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 0 1 36616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 0 1 36702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 0 1 36788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 0 1 36874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 0 1 36960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 0 1 37046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 0 1 37132 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 0 1 37218 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 0 1 37304 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 37390 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 0 1 39110 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 0 1 39196 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 0 1 39282 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 0 1 39368 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 0 1 39454 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 0 1 39540 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 0 1 39626 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 0 1 39712 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 0 1 39798 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 0 1 39884 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 0 1 39970 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 0 1 40056 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 0 1 40142 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 0 1 40228 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 0 1 40314 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 0 1 40400 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 0 1 40486 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 0 1 40572 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 0 1 40658 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 0 1 40744 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 0 1 40830 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 0 1 40916 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 0 1 41002 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 0 1 41088 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 0 1 41174 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 0 1 41260 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 0 1 41346 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 0 1 41432 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 0 1 41518 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 0 1 41604 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 0 1 41690 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 0 1 41776 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 41862 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 0 1 43582 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 0 1 43668 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 0 1 43754 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 50290 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 -544 6616 1016 8176 0 nReset
rlabel metal4 -544 11776 1016 13336 0 Clock
rlabel metal4 -544 16936 1016 18496 0 Test
rlabel metal4 -544 22096 1016 23656 0 SDI
rlabel metal4 -544 27256 1016 28816 0 Vdd!
rlabel metal4 -544 32416 1016 33976 0 SDO
rlabel metal4 -544 37576 1016 39136 0 RnW
rlabel metal4 -544 42736 1016 44296 0 nOE
rlabel metal4 6166 49274 7726 50834 0 nWait
rlabel metal4 10638 49274 12198 50834 0 nME
rlabel metal4 15110 49274 16670 50834 0 ALE
rlabel metal4 19582 49274 21142 50834 0 Data[15]
rlabel metal4 24054 49274 25614 50834 0 gnde!
rlabel metal4 28526 49274 30086 50834 0 Data[14]
rlabel metal4 32998 49274 34558 50834 0 Data[13]
rlabel metal4 37470 49274 39030 50834 0 Data[12]
rlabel metal4 41942 49274 43502 50834 0 vdde!
rlabel metal4 48652 42736 50212 44296 0 Data[11]
rlabel metal4 48652 37576 50212 39136 0 Data[10]
rlabel metal4 48652 32416 50212 33976 0 Data[9]
rlabel metal4 48652 27256 50212 28816 0 GND!
rlabel metal4 48652 22096 50212 23656 0 gnde!
rlabel metal4 48652 16936 50212 18496 0 Data[8]
rlabel metal4 48652 11776 50212 13336 0 Data[7]
rlabel metal4 48652 6616 50212 8176 0 Data[6]
rlabel metal4 41942 78 43502 1638 0 gnde!
rlabel metal4 37470 78 39030 1638 0 Data[5]
rlabel metal4 32998 78 34558 1638 0 Data[4]
rlabel metal4 28526 78 30086 1638 0 Data[3]
rlabel metal4 24054 78 25614 1638 0 vdde!
rlabel metal4 19582 78 21142 1638 0 Data[2]
rlabel metal4 15110 78 16670 1638 0 Data[1]
rlabel metal4 10638 78 12198 1638 0 Data[0]
rlabel metal4 6166 78 7726 1638 0 nIRQ
<< end >>
