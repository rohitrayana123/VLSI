../../../Design/Implementation/verilog/behavioural/trisreg.sv