magic
tech c035u
timestamp 1394541067
<< metal1 >>
rect 6911 16721 6945 16731
rect 6959 16721 6993 16731
rect 7007 16721 7041 16731
rect 7055 16721 7089 16731
rect 7103 16721 7137 16731
rect 7151 16721 7185 16731
rect 7199 16721 7233 16731
rect 7247 16721 7545 16731
rect 7559 16721 7593 16731
rect 7607 16721 7641 16731
rect 7655 16721 7689 16731
rect 7703 16721 8001 16731
rect 8015 16721 8049 16731
rect 8063 16721 8361 16731
rect 1345 16573 1427 16574
rect 0 16564 1474 16573
rect 0 16563 1355 16564
rect 1417 16563 1474 16564
rect 1345 16551 1427 16552
rect 0 16542 1474 16551
rect 0 16541 1355 16542
rect 1417 16541 1474 16542
rect 9178 15722 9509 15732
rect 1342 15531 1426 15532
rect 0 15522 1474 15531
rect 0 15521 1352 15522
rect 1416 15521 1474 15522
rect 1342 15509 1426 15510
rect 0 15500 1474 15509
rect 0 15499 1352 15500
rect 1416 15499 1474 15500
rect 9178 14680 9509 14690
rect 1343 14489 1425 14490
rect 0 14480 1474 14489
rect 0 14479 1353 14480
rect 1415 14479 1474 14480
rect 1343 14467 1425 14468
rect 0 14458 1474 14467
rect 0 14457 1353 14458
rect 1415 14457 1474 14458
rect 9178 13638 9509 13648
rect 1346 13447 1428 13448
rect 0 13438 1474 13447
rect 0 13437 1356 13438
rect 1418 13437 1474 13438
rect 1346 13425 1428 13426
rect 0 13416 1474 13425
rect 0 13415 1356 13416
rect 1418 13415 1474 13416
rect 9178 12596 9509 12606
rect 1345 12405 1425 12406
rect 0 12396 1474 12405
rect 0 12395 1355 12396
rect 1415 12395 1474 12396
rect 1345 12383 1425 12384
rect 0 12374 1474 12383
rect 0 12373 1355 12374
rect 1415 12373 1474 12374
rect 9178 11554 9509 11564
rect 1345 11363 1425 11364
rect 0 11354 1474 11363
rect 0 11353 1355 11354
rect 1415 11353 1474 11354
rect 1345 11341 1425 11342
rect 0 11332 1474 11341
rect 0 11331 1355 11332
rect 1415 11331 1474 11332
rect 9178 10512 9509 10522
rect 1344 10321 1428 10322
rect 0 10312 1474 10321
rect 0 10311 1354 10312
rect 1418 10311 1474 10312
rect 1344 10299 1428 10300
rect 0 10290 1474 10299
rect 0 10289 1354 10290
rect 1418 10289 1474 10290
rect 9178 9470 9509 9480
rect 1344 9279 1426 9280
rect 0 9270 1474 9279
rect 0 9269 1354 9270
rect 1416 9269 1474 9270
rect 1344 9257 1426 9258
rect 0 9248 1474 9257
rect 0 9247 1354 9248
rect 1416 9247 1474 9248
rect 9178 8428 9509 8438
rect 1345 8237 1430 8238
rect 0 8228 1474 8237
rect 0 8227 1355 8228
rect 1420 8227 1474 8228
rect 1345 8215 1430 8216
rect 0 8206 1474 8215
rect 0 8205 1355 8206
rect 1420 8205 1474 8206
rect 9178 7386 9509 7396
rect 1344 7195 1428 7196
rect 0 7186 1474 7195
rect 0 7185 1354 7186
rect 1418 7185 1474 7186
rect 1344 7173 1428 7174
rect 0 7164 1474 7173
rect 0 7163 1354 7164
rect 1418 7163 1474 7164
rect 9178 6344 9509 6354
rect 1345 6153 1437 6154
rect 0 6144 1474 6153
rect 0 6143 1355 6144
rect 1427 6143 1474 6144
rect 1345 6131 1437 6132
rect 0 6122 1474 6131
rect 0 6121 1355 6122
rect 1427 6121 1474 6122
rect 9178 5302 9509 5312
rect 1339 5111 1424 5112
rect 0 5102 1474 5111
rect 0 5101 1349 5102
rect 1414 5101 1474 5102
rect 1339 5089 1425 5090
rect 0 5080 1474 5089
rect 0 5079 1349 5080
rect 1415 5079 1474 5080
rect 9178 4260 9509 4270
rect 1344 4069 1426 4070
rect 0 4060 1474 4069
rect 0 4059 1354 4060
rect 1416 4059 1474 4060
rect 1344 4047 1426 4048
rect 0 4038 1474 4047
rect 0 4037 1354 4038
rect 1416 4037 1474 4038
rect 9178 3218 9509 3228
rect 1346 3027 1426 3028
rect 0 3018 1474 3027
rect 0 3017 1356 3018
rect 1416 3017 1474 3018
rect 1346 3005 1426 3006
rect 0 2996 1474 3005
rect 0 2995 1356 2996
rect 1416 2995 1474 2996
rect 9178 2176 9509 2186
rect 1346 1985 1426 1986
rect 0 1976 1474 1985
rect 0 1975 1356 1976
rect 1416 1975 1474 1976
rect 1346 1963 1426 1964
rect 0 1954 1474 1963
rect 0 1953 1356 1954
rect 1416 1953 1474 1954
rect 9178 1134 9509 1144
rect 1346 943 1430 944
rect 0 934 1474 943
rect 0 933 1356 934
rect 1420 933 1474 934
rect 1346 921 1430 922
rect 0 912 1474 921
rect 0 911 1356 912
rect 1420 911 1474 912
rect 9178 92 9509 102
rect 1511 24 2457 34
rect 2471 24 5121 34
rect 5135 24 5169 34
rect 5183 24 5217 34
rect 5231 24 5265 34
rect 5279 24 5313 34
rect 5327 24 5361 34
rect 5375 24 5409 34
rect 5423 24 5457 34
rect 5471 24 5769 34
rect 5783 24 5817 34
rect 5831 24 5865 34
rect 5879 24 5913 34
rect 5927 24 6225 34
rect 6239 24 6273 34
rect 6287 24 6657 34
rect 1991 2 2169 12
<< m2contact >>
rect 6897 16719 6911 16733
rect 6945 16719 6959 16733
rect 6993 16719 7007 16733
rect 7041 16719 7055 16733
rect 7089 16719 7103 16733
rect 7137 16719 7151 16733
rect 7185 16719 7199 16733
rect 7233 16719 7247 16733
rect 7545 16719 7559 16733
rect 7593 16719 7607 16733
rect 7641 16719 7655 16733
rect 7689 16719 7703 16733
rect 8001 16719 8015 16733
rect 8049 16719 8063 16733
rect 8361 16719 8375 16733
rect 1497 22 1511 36
rect 2457 22 2471 36
rect 5121 22 5135 36
rect 5169 22 5183 36
rect 5217 22 5231 36
rect 5265 22 5279 36
rect 5313 22 5327 36
rect 5361 22 5375 36
rect 5409 22 5423 36
rect 5457 22 5471 36
rect 5769 22 5783 36
rect 5817 22 5831 36
rect 5865 22 5879 36
rect 5913 22 5927 36
rect 6225 22 6239 36
rect 6273 22 6287 36
rect 6657 22 6671 36
rect 1977 0 1991 14
rect 2169 0 2183 14
<< metal2 >>
rect 10 16536 210 16785
rect 226 16536 238 16785
rect 250 16536 262 16785
rect 274 16536 286 16785
rect 298 16536 310 16785
rect 1546 16713 1558 16785
rect 1810 16713 1822 16785
rect 1978 16713 1990 16785
rect 2146 16713 2158 16785
rect 2170 16713 2182 16785
rect 2242 16713 2254 16785
rect 2458 16713 2470 16785
rect 2602 16713 2614 16785
rect 2938 16713 2950 16785
rect 3298 16713 3310 16785
rect 3706 16713 3718 16785
rect 4042 16713 4054 16785
rect 4354 16713 4366 16785
rect 4690 16713 4702 16785
rect 4810 16713 4822 16785
rect 4858 16713 4870 16785
rect 5026 16713 5038 16785
rect 6826 16713 6838 16785
rect 6851 16713 6863 16785
rect 6898 16713 6910 16719
rect 6946 16713 6958 16719
rect 6994 16713 7006 16719
rect 7042 16713 7054 16719
rect 7090 16713 7102 16719
rect 7138 16713 7150 16719
rect 7186 16713 7198 16719
rect 7234 16713 7246 16719
rect 7474 16713 7486 16785
rect 7690 16733 7702 16785
rect 7546 16713 7558 16719
rect 7594 16713 7606 16719
rect 7642 16713 7654 16719
rect 7690 16713 7702 16719
rect 7930 16713 7942 16785
rect 8002 16713 8014 16719
rect 8050 16713 8062 16719
rect 8290 16713 8302 16785
rect 8362 16713 8374 16719
rect 8650 16713 8662 16785
rect 8818 16713 8830 16785
rect 9058 16713 9070 16785
rect 9298 16536 9498 16785
rect 10 15494 210 15737
rect 226 15494 238 15737
rect 250 15494 262 15737
rect 274 15494 286 15737
rect 298 15494 310 15737
rect 9298 15494 9498 15737
rect 10 14452 210 14695
rect 226 14452 238 14695
rect 250 14452 262 14695
rect 274 14452 286 14695
rect 298 14452 310 14695
rect 9298 14452 9498 14695
rect 10 13410 210 13653
rect 226 13410 238 13653
rect 250 13410 262 13653
rect 274 13410 286 13653
rect 298 13410 310 13653
rect 9298 13410 9498 13653
rect 10 12368 210 12611
rect 226 12368 238 12611
rect 250 12368 262 12611
rect 274 12368 286 12611
rect 298 12368 310 12611
rect 9298 12368 9498 12611
rect 10 11326 210 11569
rect 226 11326 238 11569
rect 250 11326 262 11569
rect 274 11326 286 11569
rect 298 11326 310 11569
rect 9298 11326 9498 11569
rect 10 10284 210 10527
rect 226 10284 238 10527
rect 250 10284 262 10527
rect 274 10284 286 10527
rect 298 10284 310 10527
rect 9298 10284 9498 10527
rect 10 9242 210 9485
rect 226 9242 238 9485
rect 250 9242 262 9485
rect 274 9242 286 9485
rect 298 9242 310 9485
rect 9298 9242 9498 9485
rect 10 8200 210 8443
rect 226 8200 238 8443
rect 250 8200 262 8443
rect 274 8200 286 8443
rect 298 8200 310 8443
rect 9298 8200 9498 8443
rect 10 7158 210 7401
rect 226 7158 238 7401
rect 250 7158 262 7401
rect 274 7158 286 7401
rect 298 7158 310 7401
rect 9298 7158 9498 7401
rect 10 6116 210 6359
rect 226 6116 238 6359
rect 250 6116 262 6359
rect 274 6116 286 6359
rect 298 6116 310 6359
rect 9298 6116 9498 6359
rect 10 5074 210 5317
rect 226 5074 238 5317
rect 250 5074 262 5317
rect 274 5074 286 5317
rect 298 5074 310 5317
rect 9298 5074 9498 5317
rect 10 4032 210 4275
rect 226 4032 238 4275
rect 250 4032 262 4275
rect 274 4032 286 4275
rect 298 4032 310 4275
rect 9298 4032 9498 4275
rect 10 2990 210 3233
rect 226 2990 238 3233
rect 250 2990 262 3233
rect 274 2990 286 3233
rect 298 2990 310 3233
rect 9298 2990 9498 3233
rect 10 1948 210 2191
rect 226 1948 238 2191
rect 250 1948 262 2191
rect 274 1948 286 2191
rect 298 1948 310 2191
rect 9298 1948 9498 2191
rect 10 906 210 1149
rect 226 906 238 1149
rect 250 906 262 1149
rect 274 906 286 1149
rect 298 906 310 1149
rect 9298 906 9498 1149
rect 1498 36 1510 41
rect 1978 14 1990 41
rect 2170 14 2182 41
rect 2458 36 2470 41
rect 5122 36 5134 41
rect 5170 36 5182 41
rect 5218 36 5230 41
rect 5266 36 5278 41
rect 5314 36 5326 41
rect 5362 36 5374 41
rect 5410 36 5422 41
rect 5458 36 5470 41
rect 5770 36 5782 41
rect 5818 36 5830 41
rect 5866 36 5878 41
rect 5914 36 5926 41
rect 6226 36 6238 41
rect 6274 36 6286 41
rect 6658 36 6670 41
use leftbuf leftbuf_15
timestamp 1386242881
transform 1 0 10 0 1 15737
box 0 0 1464 799
use LLIcell_U LLIcell_U_7
timestamp 1393855556
transform 1 0 8770 0 1 15671
box 0 0 192 1042
use ALUSlice ALUSlice_15
timestamp 1394540006
transform 1 0 1474 0 1 15671
box 0 0 7704 1042
use rightend rightend_15
timestamp 1386235834
transform 1 0 9178 0 1 15737
box 0 0 320 799
use leftbuf leftbuf_14
timestamp 1386242881
transform 1 0 10 0 1 14695
box 0 0 1464 799
use LLIcell_U LLIcell_U_6
timestamp 1393855556
transform 1 0 8770 0 1 14629
box 0 0 192 1042
use ALUSlice ALUSlice_14
timestamp 1394540006
transform 1 0 1474 0 1 14629
box 0 0 7704 1042
use rightend rightend_14
timestamp 1386235834
transform 1 0 9178 0 1 14695
box 0 0 320 799
use leftbuf leftbuf_13
timestamp 1386242881
transform 1 0 10 0 1 13653
box 0 0 1464 799
use LLIcell_U LLIcell_U_5
timestamp 1393855556
transform 1 0 8770 0 1 13587
box 0 0 192 1042
use ALUSlice ALUSlice_13
timestamp 1394540006
transform 1 0 1474 0 1 13587
box 0 0 7704 1042
use rightend rightend_13
timestamp 1386235834
transform 1 0 9178 0 1 13653
box 0 0 320 799
use leftbuf leftbuf_12
timestamp 1386242881
transform 1 0 10 0 1 12611
box 0 0 1464 799
use LLIcell_U LLIcell_U_4
timestamp 1393855556
transform 1 0 8770 0 1 12545
box 0 0 192 1042
use ALUSlice ALUSlice_12
timestamp 1394540006
transform 1 0 1474 0 1 12545
box 0 0 7704 1042
use rightend rightend_12
timestamp 1386235834
transform 1 0 9178 0 1 12611
box 0 0 320 799
use leftbuf leftbuf_11
timestamp 1386242881
transform 1 0 10 0 1 11569
box 0 0 1464 799
use LLIcell_U LLIcell_U_3
timestamp 1393855556
transform 1 0 8770 0 1 11503
box 0 0 192 1042
use ALUSlice ALUSlice_11
timestamp 1394540006
transform 1 0 1474 0 1 11503
box 0 0 7704 1042
use rightend rightend_11
timestamp 1386235834
transform 1 0 9178 0 1 11569
box 0 0 320 799
use leftbuf leftbuf_10
timestamp 1386242881
transform 1 0 10 0 1 10527
box 0 0 1464 799
use LLIcell_U LLIcell_U_2
timestamp 1393855556
transform 1 0 8770 0 1 10461
box 0 0 192 1042
use ALUSlice ALUSlice_10
timestamp 1394540006
transform 1 0 1474 0 1 10461
box 0 0 7704 1042
use rightend rightend_10
timestamp 1386235834
transform 1 0 9178 0 1 10527
box 0 0 320 799
use leftbuf leftbuf_9
timestamp 1386242881
transform 1 0 10 0 1 9485
box 0 0 1464 799
use LLIcell_U LLIcell_U_1
timestamp 1393855556
transform 1 0 8770 0 1 9419
box 0 0 192 1042
use ALUSlice ALUSlice_9
timestamp 1394540006
transform 1 0 1474 0 1 9419
box 0 0 7704 1042
use rightend rightend_9
timestamp 1386235834
transform 1 0 9178 0 1 9485
box 0 0 320 799
use leftbuf leftbuf_8
timestamp 1386242881
transform 1 0 10 0 1 8443
box 0 0 1464 799
use LLIcell_U LLIcell_U_0
timestamp 1393855556
transform 1 0 8770 0 1 8377
box 0 0 192 1042
use ALUSlice ALUSlice_8
timestamp 1394540006
transform 1 0 1474 0 1 8377
box 0 0 7704 1042
use rightend rightend_8
timestamp 1386235834
transform 1 0 9178 0 1 8443
box 0 0 320 799
use leftbuf leftbuf_7
timestamp 1386242881
transform 1 0 10 0 1 7401
box 0 0 1464 799
use LLIcell_L LLIcell_L_3
timestamp 1394447900
transform 1 0 8770 0 1 7335
box 0 0 192 1042
use ALUSlice ALUSlice_7
timestamp 1394540006
transform 1 0 1474 0 1 7335
box 0 0 7704 1042
use rightend rightend_7
timestamp 1386235834
transform 1 0 9178 0 1 7401
box 0 0 320 799
use leftbuf leftbuf_6
timestamp 1386242881
transform 1 0 10 0 1 6359
box 0 0 1464 799
use LLIcell_L LLIcell_L_7
timestamp 1394447900
transform 1 0 8770 0 1 6293
box 0 0 192 1042
use ALUSlice ALUSlice_6
timestamp 1394540006
transform 1 0 1474 0 1 6293
box 0 0 7704 1042
use rightend rightend_6
timestamp 1386235834
transform 1 0 9178 0 1 6359
box 0 0 320 799
use leftbuf leftbuf_5
timestamp 1386242881
transform 1 0 10 0 1 5317
box 0 0 1464 799
use LLIcell_L LLIcell_L_6
timestamp 1394447900
transform 1 0 8770 0 1 5251
box 0 0 192 1042
use ALUSlice ALUSlice_5
timestamp 1394540006
transform 1 0 1474 0 1 5251
box 0 0 7704 1042
use rightend rightend_5
timestamp 1386235834
transform 1 0 9178 0 1 5317
box 0 0 320 799
use leftbuf leftbuf_4
timestamp 1386242881
transform 1 0 10 0 1 4275
box 0 0 1464 799
use LLIcell_L LLIcell_L_5
timestamp 1394447900
transform 1 0 8770 0 1 4209
box 0 0 192 1042
use ALUSlice ALUSlice_4
timestamp 1394540006
transform 1 0 1474 0 1 4209
box 0 0 7704 1042
use rightend rightend_4
timestamp 1386235834
transform 1 0 9178 0 1 4275
box 0 0 320 799
use leftbuf leftbuf_3
timestamp 1386242881
transform 1 0 10 0 1 3233
box 0 0 1464 799
use LLIcell_L LLIcell_L_4
timestamp 1394447900
transform 1 0 8770 0 1 3167
box 0 0 192 1042
use ALUSlice ALUSlice_3
timestamp 1394540006
transform 1 0 1474 0 1 3167
box 0 0 7704 1042
use rightend rightend_3
timestamp 1386235834
transform 1 0 9178 0 1 3233
box 0 0 320 799
use leftbuf leftbuf_2
timestamp 1386242881
transform 1 0 10 0 1 2191
box 0 0 1464 799
use LLIcell_L LLIcell_L_2
timestamp 1394447900
transform 1 0 8770 0 1 2125
box 0 0 192 1042
use ALUSlice ALUSlice_2
timestamp 1394540006
transform 1 0 1474 0 1 2125
box 0 0 7704 1042
use rightend rightend_2
timestamp 1386235834
transform 1 0 9178 0 1 2191
box 0 0 320 799
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 10 0 1 1149
box 0 0 1464 799
use LLIcell_L LLIcell_L_1
timestamp 1394447900
transform 1 0 8770 0 1 1083
box 0 0 192 1042
use ALUSlice ALUSlice_1
timestamp 1394540006
transform 1 0 1474 0 1 1083
box 0 0 7704 1042
use rightend rightend_1
timestamp 1386235834
transform 1 0 9178 0 1 1149
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 10 0 1 107
box 0 0 1464 799
use LLIcell_L LLIcell_L_0
timestamp 1394447900
transform 1 0 8770 0 1 41
box 0 0 192 1042
use ALUSlice ALUSlice_0
timestamp 1394540006
transform 1 0 1474 0 1 41
box 0 0 7704 1042
use rightend rightend_0
timestamp 1386235834
transform 1 0 9178 0 1 107
box 0 0 320 799
<< labels >>
rlabel metal2 1978 16785 1990 16785 5 CIn
rlabel metal2 2242 16785 2254 16785 5 Sum
rlabel metal2 2170 16785 2182 16785 5 COut
rlabel metal2 4858 16785 4870 16785 5 ShB
rlabel metal2 4690 16785 4702 16785 5 NOR
rlabel metal2 4354 16785 4366 16785 5 NAND
rlabel metal2 4042 16785 4054 16785 5 NOT
rlabel metal2 3706 16785 3718 16785 5 XOR
rlabel metal2 3298 16785 3310 16785 5 OR
rlabel metal2 2938 16785 2950 16785 5 AND
rlabel metal2 1810 16785 1822 16785 5 SUB
rlabel metal2 2458 16785 2470 16785 5 nZ
rlabel metal2 2602 16785 2614 16785 5 FAOut
rlabel metal2 5026 16785 5038 16785 5 ShL
rlabel metal2 2146 16785 2158 16785 5 CIn_Slice
rlabel metal2 4810 16785 4822 16785 5 Sign
rlabel metal2 1546 16785 1558 16785 5 ZeroA
rlabel metal2 10 16785 210 16785 5 Vdd!
rlabel metal2 226 16785 238 16785 5 SDO
rlabel metal2 250 16785 262 16785 5 Test
rlabel metal2 274 16785 286 16785 5 Clock
rlabel metal2 298 16785 310 16785 5 nReset
rlabel metal1 0 911 0 921 3 A[0]
rlabel metal1 0 933 0 943 3 B[0]
rlabel metal1 0 1953 0 1963 3 A[1]
rlabel metal1 0 1975 0 1984 3 B[1]
rlabel metal1 0 2995 0 3005 3 A[2]
rlabel metal1 0 3017 0 3027 3 B[2]
rlabel metal1 0 4059 0 4069 3 B[3]
rlabel metal1 0 4037 0 4047 3 A[3]
rlabel metal1 0 5101 0 5111 3 B[4]
rlabel metal1 0 5079 0 5089 3 A[4]
rlabel metal1 0 6121 0 6131 3 A[5]
rlabel metal1 0 6143 0 6153 3 B[5]
rlabel metal1 0 7185 0 7195 3 B[6]
rlabel metal1 0 7163 0 7173 3 A[6]
rlabel metal1 0 8227 0 8237 3 B[7]
rlabel metal1 0 8205 0 8215 3 A[7]
rlabel metal1 0 9269 0 9279 3 B[8]
rlabel metal1 0 9247 0 9257 3 A[8]
rlabel metal1 0 10311 0 10321 3 B[9]
rlabel metal1 0 10289 0 10299 3 A[9]
rlabel metal1 0 11353 0 11363 3 B[10]
rlabel metal1 0 11331 0 11341 3 A[10]
rlabel metal1 0 12395 0 12405 3 B[11]
rlabel metal1 0 12373 0 12383 3 A[11]
rlabel metal1 0 13415 0 13425 3 A[12]
rlabel metal1 0 13437 0 13447 3 B[12]
rlabel metal1 0 14457 0 14467 3 A[13]
rlabel metal1 0 14479 0 14489 3 B[13]
rlabel metal1 0 15521 0 15531 3 B[14]
rlabel metal1 0 15499 0 15509 3 A[14]
rlabel metal1 0 16563 0 16573 3 B[15]
rlabel metal1 0 16541 0 16551 3 A[15]
rlabel metal1 9509 15722 9509 15732 7 ALUOut[15]
rlabel metal1 9509 14680 9509 14690 7 ALUOut[14]
rlabel metal1 9509 13638 9509 13648 7 ALUOut[13]
rlabel metal1 9509 12596 9509 12606 7 ALUOut[12]
rlabel metal1 9509 11554 9509 11564 7 ALUOut[11]
rlabel metal1 9509 10512 9509 10522 7 ALUOut[10]
rlabel metal1 9509 6344 9509 6354 7 ALUOut[6]
rlabel metal1 9509 5302 9509 5312 7 ALUOut[5]
rlabel metal1 9509 4260 9509 4270 7 ALUOut[4]
rlabel metal1 9509 3218 9509 3228 7 ALUOut[3]
rlabel metal1 9509 2176 9509 2186 7 ALUOut[2]
rlabel metal1 9509 1134 9509 1144 7 ALUOut[1]
rlabel metal1 9509 92 9509 102 7 ALUOut[0]
rlabel metal2 9298 16785 9498 16785 5 GND!
rlabel metal2 9058 16785 9070 16785 5 ALUEnable
rlabel metal2 8818 16785 8830 16785 5 LLI
rlabel metal2 8650 16785 8662 16785 5 ShOut
rlabel metal2 7930 16785 7942 16785 5 Sh2
rlabel metal2 8290 16785 8302 16785 5 Sh1
rlabel metal2 7690 16785 7702 16785 5 ShSignIn
rlabel metal2 7474 16785 7486 16785 5 Sh4
rlabel metal2 6826 16785 6838 16785 5 Sh8
rlabel metal2 6851 16785 6863 16785 5 ShR
rlabel metal1 9509 7386 9509 7396 7 ALUOut[7]
rlabel metal1 9509 8428 9509 8438 7 ALUOut[8]
rlabel metal1 9509 9470 9509 9480 7 ALUOut[9]
<< end >>
