magic
tech c035u
timestamp 1395705526
<< pwell >>
rect 26955 1238 27435 1263
<< metal1 >>
rect 15952 8276 15970 8290
rect 18796 8278 18914 8288
rect 15616 8254 20510 8264
rect 14824 8230 17102 8240
rect 18688 8230 27434 8240
rect 14680 8206 25622 8216
rect 9952 8180 9970 8194
rect 11944 8182 27242 8192
rect 5992 8156 6010 8170
rect 6976 8156 6994 8170
rect 9832 8158 21362 8168
rect 4096 8134 7646 8144
rect 9352 8134 27050 8144
rect 27316 8134 27410 8144
rect 2224 8110 4190 8120
rect 4744 8110 5054 8120
rect 5536 8110 27482 8120
rect 1720 8086 2462 8096
rect 2968 8086 12830 8096
rect 12928 8086 23918 8096
rect 24568 8086 27530 8096
rect 84 8062 26114 8072
rect 84 8038 11066 8048
rect 11656 8038 22214 8048
rect 22360 8038 23066 8048
rect 27520 8038 27853 8048
rect 2152 8014 13634 8024
rect 13648 8014 18806 8024
rect 19624 8014 27458 8024
rect 27496 8014 27853 8024
rect 2440 7990 6578 8000
rect 6688 7990 24770 8000
rect 27472 7990 27853 8000
rect 4168 7966 6986 7976
rect 8488 7966 10238 7976
rect 12808 7966 14138 7976
rect 14536 7966 19250 7976
rect 20224 7964 20242 7978
rect 27448 7966 27853 7976
rect 15388 7942 16370 7952
rect 16888 7940 16906 7954
rect 18112 7942 27506 7952
rect 27544 7942 27853 7952
rect 13696 7109 13802 7119
rect 14680 7109 14714 7119
rect 13528 7085 17138 7095
rect 13384 7061 15722 7071
rect 16480 7061 26378 7071
rect 13336 7037 13658 7047
rect 14632 7037 25538 7047
rect 12880 7013 13706 7023
rect 13720 7013 18098 7023
rect 12832 6989 12866 6999
rect 13000 6989 26426 6999
rect 12640 6965 22730 6975
rect 25576 6965 25778 6975
rect 12112 6941 12170 6951
rect 12592 6941 17954 6951
rect 17968 6941 25562 6951
rect 11968 6917 15986 6927
rect 16288 6917 19778 6927
rect 11176 6893 19538 6903
rect 19720 6893 25706 6903
rect 10840 6869 15002 6879
rect 15016 6869 19706 6879
rect 10696 6845 14114 6855
rect 14128 6845 24698 6855
rect 10384 6821 23306 6831
rect 10336 6797 23138 6807
rect 10144 6773 16658 6783
rect 17584 6773 17594 6783
rect 9784 6749 27434 6759
rect 9352 6725 27146 6735
rect 9328 6701 21698 6711
rect 8344 6677 9770 6687
rect 10048 6677 18578 6687
rect 18592 6677 26042 6687
rect 8344 6653 8474 6663
rect 8560 6653 11690 6663
rect 11704 6653 21602 6663
rect 8296 6629 13946 6639
rect 13960 6629 24482 6639
rect 8248 6605 21410 6615
rect 8224 6581 21362 6591
rect 8152 6557 8378 6567
rect 8440 6557 24986 6567
rect 7768 6533 9914 6543
rect 9928 6533 10850 6543
rect 10864 6533 20042 6543
rect 7696 6509 18722 6519
rect 18736 6509 26570 6519
rect 7672 6485 12290 6495
rect 12304 6485 27362 6495
rect 7576 6461 25850 6471
rect 7528 6437 9698 6447
rect 9712 6437 12530 6447
rect 12544 6437 15434 6447
rect 15712 6437 23618 6447
rect 7528 6413 22754 6423
rect 7480 6389 20258 6399
rect 7432 6365 23210 6375
rect 23224 6365 24494 6375
rect 7384 6341 9362 6351
rect 9880 6341 15578 6351
rect 15592 6341 20906 6351
rect 20920 6341 24602 6351
rect 7336 6317 7922 6327
rect 8056 6317 8666 6327
rect 8896 6317 19298 6327
rect 7312 6293 17570 6303
rect 7096 6269 11498 6279
rect 11512 6269 17642 6279
rect 17656 6269 19322 6279
rect 19336 6269 21578 6279
rect 21592 6269 22418 6279
rect 7072 6245 21146 6255
rect 7024 6221 11258 6231
rect 11392 6221 11954 6231
rect 12064 6221 12074 6231
rect 12160 6221 12314 6231
rect 12328 6221 17042 6231
rect 17056 6221 24410 6231
rect 6928 6197 14018 6207
rect 14032 6197 27194 6207
rect 6880 6173 10226 6183
rect 10240 6173 14906 6183
rect 14920 6173 20522 6183
rect 23104 6173 23366 6183
rect 23488 6173 25946 6183
rect 6880 6149 15674 6159
rect 16048 6149 23474 6159
rect 6832 6125 12434 6135
rect 12568 6125 12650 6135
rect 12736 6125 23090 6135
rect 23104 6125 24842 6135
rect 6784 6101 7034 6111
rect 7048 6101 19418 6111
rect 6712 6077 25082 6087
rect 6664 6053 7130 6063
rect 7144 6053 8498 6063
rect 8512 6053 10442 6063
rect 10456 6053 13682 6063
rect 14272 6053 16898 6063
rect 6616 6029 22802 6039
rect 6592 6005 6698 6015
rect 6760 6005 15650 6015
rect 15664 6005 19178 6015
rect 19192 6005 22658 6015
rect 22672 6005 25634 6015
rect 6568 5981 10466 5991
rect 10480 5981 20018 5991
rect 20032 5981 22346 5991
rect 6424 5957 8882 5967
rect 8896 5957 19370 5967
rect 6376 5933 10538 5943
rect 10600 5933 10802 5943
rect 10912 5933 15266 5943
rect 15280 5933 23162 5943
rect 6352 5909 7946 5919
rect 7960 5909 12026 5919
rect 12040 5909 13754 5919
rect 13768 5909 13970 5919
rect 13984 5909 17210 5919
rect 17224 5909 21338 5919
rect 21352 5909 26306 5919
rect 26320 5909 26954 5919
rect 6328 5885 6338 5895
rect 6352 5885 12122 5895
rect 12136 5885 14378 5895
rect 14392 5885 15458 5895
rect 15472 5885 16682 5895
rect 16696 5885 22274 5895
rect 22288 5885 25730 5895
rect 25744 5885 26426 5895
rect 6304 5861 7370 5871
rect 7384 5861 18290 5871
rect 18304 5861 21314 5871
rect 21328 5861 21530 5871
rect 21544 5861 24434 5871
rect 6232 5837 9314 5847
rect 9736 5837 17810 5847
rect 19240 5837 19250 5847
rect 19936 5837 19946 5847
rect 6184 5813 6218 5823
rect 6280 5813 9794 5823
rect 9808 5813 21290 5823
rect 6136 5789 16466 5799
rect 19072 5789 27002 5799
rect 5872 5765 7394 5775
rect 7408 5765 12794 5775
rect 12856 5765 21098 5775
rect 5824 5741 9506 5751
rect 9520 5741 10130 5751
rect 10144 5741 21554 5751
rect 5800 5717 7802 5727
rect 7936 5717 9554 5727
rect 9568 5717 11834 5727
rect 11848 5717 12266 5727
rect 12520 5717 16010 5727
rect 16240 5717 17306 5727
rect 19048 5717 19070 5727
rect 19216 5717 20546 5727
rect 5752 5693 6890 5703
rect 6904 5693 8090 5703
rect 8104 5693 9650 5703
rect 9664 5693 22562 5703
rect 5752 5669 23522 5679
rect 5728 5645 7154 5655
rect 7168 5645 8738 5655
rect 8752 5645 16970 5655
rect 16984 5645 27098 5655
rect 5704 5621 5714 5631
rect 5776 5621 25418 5631
rect 5656 5597 8834 5607
rect 9280 5597 17354 5607
rect 18856 5597 25370 5607
rect 5248 5573 16538 5583
rect 16840 5573 19106 5583
rect 19120 5573 19634 5583
rect 19648 5573 23882 5583
rect 5176 5549 19346 5559
rect 19504 5549 24290 5559
rect 5080 5525 5210 5535
rect 5224 5525 22922 5535
rect 5056 5501 7250 5511
rect 7312 5501 8306 5511
rect 8320 5501 21050 5511
rect 21064 5501 27050 5511
rect 5008 5477 6602 5487
rect 6616 5477 17090 5487
rect 17392 5477 17474 5487
rect 18640 5477 20282 5487
rect 5008 5453 22778 5463
rect 4936 5429 8066 5439
rect 8080 5429 12002 5439
rect 12016 5429 14666 5439
rect 14680 5429 17234 5439
rect 17248 5429 21914 5439
rect 4864 5405 9074 5415
rect 9088 5405 9386 5415
rect 9400 5405 19202 5415
rect 19216 5405 23642 5415
rect 4792 5381 17258 5391
rect 17272 5381 17858 5391
rect 18256 5381 18386 5391
rect 18544 5381 20402 5391
rect 4792 5357 20738 5367
rect 4744 5333 6002 5343
rect 6016 5333 9434 5343
rect 9448 5333 13346 5343
rect 13360 5333 13874 5343
rect 13888 5333 15770 5343
rect 15784 5333 18266 5343
rect 18280 5333 21866 5343
rect 4720 5309 26930 5319
rect 4696 5285 8858 5295
rect 9208 5285 13994 5295
rect 14008 5285 21410 5295
rect 21424 5285 22130 5295
rect 4672 5261 4826 5271
rect 4888 5261 9122 5271
rect 9184 5261 9338 5271
rect 9688 5261 21818 5271
rect 21832 5261 22034 5271
rect 22048 5261 25970 5271
rect 25984 5261 26378 5271
rect 4648 5237 11018 5247
rect 11032 5237 11450 5247
rect 11464 5237 12554 5247
rect 12568 5237 18986 5247
rect 19000 5237 25322 5247
rect 4576 5213 11714 5223
rect 11776 5213 13538 5223
rect 14080 5213 16730 5223
rect 16744 5213 17594 5223
rect 17608 5213 23930 5223
rect 23944 5213 26594 5223
rect 4504 5189 6194 5199
rect 6208 5189 14474 5199
rect 14488 5189 14738 5199
rect 14872 5189 15458 5199
rect 15472 5189 20354 5199
rect 20800 5189 22154 5199
rect 4408 5165 22754 5175
rect 22768 5165 25514 5175
rect 4360 5141 9290 5151
rect 9640 5141 16490 5151
rect 16720 5141 16802 5151
rect 17032 5141 20762 5151
rect 4264 5117 13226 5127
rect 13288 5117 25898 5127
rect 4264 5093 15842 5103
rect 15952 5093 21110 5103
rect 21124 5093 23570 5103
rect 4192 5069 6506 5079
rect 6520 5069 10106 5079
rect 10120 5069 12578 5079
rect 12592 5069 12674 5079
rect 12688 5069 13970 5079
rect 13984 5069 21002 5079
rect 21016 5069 22298 5079
rect 22312 5069 23882 5079
rect 23896 5069 26354 5079
rect 4120 5045 22970 5055
rect 3952 5021 8522 5031
rect 8536 5021 10226 5031
rect 10240 5021 15794 5031
rect 15808 5021 22970 5031
rect 3904 4997 4082 5007
rect 4096 4997 6842 5007
rect 6856 4997 12218 5007
rect 12232 4997 12818 5007
rect 12832 4997 19922 5007
rect 19936 4997 20618 5007
rect 20632 4997 24194 5007
rect 24208 4997 26762 5007
rect 3832 4973 7538 4983
rect 7600 4973 26450 4983
rect 3808 4949 19466 4959
rect 19672 4949 19730 4959
rect 19912 4949 20474 4959
rect 20728 4949 20786 4959
rect 21688 4949 21722 4959
rect 22624 4949 22934 4959
rect 3520 4925 10106 4935
rect 10120 4925 10970 4935
rect 10984 4925 13442 4935
rect 13456 4925 20954 4935
rect 20968 4925 21674 4935
rect 21688 4925 22322 4935
rect 22336 4925 25082 4935
rect 25096 4925 25466 4935
rect 3448 4901 8618 4911
rect 8632 4901 16706 4911
rect 16720 4901 22850 4911
rect 3376 4877 4850 4887
rect 4864 4877 7106 4887
rect 7120 4877 9746 4887
rect 9760 4877 18962 4887
rect 18976 4877 19226 4887
rect 19240 4877 19850 4887
rect 19864 4877 22610 4887
rect 22624 4877 23450 4887
rect 23464 4877 23786 4887
rect 23800 4877 26090 4887
rect 3304 4853 8978 4863
rect 9088 4853 13034 4863
rect 13096 4853 20162 4863
rect 20512 4853 22826 4863
rect 3160 4829 25922 4839
rect 3112 4805 16082 4815
rect 16192 4805 20714 4815
rect 3064 4781 21458 4791
rect 3040 4757 19034 4767
rect 19048 4757 20834 4767
rect 20848 4757 25202 4767
rect 2944 4733 8786 4743
rect 8944 4733 21242 4743
rect 22648 4733 23174 4743
rect 2920 4709 14954 4719
rect 14968 4709 16322 4719
rect 16600 4709 23210 4719
rect 2848 4685 7226 4695
rect 7240 4685 24770 4695
rect 24784 4685 27122 4695
rect 2824 4661 5330 4671
rect 5344 4661 5690 4671
rect 5704 4661 5882 4671
rect 5896 4661 5954 4671
rect 5968 4661 10610 4671
rect 10624 4661 12098 4671
rect 12112 4661 24962 4671
rect 2752 4637 4514 4647
rect 4528 4637 5930 4647
rect 5944 4637 10250 4647
rect 10264 4637 12026 4647
rect 12040 4637 12194 4647
rect 12208 4637 12914 4647
rect 12928 4637 13826 4647
rect 13840 4637 18362 4647
rect 18376 4637 22994 4647
rect 23824 4637 25610 4647
rect 2680 4613 23018 4623
rect 23128 4613 23498 4623
rect 23560 4613 23834 4623
rect 24160 4613 26858 4623
rect 2632 4589 10754 4599
rect 10768 4589 24890 4599
rect 24904 4589 26786 4599
rect 2608 4565 24170 4575
rect 25144 4565 25178 4575
rect 25288 4565 25298 4575
rect 25672 4565 25682 4575
rect 26008 4565 27853 4575
rect 2536 4541 7850 4551
rect 7864 4541 7970 4551
rect 7984 4541 9026 4551
rect 9040 4541 9890 4551
rect 9904 4541 20378 4551
rect 20392 4541 20834 4551
rect 20848 4541 26810 4551
rect 2488 4517 3530 4527
rect 3544 4517 10010 4527
rect 10024 4517 15290 4527
rect 15304 4517 24434 4527
rect 25336 4517 25370 4527
rect 26824 4517 27050 4527
rect 2416 4493 5618 4503
rect 5632 4493 5666 4503
rect 5680 4493 8594 4503
rect 8608 4493 9674 4503
rect 9688 4493 13010 4503
rect 13024 4493 13370 4503
rect 13384 4493 17186 4503
rect 17200 4493 18410 4503
rect 18424 4493 20594 4503
rect 20608 4493 26642 4503
rect 2392 4469 11426 4479
rect 11440 4469 16754 4479
rect 16768 4469 18314 4479
rect 18328 4469 26498 4479
rect 2344 4445 10730 4455
rect 10792 4445 13442 4455
rect 13504 4445 16802 4455
rect 17224 4445 21074 4455
rect 21328 4445 24578 4455
rect 26512 4445 26642 4455
rect 2320 4421 3770 4431
rect 3784 4421 4034 4431
rect 4048 4421 7274 4431
rect 7288 4421 10562 4431
rect 10576 4421 15362 4431
rect 15376 4421 16682 4431
rect 16696 4421 23114 4431
rect 23128 4421 25130 4431
rect 25144 4421 27314 4431
rect 2296 4397 14090 4407
rect 14200 4397 14810 4407
rect 15136 4397 24026 4407
rect 24400 4397 26978 4407
rect 2248 4373 4226 4383
rect 4240 4373 5282 4383
rect 5416 4373 19442 4383
rect 19600 4373 20210 4383
rect 20656 4373 25178 4383
rect 2224 4349 6578 4359
rect 6592 4349 9602 4359
rect 9616 4349 17066 4359
rect 17080 4349 18266 4359
rect 18280 4349 19322 4359
rect 19336 4349 22994 4359
rect 23008 4349 23282 4359
rect 23296 4349 24122 4359
rect 24136 4349 24338 4359
rect 24352 4349 24554 4359
rect 24568 4349 26402 4359
rect 2200 4325 3866 4335
rect 3880 4325 4298 4335
rect 4312 4325 8186 4335
rect 8200 4325 12362 4335
rect 12376 4325 13850 4335
rect 13864 4325 14258 4335
rect 14272 4325 23786 4335
rect 24352 4325 24494 4335
rect 26416 4325 26450 4335
rect 2104 4301 13322 4311
rect 13336 4301 19562 4311
rect 19576 4301 26906 4311
rect 2080 4277 8570 4287
rect 8584 4277 10178 4287
rect 10312 4277 26834 4287
rect 2008 4253 10322 4263
rect 10336 4253 12122 4263
rect 12136 4253 12890 4263
rect 12904 4253 20054 4263
rect 20068 4253 21194 4263
rect 21208 4253 23810 4263
rect 23824 4253 26186 4263
rect 1984 4229 3002 4239
rect 3016 4229 3266 4239
rect 3280 4229 8858 4239
rect 8872 4229 10634 4239
rect 10648 4229 20114 4239
rect 20128 4229 21650 4239
rect 21664 4229 25394 4239
rect 1960 4205 5594 4215
rect 5608 4205 18074 4215
rect 18088 4205 21242 4215
rect 21256 4205 22898 4215
rect 22912 4205 26066 4215
rect 1912 4181 23954 4191
rect 25408 4181 25418 4191
rect 1864 4157 3218 4167
rect 3232 4157 3698 4167
rect 3712 4157 4634 4167
rect 4648 4157 6170 4167
rect 6184 4157 7874 4167
rect 7888 4157 9146 4167
rect 9160 4157 11930 4167
rect 11944 4157 13922 4167
rect 13936 4157 18602 4167
rect 18616 4157 20138 4167
rect 20152 4157 21194 4167
rect 21208 4157 22394 4167
rect 22408 4157 22538 4167
rect 22552 4157 26042 4167
rect 1840 4133 8906 4143
rect 8920 4133 11618 4143
rect 11872 4133 24458 4143
rect 1768 4109 2690 4119
rect 2704 4109 6098 4119
rect 6112 4109 6650 4119
rect 6664 4109 6962 4119
rect 6976 4109 8114 4119
rect 8128 4109 9482 4119
rect 9496 4109 17114 4119
rect 17128 4109 17882 4119
rect 18184 4109 18674 4119
rect 19000 4109 19178 4119
rect 19576 4109 19802 4119
rect 19864 4109 20330 4119
rect 20944 4109 21482 4119
rect 22072 4109 23762 4119
rect 1744 4085 3386 4095
rect 3400 4085 3482 4095
rect 3496 4085 4010 4095
rect 4024 4085 4202 4095
rect 4216 4085 11210 4095
rect 11224 4085 11810 4095
rect 11824 4085 14042 4095
rect 14056 4085 15410 4095
rect 15424 4085 18242 4095
rect 18256 4085 18458 4095
rect 18472 4085 19394 4095
rect 19408 4085 19970 4095
rect 19984 4085 25346 4095
rect 25360 4085 25442 4095
rect 25456 4085 26162 4095
rect 1720 4061 6530 4071
rect 6544 4061 13010 4071
rect 13024 4061 14882 4071
rect 14896 4061 15482 4071
rect 15496 4061 26666 4071
rect 1672 4037 9986 4047
rect 10072 4037 17690 4047
rect 19816 4037 27026 4047
rect 1648 4013 3218 4023
rect 3232 4013 7442 4023
rect 7456 4013 7730 4023
rect 7744 4013 7994 4023
rect 8008 4013 12698 4023
rect 12712 4013 18482 4023
rect 18496 4013 20858 4023
rect 20872 4013 21698 4023
rect 22720 4013 23366 4023
rect 25456 4013 27410 4023
rect 1624 3989 4610 3999
rect 4624 3989 13634 3999
rect 13648 3989 18050 3999
rect 19984 3989 20054 3999
rect 20152 3989 25034 3999
rect 84 3965 8138 3975
rect 8152 3965 16994 3975
rect 17320 3965 21434 3975
rect 22816 3965 23306 3975
rect 84 3941 9410 3951
rect 9616 3941 9818 3951
rect 9904 3941 9914 3951
rect 10096 3941 22010 3951
rect 22024 3941 26618 3951
rect 1624 3917 9170 3927
rect 9184 3917 13898 3927
rect 14080 3917 14138 3927
rect 15232 3917 15602 3927
rect 15688 3917 15722 3927
rect 16288 3917 17522 3927
rect 20872 3917 21002 3927
rect 21352 3917 23498 3927
rect 1648 3893 3554 3903
rect 3568 3893 4946 3903
rect 4960 3893 5978 3903
rect 5992 3893 9458 3903
rect 9472 3893 14690 3903
rect 14704 3893 16154 3903
rect 16168 3893 26258 3903
rect 1792 3869 26666 3879
rect 2032 3845 8306 3855
rect 9016 3845 19682 3855
rect 20968 3845 21110 3855
rect 21376 3845 21938 3855
rect 23296 3845 27853 3855
rect 2176 3821 9242 3831
rect 9256 3821 21170 3831
rect 2224 3797 3242 3807
rect 3256 3797 5426 3807
rect 5440 3797 6818 3807
rect 6832 3797 9578 3807
rect 9592 3797 13418 3807
rect 13432 3797 13898 3807
rect 13912 3797 19778 3807
rect 19792 3797 20090 3807
rect 20104 3797 21554 3807
rect 21568 3797 22634 3807
rect 22648 3797 24650 3807
rect 24664 3797 25826 3807
rect 2440 3773 13586 3783
rect 15424 3773 15434 3783
rect 16528 3773 23402 3783
rect 2512 3749 6626 3759
rect 6640 3749 7154 3759
rect 7168 3749 12002 3759
rect 12016 3749 13658 3759
rect 13672 3749 19874 3759
rect 19888 3749 21026 3759
rect 2584 3725 5114 3735
rect 5128 3725 11330 3735
rect 11608 3725 13802 3735
rect 16768 3725 25778 3735
rect 2608 3701 3602 3711
rect 3616 3701 11354 3711
rect 11368 3701 15194 3711
rect 15208 3701 22178 3711
rect 22192 3701 22346 3711
rect 22360 3701 26258 3711
rect 2656 3677 23666 3687
rect 2704 3653 5450 3663
rect 5512 3653 9266 3663
rect 9280 3653 18146 3663
rect 18160 3653 19106 3663
rect 19120 3653 24530 3663
rect 24544 3653 25274 3663
rect 2872 3629 26234 3639
rect 3280 3605 4418 3615
rect 4432 3605 8114 3615
rect 8128 3605 9050 3615
rect 9064 3605 10946 3615
rect 10960 3605 13130 3615
rect 13144 3605 17522 3615
rect 17536 3605 22250 3615
rect 24544 3605 24698 3615
rect 3328 3581 9578 3591
rect 9760 3581 12866 3591
rect 13072 3581 22490 3591
rect 3424 3557 20450 3567
rect 20464 3557 22934 3567
rect 3472 3533 3674 3543
rect 3688 3533 24626 3543
rect 3592 3509 13394 3519
rect 13480 3509 16058 3519
rect 17464 3509 24314 3519
rect 24328 3509 26474 3519
rect 3616 3485 23426 3495
rect 3640 3461 11282 3471
rect 11824 3461 17498 3471
rect 20464 3461 20474 3471
rect 3712 3437 16874 3447
rect 3736 3413 7586 3423
rect 7648 3413 10826 3423
rect 10840 3413 12050 3423
rect 12064 3413 17330 3423
rect 3760 3389 17162 3399
rect 17176 3389 19154 3399
rect 3808 3365 10442 3375
rect 10456 3365 19010 3375
rect 19168 3365 25106 3375
rect 3880 3341 8954 3351
rect 8968 3341 26546 3351
rect 3928 3317 5906 3327
rect 5920 3317 8714 3327
rect 8728 3317 8834 3327
rect 8848 3317 21530 3327
rect 21544 3317 21722 3327
rect 4000 3293 7034 3303
rect 7048 3293 12170 3303
rect 12184 3293 12626 3303
rect 12640 3293 17378 3303
rect 4024 3269 5714 3279
rect 5728 3269 8978 3279
rect 8992 3269 19070 3279
rect 19084 3269 19442 3279
rect 19456 3269 19658 3279
rect 19672 3269 20666 3279
rect 20680 3269 22442 3279
rect 4072 3245 10466 3255
rect 10480 3245 23858 3255
rect 23872 3245 24098 3255
rect 4120 3221 6914 3231
rect 6928 3221 10514 3231
rect 10528 3221 20594 3231
rect 20608 3221 23066 3231
rect 4336 3197 6122 3207
rect 6208 3197 21794 3207
rect 4360 3173 6218 3183
rect 6232 3173 13730 3183
rect 13744 3173 19754 3183
rect 21808 3173 21818 3183
rect 4432 3149 12602 3159
rect 12616 3149 14234 3159
rect 14248 3149 14930 3159
rect 14944 3149 24026 3159
rect 4456 3125 13514 3135
rect 16888 3125 16898 3135
rect 4552 3101 6314 3111
rect 6328 3101 6698 3111
rect 6712 3101 8642 3111
rect 8656 3101 13034 3111
rect 13048 3101 20258 3111
rect 20272 3101 26690 3111
rect 4576 3077 6386 3087
rect 6400 3077 6986 3087
rect 7000 3077 7490 3087
rect 7504 3077 8738 3087
rect 8752 3077 8762 3087
rect 8776 3077 17474 3087
rect 17488 3077 17666 3087
rect 17680 3077 19130 3087
rect 19144 3077 19346 3087
rect 19360 3077 22514 3087
rect 4672 3053 10586 3063
rect 10600 3053 12962 3063
rect 12976 3053 16946 3063
rect 16960 3053 17402 3063
rect 17416 3053 19994 3063
rect 20008 3053 25226 3063
rect 4744 3029 7658 3039
rect 7672 3029 11306 3039
rect 11320 3029 23906 3039
rect 4768 3005 7730 3015
rect 7744 3005 26522 3015
rect 4840 2981 6482 2991
rect 6496 2981 22874 2991
rect 22888 2981 23690 2991
rect 5128 2957 25154 2967
rect 5200 2933 12146 2943
rect 12208 2933 12290 2943
rect 12448 2933 12530 2943
rect 12736 2933 18866 2943
rect 19144 2933 19610 2943
rect 5536 2909 6674 2919
rect 6688 2909 25514 2919
rect 5560 2885 16826 2895
rect 16960 2885 17354 2895
rect 5728 2861 16418 2871
rect 16432 2861 16778 2871
rect 16792 2861 20522 2871
rect 20536 2861 24074 2871
rect 24088 2861 26738 2871
rect 5824 2837 8018 2847
rect 8032 2837 13202 2847
rect 13216 2837 20306 2847
rect 26752 2837 26954 2847
rect 6016 2813 14282 2823
rect 14296 2813 15026 2823
rect 15040 2813 16922 2823
rect 16936 2813 17426 2823
rect 17440 2813 19514 2823
rect 19528 2813 21602 2823
rect 6040 2789 19514 2799
rect 20320 2789 20354 2799
rect 6088 2765 8066 2775
rect 8200 2765 23174 2775
rect 6232 2741 7178 2751
rect 7192 2741 7778 2751
rect 7792 2741 15386 2751
rect 15400 2741 17282 2751
rect 17296 2741 18386 2751
rect 18400 2741 21074 2751
rect 21088 2741 21218 2751
rect 21232 2741 23330 2751
rect 23344 2741 23354 2751
rect 6472 2717 14138 2727
rect 16936 2717 17330 2727
rect 23344 2717 23618 2727
rect 6544 2693 16346 2703
rect 16360 2693 19250 2703
rect 19264 2693 23522 2703
rect 6688 2669 16562 2679
rect 16576 2669 19730 2679
rect 6736 2645 8522 2655
rect 8536 2645 14714 2655
rect 6784 2621 12650 2631
rect 12664 2621 17978 2631
rect 7096 2597 9098 2607
rect 9112 2597 10370 2607
rect 10384 2597 13106 2607
rect 13168 2597 23978 2607
rect 7120 2573 7130 2583
rect 7216 2573 13346 2583
rect 13360 2573 16130 2583
rect 16144 2573 23042 2583
rect 23056 2573 26882 2583
rect 7720 2549 9530 2559
rect 9544 2549 11546 2559
rect 11560 2549 23234 2559
rect 23248 2549 26306 2559
rect 7768 2525 27410 2535
rect 7816 2501 22682 2511
rect 7864 2477 25802 2487
rect 7984 2453 8402 2463
rect 8656 2453 11234 2463
rect 11920 2453 12242 2463
rect 12256 2453 17762 2463
rect 8032 2429 10946 2439
rect 10960 2429 19946 2439
rect 8248 2405 23258 2415
rect 23272 2405 24362 2415
rect 8272 2381 9554 2391
rect 9568 2381 11570 2391
rect 11584 2381 23594 2391
rect 24376 2381 24602 2391
rect 8968 2357 9218 2367
rect 9232 2357 12482 2367
rect 12784 2357 15866 2367
rect 9064 2333 9698 2343
rect 9712 2333 24722 2343
rect 9232 2309 13778 2319
rect 9256 2285 9290 2295
rect 9376 2285 13610 2295
rect 13792 2285 24674 2295
rect 24688 2285 25586 2295
rect 9424 2261 11138 2271
rect 11152 2261 11162 2271
rect 11176 2261 20978 2271
rect 20992 2261 24242 2271
rect 24256 2261 26522 2271
rect 9472 2237 9794 2247
rect 10192 2237 12458 2247
rect 12808 2237 13562 2247
rect 13624 2237 21746 2247
rect 21760 2237 26210 2247
rect 10360 2213 14402 2223
rect 10408 2189 24722 2199
rect 10504 2165 21290 2175
rect 10576 2141 10610 2151
rect 10672 2141 17618 2151
rect 17632 2141 25298 2151
rect 10912 2117 18770 2127
rect 10984 2093 11066 2103
rect 11128 2093 21458 2103
rect 11152 2069 12074 2079
rect 12088 2069 16250 2079
rect 16264 2069 18338 2079
rect 18352 2069 19898 2079
rect 19912 2069 22874 2079
rect 22888 2069 27338 2079
rect 13120 2045 18890 2055
rect 18904 2045 20882 2055
rect 13264 2021 22514 2031
rect 13480 1997 21986 2007
rect 22000 1997 25754 2007
rect 27448 1997 27853 2007
rect 13552 1973 15050 1983
rect 27424 1973 27853 1983
rect 26955 1944 27435 1954
rect 26955 1921 27435 1931
rect 26955 1883 27435 1908
rect 26955 1238 27435 1263
rect 16432 1140 23378 1150
rect 15880 1116 18842 1126
rect 14584 1092 23954 1102
rect 13216 1068 22922 1078
rect 13168 1044 14594 1054
rect 14800 1044 23426 1054
rect 23440 1044 24482 1054
rect 12688 1020 23738 1030
rect 12328 996 18098 1006
rect 11056 972 17114 982
rect 10936 948 13850 958
rect 14464 948 21122 958
rect 10864 924 23906 934
rect 10720 900 19274 910
rect 10024 876 18194 886
rect 10000 852 13730 862
rect 14368 852 16610 862
rect 9952 828 24122 838
rect 9520 804 21626 814
rect 22576 804 23642 814
rect 9136 780 22778 790
rect 8800 756 14930 766
rect 14944 756 19418 766
rect 20224 756 20690 766
rect 22480 756 26882 766
rect 7336 732 15698 742
rect 15760 732 16442 742
rect 20176 732 24602 742
rect 7240 708 13802 718
rect 14056 708 17690 718
rect 18016 708 20498 718
rect 20632 706 20650 720
rect 22216 708 27853 718
rect 6976 684 16850 694
rect 17920 684 23690 694
rect 6424 660 24002 670
rect 6256 636 12338 646
rect 12400 636 17498 646
rect 17752 636 26690 646
rect 6112 612 11186 622
rect 11248 612 26450 622
rect 5992 588 8714 598
rect 8728 588 15506 598
rect 15520 588 20042 598
rect 20056 588 20402 598
rect 20416 588 24242 598
rect 5944 564 7682 574
rect 8296 564 9818 574
rect 9880 564 15074 574
rect 15160 564 23186 574
rect 23200 564 26930 574
rect 5848 540 19754 550
rect 5488 516 6746 526
rect 6952 516 20978 526
rect 4960 492 6026 502
rect 6088 492 7418 502
rect 7480 492 20090 502
rect 4936 468 20546 478
rect 4888 444 23714 454
rect 4600 420 20426 430
rect 4480 396 20378 406
rect 20392 396 24266 406
rect 4216 372 14306 382
rect 14536 372 17066 382
rect 4168 348 10034 358
rect 10648 348 10682 358
rect 10768 348 15170 358
rect 15328 348 15554 358
rect 15640 348 26954 358
rect 3688 324 4298 334
rect 4312 324 10274 334
rect 10288 324 22106 334
rect 3664 300 21002 310
rect 3544 276 16994 286
rect 2872 252 14618 262
rect 14848 252 26594 262
rect 2752 228 26642 238
rect 2536 204 26618 214
rect 2488 180 8426 190
rect 8560 180 16802 190
rect 1816 156 7610 166
rect 8044 156 22706 166
rect 1696 132 11018 142
rect 11104 132 20738 142
rect 84 108 19850 118
rect 84 84 2354 94
rect 2416 84 18434 94
rect 2632 60 27853 70
rect 4144 36 8066 46
rect 8392 36 24074 46
rect 26944 36 27853 46
rect 11968 12 26930 22
rect 26968 12 27853 22
<< m2contact >>
rect 15938 8276 15952 8290
rect 18782 8276 18796 8290
rect 18914 8276 18928 8290
rect 15602 8252 15616 8266
rect 20510 8252 20524 8266
rect 14810 8228 14824 8242
rect 17102 8228 17116 8242
rect 18674 8228 18688 8242
rect 27434 8228 27448 8242
rect 14666 8204 14680 8218
rect 25622 8204 25636 8218
rect 9938 8180 9952 8194
rect 11930 8180 11944 8194
rect 27242 8180 27256 8194
rect 5978 8156 5992 8170
rect 6962 8156 6976 8170
rect 9818 8156 9832 8170
rect 21362 8156 21376 8170
rect 4082 8132 4096 8146
rect 7646 8132 7660 8146
rect 9338 8132 9352 8146
rect 27050 8132 27064 8146
rect 27302 8132 27316 8146
rect 27410 8132 27424 8146
rect 2210 8108 2224 8122
rect 4190 8108 4204 8122
rect 4730 8108 4744 8122
rect 5054 8108 5068 8122
rect 5522 8108 5536 8122
rect 27482 8108 27496 8122
rect 1706 8084 1720 8098
rect 2462 8084 2476 8098
rect 2954 8084 2968 8098
rect 12830 8084 12844 8098
rect 12914 8084 12928 8098
rect 23918 8084 23932 8098
rect 24554 8084 24568 8098
rect 27530 8084 27544 8098
rect 70 8060 84 8074
rect 26114 8060 26128 8074
rect 70 8036 84 8050
rect 11066 8036 11080 8050
rect 11642 8036 11656 8050
rect 22214 8036 22228 8050
rect 22346 8036 22360 8050
rect 23066 8036 23080 8050
rect 27506 8036 27520 8050
rect 27853 8036 27867 8050
rect 2138 8012 2152 8026
rect 13634 8012 13648 8026
rect 18806 8012 18820 8026
rect 19610 8012 19624 8026
rect 27458 8012 27472 8026
rect 27482 8012 27496 8026
rect 27853 8012 27867 8026
rect 2426 7988 2440 8002
rect 6578 7988 6592 8002
rect 6674 7988 6688 8002
rect 24770 7988 24784 8002
rect 27458 7988 27472 8002
rect 27853 7988 27867 8002
rect 4154 7964 4168 7978
rect 6986 7964 7000 7978
rect 8474 7964 8488 7978
rect 10238 7964 10252 7978
rect 12794 7964 12808 7978
rect 14138 7964 14152 7978
rect 14522 7964 14536 7978
rect 19250 7964 19264 7978
rect 20210 7964 20224 7978
rect 27434 7964 27448 7978
rect 27853 7964 27867 7978
rect 15374 7940 15388 7954
rect 16370 7940 16384 7954
rect 16874 7940 16888 7954
rect 18098 7940 18112 7954
rect 27506 7940 27520 7954
rect 27530 7940 27544 7954
rect 27853 7940 27867 7954
rect 13682 7107 13696 7121
rect 13802 7107 13816 7121
rect 14666 7107 14680 7121
rect 14714 7107 14728 7121
rect 13514 7083 13528 7097
rect 17138 7083 17152 7097
rect 13370 7059 13384 7073
rect 15722 7059 15736 7073
rect 16466 7059 16480 7073
rect 26378 7059 26392 7073
rect 13322 7035 13336 7049
rect 13658 7035 13672 7049
rect 14618 7035 14632 7049
rect 25538 7035 25552 7049
rect 12866 7011 12880 7025
rect 13706 7011 13720 7025
rect 18098 7011 18112 7025
rect 12818 6987 12832 7001
rect 12866 6987 12880 7001
rect 12986 6987 13000 7001
rect 26426 6987 26440 7001
rect 12626 6963 12640 6977
rect 22730 6963 22744 6977
rect 25562 6963 25576 6977
rect 25778 6963 25792 6977
rect 12098 6939 12112 6953
rect 12170 6939 12184 6953
rect 12578 6939 12592 6953
rect 17954 6939 17968 6953
rect 25562 6939 25576 6953
rect 11954 6915 11968 6929
rect 15986 6915 16000 6929
rect 16274 6915 16288 6929
rect 19778 6915 19792 6929
rect 11162 6891 11176 6905
rect 19538 6891 19552 6905
rect 19706 6891 19720 6905
rect 25706 6891 25720 6905
rect 10826 6867 10840 6881
rect 15002 6867 15016 6881
rect 19706 6867 19720 6881
rect 10682 6843 10696 6857
rect 14114 6843 14128 6857
rect 24698 6843 24712 6857
rect 10370 6819 10384 6833
rect 23306 6819 23320 6833
rect 10322 6795 10336 6809
rect 23138 6795 23152 6809
rect 10130 6771 10144 6785
rect 16658 6771 16672 6785
rect 17570 6771 17584 6785
rect 17594 6771 17608 6785
rect 9770 6747 9784 6761
rect 27434 6747 27448 6761
rect 9338 6723 9352 6737
rect 27146 6723 27160 6737
rect 9314 6699 9328 6713
rect 21698 6699 21712 6713
rect 8330 6675 8344 6689
rect 9770 6675 9784 6689
rect 10034 6675 10048 6689
rect 18578 6675 18592 6689
rect 26042 6675 26056 6689
rect 8330 6651 8344 6665
rect 8474 6651 8488 6665
rect 8546 6651 8560 6665
rect 11690 6651 11704 6665
rect 21602 6651 21616 6665
rect 8282 6627 8296 6641
rect 13946 6627 13960 6641
rect 24482 6627 24496 6641
rect 8234 6603 8248 6617
rect 21410 6603 21424 6617
rect 8210 6579 8224 6593
rect 21362 6579 21376 6593
rect 8138 6555 8152 6569
rect 8378 6555 8392 6569
rect 8426 6555 8440 6569
rect 24986 6555 25000 6569
rect 7754 6531 7768 6545
rect 9914 6531 9928 6545
rect 10850 6531 10864 6545
rect 20042 6531 20056 6545
rect 7682 6507 7696 6521
rect 18722 6507 18736 6521
rect 26570 6507 26584 6521
rect 7658 6483 7672 6497
rect 12290 6483 12304 6497
rect 27362 6483 27376 6497
rect 7562 6459 7576 6473
rect 25850 6459 25864 6473
rect 7514 6435 7528 6449
rect 9698 6435 9712 6449
rect 12530 6435 12544 6449
rect 15434 6435 15448 6449
rect 15698 6435 15712 6449
rect 23618 6435 23632 6449
rect 7514 6411 7528 6425
rect 22754 6411 22768 6425
rect 7466 6387 7480 6401
rect 20258 6387 20272 6401
rect 7418 6363 7432 6377
rect 23210 6363 23224 6377
rect 24494 6363 24508 6377
rect 7370 6339 7384 6353
rect 9362 6339 9376 6353
rect 9866 6339 9880 6353
rect 15578 6339 15592 6353
rect 20906 6339 20920 6353
rect 24602 6339 24616 6353
rect 7322 6315 7336 6329
rect 7922 6315 7936 6329
rect 8042 6315 8056 6329
rect 8666 6315 8680 6329
rect 8882 6315 8896 6329
rect 19298 6315 19312 6329
rect 7298 6291 7312 6305
rect 17570 6291 17584 6305
rect 7082 6267 7096 6281
rect 11498 6267 11512 6281
rect 17642 6267 17656 6281
rect 19322 6267 19336 6281
rect 21578 6267 21592 6281
rect 22418 6267 22432 6281
rect 7058 6243 7072 6257
rect 21146 6243 21160 6257
rect 7010 6219 7024 6233
rect 11258 6219 11272 6233
rect 11378 6219 11392 6233
rect 11954 6219 11968 6233
rect 12050 6219 12064 6233
rect 12074 6219 12088 6233
rect 12146 6219 12160 6233
rect 12314 6219 12328 6233
rect 17042 6219 17056 6233
rect 24410 6219 24424 6233
rect 6914 6195 6928 6209
rect 14018 6195 14032 6209
rect 27194 6195 27208 6209
rect 6866 6171 6880 6185
rect 10226 6171 10240 6185
rect 14906 6171 14920 6185
rect 20522 6171 20536 6185
rect 23090 6171 23104 6185
rect 23366 6171 23380 6185
rect 23474 6171 23488 6185
rect 25946 6171 25960 6185
rect 6866 6147 6880 6161
rect 15674 6147 15688 6161
rect 16034 6147 16048 6161
rect 23474 6147 23488 6161
rect 6818 6123 6832 6137
rect 12434 6123 12448 6137
rect 12554 6123 12568 6137
rect 12650 6123 12664 6137
rect 12722 6123 12736 6137
rect 23090 6123 23104 6137
rect 24842 6123 24856 6137
rect 6770 6099 6784 6113
rect 7034 6099 7048 6113
rect 19418 6099 19432 6113
rect 6698 6075 6712 6089
rect 25082 6075 25096 6089
rect 6650 6051 6664 6065
rect 7130 6051 7144 6065
rect 8498 6051 8512 6065
rect 10442 6051 10456 6065
rect 13682 6051 13696 6065
rect 14258 6051 14272 6065
rect 16898 6051 16912 6065
rect 6602 6027 6616 6041
rect 22802 6027 22816 6041
rect 6578 6003 6592 6017
rect 6698 6003 6712 6017
rect 6746 6003 6760 6017
rect 15650 6003 15664 6017
rect 19178 6003 19192 6017
rect 22658 6003 22672 6017
rect 25634 6003 25648 6017
rect 6554 5979 6568 5993
rect 10466 5979 10480 5993
rect 20018 5979 20032 5993
rect 22346 5979 22360 5993
rect 6410 5955 6424 5969
rect 8882 5955 8896 5969
rect 19370 5955 19384 5969
rect 6362 5931 6376 5945
rect 10538 5931 10552 5945
rect 10586 5931 10600 5945
rect 10802 5931 10816 5945
rect 10898 5931 10912 5945
rect 15266 5931 15280 5945
rect 23162 5931 23176 5945
rect 6338 5907 6352 5921
rect 7946 5907 7960 5921
rect 12026 5907 12040 5921
rect 13754 5907 13768 5921
rect 13970 5907 13984 5921
rect 17210 5907 17224 5921
rect 21338 5907 21352 5921
rect 26306 5907 26320 5921
rect 26954 5907 26968 5921
rect 6314 5883 6328 5897
rect 6338 5883 6352 5897
rect 12122 5883 12136 5897
rect 14378 5883 14392 5897
rect 15458 5883 15472 5897
rect 16682 5883 16696 5897
rect 22274 5883 22288 5897
rect 25730 5883 25744 5897
rect 26426 5883 26440 5897
rect 6290 5859 6304 5873
rect 7370 5859 7384 5873
rect 18290 5859 18304 5873
rect 21314 5859 21328 5873
rect 21530 5859 21544 5873
rect 24434 5859 24448 5873
rect 6218 5835 6232 5849
rect 9314 5835 9328 5849
rect 9722 5835 9736 5849
rect 17810 5835 17824 5849
rect 19226 5835 19240 5849
rect 19250 5835 19264 5849
rect 19922 5835 19936 5849
rect 19946 5835 19960 5849
rect 6170 5811 6184 5825
rect 6218 5811 6232 5825
rect 6266 5811 6280 5825
rect 9794 5811 9808 5825
rect 21290 5811 21304 5825
rect 6122 5787 6136 5801
rect 16466 5787 16480 5801
rect 19058 5787 19072 5801
rect 27002 5787 27016 5801
rect 5858 5763 5872 5777
rect 7394 5763 7408 5777
rect 12794 5763 12808 5777
rect 12842 5763 12856 5777
rect 21098 5763 21112 5777
rect 5810 5739 5824 5753
rect 9506 5739 9520 5753
rect 10130 5739 10144 5753
rect 21554 5739 21568 5753
rect 5786 5715 5800 5729
rect 7802 5715 7816 5729
rect 7922 5715 7936 5729
rect 9554 5715 9568 5729
rect 11834 5715 11848 5729
rect 12266 5715 12280 5729
rect 12506 5715 12520 5729
rect 16010 5715 16024 5729
rect 16226 5715 16240 5729
rect 17306 5715 17320 5729
rect 19034 5715 19048 5729
rect 19070 5715 19084 5729
rect 19202 5715 19216 5729
rect 20546 5715 20560 5729
rect 5738 5691 5752 5705
rect 6890 5691 6904 5705
rect 8090 5691 8104 5705
rect 9650 5691 9664 5705
rect 22562 5691 22576 5705
rect 5738 5667 5752 5681
rect 23522 5667 23536 5681
rect 5714 5643 5728 5657
rect 7154 5643 7168 5657
rect 8738 5643 8752 5657
rect 16970 5643 16984 5657
rect 27098 5643 27112 5657
rect 5690 5619 5704 5633
rect 5714 5619 5728 5633
rect 5762 5619 5776 5633
rect 25418 5619 25432 5633
rect 5642 5595 5656 5609
rect 8834 5595 8848 5609
rect 9266 5595 9280 5609
rect 17354 5595 17368 5609
rect 18842 5595 18856 5609
rect 25370 5595 25384 5609
rect 5234 5571 5248 5585
rect 16538 5571 16552 5585
rect 16826 5571 16840 5585
rect 19106 5571 19120 5585
rect 19634 5571 19648 5585
rect 23882 5571 23896 5585
rect 5162 5547 5176 5561
rect 19346 5547 19360 5561
rect 19490 5547 19504 5561
rect 24290 5547 24304 5561
rect 5066 5523 5080 5537
rect 5210 5523 5224 5537
rect 22922 5523 22936 5537
rect 5042 5499 5056 5513
rect 7250 5499 7264 5513
rect 7298 5499 7312 5513
rect 8306 5499 8320 5513
rect 21050 5499 21064 5513
rect 27050 5499 27064 5513
rect 4994 5475 5008 5489
rect 6602 5475 6616 5489
rect 17090 5475 17104 5489
rect 17378 5475 17392 5489
rect 17474 5475 17488 5489
rect 18626 5475 18640 5489
rect 20282 5475 20296 5489
rect 4994 5451 5008 5465
rect 22778 5451 22792 5465
rect 4922 5427 4936 5441
rect 8066 5427 8080 5441
rect 12002 5427 12016 5441
rect 14666 5427 14680 5441
rect 17234 5427 17248 5441
rect 21914 5427 21928 5441
rect 4850 5403 4864 5417
rect 9074 5403 9088 5417
rect 9386 5403 9400 5417
rect 19202 5403 19216 5417
rect 23642 5403 23656 5417
rect 4778 5379 4792 5393
rect 17258 5379 17272 5393
rect 17858 5379 17872 5393
rect 18242 5379 18256 5393
rect 18386 5379 18400 5393
rect 18530 5379 18544 5393
rect 20402 5379 20416 5393
rect 4778 5355 4792 5369
rect 20738 5355 20752 5369
rect 4730 5331 4744 5345
rect 6002 5331 6016 5345
rect 9434 5331 9448 5345
rect 13346 5331 13360 5345
rect 13874 5331 13888 5345
rect 15770 5331 15784 5345
rect 18266 5331 18280 5345
rect 21866 5331 21880 5345
rect 4706 5307 4720 5321
rect 26930 5307 26944 5321
rect 4682 5283 4696 5297
rect 8858 5283 8872 5297
rect 9194 5283 9208 5297
rect 13994 5283 14008 5297
rect 21410 5283 21424 5297
rect 22130 5283 22144 5297
rect 4658 5259 4672 5273
rect 4826 5259 4840 5273
rect 4874 5259 4888 5273
rect 9122 5259 9136 5273
rect 9170 5259 9184 5273
rect 9338 5259 9352 5273
rect 9674 5259 9688 5273
rect 21818 5259 21832 5273
rect 22034 5259 22048 5273
rect 25970 5259 25984 5273
rect 26378 5259 26392 5273
rect 4634 5235 4648 5249
rect 11018 5235 11032 5249
rect 11450 5235 11464 5249
rect 12554 5235 12568 5249
rect 18986 5235 19000 5249
rect 25322 5235 25336 5249
rect 4562 5211 4576 5225
rect 11714 5211 11728 5225
rect 11762 5211 11776 5225
rect 13538 5211 13552 5225
rect 14066 5211 14080 5225
rect 16730 5211 16744 5225
rect 17594 5211 17608 5225
rect 23930 5211 23944 5225
rect 26594 5211 26608 5225
rect 4490 5187 4504 5201
rect 6194 5187 6208 5201
rect 14474 5187 14488 5201
rect 14738 5187 14752 5201
rect 14858 5187 14872 5201
rect 15458 5187 15472 5201
rect 20354 5187 20368 5201
rect 20786 5187 20800 5201
rect 22154 5187 22168 5201
rect 4394 5163 4408 5177
rect 22754 5163 22768 5177
rect 25514 5163 25528 5177
rect 4346 5139 4360 5153
rect 9290 5139 9304 5153
rect 9626 5139 9640 5153
rect 16490 5139 16504 5153
rect 16706 5139 16720 5153
rect 16802 5139 16816 5153
rect 17018 5139 17032 5153
rect 20762 5139 20776 5153
rect 4250 5115 4264 5129
rect 13226 5115 13240 5129
rect 13274 5115 13288 5129
rect 25898 5115 25912 5129
rect 4250 5091 4264 5105
rect 15842 5091 15856 5105
rect 15938 5091 15952 5105
rect 21110 5091 21124 5105
rect 23570 5091 23584 5105
rect 4178 5067 4192 5081
rect 6506 5067 6520 5081
rect 10106 5067 10120 5081
rect 12578 5067 12592 5081
rect 12674 5067 12688 5081
rect 13970 5067 13984 5081
rect 21002 5067 21016 5081
rect 22298 5067 22312 5081
rect 23882 5067 23896 5081
rect 26354 5067 26368 5081
rect 4106 5043 4120 5057
rect 22970 5043 22984 5057
rect 3938 5019 3952 5033
rect 8522 5019 8536 5033
rect 10226 5019 10240 5033
rect 15794 5019 15808 5033
rect 22970 5019 22984 5033
rect 3890 4995 3904 5009
rect 4082 4995 4096 5009
rect 6842 4995 6856 5009
rect 12218 4995 12232 5009
rect 12818 4995 12832 5009
rect 19922 4995 19936 5009
rect 20618 4995 20632 5009
rect 24194 4995 24208 5009
rect 26762 4995 26776 5009
rect 3818 4971 3832 4985
rect 7538 4971 7552 4985
rect 7586 4971 7600 4985
rect 26450 4971 26464 4985
rect 3794 4947 3808 4961
rect 19466 4947 19480 4961
rect 19658 4947 19672 4961
rect 19730 4947 19744 4961
rect 19898 4947 19912 4961
rect 20474 4947 20488 4961
rect 20714 4947 20728 4961
rect 20786 4947 20800 4961
rect 21674 4947 21688 4961
rect 21722 4947 21736 4961
rect 22610 4947 22624 4961
rect 22934 4947 22948 4961
rect 3506 4923 3520 4937
rect 10106 4923 10120 4937
rect 10970 4923 10984 4937
rect 13442 4923 13456 4937
rect 20954 4923 20968 4937
rect 21674 4923 21688 4937
rect 22322 4923 22336 4937
rect 25082 4923 25096 4937
rect 25466 4923 25480 4937
rect 3434 4899 3448 4913
rect 8618 4899 8632 4913
rect 16706 4899 16720 4913
rect 22850 4899 22864 4913
rect 3362 4875 3376 4889
rect 4850 4875 4864 4889
rect 7106 4875 7120 4889
rect 9746 4875 9760 4889
rect 18962 4875 18976 4889
rect 19226 4875 19240 4889
rect 19850 4875 19864 4889
rect 22610 4875 22624 4889
rect 23450 4875 23464 4889
rect 23786 4875 23800 4889
rect 26090 4875 26104 4889
rect 3290 4851 3304 4865
rect 8978 4851 8992 4865
rect 9074 4851 9088 4865
rect 13034 4851 13048 4865
rect 13082 4851 13096 4865
rect 20162 4851 20176 4865
rect 20498 4851 20512 4865
rect 22826 4851 22840 4865
rect 3146 4827 3160 4841
rect 25922 4827 25936 4841
rect 3098 4803 3112 4817
rect 16082 4803 16096 4817
rect 16178 4803 16192 4817
rect 20714 4803 20728 4817
rect 3050 4779 3064 4793
rect 21458 4779 21472 4793
rect 3026 4755 3040 4769
rect 19034 4755 19048 4769
rect 20834 4755 20848 4769
rect 25202 4755 25216 4769
rect 2930 4731 2944 4745
rect 8786 4731 8800 4745
rect 8930 4731 8944 4745
rect 21242 4731 21256 4745
rect 22634 4731 22648 4745
rect 23174 4731 23188 4745
rect 2906 4707 2920 4721
rect 14954 4707 14968 4721
rect 16322 4707 16336 4721
rect 16586 4707 16600 4721
rect 23210 4707 23224 4721
rect 2834 4683 2848 4697
rect 7226 4683 7240 4697
rect 24770 4683 24784 4697
rect 27122 4683 27136 4697
rect 2810 4659 2824 4673
rect 5330 4659 5344 4673
rect 5690 4659 5704 4673
rect 5882 4659 5896 4673
rect 5954 4659 5968 4673
rect 10610 4659 10624 4673
rect 12098 4659 12112 4673
rect 24962 4659 24976 4673
rect 2738 4635 2752 4649
rect 4514 4635 4528 4649
rect 5930 4635 5944 4649
rect 10250 4635 10264 4649
rect 12026 4635 12040 4649
rect 12194 4635 12208 4649
rect 12914 4635 12928 4649
rect 13826 4635 13840 4649
rect 18362 4635 18376 4649
rect 22994 4635 23008 4649
rect 23810 4635 23824 4649
rect 25610 4635 25624 4649
rect 2666 4611 2680 4625
rect 23018 4611 23032 4625
rect 23114 4611 23128 4625
rect 23498 4611 23512 4625
rect 23546 4611 23560 4625
rect 23834 4611 23848 4625
rect 24146 4611 24160 4625
rect 26858 4611 26872 4625
rect 2618 4587 2632 4601
rect 10754 4587 10768 4601
rect 24890 4587 24904 4601
rect 26786 4587 26800 4601
rect 2594 4563 2608 4577
rect 24170 4563 24184 4577
rect 25130 4563 25144 4577
rect 25178 4563 25192 4577
rect 25274 4563 25288 4577
rect 25298 4563 25312 4577
rect 25658 4563 25672 4577
rect 25682 4563 25696 4577
rect 25994 4563 26008 4577
rect 27853 4563 27867 4577
rect 2522 4539 2536 4553
rect 7850 4539 7864 4553
rect 7970 4539 7984 4553
rect 9026 4539 9040 4553
rect 9890 4539 9904 4553
rect 20378 4539 20392 4553
rect 20834 4539 20848 4553
rect 26810 4539 26824 4553
rect 2474 4515 2488 4529
rect 3530 4515 3544 4529
rect 10010 4515 10024 4529
rect 15290 4515 15304 4529
rect 24434 4515 24448 4529
rect 25322 4515 25336 4529
rect 25370 4515 25384 4529
rect 26810 4515 26824 4529
rect 27050 4515 27064 4529
rect 2402 4491 2416 4505
rect 5618 4491 5632 4505
rect 5666 4491 5680 4505
rect 8594 4491 8608 4505
rect 9674 4491 9688 4505
rect 13010 4491 13024 4505
rect 13370 4491 13384 4505
rect 17186 4491 17200 4505
rect 18410 4491 18424 4505
rect 20594 4491 20608 4505
rect 26642 4491 26656 4505
rect 2378 4467 2392 4481
rect 11426 4467 11440 4481
rect 16754 4467 16768 4481
rect 18314 4467 18328 4481
rect 26498 4467 26512 4481
rect 2330 4443 2344 4457
rect 10730 4443 10744 4457
rect 10778 4443 10792 4457
rect 13442 4443 13456 4457
rect 13490 4443 13504 4457
rect 16802 4443 16816 4457
rect 17210 4443 17224 4457
rect 21074 4443 21088 4457
rect 21314 4443 21328 4457
rect 24578 4443 24592 4457
rect 26498 4443 26512 4457
rect 26642 4443 26656 4457
rect 2306 4419 2320 4433
rect 3770 4419 3784 4433
rect 4034 4419 4048 4433
rect 7274 4419 7288 4433
rect 10562 4419 10576 4433
rect 15362 4419 15376 4433
rect 16682 4419 16696 4433
rect 23114 4419 23128 4433
rect 25130 4419 25144 4433
rect 27314 4419 27328 4433
rect 2282 4395 2296 4409
rect 14090 4395 14104 4409
rect 14186 4395 14200 4409
rect 14810 4395 14824 4409
rect 15122 4395 15136 4409
rect 24026 4395 24040 4409
rect 24386 4395 24400 4409
rect 26978 4395 26992 4409
rect 2234 4371 2248 4385
rect 4226 4371 4240 4385
rect 5282 4371 5296 4385
rect 5402 4371 5416 4385
rect 19442 4371 19456 4385
rect 19586 4371 19600 4385
rect 20210 4371 20224 4385
rect 20642 4371 20656 4385
rect 25178 4371 25192 4385
rect 2210 4347 2224 4361
rect 6578 4347 6592 4361
rect 9602 4347 9616 4361
rect 17066 4347 17080 4361
rect 18266 4347 18280 4361
rect 19322 4347 19336 4361
rect 22994 4347 23008 4361
rect 23282 4347 23296 4361
rect 24122 4347 24136 4361
rect 24338 4347 24352 4361
rect 24554 4347 24568 4361
rect 26402 4347 26416 4361
rect 2186 4323 2200 4337
rect 3866 4323 3880 4337
rect 4298 4323 4312 4337
rect 8186 4323 8200 4337
rect 12362 4323 12376 4337
rect 13850 4323 13864 4337
rect 14258 4323 14272 4337
rect 23786 4323 23800 4337
rect 24338 4323 24352 4337
rect 24494 4323 24508 4337
rect 26402 4323 26416 4337
rect 26450 4323 26464 4337
rect 2090 4299 2104 4313
rect 13322 4299 13336 4313
rect 19562 4299 19576 4313
rect 26906 4299 26920 4313
rect 2066 4275 2080 4289
rect 8570 4275 8584 4289
rect 10178 4275 10192 4289
rect 10298 4275 10312 4289
rect 26834 4275 26848 4289
rect 1994 4251 2008 4265
rect 10322 4251 10336 4265
rect 12122 4251 12136 4265
rect 12890 4251 12904 4265
rect 20054 4251 20068 4265
rect 21194 4251 21208 4265
rect 23810 4251 23824 4265
rect 26186 4251 26200 4265
rect 1970 4227 1984 4241
rect 3002 4227 3016 4241
rect 3266 4227 3280 4241
rect 8858 4227 8872 4241
rect 10634 4227 10648 4241
rect 20114 4227 20128 4241
rect 21650 4227 21664 4241
rect 25394 4227 25408 4241
rect 1946 4203 1960 4217
rect 5594 4203 5608 4217
rect 18074 4203 18088 4217
rect 21242 4203 21256 4217
rect 22898 4203 22912 4217
rect 26066 4203 26080 4217
rect 1898 4179 1912 4193
rect 23954 4179 23968 4193
rect 25394 4179 25408 4193
rect 25418 4179 25432 4193
rect 1850 4155 1864 4169
rect 3218 4155 3232 4169
rect 3698 4155 3712 4169
rect 4634 4155 4648 4169
rect 6170 4155 6184 4169
rect 7874 4155 7888 4169
rect 9146 4155 9160 4169
rect 11930 4155 11944 4169
rect 13922 4155 13936 4169
rect 18602 4155 18616 4169
rect 20138 4155 20152 4169
rect 21194 4155 21208 4169
rect 22394 4155 22408 4169
rect 22538 4155 22552 4169
rect 26042 4155 26056 4169
rect 1826 4131 1840 4145
rect 8906 4131 8920 4145
rect 11618 4131 11632 4145
rect 11858 4131 11872 4145
rect 24458 4131 24472 4145
rect 1754 4107 1768 4121
rect 2690 4107 2704 4121
rect 6098 4107 6112 4121
rect 6650 4107 6664 4121
rect 6962 4107 6976 4121
rect 8114 4107 8128 4121
rect 9482 4107 9496 4121
rect 17114 4107 17128 4121
rect 17882 4107 17896 4121
rect 18170 4107 18184 4121
rect 18674 4107 18688 4121
rect 18986 4107 19000 4121
rect 19178 4107 19192 4121
rect 19562 4107 19576 4121
rect 19802 4107 19816 4121
rect 19850 4107 19864 4121
rect 20330 4107 20344 4121
rect 20930 4107 20944 4121
rect 21482 4107 21496 4121
rect 22058 4107 22072 4121
rect 23762 4107 23776 4121
rect 1730 4083 1744 4097
rect 3386 4083 3400 4097
rect 3482 4083 3496 4097
rect 4010 4083 4024 4097
rect 4202 4083 4216 4097
rect 11210 4083 11224 4097
rect 11810 4083 11824 4097
rect 14042 4083 14056 4097
rect 15410 4083 15424 4097
rect 18242 4083 18256 4097
rect 18458 4083 18472 4097
rect 19394 4083 19408 4097
rect 19970 4083 19984 4097
rect 25346 4083 25360 4097
rect 25442 4083 25456 4097
rect 26162 4083 26176 4097
rect 1706 4059 1720 4073
rect 6530 4059 6544 4073
rect 13010 4059 13024 4073
rect 14882 4059 14896 4073
rect 15482 4059 15496 4073
rect 26666 4059 26680 4073
rect 1658 4035 1672 4049
rect 9986 4035 10000 4049
rect 10058 4035 10072 4049
rect 17690 4035 17704 4049
rect 19802 4035 19816 4049
rect 27026 4035 27040 4049
rect 1634 4011 1648 4025
rect 3218 4011 3232 4025
rect 7442 4011 7456 4025
rect 7730 4011 7744 4025
rect 7994 4011 8008 4025
rect 12698 4011 12712 4025
rect 18482 4011 18496 4025
rect 20858 4011 20872 4025
rect 21698 4011 21712 4025
rect 22706 4011 22720 4025
rect 23366 4011 23380 4025
rect 25442 4011 25456 4025
rect 27410 4011 27424 4025
rect 1610 3987 1624 4001
rect 4610 3987 4624 4001
rect 13634 3987 13648 4001
rect 18050 3987 18064 4001
rect 19970 3987 19984 4001
rect 20054 3987 20068 4001
rect 20138 3987 20152 4001
rect 25034 3987 25048 4001
rect 70 3963 84 3977
rect 8138 3963 8152 3977
rect 16994 3963 17008 3977
rect 17306 3963 17320 3977
rect 21434 3963 21448 3977
rect 22802 3963 22816 3977
rect 23306 3963 23320 3977
rect 70 3939 84 3953
rect 9410 3939 9424 3953
rect 9602 3939 9616 3953
rect 9818 3939 9832 3953
rect 9890 3939 9904 3953
rect 9914 3939 9928 3953
rect 10082 3939 10096 3953
rect 22010 3939 22024 3953
rect 26618 3939 26632 3953
rect 1610 3915 1624 3929
rect 9170 3915 9184 3929
rect 13898 3915 13912 3929
rect 14066 3915 14080 3929
rect 14138 3915 14152 3929
rect 15218 3915 15232 3929
rect 15602 3915 15616 3929
rect 15674 3915 15688 3929
rect 15722 3915 15736 3929
rect 16274 3915 16288 3929
rect 17522 3915 17536 3929
rect 20858 3915 20872 3929
rect 21002 3915 21016 3929
rect 21338 3915 21352 3929
rect 23498 3915 23512 3929
rect 1634 3891 1648 3905
rect 3554 3891 3568 3905
rect 4946 3891 4960 3905
rect 5978 3891 5992 3905
rect 9458 3891 9472 3905
rect 14690 3891 14704 3905
rect 16154 3891 16168 3905
rect 26258 3891 26272 3905
rect 1778 3867 1792 3881
rect 26666 3867 26680 3881
rect 2018 3843 2032 3857
rect 8306 3843 8320 3857
rect 9002 3843 9016 3857
rect 19682 3843 19696 3857
rect 20954 3843 20968 3857
rect 21110 3843 21124 3857
rect 21362 3843 21376 3857
rect 21938 3843 21952 3857
rect 23282 3843 23296 3857
rect 27853 3843 27867 3857
rect 2162 3819 2176 3833
rect 9242 3819 9256 3833
rect 21170 3819 21184 3833
rect 2210 3795 2224 3809
rect 3242 3795 3256 3809
rect 5426 3795 5440 3809
rect 6818 3795 6832 3809
rect 9578 3795 9592 3809
rect 13418 3795 13432 3809
rect 13898 3795 13912 3809
rect 19778 3795 19792 3809
rect 20090 3795 20104 3809
rect 21554 3795 21568 3809
rect 22634 3795 22648 3809
rect 24650 3795 24664 3809
rect 25826 3795 25840 3809
rect 2426 3771 2440 3785
rect 13586 3771 13600 3785
rect 15410 3771 15424 3785
rect 15434 3771 15448 3785
rect 16514 3771 16528 3785
rect 23402 3771 23416 3785
rect 2498 3747 2512 3761
rect 6626 3747 6640 3761
rect 7154 3747 7168 3761
rect 12002 3747 12016 3761
rect 13658 3747 13672 3761
rect 19874 3747 19888 3761
rect 21026 3747 21040 3761
rect 2570 3723 2584 3737
rect 5114 3723 5128 3737
rect 11330 3723 11344 3737
rect 11594 3723 11608 3737
rect 13802 3723 13816 3737
rect 16754 3723 16768 3737
rect 25778 3723 25792 3737
rect 2594 3699 2608 3713
rect 3602 3699 3616 3713
rect 11354 3699 11368 3713
rect 15194 3699 15208 3713
rect 22178 3699 22192 3713
rect 22346 3699 22360 3713
rect 26258 3699 26272 3713
rect 2642 3675 2656 3689
rect 23666 3675 23680 3689
rect 2690 3651 2704 3665
rect 5450 3651 5464 3665
rect 5498 3651 5512 3665
rect 9266 3651 9280 3665
rect 18146 3651 18160 3665
rect 19106 3651 19120 3665
rect 24530 3651 24544 3665
rect 25274 3651 25288 3665
rect 2858 3627 2872 3641
rect 26234 3627 26248 3641
rect 3266 3603 3280 3617
rect 4418 3603 4432 3617
rect 8114 3603 8128 3617
rect 9050 3603 9064 3617
rect 10946 3603 10960 3617
rect 13130 3603 13144 3617
rect 17522 3603 17536 3617
rect 22250 3603 22264 3617
rect 24530 3603 24544 3617
rect 24698 3603 24712 3617
rect 3314 3579 3328 3593
rect 9578 3579 9592 3593
rect 9746 3579 9760 3593
rect 12866 3579 12880 3593
rect 13058 3579 13072 3593
rect 22490 3579 22504 3593
rect 3410 3555 3424 3569
rect 20450 3555 20464 3569
rect 22934 3555 22948 3569
rect 3458 3531 3472 3545
rect 3674 3531 3688 3545
rect 24626 3531 24640 3545
rect 3578 3507 3592 3521
rect 13394 3507 13408 3521
rect 13466 3507 13480 3521
rect 16058 3507 16072 3521
rect 17450 3507 17464 3521
rect 24314 3507 24328 3521
rect 26474 3507 26488 3521
rect 3602 3483 3616 3497
rect 23426 3483 23440 3497
rect 3626 3459 3640 3473
rect 11282 3459 11296 3473
rect 11810 3459 11824 3473
rect 17498 3459 17512 3473
rect 20450 3459 20464 3473
rect 20474 3459 20488 3473
rect 3698 3435 3712 3449
rect 16874 3435 16888 3449
rect 3722 3411 3736 3425
rect 7586 3411 7600 3425
rect 7634 3411 7648 3425
rect 10826 3411 10840 3425
rect 12050 3411 12064 3425
rect 17330 3411 17344 3425
rect 3746 3387 3760 3401
rect 17162 3387 17176 3401
rect 19154 3387 19168 3401
rect 3794 3363 3808 3377
rect 10442 3363 10456 3377
rect 19010 3363 19024 3377
rect 19154 3363 19168 3377
rect 25106 3363 25120 3377
rect 3866 3339 3880 3353
rect 8954 3339 8968 3353
rect 26546 3339 26560 3353
rect 3914 3315 3928 3329
rect 5906 3315 5920 3329
rect 8714 3315 8728 3329
rect 8834 3315 8848 3329
rect 21530 3315 21544 3329
rect 21722 3315 21736 3329
rect 3986 3291 4000 3305
rect 7034 3291 7048 3305
rect 12170 3291 12184 3305
rect 12626 3291 12640 3305
rect 17378 3291 17392 3305
rect 4010 3267 4024 3281
rect 5714 3267 5728 3281
rect 8978 3267 8992 3281
rect 19070 3267 19084 3281
rect 19442 3267 19456 3281
rect 19658 3267 19672 3281
rect 20666 3267 20680 3281
rect 22442 3267 22456 3281
rect 4058 3243 4072 3257
rect 10466 3243 10480 3257
rect 23858 3243 23872 3257
rect 24098 3243 24112 3257
rect 4106 3219 4120 3233
rect 6914 3219 6928 3233
rect 10514 3219 10528 3233
rect 20594 3219 20608 3233
rect 23066 3219 23080 3233
rect 4322 3195 4336 3209
rect 6122 3195 6136 3209
rect 6194 3195 6208 3209
rect 21794 3195 21808 3209
rect 4346 3171 4360 3185
rect 6218 3171 6232 3185
rect 13730 3171 13744 3185
rect 19754 3171 19768 3185
rect 21794 3171 21808 3185
rect 21818 3171 21832 3185
rect 4418 3147 4432 3161
rect 12602 3147 12616 3161
rect 14234 3147 14248 3161
rect 14930 3147 14944 3161
rect 24026 3147 24040 3161
rect 4442 3123 4456 3137
rect 13514 3123 13528 3137
rect 16874 3123 16888 3137
rect 16898 3123 16912 3137
rect 4538 3099 4552 3113
rect 6314 3099 6328 3113
rect 6698 3099 6712 3113
rect 8642 3099 8656 3113
rect 13034 3099 13048 3113
rect 20258 3099 20272 3113
rect 26690 3099 26704 3113
rect 4562 3075 4576 3089
rect 6386 3075 6400 3089
rect 6986 3075 7000 3089
rect 7490 3075 7504 3089
rect 8738 3075 8752 3089
rect 8762 3075 8776 3089
rect 17474 3075 17488 3089
rect 17666 3075 17680 3089
rect 19130 3075 19144 3089
rect 19346 3075 19360 3089
rect 22514 3075 22528 3089
rect 4658 3051 4672 3065
rect 10586 3051 10600 3065
rect 12962 3051 12976 3065
rect 16946 3051 16960 3065
rect 17402 3051 17416 3065
rect 19994 3051 20008 3065
rect 25226 3051 25240 3065
rect 4730 3027 4744 3041
rect 7658 3027 7672 3041
rect 11306 3027 11320 3041
rect 23906 3027 23920 3041
rect 4754 3003 4768 3017
rect 7730 3003 7744 3017
rect 26522 3003 26536 3017
rect 4826 2979 4840 2993
rect 6482 2979 6496 2993
rect 22874 2979 22888 2993
rect 23690 2979 23704 2993
rect 5114 2955 5128 2969
rect 25154 2955 25168 2969
rect 5186 2931 5200 2945
rect 12146 2931 12160 2945
rect 12194 2931 12208 2945
rect 12290 2931 12304 2945
rect 12434 2931 12448 2945
rect 12530 2931 12544 2945
rect 12722 2931 12736 2945
rect 18866 2931 18880 2945
rect 19130 2931 19144 2945
rect 19610 2931 19624 2945
rect 5522 2907 5536 2921
rect 6674 2907 6688 2921
rect 25514 2907 25528 2921
rect 5546 2883 5560 2897
rect 16826 2883 16840 2897
rect 16946 2883 16960 2897
rect 17354 2883 17368 2897
rect 5714 2859 5728 2873
rect 16418 2859 16432 2873
rect 16778 2859 16792 2873
rect 20522 2859 20536 2873
rect 24074 2859 24088 2873
rect 26738 2859 26752 2873
rect 5810 2835 5824 2849
rect 8018 2835 8032 2849
rect 13202 2835 13216 2849
rect 20306 2835 20320 2849
rect 26738 2835 26752 2849
rect 26954 2835 26968 2849
rect 6002 2811 6016 2825
rect 14282 2811 14296 2825
rect 15026 2811 15040 2825
rect 16922 2811 16936 2825
rect 17426 2811 17440 2825
rect 19514 2811 19528 2825
rect 21602 2811 21616 2825
rect 6026 2787 6040 2801
rect 19514 2787 19528 2801
rect 20306 2787 20320 2801
rect 20354 2787 20368 2801
rect 6074 2763 6088 2777
rect 8066 2763 8080 2777
rect 8186 2763 8200 2777
rect 23174 2763 23188 2777
rect 6218 2739 6232 2753
rect 7178 2739 7192 2753
rect 7778 2739 7792 2753
rect 15386 2739 15400 2753
rect 17282 2739 17296 2753
rect 18386 2739 18400 2753
rect 21074 2739 21088 2753
rect 21218 2739 21232 2753
rect 23330 2739 23344 2753
rect 23354 2739 23368 2753
rect 6458 2715 6472 2729
rect 14138 2715 14152 2729
rect 16922 2715 16936 2729
rect 17330 2715 17344 2729
rect 23330 2715 23344 2729
rect 23618 2715 23632 2729
rect 6530 2691 6544 2705
rect 16346 2691 16360 2705
rect 19250 2691 19264 2705
rect 23522 2691 23536 2705
rect 6674 2667 6688 2681
rect 16562 2667 16576 2681
rect 19730 2667 19744 2681
rect 6722 2643 6736 2657
rect 8522 2643 8536 2657
rect 14714 2643 14728 2657
rect 6770 2619 6784 2633
rect 12650 2619 12664 2633
rect 17978 2619 17992 2633
rect 7082 2595 7096 2609
rect 9098 2595 9112 2609
rect 10370 2595 10384 2609
rect 13106 2595 13120 2609
rect 13154 2595 13168 2609
rect 23978 2595 23992 2609
rect 7106 2571 7120 2585
rect 7130 2571 7144 2585
rect 7202 2571 7216 2585
rect 13346 2571 13360 2585
rect 16130 2571 16144 2585
rect 23042 2571 23056 2585
rect 26882 2571 26896 2585
rect 7706 2547 7720 2561
rect 9530 2547 9544 2561
rect 11546 2547 11560 2561
rect 23234 2547 23248 2561
rect 26306 2547 26320 2561
rect 7754 2523 7768 2537
rect 27410 2523 27424 2537
rect 7802 2499 7816 2513
rect 22682 2499 22696 2513
rect 7850 2475 7864 2489
rect 25802 2475 25816 2489
rect 7970 2451 7984 2465
rect 8402 2451 8416 2465
rect 8642 2451 8656 2465
rect 11234 2451 11248 2465
rect 11906 2451 11920 2465
rect 12242 2451 12256 2465
rect 17762 2451 17776 2465
rect 8018 2427 8032 2441
rect 10946 2427 10960 2441
rect 19946 2427 19960 2441
rect 8234 2403 8248 2417
rect 23258 2403 23272 2417
rect 24362 2403 24376 2417
rect 8258 2379 8272 2393
rect 9554 2379 9568 2393
rect 11570 2379 11584 2393
rect 23594 2379 23608 2393
rect 24362 2379 24376 2393
rect 24602 2379 24616 2393
rect 8954 2355 8968 2369
rect 9218 2355 9232 2369
rect 12482 2355 12496 2369
rect 12770 2355 12784 2369
rect 15866 2355 15880 2369
rect 9050 2331 9064 2345
rect 9698 2331 9712 2345
rect 24722 2331 24736 2345
rect 9218 2307 9232 2321
rect 13778 2307 13792 2321
rect 9242 2283 9256 2297
rect 9290 2283 9304 2297
rect 9362 2283 9376 2297
rect 13610 2283 13624 2297
rect 13778 2283 13792 2297
rect 24674 2283 24688 2297
rect 25586 2283 25600 2297
rect 9410 2259 9424 2273
rect 11138 2259 11152 2273
rect 11162 2259 11176 2273
rect 20978 2259 20992 2273
rect 24242 2259 24256 2273
rect 26522 2259 26536 2273
rect 9458 2235 9472 2249
rect 9794 2235 9808 2249
rect 10178 2235 10192 2249
rect 12458 2235 12472 2249
rect 12794 2235 12808 2249
rect 13562 2235 13576 2249
rect 13610 2235 13624 2249
rect 21746 2235 21760 2249
rect 26210 2235 26224 2249
rect 10346 2211 10360 2225
rect 14402 2211 14416 2225
rect 10394 2187 10408 2201
rect 24722 2187 24736 2201
rect 10490 2163 10504 2177
rect 21290 2163 21304 2177
rect 10562 2139 10576 2153
rect 10610 2139 10624 2153
rect 10658 2139 10672 2153
rect 17618 2139 17632 2153
rect 25298 2139 25312 2153
rect 10898 2115 10912 2129
rect 18770 2115 18784 2129
rect 10970 2091 10984 2105
rect 11066 2091 11080 2105
rect 11114 2091 11128 2105
rect 21458 2091 21472 2105
rect 11138 2067 11152 2081
rect 12074 2067 12088 2081
rect 16250 2067 16264 2081
rect 18338 2067 18352 2081
rect 19898 2067 19912 2081
rect 22874 2067 22888 2081
rect 27338 2067 27352 2081
rect 13106 2043 13120 2057
rect 18890 2043 18904 2057
rect 20882 2043 20896 2057
rect 13250 2019 13264 2033
rect 22514 2019 22528 2033
rect 13466 1995 13480 2009
rect 21986 1995 22000 2009
rect 25754 1995 25768 2009
rect 27434 1995 27448 2009
rect 27853 1995 27867 2009
rect 13538 1971 13552 1985
rect 15050 1971 15064 1985
rect 27410 1971 27424 1985
rect 27853 1971 27867 1985
rect 16418 1138 16432 1152
rect 23378 1138 23392 1152
rect 15866 1114 15880 1128
rect 18842 1114 18856 1128
rect 14570 1090 14584 1104
rect 23954 1090 23968 1104
rect 13202 1066 13216 1080
rect 22922 1066 22936 1080
rect 13154 1042 13168 1056
rect 14594 1042 14608 1056
rect 14786 1042 14800 1056
rect 23426 1042 23440 1056
rect 24482 1042 24496 1056
rect 12674 1018 12688 1032
rect 23738 1018 23752 1032
rect 12314 994 12328 1008
rect 18098 994 18112 1008
rect 11042 970 11056 984
rect 17114 970 17128 984
rect 10922 946 10936 960
rect 13850 946 13864 960
rect 14450 946 14464 960
rect 21122 946 21136 960
rect 10850 922 10864 936
rect 23906 922 23920 936
rect 10706 898 10720 912
rect 19274 898 19288 912
rect 10010 874 10024 888
rect 18194 874 18208 888
rect 9986 850 10000 864
rect 13730 850 13744 864
rect 14354 850 14368 864
rect 16610 850 16624 864
rect 9938 826 9952 840
rect 24122 826 24136 840
rect 9506 802 9520 816
rect 21626 802 21640 816
rect 22562 802 22576 816
rect 23642 802 23656 816
rect 9122 778 9136 792
rect 22778 778 22792 792
rect 8786 754 8800 768
rect 14930 754 14944 768
rect 19418 754 19432 768
rect 20210 754 20224 768
rect 20690 754 20704 768
rect 22466 754 22480 768
rect 26882 754 26896 768
rect 7322 730 7336 744
rect 15698 730 15712 744
rect 15746 730 15760 744
rect 16442 730 16456 744
rect 20162 730 20176 744
rect 24602 730 24616 744
rect 7226 706 7240 720
rect 13802 706 13816 720
rect 14042 706 14056 720
rect 17690 706 17704 720
rect 18002 706 18016 720
rect 20498 706 20512 720
rect 20618 706 20632 720
rect 22202 706 22216 720
rect 27853 706 27867 720
rect 6962 682 6976 696
rect 16850 682 16864 696
rect 17906 682 17920 696
rect 23690 682 23704 696
rect 6410 658 6424 672
rect 24002 658 24016 672
rect 6242 634 6256 648
rect 12338 634 12352 648
rect 12386 634 12400 648
rect 17498 634 17512 648
rect 17738 634 17752 648
rect 26690 634 26704 648
rect 6098 610 6112 624
rect 11186 610 11200 624
rect 11234 610 11248 624
rect 26450 610 26464 624
rect 5978 586 5992 600
rect 8714 586 8728 600
rect 15506 586 15520 600
rect 20042 586 20056 600
rect 20402 586 20416 600
rect 24242 586 24256 600
rect 5930 562 5944 576
rect 7682 562 7696 576
rect 8282 562 8296 576
rect 9818 562 9832 576
rect 9866 562 9880 576
rect 15074 562 15088 576
rect 15146 562 15160 576
rect 23186 562 23200 576
rect 26930 562 26944 576
rect 5834 538 5848 552
rect 19754 538 19768 552
rect 5474 514 5488 528
rect 6746 514 6760 528
rect 6938 514 6952 528
rect 20978 514 20992 528
rect 4946 490 4960 504
rect 6026 490 6040 504
rect 6074 490 6088 504
rect 7418 490 7432 504
rect 7466 490 7480 504
rect 20090 490 20104 504
rect 4922 466 4936 480
rect 20546 466 20560 480
rect 4874 442 4888 456
rect 23714 442 23728 456
rect 4586 418 4600 432
rect 20426 418 20440 432
rect 4466 394 4480 408
rect 20378 394 20392 408
rect 24266 394 24280 408
rect 4202 370 4216 384
rect 14306 370 14320 384
rect 14522 370 14536 384
rect 17066 370 17080 384
rect 4154 346 4168 360
rect 10034 346 10048 360
rect 10634 346 10648 360
rect 10682 346 10696 360
rect 10754 346 10768 360
rect 15170 346 15184 360
rect 15314 346 15328 360
rect 15554 346 15568 360
rect 15626 346 15640 360
rect 26954 346 26968 360
rect 3674 322 3688 336
rect 4298 322 4312 336
rect 10274 322 10288 336
rect 22106 322 22120 336
rect 3650 298 3664 312
rect 21002 298 21016 312
rect 3530 274 3544 288
rect 16994 274 17008 288
rect 2858 250 2872 264
rect 14618 250 14632 264
rect 14834 250 14848 264
rect 26594 250 26608 264
rect 2738 226 2752 240
rect 26642 226 26656 240
rect 2522 202 2536 216
rect 26618 202 26632 216
rect 2474 178 2488 192
rect 8426 178 8440 192
rect 8546 178 8560 192
rect 16802 178 16816 192
rect 1802 154 1816 168
rect 7610 154 7624 168
rect 8030 154 8044 168
rect 22706 154 22720 168
rect 1682 130 1696 144
rect 11018 130 11032 144
rect 11090 130 11104 144
rect 20738 130 20752 144
rect 70 106 84 120
rect 19850 106 19864 120
rect 70 82 84 96
rect 2354 82 2368 96
rect 2402 82 2416 96
rect 18434 82 18448 96
rect 2618 58 2632 72
rect 27853 58 27867 72
rect 4130 34 4144 48
rect 8066 34 8080 48
rect 8378 34 8392 48
rect 24074 34 24088 48
rect 26930 34 26944 48
rect 27853 34 27867 48
rect 11954 10 11968 24
rect 26930 10 26944 24
rect 26954 10 26968 24
rect 27853 10 27867 24
<< metal2 >>
rect 0 8061 70 8073
rect 0 8037 70 8049
rect 123 7930 323 8300
rect 339 7930 351 8300
rect 363 7930 375 8300
rect 387 7930 399 8300
rect 411 7930 423 8300
rect 1707 7930 1719 8084
rect 2139 7930 2151 8012
rect 2211 7930 2223 8108
rect 2427 8002 2439 8300
rect 2463 8098 2475 8300
rect 2955 7930 2967 8084
rect 4083 7930 4095 8132
rect 4155 7978 4167 8300
rect 4191 8122 4203 8300
rect 5055 8122 5067 8300
rect 5991 8170 6003 8300
rect 6975 8170 6987 8300
rect 5992 8156 6010 8170
rect 6976 8156 6994 8170
rect 4731 7930 4743 8108
rect 5523 7930 5535 8108
rect 5979 7930 5991 8156
rect 6579 7930 6591 7988
rect 6675 7930 6687 7988
rect 6963 7930 6975 8156
rect 7647 8146 7659 8300
rect 9339 8146 9351 8300
rect 9951 8194 9963 8300
rect 9952 8180 9970 8194
rect 6987 7930 6999 7964
rect 8475 7930 8487 7964
rect 9819 7930 9831 8156
rect 9939 7930 9951 8180
rect 10239 7978 10251 8300
rect 11931 8194 11943 8300
rect 11067 7930 11079 8036
rect 11643 7930 11655 8036
rect 12795 7978 12807 8300
rect 12831 8098 12843 8300
rect 12915 7930 12927 8084
rect 13635 7930 13647 8012
rect 14523 7978 14535 8300
rect 14139 7930 14151 7964
rect 14667 7930 14679 8204
rect 14811 7930 14823 8228
rect 15375 7954 15387 8300
rect 15951 8290 15963 8300
rect 15952 8276 15970 8290
rect 15603 7930 15615 8252
rect 15939 7930 15951 8276
rect 16887 7954 16899 8300
rect 17103 8242 17115 8300
rect 18783 8290 18795 8300
rect 16888 7940 16906 7954
rect 16371 7930 16383 7940
rect 16875 7930 16887 7940
rect 18099 7930 18111 7940
rect 18675 7930 18687 8228
rect 18807 8026 18819 8300
rect 18915 7930 18927 8276
rect 19251 7930 19263 7964
rect 19611 7930 19623 8012
rect 20223 7978 20235 8300
rect 20511 8266 20523 8300
rect 21363 8170 21375 8300
rect 22215 8050 22227 8300
rect 23067 8050 23079 8300
rect 23919 8098 23931 8300
rect 20224 7964 20242 7978
rect 20211 7930 20223 7964
rect 22347 7930 22359 8036
rect 24555 7930 24567 8084
rect 24771 8002 24783 8300
rect 25623 8218 25635 8300
rect 26115 7930 26127 8060
rect 27051 7930 27063 8132
rect 27243 7930 27255 8180
rect 27303 8146 27315 8300
rect 27411 7930 27423 8132
rect 27435 7978 27447 8228
rect 27555 8178 27756 8300
rect 27483 8026 27495 8108
rect 27459 8002 27471 8012
rect 27507 7954 27519 8036
rect 27531 7954 27543 8084
rect 27555 7930 27755 8178
rect 27867 8037 27937 8049
rect 27867 8013 27937 8025
rect 27867 7989 27937 8001
rect 27867 7965 27937 7977
rect 27867 7941 27937 7953
rect 0 3964 70 3976
rect 0 3940 70 3952
rect 123 1961 323 7131
rect 339 1961 351 7131
rect 363 1961 375 7131
rect 387 1961 399 7131
rect 411 1961 423 7131
rect 1611 4001 1623 7131
rect 1635 4025 1647 7131
rect 1659 4049 1671 7131
rect 1707 4073 1719 7131
rect 1731 4097 1743 7131
rect 1755 4121 1767 7131
rect 1611 1961 1623 3915
rect 1635 1961 1647 3891
rect 1779 3881 1791 7131
rect 1827 4145 1839 7131
rect 1851 4169 1863 7131
rect 1899 4193 1911 7131
rect 1947 4217 1959 7131
rect 1971 4241 1983 7131
rect 1995 4265 2007 7131
rect 2019 3857 2031 7131
rect 2067 4289 2079 7131
rect 2091 4313 2103 7131
rect 2187 4337 2199 7131
rect 2211 4361 2223 7131
rect 2235 4385 2247 7131
rect 2283 4409 2295 7131
rect 2307 4433 2319 7131
rect 2331 4457 2343 7131
rect 2379 4481 2391 7131
rect 2403 4505 2415 7131
rect 2163 1961 2175 3819
rect 2211 1961 2223 3795
rect 2427 3785 2439 7131
rect 2475 4529 2487 7131
rect 2523 4553 2535 7131
rect 2595 4577 2607 7131
rect 2619 4601 2631 7131
rect 2499 1961 2511 3747
rect 2571 1961 2583 3723
rect 2595 1961 2607 3699
rect 2643 3689 2655 7131
rect 2667 1961 2679 4611
rect 2691 4121 2703 7131
rect 2739 4649 2751 7131
rect 2811 4673 2823 7131
rect 2835 4697 2847 7131
rect 2691 1961 2703 3651
rect 2859 3641 2871 7131
rect 2907 4721 2919 7131
rect 2931 4745 2943 7131
rect 3003 4241 3015 7131
rect 3027 4769 3039 7131
rect 3051 4793 3063 7131
rect 3099 4817 3111 7131
rect 3147 4841 3159 7131
rect 3219 4169 3231 7131
rect 3219 1961 3231 4011
rect 3243 3809 3255 7131
rect 3267 4241 3279 7131
rect 3291 4865 3303 7131
rect 3267 1961 3279 3603
rect 3315 3593 3327 7131
rect 3363 4889 3375 7131
rect 3387 4097 3399 7131
rect 3435 4913 3447 7131
rect 3483 4097 3495 7131
rect 3507 4937 3519 7131
rect 3531 4529 3543 7131
rect 3411 1961 3423 3555
rect 3459 1961 3471 3531
rect 3555 1961 3567 3891
rect 3579 3521 3591 7131
rect 3603 3713 3615 7131
rect 3603 1961 3615 3483
rect 3627 3473 3639 7131
rect 3675 3545 3687 7131
rect 3699 4169 3711 7131
rect 3699 1961 3711 3435
rect 3723 3425 3735 7131
rect 3771 4433 3783 7131
rect 3795 4961 3807 7131
rect 3819 4985 3831 7131
rect 3867 4337 3879 7131
rect 3891 5009 3903 7131
rect 3939 5033 3951 7131
rect 4011 4097 4023 7131
rect 4035 4433 4047 7131
rect 4083 5009 4095 7131
rect 4107 5057 4119 7131
rect 4179 5081 4191 7131
rect 4203 4097 4215 7131
rect 4251 5129 4263 7131
rect 3747 1961 3759 3387
rect 3795 1961 3807 3363
rect 3867 1961 3879 3339
rect 3915 1961 3927 3315
rect 3987 1961 3999 3291
rect 4011 1961 4023 3267
rect 4059 1961 4071 3243
rect 4107 1961 4119 3219
rect 4227 1961 4239 4371
rect 4251 1961 4263 5091
rect 4299 4337 4311 7131
rect 4323 3209 4335 7131
rect 4347 5153 4359 7131
rect 4395 5177 4407 7131
rect 4419 3617 4431 7131
rect 4347 1961 4359 3171
rect 4419 1961 4431 3147
rect 4443 3137 4455 7131
rect 4491 5201 4503 7131
rect 4515 4649 4527 7131
rect 4563 5225 4575 7131
rect 4611 4001 4623 7131
rect 4635 5249 4647 7131
rect 4659 5273 4671 7131
rect 4707 5321 4719 7131
rect 4731 5345 4743 7131
rect 4779 5393 4791 7131
rect 4539 1961 4551 3099
rect 4563 1961 4575 3075
rect 4635 1961 4647 4155
rect 4659 1961 4671 3051
rect 4683 1961 4695 5283
rect 4731 1961 4743 3027
rect 4755 1961 4767 3003
rect 4779 1961 4791 5355
rect 4827 5273 4839 7131
rect 4851 5417 4863 7131
rect 4875 5273 4887 7131
rect 4923 5441 4935 7131
rect 4827 1961 4839 2979
rect 4851 1961 4863 4875
rect 4947 3905 4959 7131
rect 4995 5489 5007 7131
rect 5043 5513 5055 7131
rect 5067 5537 5079 7131
rect 4995 1961 5007 5451
rect 5115 3737 5127 7131
rect 5163 5561 5175 7131
rect 5115 1961 5127 2955
rect 5187 2945 5199 7131
rect 5211 5537 5223 7131
rect 5235 5585 5247 7131
rect 5283 4385 5295 7131
rect 5331 4673 5343 7131
rect 5403 4385 5415 7131
rect 5427 3809 5439 7131
rect 5451 3665 5463 7131
rect 5499 3665 5511 7131
rect 5523 1961 5535 2907
rect 5547 2897 5559 7131
rect 5595 4217 5607 7131
rect 5619 4505 5631 7131
rect 5643 5609 5655 7131
rect 5691 5633 5703 7131
rect 5715 5657 5727 7131
rect 5739 5705 5751 7131
rect 5667 1961 5679 4491
rect 5691 1961 5703 4659
rect 5715 3281 5727 5619
rect 5715 1961 5727 2859
rect 5739 1961 5751 5667
rect 5763 5633 5775 7131
rect 5811 5753 5823 7131
rect 5859 5777 5871 7131
rect 5787 1961 5799 5715
rect 5811 1961 5823 2835
rect 5883 1961 5895 4659
rect 5931 4649 5943 7131
rect 5955 4673 5967 7131
rect 5979 3905 5991 7131
rect 6003 5345 6015 7131
rect 5907 1961 5919 3315
rect 6003 1961 6015 2811
rect 6027 2801 6039 7131
rect 6075 2777 6087 7131
rect 6099 4121 6111 7131
rect 6123 5801 6135 7131
rect 6171 5825 6183 7131
rect 6195 5201 6207 7131
rect 6219 5849 6231 7131
rect 6267 5825 6279 7131
rect 6291 5873 6303 7131
rect 6315 5897 6327 7131
rect 6339 5921 6351 7131
rect 6363 5945 6375 7131
rect 6411 5969 6423 7131
rect 6123 1961 6135 3195
rect 6171 1961 6183 4155
rect 6195 1961 6207 3195
rect 6219 3185 6231 5811
rect 6219 1961 6231 2739
rect 6315 1961 6327 3099
rect 6339 1961 6351 5883
rect 6387 1961 6399 3075
rect 6459 2729 6471 7131
rect 6483 1961 6495 2979
rect 6507 1961 6519 5067
rect 6531 4073 6543 7131
rect 6555 5993 6567 7131
rect 6579 6017 6591 7131
rect 6603 6041 6615 7131
rect 6651 6065 6663 7131
rect 6531 1961 6543 2691
rect 6579 1961 6591 4347
rect 6603 1961 6615 5475
rect 6627 1961 6639 3747
rect 6651 1961 6663 4107
rect 6675 2921 6687 7131
rect 6699 6089 6711 7131
rect 6747 6017 6759 7131
rect 6771 6113 6783 7131
rect 6819 6137 6831 7131
rect 6867 6185 6879 7131
rect 6699 3113 6711 6003
rect 6675 1961 6687 2667
rect 6723 1961 6735 2643
rect 6771 1961 6783 2619
rect 6819 1961 6831 3795
rect 6843 1961 6855 4995
rect 6867 1961 6879 6147
rect 6891 5705 6903 7131
rect 6915 6209 6927 7131
rect 6963 4121 6975 7131
rect 6915 1961 6927 3219
rect 6987 3089 6999 7131
rect 7011 1961 7023 6219
rect 7035 6113 7047 7131
rect 7083 6281 7095 7131
rect 7035 1961 7047 3291
rect 7059 1961 7071 6243
rect 7107 4889 7119 7131
rect 7083 1961 7095 2595
rect 7131 2585 7143 6051
rect 7155 5657 7167 7131
rect 7107 1961 7119 2571
rect 7155 1961 7167 3747
rect 7179 1961 7191 2739
rect 7203 2585 7215 7131
rect 7227 4697 7239 7131
rect 7251 5513 7263 7131
rect 7299 6305 7311 7131
rect 7323 6329 7335 7131
rect 7371 6353 7383 7131
rect 7419 6377 7431 7131
rect 7275 1961 7287 4419
rect 7299 1961 7311 5499
rect 7371 1961 7383 5859
rect 7395 1961 7407 5763
rect 7443 4025 7455 7131
rect 7467 6401 7479 7131
rect 7515 6449 7527 7131
rect 7491 1961 7503 3075
rect 7515 1961 7527 6411
rect 7539 4985 7551 7131
rect 7563 1961 7575 6459
rect 7587 4985 7599 7131
rect 7635 3425 7647 7131
rect 7659 6497 7671 7131
rect 7683 6521 7695 7131
rect 7731 4025 7743 7131
rect 7755 6545 7767 7131
rect 7587 1961 7599 3411
rect 7659 1961 7671 3027
rect 7707 1961 7719 2547
rect 7731 1961 7743 3003
rect 7779 2753 7791 7131
rect 7803 5729 7815 7131
rect 7851 4553 7863 7131
rect 7875 4169 7887 7131
rect 7923 6329 7935 7131
rect 7755 1961 7767 2523
rect 7803 1961 7815 2499
rect 7851 1961 7863 2475
rect 7923 1961 7935 5715
rect 7947 1961 7959 5907
rect 7971 4553 7983 7131
rect 7995 4025 8007 7131
rect 8019 2849 8031 7131
rect 7971 1961 7983 2451
rect 8019 1961 8031 2427
rect 8043 1961 8055 6315
rect 8067 5441 8079 7131
rect 8091 5705 8103 7131
rect 8115 4121 8127 7131
rect 8139 6569 8151 7131
rect 8187 4337 8199 7131
rect 8211 6593 8223 7131
rect 8235 6617 8247 7131
rect 8283 6641 8295 7131
rect 8307 5513 8319 7131
rect 8331 6689 8343 7131
rect 8067 1961 8079 2763
rect 8115 1961 8127 3603
rect 8139 1961 8151 3963
rect 8187 1961 8199 2763
rect 8235 1961 8247 2403
rect 8259 1961 8271 2379
rect 8307 1961 8319 3843
rect 8331 1961 8343 6651
rect 8379 6569 8391 7131
rect 8403 2465 8415 7131
rect 8427 6569 8439 7131
rect 8475 6665 8487 7131
rect 8499 1961 8511 6051
rect 8523 5033 8535 7131
rect 8547 6665 8559 7131
rect 8571 4289 8583 7131
rect 8619 4913 8631 7131
rect 8523 1961 8535 2643
rect 8595 1961 8607 4491
rect 8643 3113 8655 7131
rect 8667 6329 8679 7131
rect 8715 3329 8727 7131
rect 8739 5657 8751 7131
rect 8763 3089 8775 7131
rect 8787 4745 8799 7131
rect 8835 5609 8847 7131
rect 8859 5297 8871 7131
rect 8883 6329 8895 7131
rect 8643 1961 8655 2451
rect 8739 1961 8751 3075
rect 8835 1961 8847 3315
rect 8859 1961 8871 4227
rect 8883 1961 8895 5955
rect 8931 4745 8943 7131
rect 8907 1961 8919 4131
rect 8955 3353 8967 7131
rect 8979 4865 8991 7131
rect 9027 4553 9039 7131
rect 8955 1961 8967 2355
rect 8979 1961 8991 3267
rect 9003 1961 9015 3843
rect 9051 3617 9063 7131
rect 9075 5417 9087 7131
rect 9123 5273 9135 7131
rect 9051 1961 9063 2331
rect 9075 1961 9087 4851
rect 9147 4169 9159 7131
rect 9171 5273 9183 7131
rect 9099 1961 9111 2595
rect 9171 1961 9183 3915
rect 9195 1961 9207 5283
rect 9219 2369 9231 7131
rect 9243 3833 9255 7131
rect 9267 5609 9279 7131
rect 9315 6713 9327 7131
rect 9339 6737 9351 7131
rect 9363 6353 9375 7131
rect 9219 1961 9231 2307
rect 9243 1961 9255 2283
rect 9267 1961 9279 3651
rect 9291 2297 9303 5139
rect 9315 1961 9327 5835
rect 9387 5417 9399 7131
rect 9339 1961 9351 5259
rect 9411 3953 9423 7131
rect 9363 1961 9375 2283
rect 9411 1961 9423 2259
rect 9435 1961 9447 5331
rect 9459 3905 9471 7131
rect 9483 4121 9495 7131
rect 9507 5753 9519 7131
rect 9555 5729 9567 7131
rect 9579 3809 9591 7131
rect 9603 4361 9615 7131
rect 9627 5153 9639 7131
rect 9459 1961 9471 2235
rect 9531 1961 9543 2547
rect 9555 1961 9567 2379
rect 9579 1961 9591 3579
rect 9603 1961 9615 3939
rect 9651 1961 9663 5691
rect 9675 5273 9687 7131
rect 9699 6449 9711 7131
rect 9723 5849 9735 7131
rect 9747 4889 9759 7131
rect 9771 6761 9783 7131
rect 9675 1961 9687 4491
rect 9699 1961 9711 2331
rect 9747 1961 9759 3579
rect 9771 1961 9783 6675
rect 9795 2249 9807 5811
rect 9819 3953 9831 7131
rect 9867 6353 9879 7131
rect 9891 4553 9903 7131
rect 9915 3953 9927 6531
rect 9987 4049 9999 7131
rect 10011 4529 10023 7131
rect 10035 6689 10047 7131
rect 9891 1961 9903 3939
rect 10059 1961 10071 4035
rect 10083 3953 10095 7131
rect 10107 5081 10119 7131
rect 10131 6785 10143 7131
rect 10107 1961 10119 4923
rect 10131 1961 10143 5739
rect 10179 4289 10191 7131
rect 10227 6185 10239 7131
rect 10179 1961 10191 2235
rect 10227 1961 10239 5019
rect 10251 1961 10263 4635
rect 10299 4289 10311 7131
rect 10323 6809 10335 7131
rect 10323 1961 10335 4251
rect 10347 2225 10359 7131
rect 10371 6833 10383 7131
rect 10371 1961 10383 2595
rect 10395 2201 10407 7131
rect 10443 6065 10455 7131
rect 10467 5993 10479 7131
rect 10443 1961 10455 3363
rect 10467 1961 10479 3243
rect 10491 2177 10503 7131
rect 10539 5945 10551 7131
rect 10563 4433 10575 7131
rect 10587 5945 10599 7131
rect 10515 1961 10527 3219
rect 10563 1961 10575 2139
rect 10587 1961 10599 3051
rect 10611 2153 10623 4659
rect 10635 4241 10647 7131
rect 10659 2153 10671 7131
rect 10683 6857 10695 7131
rect 10731 4457 10743 7131
rect 10755 4601 10767 7131
rect 10779 4457 10791 7131
rect 10827 6881 10839 7131
rect 10851 6545 10863 7131
rect 10899 5945 10911 7131
rect 10803 1961 10815 5931
rect 10947 3617 10959 7131
rect 10971 4937 10983 7131
rect 11019 5249 11031 7131
rect 10827 1961 10839 3411
rect 10899 1961 10911 2115
rect 10947 1961 10959 2427
rect 11067 2105 11079 7131
rect 11115 2105 11127 7131
rect 11139 2273 11151 7131
rect 11163 6905 11175 7131
rect 11211 4097 11223 7131
rect 11235 2465 11247 7131
rect 11259 6233 11271 7131
rect 10971 1961 10983 2091
rect 11139 1961 11151 2067
rect 11163 1961 11175 2259
rect 11283 1961 11295 3459
rect 11307 3041 11319 7131
rect 11331 3737 11343 7131
rect 11355 3713 11367 7131
rect 11379 6233 11391 7131
rect 11427 4481 11439 7131
rect 11451 5249 11463 7131
rect 11499 6281 11511 7131
rect 11547 2561 11559 7131
rect 11571 2393 11583 7131
rect 11595 3737 11607 7131
rect 11619 4145 11631 7131
rect 11691 6665 11703 7131
rect 11715 5225 11727 7131
rect 11763 5225 11775 7131
rect 11811 4097 11823 7131
rect 11835 5729 11847 7131
rect 11859 4145 11871 7131
rect 11811 1961 11823 3459
rect 11907 2465 11919 7131
rect 11931 4169 11943 7131
rect 11955 6929 11967 7131
rect 11955 1961 11967 6219
rect 12003 5441 12015 7131
rect 12027 5921 12039 7131
rect 12051 6233 12063 7131
rect 12099 6953 12111 7131
rect 12003 1961 12015 3747
rect 12027 1961 12039 4635
rect 12051 1961 12063 3411
rect 12075 2081 12087 6219
rect 12123 5897 12135 7131
rect 12147 6233 12159 7131
rect 12099 1961 12111 4659
rect 12123 1961 12135 4251
rect 12171 3305 12183 6939
rect 12195 4649 12207 7131
rect 12219 5009 12231 7131
rect 12267 5729 12279 7131
rect 12291 2945 12303 6483
rect 12315 6233 12327 7131
rect 12363 4337 12375 7131
rect 12435 6137 12447 7131
rect 12147 1961 12159 2931
rect 12195 1961 12207 2931
rect 12243 1961 12255 2451
rect 12435 1961 12447 2931
rect 12459 2249 12471 7131
rect 12507 5729 12519 7131
rect 12531 2945 12543 6435
rect 12555 6137 12567 7131
rect 12579 6953 12591 7131
rect 12483 1961 12495 2355
rect 12555 1961 12567 5235
rect 12579 1961 12591 5067
rect 12603 3161 12615 7131
rect 12627 6977 12639 7131
rect 12627 1961 12639 3291
rect 12651 2633 12663 6123
rect 12675 5081 12687 7131
rect 12699 4025 12711 7131
rect 12723 6137 12735 7131
rect 12723 1961 12735 2931
rect 12771 2369 12783 7131
rect 12795 5777 12807 7131
rect 12819 7001 12831 7131
rect 12867 7025 12879 7131
rect 12987 7001 12999 7131
rect 12795 1961 12807 2235
rect 12819 1961 12831 4995
rect 12843 1961 12855 5763
rect 12867 3593 12879 6987
rect 12891 1961 12903 4251
rect 12915 1961 12927 4635
rect 13011 4505 13023 7131
rect 13035 4865 13047 7131
rect 13083 4865 13095 7131
rect 12963 1961 12975 3051
rect 13011 1961 13023 4059
rect 13035 1961 13047 3099
rect 13059 1961 13071 3579
rect 13107 2609 13119 7131
rect 13107 1961 13119 2043
rect 13131 1961 13143 3603
rect 13155 2609 13167 7131
rect 13203 2849 13215 7131
rect 13227 1961 13239 5115
rect 13251 2033 13263 7131
rect 13323 7049 13335 7131
rect 13347 5345 13359 7131
rect 13371 7073 13383 7131
rect 13275 1961 13287 5115
rect 13323 1961 13335 4299
rect 13347 1961 13359 2571
rect 13371 1961 13383 4491
rect 13419 3809 13431 7131
rect 13443 4937 13455 7131
rect 13395 1961 13407 3507
rect 13443 1961 13455 4443
rect 13467 3521 13479 7131
rect 13515 7097 13527 7131
rect 13539 5225 13551 7131
rect 13467 1961 13479 1995
rect 13491 1961 13503 4443
rect 13515 1961 13527 3123
rect 13563 2249 13575 7131
rect 13539 1961 13551 1971
rect 13587 1961 13599 3771
rect 13611 2297 13623 7131
rect 13683 7121 13695 7131
rect 13611 1961 13623 2235
rect 13635 1961 13647 3987
rect 13659 3761 13671 7035
rect 13683 1961 13695 6051
rect 13707 1961 13719 7011
rect 13731 3185 13743 7131
rect 13755 5921 13767 7131
rect 13779 2321 13791 7131
rect 13803 3737 13815 7107
rect 13827 4649 13839 7131
rect 13851 4337 13863 7131
rect 13875 5345 13887 7131
rect 13899 3929 13911 7131
rect 13947 6641 13959 7131
rect 13971 5921 13983 7131
rect 13995 5297 14007 7131
rect 13779 1961 13791 2283
rect 13899 1961 13911 3795
rect 13923 1961 13935 4155
rect 13971 1961 13983 5067
rect 14019 1961 14031 6195
rect 14043 4097 14055 7131
rect 14067 5225 14079 7131
rect 14091 4409 14103 7131
rect 14067 1961 14079 3915
rect 14115 1961 14127 6843
rect 14139 3929 14151 7131
rect 14259 6065 14271 7131
rect 14619 7049 14631 7131
rect 14667 7121 14679 7131
rect 14139 1961 14151 2715
rect 14187 1961 14199 4395
rect 14235 1961 14247 3147
rect 14259 1961 14271 4323
rect 14283 1961 14295 2811
rect 14379 1961 14391 5883
rect 14403 1961 14415 2211
rect 14475 1961 14487 5187
rect 14667 1961 14679 5427
rect 14691 1961 14703 3891
rect 14715 2657 14727 7107
rect 14739 1961 14751 5187
rect 14811 4409 14823 7131
rect 14859 5201 14871 7131
rect 14883 4073 14895 7131
rect 14907 1961 14919 6171
rect 14931 3161 14943 7131
rect 14955 1961 14967 4707
rect 15003 1961 15015 6867
rect 15027 1961 15039 2811
rect 15051 1985 15063 7131
rect 15123 1961 15135 4395
rect 15195 1961 15207 3699
rect 15219 1961 15231 3915
rect 15267 1961 15279 5931
rect 15291 1961 15303 4515
rect 15363 1961 15375 4419
rect 15411 4097 15423 7131
rect 15435 3785 15447 6435
rect 15459 5897 15471 7131
rect 15387 1961 15399 2739
rect 15411 1961 15423 3771
rect 15459 1961 15471 5187
rect 15483 1961 15495 4059
rect 15579 1961 15591 6339
rect 15603 3929 15615 7131
rect 15651 6017 15663 7131
rect 15675 6161 15687 7131
rect 15699 6449 15711 7131
rect 15723 3929 15735 7059
rect 15771 5345 15783 7131
rect 15795 5033 15807 7131
rect 15843 5105 15855 7131
rect 15675 1961 15687 3915
rect 15867 2369 15879 7131
rect 15939 5105 15951 7131
rect 15987 6929 15999 7131
rect 16011 5729 16023 7131
rect 16035 6161 16047 7131
rect 16059 3521 16071 7131
rect 16083 4817 16095 7131
rect 16131 2585 16143 7131
rect 16155 3905 16167 7131
rect 16179 4817 16191 7131
rect 16227 5729 16239 7131
rect 16251 2081 16263 7131
rect 16275 6929 16287 7131
rect 16323 4721 16335 7131
rect 16275 1961 16287 3915
rect 16347 2705 16359 7131
rect 16419 2873 16431 7131
rect 16467 7073 16479 7131
rect 16467 1961 16479 5787
rect 16539 5585 16551 7131
rect 16491 1961 16503 5139
rect 16587 4721 16599 7131
rect 16659 6785 16671 7131
rect 16683 5897 16695 7131
rect 16707 5153 16719 7131
rect 16515 1961 16527 3771
rect 16563 1961 16575 2667
rect 16683 1961 16695 4419
rect 16707 1961 16719 4899
rect 16731 1961 16743 5211
rect 16755 4481 16767 7131
rect 16755 1961 16767 3723
rect 16779 2873 16791 7131
rect 16827 5585 16839 7131
rect 16803 4457 16815 5139
rect 16875 3449 16887 7131
rect 16899 3137 16911 6051
rect 16827 1961 16839 2883
rect 16875 1961 16887 3123
rect 16923 2825 16935 7131
rect 16947 3065 16959 7131
rect 16971 5657 16983 7131
rect 16995 3977 17007 7131
rect 17019 5153 17031 7131
rect 16923 1961 16935 2715
rect 16947 1961 16959 2883
rect 17043 1961 17055 6219
rect 17067 4361 17079 7131
rect 17091 5489 17103 7131
rect 17115 4121 17127 7131
rect 17139 7097 17151 7131
rect 17211 5921 17223 7131
rect 17235 5441 17247 7131
rect 17163 1961 17175 3387
rect 17187 1961 17199 4491
rect 17211 1961 17223 4443
rect 17259 1961 17271 5379
rect 17283 2753 17295 7131
rect 17307 5729 17319 7131
rect 17307 1961 17319 3963
rect 17331 2729 17343 3411
rect 17355 2897 17367 5595
rect 17379 5489 17391 7131
rect 17379 1961 17391 3291
rect 17403 1961 17415 3051
rect 17427 2825 17439 7131
rect 17451 1961 17463 3507
rect 17475 3089 17487 5475
rect 17499 3473 17511 7131
rect 17523 3929 17535 7131
rect 17571 6785 17583 7131
rect 17523 1961 17535 3603
rect 17571 1961 17583 6291
rect 17595 5225 17607 6771
rect 17619 1961 17631 2139
rect 17643 1961 17655 6267
rect 17691 4049 17703 7131
rect 18099 7025 18111 7131
rect 17667 1961 17679 3075
rect 17763 1961 17775 2451
rect 17811 1961 17823 5835
rect 17859 1961 17871 5379
rect 17883 1961 17895 4107
rect 17955 1961 17967 6939
rect 18243 5393 18255 7131
rect 18267 5345 18279 7131
rect 18291 5873 18303 7131
rect 17979 1961 17991 2619
rect 18051 1961 18063 3987
rect 18075 1961 18087 4203
rect 18147 1961 18159 3651
rect 18171 1961 18183 4107
rect 18243 1961 18255 4083
rect 18267 1961 18279 4347
rect 18315 1961 18327 4467
rect 18339 2081 18351 7131
rect 18363 4649 18375 7131
rect 18387 2753 18399 5379
rect 18411 4505 18423 7131
rect 18459 4097 18471 7131
rect 18483 4025 18495 7131
rect 18531 5393 18543 7131
rect 18579 6689 18591 7131
rect 18603 4169 18615 7131
rect 18627 5489 18639 7131
rect 18675 4121 18687 7131
rect 18723 6521 18735 7131
rect 18771 2129 18783 7131
rect 18843 5609 18855 7131
rect 18867 2945 18879 7131
rect 18891 2057 18903 7131
rect 18963 4889 18975 7131
rect 18987 5249 18999 7131
rect 18987 1961 18999 4107
rect 19011 3377 19023 7131
rect 19035 5729 19047 7131
rect 19059 5801 19071 7131
rect 19035 1961 19047 4755
rect 19071 3281 19083 5715
rect 19107 5585 19119 7131
rect 19107 1961 19119 3651
rect 19131 3089 19143 7131
rect 19155 3401 19167 7131
rect 19179 4121 19191 6003
rect 19203 5729 19215 7131
rect 19227 5849 19239 7131
rect 19299 6329 19311 7131
rect 19323 6281 19335 7131
rect 19131 1961 19143 2931
rect 19155 1961 19167 3363
rect 19203 1961 19215 5403
rect 19227 1961 19239 4875
rect 19251 2705 19263 5835
rect 19347 5561 19359 7131
rect 19323 1961 19335 4347
rect 19347 1961 19359 3075
rect 19371 1961 19383 5955
rect 19395 4097 19407 7131
rect 19419 6113 19431 7131
rect 19443 4385 19455 7131
rect 19491 5561 19503 7131
rect 19443 1961 19455 3267
rect 19467 1961 19479 4947
rect 19515 2825 19527 7131
rect 19515 1961 19527 2787
rect 19539 1961 19551 6891
rect 19563 4313 19575 7131
rect 19563 1961 19575 4107
rect 19587 1961 19599 4371
rect 19611 2945 19623 7131
rect 19635 1961 19647 5571
rect 19659 4961 19671 7131
rect 19683 3857 19695 7131
rect 19707 6905 19719 7131
rect 19659 1961 19671 3267
rect 19707 1961 19719 6867
rect 19731 2681 19743 4947
rect 19755 3185 19767 7131
rect 19779 6929 19791 7131
rect 19803 4121 19815 7131
rect 19851 4889 19863 7131
rect 19779 1961 19791 3795
rect 19803 1961 19815 4035
rect 19851 1961 19863 4107
rect 19875 3761 19887 7131
rect 19899 4961 19911 7131
rect 19923 5849 19935 7131
rect 19899 1961 19911 2067
rect 19923 1961 19935 4995
rect 19947 2441 19959 5835
rect 19971 4097 19983 7131
rect 19971 1961 19983 3987
rect 19995 3065 20007 7131
rect 20043 6545 20055 7131
rect 20019 1961 20031 5979
rect 20055 4001 20067 4251
rect 20091 3809 20103 7131
rect 20115 4241 20127 7131
rect 20139 4169 20151 7131
rect 20163 4865 20175 7131
rect 20211 4385 20223 7131
rect 20259 6401 20271 7131
rect 20283 5489 20295 7131
rect 20139 1961 20151 3987
rect 20259 1961 20271 3099
rect 20307 2849 20319 7131
rect 20331 4121 20343 7131
rect 20355 2801 20367 5187
rect 20379 4553 20391 7131
rect 20403 5393 20415 7131
rect 20451 3569 20463 7131
rect 20475 3473 20487 4947
rect 20499 4865 20511 7131
rect 20523 6185 20535 7131
rect 20547 5729 20559 7131
rect 20595 4505 20607 7131
rect 20619 5009 20631 7131
rect 20307 1961 20319 2787
rect 20451 1961 20463 3459
rect 20523 1961 20535 2859
rect 20595 1961 20607 3219
rect 20643 1961 20655 4371
rect 20667 3281 20679 7131
rect 20715 4961 20727 7131
rect 20739 5369 20751 7131
rect 20787 5201 20799 7131
rect 20715 1961 20727 4803
rect 20763 1961 20775 5139
rect 20787 1961 20799 4947
rect 20835 4769 20847 7131
rect 20835 1961 20847 4539
rect 20859 4025 20871 7131
rect 20907 6353 20919 7131
rect 20955 4937 20967 7131
rect 20859 1961 20871 3915
rect 20883 1961 20895 2043
rect 20931 1961 20943 4107
rect 20955 1961 20967 3843
rect 20979 2273 20991 7131
rect 21003 3929 21015 5067
rect 21027 3761 21039 7131
rect 21051 1961 21063 5499
rect 21075 4457 21087 7131
rect 21099 5777 21111 7131
rect 21147 6257 21159 7131
rect 21111 3857 21123 5091
rect 21195 4265 21207 7131
rect 21075 1961 21087 2739
rect 21171 1961 21183 3819
rect 21195 1961 21207 4155
rect 21219 2753 21231 7131
rect 21243 4745 21255 7131
rect 21291 5825 21303 7131
rect 21315 5873 21327 7131
rect 21339 5921 21351 7131
rect 21363 6593 21375 7131
rect 21411 6617 21423 7131
rect 21243 1961 21255 4203
rect 21291 1961 21303 2163
rect 21315 1961 21327 4443
rect 21339 1961 21351 3915
rect 21363 1961 21375 3843
rect 21411 1961 21423 5283
rect 21435 3977 21447 7131
rect 21459 4793 21471 7131
rect 21483 4121 21495 7131
rect 21531 5873 21543 7131
rect 21555 5753 21567 7131
rect 21603 6665 21615 7131
rect 21459 1961 21471 2091
rect 21531 1961 21543 3315
rect 21555 1961 21567 3795
rect 21579 1961 21591 6267
rect 21651 4241 21663 7131
rect 21675 4961 21687 7131
rect 21699 6713 21711 7131
rect 21603 1961 21615 2811
rect 21675 1961 21687 4923
rect 21699 1961 21711 4011
rect 21723 3329 21735 4947
rect 21747 2249 21759 7131
rect 21795 3209 21807 7131
rect 21819 3185 21831 5259
rect 21795 1961 21807 3171
rect 21867 1961 21879 5331
rect 21915 1961 21927 5427
rect 21939 3857 21951 7131
rect 22347 5993 22359 7131
rect 21987 1961 21999 1995
rect 22011 1961 22023 3939
rect 22035 1961 22047 5259
rect 22059 1961 22071 4107
rect 22131 1961 22143 5283
rect 22155 1961 22167 5187
rect 22179 1961 22191 3699
rect 22251 1961 22263 3603
rect 22275 1961 22287 5883
rect 22299 1961 22311 5067
rect 22323 1961 22335 4923
rect 22347 1961 22359 3699
rect 22395 1961 22407 4155
rect 22419 1961 22431 6267
rect 22491 3593 22503 7131
rect 22443 1961 22455 3267
rect 22515 3089 22527 7131
rect 22563 5705 22575 7131
rect 22611 4961 22623 7131
rect 22515 1961 22527 2019
rect 22539 1961 22551 4155
rect 22611 1961 22623 4875
rect 22635 4745 22647 7131
rect 22635 1961 22647 3795
rect 22659 1961 22671 6003
rect 22683 2513 22695 7131
rect 22731 6977 22743 7131
rect 22755 6425 22767 7131
rect 22779 5465 22791 7131
rect 22803 6041 22815 7131
rect 22707 1961 22719 4011
rect 22755 1961 22767 5163
rect 22827 4865 22839 7131
rect 22803 1961 22815 3963
rect 22851 1961 22863 4899
rect 22875 2993 22887 7131
rect 22899 4217 22911 7131
rect 22923 5537 22935 7131
rect 22971 5057 22983 7131
rect 22935 3569 22947 4947
rect 22875 1961 22887 2067
rect 22971 1961 22983 5019
rect 22995 4649 23007 7131
rect 23019 4625 23031 7131
rect 22995 1961 23007 4347
rect 23067 3233 23079 7131
rect 23091 6185 23103 7131
rect 23043 1961 23055 2571
rect 23091 1961 23103 6123
rect 23115 4625 23127 7131
rect 23115 1961 23127 4419
rect 23139 1961 23151 6795
rect 23163 5945 23175 7131
rect 23211 6377 23223 7131
rect 23175 2777 23187 4731
rect 23211 1961 23223 4707
rect 23283 4361 23295 7131
rect 23307 3977 23319 6819
rect 23235 1961 23247 2547
rect 23259 1961 23271 2403
rect 23283 1961 23295 3843
rect 23331 2753 23343 7131
rect 23367 4025 23379 6171
rect 23403 3785 23415 7131
rect 23427 3497 23439 7131
rect 23475 6185 23487 7131
rect 23331 1961 23343 2715
rect 23355 1961 23367 2739
rect 23451 1961 23463 4875
rect 23475 1961 23487 6147
rect 23523 5681 23535 7131
rect 23547 4625 23559 7131
rect 23499 3929 23511 4611
rect 23523 1961 23535 2691
rect 23571 1961 23583 5091
rect 23595 2393 23607 7131
rect 23619 2729 23631 6435
rect 23643 5417 23655 7131
rect 23667 1961 23679 3675
rect 23691 2993 23703 7131
rect 23763 4121 23775 7131
rect 23787 4889 23799 7131
rect 23811 4649 23823 7131
rect 23787 1961 23799 4323
rect 23811 1961 23823 4251
rect 23835 1961 23847 4611
rect 23859 3257 23871 7131
rect 23883 5585 23895 7131
rect 23883 1961 23895 5067
rect 23907 3041 23919 7131
rect 23931 1961 23943 5211
rect 23955 4193 23967 7131
rect 23979 2609 23991 7131
rect 24027 4409 24039 7131
rect 24027 1961 24039 3147
rect 24075 2873 24087 7131
rect 24099 3257 24111 7131
rect 24123 4361 24135 7131
rect 24147 4625 24159 7131
rect 24195 5009 24207 7131
rect 24171 1961 24183 4563
rect 24243 2273 24255 7131
rect 24291 1961 24303 5547
rect 24315 3521 24327 7131
rect 24339 4361 24351 7131
rect 24339 1961 24351 4323
rect 24363 2417 24375 7131
rect 24411 6233 24423 7131
rect 24435 5873 24447 7131
rect 24483 6641 24495 7131
rect 24363 1961 24375 2379
rect 24387 1961 24399 4395
rect 24435 1961 24447 4515
rect 24495 4337 24507 6363
rect 24459 1961 24471 4131
rect 24531 3665 24543 7131
rect 24579 4457 24591 7131
rect 24531 1961 24543 3603
rect 24555 1961 24567 4347
rect 24603 2393 24615 6339
rect 24627 3545 24639 7131
rect 24651 3809 24663 7131
rect 24675 2297 24687 7131
rect 24699 3617 24711 6843
rect 24723 2345 24735 7131
rect 24771 4697 24783 7131
rect 24843 6137 24855 7131
rect 24891 4601 24903 7131
rect 24963 4673 24975 7131
rect 24987 6569 24999 7131
rect 25035 4001 25047 7131
rect 25083 6089 25095 7131
rect 24723 1961 24735 2187
rect 25083 1961 25095 4923
rect 25107 3377 25119 7131
rect 25131 4577 25143 7131
rect 25131 1961 25143 4419
rect 25155 2969 25167 7131
rect 25203 4769 25215 7131
rect 25179 4385 25191 4563
rect 25227 3065 25239 7131
rect 25275 4577 25287 7131
rect 25323 5249 25335 7131
rect 25275 1961 25287 3651
rect 25299 2153 25311 4563
rect 25323 1961 25335 4515
rect 25347 4097 25359 7131
rect 25371 4529 25383 5595
rect 25395 4241 25407 7131
rect 25419 4193 25431 5619
rect 25395 1961 25407 4179
rect 25443 4097 25455 7131
rect 25467 4937 25479 7131
rect 25515 5177 25527 7131
rect 25443 1961 25455 4011
rect 25515 1961 25527 2907
rect 25539 1961 25551 7035
rect 25563 6977 25575 7131
rect 25563 1961 25575 6939
rect 25587 2297 25599 7131
rect 25611 4649 25623 7131
rect 25635 6017 25647 7131
rect 25659 4577 25671 7131
rect 25707 6905 25719 7131
rect 25731 5897 25743 7131
rect 25683 1961 25695 4563
rect 25755 2009 25767 7131
rect 25779 3737 25791 6963
rect 25803 2489 25815 7131
rect 25827 3809 25839 7131
rect 25851 6473 25863 7131
rect 25899 5129 25911 7131
rect 25923 4841 25935 7131
rect 25947 6185 25959 7131
rect 25971 5273 25983 7131
rect 25995 4577 26007 7131
rect 26043 6689 26055 7131
rect 26067 4217 26079 7131
rect 26043 1961 26055 4155
rect 26091 1961 26103 4875
rect 26163 4097 26175 7131
rect 26187 4265 26199 7131
rect 26211 2249 26223 7131
rect 26259 3905 26271 7131
rect 26307 5921 26319 7131
rect 26379 7073 26391 7131
rect 26235 1961 26247 3627
rect 26259 1961 26271 3699
rect 26307 1961 26319 2547
rect 26355 1961 26367 5067
rect 26379 1961 26391 5259
rect 26403 4361 26415 7131
rect 26427 7001 26439 7131
rect 26403 1961 26415 4323
rect 26427 1961 26439 5883
rect 26451 4337 26463 4971
rect 26475 3521 26487 7131
rect 26499 4481 26511 7131
rect 26499 1961 26511 4443
rect 26523 3017 26535 7131
rect 26571 6521 26583 7131
rect 26595 5225 26607 7131
rect 26619 3953 26631 7131
rect 26643 4457 26655 4491
rect 26667 4073 26679 7131
rect 26523 1961 26535 2259
rect 26547 1961 26559 3339
rect 26667 1961 26679 3867
rect 26691 3113 26703 7131
rect 26739 2873 26751 7131
rect 26739 1961 26751 2835
rect 26763 1961 26775 4995
rect 26787 4601 26799 7131
rect 26811 4553 26823 7131
rect 26811 1961 26823 4515
rect 26835 4289 26847 7131
rect 26859 1961 26871 4611
rect 26883 2585 26895 7131
rect 26907 4313 26919 7131
rect 26931 5321 26943 7131
rect 26955 2849 26967 5907
rect 26979 4409 26991 7131
rect 27003 5801 27015 7131
rect 27027 4049 27039 7131
rect 27099 5657 27111 7131
rect 27051 4529 27063 5499
rect 27123 4697 27135 7131
rect 27147 6737 27159 7131
rect 27195 6209 27207 7131
rect 27315 4433 27327 7131
rect 27339 2081 27351 7131
rect 27363 6497 27375 7131
rect 27411 4025 27423 7131
rect 27411 1985 27423 2523
rect 27435 2009 27447 6747
rect 27555 1961 27755 7131
rect 27867 4564 27937 4576
rect 27867 3844 27937 3856
rect 27867 1996 27937 2008
rect 27867 1972 27937 1984
rect 0 107 70 119
rect 0 83 70 95
rect 123 0 323 1162
rect 339 0 351 1162
rect 363 0 375 1162
rect 387 0 399 1162
rect 411 0 423 1162
rect 1683 144 1695 1162
rect 1803 168 1815 1162
rect 2355 96 2367 1162
rect 2403 96 2415 1162
rect 2475 192 2487 1162
rect 2523 216 2535 1162
rect 2619 72 2631 1162
rect 2739 240 2751 1162
rect 2859 264 2871 1162
rect 3531 288 3543 1162
rect 3651 312 3663 1162
rect 3675 336 3687 1162
rect 4131 48 4143 1162
rect 4155 360 4167 1162
rect 4203 384 4215 1162
rect 4299 336 4311 1162
rect 4467 408 4479 1162
rect 4587 432 4599 1162
rect 4875 456 4887 1162
rect 4923 480 4935 1162
rect 4947 504 4959 1162
rect 5475 528 5487 1162
rect 5835 552 5847 1162
rect 5931 576 5943 1162
rect 5979 600 5991 1162
rect 6027 504 6039 1162
rect 6075 504 6087 1162
rect 6099 624 6111 1162
rect 6243 648 6255 1162
rect 6411 672 6423 1162
rect 6747 528 6759 1162
rect 6939 528 6951 1162
rect 6963 696 6975 1162
rect 7227 720 7239 1162
rect 7323 744 7335 1162
rect 7419 504 7431 1162
rect 7467 504 7479 1162
rect 7611 168 7623 1162
rect 7683 576 7695 1162
rect 8283 576 8295 1162
rect 8031 0 8043 154
rect 8379 48 8391 1162
rect 8427 192 8439 1162
rect 8547 192 8559 1162
rect 8715 600 8727 1162
rect 8787 768 8799 1162
rect 9123 792 9135 1162
rect 9507 816 9519 1162
rect 9819 576 9831 1162
rect 9867 576 9879 1162
rect 9939 840 9951 1162
rect 9987 864 9999 1162
rect 10011 888 10023 1162
rect 10035 360 10047 1162
rect 10275 336 10287 1162
rect 10635 360 10647 1162
rect 10683 360 10695 1162
rect 10707 912 10719 1162
rect 10755 360 10767 1162
rect 10851 936 10863 1162
rect 10923 960 10935 1162
rect 11019 144 11031 1162
rect 11043 984 11055 1162
rect 11091 144 11103 1162
rect 11187 624 11199 1162
rect 11235 624 11247 1162
rect 8067 0 8079 34
rect 11955 24 11967 1162
rect 12315 1008 12327 1162
rect 12339 648 12351 1162
rect 12387 648 12399 1162
rect 12675 1032 12687 1162
rect 13155 1056 13167 1162
rect 13203 1080 13215 1162
rect 13731 864 13743 1162
rect 13803 720 13815 1162
rect 13851 960 13863 1162
rect 14043 720 14055 1162
rect 14307 384 14319 1162
rect 14355 864 14367 1162
rect 14451 960 14463 1162
rect 14523 384 14535 1162
rect 14571 1104 14583 1162
rect 14595 1056 14607 1162
rect 14619 264 14631 1162
rect 14787 1056 14799 1162
rect 14835 264 14847 1162
rect 14931 768 14943 1162
rect 15075 576 15087 1162
rect 15147 576 15159 1162
rect 15171 360 15183 1162
rect 15315 360 15327 1162
rect 15507 600 15519 1162
rect 15555 360 15567 1162
rect 15627 360 15639 1162
rect 15699 744 15711 1162
rect 15747 744 15759 1162
rect 15867 1128 15879 1162
rect 16419 1152 16431 1162
rect 16443 744 16455 1162
rect 16611 864 16623 1162
rect 16803 192 16815 1162
rect 16851 696 16863 1162
rect 16995 288 17007 1162
rect 17067 384 17079 1162
rect 17115 984 17127 1162
rect 17499 648 17511 1162
rect 17691 720 17703 1162
rect 17739 648 17751 1162
rect 17907 696 17919 1162
rect 18003 720 18015 1162
rect 18099 1008 18111 1162
rect 18195 888 18207 1162
rect 18435 96 18447 1162
rect 18843 1128 18855 1162
rect 19275 912 19287 1162
rect 19419 768 19431 1162
rect 19755 552 19767 1162
rect 19851 120 19863 1162
rect 20043 600 20055 1162
rect 20091 504 20103 1162
rect 20163 744 20175 1162
rect 20211 768 20223 1162
rect 20379 408 20391 1162
rect 20403 600 20415 1162
rect 20427 432 20439 1162
rect 20499 720 20511 1162
rect 20547 480 20559 1162
rect 20619 720 20631 1162
rect 20691 768 20703 1162
rect 20632 706 20650 720
rect 20631 0 20643 706
rect 20739 144 20751 1162
rect 20979 0 20991 514
rect 21003 312 21015 1162
rect 21123 960 21135 1162
rect 21627 816 21639 1162
rect 22107 336 22119 1162
rect 22203 720 22215 1162
rect 22467 768 22479 1162
rect 22563 816 22575 1162
rect 22707 168 22719 1162
rect 22779 792 22791 1162
rect 22923 1080 22935 1162
rect 23187 576 23199 1162
rect 23379 1152 23391 1162
rect 23427 1056 23439 1162
rect 23643 816 23655 1162
rect 23691 696 23703 1162
rect 23715 456 23727 1162
rect 23739 1032 23751 1162
rect 23907 936 23919 1162
rect 23955 1104 23967 1162
rect 24003 672 24015 1162
rect 24075 48 24087 1162
rect 24123 840 24135 1162
rect 24243 600 24255 1162
rect 24267 408 24279 1162
rect 24483 1056 24495 1162
rect 24603 744 24615 1162
rect 26451 624 26463 1162
rect 26595 264 26607 1162
rect 26619 216 26631 1162
rect 26643 240 26655 1162
rect 26691 648 26703 1162
rect 26883 768 26895 1162
rect 26931 576 26943 1162
rect 26931 24 26943 34
rect 26955 24 26967 346
rect 27555 0 27755 1162
rect 27867 707 27937 719
rect 27867 59 27937 71
rect 27867 35 27937 47
rect 27867 11 27937 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7131
box 0 0 1464 799
use nand2 g8291
timestamp 1386234792
transform 1 0 1587 0 1 7131
box 0 0 96 799
use nand3 g8060
timestamp 1386234893
transform 1 0 1683 0 1 7131
box 0 0 120 799
use nor2 g8182
timestamp 1386235306
transform 1 0 1803 0 1 7131
box 0 0 120 799
use nand3 g8066
timestamp 1386234893
transform 1 0 1923 0 1 7131
box 0 0 120 799
use nor2 g8169
timestamp 1386235306
transform 1 0 2043 0 1 7131
box 0 0 120 799
use nand2 g8107
timestamp 1386234792
transform 1 0 2163 0 1 7131
box 0 0 96 799
use nand2 g8229
timestamp 1386234792
transform 1 0 2259 0 1 7131
box 0 0 96 799
use nand2 g8313
timestamp 1386234792
transform 1 0 2355 0 1 7131
box 0 0 96 799
use inv g8039
timestamp 1386238110
transform 1 0 2451 0 1 7131
box 0 0 120 799
use nand2 g8344
timestamp 1386234792
transform 1 0 2571 0 1 7131
box 0 0 96 799
use inv g8123
timestamp 1386238110
transform 1 0 2667 0 1 7131
box 0 0 120 799
use nand2 g8046
timestamp 1386234792
transform 1 0 2787 0 1 7131
box 0 0 96 799
use nand2 g8222
timestamp 1386234792
transform 1 0 2883 0 1 7131
box 0 0 96 799
use nand2 g8098
timestamp 1386234792
transform 1 0 2979 0 1 7131
box 0 0 96 799
use inv g8102
timestamp 1386238110
transform 1 0 3075 0 1 7131
box 0 0 120 799
use nand4 g8327
timestamp 1386234936
transform 1 0 3195 0 1 7131
box 0 0 144 799
use and2 g8314
timestamp 1386234845
transform 1 0 3339 0 1 7131
box 0 0 120 799
use nand2 g8012
timestamp 1386234792
transform 1 0 3459 0 1 7131
box 0 0 96 799
use nand2 g8187
timestamp 1386234792
transform 1 0 3555 0 1 7131
box 0 0 96 799
use nand2 g8135
timestamp 1386234792
transform 1 0 3651 0 1 7131
box 0 0 96 799
use nand2 g8171
timestamp 1386234792
transform 1 0 3747 0 1 7131
box 0 0 96 799
use and2 g8295
timestamp 1386234845
transform 1 0 3843 0 1 7131
box 0 0 120 799
use mux2 g8287
timestamp 1386235218
transform 1 0 3963 0 1 7131
box 0 0 192 799
use nor2 g8154
timestamp 1386235306
transform 1 0 4155 0 1 7131
box 0 0 120 799
use nand2 g8276
timestamp 1386234792
transform 1 0 4275 0 1 7131
box 0 0 96 799
use nand2 g8261
timestamp 1386234792
transform 1 0 4371 0 1 7131
box 0 0 96 799
use and2 g8130
timestamp 1386234845
transform 1 0 4467 0 1 7131
box 0 0 120 799
use nand2 g8027
timestamp 1386234792
transform 1 0 4587 0 1 7131
box 0 0 96 799
use nor2 g8082
timestamp 1386235306
transform 1 0 4683 0 1 7131
box 0 0 120 799
use nand2 g8318
timestamp 1386234792
transform 1 0 4803 0 1 7131
box 0 0 96 799
use nor2 g8035
timestamp 1386235306
transform 1 0 4899 0 1 7131
box 0 0 120 799
use and2 g8019
timestamp 1386234845
transform 1 0 5019 0 1 7131
box 0 0 120 799
use nand3 g8168
timestamp 1386234893
transform 1 0 5139 0 1 7131
box 0 0 120 799
use inv g8238
timestamp 1386238110
transform 1 0 5259 0 1 7131
box 0 0 120 799
use nand2 g7989
timestamp 1386234792
transform 1 0 5379 0 1 7131
box 0 0 96 799
use nand2 g8225
timestamp 1386234792
transform 1 0 5475 0 1 7131
box 0 0 96 799
use nand2 g8143
timestamp 1386234792
transform 1 0 5571 0 1 7131
box 0 0 96 799
use nand3 g8333
timestamp 1386234893
transform 1 0 5667 0 1 7131
box 0 0 120 799
use inv g2
timestamp 1386238110
transform 1 0 5787 0 1 7131
box 0 0 120 799
use nand4 g8042
timestamp 1386234936
transform 1 0 5907 0 1 7131
box 0 0 144 799
use nand2 g8069
timestamp 1386234792
transform 1 0 6051 0 1 7131
box 0 0 96 799
use nand2 g8149
timestamp 1386234792
transform 1 0 6147 0 1 7131
box 0 0 96 799
use nand4 g8338
timestamp 1386234936
transform 1 0 6243 0 1 7131
box 0 0 144 799
use inv g8280
timestamp 1386238110
transform 1 0 6387 0 1 7131
box 0 0 120 799
use nand3 g7985
timestamp 1386234893
transform 1 0 6507 0 1 7131
box 0 0 120 799
use nand2 g8249
timestamp 1386234792
transform 1 0 6627 0 1 7131
box 0 0 96 799
use nor2 g8064
timestamp 1386235306
transform 1 0 6723 0 1 7131
box 0 0 120 799
use nand2 g8310
timestamp 1386234792
transform 1 0 6843 0 1 7131
box 0 0 96 799
use nor2 g8235
timestamp 1386235306
transform 1 0 6939 0 1 7131
box 0 0 120 799
use and2 g8058
timestamp 1386234845
transform 1 0 7059 0 1 7131
box 0 0 120 799
use nand2 g8009
timestamp 1386234792
transform 1 0 7179 0 1 7131
box 0 0 96 799
use nor2 g8055
timestamp 1386235306
transform 1 0 7275 0 1 7131
box 0 0 120 799
use nand2 g8088
timestamp 1386234792
transform 1 0 7395 0 1 7131
box 0 0 96 799
use and2 g8214
timestamp 1386234845
transform 1 0 7491 0 1 7131
box 0 0 120 799
use nand2 g8056
timestamp 1386234792
transform 1 0 7611 0 1 7131
box 0 0 96 799
use nand3 g8281
timestamp 1386234893
transform 1 0 7707 0 1 7131
box 0 0 120 799
use and2 g8269
timestamp 1386234845
transform 1 0 7827 0 1 7131
box 0 0 120 799
use nand2 g8183
timestamp 1386234792
transform 1 0 7947 0 1 7131
box 0 0 96 799
use nand3 g8170
timestamp 1386234893
transform 1 0 8043 0 1 7131
box 0 0 120 799
use nand2 g8124
timestamp 1386234792
transform 1 0 8163 0 1 7131
box 0 0 96 799
use nand2 g8106
timestamp 1386234792
transform 1 0 8259 0 1 7131
box 0 0 96 799
use nand2 g8119
timestamp 1386234792
transform 1 0 8355 0 1 7131
box 0 0 96 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 8451 0 1 7131
box 0 0 48 799
use nand2 g8275
timestamp 1386234792
transform 1 0 8499 0 1 7131
box 0 0 96 799
use nand2 g8146
timestamp 1386234792
transform 1 0 8595 0 1 7131
box 0 0 96 799
use nand3 g8127
timestamp 1386234893
transform 1 0 8691 0 1 7131
box 0 0 120 799
use nand2 g8155
timestamp 1386234792
transform 1 0 8811 0 1 7131
box 0 0 96 799
use nand2 g8290
timestamp 1386234792
transform 1 0 8907 0 1 7131
box 0 0 96 799
use nand2 g8033
timestamp 1386234792
transform 1 0 9003 0 1 7131
box 0 0 96 799
use nand2 g8252
timestamp 1386234792
transform 1 0 9099 0 1 7131
box 0 0 96 799
use nand2 g7978
timestamp 1386234792
transform 1 0 9195 0 1 7131
box 0 0 96 799
use nand4 g8334
timestamp 1386234936
transform 1 0 9291 0 1 7131
box 0 0 144 799
use nand2 g8244
timestamp 1386234792
transform 1 0 9435 0 1 7131
box 0 0 96 799
use nand3 g7972
timestamp 1386234893
transform 1 0 9531 0 1 7131
box 0 0 120 799
use nand4 g8240
timestamp 1386234936
transform 1 0 9651 0 1 7131
box 0 0 144 799
use rowcrosser PcWe
timestamp 1386086759
transform 1 0 9795 0 1 7131
box 0 0 48 799
use and2 g8054
timestamp 1386234845
transform 1 0 9843 0 1 7131
box 0 0 120 799
use nand2 g8139
timestamp 1386234792
transform 1 0 9963 0 1 7131
box 0 0 96 799
use nand2 g8118
timestamp 1386234792
transform 1 0 10059 0 1 7131
box 0 0 96 799
use inv g8023
timestamp 1386238110
transform 1 0 10155 0 1 7131
box 0 0 120 799
use nand4 g7981
timestamp 1386234936
transform 1 0 10275 0 1 7131
box 0 0 144 799
use nand2 g8111
timestamp 1386234792
transform 1 0 10419 0 1 7131
box 0 0 96 799
use nand2 g8120
timestamp 1386234792
transform 1 0 10515 0 1 7131
box 0 0 96 799
use nand2 g8091
timestamp 1386234792
transform 1 0 10611 0 1 7131
box 0 0 96 799
use nand2 g8134
timestamp 1386234792
transform 1 0 10707 0 1 7131
box 0 0 96 799
use nor2 g8320
timestamp 1386235306
transform 1 0 10803 0 1 7131
box 0 0 120 799
use nor2 g8050
timestamp 1386235306
transform 1 0 10923 0 1 7131
box 0 0 120 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 11043 0 1 7131
box 0 0 48 799
use nand2 g8218
timestamp 1386234792
transform 1 0 11091 0 1 7131
box 0 0 96 799
use nand2 g7995
timestamp 1386234792
transform 1 0 11187 0 1 7131
box 0 0 96 799
use nand3 g8284
timestamp 1386234893
transform 1 0 11283 0 1 7131
box 0 0 120 799
use and2 g7964
timestamp 1386234845
transform 1 0 11403 0 1 7131
box 0 0 120 799
use nand4 g8198
timestamp 1386234936
transform 1 0 11523 0 1 7131
box 0 0 144 799
use nor2 g8272
timestamp 1386235306
transform 1 0 11667 0 1 7131
box 0 0 120 799
use nand2 g8199
timestamp 1386234792
transform 1 0 11787 0 1 7131
box 0 0 96 799
use nand2 g8306
timestamp 1386234792
transform 1 0 11883 0 1 7131
box 0 0 96 799
use nand2 g8221
timestamp 1386234792
transform 1 0 11979 0 1 7131
box 0 0 96 799
use nand2 g8319
timestamp 1386234792
transform 1 0 12075 0 1 7131
box 0 0 96 799
use nor2 g8220
timestamp 1386235306
transform 1 0 12171 0 1 7131
box 0 0 120 799
use inv g8194
timestamp 1386238110
transform 1 0 12291 0 1 7131
box 0 0 120 799
use nor2 g8230
timestamp 1386235306
transform 1 0 12411 0 1 7131
box 0 0 120 799
use nand3 g8271
timestamp 1386234893
transform 1 0 12531 0 1 7131
box 0 0 120 799
use nand2 g8004
timestamp 1386234792
transform 1 0 12651 0 1 7131
box 0 0 96 799
use nand2 rm_assigns_buf_StatusReg_1
timestamp 1386234792
transform 1 0 12747 0 1 7131
box 0 0 96 799
use buffer g8209
timestamp 1386236986
transform 1 0 12843 0 1 7131
box 0 0 120 799
use nand2 g8103
timestamp 1386234792
transform 1 0 12963 0 1 7131
box 0 0 96 799
use nor2 g8268
timestamp 1386235306
transform 1 0 13059 0 1 7131
box 0 0 120 799
use inv g8283
timestamp 1386238110
transform 1 0 13179 0 1 7131
box 0 0 120 799
use nand2 g8321
timestamp 1386234792
transform 1 0 13299 0 1 7131
box 0 0 96 799
use nand2 g8180
timestamp 1386234792
transform 1 0 13395 0 1 7131
box 0 0 96 799
use nand2 g8005
timestamp 1386234792
transform 1 0 13491 0 1 7131
box 0 0 96 799
use nor2 g8052
timestamp 1386235306
transform 1 0 13587 0 1 7131
box 0 0 120 799
use nand2 g8136
timestamp 1386234792
transform 1 0 13707 0 1 7131
box 0 0 96 799
use nand3 g8110
timestamp 1386234893
transform 1 0 13803 0 1 7131
box 0 0 120 799
use nand2 g8153
timestamp 1386234792
transform 1 0 13923 0 1 7131
box 0 0 96 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 14019 0 1 7131
box 0 0 96 799
use rowcrosser AluWe
timestamp 1386086759
transform 1 0 14115 0 1 7131
box 0 0 48 799
use scandtype g8308
timestamp 1386241841
transform 1 0 14163 0 1 7131
box 0 0 624 799
use rowcrosser LrWe
timestamp 1386086759
transform 1 0 14787 0 1 7131
box 0 0 48 799
use nor2 stateSub_reg_91_2_93_
timestamp 1386235306
transform 1 0 14835 0 1 7131
box 0 0 120 799
use scandtype g8294
timestamp 1386241841
transform 1 0 14955 0 1 7131
box 0 0 624 799
use rowcrosser g8048
timestamp 1386086759
transform 1 0 15579 0 1 7131
box 0 0 48 799
use nand2 g8024
timestamp 1386234792
transform 1 0 15627 0 1 7131
box 0 0 96 799
use mux2 g8099
timestamp 1386235218
transform 1 0 15723 0 1 7131
box 0 0 192 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 15915 0 1 7131
box 0 0 48 799
use nand4 g8057
timestamp 1386234936
transform 1 0 15963 0 1 7131
box 0 0 144 799
use nand2 g8190
timestamp 1386234792
transform 1 0 16107 0 1 7131
box 0 0 96 799
use nand2 g8045
timestamp 1386234792
transform 1 0 16203 0 1 7131
box 0 0 96 799
use nand2 g8304
timestamp 1386234792
transform 1 0 16299 0 1 7131
box 0 0 96 799
use inv g8018
timestamp 1386238110
transform 1 0 16395 0 1 7131
box 0 0 120 799
use inv g8092
timestamp 1386238110
transform 1 0 16515 0 1 7131
box 0 0 120 799
use nand2 g8277
timestamp 1386234792
transform 1 0 16635 0 1 7131
box 0 0 96 799
use and2 g8081
timestamp 1386234845
transform 1 0 16731 0 1 7131
box 0 0 120 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 16851 0 1 7131
box 0 0 48 799
use nand4 g8243
timestamp 1386234936
transform 1 0 16899 0 1 7131
box 0 0 144 799
use nand3 g8296
timestamp 1386234893
transform 1 0 17043 0 1 7131
box 0 0 120 799
use mux2 g8348
timestamp 1386235218
transform 1 0 17163 0 1 7131
box 0 0 192 799
use inv g8234
timestamp 1386238110
transform 1 0 17355 0 1 7131
box 0 0 120 799
use and2 StatusReg_reg_91_1_93_
timestamp 1386234845
transform 1 0 17475 0 1 7131
box 0 0 120 799
use scandtype g8324
timestamp 1386241841
transform 1 0 17595 0 1 7131
box 0 0 624 799
use nand2 g8293
timestamp 1386234792
transform 1 0 18219 0 1 7131
box 0 0 96 799
use nor2 g8312
timestamp 1386235306
transform 1 0 18315 0 1 7131
box 0 0 120 799
use and2 g8028
timestamp 1386234845
transform 1 0 18435 0 1 7131
box 0 0 120 799
use nand2 g8213
timestamp 1386234792
transform 1 0 18555 0 1 7131
box 0 0 96 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 18651 0 1 7131
box 0 0 48 799
use inv g7963
timestamp 1386238110
transform 1 0 18699 0 1 7131
box 0 0 120 799
use nand3 g8096
timestamp 1386234893
transform 1 0 18819 0 1 7131
box 0 0 120 799
use nand4 g8212
timestamp 1386234936
transform 1 0 18939 0 1 7131
box 0 0 144 799
use nand2 g8015
timestamp 1386234792
transform 1 0 19083 0 1 7131
box 0 0 96 799
use nand2 g8084
timestamp 1386234792
transform 1 0 19179 0 1 7131
box 0 0 96 799
use nand2 g8265
timestamp 1386234792
transform 1 0 19275 0 1 7131
box 0 0 96 799
use nand2 g8200
timestamp 1386234792
transform 1 0 19371 0 1 7131
box 0 0 96 799
use and2 g8108
timestamp 1386234845
transform 1 0 19467 0 1 7131
box 0 0 120 799
use rowcrosser StatusRegEn
timestamp 1386086759
transform 1 0 19587 0 1 7131
box 0 0 48 799
use nand2 g8049
timestamp 1386234792
transform 1 0 19635 0 1 7131
box 0 0 96 799
use nand2 g8144
timestamp 1386234792
transform 1 0 19731 0 1 7131
box 0 0 96 799
use nand3 g8159
timestamp 1386234893
transform 1 0 19827 0 1 7131
box 0 0 120 799
use and2 g8177
timestamp 1386234845
transform 1 0 19947 0 1 7131
box 0 0 120 799
use nand3 g7996
timestamp 1386234893
transform 1 0 20067 0 1 7131
box 0 0 120 799
use rowcrosser PcSel_91_2_93_
timestamp 1386086759
transform 1 0 20187 0 1 7131
box 0 0 48 799
use nand3 g8251
timestamp 1386234893
transform 1 0 20235 0 1 7131
box 0 0 120 799
use nor2 g8036
timestamp 1386235306
transform 1 0 20355 0 1 7131
box 0 0 120 799
use nand2 g8226
timestamp 1386234792
transform 1 0 20475 0 1 7131
box 0 0 96 799
use and2 g7979
timestamp 1386234845
transform 1 0 20571 0 1 7131
box 0 0 120 799
use nor2 g8264
timestamp 1386235306
transform 1 0 20691 0 1 7131
box 0 0 120 799
use and2 g8332
timestamp 1386234845
transform 1 0 20811 0 1 7131
box 0 0 120 799
use nor2 g8089
timestamp 1386235306
transform 1 0 20931 0 1 7131
box 0 0 120 799
use and2 g8206
timestamp 1386234845
transform 1 0 21051 0 1 7131
box 0 0 120 799
use nand2 g8237
timestamp 1386234792
transform 1 0 21171 0 1 7131
box 0 0 96 799
use nand3 g8016
timestamp 1386234893
transform 1 0 21267 0 1 7131
box 0 0 120 799
use nand3 g8278
timestamp 1386234893
transform 1 0 21387 0 1 7131
box 0 0 120 799
use nor2 g8181
timestamp 1386235306
transform 1 0 21507 0 1 7131
box 0 0 120 799
use nand2 g8216
timestamp 1386234792
transform 1 0 21627 0 1 7131
box 0 0 96 799
use inv StatusReg_reg_91_0_93_
timestamp 1386238110
transform 1 0 21723 0 1 7131
box 0 0 120 799
use scandtype g8253
timestamp 1386241841
transform 1 0 21843 0 1 7131
box 0 0 624 799
use nor2 g8186
timestamp 1386235306
transform 1 0 22467 0 1 7131
box 0 0 120 799
use nor2 g8090
timestamp 1386235306
transform 1 0 22587 0 1 7131
box 0 0 120 799
use nand4 g8223
timestamp 1386234936
transform 1 0 22707 0 1 7131
box 0 0 144 799
use nand2 g8195
timestamp 1386234792
transform 1 0 22851 0 1 7131
box 0 0 96 799
use nand2 g8077
timestamp 1386234792
transform 1 0 22947 0 1 7131
box 0 0 96 799
use nand2 g8133
timestamp 1386234792
transform 1 0 23043 0 1 7131
box 0 0 96 799
use inv g8341
timestamp 1386238110
transform 1 0 23139 0 1 7131
box 0 0 120 799
use inv g7971
timestamp 1386238110
transform 1 0 23259 0 1 7131
box 0 0 120 799
use nor2 g8041
timestamp 1386235306
transform 1 0 23379 0 1 7131
box 0 0 120 799
use and2 g8289
timestamp 1386234845
transform 1 0 23499 0 1 7131
box 0 0 120 799
use inv g8002
timestamp 1386238110
transform 1 0 23619 0 1 7131
box 0 0 120 799
use nand2 g8128
timestamp 1386234792
transform 1 0 23739 0 1 7131
box 0 0 96 799
use nand2 g8029
timestamp 1386234792
transform 1 0 23835 0 1 7131
box 0 0 96 799
use nor2 g8100
timestamp 1386235306
transform 1 0 23931 0 1 7131
box 0 0 120 799
use nand3 g8350
timestamp 1386234893
transform 1 0 24051 0 1 7131
box 0 0 120 799
use inv g8117
timestamp 1386238110
transform 1 0 24171 0 1 7131
box 0 0 120 799
use nand2 g8167
timestamp 1386234792
transform 1 0 24291 0 1 7131
box 0 0 96 799
use nor2 g7982
timestamp 1386235306
transform 1 0 24387 0 1 7131
box 0 0 120 799
use nand2 g8191
timestamp 1386234792
transform 1 0 24507 0 1 7131
box 0 0 96 799
use nand2 g8227
timestamp 1386234792
transform 1 0 24603 0 1 7131
box 0 0 96 799
use inv g8270
timestamp 1386238110
transform 1 0 24699 0 1 7131
box 0 0 120 799
use inv g8073
timestamp 1386238110
transform 1 0 24819 0 1 7131
box 0 0 120 799
use and2 g7967
timestamp 1386234845
transform 1 0 24939 0 1 7131
box 0 0 120 799
use nand3 g8163
timestamp 1386234893
transform 1 0 25059 0 1 7131
box 0 0 120 799
use and2 g8273
timestamp 1386234845
transform 1 0 25179 0 1 7131
box 0 0 120 799
use and2 g8337
timestamp 1386234845
transform 1 0 25299 0 1 7131
box 0 0 120 799
use nor2 g7969
timestamp 1386235306
transform 1 0 25419 0 1 7131
box 0 0 120 799
use nand4 g8051
timestamp 1386234936
transform 1 0 25539 0 1 7131
box 0 0 144 799
use nand2 g8147
timestamp 1386234792
transform 1 0 25683 0 1 7131
box 0 0 96 799
use nand2 g7955
timestamp 1386234792
transform 1 0 25779 0 1 7131
box 0 0 96 799
use nand4 g8030
timestamp 1386234936
transform 1 0 25875 0 1 7131
box 0 0 144 799
use and2 g8217
timestamp 1386234845
transform 1 0 26019 0 1 7131
box 0 0 120 799
use nand2 g8353
timestamp 1386234792
transform 1 0 26139 0 1 7131
box 0 0 96 799
use inv g8248
timestamp 1386238110
transform 1 0 26235 0 1 7131
box 0 0 120 799
use nand2 g8114
timestamp 1386234792
transform 1 0 26355 0 1 7131
box 0 0 96 799
use nand2 g8174
timestamp 1386234792
transform 1 0 26451 0 1 7131
box 0 0 96 799
use nand2 g8305
timestamp 1386234792
transform 1 0 26547 0 1 7131
box 0 0 96 799
use nor2 g8241
timestamp 1386235306
transform 1 0 26643 0 1 7131
box 0 0 120 799
use nand2 g8067
timestamp 1386234792
transform 1 0 26763 0 1 7131
box 0 0 96 799
use nand2 g7990
timestamp 1386234792
transform 1 0 26859 0 1 7131
box 0 0 96 799
use nand3 g8158
timestamp 1386234893
transform 1 0 26955 0 1 7131
box 0 0 120 799
use nand2 g8063
timestamp 1386234792
transform 1 0 27075 0 1 7131
box 0 0 96 799
use inv g8257
timestamp 1386238110
transform 1 0 27171 0 1 7131
box 0 0 120 799
use nand2 Op2Sel_91_0_93_
timestamp 1386234792
transform 1 0 27291 0 1 7131
box 0 0 96 799
use rowcrosser Op2Sel_91_1_93_
timestamp 1386086759
transform 1 0 27387 0 1 7131
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27435 0 1 7131
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 1162
box 0 0 1464 799
use nor2 stateSub_reg_91_0_93_
timestamp 1386235306
transform 1 0 1587 0 1 1162
box 0 0 120 799
use scandtype g8352
timestamp 1386241841
transform 1 0 1707 0 1 1162
box 0 0 624 799
use inv g8150
timestamp 1386238110
transform 1 0 2331 0 1 1162
box 0 0 120 799
use nand2 g8020
timestamp 1386234792
transform 1 0 2451 0 1 1162
box 0 0 96 799
use nand2 g8178
timestamp 1386234792
transform 1 0 2547 0 1 1162
box 0 0 96 799
use and2 state_reg_91_1_93_
timestamp 1386234845
transform 1 0 2643 0 1 1162
box 0 0 120 799
use scandtype g8250
timestamp 1386241841
transform 1 0 2763 0 1 1162
box 0 0 624 799
use inv g8148
timestamp 1386238110
transform 1 0 3387 0 1 1162
box 0 0 120 799
use nor2 g7976
timestamp 1386235306
transform 1 0 3507 0 1 1162
box 0 0 120 799
use nand2 g8211
timestamp 1386234792
transform 1 0 3627 0 1 1162
box 0 0 96 799
use inv g8196
timestamp 1386238110
transform 1 0 3723 0 1 1162
box 0 0 120 799
use inv g8175
timestamp 1386238110
transform 1 0 3843 0 1 1162
box 0 0 120 799
use and2 g8078
timestamp 1386234845
transform 1 0 3963 0 1 1162
box 0 0 120 799
use nand2 g8093
timestamp 1386234792
transform 1 0 4083 0 1 1162
box 0 0 96 799
use nand2 g8104
timestamp 1386234792
transform 1 0 4179 0 1 1162
box 0 0 96 799
use inv g8307
timestamp 1386238110
transform 1 0 4275 0 1 1162
box 0 0 120 799
use inv g8335
timestamp 1386238110
transform 1 0 4395 0 1 1162
box 0 0 120 799
use nand2 g8160
timestamp 1386234792
transform 1 0 4515 0 1 1162
box 0 0 96 799
use nand2 g8076
timestamp 1386234792
transform 1 0 4611 0 1 1162
box 0 0 96 799
use nand2 g8224
timestamp 1386234792
transform 1 0 4707 0 1 1162
box 0 0 96 799
use nand2 g8161
timestamp 1386234792
transform 1 0 4803 0 1 1162
box 0 0 96 799
use and2 StatusReg_reg_91_2_93_
timestamp 1386234845
transform 1 0 4899 0 1 1162
box 0 0 120 799
use scandtype g8094
timestamp 1386241841
transform 1 0 5019 0 1 1162
box 0 0 624 799
use nand3 g8037
timestamp 1386234893
transform 1 0 5643 0 1 1162
box 0 0 120 799
use nand2 g8121
timestamp 1386234792
transform 1 0 5763 0 1 1162
box 0 0 96 799
use nand2 g8266
timestamp 1386234792
transform 1 0 5859 0 1 1162
box 0 0 96 799
use nand2 g8189
timestamp 1386234792
transform 1 0 5955 0 1 1162
box 0 0 96 799
use nand2 g8125
timestamp 1386234792
transform 1 0 6051 0 1 1162
box 0 0 96 799
use nand3 g8297
timestamp 1386234893
transform 1 0 6147 0 1 1162
box 0 0 120 799
use mux2 g8232
timestamp 1386235218
transform 1 0 6267 0 1 1162
box 0 0 192 799
use nand2 g8152
timestamp 1386234792
transform 1 0 6459 0 1 1162
box 0 0 96 799
use nand4 g8303
timestamp 1386234936
transform 1 0 6555 0 1 1162
box 0 0 144 799
use nand2 g8328
timestamp 1386234792
transform 1 0 6699 0 1 1162
box 0 0 96 799
use nand2 g8080
timestamp 1386234792
transform 1 0 6795 0 1 1162
box 0 0 96 799
use nand2 g7997
timestamp 1386234792
transform 1 0 6891 0 1 1162
box 0 0 96 799
use nand4 g8267
timestamp 1386234936
transform 1 0 6987 0 1 1162
box 0 0 144 799
use and2 g8282
timestamp 1386234845
transform 1 0 7131 0 1 1162
box 0 0 120 799
use nand2 g8274
timestamp 1386234792
transform 1 0 7251 0 1 1162
box 0 0 96 799
use nand2 g8236
timestamp 1386234792
transform 1 0 7347 0 1 1162
box 0 0 96 799
use nand2 g8101
timestamp 1386234792
transform 1 0 7443 0 1 1162
box 0 0 96 799
use nand2 g8011
timestamp 1386234792
transform 1 0 7539 0 1 1162
box 0 0 96 799
use nand4 g8185
timestamp 1386234936
transform 1 0 7635 0 1 1162
box 0 0 144 799
use inv g8255
timestamp 1386238110
transform 1 0 7779 0 1 1162
box 0 0 120 799
use nand2 g8086
timestamp 1386234792
transform 1 0 7899 0 1 1162
box 0 0 96 799
use nand2 g8301
timestamp 1386234792
transform 1 0 7995 0 1 1162
box 0 0 96 799
use nor2 g7962
timestamp 1386235306
transform 1 0 8091 0 1 1162
box 0 0 120 799
use nand4 g8192
timestamp 1386234936
transform 1 0 8211 0 1 1162
box 0 0 144 799
use inv g7988
timestamp 1386238110
transform 1 0 8355 0 1 1162
box 0 0 120 799
use nand2 g8292
timestamp 1386234792
transform 1 0 8475 0 1 1162
box 0 0 96 799
use inv g8254
timestamp 1386238110
transform 1 0 8571 0 1 1162
box 0 0 120 799
use nor2 g8116
timestamp 1386235306
transform 1 0 8691 0 1 1162
box 0 0 120 799
use nand3 g8166
timestamp 1386234893
transform 1 0 8811 0 1 1162
box 0 0 120 799
use nand2 g8145
timestamp 1386234792
transform 1 0 8931 0 1 1162
box 0 0 96 799
use nand3 g8001
timestamp 1386234893
transform 1 0 9027 0 1 1162
box 0 0 120 799
use nand4 g8014
timestamp 1386234936
transform 1 0 9147 0 1 1162
box 0 0 144 799
use nand2 g8315
timestamp 1386234792
transform 1 0 9291 0 1 1162
box 0 0 96 799
use nand2 g7998
timestamp 1386234792
transform 1 0 9387 0 1 1162
box 0 0 96 799
use nand4 g8228
timestamp 1386234936
transform 1 0 9483 0 1 1162
box 0 0 144 799
use nand2 g7987
timestamp 1386234792
transform 1 0 9627 0 1 1162
box 0 0 96 799
use and2 g8072
timestamp 1386234845
transform 1 0 9723 0 1 1162
box 0 0 120 799
use nor2 g7966
timestamp 1386235306
transform 1 0 9843 0 1 1162
box 0 0 120 799
use nand3 g8279
timestamp 1386234893
transform 1 0 9963 0 1 1162
box 0 0 120 799
use nor2 g8105
timestamp 1386235306
transform 1 0 10083 0 1 1162
box 0 0 120 799
use nand2 g8259
timestamp 1386234792
transform 1 0 10203 0 1 1162
box 0 0 96 799
use inv g8129
timestamp 1386238110
transform 1 0 10299 0 1 1162
box 0 0 120 799
use and2 g8122
timestamp 1386234845
transform 1 0 10419 0 1 1162
box 0 0 120 799
use and2 g8059
timestamp 1386234845
transform 1 0 10539 0 1 1162
box 0 0 120 799
use nor2 g8062
timestamp 1386235306
transform 1 0 10659 0 1 1162
box 0 0 120 799
use nand2 g8097
timestamp 1386234792
transform 1 0 10779 0 1 1162
box 0 0 96 799
use nand3 g8025
timestamp 1386234893
transform 1 0 10875 0 1 1162
box 0 0 120 799
use nor2 g8247
timestamp 1386235306
transform 1 0 10995 0 1 1162
box 0 0 120 799
use nand2 IntStatus_reg
timestamp 1386234792
transform 1 0 11115 0 1 1162
box 0 0 96 799
use scanreg g8263
timestamp 1386241447
transform 1 0 11211 0 1 1162
box 0 0 720 799
use rowcrosser SysBus_91_0_93_
timestamp 1386086759
transform 1 0 11931 0 1 1162
box 0 0 48 799
use nand2 g8131
timestamp 1386234792
transform 1 0 11979 0 1 1162
box 0 0 96 799
use nand2 g8256
timestamp 1386234792
transform 1 0 12075 0 1 1162
box 0 0 96 799
use inv g8087
timestamp 1386238110
transform 1 0 12171 0 1 1162
box 0 0 120 799
use and2 g8322
timestamp 1386234845
transform 1 0 12291 0 1 1162
box 0 0 120 799
use inv g8286
timestamp 1386238110
transform 1 0 12411 0 1 1162
box 0 0 120 799
use and2 g7991
timestamp 1386234845
transform 1 0 12531 0 1 1162
box 0 0 120 799
use inv g8137
timestamp 1386238110
transform 1 0 12651 0 1 1162
box 0 0 120 799
use nand2 g8201
timestamp 1386234792
transform 1 0 12771 0 1 1162
box 0 0 96 799
use and2 g8331
timestamp 1386234845
transform 1 0 12867 0 1 1162
box 0 0 120 799
use nand2 g8242
timestamp 1386234792
transform 1 0 12987 0 1 1162
box 0 0 96 799
use nand2 g8207
timestamp 1386234792
transform 1 0 13083 0 1 1162
box 0 0 96 799
use nor2 g8044
timestamp 1386235306
transform 1 0 13179 0 1 1162
box 0 0 120 799
use nand3 g8006
timestamp 1386234893
transform 1 0 13299 0 1 1162
box 0 0 120 799
use nand4 g8173
timestamp 1386234936
transform 1 0 13419 0 1 1162
box 0 0 144 799
use nand2 g7983
timestamp 1386234792
transform 1 0 13563 0 1 1162
box 0 0 96 799
use nand2 g8157
timestamp 1386234792
transform 1 0 13659 0 1 1162
box 0 0 96 799
use nor2 g8325
timestamp 1386235306
transform 1 0 13755 0 1 1162
box 0 0 120 799
use nor2 g8040
timestamp 1386235306
transform 1 0 13875 0 1 1162
box 0 0 120 799
use nand2 g8068
timestamp 1386234792
transform 1 0 13995 0 1 1162
box 0 0 96 799
use nor2 g8140
timestamp 1386235306
transform 1 0 14091 0 1 1162
box 0 0 120 799
use nand3 g8141
timestamp 1386234893
transform 1 0 14211 0 1 1162
box 0 0 120 799
use nand2 g8210
timestamp 1386234792
transform 1 0 14331 0 1 1162
box 0 0 96 799
use nor2 g8003
timestamp 1386235306
transform 1 0 14427 0 1 1162
box 0 0 120 799
use nand2 g8317
timestamp 1386234792
transform 1 0 14547 0 1 1162
box 0 0 96 799
use and2 g8203
timestamp 1386234845
transform 1 0 14643 0 1 1162
box 0 0 120 799
use inv g8065
timestamp 1386238110
transform 1 0 14763 0 1 1162
box 0 0 120 799
use nand2 g8113
timestamp 1386234792
transform 1 0 14883 0 1 1162
box 0 0 96 799
use and2 g7977
timestamp 1386234845
transform 1 0 14979 0 1 1162
box 0 0 120 799
use nand4 g8070
timestamp 1386234936
transform 1 0 15099 0 1 1162
box 0 0 144 799
use nand2 g8323
timestamp 1386234792
transform 1 0 15243 0 1 1162
box 0 0 96 799
use nand2 g8309
timestamp 1386234792
transform 1 0 15339 0 1 1162
box 0 0 96 799
use nand2 g8038
timestamp 1386234792
transform 1 0 15435 0 1 1162
box 0 0 96 799
use and2 g8233
timestamp 1386234845
transform 1 0 15531 0 1 1162
box 0 0 120 799
use and2 IRQ2_reg
timestamp 1386234845
transform 1 0 15651 0 1 1162
box 0 0 120 799
use scandtype g7980
timestamp 1386241841
transform 1 0 15771 0 1 1162
box 0 0 624 799
use nand4 g8151
timestamp 1386234936
transform 1 0 16395 0 1 1162
box 0 0 144 799
use inv g8138
timestamp 1386238110
transform 1 0 16539 0 1 1162
box 0 0 120 799
use nand3 g7968
timestamp 1386234893
transform 1 0 16659 0 1 1162
box 0 0 120 799
use nand3 g8188
timestamp 1386234893
transform 1 0 16779 0 1 1162
box 0 0 120 799
use and2 g8176
timestamp 1386234845
transform 1 0 16899 0 1 1162
box 0 0 120 799
use nor2 g8172
timestamp 1386235306
transform 1 0 17019 0 1 1162
box 0 0 120 799
use nand2 g8026
timestamp 1386234792
transform 1 0 17139 0 1 1162
box 0 0 96 799
use inv g8162
timestamp 1386238110
transform 1 0 17235 0 1 1162
box 0 0 120 799
use and2 g8031
timestamp 1386234845
transform 1 0 17355 0 1 1162
box 0 0 120 799
use nor2 g8095
timestamp 1386235306
transform 1 0 17475 0 1 1162
box 0 0 120 799
use nand3 g8008
timestamp 1386234893
transform 1 0 17595 0 1 1162
box 0 0 120 799
use nor2 g8013
timestamp 1386235306
transform 1 0 17715 0 1 1162
box 0 0 120 799
use nand2 g8299
timestamp 1386234792
transform 1 0 17835 0 1 1162
box 0 0 96 799
use nand2 g8126
timestamp 1386234792
transform 1 0 17931 0 1 1162
box 0 0 96 799
use nand2 g7984
timestamp 1386234792
transform 1 0 18027 0 1 1162
box 0 0 96 799
use nand2 g8326
timestamp 1386234792
transform 1 0 18123 0 1 1162
box 0 0 96 799
use and2 IRQ1_reg
timestamp 1386234845
transform 1 0 18219 0 1 1162
box 0 0 120 799
use scandtype g8329
timestamp 1386241841
transform 1 0 18339 0 1 1162
box 0 0 624 799
use inv g7986
timestamp 1386238110
transform 1 0 18963 0 1 1162
box 0 0 120 799
use nand2 g8205
timestamp 1386234792
transform 1 0 19083 0 1 1162
box 0 0 96 799
use nor2 g8339
timestamp 1386235306
transform 1 0 19179 0 1 1162
box 0 0 120 799
use nand2 g8164
timestamp 1386234792
transform 1 0 19299 0 1 1162
box 0 0 96 799
use nand2 g8017
timestamp 1386234792
transform 1 0 19395 0 1 1162
box 0 0 96 799
use nand3 g8165
timestamp 1386234893
transform 1 0 19491 0 1 1162
box 0 0 120 799
use and2 g8010
timestamp 1386234845
transform 1 0 19611 0 1 1162
box 0 0 120 799
use nand2 g8260
timestamp 1386234792
transform 1 0 19731 0 1 1162
box 0 0 96 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 19827 0 1 1162
box 0 0 48 799
use nor2 g8245
timestamp 1386235306
transform 1 0 19875 0 1 1162
box 0 0 120 799
use nor2 g8034
timestamp 1386235306
transform 1 0 19995 0 1 1162
box 0 0 120 799
use nor2 g8351
timestamp 1386235306
transform 1 0 20115 0 1 1162
box 0 0 120 799
use inv g8215
timestamp 1386238110
transform 1 0 20235 0 1 1162
box 0 0 120 799
use nand3 g8239
timestamp 1386234893
transform 1 0 20355 0 1 1162
box 0 0 120 799
use nand2 g8079
timestamp 1386234792
transform 1 0 20475 0 1 1162
box 0 0 96 799
use nand2 g7999
timestamp 1386234792
transform 1 0 20571 0 1 1162
box 0 0 96 799
use nand4 g8288
timestamp 1386234936
transform 1 0 20667 0 1 1162
box 0 0 144 799
use nand2 g8007
timestamp 1386234792
transform 1 0 20811 0 1 1162
box 0 0 96 799
use nor2 g8262
timestamp 1386235306
transform 1 0 20907 0 1 1162
box 0 0 120 799
use and2 g8311
timestamp 1386234845
transform 1 0 21027 0 1 1162
box 0 0 120 799
use and2 g7965
timestamp 1386234845
transform 1 0 21147 0 1 1162
box 0 0 120 799
use nand3 g8109
timestamp 1386234893
transform 1 0 21267 0 1 1162
box 0 0 120 799
use inv g8085
timestamp 1386238110
transform 1 0 21387 0 1 1162
box 0 0 120 799
use nand4 g8298
timestamp 1386234936
transform 1 0 21507 0 1 1162
box 0 0 144 799
use xor2 g8346
timestamp 1386237344
transform 1 0 21651 0 1 1162
box 0 0 192 799
use inv g8021
timestamp 1386238110
transform 1 0 21843 0 1 1162
box 0 0 120 799
use nand3 g7961
timestamp 1386234893
transform 1 0 21963 0 1 1162
box 0 0 120 799
use nand4 g8184
timestamp 1386234936
transform 1 0 22083 0 1 1162
box 0 0 144 799
use nand4 g8132
timestamp 1386234936
transform 1 0 22227 0 1 1162
box 0 0 144 799
use nand3 g8219
timestamp 1386234893
transform 1 0 22371 0 1 1162
box 0 0 120 799
use nand2 g8330
timestamp 1386234792
transform 1 0 22491 0 1 1162
box 0 0 96 799
use nand2 g8061
timestamp 1386234792
transform 1 0 22587 0 1 1162
box 0 0 96 799
use rowcrosser nWE
timestamp 1386086759
transform 1 0 22683 0 1 1162
box 0 0 48 799
use nand2 g8258
timestamp 1386234792
transform 1 0 22731 0 1 1162
box 0 0 96 799
use and2 g8115
timestamp 1386234845
transform 1 0 22827 0 1 1162
box 0 0 120 799
use and2 g8202
timestamp 1386234845
transform 1 0 22947 0 1 1162
box 0 0 120 799
use nand2 g7973
timestamp 1386234792
transform 1 0 23067 0 1 1162
box 0 0 96 799
use nand4 g8208
timestamp 1386234936
transform 1 0 23163 0 1 1162
box 0 0 144 799
use nand2 g8156
timestamp 1386234792
transform 1 0 23307 0 1 1162
box 0 0 96 799
use nand2 g8231
timestamp 1386234792
transform 1 0 23403 0 1 1162
box 0 0 96 799
use inv g7992
timestamp 1386238110
transform 1 0 23499 0 1 1162
box 0 0 120 799
use nand4 g8179
timestamp 1386234936
transform 1 0 23619 0 1 1162
box 0 0 144 799
use nand2 g8022
timestamp 1386234792
transform 1 0 23763 0 1 1162
box 0 0 96 799
use nand3 g8193
timestamp 1386234893
transform 1 0 23859 0 1 1162
box 0 0 120 799
use nor2 g8071
timestamp 1386235306
transform 1 0 23979 0 1 1162
box 0 0 120 799
use inv g8285
timestamp 1386238110
transform 1 0 24099 0 1 1162
box 0 0 120 799
use nand2 g8083
timestamp 1386234792
transform 1 0 24219 0 1 1162
box 0 0 96 799
use nand2 g8204
timestamp 1386234792
transform 1 0 24315 0 1 1162
box 0 0 96 799
use nand2 g8053
timestamp 1386234792
transform 1 0 24411 0 1 1162
box 0 0 96 799
use nor2 state_reg_91_0_93_
timestamp 1386235306
transform 1 0 24507 0 1 1162
box 0 0 120 799
use scandtype g8000
timestamp 1386241841
transform 1 0 24627 0 1 1162
box 0 0 624 799
use inv g8142
timestamp 1386238110
transform 1 0 25251 0 1 1162
box 0 0 120 799
use inv g8302
timestamp 1386238110
transform 1 0 25371 0 1 1162
box 0 0 120 799
use nand2 stateSub_reg_91_1_93_
timestamp 1386234792
transform 1 0 25491 0 1 1162
box 0 0 96 799
use scandtype g8075
timestamp 1386241841
transform 1 0 25587 0 1 1162
box 0 0 624 799
use and2 g7994
timestamp 1386234845
transform 1 0 26211 0 1 1162
box 0 0 120 799
use nand4 g8197
timestamp 1386234936
transform 1 0 26331 0 1 1162
box 0 0 144 799
use nand2 g8032
timestamp 1386234792
transform 1 0 26475 0 1 1162
box 0 0 96 799
use nand4 g8316
timestamp 1386234936
transform 1 0 26571 0 1 1162
box 0 0 144 799
use nor2 g8043
timestamp 1386235306
transform 1 0 26715 0 1 1162
box 0 0 120 799
use and2 AluOR_91_1_93_
timestamp 1386234845
transform 1 0 26835 0 1 1162
box 0 0 120 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27435 0 1 1162
box 0 0 320 799
<< labels >>
rlabel m2contact 27537 8091 27537 8091 6 Flags[0]
rlabel m2contact 27537 7947 27537 7947 6 Flags[0]
rlabel m2contact 27513 8043 27513 8043 6 CFlag
rlabel m2contact 27513 7947 27513 7947 6 CFlag
rlabel m2contact 27489 8115 27489 8115 6 Flags[3]
rlabel m2contact 27489 8019 27489 8019 6 Flags[3]
rlabel m2contact 27465 8019 27465 8019 6 Flags[2]
rlabel m2contact 27465 7995 27465 7995 6 Flags[2]
rlabel m2contact 27441 8235 27441 8235 6 Flags[1]
rlabel m2contact 27441 7971 27441 7971 6 Flags[1]
rlabel m2contact 27417 8139 27417 8139 6 StatusRegEn
rlabel m2contact 27309 8139 27309 8139 6 StatusRegEn
rlabel m2contact 27249 8187 27249 8187 6 LrSel
rlabel m2contact 27057 8139 27057 8139 6 MemEn
rlabel m2contact 26121 8067 26121 8067 6 ALE
rlabel m2contact 25629 8211 25629 8211 6 StatusReg[3]
rlabel m2contact 24777 7995 24777 7995 6 StatusReg[2]
rlabel m2contact 24561 8091 24561 8091 6 Flags[0]
rlabel m2contact 23925 8091 23925 8091 6 StatusReg[1]
rlabel m2contact 23073 8043 23073 8043 6 StatusReg[0]
rlabel m2contact 22353 8043 22353 8043 6 StatusReg[0]
rlabel m2contact 22221 8043 22221 8043 6 AluEn
rlabel m2contact 21369 8163 21369 8163 6 AluWe
rlabel m2contact 20517 8259 20517 8259 6 Op2Sel[1]
rlabel metal2 20235 7971 20235 7971 6 Op2Sel[0]
rlabel m2contact 20217 7971 20217 7971 6 Op2Sel[0]
rlabel m2contact 19617 8019 19617 8019 6 Flags[2]
rlabel m2contact 19257 7971 19257 7971 6 PcSel[0]
rlabel m2contact 18921 8283 18921 8283 6 PcEn
rlabel m2contact 18813 8019 18813 8019 6 Op1Sel
rlabel m2contact 18789 8283 18789 8283 6 PcEn
rlabel m2contact 18681 8235 18681 8235 6 Flags[1]
rlabel m2contact 18105 7947 18105 7947 6 CFlag
rlabel m2contact 17109 8235 17109 8235 6 WdSel
rlabel metal2 16899 7947 16899 7947 6 PcWe
rlabel m2contact 16881 7947 16881 7947 6 PcWe
rlabel m2contact 16377 7947 16377 7947 6 PcSel[1]
rlabel metal2 15963 8283 15963 8283 6 PcSel[2]
rlabel m2contact 15945 8283 15945 8283 6 PcSel[2]
rlabel m2contact 15609 8259 15609 8259 6 Op2Sel[1]
rlabel m2contact 15381 7947 15381 7947 6 PcSel[1]
rlabel m2contact 14817 8235 14817 8235 6 WdSel
rlabel m2contact 14673 8211 14673 8211 6 StatusReg[3]
rlabel m2contact 14529 7971 14529 7971 6 PcSel[0]
rlabel m2contact 14145 7971 14145 7971 4 LrWe
rlabel m2contact 13641 8019 13641 8019 4 Op1Sel
rlabel m2contact 12921 8091 12921 8091 4 StatusReg[1]
rlabel m2contact 12837 8091 12837 8091 4 LrEn
rlabel m2contact 12801 7971 12801 7971 4 LrWe
rlabel m2contact 11937 8187 11937 8187 4 LrSel
rlabel m2contact 11649 8043 11649 8043 4 AluEn
rlabel m2contact 11073 8043 11073 8043 4 nME
rlabel m2contact 10245 7971 10245 7971 4 ImmSel
rlabel metal2 9963 8187 9963 8187 4 IrWe
rlabel m2contact 9945 8187 9945 8187 4 IrWe
rlabel m2contact 9825 8163 9825 8163 4 AluWe
rlabel m2contact 9345 8139 9345 8139 4 MemEn
rlabel m2contact 8481 7971 8481 7971 4 ImmSel
rlabel m2contact 7653 8139 7653 8139 4 OpcodeCondIn[7]
rlabel m2contact 6993 7971 6993 7971 4 OpcodeCondIn[2]
rlabel metal2 6987 8163 6987 8163 4 OpcodeCondIn[6]
rlabel m2contact 6969 8163 6969 8163 4 OpcodeCondIn[6]
rlabel m2contact 6681 7995 6681 7995 4 StatusReg[2]
rlabel m2contact 6585 7995 6585 7995 4 OpcodeCondIn[0]
rlabel metal2 6003 8163 6003 8163 4 OpcodeCondIn[5]
rlabel m2contact 5985 8163 5985 8163 4 OpcodeCondIn[5]
rlabel m2contact 5529 8115 5529 8115 4 Flags[3]
rlabel m2contact 5061 8115 5061 8115 4 OpcodeCondIn[4]
rlabel m2contact 4737 8115 4737 8115 4 OpcodeCondIn[4]
rlabel m2contact 4197 8115 4197 8115 4 OpcodeCondIn[3]
rlabel m2contact 4161 7971 4161 7971 4 OpcodeCondIn[2]
rlabel m2contact 4089 8139 4089 8139 4 OpcodeCondIn[7]
rlabel m2contact 2961 8091 2961 8091 4 LrEn
rlabel m2contact 2469 8091 2469 8091 4 OpcodeCondIn[1]
rlabel m2contact 2433 7995 2433 7995 4 OpcodeCondIn[0]
rlabel m2contact 2217 8115 2217 8115 4 OpcodeCondIn[3]
rlabel m2contact 2145 8019 2145 8019 4 Op1Sel
rlabel m2contact 1713 8091 1713 8091 4 OpcodeCondIn[1]
rlabel m2contact 27441 6754 27441 6754 6 RwSel[0]
rlabel m2contact 27441 2002 27441 2002 6 RwSel[0]
rlabel m2contact 27417 2530 27417 2530 6 RwSel[1]
rlabel m2contact 27417 1978 27417 1978 6 RwSel[1]
rlabel m2contact 27417 4018 27417 4018 6 StatusRegEn
rlabel m2contact 27369 6490 27369 6490 6 n_56
rlabel m2contact 27345 2074 27345 2074 6 n_42
rlabel m2contact 27321 4426 27321 4426 6 state[0]
rlabel m2contact 27201 6202 27201 6202 6 n_317
rlabel m2contact 27153 6730 27153 6730 6 n_167
rlabel m2contact 27129 4690 27129 4690 6 n_267
rlabel m2contact 27105 5650 27105 5650 6 n_166
rlabel m2contact 27057 5506 27057 5506 6 n_45
rlabel m2contact 27057 4522 27057 4522 6 n_45
rlabel m2contact 27033 4042 27033 4042 6 n_316
rlabel m2contact 27009 5794 27009 5794 6 n_180
rlabel m2contact 26985 4402 26985 4402 6 n_278
rlabel m2contact 26961 5914 26961 5914 6 n_215
rlabel m2contact 26961 2842 26961 2842 6 n_215
rlabel m2contact 26937 5314 26937 5314 6 n_281
rlabel m2contact 26913 4306 26913 4306 6 n_282
rlabel m2contact 26889 2578 26889 2578 6 n_284
rlabel m2contact 26865 4618 26865 4618 6 n_233
rlabel m2contact 26841 4282 26841 4282 6 n_128
rlabel m2contact 26817 4522 26817 4522 6 n_45
rlabel m2contact 26817 4546 26817 4546 6 n_102
rlabel m2contact 26793 4594 26793 4594 6 n_237
rlabel m2contact 26769 5002 26769 5002 6 OpcodeCondIn[7]
rlabel m2contact 26745 2842 26745 2842 6 n_215
rlabel m2contact 26745 2866 26745 2866 6 n_232
rlabel m2contact 26697 3106 26697 3106 6 OpcodeCondIn[0]
rlabel m2contact 26673 3874 26673 3874 6 n_17
rlabel m2contact 26673 4066 26673 4066 6 OpcodeCondIn[1]
rlabel m2contact 26649 4498 26649 4498 6 n_274
rlabel m2contact 26649 4450 26649 4450 6 n_274
rlabel m2contact 26625 3946 26625 3946 6 n_196
rlabel m2contact 26601 5218 26601 5218 6 n_171
rlabel m2contact 26577 6514 26577 6514 6 n_124
rlabel m2contact 26553 3346 26553 3346 6 n_117
rlabel m2contact 26529 2266 26529 2266 6 n_96
rlabel m2contact 26529 3010 26529 3010 6 n_253
rlabel m2contact 26505 4450 26505 4450 6 n_274
rlabel m2contact 26505 4474 26505 4474 6 n_84
rlabel m2contact 26481 3514 26481 3514 6 n_212
rlabel m2contact 26457 4978 26457 4978 6 n_241
rlabel m2contact 26457 4330 26457 4330 6 n_241
rlabel m2contact 26433 6994 26433 6994 6 n_31
rlabel m2contact 26433 5890 26433 5890 6 stateSub[2]
rlabel m2contact 26409 4330 26409 4330 6 n_241
rlabel m2contact 26409 4354 26409 4354 6 OpcodeCondIn[3]
rlabel m2contact 26385 7066 26385 7066 6 n_16
rlabel m2contact 26385 5266 26385 5266 6 n_323
rlabel m2contact 26361 5074 26361 5074 6 n_243
rlabel m2contact 26313 2554 26313 2554 6 n_373
rlabel m2contact 26313 5914 26313 5914 6 n_215
rlabel m2contact 26265 3706 26265 3706 6 n_359
rlabel m2contact 26265 3898 26265 3898 6 OpcodeCondIn[5]
rlabel m2contact 26241 3634 26241 3634 6 n_268
rlabel m2contact 26217 2242 26217 2242 6 n_109
rlabel m2contact 26193 4258 26193 4258 6 n_162
rlabel m2contact 26169 4090 26169 4090 6 n_151
rlabel m2contact 26097 4882 26097 4882 6 stateSub[1]
rlabel m2contact 26073 4210 26073 4210 6 n_204
rlabel m2contact 26049 6682 26049 6682 6 n_304
rlabel m2contact 26049 4162 26049 4162 6 n_309
rlabel m2contact 26001 4570 26001 4570 6 Rs1Sel[0]
rlabel m2contact 25977 5266 25977 5266 6 n_323
rlabel m2contact 25953 6178 25953 6178 6 n_338
rlabel m2contact 25929 4834 25929 4834 6 n_234
rlabel m2contact 25905 5122 25905 5122 6 n_92
rlabel m2contact 25857 6466 25857 6466 6 n_192
rlabel m2contact 25833 3802 25833 3802 6 stateSub[0]
rlabel m2contact 25809 2482 25809 2482 6 n_136
rlabel m2contact 25785 6970 25785 6970 6 n_172
rlabel m2contact 25785 3730 25785 3730 6 n_172
rlabel m2contact 25761 2002 25761 2002 6 n_294
rlabel m2contact 25737 5890 25737 5890 6 stateSub[2]
rlabel m2contact 25713 6898 25713 6898 6 n_217
rlabel m2contact 25689 4570 25689 4570 6 n_369
rlabel m2contact 25665 4570 25665 4570 6 n_369
rlabel m2contact 25641 6010 25641 6010 6 n_23
rlabel m2contact 25617 4642 25617 4642 6 n_331
rlabel m2contact 25593 2290 25593 2290 6 n_190
rlabel m2contact 25569 6970 25569 6970 6 n_172
rlabel m2contact 25569 6946 25569 6946 6 n_40
rlabel m2contact 25545 7042 25545 7042 6 n_499
rlabel m2contact 25521 2914 25521 2914 6 StatusReg[2]
rlabel m2contact 25521 5170 25521 5170 6 n_47
rlabel m2contact 25473 4930 25473 4930 6 n_26
rlabel m2contact 25449 4018 25449 4018 6 StatusRegEn
rlabel m2contact 25449 4090 25449 4090 6 n_151
rlabel m2contact 25425 5626 25425 5626 6 n_160
rlabel m2contact 25425 4186 25425 4186 6 n_160
rlabel m2contact 25401 4186 25401 4186 6 n_160
rlabel m2contact 25401 4234 25401 4234 6 n_211
rlabel m2contact 25377 5602 25377 5602 6 n_362
rlabel m2contact 25377 4522 25377 4522 6 n_362
rlabel m2contact 25353 4090 25353 4090 6 n_151
rlabel m2contact 25329 4522 25329 4522 6 n_362
rlabel m2contact 25329 5242 25329 5242 6 n_179
rlabel m2contact 25305 4570 25305 4570 6 n_181
rlabel m2contact 25305 2146 25305 2146 6 n_181
rlabel m2contact 25281 4570 25281 4570 6 n_181
rlabel m2contact 25281 3658 25281 3658 6 n_367
rlabel m2contact 25233 3058 25233 3058 6 n_157
rlabel m2contact 25209 4762 25209 4762 6 n_87
rlabel m2contact 25185 4570 25185 4570 6 n_249
rlabel m2contact 25185 4378 25185 4378 6 n_249
rlabel m2contact 25161 2962 25161 2962 6 n_387
rlabel m2contact 25137 4570 25137 4570 6 n_249
rlabel m2contact 25137 4426 25137 4426 6 state[0]
rlabel m2contact 25113 3370 25113 3370 6 n_366
rlabel m2contact 25089 6082 25089 6082 6 n_340
rlabel m2contact 25089 4930 25089 4930 6 n_26
rlabel m2contact 25041 3994 25041 3994 6 n_257
rlabel m2contact 24993 6562 24993 6562 6 n_156
rlabel m2contact 24969 4666 24969 4666 6 n_273
rlabel m2contact 24897 4594 24897 4594 6 n_237
rlabel m2contact 24849 6130 24849 6130 6 n_79
rlabel m2contact 24777 4690 24777 4690 6 n_267
rlabel m2contact 24729 2194 24729 2194 6 n_293
rlabel m2contact 24729 2338 24729 2338 6 n_107
rlabel m2contact 24705 6850 24705 6850 6 n_261
rlabel m2contact 24705 3610 24705 3610 6 n_261
rlabel m2contact 24681 2290 24681 2290 6 n_190
rlabel m2contact 24657 3802 24657 3802 6 stateSub[0]
rlabel m2contact 24633 3538 24633 3538 6 n_134
rlabel m2contact 24609 6346 24609 6346 6 n_276
rlabel m2contact 24609 2386 24609 2386 6 n_276
rlabel m2contact 24585 4450 24585 4450 6 n_370
rlabel m2contact 24561 4354 24561 4354 6 OpcodeCondIn[3]
rlabel m2contact 24537 3610 24537 3610 6 n_261
rlabel m2contact 24537 3658 24537 3658 6 n_367
rlabel m2contact 24501 6370 24501 6370 6 n_277
rlabel m2contact 24501 4330 24501 4330 6 n_277
rlabel m2contact 24489 6634 24489 6634 6 n_209
rlabel m2contact 24465 4138 24465 4138 6 n_53
rlabel m2contact 24441 5866 24441 5866 6 n_74
rlabel m2contact 24441 4522 24441 4522 6 n_259
rlabel m2contact 24417 6226 24417 6226 6 n_138
rlabel m2contact 24393 4402 24393 4402 6 n_278
rlabel m2contact 24369 2386 24369 2386 6 n_276
rlabel m2contact 24369 2410 24369 2410 6 n_372
rlabel m2contact 24345 4330 24345 4330 6 n_277
rlabel m2contact 24345 4354 24345 4354 6 OpcodeCondIn[3]
rlabel m2contact 24321 3514 24321 3514 6 n_212
rlabel m2contact 24297 5554 24297 5554 6 n_77
rlabel m2contact 24249 2266 24249 2266 6 n_96
rlabel m2contact 24201 5002 24201 5002 6 OpcodeCondIn[7]
rlabel m2contact 24177 4570 24177 4570 6 n_280
rlabel m2contact 24153 4618 24153 4618 6 n_233
rlabel m2contact 24129 4354 24129 4354 6 OpcodeCondIn[3]
rlabel m2contact 24105 3250 24105 3250 6 n_202
rlabel m2contact 24081 2866 24081 2866 6 n_232
rlabel m2contact 24033 4402 24033 4402 6 n_291
rlabel m2contact 24033 3154 24033 3154 6 n_57
rlabel m2contact 23985 2602 23985 2602 6 n_177
rlabel m2contact 23961 4186 23961 4186 6 n_223
rlabel m2contact 23937 5218 23937 5218 6 n_171
rlabel m2contact 23913 3034 23913 3034 6 n_346
rlabel m2contact 23889 5578 23889 5578 6 n_142
rlabel m2contact 23889 5074 23889 5074 6 n_243
rlabel m2contact 23865 3250 23865 3250 6 n_202
rlabel m2contact 23841 4618 23841 4618 6 n_163
rlabel m2contact 23817 4642 23817 4642 6 n_331
rlabel m2contact 23817 4258 23817 4258 6 n_162
rlabel m2contact 23793 4882 23793 4882 6 stateSub[1]
rlabel m2contact 23793 4330 23793 4330 6 n_194
rlabel m2contact 23769 4114 23769 4114 6 n_295
rlabel m2contact 23697 2986 23697 2986 6 n_131
rlabel m2contact 23673 3682 23673 3682 6 n_322
rlabel m2contact 23649 5410 23649 5410 6 n_246
rlabel m2contact 23625 6442 23625 6442 6 n_24
rlabel m2contact 23625 2722 23625 2722 6 n_24
rlabel m2contact 23601 2386 23601 2386 6 n_381
rlabel m2contact 23577 5098 23577 5098 6 PcSel[2]
rlabel m2contact 23553 4618 23553 4618 6 n_163
rlabel m2contact 23529 2698 23529 2698 6 n_332
rlabel m2contact 23529 5674 23529 5674 6 n_275
rlabel m2contact 23505 4618 23505 4618 6 n_252
rlabel m2contact 23505 3922 23505 3922 6 n_252
rlabel m2contact 23481 6178 23481 6178 6 n_338
rlabel m2contact 23481 6154 23481 6154 6 n_153
rlabel m2contact 23457 4882 23457 4882 6 stateSub[1]
rlabel m2contact 23433 3490 23433 3490 6 n_169
rlabel m2contact 23409 3778 23409 3778 6 n_320
rlabel m2contact 23373 6178 23373 6178 6 SysBus[0]
rlabel m2contact 23373 4018 23373 4018 6 SysBus[0]
rlabel m2contact 23361 2746 23361 2746 6 n_207
rlabel m2contact 23337 2722 23337 2722 6 n_24
rlabel m2contact 23337 2746 23337 2746 6 n_207
rlabel m2contact 23313 6826 23313 6826 6 n_221
rlabel m2contact 23313 3970 23313 3970 6 n_221
rlabel m2contact 23289 3850 23289 3850 6 Rs1Sel[1]
rlabel m2contact 23289 4354 23289 4354 6 OpcodeCondIn[3]
rlabel m2contact 23265 2410 23265 2410 6 n_372
rlabel m2contact 23241 2554 23241 2554 6 n_373
rlabel m2contact 23217 4714 23217 4714 6 n_327
rlabel m2contact 23217 6370 23217 6370 6 n_277
rlabel m2contact 23181 4738 23181 4738 6 n_6
rlabel m2contact 23181 2770 23181 2770 6 n_6
rlabel m2contact 23169 5938 23169 5938 6 n_227
rlabel m2contact 23145 6802 23145 6802 6 n_93
rlabel m2contact 23121 4618 23121 4618 6 n_252
rlabel m2contact 23121 4426 23121 4426 6 state[0]
rlabel m2contact 23097 6178 23097 6178 6 SysBus[0]
rlabel m2contact 23097 6130 23097 6130 6 n_79
rlabel m2contact 23073 3226 23073 3226 6 n_250
rlabel m2contact 23049 2578 23049 2578 6 n_284
rlabel m2contact 23025 4618 23025 4618 6 n_67
rlabel m2contact 23001 4642 23001 4642 6 n_229
rlabel m2contact 23001 4354 23001 4354 6 OpcodeCondIn[3]
rlabel m2contact 22977 5050 22977 5050 6 n_22
rlabel m2contact 22977 5026 22977 5026 6 n_230
rlabel m2contact 22941 4954 22941 4954 6 n_80
rlabel m2contact 22941 3562 22941 3562 6 n_80
rlabel m2contact 22929 5530 22929 5530 6 n_314
rlabel m2contact 22905 4210 22905 4210 6 n_204
rlabel m2contact 22881 2074 22881 2074 6 n_42
rlabel m2contact 22881 2986 22881 2986 6 n_131
rlabel m2contact 22857 4906 22857 4906 6 n_49
rlabel m2contact 22833 4858 22833 4858 6 n_220
rlabel m2contact 22809 3970 22809 3970 6 n_221
rlabel m2contact 22809 6034 22809 6034 6 n_11
rlabel m2contact 22785 5458 22785 5458 6 n_147
rlabel m2contact 22761 6418 22761 6418 6 n_81
rlabel m2contact 22761 5170 22761 5170 6 n_47
rlabel m2contact 22737 6970 22737 6970 6 n_58
rlabel m2contact 22713 4018 22713 4018 6 SysBus[0]
rlabel m2contact 22689 2506 22689 2506 6 n_120
rlabel m2contact 22665 6010 22665 6010 6 n_23
rlabel m2contact 22641 4738 22641 4738 6 n_6
rlabel m2contact 22641 3802 22641 3802 6 stateSub[0]
rlabel m2contact 22617 4954 22617 4954 6 n_80
rlabel m2contact 22617 4882 22617 4882 6 stateSub[1]
rlabel m2contact 22569 5698 22569 5698 6 n_159
rlabel m2contact 22545 4162 22545 4162 6 n_309
rlabel m2contact 22521 2026 22521 2026 6 n_104
rlabel m2contact 22521 3082 22521 3082 6 OpcodeCondIn[2]
rlabel m2contact 22497 3586 22497 3586 6 n_3
rlabel m2contact 22449 3274 22449 3274 6 n_174
rlabel m2contact 22425 6274 22425 6274 6 n_186
rlabel m2contact 22401 4162 22401 4162 6 n_309
rlabel m2contact 22353 5986 22353 5986 6 StatusReg[0]
rlabel m2contact 22353 3706 22353 3706 6 n_359
rlabel m2contact 22329 4930 22329 4930 6 n_26
rlabel m2contact 22305 5074 22305 5074 6 n_243
rlabel m2contact 22281 5890 22281 5890 6 stateSub[2]
rlabel m2contact 22257 3610 22257 3610 6 state[1]
rlabel m2contact 22185 3706 22185 3706 6 n_359
rlabel m2contact 22161 5194 22161 5194 6 n_371
rlabel m2contact 22137 5290 22137 5290 6 n_354
rlabel m2contact 22065 4114 22065 4114 6 n_295
rlabel m2contact 22041 5266 22041 5266 6 n_323
rlabel m2contact 22017 3946 22017 3946 6 n_196
rlabel m2contact 21993 2002 21993 2002 6 n_294
rlabel m2contact 21945 3850 21945 3850 6 n_389
rlabel m2contact 21921 5434 21921 5434 6 n_20
rlabel m2contact 21873 5338 21873 5338 6 OpcodeCondIn[4]
rlabel m2contact 21825 5266 21825 5266 6 n_323
rlabel m2contact 21825 3178 21825 3178 6 n_323
rlabel m2contact 21801 3178 21801 3178 6 n_323
rlabel m2contact 21801 3202 21801 3202 6 n_110
rlabel m2contact 21753 2242 21753 2242 6 n_109
rlabel m2contact 21729 4954 21729 4954 6 n_187
rlabel m2contact 21729 3322 21729 3322 6 n_187
rlabel m2contact 21705 6706 21705 6706 6 n_161
rlabel m2contact 21705 4018 21705 4018 6 n_225
rlabel m2contact 21681 4954 21681 4954 6 n_187
rlabel m2contact 21681 4930 21681 4930 6 n_26
rlabel m2contact 21657 4234 21657 4234 6 n_211
rlabel m2contact 21609 6658 21609 6658 6 n_94
rlabel m2contact 21609 2818 21609 2818 6 n_193
rlabel m2contact 21585 6274 21585 6274 6 n_186
rlabel m2contact 21561 5746 21561 5746 6 n_25
rlabel m2contact 21561 3802 21561 3802 6 stateSub[0]
rlabel m2contact 21537 5866 21537 5866 6 n_74
rlabel m2contact 21537 3322 21537 3322 6 n_187
rlabel m2contact 21489 4114 21489 4114 6 n_364
rlabel m2contact 21465 2098 21465 2098 6 n_228
rlabel m2contact 21465 4786 21465 4786 6 n_88
rlabel m2contact 21441 3970 21441 3970 6 n_326
rlabel m2contact 21417 5290 21417 5290 6 n_354
rlabel m2contact 21417 6610 21417 6610 6 n_165
rlabel m2contact 21369 3850 21369 3850 6 n_389
rlabel m2contact 21369 6586 21369 6586 6 n_75
rlabel m2contact 21345 3922 21345 3922 6 n_252
rlabel m2contact 21345 5914 21345 5914 6 n_215
rlabel m2contact 21321 4450 21321 4450 6 n_370
rlabel m2contact 21321 5866 21321 5866 6 n_74
rlabel m2contact 21297 2170 21297 2170 6 n_344
rlabel m2contact 21297 5818 21297 5818 6 n_72
rlabel m2contact 21249 4738 21249 4738 6 n_83
rlabel m2contact 21249 4210 21249 4210 6 n_204
rlabel m2contact 21225 2746 21225 2746 6 n_207
rlabel m2contact 21201 4258 21201 4258 6 n_162
rlabel m2contact 21201 4162 21201 4162 6 n_309
rlabel m2contact 21177 3826 21177 3826 6 n_14
rlabel m2contact 21153 6250 21153 6250 6 n_239
rlabel m2contact 21117 5098 21117 5098 6 PcSel[2]
rlabel m2contact 21117 3850 21117 3850 6 PcSel[2]
rlabel m2contact 21105 5770 21105 5770 6 n_198
rlabel m2contact 21081 4450 21081 4450 6 n_140
rlabel m2contact 21081 2746 21081 2746 6 n_207
rlabel m2contact 21057 5506 21057 5506 6 n_45
rlabel m2contact 21033 3754 21033 3754 6 n_126
rlabel m2contact 21009 5074 21009 5074 6 n_243
rlabel m2contact 21009 3922 21009 3922 6 n_243
rlabel m2contact 20985 2266 20985 2266 6 n_96
rlabel m2contact 20961 3850 20961 3850 6 PcSel[2]
rlabel m2contact 20961 4930 20961 4930 6 n_26
rlabel m2contact 20937 4114 20937 4114 6 n_364
rlabel m2contact 20913 6346 20913 6346 6 n_276
rlabel m2contact 20889 2050 20889 2050 6 n_105
rlabel m2contact 20865 3922 20865 3922 6 n_243
rlabel m2contact 20865 4018 20865 4018 6 n_225
rlabel m2contact 20841 4762 20841 4762 6 n_87
rlabel m2contact 20841 4546 20841 4546 6 n_102
rlabel m2contact 20793 5194 20793 5194 6 n_371
rlabel m2contact 20793 4954 20793 4954 6 n_355
rlabel m2contact 20769 5146 20769 5146 6 n_158
rlabel m2contact 20745 5362 20745 5362 6 n_254
rlabel m2contact 20721 4954 20721 4954 6 n_355
rlabel m2contact 20721 4810 20721 4810 6 n_285
rlabel m2contact 20673 3274 20673 3274 6 n_174
rlabel m2contact 20649 4378 20649 4378 6 n_249
rlabel m2contact 20625 5002 20625 5002 6 OpcodeCondIn[7]
rlabel m2contact 20601 3226 20601 3226 6 n_250
rlabel m2contact 20601 4498 20601 4498 6 n_274
rlabel m2contact 20553 5722 20553 5722 6 n_307
rlabel m2contact 20529 6178 20529 6178 6 n_297
rlabel m2contact 20529 2866 20529 2866 6 n_232
rlabel m2contact 20505 4858 20505 4858 6 n_220
rlabel m2contact 20481 4954 20481 4954 6 n_65
rlabel m2contact 20481 3466 20481 3466 6 n_65
rlabel m2contact 20457 3466 20457 3466 6 n_65
rlabel m2contact 20457 3562 20457 3562 6 n_80
rlabel m2contact 20409 5386 20409 5386 6 n_13
rlabel m2contact 20385 4546 20385 4546 6 n_102
rlabel m2contact 20361 5194 20361 5194 6 n_12
rlabel m2contact 20361 2794 20361 2794 6 n_12
rlabel m2contact 20337 4114 20337 4114 6 nWE
rlabel m2contact 20313 2794 20313 2794 6 n_12
rlabel m2contact 20313 2842 20313 2842 6 n_289
rlabel m2contact 20289 5482 20289 5482 6 n_312
rlabel m2contact 20265 6394 20265 6394 6 n_286
rlabel m2contact 20265 3106 20265 3106 6 OpcodeCondIn[0]
rlabel m2contact 20217 4378 20217 4378 6 Op2Sel[0]
rlabel m2contact 20169 4858 20169 4858 6 n_123
rlabel m2contact 20145 3994 20145 3994 6 n_257
rlabel m2contact 20145 4162 20145 4162 6 n_309
rlabel m2contact 20121 4234 20121 4234 6 n_211
rlabel m2contact 20097 3802 20097 3802 6 stateSub[0]
rlabel m2contact 20061 4258 20061 4258 6 n_162
rlabel m2contact 20061 3994 20061 3994 6 n_162
rlabel m2contact 20049 6538 20049 6538 6 n_224
rlabel m2contact 20025 5986 20025 5986 6 StatusReg[0]
rlabel m2contact 20001 3058 20001 3058 6 n_157
rlabel m2contact 19977 3994 19977 3994 6 n_162
rlabel m2contact 19977 4090 19977 4090 6 n_151
rlabel m2contact 19953 5842 19953 5842 6 n_184
rlabel m2contact 19953 2434 19953 2434 6 n_184
rlabel m2contact 19929 5842 19929 5842 6 n_184
rlabel m2contact 19929 5002 19929 5002 6 OpcodeCondIn[7]
rlabel m2contact 19905 4954 19905 4954 6 n_65
rlabel m2contact 19905 2074 19905 2074 6 n_42
rlabel m2contact 19881 3754 19881 3754 6 n_126
rlabel m2contact 19857 4114 19857 4114 6 nWE
rlabel m2contact 19857 4882 19857 4882 6 stateSub[1]
rlabel m2contact 19809 4042 19809 4042 6 n_316
rlabel m2contact 19809 4114 19809 4114 6 n_302
rlabel m2contact 19785 6922 19785 6922 6 n_70
rlabel m2contact 19785 3802 19785 3802 6 stateSub[0]
rlabel m2contact 19761 3178 19761 3178 6 n_299
rlabel m2contact 19737 4954 19737 4954 6 n_99
rlabel m2contact 19737 2674 19737 2674 6 n_99
rlabel m2contact 19713 6898 19713 6898 6 n_217
rlabel m2contact 19713 6874 19713 6874 6 n_200
rlabel m2contact 19689 3850 19689 3850 6 n_141
rlabel m2contact 19665 4954 19665 4954 6 n_99
rlabel m2contact 19665 3274 19665 3274 6 n_174
rlabel m2contact 19641 5578 19641 5578 6 n_142
rlabel m2contact 19617 2938 19617 2938 6 Flags[2]
rlabel m2contact 19593 4378 19593 4378 6 Op2Sel[0]
rlabel m2contact 19569 4114 19569 4114 6 n_302
rlabel m2contact 19569 4306 19569 4306 6 n_282
rlabel m2contact 19545 6898 19545 6898 6 n_287
rlabel m2contact 19521 2794 19521 2794 6 n_501
rlabel m2contact 19521 2818 19521 2818 6 n_193
rlabel m2contact 19497 5554 19497 5554 6 n_77
rlabel m2contact 19473 4954 19473 4954 6 n_144
rlabel m2contact 19449 4378 19449 4378 6 n_28
rlabel m2contact 19449 3274 19449 3274 6 n_174
rlabel m2contact 19425 6106 19425 6106 6 n_18
rlabel m2contact 19401 4090 19401 4090 6 n_151
rlabel m2contact 19377 5962 19377 5962 6 n_9
rlabel m2contact 19353 5554 19353 5554 6 n_245
rlabel m2contact 19353 3082 19353 3082 6 OpcodeCondIn[2]
rlabel m2contact 19329 6274 19329 6274 6 n_186
rlabel m2contact 19329 4354 19329 4354 6 OpcodeCondIn[3]
rlabel m2contact 19305 6322 19305 6322 6 n_203
rlabel m2contact 19257 5842 19257 5842 6 n_332
rlabel m2contact 19257 2698 19257 2698 6 n_332
rlabel m2contact 19233 5842 19233 5842 6 n_332
rlabel m2contact 19233 4882 19233 4882 6 stateSub[1]
rlabel m2contact 19209 5722 19209 5722 6 n_307
rlabel m2contact 19209 5410 19209 5410 6 n_246
rlabel m2contact 19185 6010 19185 6010 6 n_23
rlabel m2contact 19185 4114 19185 4114 6 n_23
rlabel m2contact 19161 3370 19161 3370 6 n_366
rlabel m2contact 19161 3394 19161 3394 6 n_111
rlabel m2contact 19137 2938 19137 2938 6 Flags[2]
rlabel m2contact 19137 3082 19137 3082 6 OpcodeCondIn[2]
rlabel m2contact 19113 5578 19113 5578 6 n_142
rlabel m2contact 19113 3658 19113 3658 6 n_367
rlabel m2contact 19077 5722 19077 5722 6 n_174
rlabel m2contact 19077 3274 19077 3274 6 n_174
rlabel m2contact 19065 5794 19065 5794 6 n_180
rlabel m2contact 19041 5722 19041 5722 6 n_174
rlabel m2contact 19041 4762 19041 4762 6 n_87
rlabel m2contact 19017 3370 19017 3370 6 n_178
rlabel m2contact 18993 4114 18993 4114 6 n_23
rlabel m2contact 18993 5242 18993 5242 6 n_179
rlabel m2contact 18969 4882 18969 4882 6 stateSub[1]
rlabel m2contact 18897 2050 18897 2050 6 n_105
rlabel m2contact 18873 2938 18873 2938 6 n_378
rlabel m2contact 18849 5602 18849 5602 6 n_362
rlabel m2contact 18777 2122 18777 2122 6 n_125
rlabel m2contact 18729 6514 18729 6514 6 n_124
rlabel m2contact 18681 4114 18681 4114 6 Flags[1]
rlabel m2contact 18633 5482 18633 5482 6 n_312
rlabel m2contact 18609 4162 18609 4162 6 n_309
rlabel m2contact 18585 6682 18585 6682 6 n_304
rlabel m2contact 18537 5386 18537 5386 6 n_13
rlabel m2contact 18489 4018 18489 4018 6 n_225
rlabel m2contact 18465 4090 18465 4090 6 n_151
rlabel m2contact 18417 4498 18417 4498 6 n_274
rlabel m2contact 18393 5386 18393 5386 6 n_207
rlabel m2contact 18393 2746 18393 2746 6 n_207
rlabel m2contact 18369 4642 18369 4642 6 n_229
rlabel m2contact 18345 2074 18345 2074 6 n_42
rlabel m2contact 18321 4474 18321 4474 6 n_84
rlabel m2contact 18297 5866 18297 5866 6 n_74
rlabel m2contact 18273 5338 18273 5338 6 OpcodeCondIn[4]
rlabel m2contact 18273 4354 18273 4354 6 OpcodeCondIn[3]
rlabel m2contact 18249 5386 18249 5386 6 n_207
rlabel m2contact 18249 4090 18249 4090 6 n_151
rlabel m2contact 18177 4114 18177 4114 6 Flags[1]
rlabel m2contact 18153 3658 18153 3658 6 n_367
rlabel m2contact 18105 7018 18105 7018 6 CFlag
rlabel m2contact 18081 4210 18081 4210 6 n_204
rlabel m2contact 18057 3994 18057 3994 6 n_205
rlabel m2contact 17985 2626 17985 2626 6 n_39
rlabel m2contact 17961 6946 17961 6946 6 n_40
rlabel m2contact 17889 4114 17889 4114 6 OpcodeCondIn[6]
rlabel m2contact 17865 5386 17865 5386 6 n_325
rlabel m2contact 17817 5842 17817 5842 6 n_263
rlabel m2contact 17769 2458 17769 2458 6 n_115
rlabel m2contact 17697 4042 17697 4042 6 n_388
rlabel m2contact 17673 3082 17673 3082 6 OpcodeCondIn[2]
rlabel m2contact 17649 6274 17649 6274 6 n_186
rlabel m2contact 17625 2146 17625 2146 6 n_181
rlabel m2contact 17601 6778 17601 6778 6 n_171
rlabel m2contact 17601 5218 17601 5218 6 n_171
rlabel m2contact 17577 6778 17577 6778 6 n_171
rlabel m2contact 17577 6298 17577 6298 6 n_311
rlabel m2contact 17529 3922 17529 3922 6 IRQ2
rlabel m2contact 17529 3610 17529 3610 6 state[1]
rlabel m2contact 17505 3466 17505 3466 6 IntStatus
rlabel m2contact 17481 5482 17481 5482 6 OpcodeCondIn[2]
rlabel m2contact 17481 3082 17481 3082 6 OpcodeCondIn[2]
rlabel m2contact 17457 3514 17457 3514 6 n_212
rlabel m2contact 17433 2818 17433 2818 6 n_193
rlabel m2contact 17409 3058 17409 3058 6 n_157
rlabel m2contact 17385 5482 17385 5482 6 OpcodeCondIn[2]
rlabel m2contact 17385 3298 17385 3298 6 n_145
rlabel m2contact 17361 5602 17361 5602 6 n_60
rlabel m2contact 17361 2890 17361 2890 6 n_60
rlabel m2contact 17337 3418 17337 3418 6 n_118
rlabel m2contact 17337 2722 17337 2722 6 n_118
rlabel m2contact 17313 3970 17313 3970 6 n_326
rlabel m2contact 17313 5722 17313 5722 6 n_21
rlabel m2contact 17289 2746 17289 2746 6 n_207
rlabel m2contact 17265 5386 17265 5386 6 n_325
rlabel m2contact 17241 5434 17241 5434 6 n_20
rlabel m2contact 17217 4450 17217 4450 6 n_140
rlabel m2contact 17217 5914 17217 5914 6 n_215
rlabel m2contact 17193 4498 17193 4498 6 n_274
rlabel m2contact 17169 3394 17169 3394 6 n_111
rlabel m2contact 17145 7090 17145 7090 6 n_76
rlabel m2contact 17121 4114 17121 4114 6 OpcodeCondIn[6]
rlabel m2contact 17097 5482 17097 5482 6 n_71
rlabel m2contact 17073 4354 17073 4354 6 OpcodeCondIn[3]
rlabel m2contact 17049 6226 17049 6226 6 n_138
rlabel m2contact 17025 5146 17025 5146 6 n_158
rlabel m2contact 17001 3970 17001 3970 6 nWait
rlabel m2contact 16977 5650 16977 5650 6 n_166
rlabel m2contact 16953 2890 16953 2890 6 n_60
rlabel m2contact 16953 3058 16953 3058 6 n_157
rlabel m2contact 16929 2722 16929 2722 6 n_118
rlabel m2contact 16929 2818 16929 2818 6 n_193
rlabel m2contact 16905 6058 16905 6058 6 n_383
rlabel m2contact 16905 3130 16905 3130 6 n_383
rlabel m2contact 16881 3130 16881 3130 6 n_383
rlabel m2contact 16881 3442 16881 3442 6 PcWe
rlabel m2contact 16833 5578 16833 5578 6 n_142
rlabel m2contact 16833 2890 16833 2890 6 n_363
rlabel m2contact 16809 5146 16809 5146 6 n_236
rlabel m2contact 16809 4450 16809 4450 6 n_236
rlabel m2contact 16785 2866 16785 2866 6 n_232
rlabel m2contact 16761 3730 16761 3730 6 n_172
rlabel m2contact 16761 4474 16761 4474 6 n_84
rlabel m2contact 16737 5218 16737 5218 6 n_171
rlabel m2contact 16713 5146 16713 5146 6 n_236
rlabel m2contact 16713 4906 16713 4906 6 n_49
rlabel m2contact 16689 5890 16689 5890 6 stateSub[2]
rlabel m2contact 16689 4426 16689 4426 6 state[0]
rlabel m2contact 16665 6778 16665 6778 6 n_197
rlabel m2contact 16593 4714 16593 4714 6 n_327
rlabel m2contact 16569 2674 16569 2674 6 n_99
rlabel m2contact 16545 5578 16545 5578 6 n_315
rlabel m2contact 16521 3778 16521 3778 6 n_320
rlabel m2contact 16497 5146 16497 5146 6 n_34
rlabel m2contact 16473 7066 16473 7066 6 n_16
rlabel m2contact 16473 5794 16473 5794 6 n_266
rlabel m2contact 16425 2866 16425 2866 6 n_232
rlabel m2contact 16353 2698 16353 2698 6 n_332
rlabel m2contact 16329 4714 16329 4714 6 n_334
rlabel m2contact 16281 3922 16281 3922 6 IRQ2
rlabel m2contact 16281 6922 16281 6922 6 n_70
rlabel m2contact 16257 2074 16257 2074 6 n_42
rlabel m2contact 16233 5722 16233 5722 6 n_21
rlabel m2contact 16185 4810 16185 4810 6 n_285
rlabel m2contact 16161 3898 16161 3898 6 OpcodeCondIn[5]
rlabel m2contact 16137 2578 16137 2578 6 n_284
rlabel m2contact 16089 4810 16089 4810 6 n_219
rlabel m2contact 16065 3514 16065 3514 6 n_8
rlabel m2contact 16041 6154 16041 6154 6 n_153
rlabel m2contact 16017 5722 16017 5722 6 n_68
rlabel m2contact 15993 6922 15993 6922 6 n_116
rlabel m2contact 15945 5098 15945 5098 6 PcSel[2]
rlabel m2contact 15873 2362 15873 2362 6 n_313
rlabel m2contact 15849 5098 15849 5098 6 n_235
rlabel m2contact 15801 5026 15801 5026 6 n_230
rlabel m2contact 15777 5338 15777 5338 6 OpcodeCondIn[4]
rlabel m2contact 15729 7066 15729 7066 6 n_44
rlabel m2contact 15729 3922 15729 3922 6 n_44
rlabel m2contact 15705 6442 15705 6442 6 n_24
rlabel m2contact 15681 3922 15681 3922 6 n_44
rlabel m2contact 15681 6154 15681 6154 6 n_4
rlabel m2contact 15657 6010 15657 6010 6 n_23
rlabel m2contact 15609 3922 15609 3922 6 Op2Sel[1]
rlabel m2contact 15585 6346 15585 6346 6 n_276
rlabel m2contact 15489 4066 15489 4066 6 OpcodeCondIn[1]
rlabel m2contact 15465 5194 15465 5194 6 n_12
rlabel m2contact 15465 5890 15465 5890 6 stateSub[2]
rlabel m2contact 15441 6442 15441 6442 6 n_240
rlabel m2contact 15441 3778 15441 3778 6 n_240
rlabel m2contact 15417 3778 15417 3778 6 n_240
rlabel m2contact 15417 4090 15417 4090 6 n_151
rlabel m2contact 15393 2746 15393 2746 6 n_207
rlabel m2contact 15369 4426 15369 4426 6 state[0]
rlabel m2contact 15297 4522 15297 4522 6 n_259
rlabel m2contact 15273 5938 15273 5938 6 n_227
rlabel m2contact 15225 3922 15225 3922 6 Op2Sel[1]
rlabel m2contact 15201 3706 15201 3706 6 n_359
rlabel m2contact 15129 4402 15129 4402 6 n_291
rlabel m2contact 15057 1978 15057 1978 6 n_319
rlabel m2contact 15033 2818 15033 2818 6 n_193
rlabel m2contact 15009 6874 15009 6874 6 n_200
rlabel m2contact 14961 4714 14961 4714 6 n_334
rlabel m2contact 14937 3154 14937 3154 6 n_57
rlabel m2contact 14913 6178 14913 6178 6 n_297
rlabel m2contact 14889 4066 14889 4066 6 OpcodeCondIn[1]
rlabel m2contact 14865 5194 14865 5194 6 n_12
rlabel m2contact 14817 4402 14817 4402 6 WdSel
rlabel m2contact 14745 5194 14745 5194 6 n_89
rlabel m2contact 14721 7114 14721 7114 6 StatusReg[3]
rlabel m2contact 14721 2650 14721 2650 6 StatusReg[3]
rlabel m2contact 14697 3898 14697 3898 6 OpcodeCondIn[5]
rlabel m2contact 14673 7114 14673 7114 6 StatusReg[3]
rlabel m2contact 14673 5434 14673 5434 6 n_20
rlabel m2contact 14625 7042 14625 7042 6 n_499
rlabel m2contact 14481 5194 14481 5194 6 n_89
rlabel m2contact 14409 2218 14409 2218 6 n_130
rlabel m2contact 14385 5890 14385 5890 6 stateSub[2]
rlabel m2contact 14289 2818 14289 2818 6 n_193
rlabel m2contact 14265 6058 14265 6058 6 n_383
rlabel m2contact 14265 4330 14265 4330 6 n_194
rlabel m2contact 14241 3154 14241 3154 6 n_57
rlabel m2contact 14193 4402 14193 4402 4 WdSel
rlabel m2contact 14145 3922 14145 3922 4 LrWe
rlabel m2contact 14145 2722 14145 2722 4 n_10
rlabel m2contact 14121 6850 14121 6850 4 n_261
rlabel m2contact 14097 4402 14097 4402 4 n_155
rlabel m2contact 14073 3922 14073 3922 4 LrWe
rlabel m2contact 14073 5218 14073 5218 4 n_171
rlabel m2contact 14049 4090 14049 4090 4 n_151
rlabel m2contact 14025 6202 14025 6202 4 n_317
rlabel m2contact 14001 5290 14001 5290 4 n_354
rlabel m2contact 13977 5914 13977 5914 4 n_215
rlabel m2contact 13977 5074 13977 5074 4 n_243
rlabel m2contact 13953 6634 13953 6634 4 n_209
rlabel m2contact 13929 4162 13929 4162 4 n_309
rlabel m2contact 13905 3802 13905 3802 4 stateSub[0]
rlabel m2contact 13905 3922 13905 3922 4 n_255
rlabel m2contact 13881 5338 13881 5338 4 OpcodeCondIn[4]
rlabel m2contact 13857 4330 13857 4330 4 n_194
rlabel m2contact 13833 4642 13833 4642 4 n_229
rlabel m2contact 13809 7114 13809 7114 4 n_357
rlabel m2contact 13809 3730 13809 3730 4 n_357
rlabel m2contact 13785 2290 13785 2290 4 n_190
rlabel m2contact 13785 2314 13785 2314 4 n_300
rlabel m2contact 13761 5914 13761 5914 4 n_215
rlabel m2contact 13737 3178 13737 3178 4 n_299
rlabel m2contact 13713 7018 13713 7018 4 CFlag
rlabel m2contact 13689 7114 13689 7114 4 n_357
rlabel m2contact 13689 6058 13689 6058 4 n_342
rlabel m2contact 13665 7042 13665 7042 4 n_126
rlabel m2contact 13665 3754 13665 3754 4 n_126
rlabel m2contact 13641 3994 13641 3994 4 n_205
rlabel m2contact 13617 2242 13617 2242 4 n_109
rlabel m2contact 13617 2290 13617 2290 4 n_328
rlabel m2contact 13593 3778 13593 3778 4 n_85
rlabel m2contact 13569 2242 13569 2242 4 n_137
rlabel m2contact 13545 1978 13545 1978 4 n_319
rlabel m2contact 13545 5218 13545 5218 4 n_95
rlabel m2contact 13521 7090 13521 7090 4 n_76
rlabel m2contact 13521 3130 13521 3130 4 n_48
rlabel m2contact 13497 4450 13497 4450 4 n_236
rlabel m2contact 13473 2002 13473 2002 4 n_294
rlabel m2contact 13473 3514 13473 3514 4 n_8
rlabel m2contact 13449 4450 13449 4450 4 n_238
rlabel m2contact 13449 4930 13449 4930 4 n_26
rlabel m2contact 13425 3802 13425 3802 4 stateSub[0]
rlabel m2contact 13401 3514 13401 3514 4 n_306
rlabel m2contact 13377 7066 13377 7066 4 n_44
rlabel m2contact 13377 4498 13377 4498 4 n_274
rlabel m2contact 13353 2578 13353 2578 4 n_284
rlabel m2contact 13353 5338 13353 5338 4 OpcodeCondIn[4]
rlabel m2contact 13329 7042 13329 7042 4 n_126
rlabel m2contact 13329 4306 13329 4306 4 n_282
rlabel m2contact 13281 5122 13281 5122 4 n_92
rlabel m2contact 13257 2026 13257 2026 4 n_104
rlabel m2contact 13233 5122 13233 5122 4 n_38
rlabel m2contact 13209 2842 13209 2842 4 n_289
rlabel m2contact 13161 2602 13161 2602 4 n_177
rlabel m2contact 13137 3610 13137 3610 4 state[1]
rlabel m2contact 13113 2050 13113 2050 4 n_105
rlabel m2contact 13113 2602 13113 2602 4 n_176
rlabel m2contact 13089 4858 13089 4858 4 n_123
rlabel m2contact 13065 3586 13065 3586 4 n_3
rlabel m2contact 13041 4858 13041 4858 4 n_91
rlabel m2contact 13041 3106 13041 3106 4 OpcodeCondIn[0]
rlabel m2contact 13017 4498 13017 4498 4 n_274
rlabel m2contact 13017 4066 13017 4066 4 OpcodeCondIn[1]
rlabel m2contact 12993 6994 12993 6994 4 n_31
rlabel m2contact 12969 3058 12969 3058 4 n_157
rlabel m2contact 12921 4642 12921 4642 4 n_229
rlabel m2contact 12897 4258 12897 4258 4 n_162
rlabel m2contact 12873 7018 12873 7018 4 CFlag
rlabel m2contact 12873 6994 12873 6994 4 n_345
rlabel m2contact 12873 3586 12873 3586 4 n_345
rlabel m2contact 12849 5770 12849 5770 4 n_198
rlabel m2contact 12825 6994 12825 6994 4 n_345
rlabel m2contact 12825 5002 12825 5002 4 OpcodeCondIn[7]
rlabel m2contact 12801 2242 12801 2242 4 n_137
rlabel m2contact 12801 5770 12801 5770 4 n_51
rlabel m2contact 12777 2362 12777 2362 4 n_313
rlabel m2contact 12729 2938 12729 2938 4 n_378
rlabel m2contact 12729 6130 12729 6130 4 n_79
rlabel m2contact 12705 4018 12705 4018 4 n_225
rlabel m2contact 12681 5074 12681 5074 4 n_243
rlabel m2contact 12657 6130 12657 6130 4 n_39
rlabel m2contact 12657 2626 12657 2626 4 n_39
rlabel m2contact 12633 6970 12633 6970 4 n_58
rlabel m2contact 12633 3298 12633 3298 4 n_145
rlabel m2contact 12609 3154 12609 3154 4 n_57
rlabel m2contact 12585 6946 12585 6946 4 n_40
rlabel m2contact 12585 5074 12585 5074 4 n_243
rlabel m2contact 12561 6130 12561 6130 4 n_39
rlabel m2contact 12561 5242 12561 5242 4 n_179
rlabel m2contact 12537 6442 12537 6442 4 n_240
rlabel m2contact 12537 2938 12537 2938 4 n_240
rlabel m2contact 12513 5722 12513 5722 4 n_68
rlabel m2contact 12489 2362 12489 2362 4 n_59
rlabel m2contact 12465 2242 12465 2242 4 n_27
rlabel m2contact 12441 2938 12441 2938 4 n_240
rlabel m2contact 12441 6130 12441 6130 4 n_19
rlabel m2contact 12369 4330 12369 4330 4 n_194
rlabel m2contact 12321 6226 12321 6226 4 n_138
rlabel m2contact 12297 6490 12297 6490 4 n_56
rlabel m2contact 12297 2938 12297 2938 4 n_56
rlabel m2contact 12273 5722 12273 5722 4 n_33
rlabel m2contact 12249 2458 12249 2458 4 n_115
rlabel m2contact 12225 5002 12225 5002 4 OpcodeCondIn[7]
rlabel m2contact 12201 2938 12201 2938 4 n_56
rlabel m2contact 12201 4642 12201 4642 4 n_229
rlabel m2contact 12177 6946 12177 6946 4 n_145
rlabel m2contact 12177 3298 12177 3298 4 n_145
rlabel m2contact 12153 6226 12153 6226 4 n_138
rlabel m2contact 12153 2938 12153 2938 4 n_265
rlabel m2contact 12129 5890 12129 5890 4 stateSub[2]
rlabel m2contact 12129 4258 12129 4258 4 n_162
rlabel m2contact 12105 6946 12105 6946 4 n_145
rlabel m2contact 12105 4666 12105 4666 4 n_273
rlabel m2contact 12081 6226 12081 6226 4 n_42
rlabel m2contact 12081 2074 12081 2074 4 n_42
rlabel m2contact 12057 6226 12057 6226 4 n_42
rlabel m2contact 12057 3418 12057 3418 4 n_118
rlabel m2contact 12033 5914 12033 5914 4 n_215
rlabel m2contact 12033 4642 12033 4642 4 n_229
rlabel m2contact 12009 5434 12009 5434 4 n_20
rlabel m2contact 12009 3754 12009 3754 4 n_126
rlabel m2contact 11961 6922 11961 6922 4 n_116
rlabel m2contact 11961 6226 11961 6226 4 AluOR[1]
rlabel m2contact 11937 4162 11937 4162 4 n_309
rlabel m2contact 11913 2458 11913 2458 4 n_115
rlabel m2contact 11865 4138 11865 4138 4 n_53
rlabel m2contact 11841 5722 11841 5722 4 n_33
rlabel m2contact 11817 3466 11817 3466 4 IntStatus
rlabel m2contact 11817 4090 11817 4090 4 n_151
rlabel m2contact 11769 5218 11769 5218 4 n_95
rlabel m2contact 11721 5218 11721 5218 4 n_37
rlabel m2contact 11697 6658 11697 6658 4 n_94
rlabel m2contact 11625 4138 11625 4138 4 n_222
rlabel m2contact 11601 3730 11601 3730 4 n_357
rlabel m2contact 11577 2386 11577 2386 4 n_381
rlabel m2contact 11553 2554 11553 2554 4 n_373
rlabel m2contact 11505 6274 11505 6274 4 n_186
rlabel m2contact 11457 5242 11457 5242 4 n_179
rlabel m2contact 11433 4474 11433 4474 4 n_84
rlabel m2contact 11385 6226 11385 6226 4 AluOR[1]
rlabel m2contact 11361 3706 11361 3706 4 n_359
rlabel m2contact 11337 3730 11337 3730 4 n_352
rlabel m2contact 11313 3034 11313 3034 4 n_346
rlabel m2contact 11289 3466 11289 3466 4 n_329
rlabel m2contact 11265 6226 11265 6226 4 n_108
rlabel m2contact 11241 2458 11241 2458 4 n_62
rlabel m2contact 11217 4090 11217 4090 4 n_151
rlabel m2contact 11169 6898 11169 6898 4 n_287
rlabel m2contact 11169 2266 11169 2266 4 n_96
rlabel m2contact 11145 2074 11145 2074 4 n_42
rlabel m2contact 11145 2266 11145 2266 4 n_96
rlabel m2contact 11121 2098 11121 2098 4 n_228
rlabel m2contact 11073 2098 11073 2098 4 nME
rlabel m2contact 11025 5242 11025 5242 4 n_179
rlabel m2contact 10977 2098 10977 2098 4 nME
rlabel m2contact 10977 4930 10977 4930 4 n_26
rlabel m2contact 10953 2434 10953 2434 4 n_184
rlabel m2contact 10953 3610 10953 3610 4 state[1]
rlabel m2contact 10905 2122 10905 2122 4 n_125
rlabel m2contact 10905 5938 10905 5938 4 n_227
rlabel m2contact 10857 6538 10857 6538 4 n_224
rlabel m2contact 10833 6874 10833 6874 4 n_200
rlabel m2contact 10833 3418 10833 3418 4 n_118
rlabel m2contact 10809 5938 10809 5938 4 n_129
rlabel m2contact 10785 4450 10785 4450 4 n_238
rlabel m2contact 10761 4594 10761 4594 4 n_237
rlabel m2contact 10737 4450 10737 4450 4 n_216
rlabel m2contact 10689 6850 10689 6850 4 n_261
rlabel m2contact 10665 2146 10665 2146 4 n_181
rlabel m2contact 10641 4234 10641 4234 4 n_211
rlabel m2contact 10617 4666 10617 4666 4 n_273
rlabel m2contact 10617 2146 10617 2146 4 n_273
rlabel m2contact 10593 5938 10593 5938 4 n_129
rlabel m2contact 10593 3058 10593 3058 4 n_157
rlabel m2contact 10569 2146 10569 2146 4 n_273
rlabel m2contact 10569 4426 10569 4426 4 state[0]
rlabel m2contact 10545 5938 10545 5938 4 n_73
rlabel m2contact 10521 3226 10521 3226 4 n_250
rlabel m2contact 10497 2170 10497 2170 4 n_344
rlabel m2contact 10473 5986 10473 5986 4 StatusReg[0]
rlabel m2contact 10473 3250 10473 3250 4 n_202
rlabel m2contact 10449 6058 10449 6058 4 n_342
rlabel m2contact 10449 3370 10449 3370 4 n_178
rlabel m2contact 10401 2194 10401 2194 4 n_293
rlabel m2contact 10377 6826 10377 6826 4 n_221
rlabel m2contact 10377 2602 10377 2602 4 n_176
rlabel m2contact 10353 2218 10353 2218 4 n_130
rlabel m2contact 10329 6802 10329 6802 4 n_93
rlabel m2contact 10329 4258 10329 4258 4 n_162
rlabel m2contact 10305 4282 10305 4282 4 n_128
rlabel m2contact 10257 4642 10257 4642 4 n_229
rlabel m2contact 10233 6178 10233 6178 4 n_297
rlabel m2contact 10233 5026 10233 5026 4 n_230
rlabel m2contact 10185 2242 10185 2242 4 n_27
rlabel m2contact 10185 4282 10185 4282 4 n_271
rlabel m2contact 10137 6778 10137 6778 4 n_197
rlabel m2contact 10137 5746 10137 5746 4 n_25
rlabel m2contact 10113 5074 10113 5074 4 n_243
rlabel m2contact 10113 4930 10113 4930 4 n_26
rlabel m2contact 10089 3946 10089 3946 4 n_196
rlabel m2contact 10065 4042 10065 4042 4 n_388
rlabel m2contact 10041 6682 10041 6682 4 n_304
rlabel m2contact 10017 4522 10017 4522 4 n_259
rlabel m2contact 9993 4042 9993 4042 4 n_214
rlabel m2contact 9921 6538 9921 6538 4 n_224
rlabel m2contact 9921 3946 9921 3946 4 n_224
rlabel m2contact 9897 3946 9897 3946 4 n_224
rlabel m2contact 9897 4546 9897 4546 4 n_102
rlabel m2contact 9873 6346 9873 6346 4 n_276
rlabel m2contact 9825 3946 9825 3946 4 AluWe
rlabel m2contact 9801 5818 9801 5818 4 n_72
rlabel m2contact 9801 2242 9801 2242 4 n_72
rlabel m2contact 9777 6754 9777 6754 4 RwSel[0]
rlabel m2contact 9777 6682 9777 6682 4 n_210
rlabel m2contact 9753 3586 9753 3586 4 n_345
rlabel m2contact 9753 4882 9753 4882 4 stateSub[1]
rlabel m2contact 9729 5842 9729 5842 4 n_263
rlabel m2contact 9705 2338 9705 2338 4 n_107
rlabel m2contact 9705 6442 9705 6442 4 n_240
rlabel m2contact 9681 5266 9681 5266 4 n_323
rlabel m2contact 9681 4498 9681 4498 4 n_274
rlabel m2contact 9657 5698 9657 5698 4 n_159
rlabel m2contact 9633 5146 9633 5146 4 n_34
rlabel m2contact 9609 3946 9609 3946 4 AluWe
rlabel m2contact 9609 4354 9609 4354 4 OpcodeCondIn[3]
rlabel m2contact 9585 3586 9585 3586 4 n_231
rlabel m2contact 9585 3802 9585 3802 4 stateSub[0]
rlabel m2contact 9561 2386 9561 2386 4 n_381
rlabel m2contact 9561 5722 9561 5722 4 n_33
rlabel m2contact 9537 2554 9537 2554 4 n_373
rlabel m2contact 9513 5746 9513 5746 4 n_25
rlabel m2contact 9489 4114 9489 4114 4 OpcodeCondIn[6]
rlabel m2contact 9465 2242 9465 2242 4 n_72
rlabel m2contact 9465 3898 9465 3898 4 OpcodeCondIn[5]
rlabel m2contact 9441 5338 9441 5338 4 OpcodeCondIn[4]
rlabel m2contact 9417 2266 9417 2266 4 n_96
rlabel m2contact 9417 3946 9417 3946 4 nOE
rlabel m2contact 9393 5410 9393 5410 4 n_246
rlabel m2contact 9369 2290 9369 2290 4 n_328
rlabel m2contact 9369 6346 9369 6346 4 n_330
rlabel m2contact 9345 6730 9345 6730 4 n_167
rlabel m2contact 9345 5266 9345 5266 4 n_310
rlabel m2contact 9321 6706 9321 6706 4 n_161
rlabel m2contact 9321 5842 9321 5842 4 n_296
rlabel m2contact 9297 5146 9297 5146 4 n_168
rlabel m2contact 9297 2290 9297 2290 4 n_168
rlabel m2contact 9273 5602 9273 5602 4 n_60
rlabel m2contact 9273 3658 9273 3658 4 n_367
rlabel m2contact 9249 2290 9249 2290 4 n_168
rlabel m2contact 9249 3826 9249 3826 4 n_14
rlabel m2contact 9225 2314 9225 2314 4 n_300
rlabel m2contact 9225 2362 9225 2362 4 n_59
rlabel m2contact 9201 5290 9201 5290 4 n_354
rlabel m2contact 9177 5266 9177 5266 4 n_310
rlabel m2contact 9177 3922 9177 3922 4 n_255
rlabel m2contact 9153 4162 9153 4162 4 n_309
rlabel m2contact 9129 5266 9129 5266 4 n_247
rlabel m2contact 9105 2602 9105 2602 4 n_176
rlabel m2contact 9081 4858 9081 4858 4 n_91
rlabel m2contact 9081 5410 9081 5410 4 n_246
rlabel m2contact 9057 2338 9057 2338 4 n_107
rlabel m2contact 9057 3610 9057 3610 4 state[1]
rlabel m2contact 9033 4546 9033 4546 4 n_102
rlabel m2contact 9009 3850 9009 3850 4 n_141
rlabel m2contact 8985 3274 8985 3274 4 n_174
rlabel m2contact 8985 4858 8985 4858 4 n_154
rlabel m2contact 8961 2362 8961 2362 4 n_59
rlabel m2contact 8961 3346 8961 3346 4 n_117
rlabel m2contact 8937 4738 8937 4738 4 n_83
rlabel m2contact 8913 4138 8913 4138 4 n_222
rlabel m2contact 8889 6322 8889 6322 4 n_203
rlabel m2contact 8889 5962 8889 5962 4 n_9
rlabel m2contact 8865 5290 8865 5290 4 n_149
rlabel m2contact 8865 4234 8865 4234 4 n_211
rlabel m2contact 8841 5602 8841 5602 4 n_86
rlabel m2contact 8841 3322 8841 3322 4 n_187
rlabel m2contact 8793 4738 8793 4738 4 n_170
rlabel m2contact 8769 3082 8769 3082 4 OpcodeCondIn[2]
rlabel m2contact 8745 5650 8745 5650 4 n_166
rlabel m2contact 8745 3082 8745 3082 4 OpcodeCondIn[2]
rlabel m2contact 8721 3322 8721 3322 4 n_187
rlabel m2contact 8673 6322 8673 6322 4 n_50
rlabel m2contact 8649 2458 8649 2458 4 n_62
rlabel m2contact 8649 3106 8649 3106 4 OpcodeCondIn[0]
rlabel m2contact 8625 4906 8625 4906 4 n_49
rlabel m2contact 8601 4498 8601 4498 4 n_274
rlabel m2contact 8577 4282 8577 4282 4 n_271
rlabel m2contact 8553 6658 8553 6658 4 n_94
rlabel m2contact 8529 2650 8529 2650 4 StatusReg[3]
rlabel m2contact 8529 5026 8529 5026 4 n_230
rlabel m2contact 8505 6058 8505 6058 4 n_342
rlabel m2contact 8481 6658 8481 6658 4 ImmSel
rlabel m2contact 8433 6562 8433 6562 4 n_156
rlabel m2contact 8409 2458 8409 2458 4 n_30
rlabel m2contact 8385 6562 8385 6562 4 n_97
rlabel m2contact 8337 6682 8337 6682 4 n_210
rlabel m2contact 8337 6658 8337 6658 4 ImmSel
rlabel m2contact 8313 5506 8313 5506 4 n_45
rlabel m2contact 8313 3850 8313 3850 4 n_121
rlabel m2contact 8289 6634 8289 6634 4 n_209
rlabel m2contact 8265 2386 8265 2386 4 n_381
rlabel m2contact 8241 2410 8241 2410 4 n_372
rlabel m2contact 8241 6610 8241 6610 4 n_165
rlabel m2contact 8217 6586 8217 6586 4 n_75
rlabel m2contact 8193 2770 8193 2770 4 n_6
rlabel m2contact 8193 4330 8193 4330 4 n_194
rlabel m2contact 8145 6562 8145 6562 4 n_97
rlabel m2contact 8145 3970 8145 3970 4 nWait
rlabel m2contact 8121 3610 8121 3610 4 state[1]
rlabel m2contact 8121 4114 8121 4114 4 OpcodeCondIn[6]
rlabel m2contact 8097 5698 8097 5698 4 n_159
rlabel m2contact 8073 2770 8073 2770 4 n_185
rlabel m2contact 8073 5434 8073 5434 4 n_20
rlabel m2contact 8049 6322 8049 6322 4 n_50
rlabel m2contact 8025 2434 8025 2434 4 n_184
rlabel m2contact 8025 2842 8025 2842 4 n_289
rlabel m2contact 8001 4018 8001 4018 4 n_225
rlabel m2contact 7977 2458 7977 2458 4 n_30
rlabel m2contact 7977 4546 7977 4546 4 n_102
rlabel m2contact 7953 5914 7953 5914 4 n_215
rlabel m2contact 7929 5722 7929 5722 4 n_33
rlabel m2contact 7929 6322 7929 6322 4 n_78
rlabel m2contact 7881 4162 7881 4162 4 n_309
rlabel m2contact 7857 2482 7857 2482 4 n_136
rlabel m2contact 7857 4546 7857 4546 4 n_102
rlabel m2contact 7809 2506 7809 2506 4 n_120
rlabel m2contact 7809 5722 7809 5722 4 n_226
rlabel m2contact 7785 2746 7785 2746 4 n_207
rlabel m2contact 7761 6538 7761 6538 4 n_224
rlabel m2contact 7761 2530 7761 2530 4 RwSel[1]
rlabel m2contact 7737 3010 7737 3010 4 n_253
rlabel m2contact 7737 4018 7737 4018 4 n_225
rlabel m2contact 7713 2554 7713 2554 4 n_373
rlabel m2contact 7689 6514 7689 6514 4 n_124
rlabel m2contact 7665 6490 7665 6490 4 n_56
rlabel m2contact 7665 3034 7665 3034 4 n_346
rlabel m2contact 7641 3418 7641 3418 4 n_118
rlabel m2contact 7593 4978 7593 4978 4 n_241
rlabel m2contact 7593 3418 7593 3418 4 n_135
rlabel m2contact 7569 6466 7569 6466 4 n_192
rlabel m2contact 7545 4978 7545 4978 4 n_199
rlabel m2contact 7521 6442 7521 6442 4 n_240
rlabel m2contact 7521 6418 7521 6418 4 n_81
rlabel m2contact 7497 3082 7497 3082 4 OpcodeCondIn[2]
rlabel m2contact 7473 6394 7473 6394 4 n_286
rlabel m2contact 7449 4018 7449 4018 4 n_225
rlabel m2contact 7425 6370 7425 6370 4 n_277
rlabel m2contact 7401 5770 7401 5770 4 n_51
rlabel m2contact 7377 6346 7377 6346 4 n_330
rlabel m2contact 7377 5866 7377 5866 4 n_74
rlabel m2contact 7329 6322 7329 6322 4 n_78
rlabel m2contact 7305 6298 7305 6298 4 n_311
rlabel m2contact 7305 5506 7305 5506 4 n_45
rlabel m2contact 7281 4426 7281 4426 4 state[0]
rlabel m2contact 7257 5506 7257 5506 4 n_283
rlabel m2contact 7233 4690 7233 4690 4 n_267
rlabel m2contact 7209 2578 7209 2578 4 n_284
rlabel m2contact 7185 2746 7185 2746 4 n_207
rlabel m2contact 7161 5650 7161 5650 4 n_166
rlabel m2contact 7161 3754 7161 3754 4 n_126
rlabel m2contact 7137 6058 7137 6058 4 n_342
rlabel m2contact 7137 2578 7137 2578 4 n_342
rlabel m2contact 7113 2578 7113 2578 4 n_342
rlabel m2contact 7113 4882 7113 4882 4 stateSub[1]
rlabel m2contact 7089 6274 7089 6274 4 n_186
rlabel m2contact 7089 2602 7089 2602 4 n_176
rlabel m2contact 7065 6250 7065 6250 4 n_239
rlabel m2contact 7041 6106 7041 6106 4 n_18
rlabel m2contact 7041 3298 7041 3298 4 n_145
rlabel m2contact 7017 6226 7017 6226 4 n_108
rlabel m2contact 6993 3082 6993 3082 4 OpcodeCondIn[2]
rlabel m2contact 6969 4114 6969 4114 4 OpcodeCondIn[6]
rlabel m2contact 6921 6202 6921 6202 4 n_317
rlabel m2contact 6921 3226 6921 3226 4 n_250
rlabel m2contact 6897 5698 6897 5698 4 n_159
rlabel m2contact 6873 6178 6873 6178 4 n_297
rlabel m2contact 6873 6154 6873 6154 4 n_4
rlabel m2contact 6849 5002 6849 5002 4 OpcodeCondIn[7]
rlabel m2contact 6825 6130 6825 6130 4 n_19
rlabel m2contact 6825 3802 6825 3802 4 stateSub[0]
rlabel m2contact 6777 2626 6777 2626 4 n_39
rlabel m2contact 6777 6106 6777 6106 4 n_18
rlabel m2contact 6753 6010 6753 6010 4 n_23
rlabel m2contact 6729 2650 6729 2650 4 StatusReg[3]
rlabel m2contact 6705 6082 6705 6082 4 n_340
rlabel m2contact 6705 6010 6705 6010 4 OpcodeCondIn[0]
rlabel m2contact 6705 3106 6705 3106 4 OpcodeCondIn[0]
rlabel m2contact 6681 2674 6681 2674 4 n_99
rlabel m2contact 6681 2914 6681 2914 4 StatusReg[2]
rlabel m2contact 6657 6058 6657 6058 4 n_342
rlabel m2contact 6657 4114 6657 4114 4 OpcodeCondIn[6]
rlabel m2contact 6633 3754 6633 3754 4 n_126
rlabel m2contact 6609 6034 6609 6034 4 n_11
rlabel m2contact 6609 5482 6609 5482 4 n_71
rlabel m2contact 6585 6010 6585 6010 4 OpcodeCondIn[0]
rlabel m2contact 6585 4354 6585 4354 4 OpcodeCondIn[3]
rlabel m2contact 6561 5986 6561 5986 4 StatusReg[0]
rlabel m2contact 6537 2698 6537 2698 4 n_332
rlabel m2contact 6537 4066 6537 4066 4 OpcodeCondIn[1]
rlabel m2contact 6513 5074 6513 5074 4 n_243
rlabel m2contact 6489 2986 6489 2986 4 n_131
rlabel m2contact 6465 2722 6465 2722 4 n_10
rlabel m2contact 6417 5962 6417 5962 4 n_9
rlabel m2contact 6393 3082 6393 3082 4 OpcodeCondIn[2]
rlabel m2contact 6369 5938 6369 5938 4 n_73
rlabel m2contact 6345 5914 6345 5914 4 n_215
rlabel m2contact 6345 5890 6345 5890 4 stateSub[2]
rlabel m2contact 6321 5890 6321 5890 4 stateSub[2]
rlabel m2contact 6321 3106 6321 3106 4 OpcodeCondIn[0]
rlabel m2contact 6297 5866 6297 5866 4 n_74
rlabel m2contact 6273 5818 6273 5818 4 n_72
rlabel m2contact 6225 5842 6225 5842 4 n_296
rlabel m2contact 6225 2746 6225 2746 4 n_207
rlabel m2contact 6225 5818 6225 5818 4 n_299
rlabel m2contact 6225 3178 6225 3178 4 n_299
rlabel m2contact 6201 3202 6201 3202 4 n_110
rlabel m2contact 6201 5194 6201 5194 4 n_89
rlabel m2contact 6177 5818 6177 5818 4 n_299
rlabel m2contact 6177 4162 6177 4162 4 n_309
rlabel m2contact 6129 5794 6129 5794 4 n_266
rlabel m2contact 6129 3202 6129 3202 4 n_98
rlabel m2contact 6105 4114 6105 4114 4 OpcodeCondIn[6]
rlabel m2contact 6081 2770 6081 2770 4 n_185
rlabel m2contact 6033 2794 6033 2794 4 n_501
rlabel m2contact 6009 2818 6009 2818 4 n_193
rlabel m2contact 6009 5338 6009 5338 4 OpcodeCondIn[4]
rlabel m2contact 5985 3898 5985 3898 4 OpcodeCondIn[5]
rlabel m2contact 5961 4666 5961 4666 4 n_273
rlabel m2contact 5937 4642 5937 4642 4 n_229
rlabel m2contact 5913 3322 5913 3322 4 n_187
rlabel m2contact 5889 4666 5889 4666 4 n_273
rlabel m2contact 5865 5770 5865 5770 4 n_51
rlabel m2contact 5817 5746 5817 5746 4 n_25
rlabel m2contact 5817 2842 5817 2842 4 n_289
rlabel m2contact 5793 5722 5793 5722 4 n_226
rlabel m2contact 5769 5626 5769 5626 4 n_160
rlabel m2contact 5745 5698 5745 5698 4 n_159
rlabel m2contact 5745 5674 5745 5674 4 n_275
rlabel m2contact 5721 2866 5721 2866 4 n_232
rlabel m2contact 5721 5650 5721 5650 4 n_166
rlabel m2contact 5721 5626 5721 5626 4 n_174
rlabel m2contact 5721 3274 5721 3274 4 n_174
rlabel m2contact 5697 5626 5697 5626 4 n_174
rlabel m2contact 5697 4666 5697 4666 4 n_273
rlabel m2contact 5673 4498 5673 4498 4 n_274
rlabel m2contact 5649 5602 5649 5602 4 n_86
rlabel m2contact 5625 4498 5625 4498 4 n_274
rlabel m2contact 5601 4210 5601 4210 4 n_204
rlabel m2contact 5553 2890 5553 2890 4 n_363
rlabel m2contact 5529 2914 5529 2914 4 StatusReg[2]
rlabel m2contact 5505 3658 5505 3658 4 n_367
rlabel m2contact 5457 3658 5457 3658 4 n_61
rlabel m2contact 5433 3802 5433 3802 4 stateSub[0]
rlabel m2contact 5409 4378 5409 4378 4 n_28
rlabel m2contact 5337 4666 5337 4666 4 n_273
rlabel m2contact 5289 4378 5289 4378 4 n_189
rlabel m2contact 5241 5578 5241 5578 4 n_315
rlabel m2contact 5217 5530 5217 5530 4 n_314
rlabel m2contact 5193 2938 5193 2938 4 n_265
rlabel m2contact 5169 5554 5169 5554 4 n_245
rlabel m2contact 5121 2962 5121 2962 4 n_387
rlabel m2contact 5121 3730 5121 3730 4 n_352
rlabel m2contact 5073 5530 5073 5530 4 n_314
rlabel m2contact 5049 5506 5049 5506 4 n_283
rlabel m2contact 5001 5482 5001 5482 4 n_71
rlabel m2contact 5001 5458 5001 5458 4 n_147
rlabel m2contact 4953 3898 4953 3898 4 OpcodeCondIn[5]
rlabel m2contact 4929 5434 4929 5434 4 n_20
rlabel m2contact 4881 5266 4881 5266 4 n_247
rlabel m2contact 4857 5410 4857 5410 4 n_246
rlabel m2contact 4857 4882 4857 4882 4 stateSub[1]
rlabel m2contact 4833 2986 4833 2986 4 n_131
rlabel m2contact 4833 5266 4833 5266 4 n_201
rlabel m2contact 4785 5386 4785 5386 4 n_325
rlabel m2contact 4785 5362 4785 5362 4 n_254
rlabel m2contact 4761 3010 4761 3010 4 n_253
rlabel m2contact 4737 3034 4737 3034 4 n_346
rlabel m2contact 4737 5338 4737 5338 4 OpcodeCondIn[4]
rlabel m2contact 4713 5314 4713 5314 4 n_281
rlabel m2contact 4689 5290 4689 5290 4 n_149
rlabel m2contact 4665 3058 4665 3058 4 n_157
rlabel m2contact 4665 5266 4665 5266 4 n_201
rlabel m2contact 4641 5242 4641 5242 4 n_179
rlabel m2contact 4641 4162 4641 4162 4 n_309
rlabel m2contact 4617 3994 4617 3994 4 n_205
rlabel m2contact 4569 3082 4569 3082 4 OpcodeCondIn[2]
rlabel m2contact 4569 5218 4569 5218 4 n_37
rlabel m2contact 4545 3106 4545 3106 4 OpcodeCondIn[0]
rlabel m2contact 4521 4642 4521 4642 4 n_229
rlabel m2contact 4497 5194 4497 5194 4 n_89
rlabel m2contact 4449 3130 4449 3130 4 n_48
rlabel m2contact 4425 3154 4425 3154 4 n_57
rlabel m2contact 4425 3610 4425 3610 4 state[1]
rlabel m2contact 4401 5170 4401 5170 4 n_47
rlabel m2contact 4353 5146 4353 5146 4 n_168
rlabel m2contact 4353 3178 4353 3178 4 n_299
rlabel m2contact 4329 3202 4329 3202 4 n_98
rlabel m2contact 4305 4330 4305 4330 4 n_194
rlabel m2contact 4257 5122 4257 5122 4 n_38
rlabel m2contact 4257 5098 4257 5098 4 n_235
rlabel m2contact 4233 4378 4233 4378 4 n_189
rlabel m2contact 4209 4090 4209 4090 4 n_151
rlabel m2contact 4185 5074 4185 5074 4 n_243
rlabel m2contact 4113 3226 4113 3226 4 n_250
rlabel m2contact 4113 5050 4113 5050 4 n_22
rlabel m2contact 4089 5002 4089 5002 4 OpcodeCondIn[7]
rlabel m2contact 4065 3250 4065 3250 4 n_202
rlabel m2contact 4041 4426 4041 4426 4 state[0]
rlabel m2contact 4017 3274 4017 3274 4 n_174
rlabel m2contact 4017 4090 4017 4090 4 n_151
rlabel m2contact 3993 3298 3993 3298 4 n_145
rlabel m2contact 3945 5026 3945 5026 4 n_230
rlabel m2contact 3921 3322 3921 3322 4 n_187
rlabel m2contact 3897 5002 3897 5002 4 OpcodeCondIn[7]
rlabel m2contact 3873 3346 3873 3346 4 n_117
rlabel m2contact 3873 4330 3873 4330 4 n_194
rlabel m2contact 3825 4978 3825 4978 4 n_199
rlabel m2contact 3801 4954 3801 4954 4 n_144
rlabel m2contact 3801 3370 3801 3370 4 n_178
rlabel m2contact 3777 4426 3777 4426 4 state[0]
rlabel m2contact 3753 3394 3753 3394 4 n_111
rlabel m2contact 3729 3418 3729 3418 4 n_135
rlabel m2contact 3705 3442 3705 3442 4 PcWe
rlabel m2contact 3705 4162 3705 4162 4 n_309
rlabel m2contact 3681 3538 3681 3538 4 n_134
rlabel m2contact 3633 3466 3633 3466 4 n_329
rlabel m2contact 3609 3490 3609 3490 4 n_169
rlabel m2contact 3609 3706 3609 3706 4 n_359
rlabel m2contact 3585 3514 3585 3514 4 n_306
rlabel m2contact 3561 3898 3561 3898 4 OpcodeCondIn[5]
rlabel m2contact 3537 4522 3537 4522 4 n_259
rlabel m2contact 3513 4930 3513 4930 4 n_26
rlabel m2contact 3489 4090 3489 4090 4 n_151
rlabel m2contact 3465 3538 3465 3538 4 n_134
rlabel m2contact 3441 4906 3441 4906 4 n_49
rlabel m2contact 3417 3562 3417 3562 4 n_80
rlabel m2contact 3393 4090 3393 4090 4 n_151
rlabel m2contact 3369 4882 3369 4882 4 stateSub[1]
rlabel m2contact 3321 3586 3321 3586 4 n_231
rlabel m2contact 3297 4858 3297 4858 4 n_154
rlabel m2contact 3273 3610 3273 3610 4 state[1]
rlabel m2contact 3273 4234 3273 4234 4 n_211
rlabel m2contact 3249 3802 3249 3802 4 stateSub[0]
rlabel m2contact 3225 4162 3225 4162 4 n_309
rlabel m2contact 3225 4018 3225 4018 4 n_225
rlabel m2contact 3153 4834 3153 4834 4 n_234
rlabel m2contact 3105 4810 3105 4810 4 n_219
rlabel m2contact 3057 4786 3057 4786 4 n_88
rlabel m2contact 3033 4762 3033 4762 4 n_87
rlabel m2contact 3009 4234 3009 4234 4 n_211
rlabel m2contact 2937 4738 2937 4738 4 n_170
rlabel m2contact 2913 4714 2913 4714 4 n_334
rlabel m2contact 2865 3634 2865 3634 4 n_268
rlabel m2contact 2841 4690 2841 4690 4 n_267
rlabel m2contact 2817 4666 2817 4666 4 n_273
rlabel m2contact 2745 4642 2745 4642 4 n_229
rlabel m2contact 2697 3658 2697 3658 4 n_61
rlabel m2contact 2697 4114 2697 4114 4 OpcodeCondIn[6]
rlabel m2contact 2673 4618 2673 4618 4 n_67
rlabel m2contact 2649 3682 2649 3682 4 n_322
rlabel m2contact 2625 4594 2625 4594 4 n_237
rlabel m2contact 2601 4570 2601 4570 4 n_280
rlabel m2contact 2601 3706 2601 3706 4 n_359
rlabel m2contact 2577 3730 2577 3730 4 n_352
rlabel m2contact 2529 4546 2529 4546 4 n_102
rlabel m2contact 2505 3754 2505 3754 4 n_126
rlabel m2contact 2481 4522 2481 4522 4 n_259
rlabel m2contact 2433 3778 2433 3778 4 n_85
rlabel m2contact 2409 4498 2409 4498 4 n_274
rlabel m2contact 2385 4474 2385 4474 4 n_84
rlabel m2contact 2337 4450 2337 4450 4 n_216
rlabel m2contact 2313 4426 2313 4426 4 state[0]
rlabel m2contact 2289 4402 2289 4402 4 n_155
rlabel m2contact 2241 4378 2241 4378 4 n_189
rlabel m2contact 2217 3802 2217 3802 4 stateSub[0]
rlabel m2contact 2217 4354 2217 4354 4 OpcodeCondIn[3]
rlabel m2contact 2193 4330 2193 4330 4 n_194
rlabel m2contact 2169 3826 2169 3826 4 n_14
rlabel m2contact 2097 4306 2097 4306 4 n_282
rlabel m2contact 2073 4282 2073 4282 4 n_271
rlabel m2contact 2025 3850 2025 3850 4 n_121
rlabel m2contact 2001 4258 2001 4258 4 n_162
rlabel m2contact 1977 4234 1977 4234 4 n_211
rlabel m2contact 1953 4210 1953 4210 4 n_204
rlabel m2contact 1905 4186 1905 4186 4 n_223
rlabel m2contact 1857 4162 1857 4162 4 n_309
rlabel m2contact 1833 4138 1833 4138 4 n_222
rlabel m2contact 1785 3874 1785 3874 4 n_17
rlabel m2contact 1761 4114 1761 4114 4 OpcodeCondIn[6]
rlabel m2contact 1737 4090 1737 4090 4 n_151
rlabel m2contact 1713 4066 1713 4066 4 OpcodeCondIn[1]
rlabel m2contact 1665 4042 1665 4042 4 n_214
rlabel m2contact 1641 4018 1641 4018 4 n_225
rlabel m2contact 1641 3898 1641 3898 4 OpcodeCondIn[5]
rlabel m2contact 1617 3922 1617 3922 4 n_255
rlabel m2contact 1617 3994 1617 3994 4 n_205
rlabel m2contact 26961 353 26961 353 8 ENB
rlabel m2contact 26961 17 26961 17 8 ENB
rlabel m2contact 26937 41 26937 41 8 AluOR[1]
rlabel m2contact 26937 17 26937 17 8 AluOR[1]
rlabel m2contact 26937 569 26937 569 8 n_350
rlabel m2contact 26889 761 26889 761 8 n_175
rlabel m2contact 26697 641 26697 641 8 n_218
rlabel m2contact 26649 233 26649 233 8 n_122
rlabel m2contact 26625 209 26625 209 8 n_127
rlabel m2contact 26601 257 26601 257 8 n_114
rlabel m2contact 26457 617 26457 617 8 n_324
rlabel m2contact 24609 737 24609 737 8 n_264
rlabel m2contact 24489 1049 24489 1049 6 n_113
rlabel m2contact 24273 401 24273 401 8 n_64
rlabel m2contact 24249 593 24249 593 8 n_63
rlabel m2contact 24129 833 24129 833 6 n_258
rlabel m2contact 24081 41 24081 41 8 n_36
rlabel m2contact 24009 665 24009 665 8 n_15
rlabel m2contact 23961 1097 23961 1097 6 n_244
rlabel m2contact 23913 929 23913 929 6 n_164
rlabel m2contact 23745 1025 23745 1025 6 n_376
rlabel m2contact 23721 449 23721 449 8 n_132
rlabel m2contact 23697 689 23697 689 8 n_341
rlabel m2contact 23649 809 23649 809 6 n_133
rlabel m2contact 23433 1049 23433 1049 6 n_113
rlabel m2contact 23385 1145 23385 1145 6 n_66
rlabel m2contact 23193 569 23193 569 8 n_350
rlabel m2contact 22929 1073 22929 1073 6 n_35
rlabel m2contact 22785 785 22785 785 8 n_173
rlabel m2contact 22713 161 22713 161 8 SysBus[0]
rlabel m2contact 22569 809 22569 809 6 n_133
rlabel m2contact 22473 761 22473 761 8 n_175
rlabel m2contact 22209 713 22209 713 8 RegWe
rlabel m2contact 22113 329 22113 329 8 n_384
rlabel m2contact 21633 809 21633 809 6 n_188
rlabel m2contact 21129 953 21129 953 6 n_29
rlabel m2contact 21009 305 21009 305 8 n_380
rlabel m2contact 20985 521 20985 521 8 SysBus[3]
rlabel m2contact 20745 137 20745 137 8 n_292
rlabel m2contact 20697 761 20697 761 8 n_308
rlabel metal2 20643 713 20643 713 8 SysBus[2]
rlabel m2contact 20625 713 20625 713 8 SysBus[2]
rlabel m2contact 20553 473 20553 473 8 n_101
rlabel m2contact 20505 713 20505 713 8 n_41
rlabel m2contact 20433 425 20433 425 8 n_7
rlabel m2contact 20409 593 20409 593 8 n_63
rlabel m2contact 20385 401 20385 401 8 n_64
rlabel m2contact 20217 761 20217 761 8 n_308
rlabel m2contact 20169 737 20169 737 8 n_264
rlabel m2contact 20097 497 20097 497 8 n_32
rlabel m2contact 20049 593 20049 593 8 n_63
rlabel m2contact 19857 113 19857 113 8 nWE
rlabel m2contact 19761 545 19761 545 8 n_290
rlabel m2contact 19425 761 19425 761 8 n_143
rlabel m2contact 19281 905 19281 905 6 n_112
rlabel m2contact 18849 1121 18849 1121 6 IRQ1
rlabel m2contact 18441 89 18441 89 8 n_0
rlabel m2contact 18201 881 18201 881 6 n_368
rlabel m2contact 18105 1001 18105 1001 6 n_206
rlabel m2contact 18009 713 18009 713 8 n_41
rlabel m2contact 17913 689 17913 689 8 n_341
rlabel m2contact 17745 641 17745 641 8 n_218
rlabel m2contact 17697 713 17697 713 8 n_182
rlabel m2contact 17505 641 17505 641 8 n_242
rlabel m2contact 17121 977 17121 977 6 n_139
rlabel m2contact 17073 377 17073 377 8 n_90
rlabel m2contact 17001 281 17001 281 8 n_119
rlabel m2contact 16857 689 16857 689 8 n_248
rlabel m2contact 16809 185 16809 185 8 n_339
rlabel m2contact 16617 857 16617 857 6 n_100
rlabel m2contact 16449 737 16449 737 8 n_82
rlabel m2contact 16425 1145 16425 1145 6 n_66
rlabel m2contact 15873 1121 15873 1121 6 IRQ1
rlabel m2contact 15753 737 15753 737 8 n_82
rlabel m2contact 15705 737 15705 737 8 n_46
rlabel m2contact 15633 353 15633 353 8 ENB
rlabel m2contact 15561 353 15561 353 8 n_260
rlabel m2contact 15513 593 15513 593 8 n_63
rlabel m2contact 15321 353 15321 353 8 n_260
rlabel m2contact 15177 353 15177 353 8 n_298
rlabel m2contact 15153 569 15153 569 8 n_350
rlabel m2contact 15081 569 15081 569 8 n_213
rlabel m2contact 14937 761 14937 761 8 n_143
rlabel m2contact 14841 257 14841 257 8 n_114
rlabel m2contact 14793 1049 14793 1049 6 n_113
rlabel m2contact 14625 257 14625 257 8 n_301
rlabel m2contact 14601 1049 14601 1049 6 n_106
rlabel m2contact 14577 1097 14577 1097 6 n_244
rlabel m2contact 14529 377 14529 377 8 n_90
rlabel m2contact 14457 953 14457 953 6 n_29
rlabel m2contact 14361 857 14361 857 6 n_100
rlabel m2contact 14313 377 14313 377 8 n_195
rlabel m2contact 14049 713 14049 713 2 n_182
rlabel m2contact 13857 953 13857 953 4 n_191
rlabel m2contact 13809 713 13809 713 2 n_54
rlabel m2contact 13737 857 13737 857 4 n_343
rlabel m2contact 13209 1073 13209 1073 4 n_35
rlabel m2contact 13161 1049 13161 1049 4 n_106
rlabel m2contact 12681 1025 12681 1025 4 n_376
rlabel m2contact 12393 641 12393 641 2 n_242
rlabel m2contact 12345 641 12345 641 2 n_208
rlabel m2contact 12321 1001 12321 1001 4 n_206
rlabel m2contact 11961 17 11961 17 2 AluOR[1]
rlabel m2contact 11241 617 11241 617 2 n_324
rlabel m2contact 11193 617 11193 617 2 n_43
rlabel m2contact 11097 137 11097 137 2 n_292
rlabel m2contact 11049 977 11049 977 4 n_139
rlabel m2contact 11025 137 11025 137 2 n_256
rlabel m2contact 10929 953 10929 953 4 n_191
rlabel m2contact 10857 929 10857 929 4 n_164
rlabel m2contact 10761 353 10761 353 2 n_298
rlabel m2contact 10713 905 10713 905 4 n_112
rlabel m2contact 10689 353 10689 353 2 n_269
rlabel m2contact 10641 353 10641 353 2 n_269
rlabel m2contact 10281 329 10281 329 2 n_384
rlabel m2contact 10041 353 10041 353 2 n_251
rlabel m2contact 10017 881 10017 881 4 n_368
rlabel m2contact 9993 857 9993 857 4 n_343
rlabel m2contact 9945 833 9945 833 4 n_258
rlabel m2contact 9873 569 9873 569 2 n_213
rlabel m2contact 9825 569 9825 569 2 n_365
rlabel m2contact 9513 809 9513 809 4 n_188
rlabel m2contact 9129 785 9129 785 2 n_173
rlabel m2contact 8793 761 8793 761 2 n_143
rlabel m2contact 8721 593 8721 593 2 n_63
rlabel m2contact 8553 185 8553 185 2 n_339
rlabel m2contact 8433 185 8433 185 2 n_69
rlabel m2contact 8385 41 8385 41 2 n_36
rlabel m2contact 8289 569 8289 569 2 n_365
rlabel m2contact 8073 41 8073 41 2 SysBus[1]
rlabel m2contact 8037 161 8037 161 2 SysBus[0]
rlabel m2contact 7689 569 7689 569 2 n_270
rlabel m2contact 7617 161 7617 161 2 n_272
rlabel m2contact 7473 497 7473 497 2 n_32
rlabel m2contact 7425 497 7425 497 2 n_52
rlabel m2contact 7329 737 7329 737 2 n_46
rlabel m2contact 7233 713 7233 713 2 n_54
rlabel m2contact 6969 689 6969 689 2 n_248
rlabel m2contact 6945 521 6945 521 2 SysBus[3]
rlabel m2contact 6753 521 6753 521 2 n_500
rlabel m2contact 6417 665 6417 665 2 n_15
rlabel m2contact 6249 641 6249 641 2 n_208
rlabel m2contact 6105 617 6105 617 2 n_43
rlabel m2contact 6081 497 6081 497 2 n_52
rlabel m2contact 6033 497 6033 497 2 n_55
rlabel m2contact 5985 593 5985 593 2 n_63
rlabel m2contact 5937 569 5937 569 2 n_270
rlabel m2contact 5841 545 5841 545 2 n_290
rlabel m2contact 5481 521 5481 521 2 n_500
rlabel m2contact 4953 497 4953 497 2 n_55
rlabel m2contact 4929 473 4929 473 2 n_101
rlabel m2contact 4881 449 4881 449 2 n_132
rlabel m2contact 4593 425 4593 425 2 n_7
rlabel m2contact 4473 401 4473 401 2 n_64
rlabel m2contact 4305 329 4305 329 2 n_384
rlabel m2contact 4209 377 4209 377 2 n_195
rlabel m2contact 4161 353 4161 353 2 n_251
rlabel m2contact 4137 41 4137 41 2 SysBus[1]
rlabel m2contact 3681 329 3681 329 2 n_384
rlabel m2contact 3657 305 3657 305 2 n_380
rlabel m2contact 3537 281 3537 281 2 n_119
rlabel m2contact 2865 257 2865 257 2 n_301
rlabel m2contact 2745 233 2745 233 2 n_122
rlabel m2contact 2625 65 2625 65 2 AluOR[0]
rlabel m2contact 2529 209 2529 209 2 n_127
rlabel m2contact 2481 185 2481 185 2 n_69
rlabel m2contact 2409 89 2409 89 2 n_0
rlabel m2contact 2361 89 2361 89 2 nIRQ
rlabel m2contact 1809 161 1809 161 2 n_272
rlabel m2contact 1689 137 1689 137 2 n_256
rlabel metal2 27303 8300 27315 8300 6 StatusRegEn
rlabel metal2 25623 8300 25635 8300 6 StatusReg[3]
rlabel metal2 24771 8300 24783 8300 6 StatusReg[2]
rlabel metal2 23919 8300 23931 8300 6 StatusReg[1]
rlabel metal2 23067 8300 23079 8300 6 StatusReg[0]
rlabel metal2 22215 8300 22227 8300 6 AluEn
rlabel metal2 21363 8300 21375 8300 6 AluWe
rlabel metal2 20511 8300 20523 8300 6 Op2Sel[1]
rlabel metal2 20223 8300 20235 8300 6 Op2Sel[0]
rlabel metal2 18807 8300 18819 8300 6 Op1Sel
rlabel metal2 18783 8300 18795 8300 6 PcEn
rlabel metal2 17103 8300 17115 8300 6 WdSel
rlabel metal2 16887 8300 16899 8300 6 PcWe
rlabel metal2 15951 8300 15963 8300 6 PcSel[2]
rlabel metal2 15375 8300 15387 8300 6 PcSel[1]
rlabel metal2 14523 8300 14535 8300 6 PcSel[0]
rlabel metal2 12831 8300 12843 8300 4 LrEn
rlabel metal2 12795 8300 12807 8300 4 LrWe
rlabel metal2 11931 8300 11943 8300 4 LrSel
rlabel metal2 10239 8300 10251 8300 4 ImmSel
rlabel metal2 9951 8300 9963 8300 4 IrWe
rlabel metal2 9339 8300 9351 8300 4 MemEn
rlabel metal2 7647 8300 7659 8300 4 OpcodeCondIn[7]
rlabel metal2 6975 8300 6987 8300 4 OpcodeCondIn[6]
rlabel metal2 5991 8300 6003 8300 4 OpcodeCondIn[5]
rlabel metal2 5055 8300 5067 8300 4 OpcodeCondIn[4]
rlabel metal2 4191 8300 4203 8300 4 OpcodeCondIn[3]
rlabel metal2 4155 8300 4167 8300 4 OpcodeCondIn[2]
rlabel metal2 2463 8300 2475 8300 4 OpcodeCondIn[1]
rlabel metal2 2427 8300 2439 8300 4 OpcodeCondIn[0]
rlabel metal2 20979 0 20991 0 8 SysBus[3]
rlabel metal2 20631 0 20643 0 8 SysBus[2]
rlabel metal2 8067 0 8079 0 2 SysBus[1]
rlabel metal2 8031 0 8043 0 2 SysBus[0]
rlabel metal2 27937 707 27937 719 8 RegWe
rlabel metal2 27937 59 27937 71 8 AluOR[0]
rlabel metal2 27937 35 27937 47 8 AluOR[1]
rlabel metal2 27937 11 27937 23 8 ENB
rlabel metal2 27937 4564 27937 4576 6 Rs1Sel[0]
rlabel metal2 27937 3844 27937 3856 6 Rs1Sel[1]
rlabel metal2 27937 1996 27937 2008 6 RwSel[0]
rlabel metal2 27937 1972 27937 1984 6 RwSel[1]
rlabel metal2 27937 8037 27937 8049 6 CFlag
rlabel metal2 27937 8013 27937 8025 6 Flags[3]
rlabel metal2 27937 7989 27937 8001 6 Flags[2]
rlabel metal2 27937 7965 27937 7977 6 Flags[1]
rlabel metal2 27937 7941 27937 7953 6 Flags[0]
rlabel metal2 0 107 0 119 2 nWE
rlabel metal2 0 83 0 95 2 nIRQ
rlabel metal2 0 3964 0 3976 4 nWait
rlabel metal2 0 3940 0 3952 4 nOE
rlabel metal2 0 8061 0 8073 4 ALE
rlabel metal2 0 8037 0 8049 4 nME
rlabel metal2 27555 0 27755 0 1 GND!
rlabel space 123 0 324 0 1 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 123 8300 323 8300 5 Vdd!
rlabel metal2 339 8300 351 8300 5 SDO
rlabel metal2 363 8300 375 8300 5 Test
rlabel metal2 387 8300 399 8300 5 Clock
rlabel metal2 411 8300 423 8300 5 nReset
rlabel metal2 27555 8300 27756 8300 5 GND!
<< end >>
