magic
tech c035u
timestamp 1394475556
<< metal1 >>
rect 805 892 935 902
rect 757 870 887 880
rect 0 50 599 60
rect 613 50 743 60
rect 0 28 23 38
rect 37 28 1008 38
rect 973 6 1008 16
<< m2contact >>
rect 791 890 805 904
rect 935 890 949 904
rect 743 868 757 882
rect 887 868 901 882
rect 599 48 613 62
rect 743 48 757 62
rect 23 26 37 40
rect 959 4 973 18
<< metal2 >>
rect 72 865 84 1042
rect 744 882 756 1042
rect 792 904 804 1042
rect 744 865 756 868
rect 792 865 804 890
rect 864 865 876 1042
rect 888 865 900 868
rect 936 865 948 890
rect 24 40 36 66
rect 72 0 84 66
rect 600 62 612 66
rect 744 62 756 66
rect 792 0 804 66
rect 864 0 876 66
rect 960 18 972 66
use scanreg  scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 66
box 0 0 720 799
use rowcrosser  rowcrosser_2
timestamp 1386086759
transform 1 0 720 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_3
timestamp 1386086759
transform 1 0 768 0 1 66
box 0 0 48 799
use mux2  mux2_1
timestamp 1386235218
transform 1 0 816 0 1 66
box 0 0 192 799
<< labels >>
rlabel metal1 0 50 0 60 3 Ir
rlabel metal1 1008 6 1008 16 7 Imm
rlabel metal1 1008 28 1008 38 7 SysBus
rlabel metal1 0 28 0 38 3 SysBus
rlabel metal2 72 0 84 0 1 IrWe
rlabel metal2 792 0 804 0 1 Ext1
rlabel metal2 864 0 876 0 1 ImmSel
rlabel metal2 864 1042 876 1042 5 ImmSel
rlabel metal2 792 1042 804 1042 5 Ext1
rlabel metal2 72 1042 84 1042 5 IrWe
rlabel metal2 744 1042 756 1042 5 Ir
<< end >>
