magic
tech c035u
timestamp 1397224710
<< metal1 >>
rect 805 938 935 948
rect 757 916 887 926
rect 0 96 599 106
rect 613 96 743 106
rect 757 96 791 106
rect 0 29 23 39
rect 37 29 1008 39
rect 928 7 949 17
rect 973 7 1008 17
<< m2contact >>
rect 791 936 805 950
rect 935 936 949 950
rect 743 914 757 928
rect 887 914 901 928
rect 599 94 613 108
rect 743 94 757 108
rect 791 94 805 108
rect 23 28 37 42
rect 959 5 973 19
<< metal2 >>
rect 72 911 84 1111
rect 744 928 756 1111
rect 792 950 804 1111
rect 744 911 756 914
rect 792 911 804 936
rect 864 911 876 1111
rect 888 911 900 914
rect 936 911 948 936
rect 24 42 36 112
rect 72 0 84 112
rect 600 108 612 112
rect 744 108 756 112
rect 792 108 804 112
rect 864 0 876 112
rect 960 19 972 112
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 0 0 1 112
box 0 0 720 799
use rowcrosser rowcrosser_2
timestamp 1397224710
transform 1 0 720 0 1 112
box 0 0 48 799
use rowcrosser rowcrosser_3
timestamp 1397224710
transform 1 0 768 0 1 112
box 0 0 48 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 816 0 1 112
box 0 0 192 799
<< labels >>
rlabel metal2 864 1111 876 1111 5 ImmSel
rlabel metal2 72 1111 84 1111 5 IrWe
rlabel metal2 744 1111 756 1111 5 Ir
rlabel metal2 792 1111 804 1111 5 Ir
rlabel metal1 0 29 0 39 3 SysBus
rlabel metal1 1008 29 1008 39 7 SysBus
rlabel metal1 1008 7 1008 17 7 Imm
rlabel metal1 0 96 0 106 3 Ir
rlabel metal2 864 0 876 0 1 ImmSel
rlabel metal2 72 0 84 0 1 IrWe
<< end >>
