magic
tech c035u
timestamp 1394227191
<< metal1 >>
rect 2496 9240 4526 9250
rect 3591 9195 4861 9205
rect 1288 9115 4166 9125
rect 4745 9059 5223 9070
rect 135 9000 3803 9010
rect 3556 8922 9145 8932
rect 3316 8900 7993 8910
rect 3100 8878 6841 8888
rect 2884 8855 5690 8865
rect 2644 8831 4537 8841
rect 1095 8808 1934 8818
rect 2428 8809 3385 8819
rect 1804 8787 8929 8797
rect 1564 8763 7777 8773
rect 1348 8739 6624 8749
rect 1132 8715 5474 8725
rect 892 8691 4321 8701
rect 676 8670 3169 8680
rect 436 8646 2017 8656
rect 196 8623 865 8633
<< m2contact >>
rect 2482 9239 2496 9253
rect 4526 9239 4540 9253
rect 3577 9194 3591 9208
rect 4861 9193 4876 9207
rect 1273 9112 1288 9126
rect 4166 9115 4180 9129
rect 4726 9055 4745 9072
rect 5223 9058 5239 9073
rect 120 8999 135 9013
rect 3803 8996 3822 9014
rect 3542 8920 3556 8934
rect 9145 8920 9159 8934
rect 3302 8898 3316 8912
rect 7993 8898 8007 8912
rect 3086 8876 3100 8890
rect 6841 8875 6855 8889
rect 2870 8851 2884 8865
rect 5690 8853 5704 8867
rect 2630 8829 2644 8843
rect 4537 8829 4551 8843
rect 1081 8806 1095 8820
rect 1934 8807 1948 8821
rect 2414 8809 2428 8823
rect 3385 8807 3399 8821
rect 1790 8783 1804 8797
rect 8929 8785 8943 8799
rect 1550 8759 1564 8773
rect 7777 8762 7791 8776
rect 1334 8735 1348 8749
rect 6624 8738 6638 8752
rect 1118 8711 1132 8725
rect 5474 8713 5488 8727
rect 878 8691 892 8705
rect 4321 8689 4335 8703
rect 662 8669 676 8683
rect 3169 8667 3183 8681
rect 422 8644 436 8658
rect 2017 8646 2031 8660
rect 182 8623 196 8637
rect 865 8621 879 8635
<< metal2 >>
rect 87 10236 99 10305
rect 111 10236 123 10305
rect 135 10236 147 10305
rect 1839 10236 1851 10305
rect 1863 10236 1875 10305
rect 1887 10236 1899 10305
rect 122 8600 134 8999
rect 183 8637 195 9282
rect 423 8658 435 9282
rect 663 8683 675 9282
rect 879 8705 891 9282
rect 866 8600 878 8621
rect 1082 8600 1094 8806
rect 1119 8725 1131 9282
rect 1274 8600 1286 9112
rect 1335 8749 1347 9282
rect 1551 8773 1563 9282
rect 1791 8797 1803 9282
rect 1935 8821 1947 9282
rect 2018 8600 2030 8646
rect 2175 8631 2187 9283
rect 2415 8823 2427 9282
rect 2483 8664 2495 9239
rect 2631 8843 2643 9282
rect 2871 8865 2883 9282
rect 3087 8890 3099 9282
rect 3303 8912 3315 9282
rect 3543 8934 3555 9282
rect 2426 8652 2495 8664
rect 2175 8619 2246 8631
rect 2234 8600 2246 8619
rect 2426 8594 2438 8652
rect 3170 8600 3182 8667
rect 3386 8600 3398 8807
rect 3578 8599 3590 9194
rect 3807 9014 3819 9282
rect 4167 9129 4179 9282
rect 4527 9253 4539 9288
rect 4863 9207 4875 9283
rect 5223 9073 5235 9283
rect 5559 9098 5571 9282
rect 5895 9158 5907 9282
rect 6255 9244 6267 9282
rect 6255 9232 8006 9244
rect 5895 9146 7046 9158
rect 5559 9086 5894 9098
rect 4322 8600 4334 8689
rect 4538 8600 4550 8829
rect 4730 8595 4742 9055
rect 5474 8600 5486 8713
rect 5690 8600 5702 8853
rect 5882 8600 5894 9086
rect 6626 8600 6638 8738
rect 6842 8600 6854 8875
rect 7034 8600 7046 9146
rect 7994 8912 8006 9232
rect 7778 8600 7790 8762
rect 7994 8600 8006 8898
rect 8930 8600 8942 8785
rect 9146 8600 9158 8920
use decoder decoder_0
timestamp 1394117868
transform 1 0 63 0 1 9282
box 0 0 1752 932
use decoder decoder_1
timestamp 1394117868
transform 1 0 1815 0 1 9282
box 0 0 1752 932
use wdecoder wdecoder_0
timestamp 1394121495
transform 1 0 3687 0 1 9282
box -120 0 2592 989
use regBlock_slice regBlock_slice_0
array 0 0 9385 0 7 1075
timestamp 1394121372
transform 1 0 0 0 1 0
box 0 0 9385 1075
<< labels >>
rlabel metal2 87 10305 99 10305 5 Rs1[0]
rlabel metal2 111 10305 123 10305 5 Rs1[1]
rlabel metal2 135 10305 147 10305 5 Rs1[2]
rlabel metal2 1839 10305 1851 10305 5 Rs2[0]
rlabel metal2 1863 10305 1875 10305 5 Rs2[1]
rlabel metal2 1887 10305 1899 10305 5 Rs2[2]
<< end >>
