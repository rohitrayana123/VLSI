magic
tech c035u
timestamp 1394477934
<< checkpaint >>
rect -1300 21979 16132 21981
rect -1300 21932 16148 21979
rect -1321 17584 16148 21932
rect -1321 17537 16137 17584
rect -1300 17516 16137 17537
rect -1300 -1300 1500 17516
use slice17  slice17_0
timestamp 1394305018
transform 1 0 4334 0 1 18816
box -4329 0 10503 1795
use leftbuf_slice  leftbuf_slice_0
array 0 0 1469 0 15 1176
timestamp 1394477934
transform 1 0 0 0 1 6
box 0 -6 1469 1170
use IrAA  IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394477934
transform 1 0 1469 0 1 9519
box 0 -111 1008 1065
use IrBA  IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394477934
transform 1 0 1469 0 1 5991
box 0 -111 1008 1065
use IrBB  IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394477934
transform 1 0 1469 0 1 112
box 0 -112 1008 1064
use Datapath_slice  Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394475869
transform 1 0 2477 0 1 0
box 0 0 12364 1176
<< end >>
