magic
tech c035u
timestamp 1395325201
use control control_0
timestamp 1395324901
transform 1 0 -622 0 1 21905
box 0 0 28280 8252
use datapath datapath_0
timestamp 1394841956
transform 1 0 48 0 1 0
box -48 0 25445 21228
<< end >>
