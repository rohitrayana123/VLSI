magic
tech c035u
timestamp 1394475379
<< metal1 >>
rect 1261 915 1751 925
rect 1789 915 1943 925
rect 62 893 2626 903
rect 277 871 431 881
rect 445 871 1511 881
rect 1598 870 1895 880
rect 2616 882 2626 893
rect 1981 870 2039 880
rect 397 44 1391 54
rect 1405 44 1703 54
rect 1717 44 2903 54
<< m2contact >>
rect 1247 913 1261 927
rect 1751 913 1765 927
rect 1775 913 1789 927
rect 1943 913 1957 927
rect 48 890 62 904
rect 263 869 277 883
rect 431 869 445 883
rect 1511 869 1525 883
rect 1583 868 1598 882
rect 1895 868 1909 882
rect 1967 869 1981 883
rect 2039 868 2053 882
rect 2614 868 2629 882
rect 383 40 397 54
rect 1391 42 1405 56
rect 1703 42 1717 56
rect 2903 42 2917 56
<< metal2 >>
rect 48 865 60 890
rect 216 865 228 1042
rect 264 865 276 869
rect 360 865 372 1042
rect 432 865 444 869
rect 456 865 540 877
rect 576 865 588 1042
rect 1248 877 1260 913
rect 1104 865 1260 877
rect 1320 865 1332 1042
rect 1488 865 1500 1042
rect 1512 865 1524 869
rect 1560 865 1572 1042
rect 1584 865 1596 868
rect 1752 865 1764 913
rect 1776 865 1788 913
rect 1872 865 1884 1042
rect 1896 865 1908 868
rect 1944 865 1956 913
rect 1968 865 1980 869
rect 2040 865 2052 868
rect 2088 865 2100 1042
rect 2629 868 2772 880
rect 2616 865 2628 868
rect 2760 865 2772 868
rect 2832 865 2844 1042
rect 72 56 84 66
rect 72 44 228 56
rect 216 0 228 44
rect 360 0 372 66
rect 384 54 396 66
rect 576 0 588 66
rect 1320 0 1332 66
rect 1392 56 1404 66
rect 1488 56 1500 66
rect 1680 56 1692 66
rect 1704 56 1716 66
rect 1488 44 1692 56
rect 1488 0 1500 44
rect 1872 0 1884 66
rect 2088 0 2100 66
rect 2616 0 2628 66
rect 2832 0 2844 66
rect 2904 56 2916 66
rect 2904 0 2916 42
use halfadder  halfadder_0
timestamp 1386235204
transform 1 0 0 0 1 66
box 0 0 312 799
use mux2  mux2_2
timestamp 1386235218
transform 1 0 312 0 1 66
box 0 0 192 799
use scanreg  scanreg_0
timestamp 1386241447
transform 1 0 504 0 1 66
box 0 0 720 799
use trisbuf  trisbuf_0
timestamp 1386237216
transform 1 0 1224 0 1 66
box 0 0 216 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 1440 0 1 66
box 0 0 192 799
use mux2  mux2_1
timestamp 1386235218
transform 1 0 1632 0 1 66
box 0 0 192 799
use mux2  mux2_3
timestamp 1386235218
transform 1 0 1824 0 1 66
box 0 0 192 799
use scanreg  scanreg_1
timestamp 1386241447
transform 1 0 2016 0 1 66
box 0 0 720 799
use trisbuf  trisbuf_1
timestamp 1386237216
transform 1 0 2736 0 1 66
box 0 0 216 799
<< labels >>
rlabel metal1 1505 876 1505 876 1 Pc1
rlabel metal1 1745 920 1745 920 1 Lr
rlabel metal2 1488 1042 1500 1042 1 PcSel[0]
rlabel metal2 1320 1042 1332 1042 1 LrEn
rlabel metal2 576 1042 588 1042 1 LrWe
rlabel metal2 360 1042 372 1042 1 LrSel
rlabel metal2 216 1042 228 1042 5 PcIncCout
rlabel metal2 2832 1042 2844 1042 1 PcEn
rlabel metal2 2088 1042 2100 1042 1 PcWe
rlabel metal2 1560 1042 1572 1042 1 ALU
rlabel metal2 1872 1042 1884 1042 1 PcSel[1]
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 2088 0 2100 0 1 PcWe
rlabel metal2 2616 0 2628 0 1 Pc
rlabel metal2 2832 0 2844 0 1 PcEn
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 2904 0 2916 0 1 SysBus
<< end >>
