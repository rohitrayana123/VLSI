../../../Design/Implementation/verilog/behavioural/simple_interface.sv