../../../Design/Implementation/verilog/behavioural/regBlock.sv