magic
tech c035u
timestamp 1396394179
<< metal1 >>
rect 14 19475 14577 19485
rect 37 19451 14770 19461
rect 60 19427 14962 19437
rect 83 19403 15154 19413
rect 106 19379 15346 19389
rect 129 19355 4161 19365
rect 152 19331 4593 19341
rect 175 19307 4977 19317
rect 198 19283 4209 19293
rect 221 19259 4641 19269
rect 244 19235 5025 19245
rect 267 19211 7165 19221
rect 290 19187 7141 19197
rect 7155 19187 22353 19197
rect 313 19163 7117 19173
rect 7131 19163 22545 19173
rect 336 19139 22665 19149
rect 359 19115 22785 19125
rect 2879 17675 2890 17685
rect 14 16831 365 16841
rect 2842 16721 2890 16731
rect 25391 16721 25408 16731
rect 2842 16699 2890 16709
rect 25391 16699 25408 16709
rect 2879 16564 2890 16574
rect 37 15720 365 15730
rect 2842 15610 2890 15620
rect 25391 15610 25408 15620
rect 2842 15588 2890 15598
rect 25391 15588 25408 15598
rect 2879 15453 2890 15463
rect 60 14609 365 14619
rect 2842 14499 2890 14509
rect 25391 14499 25408 14509
rect 2842 14477 2890 14487
rect 25391 14477 25408 14487
rect 2879 14342 2890 14352
rect 83 13498 365 13508
rect 2842 13388 2890 13398
rect 25391 13388 25408 13398
rect 2842 13366 2890 13376
rect 25391 13366 25408 13376
rect 2879 13231 2890 13241
rect 106 12387 365 12397
rect 2842 12277 2890 12287
rect 25391 12277 25408 12287
rect 2842 12255 2890 12265
rect 25391 12255 25408 12265
rect 2879 12120 2890 12130
rect 129 11276 365 11286
rect 2842 11166 2890 11176
rect 25391 11166 25408 11176
rect 2842 11144 2890 11154
rect 25391 11144 25408 11154
rect 2879 11009 2890 11019
rect 152 10165 365 10175
rect 2842 10055 2890 10065
rect 25391 10055 25408 10065
rect 2842 10033 2890 10043
rect 25391 10033 25408 10043
rect 2879 9898 2890 9908
rect 175 9054 365 9064
rect 2842 8944 2890 8954
rect 25391 8944 25408 8954
rect 2842 8922 2890 8932
rect 25391 8922 25408 8932
rect 2879 8787 2890 8797
rect 198 7943 365 7953
rect 2842 7833 2890 7843
rect 25391 7833 25408 7843
rect 2842 7811 2890 7821
rect 25391 7811 25408 7821
rect 2879 7676 2890 7686
rect 221 6832 365 6842
rect 2842 6722 2890 6732
rect 25391 6722 25408 6732
rect 2842 6700 2890 6710
rect 25391 6700 25408 6710
rect 2879 6565 2890 6575
rect 244 5721 365 5731
rect 2842 5611 2890 5621
rect 25391 5611 25408 5621
rect 2842 5589 2890 5599
rect 25391 5589 25408 5599
rect 2879 5454 2890 5464
rect 267 4610 365 4620
rect 2842 4500 2890 4510
rect 25391 4500 25408 4510
rect 2842 4478 2890 4488
rect 25391 4478 25408 4488
rect 2879 4343 2890 4353
rect 290 3499 365 3509
rect 2842 3389 2890 3399
rect 25391 3389 25408 3399
rect 2842 3367 2890 3377
rect 25391 3367 25408 3377
rect 2879 3232 2890 3242
rect 313 2388 365 2398
rect 2842 2278 2890 2288
rect 25391 2278 25408 2288
rect 2842 2256 2890 2266
rect 25391 2256 25408 2266
rect 2879 2121 2890 2131
rect 336 1277 365 1287
rect 2842 1167 2890 1177
rect 25391 1167 25408 1177
rect 2842 1145 2890 1155
rect 25391 1145 25408 1155
rect 2879 1010 2890 1020
rect 359 166 365 176
rect 2842 56 2890 66
rect 25391 56 25408 66
rect 2842 34 2890 44
rect 25391 34 25408 44
rect 570 8 3105 18
rect 17063 7 19713 17
rect 19727 7 19760 17
rect 19774 7 19809 17
rect 19823 7 19857 17
rect 19871 7 19905 17
rect 19919 7 19953 17
rect 19967 7 20001 17
rect 20015 7 20049 17
rect 20063 7 20361 17
rect 20375 7 20409 17
rect 20423 7 20456 17
rect 20470 7 20505 17
rect 20519 7 20817 17
rect 20831 7 20865 17
rect 20879 7 21249 17
rect 21263 7 25186 17
<< m2contact >>
rect 0 19473 14 19487
rect 14577 19474 14591 19488
rect 23 19449 37 19463
rect 14770 19449 14784 19463
rect 46 19425 60 19439
rect 14962 19425 14976 19439
rect 69 19401 83 19415
rect 15154 19401 15168 19415
rect 92 19377 106 19391
rect 15346 19377 15360 19392
rect 115 19353 129 19367
rect 4161 19353 4175 19367
rect 138 19329 152 19343
rect 4593 19329 4607 19343
rect 161 19305 175 19319
rect 4977 19305 4991 19319
rect 184 19281 198 19295
rect 4209 19281 4223 19295
rect 207 19257 221 19271
rect 4641 19257 4655 19271
rect 230 19233 244 19247
rect 5025 19233 5039 19247
rect 253 19209 267 19223
rect 7165 19209 7179 19223
rect 276 19185 290 19199
rect 7141 19185 7155 19199
rect 22353 19185 22367 19199
rect 299 19161 313 19175
rect 7117 19161 7131 19175
rect 22545 19160 22559 19174
rect 322 19137 336 19151
rect 22665 19137 22679 19151
rect 345 19113 359 19127
rect 22785 19113 22799 19127
rect 2865 17673 2879 17687
rect 0 16829 14 16843
rect 2865 16562 2879 16576
rect 23 15718 37 15732
rect 2865 15451 2879 15465
rect 46 14607 60 14621
rect 2865 14340 2879 14354
rect 69 13496 83 13510
rect 2865 13229 2879 13243
rect 92 12385 106 12399
rect 2865 12118 2879 12132
rect 115 11274 129 11288
rect 2865 11007 2879 11021
rect 138 10163 152 10177
rect 2865 9896 2879 9910
rect 161 9052 175 9066
rect 2865 8785 2879 8799
rect 184 7941 198 7955
rect 2865 7674 2879 7688
rect 207 6830 221 6844
rect 2865 6563 2879 6577
rect 230 5719 244 5733
rect 2865 5452 2879 5466
rect 253 4608 267 4622
rect 2865 4341 2879 4355
rect 276 3497 290 3511
rect 2865 3230 2879 3244
rect 299 2386 313 2400
rect 2865 2119 2879 2133
rect 322 1275 336 1289
rect 2865 1008 2879 1022
rect 345 164 359 178
rect 556 6 570 20
rect 3105 5 3119 19
rect 17049 5 17063 19
rect 19713 5 19727 19
rect 19760 5 19774 19
rect 19809 5 19823 19
rect 19857 5 19871 19
rect 19905 5 19919 19
rect 19953 5 19967 19
rect 20001 5 20015 19
rect 20049 5 20063 19
rect 20361 5 20375 19
rect 20409 5 20423 19
rect 20456 5 20470 19
rect 20505 5 20519 19
rect 20817 5 20831 19
rect 20865 5 20879 19
rect 21249 5 21263 19
rect 25186 5 25200 19
<< metal2 >>
rect 1 16843 13 19473
rect 1 0 13 16829
rect 24 15732 36 19449
rect 24 0 36 15718
rect 47 14621 59 19425
rect 47 0 59 14607
rect 70 13510 82 19401
rect 70 0 82 13496
rect 93 12399 105 19377
rect 93 0 105 12385
rect 116 11288 128 19353
rect 116 0 128 11274
rect 139 10177 151 19329
rect 139 0 151 10163
rect 162 9066 174 19305
rect 162 0 174 9052
rect 185 7955 197 19281
rect 185 0 197 7941
rect 208 6844 220 19257
rect 208 0 220 6830
rect 231 5733 243 19233
rect 231 0 243 5719
rect 254 4622 266 19209
rect 254 0 266 4608
rect 277 3511 289 19185
rect 277 0 289 3497
rect 300 2400 312 19161
rect 300 0 312 2386
rect 323 1289 335 19137
rect 323 0 335 1275
rect 346 178 358 19113
rect 370 19105 570 19490
rect 586 19105 598 19490
rect 610 19105 622 19490
rect 634 19105 646 19490
rect 658 19105 670 19490
rect 4138 19105 4150 19490
rect 4162 19105 4174 19353
rect 4210 19105 4222 19281
rect 4378 19105 4390 19490
rect 4594 19105 4606 19329
rect 4642 19105 4654 19257
rect 4978 19105 4990 19305
rect 5026 19105 5038 19233
rect 5338 19105 5350 19490
rect 5530 19105 5542 19490
rect 6564 19105 6576 19490
rect 7118 19105 7130 19161
rect 7142 19105 7154 19185
rect 7166 19105 7178 19209
rect 14555 19105 14567 19490
rect 14579 19105 14591 19474
rect 14771 19105 14783 19449
rect 14819 19105 14831 19490
rect 14963 19105 14975 19425
rect 15155 19105 15167 19401
rect 15347 19105 15359 19377
rect 15539 19105 15551 19490
rect 17338 19105 17350 19490
rect 17530 19105 17542 19490
rect 17602 19105 17614 19490
rect 17698 19105 17710 19490
rect 22354 19105 22366 19185
rect 22546 19105 22558 19160
rect 22666 19105 22678 19137
rect 22786 19105 22798 19113
rect 25186 19105 25386 19490
rect 2866 17603 2878 17673
rect 2866 16492 2878 16562
rect 2866 15381 2878 15451
rect 2866 14270 2878 14340
rect 2866 13159 2878 13229
rect 2866 12048 2878 12118
rect 2866 10937 2878 11007
rect 2866 9826 2878 9896
rect 2866 8715 2878 8785
rect 2866 7604 2878 7674
rect 2866 6493 2878 6563
rect 2866 5382 2878 5452
rect 2866 4271 2878 4341
rect 2866 3160 2878 3230
rect 2866 2049 2878 2119
rect 2866 938 2878 1008
rect 346 0 358 164
rect 370 20 570 27
rect 370 6 556 20
rect 370 0 570 6
rect 586 0 598 27
rect 610 0 622 27
rect 634 0 646 27
rect 658 0 670 27
rect 1906 0 1918 27
rect 2698 0 2710 27
rect 3106 19 3118 27
rect 3250 0 3262 27
rect 3466 0 3478 27
rect 4210 0 4222 27
rect 4378 0 4390 27
rect 4762 0 4774 27
rect 4954 0 4966 27
rect 5170 0 5182 27
rect 5914 0 5926 27
rect 6082 0 6094 27
rect 15490 0 15502 27
rect 15682 0 15694 27
rect 15922 0 15934 27
rect 16570 21 16582 27
rect 16762 21 16774 27
rect 16570 9 16774 21
rect 17050 19 17062 27
rect 19714 19 19726 27
rect 19762 19 19774 27
rect 19810 19 19822 27
rect 19858 19 19870 27
rect 19906 19 19918 27
rect 19954 19 19966 27
rect 20002 19 20014 27
rect 20050 19 20062 27
rect 20362 19 20374 27
rect 20410 19 20422 27
rect 20458 19 20470 27
rect 20506 19 20518 27
rect 20818 19 20830 27
rect 20866 19 20878 27
rect 21250 19 21262 27
rect 23626 0 23638 27
rect 24370 0 24382 27
rect 24586 0 24598 27
rect 24730 0 24742 27
rect 24778 0 24790 27
rect 24826 0 24838 27
rect 24874 0 24886 27
rect 24946 0 24958 27
rect 25186 19 25386 27
rect 25200 5 25386 19
rect 25186 0 25386 5
use slice17 slice17_0
timestamp 1396388721
transform 1 0 370 0 1 17803
box 0 0 25016 1302
use leftbuf_slice leftbuf_slice_15
timestamp 1396389552
transform 1 0 365 0 1 16692
box 0 0 1469 1111
use IrAA IrAA_7
timestamp 1396389886
transform 1 0 1834 0 1 16692
box 0 0 1008 1111
use tielow tielow_0
timestamp 1386086605
transform 1 0 2842 0 1 16804
box 0 0 48 799
use leftbuf_slice leftbuf_slice_14
timestamp 1396389552
transform 1 0 365 0 1 15581
box 0 0 1469 1111
use IrAA IrAA_6
timestamp 1396389886
transform 1 0 1834 0 1 15581
box 0 0 1008 1111
use Datapath_slice Datapath_slice_15
timestamp 1396393905
transform 1 0 2890 0 1 16692
box 0 0 20472 1111
use LLIcell_U LLIcell_U_7
timestamp 1396390011
transform 1 0 23362 0 1 16692
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_11
timestamp 1396394092
transform 1 0 23554 0 1 16692
box 0 0 1837 1111
use tielow tielow_1
timestamp 1386086605
transform 1 0 2842 0 1 15693
box 0 0 48 799
use leftbuf_slice leftbuf_slice_13
timestamp 1396389552
transform 1 0 365 0 1 14470
box 0 0 1469 1111
use IrAA IrAA_5
timestamp 1396389886
transform 1 0 1834 0 1 14470
box 0 0 1008 1111
use Datapath_slice Datapath_slice_14
timestamp 1396393905
transform 1 0 2890 0 1 15581
box 0 0 20472 1111
use LLIcell_U LLIcell_U_6
timestamp 1396390011
transform 1 0 23362 0 1 15581
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_10
timestamp 1396394092
transform 1 0 23554 0 1 15581
box 0 0 1837 1111
use tielow tielow_2
timestamp 1386086605
transform 1 0 2842 0 1 14582
box 0 0 48 799
use leftbuf_slice leftbuf_slice_12
timestamp 1396389552
transform 1 0 365 0 1 13359
box 0 0 1469 1111
use IrAA IrAA_4
timestamp 1396389886
transform 1 0 1834 0 1 13359
box 0 0 1008 1111
use Datapath_slice Datapath_slice_13
timestamp 1396393905
transform 1 0 2890 0 1 14470
box 0 0 20472 1111
use LLIcell_U LLIcell_U_5
timestamp 1396390011
transform 1 0 23362 0 1 14470
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_9
timestamp 1396394092
transform 1 0 23554 0 1 14470
box 0 0 1837 1111
use tielow tielow_3
timestamp 1386086605
transform 1 0 2842 0 1 13471
box 0 0 48 799
use leftbuf_slice leftbuf_slice_11
timestamp 1396389552
transform 1 0 365 0 1 12248
box 0 0 1469 1111
use IrAA IrAA_3
timestamp 1396389886
transform 1 0 1834 0 1 12248
box 0 0 1008 1111
use Datapath_slice Datapath_slice_12
timestamp 1396393905
transform 1 0 2890 0 1 13359
box 0 0 20472 1111
use LLIcell_U LLIcell_U_4
timestamp 1396390011
transform 1 0 23362 0 1 13359
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_8
timestamp 1396394092
transform 1 0 23554 0 1 13359
box 0 0 1837 1111
use tielow tielow_4
timestamp 1386086605
transform 1 0 2842 0 1 12360
box 0 0 48 799
use leftbuf_slice leftbuf_slice_10
timestamp 1396389552
transform 1 0 365 0 1 11137
box 0 0 1469 1111
use IrAA IrAA_2
timestamp 1396389886
transform 1 0 1834 0 1 11137
box 0 0 1008 1111
use Datapath_slice Datapath_slice_11
timestamp 1396393905
transform 1 0 2890 0 1 12248
box 0 0 20472 1111
use LLIcell_U LLIcell_U_3
timestamp 1396390011
transform 1 0 23362 0 1 12248
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_7
timestamp 1396394092
transform 1 0 23554 0 1 12248
box 0 0 1837 1111
use tielow tielow_5
timestamp 1386086605
transform 1 0 2842 0 1 11249
box 0 0 48 799
use leftbuf_slice leftbuf_slice_9
timestamp 1396389552
transform 1 0 365 0 1 10026
box 0 0 1469 1111
use IrAA IrAA_1
timestamp 1396389886
transform 1 0 1834 0 1 10026
box 0 0 1008 1111
use Datapath_slice Datapath_slice_10
timestamp 1396393905
transform 1 0 2890 0 1 11137
box 0 0 20472 1111
use LLIcell_U LLIcell_U_2
timestamp 1396390011
transform 1 0 23362 0 1 11137
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_6
timestamp 1396394092
transform 1 0 23554 0 1 11137
box 0 0 1837 1111
use tielow tielow_6
timestamp 1386086605
transform 1 0 2842 0 1 10138
box 0 0 48 799
use leftbuf_slice leftbuf_slice_8
timestamp 1396389552
transform 1 0 365 0 1 8915
box 0 0 1469 1111
use IrAA IrAA_0
timestamp 1396389886
transform 1 0 1834 0 1 8915
box 0 0 1008 1111
use Datapath_slice Datapath_slice_9
timestamp 1396393905
transform 1 0 2890 0 1 10026
box 0 0 20472 1111
use LLIcell_U LLIcell_U_1
timestamp 1396390011
transform 1 0 23362 0 1 10026
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_5
timestamp 1396394092
transform 1 0 23554 0 1 10026
box 0 0 1837 1111
use tielow tielow_7
timestamp 1386086605
transform 1 0 2842 0 1 9027
box 0 0 48 799
use leftbuf_slice leftbuf_slice_7
timestamp 1396389552
transform 1 0 365 0 1 7804
box 0 0 1469 1111
use IrBA IrBA_2
timestamp 1396389912
transform 1 0 1834 0 1 7804
box 0 0 1008 1111
use Datapath_slice Datapath_slice_8
timestamp 1396393905
transform 1 0 2890 0 1 8915
box 0 0 20472 1111
use LLIcell_U LLIcell_U_0
timestamp 1396390011
transform 1 0 23362 0 1 8915
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_4
timestamp 1396394092
transform 1 0 23554 0 1 8915
box 0 0 1837 1111
use tielow tielow_8
timestamp 1386086605
transform 1 0 2842 0 1 7916
box 0 0 48 799
use leftbuf_slice leftbuf_slice_6
timestamp 1396389552
transform 1 0 365 0 1 6693
box 0 0 1469 1111
use IrBA IrBA_1
timestamp 1396389912
transform 1 0 1834 0 1 6693
box 0 0 1008 1111
use Datapath_slice Datapath_slice_7
timestamp 1396393905
transform 1 0 2890 0 1 7804
box 0 0 20472 1111
use LLIcell_L LLIcell_L_7
timestamp 1396390031
transform 1 0 23362 0 1 7804
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_3
timestamp 1396394092
transform 1 0 23554 0 1 7804
box 0 0 1837 1111
use tielow tielow_9
timestamp 1386086605
transform 1 0 2842 0 1 6805
box 0 0 48 799
use leftbuf_slice leftbuf_slice_5
timestamp 1396389552
transform 1 0 365 0 1 5582
box 0 0 1469 1111
use IrBA IrBA_0
timestamp 1396389912
transform 1 0 1834 0 1 5582
box 0 0 1008 1111
use Datapath_slice Datapath_slice_6
timestamp 1396393905
transform 1 0 2890 0 1 6693
box 0 0 20472 1111
use LLIcell_L LLIcell_L_6
timestamp 1396390031
transform 1 0 23362 0 1 6693
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_2
timestamp 1396394092
transform 1 0 23554 0 1 6693
box 0 0 1837 1111
use tielow tielow_10
timestamp 1386086605
transform 1 0 2842 0 1 5694
box 0 0 48 799
use leftbuf_slice leftbuf_slice_4
timestamp 1396389552
transform 1 0 365 0 1 4471
box 0 0 1469 1111
use IrBB IrBB_4
timestamp 1396389938
transform 1 0 1834 0 1 4471
box 0 0 1008 1111
use Datapath_slice Datapath_slice_5
timestamp 1396393905
transform 1 0 2890 0 1 5582
box 0 0 20472 1111
use LLIcell_L LLIcell_L_5
timestamp 1396390031
transform 1 0 23362 0 1 5582
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_1
timestamp 1396394092
transform 1 0 23554 0 1 5582
box 0 0 1837 1111
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 2842 0 1 4583
box 0 0 48 799
use leftbuf_slice leftbuf_slice_3
timestamp 1396389552
transform 1 0 365 0 1 3360
box 0 0 1469 1111
use IrBB IrBB_3
timestamp 1396389938
transform 1 0 1834 0 1 3360
box 0 0 1008 1111
use Datapath_slice Datapath_slice_4
timestamp 1396393905
transform 1 0 2890 0 1 4471
box 0 0 20472 1111
use LLIcell_L LLIcell_L_4
timestamp 1396390031
transform 1 0 23362 0 1 4471
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_0
timestamp 1396394092
transform 1 0 23554 0 1 4471
box 0 0 1837 1111
use tielow tielow_12
timestamp 1386086605
transform 1 0 2842 0 1 3472
box 0 0 48 799
use leftbuf_slice leftbuf_slice_2
timestamp 1396389552
transform 1 0 365 0 1 2249
box 0 0 1469 1111
use IrBB IrBB_2
timestamp 1396389938
transform 1 0 1834 0 1 2249
box 0 0 1008 1111
use Datapath_slice Datapath_slice_3
timestamp 1396393905
transform 1 0 2890 0 1 3360
box 0 0 20472 1111
use LLIcell_L LLIcell_L_3
timestamp 1396390031
transform 1 0 23362 0 1 3360
box 0 0 192 1111
use Datapath_end_low Datapath_end_low_3
timestamp 1396394133
transform 1 0 23554 0 1 3360
box 0 0 1837 1111
use tielow tielow_13
timestamp 1386086605
transform 1 0 2842 0 1 2361
box 0 0 48 799
use leftbuf_slice leftbuf_slice_1
timestamp 1396389552
transform 1 0 365 0 1 1138
box 0 0 1469 1111
use IrBB IrBB_1
timestamp 1396389938
transform 1 0 1834 0 1 1138
box 0 0 1008 1111
use Datapath_slice Datapath_slice_2
timestamp 1396393905
transform 1 0 2890 0 1 2249
box 0 0 20472 1111
use LLIcell_L LLIcell_L_2
timestamp 1396390031
transform 1 0 23362 0 1 2249
box 0 0 192 1111
use Datapath_end_low Datapath_end_low_2
timestamp 1396394133
transform 1 0 23554 0 1 2249
box 0 0 1837 1111
use tielow tielow_14
timestamp 1386086605
transform 1 0 2842 0 1 1250
box 0 0 48 799
use leftbuf_slice leftbuf_slice_0
timestamp 1396389552
transform 1 0 365 0 1 27
box 0 0 1469 1111
use IrBB IrBB_0
timestamp 1396389938
transform 1 0 1834 0 1 27
box 0 0 1008 1111
use Datapath_slice Datapath_slice_1
timestamp 1396393905
transform 1 0 2890 0 1 1138
box 0 0 20472 1111
use LLIcell_L LLIcell_L_1
timestamp 1396390031
transform 1 0 23362 0 1 1138
box 0 0 192 1111
use Datapath_end_low Datapath_end_low_1
timestamp 1396394133
transform 1 0 23554 0 1 1138
box 0 0 1837 1111
use tielow tielow_15
timestamp 1386086605
transform 1 0 2842 0 1 139
box 0 0 48 799
use Datapath_slice Datapath_slice_0
timestamp 1396393905
transform 1 0 2890 0 1 27
box 0 0 20472 1111
use LLIcell_L LLIcell_L_0
timestamp 1396390031
transform 1 0 23362 0 1 27
box 0 0 192 1111
use Datapath_end_low Datapath_end_low_0
timestamp 1396394133
transform 1 0 23554 0 1 27
box 0 0 1837 1111
<< labels >>
rlabel metal2 1 0 13 0 1 Ir[15]
rlabel metal2 24 0 36 0 1 Ir[14]
rlabel metal2 47 0 59 0 1 Ir[13]
rlabel metal2 70 0 82 0 1 Ir[12]
rlabel metal2 93 0 105 0 1 Ir[11]
rlabel metal2 116 0 128 0 1 Ir[10]
rlabel metal2 139 0 151 0 1 Ir[9]
rlabel metal2 162 0 174 0 1 Ir[8]
rlabel metal2 185 0 197 0 1 Ir[7]
rlabel metal2 208 0 220 0 1 Ir[6]
rlabel metal2 231 0 243 0 1 Ir[5]
rlabel metal2 254 0 266 0 1 Ir[4]
rlabel metal2 277 0 289 0 1 Ir[3]
rlabel metal2 300 0 312 0 1 Ir[2]
rlabel metal2 323 0 335 0 1 Ir[1]
rlabel metal2 346 0 358 0 1 Ir[0]
rlabel metal2 658 0 670 0 1 nReset
rlabel metal2 634 0 646 0 1 Clock
rlabel metal2 610 0 622 0 1 Test
rlabel metal2 586 0 598 0 1 SDI
rlabel metal2 370 0 570 0 1 Vdd!
rlabel metal2 24586 0 24598 0 1 MemEn
rlabel metal2 24946 0 24958 0 1 StatusRegEn
rlabel metal2 24730 0 24742 0 1 StatusReg[3]
rlabel metal2 24778 0 24790 0 1 StatusReg[2]
rlabel metal2 24826 0 24838 0 1 StatusReg[1]
rlabel metal2 24874 0 24886 0 1 StatusReg[0]
rlabel metal2 25186 0 25386 0 1 GND!
rlabel metal2 4210 0 4222 0 1 LrEn
rlabel metal2 4378 0 4390 0 1 PcSel[0]
rlabel metal2 4762 0 4774 0 1 PcSel[1]
rlabel metal2 23626 0 23638 0 1 AluWe
rlabel metal2 24370 0 24382 0 1 AluEn
rlabel metal2 5170 0 5182 0 1 PcWe
rlabel metal2 4954 0 4966 0 1 PcSel[2]
rlabel metal2 5914 0 5926 0 1 PcEn
rlabel metal2 6082 0 6094 0 1 WdSel
rlabel metal2 15490 0 15502 0 1 Op1Sel
rlabel metal2 15682 0 15694 0 1 Op2Sel[0]
rlabel metal2 15922 0 15934 0 1 Op2Sel[1]
rlabel metal2 1906 0 1918 0 1 IrWe
rlabel metal2 2698 0 2710 0 1 ImmSel
rlabel metal2 3466 0 3478 0 1 LrWe
rlabel metal2 3250 0 3262 0 1 LrSel
rlabel metal1 25408 34 25408 44 7 DataIn[0]
rlabel metal1 25408 56 25408 66 7 DataOut[0]
rlabel metal1 25408 1145 25408 1155 7 DataIn[1]
rlabel metal1 25408 1167 25408 1177 7 DataOut[1]
rlabel metal1 25408 2278 25408 2288 7 DataOut[2]
rlabel metal1 25408 2256 25408 2266 7 DataIn[2]
rlabel metal1 25408 3389 25408 3399 7 DataOut[3]
rlabel metal1 25408 3367 25408 3377 7 DataIn[3]
rlabel metal1 25408 4500 25408 4510 7 DataOut[4]
rlabel metal1 25408 4478 25408 4488 7 DataIn[4]
rlabel metal1 25408 5611 25408 5621 7 DataOut[5]
rlabel metal1 25408 5589 25408 5599 7 DataIn[5]
rlabel metal1 25408 6722 25408 6732 7 DataOut[6]
rlabel metal1 25408 6700 25408 6710 7 DataIn[6]
rlabel metal1 25408 7833 25408 7843 7 DataOut[7]
rlabel metal1 25408 7811 25408 7821 7 DataIn[7]
rlabel metal1 25408 8944 25408 8954 7 DataOut[8]
rlabel metal1 25408 8922 25408 8932 7 DataIn[8]
rlabel metal1 25408 10055 25408 10065 7 DataOut[9]
rlabel metal1 25408 10033 25408 10043 7 DataIn[9]
rlabel metal1 25408 11166 25408 11176 7 DataOut[10]
rlabel metal1 25408 11144 25408 11154 7 DataIn[10]
rlabel metal1 25408 12277 25408 12287 7 DataOut[11]
rlabel metal1 25408 12255 25408 12265 7 DataIn[11]
rlabel metal1 25408 13388 25408 13398 7 DataOut[12]
rlabel metal1 25408 13366 25408 13376 7 DataIn[12]
rlabel metal1 25408 14499 25408 14509 7 DataOut[13]
rlabel metal1 25408 14477 25408 14487 7 DataIn[13]
rlabel metal1 25408 15610 25408 15620 7 DataOut[14]
rlabel metal1 25408 15588 25408 15598 7 DataIn[14]
rlabel metal1 25408 16721 25408 16731 7 DataOut[15]
rlabel metal1 25408 16699 25408 16709 7 DataIn[15]
rlabel metal2 6 19178 6 19178 1 Ir[15]
rlabel metal2 30 19177 30 19177 1 Ir[14]
rlabel metal2 53 19177 53 19177 1 Ir[13]
rlabel metal2 76 19178 76 19178 1 Ir[12]
rlabel metal2 99 19178 99 19178 1 Ir[11]
rlabel metal2 122 19177 122 19177 1 Ir[10]
rlabel metal2 145 19178 145 19178 1 Ir[9]
rlabel metal2 168 19178 168 19178 1 Ir[8]
rlabel metal2 191 19180 191 19180 1 Ir[7]
rlabel metal2 214 19181 214 19181 1 Ir[6]
rlabel metal2 237 19182 237 19182 1 Ir[5]
rlabel metal2 260 19183 260 19183 1 Ir[4]
rlabel metal2 283 19182 283 19182 1 Ir[3]
rlabel metal2 22792 19108 22792 19108 1 Ir[0]
rlabel metal2 22671 19130 22671 19130 1 Ir[1]
rlabel metal2 22551 19155 22551 19155 1 Ir[2]
rlabel metal2 22360 19180 22360 19180 1 Ir[3]
rlabel metal2 14968 19419 14968 19419 1 Ir[13]
rlabel metal2 15161 19395 15161 19395 1 Ir[12]
rlabel metal2 15353 19370 15353 19370 1 Ir[11]
rlabel metal2 14775 19442 14775 19442 1 Ir[14]
rlabel metal2 14584 19467 14584 19467 1 Ir[15]
rlabel metal2 7122 19153 7122 19153 1 Ir[2]
rlabel metal2 7148 19177 7148 19177 1 Ir[3]
rlabel metal2 7171 19201 7171 19201 1 Ir[4]
rlabel metal2 4216 19273 4216 19273 1 Ir[7]
rlabel metal2 4167 19346 4167 19346 1 Ir[10]
rlabel metal2 4648 19250 4648 19250 1 Ir[6]
rlabel metal2 4599 19321 4599 19321 1 Ir[9]
rlabel metal2 4983 19298 4983 19298 1 Ir[8]
rlabel metal2 5033 19227 5033 19227 1 Ir[5]
rlabel metal2 6564 19490 6576 19490 5 RegWe
rlabel metal2 586 19490 598 19490 5 SDO
rlabel metal2 370 19490 570 19490 5 Vdd!
rlabel metal2 658 19490 670 19490 1 nReset
rlabel metal2 634 19490 646 19490 1 Clock
rlabel metal2 610 19490 622 19490 1 Test
rlabel metal2 17698 19490 17710 19490 5 Flags[0]
rlabel metal2 17602 19490 17614 19490 5 Flags[3]
rlabel metal2 17530 19490 17542 19490 5 Flags[1]
rlabel metal2 17338 19490 17350 19490 5 Flags[2]
rlabel metal2 14819 19490 14831 19490 5 AluOR[0]
rlabel metal2 14555 19490 14567 19490 5 AluOR[1]
rlabel metal2 15539 19490 15551 19490 5 CFlag
rlabel metal2 4138 19490 4150 19490 5 Rs1Sel[0]
rlabel metal2 4378 19490 4390 19490 5 Rs1Sel[1]
rlabel metal2 5338 19490 5350 19490 5 RwSel[0]
rlabel metal2 5530 19490 5542 19490 5 RwSel[1]
rlabel metal2 25186 19490 25386 19490 1 GND!
<< end >>
