magic
tech c035u
timestamp 1394287323
<< metal1 >>
rect 1371 900 1861 910
rect 1899 900 2053 910
rect 172 878 2736 888
rect 387 856 541 866
rect 555 856 1621 866
rect 1708 855 2005 865
rect 2726 867 2736 878
rect 2091 855 2149 865
rect 0 833 110 843
rect 3062 833 3127 843
rect 0 772 110 797
rect 3062 772 3127 797
rect 0 127 110 152
rect 3062 127 3127 152
rect 0 104 110 114
rect 3062 104 3127 114
rect 0 81 110 91
rect 3062 81 3127 91
rect 0 58 110 68
rect 3062 58 3127 68
rect 0 27 493 37
rect 507 27 1500 37
rect 1516 27 1813 37
rect 1827 27 3012 37
rect 3028 27 3127 37
<< m2contact >>
rect 1357 898 1371 912
rect 1861 898 1875 912
rect 1885 898 1899 912
rect 2053 898 2067 912
rect 158 875 172 889
rect 373 854 387 868
rect 541 854 555 868
rect 1621 854 1635 868
rect 1693 853 1708 867
rect 2005 853 2019 867
rect 2077 854 2091 868
rect 2149 853 2163 867
rect 2724 853 2739 867
rect 493 26 507 40
rect 1500 26 1516 40
rect 1813 25 1827 39
rect 3012 25 3028 39
<< metal2 >>
rect 158 850 170 875
rect 326 850 338 924
rect 374 850 386 854
rect 470 850 482 924
rect 542 850 554 854
rect 566 850 650 862
rect 686 850 698 924
rect 1358 862 1370 898
rect 1214 850 1370 862
rect 1430 850 1442 924
rect 1598 850 1610 924
rect 1622 850 1634 854
rect 1670 850 1682 924
rect 1694 850 1706 853
rect 1862 850 1874 898
rect 1886 850 1898 898
rect 1982 850 1994 924
rect 2006 850 2018 853
rect 2054 850 2066 898
rect 2078 850 2090 854
rect 2150 850 2162 853
rect 2198 850 2210 924
rect 2739 853 2882 865
rect 2726 850 2738 853
rect 2870 850 2882 853
rect 2942 850 2954 924
rect 182 41 194 51
rect 182 29 338 41
rect 326 0 338 29
rect 470 0 482 51
rect 494 40 506 51
rect 686 0 698 51
rect 1430 0 1442 51
rect 1502 40 1514 51
rect 1598 41 1610 51
rect 1790 41 1802 51
rect 1598 29 1802 41
rect 1814 39 1826 51
rect 1598 0 1610 29
rect 1982 0 1994 51
rect 2198 0 2210 51
rect 2726 0 2738 51
rect 2942 0 2954 51
rect 3014 39 3026 51
use halfadder halfadder_0
timestamp 1386235204
transform 1 0 110 0 1 51
box 0 0 312 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 422 0 1 51
box 0 0 192 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 614 0 1 51
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 1334 0 1 51
box 0 0 216 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 1550 0 1 51
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 1742 0 1 51
box 0 0 192 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 1934 0 1 51
box 0 0 192 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 2126 0 1 51
box 0 0 720 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 2846 0 1 51
box 0 0 216 799
<< labels >>
rlabel metal1 0 772 0 797 3 Vdd!
rlabel metal1 0 833 0 843 3 ScanReturn
rlabel metal1 0 58 0 68 3 nReset
rlabel metal1 0 81 0 91 3 Test
rlabel metal1 0 104 0 114 3 Clock
rlabel metal1 0 127 0 152 3 GND!
rlabel metal2 326 0 338 0 1 PcIncCin
rlabel metal2 470 0 482 0 1 LrSel
rlabel metal2 686 0 698 0 1 LrWe
rlabel metal2 1430 0 1442 0 1 LrEn
rlabel metal2 1598 0 1610 0 1 PcSel[0]
rlabel metal1 3127 772 3127 797 7 Vdd!
rlabel metal1 3127 833 3127 843 7 ScanReturn
rlabel metal1 3127 127 3127 152 7 GND!
rlabel metal1 3127 58 3127 68 7 nReset
rlabel metal1 3127 81 3127 91 7 Test
rlabel metal1 3127 104 3127 114 7 Clock
rlabel metal2 2198 0 2210 0 1 PcWe
rlabel metal2 2726 0 2738 0 1 Pc
rlabel metal2 2942 0 2954 0 1 PcEn
rlabel metal2 1982 0 1994 0 1 PcSel[1]
rlabel metal1 1615 861 1615 861 1 Pc1
rlabel metal1 1855 905 1855 905 1 Lr
rlabel metal2 1598 924 1610 924 1 PcSel[0]
rlabel metal2 1430 924 1442 924 1 LrEn
rlabel metal2 686 924 698 924 1 LrWe
rlabel metal2 470 924 482 924 1 LrSel
rlabel metal2 326 924 338 924 5 PcIncCout
rlabel metal2 2942 924 2954 924 1 PcEn
rlabel metal2 2198 924 2210 924 1 PcWe
rlabel metal2 1670 924 1682 924 1 ALU
rlabel metal2 1982 924 1994 924 1 PcSel[1]
rlabel metal1 3127 27 3127 37 7 SysBus
rlabel metal1 0 27 0 37 3 SysBus
<< end >>
