magic
tech c035u
timestamp 1394305018
use slice17  slice17_0
timestamp 1394305018
transform 1 0 4338 0 1 17245
box -4329 0 10503 1795
use Datapath_slice  Datapath_slice_0
array 0 0 14841 0 15 1079
timestamp 1394303457
transform 1 0 4 0 1 -19
box 0 0 14841 1079
<< end >>
