magic
tech c035u
timestamp 1394709079
use Datapath/datapath datapath_0
timestamp 1394643424
transform 1 0 21 0 1 19
box 0 0 25013 22218
use Control/control_ROUTED control_ROUTED_0
timestamp 1394708833
transform 1 0 -62624 0 1 -6683
box 0 -823 51336 3997
<< end >>
