magic
tech c035u
timestamp 1395690245
<< metal1 >>
rect 14 20557 14577 20567
rect 37 20533 14770 20543
rect 60 20509 14962 20519
rect 83 20485 15154 20495
rect 106 20461 15346 20471
rect 129 20437 4161 20447
rect 152 20413 4593 20423
rect 175 20389 4977 20399
rect 198 20365 4209 20375
rect 221 20341 4641 20351
rect 244 20317 5025 20327
rect 267 20293 7165 20303
rect 290 20269 7141 20279
rect 7155 20269 22353 20279
rect 313 20245 7117 20255
rect 7131 20245 22545 20255
rect 336 20221 22665 20231
rect 359 20197 22785 20207
rect 23578 18848 23770 18858
rect 3095 18737 3106 18747
rect 14 17850 365 17860
rect 3058 17784 3106 17794
rect 23578 17784 23770 17794
rect 25391 17784 25408 17794
rect 3058 17762 3106 17772
rect 3058 17718 3106 17728
rect 23578 17718 23770 17728
rect 25391 17718 25408 17728
rect 23578 17672 23770 17682
rect 3095 17561 3106 17571
rect 37 16674 365 16684
rect 3058 16608 3106 16618
rect 23578 16608 23770 16618
rect 25391 16608 25408 16618
rect 3058 16586 3106 16596
rect 3058 16542 3106 16552
rect 23578 16542 23770 16552
rect 25391 16542 25408 16552
rect 23578 16496 23770 16506
rect 3095 16385 3106 16395
rect 60 15498 365 15508
rect 3058 15432 3106 15442
rect 23578 15432 23770 15442
rect 25391 15432 25408 15442
rect 3058 15410 3106 15420
rect 3058 15366 3106 15376
rect 23578 15366 23770 15376
rect 25391 15366 25408 15376
rect 23578 15320 23770 15330
rect 3095 15209 3106 15219
rect 83 14322 365 14332
rect 3058 14256 3106 14266
rect 23578 14256 23770 14266
rect 25391 14256 25408 14266
rect 3058 14234 3106 14244
rect 3058 14190 3106 14200
rect 23578 14190 23770 14200
rect 25391 14190 25408 14200
rect 23578 14144 23770 14154
rect 3095 14033 3106 14043
rect 106 13146 365 13156
rect 3058 13080 3106 13090
rect 23578 13080 23770 13090
rect 25391 13080 25408 13090
rect 3058 13058 3106 13068
rect 3058 13014 3106 13024
rect 23578 13014 23770 13024
rect 25391 13014 25408 13024
rect 23578 12968 23770 12978
rect 3095 12857 3106 12867
rect 129 11970 365 11980
rect 3058 11904 3106 11914
rect 23578 11904 23770 11914
rect 25391 11904 25408 11914
rect 3058 11882 3106 11892
rect 3058 11838 3106 11848
rect 23578 11838 23770 11848
rect 25391 11838 25408 11848
rect 23578 11792 23770 11802
rect 3095 11681 3106 11691
rect 152 10794 365 10804
rect 3058 10728 3106 10738
rect 23578 10728 23770 10738
rect 25391 10728 25408 10738
rect 3058 10706 3106 10716
rect 3058 10662 3106 10672
rect 23578 10662 23770 10672
rect 25391 10662 25408 10672
rect 23578 10616 23770 10626
rect 3095 10505 3106 10515
rect 175 9618 365 9628
rect 3058 9552 3106 9562
rect 23578 9552 23770 9562
rect 25391 9552 25408 9562
rect 3058 9530 3106 9540
rect 3058 9486 3106 9496
rect 23578 9486 23770 9496
rect 25391 9486 25408 9496
rect 23578 9440 23770 9450
rect 3095 9329 3106 9339
rect 198 8442 365 8452
rect 3058 8376 3106 8386
rect 23578 8376 23770 8386
rect 25391 8376 25408 8386
rect 3058 8354 3106 8364
rect 3058 8310 3106 8320
rect 23578 8310 23770 8320
rect 25391 8310 25408 8320
rect 23578 8264 23770 8274
rect 3095 8153 3106 8163
rect 221 7266 365 7276
rect 3058 7200 3106 7210
rect 23578 7200 23770 7210
rect 25391 7200 25408 7210
rect 3058 7178 3106 7188
rect 3058 7134 3106 7144
rect 23578 7134 23770 7144
rect 25391 7134 25408 7144
rect 23578 7088 23770 7098
rect 3095 6977 3106 6987
rect 244 6090 365 6100
rect 3058 6024 3106 6034
rect 23578 6024 23770 6034
rect 25391 6024 25408 6034
rect 3058 6002 3106 6012
rect 3058 5958 3106 5968
rect 23578 5958 23770 5968
rect 25391 5958 25408 5968
rect 23578 5912 23770 5922
rect 3095 5801 3106 5811
rect 267 4914 365 4924
rect 3058 4848 3106 4858
rect 23578 4848 23770 4858
rect 25391 4848 25408 4858
rect 3058 4826 3106 4836
rect 3058 4782 3106 4792
rect 23578 4782 23770 4792
rect 25391 4782 25408 4792
rect 23578 4736 23770 4746
rect 3095 4625 3106 4635
rect 290 3738 365 3748
rect 3058 3672 3106 3682
rect 23578 3672 23770 3682
rect 25391 3672 25408 3682
rect 3058 3650 3106 3660
rect 3058 3606 3106 3616
rect 23578 3606 23770 3616
rect 25391 3606 25408 3616
rect 23578 3560 23770 3570
rect 3095 3449 3106 3459
rect 313 2562 365 2572
rect 3058 2496 3106 2506
rect 23578 2496 23770 2506
rect 25391 2496 25408 2506
rect 3058 2474 3106 2484
rect 3058 2430 3106 2440
rect 23578 2430 23770 2440
rect 25391 2430 25408 2440
rect 23578 2384 23770 2394
rect 3095 2273 3106 2283
rect 336 1386 365 1396
rect 3058 1320 3106 1330
rect 23578 1320 23770 1330
rect 25391 1320 25408 1330
rect 3058 1298 3106 1308
rect 3058 1254 3106 1264
rect 23578 1254 23770 1264
rect 25391 1254 25408 1264
rect 23578 1208 23770 1218
rect 3095 1097 3106 1107
rect 359 210 365 220
rect 3058 144 3106 154
rect 23578 144 23770 154
rect 25391 144 25408 154
rect 3058 122 3106 132
rect 3058 78 3106 88
rect 23578 78 23770 88
rect 25391 78 25408 88
rect 2055 29 17265 39
rect 17279 29 19929 39
rect 19943 29 19976 39
rect 19990 29 20025 39
rect 20039 29 20073 39
rect 20087 29 20121 39
rect 20135 29 20169 39
rect 20183 29 20217 39
rect 20231 29 20265 39
rect 20279 29 20577 39
rect 20591 29 20625 39
rect 20639 29 20672 39
rect 20686 29 20721 39
rect 20735 29 21033 39
rect 21047 29 21081 39
rect 21095 29 21465 39
rect 21479 29 25186 39
rect 570 8 3321 18
<< m2contact >>
rect 0 20555 14 20569
rect 14577 20556 14591 20570
rect 23 20531 37 20545
rect 14770 20531 14784 20545
rect 46 20507 60 20521
rect 14962 20507 14976 20521
rect 69 20483 83 20497
rect 15154 20483 15168 20497
rect 92 20459 106 20473
rect 15346 20459 15360 20474
rect 115 20435 129 20449
rect 4161 20435 4175 20449
rect 138 20411 152 20425
rect 4593 20411 4607 20425
rect 161 20387 175 20401
rect 4977 20387 4991 20401
rect 184 20363 198 20377
rect 4209 20363 4223 20377
rect 207 20339 221 20353
rect 4641 20339 4655 20353
rect 230 20315 244 20329
rect 5025 20315 5039 20329
rect 253 20291 267 20305
rect 7165 20291 7179 20305
rect 276 20267 290 20281
rect 7141 20267 7155 20281
rect 22353 20267 22367 20281
rect 299 20243 313 20257
rect 7117 20243 7131 20257
rect 22545 20242 22559 20256
rect 322 20219 336 20233
rect 22665 20219 22679 20233
rect 345 20195 359 20209
rect 22785 20195 22799 20209
rect 3081 18735 3095 18749
rect 0 17848 14 17862
rect 3081 17559 3095 17573
rect 23 16672 37 16686
rect 3081 16383 3095 16397
rect 46 15496 60 15510
rect 3081 15207 3095 15221
rect 69 14320 83 14334
rect 3081 14031 3095 14045
rect 92 13144 106 13158
rect 3081 12855 3095 12869
rect 115 11968 129 11982
rect 3081 11679 3095 11693
rect 138 10792 152 10806
rect 3081 10503 3095 10517
rect 161 9616 175 9630
rect 3081 9327 3095 9341
rect 184 8440 198 8454
rect 3081 8151 3095 8165
rect 207 7264 221 7278
rect 3081 6975 3095 6989
rect 230 6088 244 6102
rect 3081 5799 3095 5813
rect 253 4912 267 4926
rect 3081 4623 3095 4637
rect 276 3736 290 3750
rect 3081 3447 3095 3461
rect 299 2560 313 2574
rect 3081 2271 3095 2285
rect 322 1384 336 1398
rect 3081 1095 3095 1109
rect 345 208 359 222
rect 17265 27 17279 41
rect 19929 27 19943 41
rect 19976 27 19990 41
rect 20025 27 20039 41
rect 20073 27 20087 41
rect 20121 27 20135 41
rect 20169 27 20183 41
rect 20217 27 20231 41
rect 20265 27 20279 41
rect 20577 27 20591 41
rect 20625 27 20639 41
rect 20672 27 20686 41
rect 20721 27 20735 41
rect 21033 27 21047 41
rect 21081 27 21095 41
rect 21465 27 21479 41
rect 25186 27 25200 41
rect 556 6 570 20
rect 3321 5 3335 19
<< metal2 >>
rect 1 17862 13 20555
rect 1 0 13 17848
rect 24 16686 36 20531
rect 24 0 36 16672
rect 47 15510 59 20507
rect 47 0 59 15496
rect 70 14334 82 20483
rect 70 0 82 14320
rect 93 13158 105 20459
rect 93 0 105 13144
rect 116 11982 128 20435
rect 116 0 128 11968
rect 139 10806 151 20411
rect 139 0 151 10792
rect 162 9630 174 20387
rect 162 0 174 9616
rect 185 8454 197 20363
rect 185 0 197 8440
rect 208 7278 220 20339
rect 208 0 220 7264
rect 231 6102 243 20315
rect 231 0 243 6088
rect 254 4926 266 20291
rect 254 0 266 4912
rect 277 3750 289 20267
rect 277 0 289 3736
rect 300 2574 312 20243
rect 300 0 312 2560
rect 323 1398 335 20219
rect 323 0 335 1384
rect 346 222 358 20195
rect 370 20186 570 20572
rect 586 20186 598 20572
rect 610 20186 622 20572
rect 634 20186 646 20572
rect 658 20186 670 20572
rect 4138 20186 4150 20572
rect 4162 20186 4174 20435
rect 4210 20186 4222 20363
rect 4378 20186 4390 20572
rect 4594 20186 4606 20411
rect 4642 20186 4654 20339
rect 4978 20186 4990 20387
rect 5026 20186 5038 20315
rect 5338 20186 5350 20572
rect 5530 20186 5542 20572
rect 6564 20186 6576 20572
rect 7118 20186 7130 20243
rect 7142 20186 7154 20267
rect 7166 20186 7178 20291
rect 14555 20186 14567 20572
rect 14579 20186 14591 20556
rect 14771 20186 14783 20531
rect 14819 20186 14831 20572
rect 14963 20186 14975 20507
rect 15155 20186 15167 20483
rect 15347 20186 15359 20459
rect 15539 20186 15551 20572
rect 17338 20186 17350 20572
rect 17530 20186 17542 20572
rect 17602 20186 17614 20572
rect 17698 20186 17710 20572
rect 22354 20186 22366 20267
rect 22546 20186 22558 20242
rect 22666 20186 22678 20219
rect 22786 20186 22798 20195
rect 25186 20186 25386 20572
rect 23626 18842 23638 18865
rect 3082 18665 3094 18735
rect 23626 17666 23638 17800
rect 3082 17489 3094 17559
rect 23626 16490 23638 16624
rect 3082 16313 3094 16383
rect 23626 15314 23638 15448
rect 3082 15137 3094 15207
rect 23626 14138 23638 14272
rect 3082 13961 3094 14031
rect 23626 12962 23638 13096
rect 3082 12785 3094 12855
rect 23626 11786 23638 11920
rect 3082 11609 3094 11679
rect 23626 10610 23638 10744
rect 3082 10433 3094 10503
rect 23626 9434 23638 9568
rect 3082 9257 3094 9327
rect 23626 8258 23638 8392
rect 3082 8081 3094 8151
rect 23626 7082 23638 7216
rect 3082 6905 3094 6975
rect 23626 5906 23638 6040
rect 3082 5729 3094 5799
rect 23626 4730 23638 4864
rect 3082 4553 3094 4623
rect 23626 3554 23638 3688
rect 3082 3377 3094 3447
rect 23626 2378 23638 2512
rect 3082 2201 3094 2271
rect 23626 1202 23638 1336
rect 3082 1025 3094 1095
rect 346 0 358 208
rect 23626 49 23638 160
rect 370 20 570 49
rect 370 6 556 20
rect 370 0 570 6
rect 586 0 598 49
rect 610 0 622 49
rect 634 0 646 49
rect 658 0 670 49
rect 1930 0 1942 49
rect 2122 0 2134 49
rect 2914 0 2926 49
rect 3322 19 3334 49
rect 3466 0 3478 49
rect 3682 0 3694 49
rect 4426 0 4438 49
rect 4594 0 4606 49
rect 4978 0 4990 49
rect 5170 0 5182 49
rect 5386 0 5398 49
rect 6130 0 6142 49
rect 6298 0 6310 49
rect 15706 0 15718 49
rect 15898 0 15910 49
rect 16138 0 16150 49
rect 16786 43 16798 49
rect 16978 43 16990 49
rect 16786 31 16990 43
rect 17266 41 17278 49
rect 19930 41 19942 49
rect 19978 41 19990 49
rect 20026 41 20038 49
rect 20074 41 20086 49
rect 20122 41 20134 49
rect 20170 41 20182 49
rect 20218 41 20230 49
rect 20266 41 20278 49
rect 20578 41 20590 49
rect 20626 41 20638 49
rect 20674 41 20686 49
rect 20722 41 20734 49
rect 21034 41 21046 49
rect 21082 41 21094 49
rect 21466 41 21478 49
rect 23842 0 23854 49
rect 24586 0 24598 49
rect 24730 0 24742 49
rect 24778 0 24790 49
rect 24826 0 24838 49
rect 24874 0 24886 49
rect 24946 0 24958 49
rect 25186 41 25386 49
rect 25200 27 25386 41
rect 25186 0 25386 27
use slice17 slice17_0
timestamp 1395569125
transform 1 0 370 0 1 18865
box 0 0 25016 1321
use leftbuf_slice leftbuf_slice_0
array 0 0 1685 0 15 1176
timestamp 1395689796
transform 1 0 365 0 1 49
box 0 0 1685 1176
use IrAA IrAA_0
array 0 0 1008 0 7 1176
timestamp 1395689161
transform 1 0 2050 0 1 9568
box 0 -111 1008 1065
use tielow tielow_0
timestamp 1386086605
transform 1 0 3058 0 1 17866
box 0 0 48 799
use tielow tielow_1
timestamp 1386086605
transform 1 0 3058 0 1 16690
box 0 0 48 799
use tielow tielow_2
timestamp 1386086605
transform 1 0 3058 0 1 15514
box 0 0 48 799
use tielow tielow_3
timestamp 1386086605
transform 1 0 3058 0 1 14338
box 0 0 48 799
use tielow tielow_4
timestamp 1386086605
transform 1 0 3058 0 1 13162
box 0 0 48 799
use tielow tielow_5
timestamp 1386086605
transform 1 0 3058 0 1 11986
box 0 0 48 799
use tielow tielow_6
timestamp 1386086605
transform 1 0 3058 0 1 10810
box 0 0 48 799
use tielow tielow_7
timestamp 1386086605
transform 1 0 3058 0 1 9634
box 0 0 48 799
use IrBA IrBA_0
array 0 0 1008 0 2 1176
timestamp 1395689161
transform 1 0 2050 0 1 6040
box 0 -111 1008 1065
use tielow tielow_8
timestamp 1386086605
transform 1 0 3058 0 1 8458
box 0 0 48 799
use tielow tielow_9
timestamp 1386086605
transform 1 0 3058 0 1 7282
box 0 0 48 799
use tielow tielow_10
timestamp 1386086605
transform 1 0 3058 0 1 6106
box 0 0 48 799
use IrBB IrBB_0
array 0 0 1008 0 4 1176
timestamp 1395689161
transform 1 0 2050 0 1 161
box 0 -112 1008 1064
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 3058 0 1 4930
box 0 0 48 799
use tielow tielow_12
timestamp 1386086605
transform 1 0 3058 0 1 3754
box 0 0 48 799
use tielow tielow_13
timestamp 1386086605
transform 1 0 3058 0 1 2578
box 0 0 48 799
use tielow tielow_14
timestamp 1386086605
transform 1 0 3058 0 1 1402
box 0 0 48 799
use tielow tielow_15
timestamp 1386086605
transform 1 0 3058 0 1 226
box 0 0 48 799
use Datapath_slice Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1395690245
transform 1 0 3106 0 1 49
box 0 0 20472 1176
use LLIcell_U LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1394841956
transform 1 0 23578 0 1 9568
box 0 0 192 1042
use LLIcell_L LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23578 0 1 160
box 0 0 192 1042
use Datapath_end_high Datapath_end_high_0
array 0 0 1621 0 11 1176
timestamp 1395689161
transform 1 0 23770 0 1 4753
box 0 0 1621 1176
use Datapath_end_low Datapath_end_low_0
array 0 0 1616 0 3 1176
timestamp 1395689161
transform 1 0 23770 0 1 49
box 0 0 1621 1176
<< labels >>
rlabel metal1 23674 1214 23674 1214 1 Aluout[0]
rlabel metal2 6 20260 6 20260 1 Ir[15]
rlabel metal2 30 20259 30 20259 1 Ir[14]
rlabel metal2 53 20259 53 20259 1 Ir[13]
rlabel metal2 76 20260 76 20260 1 Ir[12]
rlabel metal2 99 20260 99 20260 1 Ir[11]
rlabel metal2 122 20259 122 20259 1 Ir[10]
rlabel metal2 145 20260 145 20260 1 Ir[9]
rlabel metal2 168 20260 168 20260 1 Ir[8]
rlabel metal2 191 20262 191 20262 1 Ir[7]
rlabel metal2 214 20263 214 20263 1 Ir[6]
rlabel metal2 237 20264 237 20264 1 Ir[5]
rlabel metal2 260 20265 260 20265 1 Ir[4]
rlabel metal2 283 20264 283 20264 1 Ir[3]
rlabel metal2 22792 20190 22792 20190 1 Ir[0]
rlabel metal2 22671 20212 22671 20212 1 Ir[1]
rlabel metal2 22551 20237 22551 20237 1 Ir[2]
rlabel metal2 22360 20262 22360 20262 1 Ir[3]
rlabel metal2 14968 20501 14968 20501 1 Ir[13]
rlabel metal2 15161 20477 15161 20477 1 Ir[12]
rlabel metal2 15353 20452 15353 20452 1 Ir[11]
rlabel metal2 14775 20524 14775 20524 1 Ir[14]
rlabel metal2 14584 20549 14584 20549 1 Ir[15]
rlabel metal2 7122 20235 7122 20235 1 Ir[2]
rlabel metal2 7148 20259 7148 20259 1 Ir[3]
rlabel metal2 7171 20283 7171 20283 1 Ir[4]
rlabel metal2 4216 20355 4216 20355 1 Ir[7]
rlabel metal2 4167 20428 4167 20428 1 Ir[10]
rlabel metal2 4648 20332 4648 20332 1 Ir[6]
rlabel metal2 4599 20403 4599 20403 1 Ir[9]
rlabel metal2 4983 20380 4983 20380 1 Ir[8]
rlabel metal2 5033 20309 5033 20309 1 Ir[5]
rlabel metal2 6564 20572 6576 20572 5 RegWe
rlabel metal2 586 20572 598 20572 5 SDO
rlabel metal2 370 20572 570 20572 5 Vdd!
rlabel metal2 658 20572 670 20572 1 nReset
rlabel metal2 634 20572 646 20572 1 Clock
rlabel metal2 610 20572 622 20572 1 Test
rlabel metal2 17698 20572 17710 20572 5 Flags[0]
rlabel metal2 17602 20572 17614 20572 5 Flags[3]
rlabel metal2 17530 20572 17542 20572 5 Flags[1]
rlabel metal2 17338 20572 17350 20572 5 Flags[2]
rlabel metal2 14819 20572 14831 20572 5 AluOR[0]
rlabel metal2 14555 20572 14567 20572 5 AluOR[1]
rlabel metal2 15539 20572 15551 20572 5 CFlag
rlabel metal2 4138 20572 4150 20572 5 Rs1Sel[0]
rlabel metal2 4378 20572 4390 20572 5 Rs1Sel[1]
rlabel metal2 5338 20572 5350 20572 5 RwSel[0]
rlabel metal2 5530 20572 5542 20572 5 RwSel[1]
rlabel metal2 3466 0 3478 0 1 LrSel
rlabel metal2 3682 0 3694 0 1 LrWe
rlabel metal2 4426 0 4438 0 1 LrEn
rlabel metal2 4594 0 4606 0 1 PcSel[0]
rlabel metal2 4978 0 4990 0 1 PcSel[1]
rlabel metal2 23842 0 23854 0 1 AluWe
rlabel metal2 24586 0 24598 0 1 AluEn
rlabel metal2 370 0 570 0 1 Vdd!
rlabel metal2 586 0 598 0 1 SDI
rlabel metal2 610 0 622 0 1 Test
rlabel metal2 634 0 646 0 1 Clock
rlabel metal2 658 0 670 0 1 nReset
rlabel metal2 2914 0 2926 0 1 ImmSel
rlabel metal2 2122 0 2134 0 1 IrWe
rlabel metal2 1930 0 1942 0 1 MemEn
rlabel metal2 5386 0 5398 0 1 PcWe
rlabel metal2 5170 0 5182 0 1 PcSel[2]
rlabel metal2 6130 0 6142 0 1 PcEn
rlabel metal2 6298 0 6310 0 1 WdSel
rlabel metal2 15706 0 15718 0 1 Op1Sel
rlabel metal2 15898 0 15910 0 1 Op2Sel[0]
rlabel metal2 16138 0 16150 0 1 Op2Sel[1]
rlabel metal2 25186 0 25386 0 1 GND!
rlabel metal2 25186 20572 25386 20572 1 GND!
rlabel metal2 24946 0 24958 0 1 StatusRegEn
rlabel metal2 24730 0 24742 0 1 StatusReg[3]
rlabel metal2 24778 0 24790 0 1 StatusReg[2]
rlabel metal2 24826 0 24838 0 1 StatusReg[1]
rlabel metal2 24874 0 24886 0 1 StatusReg[0]
rlabel metal1 25408 78 25408 88 7 DataIn[0]
rlabel metal1 25408 1254 25408 1264 7 DataIn[1]
rlabel metal1 25408 2430 25408 2440 7 DataIn[2]
rlabel metal1 25408 3606 25408 3616 7 DataIn[3]
rlabel metal1 25408 4782 25408 4792 7 DataIn[4]
rlabel metal1 25408 5958 25408 5968 7 DataIn[5]
rlabel metal1 25408 7134 25408 7144 7 DataIn[6]
rlabel metal1 25408 8310 25408 8320 7 DataIn[7]
rlabel metal1 25408 9486 25408 9496 7 DataIn[8]
rlabel metal1 25408 10662 25408 10672 7 DataIn[9]
rlabel metal1 25408 11838 25408 11848 7 DataIn[10]
rlabel metal1 25408 13014 25408 13024 7 DataIn[11]
rlabel metal1 25408 14190 25408 14200 7 DataIn[12]
rlabel metal1 25408 15366 25408 15376 7 DataIn[13]
rlabel metal1 25408 16542 25408 16552 7 DataIn[14]
rlabel metal1 25408 17718 25408 17728 7 DataIn[15]
rlabel metal1 25408 144 25408 154 7 DataOut[0]
rlabel metal1 25408 1320 25408 1330 7 DataOut[1]
rlabel metal1 25408 2496 25408 2506 7 DataOut[2]
rlabel metal1 25408 3672 25408 3682 7 DataOut[3]
rlabel metal1 25408 4848 25408 4858 7 DataOut[4]
rlabel metal1 25408 6024 25408 6034 7 DataOut[5]
rlabel metal1 25408 7200 25408 7210 7 DataOut[6]
rlabel metal1 25408 8376 25408 8386 7 DataOut[7]
rlabel metal1 25408 9552 25408 9562 7 DataOut[8]
rlabel metal1 25408 10728 25408 10738 7 DataOut[9]
rlabel metal1 25408 11904 25408 11914 7 DataOut[10]
rlabel metal1 25408 13080 25408 13090 7 DataOut[11]
rlabel metal1 25408 14256 25408 14266 7 DataOut[12]
rlabel metal1 25408 15432 25408 15442 7 DataOut[13]
rlabel metal1 25408 16608 25408 16618 7 DataOut[14]
rlabel metal1 25408 17784 25408 17794 7 DataOut[15]
rlabel metal2 346 0 358 0 1 Ir[0]
rlabel metal2 323 0 335 0 1 Ir[1]
rlabel metal2 300 0 312 0 1 Ir[2]
rlabel metal2 277 0 289 0 1 Ir[3]
rlabel metal2 254 0 266 0 1 Ir[4]
rlabel metal2 231 0 243 0 1 Ir[5]
rlabel metal2 208 0 220 0 1 Ir[6]
rlabel metal2 185 0 197 0 1 Ir[7]
rlabel metal2 162 0 174 0 1 Ir[8]
rlabel metal2 139 0 151 0 1 Ir[9]
rlabel metal2 116 0 128 0 1 Ir[10]
rlabel metal2 93 0 105 0 1 Ir[11]
rlabel metal2 70 0 82 0 1 Ir[12]
rlabel metal2 47 0 59 0 1 Ir[13]
rlabel metal2 24 0 36 0 1 Ir[14]
rlabel metal2 1 0 13 0 1 Ir[15]
<< end >>
