magic
tech c035u
timestamp 1394990419
<< error_s >>
rect 492 55899 496 55909
rect 732 55899 736 55909
rect 972 55899 976 55909
rect 1212 55899 1216 55909
rect 1452 55899 1456 55909
rect 1692 55899 1696 55909
rect 1932 55899 1936 55909
rect 2172 55899 2176 55909
rect 2412 55899 2416 55909
rect 2652 55899 2656 55909
rect 2892 55899 2896 55909
rect 3132 55899 3136 55909
rect 3372 55899 3376 55909
rect 3612 55899 3616 55909
rect 3852 55899 3856 55909
rect 4092 55899 4096 55909
rect 4332 55899 4336 55909
rect 4572 55899 4576 55909
rect 4812 55899 4816 55909
rect 7212 55899 7216 55909
rect 10092 55899 10096 55909
rect 10332 55899 10336 55909
rect 10572 55899 10576 55909
rect 10812 55899 10816 55909
rect 11052 55899 11056 55909
rect 11292 55899 11296 55909
rect 11532 55899 11536 55909
rect 11772 55899 11776 55909
rect 12012 55899 12016 55909
rect 12252 55899 12256 55909
rect 12492 55899 12496 55909
rect 12732 55899 12736 55909
rect 12972 55899 12976 55909
rect 13212 55899 13216 55909
rect 13452 55899 13456 55909
rect 13692 55899 13696 55909
rect 13932 55899 13936 55909
rect 14172 55899 14176 55909
rect 14412 55899 14416 55909
rect 14652 55899 14656 55909
rect 14892 55899 14896 55909
rect 15132 55899 15136 55909
rect 15372 55899 15376 55909
rect 15612 55899 15616 55909
rect 15852 55899 15856 55909
rect 21800 55899 21808 55909
rect 502 55870 506 55899
rect 742 55870 746 55899
rect 982 55870 986 55899
rect 1222 55870 1226 55899
rect 1462 55870 1466 55899
rect 1702 55870 1706 55899
rect 1942 55870 1946 55899
rect 2182 55870 2186 55899
rect 2422 55870 2426 55899
rect 2662 55870 2666 55899
rect 2902 55870 2906 55899
rect 3142 55870 3146 55899
rect 3382 55870 3386 55899
rect 3622 55870 3626 55899
rect 3862 55870 3866 55899
rect 4102 55870 4106 55899
rect 4342 55870 4346 55899
rect 4582 55870 4586 55899
rect 4822 55870 4826 55899
rect 7222 55870 7226 55899
rect 10102 55870 10106 55899
rect 10342 55870 10346 55899
rect 10582 55870 10586 55899
rect 10822 55870 10826 55899
rect 11062 55870 11066 55899
rect 11302 55870 11306 55899
rect 11542 55870 11546 55899
rect 11782 55870 11786 55899
rect 12022 55870 12026 55899
rect 12262 55870 12266 55899
rect 12502 55870 12506 55899
rect 12742 55870 12746 55899
rect 12982 55870 12986 55899
rect 13222 55870 13226 55899
rect 13462 55870 13466 55899
rect 13702 55870 13706 55899
rect 13942 55870 13946 55899
rect 14182 55870 14186 55899
rect 14422 55870 14426 55899
rect 14662 55870 14666 55899
rect 14902 55870 14906 55899
rect 15142 55870 15146 55899
rect 15382 55870 15386 55899
rect 15622 55870 15626 55899
rect 15862 55870 15866 55899
rect 21810 55870 21818 55899
rect -2371 48014 -2366 49150
rect -2348 48014 -2343 49150
rect -2325 49126 -2320 49150
rect -2325 49118 -2317 49126
rect -2325 49098 -2320 49118
rect -2317 49110 -2309 49118
rect -2325 49082 -2317 49098
rect -2325 49066 -2320 49082
rect -2309 49070 -2301 49082
rect -2317 49066 -2309 49070
rect -2103 49066 -2096 49068
rect -2083 49066 -2053 49068
rect -2325 49054 -2317 49066
rect -2103 49057 -2053 49066
rect -2018 49064 -2017 49070
rect -2003 49064 -2002 49066
rect -2026 49060 -2017 49064
rect -2325 49038 -2320 49054
rect -2309 49042 -2301 49054
rect -2017 49050 -2012 49060
rect -2317 49038 -2309 49042
rect -2325 49026 -2317 49038
rect -2325 49006 -2320 49026
rect -2325 48998 -2317 49006
rect -2325 48978 -2320 48998
rect -2317 48990 -2309 48998
rect -2325 48962 -2317 48978
rect -2325 48946 -2320 48962
rect -2309 48950 -2301 48962
rect -2317 48946 -2309 48950
rect -2103 48946 -2096 48948
rect -2083 48946 -2053 48948
rect -2325 48934 -2317 48946
rect -2103 48937 -2053 48946
rect -2018 48944 -2017 48950
rect -2003 48944 -2002 48946
rect -2026 48940 -2017 48944
rect -2325 48918 -2320 48934
rect -2309 48922 -2301 48934
rect -2017 48930 -2012 48940
rect -2317 48918 -2309 48922
rect -2325 48906 -2317 48918
rect -2325 48886 -2320 48906
rect -2325 48878 -2317 48886
rect -2325 48858 -2320 48878
rect -2317 48870 -2309 48878
rect -2325 48842 -2317 48858
rect -2325 48826 -2320 48842
rect -2309 48830 -2301 48842
rect -2317 48826 -2309 48830
rect -2103 48826 -2096 48828
rect -2083 48826 -2053 48828
rect -2325 48814 -2317 48826
rect -2103 48817 -2053 48826
rect -2018 48824 -2017 48830
rect -2003 48824 -2002 48826
rect -2026 48820 -2017 48824
rect -2325 48798 -2320 48814
rect -2309 48802 -2301 48814
rect -2017 48810 -2012 48820
rect -2317 48798 -2309 48802
rect -2325 48786 -2317 48798
rect -2325 48766 -2320 48786
rect -2325 48758 -2317 48766
rect -2325 48738 -2320 48758
rect -2317 48750 -2309 48758
rect -2325 48722 -2317 48738
rect -2325 48706 -2320 48722
rect -2309 48710 -2301 48722
rect -2317 48706 -2309 48710
rect -2103 48706 -2096 48708
rect -2083 48706 -2053 48708
rect -2325 48694 -2317 48706
rect -2103 48697 -2053 48706
rect -2018 48704 -2017 48710
rect -2003 48704 -2002 48706
rect -2026 48700 -2017 48704
rect -2325 48678 -2320 48694
rect -2309 48682 -2301 48694
rect -2017 48690 -2012 48700
rect -2317 48678 -2309 48682
rect -2325 48666 -2317 48678
rect -2325 48646 -2320 48666
rect -2325 48638 -2317 48646
rect -2325 48618 -2320 48638
rect -2317 48630 -2309 48638
rect -2325 48602 -2317 48618
rect -2325 48586 -2320 48602
rect -2309 48590 -2301 48602
rect -2317 48586 -2309 48590
rect -2103 48586 -2096 48588
rect -2083 48586 -2053 48588
rect -2325 48574 -2317 48586
rect -2103 48577 -2053 48586
rect -2018 48584 -2017 48590
rect -2003 48584 -2002 48586
rect -2026 48580 -2017 48584
rect -2325 48558 -2320 48574
rect -2309 48562 -2301 48574
rect -2017 48570 -2012 48580
rect -2317 48558 -2309 48562
rect -2325 48546 -2317 48558
rect -2325 48526 -2320 48546
rect -2325 48518 -2317 48526
rect -2325 48498 -2320 48518
rect -2317 48510 -2309 48518
rect -2325 48482 -2317 48498
rect -2325 48466 -2320 48482
rect -2309 48470 -2301 48482
rect -2317 48466 -2309 48470
rect -2103 48466 -2096 48468
rect -2083 48466 -2053 48468
rect -2325 48454 -2317 48466
rect -2103 48457 -2053 48466
rect -2018 48464 -2017 48470
rect -2003 48464 -2002 48466
rect -2026 48460 -2017 48464
rect -2325 48438 -2320 48454
rect -2309 48442 -2301 48454
rect -2017 48450 -2012 48460
rect -2317 48438 -2309 48442
rect -2325 48426 -2317 48438
rect -2325 48406 -2320 48426
rect -2325 48398 -2317 48406
rect -2325 48378 -2320 48398
rect -2317 48390 -2309 48398
rect -2325 48362 -2317 48378
rect -2325 48346 -2320 48362
rect -2309 48350 -2301 48362
rect -2317 48346 -2309 48350
rect -2103 48346 -2096 48348
rect -2083 48346 -2053 48348
rect -2325 48334 -2317 48346
rect -2103 48337 -2053 48346
rect -2018 48344 -2017 48350
rect -2003 48344 -2002 48346
rect -2026 48340 -2017 48344
rect -2325 48318 -2320 48334
rect -2309 48322 -2301 48334
rect -2017 48330 -2012 48340
rect -2317 48318 -2309 48322
rect -2325 48306 -2317 48318
rect -2325 48286 -2320 48306
rect -2325 48278 -2317 48286
rect -2325 48258 -2320 48278
rect -2317 48270 -2309 48278
rect -2325 48242 -2317 48258
rect -2325 48226 -2320 48242
rect -2309 48230 -2301 48242
rect -2317 48226 -2309 48230
rect -2103 48226 -2096 48228
rect -2083 48226 -2053 48228
rect -2325 48214 -2317 48226
rect -2103 48217 -2053 48226
rect -2018 48224 -2017 48230
rect -2003 48224 -2002 48226
rect -2026 48220 -2017 48224
rect -2325 48198 -2320 48214
rect -2309 48202 -2301 48214
rect -2017 48210 -2012 48220
rect -2317 48198 -2309 48202
rect -2325 48186 -2317 48198
rect -2325 48166 -2320 48186
rect -2325 48158 -2317 48166
rect -2325 48138 -2320 48158
rect -2317 48150 -2309 48158
rect -2325 48122 -2317 48138
rect -2325 48106 -2320 48122
rect -2309 48110 -2301 48122
rect -2317 48106 -2309 48110
rect -2103 48106 -2096 48108
rect -2083 48106 -2053 48108
rect -2325 48094 -2317 48106
rect -2103 48097 -2053 48106
rect -2018 48104 -2017 48110
rect -2003 48104 -2002 48106
rect -2026 48100 -2017 48104
rect -2325 48078 -2320 48094
rect -2309 48082 -2301 48094
rect -2017 48090 -2012 48100
rect -2317 48078 -2309 48082
rect -2325 48066 -2317 48078
rect -2325 48046 -2320 48066
rect -2325 48038 -2317 48046
rect -2325 48018 -2320 48038
rect -2317 48030 -2309 48038
rect -2325 48014 -2317 48018
rect -2000 48014 -1992 49140
rect -1671 49118 -1663 49126
rect -1663 49110 -1655 49118
rect -1671 49082 -1663 49098
rect -1655 49070 -1647 49082
rect -1972 49066 -1924 49068
rect -1663 49066 -1655 49070
rect -1972 49057 -1922 49066
rect -1671 49054 -1663 49066
rect -1655 49042 -1647 49054
rect -1663 49038 -1655 49042
rect -1671 49026 -1663 49038
rect -1671 48998 -1663 49006
rect -1663 48990 -1655 48998
rect -1671 48962 -1663 48978
rect -1655 48950 -1647 48962
rect -1972 48946 -1924 48948
rect -1663 48946 -1655 48950
rect -1972 48937 -1922 48946
rect -1671 48934 -1663 48946
rect -1655 48922 -1647 48934
rect -1663 48918 -1655 48922
rect -1671 48906 -1663 48918
rect -1671 48878 -1663 48886
rect -1663 48870 -1655 48878
rect -1671 48842 -1663 48858
rect -1655 48830 -1647 48842
rect -1972 48826 -1924 48828
rect -1663 48826 -1655 48830
rect -1972 48817 -1922 48826
rect -1671 48814 -1663 48826
rect -1655 48802 -1647 48814
rect -1663 48798 -1655 48802
rect -1671 48786 -1663 48798
rect -1671 48758 -1663 48766
rect -1663 48750 -1655 48758
rect -1671 48722 -1663 48738
rect -1655 48710 -1647 48722
rect -1972 48706 -1924 48708
rect -1663 48706 -1655 48710
rect -1972 48697 -1922 48706
rect -1671 48694 -1663 48706
rect -1655 48682 -1647 48694
rect -1663 48678 -1655 48682
rect -1671 48666 -1663 48678
rect -1671 48638 -1663 48646
rect -1663 48630 -1655 48638
rect -1671 48602 -1663 48618
rect -1655 48590 -1647 48602
rect -1972 48586 -1924 48588
rect -1663 48586 -1655 48590
rect -1972 48577 -1922 48586
rect -1671 48574 -1663 48586
rect -1655 48562 -1647 48574
rect -1663 48558 -1655 48562
rect -1671 48546 -1663 48558
rect -1671 48518 -1663 48526
rect -1663 48510 -1655 48518
rect -1671 48482 -1663 48498
rect -1655 48470 -1647 48482
rect -1972 48466 -1924 48468
rect -1663 48466 -1655 48470
rect -1972 48457 -1922 48466
rect -1671 48454 -1663 48466
rect -1655 48442 -1647 48454
rect -1663 48438 -1655 48442
rect -1671 48426 -1663 48438
rect -1671 48398 -1663 48406
rect -1663 48390 -1655 48398
rect -1671 48362 -1663 48378
rect -1655 48350 -1647 48362
rect -1972 48346 -1924 48348
rect -1663 48346 -1655 48350
rect -1972 48337 -1922 48346
rect -1671 48334 -1663 48346
rect -1655 48322 -1647 48334
rect -1663 48318 -1655 48322
rect -1671 48306 -1663 48318
rect -1671 48278 -1663 48286
rect -1663 48270 -1655 48278
rect -1671 48242 -1663 48258
rect -1655 48230 -1647 48242
rect -1972 48226 -1924 48228
rect -1663 48226 -1655 48230
rect -1972 48217 -1922 48226
rect -1671 48214 -1663 48226
rect -1655 48202 -1647 48214
rect -1663 48198 -1655 48202
rect -1671 48186 -1663 48198
rect -1671 48158 -1663 48166
rect -1663 48150 -1655 48158
rect -1671 48122 -1663 48138
rect -1655 48110 -1647 48122
rect -1972 48106 -1924 48108
rect -1663 48106 -1655 48110
rect -1972 48097 -1922 48106
rect -1671 48094 -1663 48106
rect -1655 48082 -1647 48094
rect -1663 48078 -1655 48082
rect -1671 48066 -1663 48078
rect -1671 48038 -1663 48046
rect -1663 48030 -1655 48038
rect -1671 48014 -1663 48018
rect -1642 48014 -1637 49150
rect -1619 48014 -1614 49150
rect 499 49133 504 49143
rect 739 49133 744 49143
rect 509 49119 514 49133
rect 749 49119 754 49133
rect -1554 49102 -1547 49115
rect -1554 49091 -1547 49092
rect -1530 49078 -1526 49112
rect -1554 49054 -1547 49067
rect -1554 49043 -1547 49044
rect -1530 49043 -1523 49067
rect -1517 49061 -1512 49071
rect -1507 49047 -1502 49061
rect -1493 49057 -1485 49061
rect -1499 49047 -1493 49057
rect -1565 48974 -1531 48975
rect -1530 48974 -1526 49043
rect -1506 48974 -1502 49047
rect 486 49043 493 49067
rect 726 49043 733 49067
rect 499 49013 504 49023
rect 739 49013 744 49023
rect 1219 49013 1224 49023
rect 1459 49013 1464 49023
rect 1699 49013 1704 49023
rect 1939 49013 1944 49023
rect 2179 49013 2184 49023
rect 2419 49013 2424 49023
rect 2659 49013 2664 49023
rect 2899 49013 2904 49023
rect 3139 49013 3144 49023
rect 3379 49013 3384 49023
rect 509 48999 514 49013
rect 749 48999 754 49013
rect 1229 48999 1234 49013
rect 1469 48999 1474 49013
rect 1709 48999 1714 49013
rect 1949 48999 1954 49013
rect 2189 48999 2194 49013
rect 2429 48999 2434 49013
rect 2669 48999 2674 49013
rect 2909 48999 2914 49013
rect 3149 48999 3154 49013
rect 3389 48999 3394 49013
rect -1493 48974 -1485 48975
rect -1565 48972 -1485 48974
rect -1530 48899 -1526 48972
rect -1506 48927 -1502 48972
rect -1499 48971 -1485 48972
rect -1493 48965 -1488 48971
rect -1483 48951 -1478 48965
rect -1517 48926 -1483 48927
rect -1482 48926 -1478 48951
rect -1469 48926 -1435 48927
rect -1517 48924 -1435 48926
rect -1517 48917 -1512 48924
rect -1506 48917 -1502 48924
rect -1507 48903 -1502 48917
rect -1530 48875 -1523 48899
rect -1517 48893 -1512 48903
rect -1507 48879 -1502 48893
rect -1554 48862 -1547 48875
rect -1554 48851 -1547 48852
rect -1541 48845 -1536 48855
rect -1530 48845 -1526 48872
rect -1531 48831 -1526 48845
rect -1541 48821 -1536 48831
rect -1531 48807 -1526 48821
rect -1565 48806 -1531 48807
rect -1530 48806 -1526 48807
rect -1506 48806 -1502 48879
rect -1482 48851 -1478 48924
rect -1475 48923 -1461 48924
rect 486 48923 493 48947
rect 726 48923 733 48947
rect 1206 48923 1213 48947
rect 1446 48923 1453 48947
rect 1686 48923 1693 48947
rect 1926 48923 1933 48947
rect 2166 48923 2173 48947
rect 2406 48923 2413 48947
rect 2646 48923 2653 48947
rect 2886 48923 2893 48947
rect 3126 48923 3133 48947
rect 3366 48923 3373 48947
rect -1458 48875 -1451 48899
rect 499 48893 504 48903
rect 739 48893 744 48903
rect 1219 48893 1224 48903
rect 1459 48893 1464 48903
rect 1699 48893 1704 48903
rect 1939 48893 1944 48903
rect 509 48879 514 48893
rect 749 48879 754 48893
rect 1229 48879 1234 48893
rect 1469 48879 1474 48893
rect 1709 48879 1714 48893
rect 1949 48879 1954 48893
rect -1482 48806 -1475 48851
rect -1458 48806 -1454 48875
rect -1435 48831 -1427 48845
rect -1434 48827 -1427 48831
rect -1434 48806 -1430 48827
rect -1421 48806 -1387 48807
rect -1565 48804 -1387 48806
rect -1530 48731 -1526 48804
rect -1506 48779 -1502 48804
rect -1499 48803 -1485 48804
rect -1482 48803 -1475 48804
rect -1506 48731 -1499 48779
rect -1530 48710 -1523 48731
rect -1506 48710 -1502 48731
rect -1482 48710 -1478 48803
rect -1469 48725 -1464 48735
rect -1458 48725 -1454 48804
rect -1459 48711 -1454 48725
rect -1469 48710 -1435 48711
rect -1547 48708 -1435 48710
rect -1547 48707 -1533 48708
rect -1554 48694 -1547 48707
rect -1530 48687 -1523 48708
rect -1541 48686 -1507 48687
rect -1506 48686 -1502 48708
rect -1482 48686 -1478 48708
rect -1469 48701 -1464 48708
rect -1459 48687 -1454 48701
rect -1458 48686 -1454 48687
rect -1434 48686 -1430 48804
rect -1427 48803 -1413 48804
rect 486 48803 493 48827
rect 726 48803 733 48827
rect 1206 48803 1213 48827
rect 1446 48803 1453 48827
rect 1686 48803 1693 48827
rect 1926 48803 1933 48827
rect -1410 48755 -1403 48779
rect 499 48773 504 48783
rect 739 48773 744 48783
rect 509 48759 514 48773
rect 749 48759 754 48773
rect -1410 48686 -1406 48755
rect -1387 48711 -1379 48725
rect -1386 48707 -1379 48711
rect -1386 48686 -1382 48707
rect -1373 48686 -1339 48687
rect -1541 48684 -1339 48686
rect -1554 48683 -1547 48684
rect -1541 48683 -1533 48684
rect -1530 48683 -1523 48684
rect -1541 48677 -1536 48683
rect -1530 48677 -1526 48683
rect -1531 48663 -1526 48677
rect -1541 48653 -1536 48663
rect -1531 48639 -1526 48653
rect -1530 48014 -1526 48639
rect -1506 48611 -1502 48684
rect -1506 48590 -1499 48611
rect -1482 48590 -1478 48684
rect -1458 48590 -1454 48684
rect -1434 48659 -1430 48684
rect -1434 48611 -1427 48659
rect -1434 48590 -1430 48611
rect -1410 48590 -1406 48684
rect -1397 48605 -1392 48615
rect -1386 48605 -1382 48684
rect -1379 48683 -1365 48684
rect 486 48683 493 48707
rect 726 48683 733 48707
rect -1387 48591 -1382 48605
rect -1362 48635 -1355 48659
rect 499 48653 504 48663
rect 509 48639 514 48653
rect -1397 48590 -1363 48591
rect -1523 48588 -1363 48590
rect -1523 48587 -1509 48588
rect -1506 48567 -1499 48588
rect -1517 48566 -1483 48567
rect -1482 48566 -1478 48588
rect -1458 48566 -1454 48588
rect -1434 48566 -1430 48588
rect -1410 48566 -1406 48588
rect -1397 48581 -1392 48588
rect -1387 48567 -1382 48581
rect -1386 48566 -1382 48567
rect -1362 48566 -1358 48635
rect -1339 48591 -1331 48605
rect -1338 48587 -1331 48591
rect -1338 48566 -1334 48587
rect -1325 48566 -1291 48567
rect -1517 48564 -1291 48566
rect -1517 48563 -1509 48564
rect -1506 48563 -1499 48564
rect -1517 48557 -1512 48563
rect -1506 48557 -1502 48563
rect -1507 48543 -1502 48557
rect -1517 48533 -1512 48543
rect -1507 48519 -1502 48533
rect -1506 48207 -1502 48519
rect -1482 48491 -1478 48564
rect -1482 48470 -1475 48491
rect -1458 48470 -1454 48564
rect -1434 48470 -1430 48564
rect -1410 48495 -1406 48564
rect -1421 48494 -1387 48495
rect -1386 48494 -1382 48564
rect -1362 48539 -1358 48564
rect -1421 48492 -1365 48494
rect -1421 48485 -1416 48492
rect -1410 48485 -1406 48492
rect -1411 48471 -1406 48485
rect -1421 48470 -1387 48471
rect -1499 48468 -1387 48470
rect -1499 48467 -1485 48468
rect -1482 48443 -1475 48468
rect -1517 48206 -1483 48207
rect -1482 48206 -1478 48443
rect -1458 48206 -1454 48468
rect -1434 48206 -1430 48468
rect -1421 48461 -1416 48468
rect -1411 48447 -1406 48461
rect -1410 48206 -1406 48447
rect -1386 48419 -1382 48492
rect -1379 48491 -1365 48492
rect -1362 48491 -1355 48539
rect -1386 48371 -1379 48419
rect -1386 48206 -1382 48371
rect -1373 48365 -1368 48375
rect -1362 48365 -1358 48491
rect -1363 48351 -1358 48365
rect -1373 48341 -1368 48351
rect -1363 48327 -1358 48341
rect -1362 48206 -1358 48327
rect -1338 48299 -1334 48564
rect -1331 48563 -1317 48564
rect 486 48563 493 48587
rect -1314 48515 -1307 48539
rect -1338 48251 -1331 48299
rect -1338 48206 -1334 48251
rect -1314 48206 -1310 48515
rect -1291 48471 -1283 48485
rect -1290 48467 -1283 48471
rect -1290 48424 -1286 48467
rect -1280 48443 -1269 48444
rect -1301 48413 -1296 48423
rect -1291 48399 -1286 48413
rect -1277 48409 -1269 48413
rect -1283 48399 -1277 48409
rect -1290 48206 -1286 48399
rect -1266 48395 -1259 48419
rect -1266 48358 -1262 48395
rect -1243 48351 -1238 48365
rect -1266 48323 -1259 48347
rect -1266 48206 -1262 48323
rect -1242 48304 -1238 48351
rect -1232 48323 -1221 48324
rect -1253 48293 -1248 48303
rect -1243 48279 -1238 48293
rect -1229 48289 -1221 48293
rect -1235 48279 -1229 48289
rect -1253 48245 -1248 48255
rect -1242 48245 -1238 48279
rect -1243 48231 -1238 48245
rect -1218 48275 -1211 48299
rect 1699 48293 1704 48303
rect 1939 48293 1944 48303
rect 2419 48293 2424 48303
rect 2659 48293 2664 48303
rect 2899 48293 2904 48303
rect 3139 48293 3144 48303
rect 1709 48279 1714 48293
rect 1949 48279 1954 48293
rect 2429 48279 2434 48293
rect 2669 48279 2674 48293
rect 2909 48279 2914 48293
rect 3149 48279 3154 48293
rect -1218 48238 -1214 48275
rect -1195 48231 -1190 48245
rect -1253 48221 -1248 48231
rect -1234 48228 -1219 48231
rect -1243 48207 -1238 48221
rect -1229 48217 -1221 48221
rect -1235 48207 -1229 48217
rect -1242 48206 -1238 48207
rect -1218 48206 -1211 48227
rect -1194 48206 -1190 48231
rect -1181 48206 -1147 48207
rect -1517 48204 -1147 48206
rect -1517 48197 -1512 48204
rect -1506 48197 -1502 48204
rect -1507 48183 -1502 48197
rect -1517 48173 -1512 48183
rect -1507 48159 -1502 48173
rect -1506 48014 -1502 48159
rect -1482 48131 -1478 48204
rect -1482 48110 -1475 48131
rect -1458 48110 -1454 48204
rect -1434 48110 -1430 48204
rect -1410 48110 -1406 48204
rect -1386 48110 -1382 48204
rect -1362 48110 -1358 48204
rect -1338 48110 -1334 48204
rect -1314 48110 -1310 48204
rect -1290 48110 -1286 48204
rect -1266 48110 -1262 48204
rect -1242 48110 -1238 48204
rect -1235 48203 -1221 48204
rect -1218 48203 -1211 48204
rect -1218 48179 -1214 48203
rect -1218 48131 -1211 48179
rect -1218 48110 -1214 48131
rect -1205 48125 -1200 48135
rect -1194 48125 -1190 48204
rect -1187 48203 -1173 48204
rect 1686 48203 1693 48227
rect 1926 48203 1933 48227
rect 2406 48203 2413 48227
rect 2646 48203 2653 48227
rect 2886 48203 2893 48227
rect 3126 48203 3133 48227
rect -1195 48111 -1190 48125
rect -1170 48155 -1163 48179
rect 1699 48173 1704 48183
rect 1709 48159 1714 48173
rect -1205 48110 -1171 48111
rect -1499 48108 -1171 48110
rect -1499 48107 -1485 48108
rect -1482 48083 -1475 48108
rect -1482 48014 -1478 48083
rect -1458 48014 -1454 48108
rect -1434 48014 -1430 48108
rect -1410 48014 -1406 48108
rect -1397 48029 -1392 48039
rect -1386 48029 -1382 48108
rect -1387 48015 -1382 48029
rect -1362 48014 -1358 48108
rect -1338 48014 -1334 48108
rect -1314 48014 -1310 48108
rect -1290 48014 -1286 48108
rect -1266 48014 -1262 48108
rect -1242 48014 -1238 48108
rect -1218 48014 -1214 48108
rect -1205 48101 -1200 48108
rect -1195 48087 -1190 48101
rect -1205 48086 -1171 48087
rect -1170 48086 -1166 48155
rect -1147 48111 -1139 48125
rect -1146 48107 -1139 48111
rect -1146 48086 -1142 48107
rect -1133 48086 -1099 48087
rect -1205 48084 -1099 48086
rect -1205 48077 -1200 48084
rect -1194 48077 -1190 48084
rect -1195 48063 -1190 48077
rect -1205 48053 -1200 48063
rect -1170 48059 -1166 48084
rect -1195 48039 -1190 48053
rect -1181 48049 -1173 48053
rect -1187 48039 -1181 48049
rect -1194 48014 -1190 48039
rect -1170 48038 -1163 48059
rect -1146 48038 -1142 48084
rect -1139 48083 -1125 48084
rect 1686 48083 1693 48107
rect -1187 48036 -1125 48038
rect -1187 48035 -1173 48036
rect -2393 48012 -1969 48014
rect -1955 48012 -1173 48014
rect -2371 47966 -2366 48012
rect -2348 47966 -2343 48012
rect -2325 48002 -2317 48012
rect -2080 48010 -1969 48012
rect -2080 48004 -2053 48010
rect -2325 47986 -2320 48002
rect -2309 47990 -2301 48002
rect -2070 47995 -2040 48002
rect -2000 47994 -1992 48010
rect -1972 48006 -1969 48010
rect -1972 48004 -1955 48006
rect -1955 47994 -1850 48003
rect -1671 48002 -1663 48012
rect -2317 47986 -2309 47990
rect -2070 47987 -2053 47993
rect -2027 47992 -1992 47994
rect -1969 47992 -1955 47993
rect -2325 47974 -2317 47986
rect -2292 47977 -2053 47986
rect -2325 47966 -2320 47974
rect -2309 47966 -2301 47974
rect -2000 47966 -1992 47992
rect -1655 47990 -1647 48002
rect -1663 47986 -1655 47990
rect -1972 47978 -1924 47985
rect -1945 47977 -1929 47978
rect -1860 47977 -1680 47986
rect -1671 47974 -1663 47986
rect -1978 47966 -1942 47967
rect -1655 47966 -1647 47974
rect -1642 47966 -1637 48012
rect -1619 47966 -1614 48012
rect -1530 47966 -1526 48012
rect -1506 47966 -1502 48012
rect -1493 47981 -1488 47991
rect -1482 47981 -1478 48012
rect -1483 47967 -1478 47981
rect -1458 47966 -1454 48012
rect -1434 47966 -1430 48012
rect -1410 47966 -1406 48012
rect -1397 47966 -1363 47967
rect -2393 47964 -1363 47966
rect -2371 47870 -2366 47964
rect -2348 47870 -2343 47964
rect -2325 47958 -2320 47964
rect -2309 47962 -2301 47964
rect -2317 47958 -2309 47962
rect -2325 47946 -2317 47958
rect -2325 47926 -2320 47946
rect -2062 47926 -2032 47927
rect -2000 47926 -1992 47964
rect -1655 47962 -1647 47964
rect -1663 47958 -1655 47962
rect -1671 47946 -1663 47958
rect -1942 47928 -1937 47940
rect -1850 47937 -1822 47938
rect -1850 47933 -1802 47937
rect -2325 47918 -2317 47926
rect -2062 47924 -1961 47926
rect -2325 47898 -2320 47918
rect -2317 47910 -2309 47918
rect -2062 47911 -2040 47922
rect -2032 47917 -1961 47924
rect -1947 47918 -1942 47926
rect -1842 47924 -1794 47927
rect -2070 47906 -2022 47910
rect -2325 47884 -2317 47898
rect -2072 47890 -2032 47891
rect -2102 47884 -2032 47890
rect -2325 47870 -2320 47884
rect -2317 47882 -2309 47884
rect -2309 47870 -2301 47882
rect -2070 47875 -2062 47880
rect -2000 47870 -1992 47917
rect -1942 47916 -1937 47918
rect -1932 47908 -1927 47916
rect -1912 47913 -1896 47919
rect -1842 47911 -1802 47922
rect -1671 47918 -1663 47926
rect -1663 47910 -1655 47918
rect -1850 47906 -1680 47910
rect -1924 47892 -1921 47894
rect -1806 47884 -1680 47890
rect -1671 47884 -1663 47898
rect -1663 47882 -1655 47884
rect -1854 47875 -1806 47880
rect -1974 47870 -1964 47871
rect -1960 47870 -1944 47872
rect -1842 47870 -1806 47873
rect -1655 47870 -1647 47882
rect -1642 47870 -1637 47964
rect -1619 47870 -1614 47964
rect -1530 47870 -1526 47964
rect -1506 47870 -1502 47964
rect -1493 47933 -1488 47943
rect -1483 47919 -1478 47933
rect -1482 47870 -1478 47919
rect -1458 47915 -1454 47964
rect -1458 47894 -1451 47915
rect -1434 47894 -1430 47964
rect -1410 47894 -1406 47964
rect -1397 47957 -1392 47964
rect -1362 47963 -1358 48012
rect -1387 47943 -1382 47957
rect -1373 47953 -1365 47957
rect -1379 47943 -1373 47953
rect -1386 47894 -1382 47943
rect -1362 47939 -1355 47963
rect -1338 47894 -1334 48012
rect -1314 47894 -1310 48012
rect -1290 47894 -1286 48012
rect -1266 47894 -1262 48012
rect -1242 47894 -1238 48012
rect -1218 47919 -1214 48012
rect -1229 47918 -1195 47919
rect -1194 47918 -1190 48012
rect -1187 48011 -1173 48012
rect -1170 47990 -1163 48036
rect -1146 47990 -1142 48036
rect -1139 48035 -1125 48036
rect -1122 48035 -1115 48059
rect -1122 47990 -1118 48035
rect -1099 47991 -1091 48005
rect -1187 47988 -1101 47990
rect -1187 47987 -1173 47988
rect -1170 47963 -1163 47988
rect -1170 47918 -1166 47963
rect -1146 47918 -1142 47988
rect -1122 47918 -1118 47988
rect -1115 47987 -1101 47988
rect -1098 47987 -1091 47991
rect -1098 47918 -1094 47987
rect -1074 47974 -1067 47987
rect -1074 47950 -1067 47964
rect -1229 47916 -1077 47918
rect -1229 47909 -1224 47916
rect -1218 47909 -1214 47916
rect -1219 47895 -1214 47909
rect -1229 47894 -1195 47895
rect -1475 47892 -1195 47894
rect -1475 47891 -1461 47892
rect -1458 47891 -1451 47892
rect -1434 47870 -1430 47892
rect -1410 47870 -1406 47892
rect -1386 47870 -1382 47892
rect -2393 47868 -1365 47870
rect -2371 47846 -2366 47868
rect -2348 47846 -2343 47868
rect -2325 47856 -2317 47868
rect -2325 47846 -2320 47856
rect -2317 47854 -2309 47856
rect -2062 47855 -2032 47862
rect -2309 47846 -2301 47854
rect -2070 47848 -2062 47855
rect -2000 47850 -1992 47868
rect -1974 47866 -1944 47868
rect -1960 47865 -1944 47866
rect -1842 47864 -1806 47868
rect -1842 47857 -1798 47862
rect -1806 47855 -1798 47857
rect -1671 47856 -1663 47868
rect -1854 47853 -1842 47855
rect -1663 47854 -1655 47856
rect -2062 47846 -2036 47848
rect -2393 47844 -2036 47846
rect -2032 47846 -2012 47848
rect -2004 47846 -1974 47850
rect -1854 47848 -1806 47853
rect -1864 47846 -1796 47847
rect -1655 47846 -1647 47854
rect -1642 47846 -1637 47868
rect -1619 47846 -1614 47868
rect -1530 47847 -1526 47868
rect -1541 47846 -1507 47847
rect -2032 47844 -1507 47846
rect -2371 47798 -2366 47844
rect -2348 47798 -2343 47844
rect -2325 47840 -2320 47844
rect -2309 47842 -2301 47844
rect -2317 47840 -2309 47842
rect -2325 47828 -2317 47840
rect -2052 47838 -2036 47840
rect -2052 47836 -2032 47838
rect -2062 47830 -2032 47836
rect -2325 47798 -2320 47828
rect -2317 47826 -2309 47828
rect -2092 47814 -2062 47816
rect -2094 47810 -2062 47814
rect -2000 47798 -1992 47844
rect -1904 47837 -1874 47844
rect -1842 47837 -1806 47844
rect -1655 47842 -1647 47844
rect -1663 47840 -1655 47842
rect -1842 47830 -1680 47836
rect -1671 47828 -1663 47840
rect -1663 47826 -1655 47828
rect -1854 47814 -1806 47816
rect -1854 47810 -1680 47814
rect -1642 47798 -1637 47844
rect -1619 47798 -1614 47844
rect -1541 47837 -1536 47844
rect -1530 47837 -1526 47844
rect -1531 47823 -1526 47837
rect -1541 47813 -1536 47823
rect -1530 47813 -1526 47823
rect -1531 47799 -1526 47813
rect -1541 47798 -1507 47799
rect -2393 47796 -1507 47798
rect -2371 47750 -2366 47796
rect -2348 47750 -2343 47796
rect -2325 47750 -2320 47796
rect -2309 47780 -2301 47790
rect -2317 47774 -2309 47780
rect -2097 47774 -2095 47783
rect -2309 47752 -2301 47762
rect -2097 47760 -2095 47764
rect -2292 47759 -2095 47760
rect -2097 47757 -2095 47759
rect -2084 47752 -2083 47795
rect -2069 47788 -2054 47790
rect -2054 47772 -2018 47774
rect -2054 47770 -2004 47772
rect -2059 47766 -2045 47770
rect -2054 47764 -2049 47766
rect -2317 47750 -2309 47752
rect -2084 47750 -2054 47752
rect -2044 47750 -2039 47764
rect -2025 47754 -2014 47760
rect -2000 47754 -1992 47796
rect -1920 47794 -1906 47796
rect -1977 47779 -1929 47785
rect -1655 47780 -1647 47790
rect -1977 47769 -1966 47779
rect -1663 47774 -1655 47780
rect -1977 47757 -1929 47759
rect -2033 47750 -1992 47754
rect -1655 47752 -1647 47762
rect -1663 47750 -1655 47752
rect -1642 47750 -1637 47796
rect -1619 47750 -1614 47796
rect -1541 47789 -1536 47796
rect -1531 47775 -1526 47789
rect -1530 47750 -1526 47775
rect -1506 47771 -1502 47868
rect -2393 47748 -1509 47750
rect -2371 47630 -2366 47748
rect -2348 47630 -2343 47748
rect -2325 47714 -2320 47748
rect -2317 47746 -2309 47748
rect -2084 47735 -2083 47748
rect -2084 47734 -2054 47735
rect -2325 47706 -2317 47714
rect -2325 47686 -2320 47706
rect -2317 47698 -2309 47706
rect -2117 47697 -2095 47707
rect -2045 47704 -2037 47718
rect -2325 47670 -2317 47686
rect -2325 47654 -2320 47670
rect -2309 47658 -2301 47670
rect -2317 47654 -2309 47658
rect -2117 47656 -2095 47663
rect -2069 47662 -2041 47670
rect -2017 47668 -2015 47670
rect -2325 47642 -2317 47654
rect -2125 47647 -2095 47654
rect -2047 47652 -2011 47654
rect -2059 47650 -2011 47652
rect -2000 47650 -1992 47748
rect -1663 47746 -1655 47748
rect -1969 47697 -1929 47709
rect -1671 47706 -1663 47714
rect -1663 47698 -1655 47706
rect -1671 47670 -1663 47686
rect -1655 47658 -1647 47670
rect -1663 47654 -1655 47658
rect -2125 47645 -2117 47647
rect -2059 47646 -2045 47650
rect -2021 47647 -1992 47650
rect -1977 47647 -1929 47654
rect -2325 47630 -2320 47642
rect -2309 47630 -2301 47642
rect -2131 47637 -2129 47642
rect -2125 47639 -2095 47645
rect -2021 47640 -2009 47644
rect -2125 47637 -2117 47639
rect -2133 47630 -2129 47637
rect -2117 47630 -2087 47637
rect -2025 47634 -2021 47640
rect -2000 47634 -1992 47647
rect -1969 47639 -1929 47645
rect -1671 47642 -1663 47654
rect -2033 47630 -1992 47634
rect -1969 47630 -1921 47637
rect -1655 47630 -1647 47642
rect -1642 47630 -1637 47748
rect -1619 47630 -1614 47748
rect -1530 47630 -1526 47748
rect -1523 47747 -1509 47748
rect -1506 47726 -1499 47771
rect -1482 47726 -1478 47868
rect -1458 47843 -1451 47867
rect -1458 47726 -1454 47843
rect -1434 47726 -1430 47868
rect -1410 47726 -1406 47868
rect -1386 47726 -1382 47868
rect -1379 47867 -1365 47868
rect -1362 47867 -1355 47891
rect -1362 47726 -1358 47867
rect -1338 47726 -1334 47892
rect -1314 47726 -1310 47892
rect -1301 47861 -1296 47871
rect -1290 47861 -1286 47892
rect -1291 47847 -1286 47861
rect -1290 47726 -1286 47847
rect -1266 47795 -1262 47892
rect -1266 47771 -1259 47795
rect -1266 47726 -1262 47771
rect -1242 47726 -1238 47892
rect -1229 47885 -1224 47892
rect -1219 47871 -1214 47885
rect -1218 47726 -1214 47871
rect -1194 47843 -1190 47916
rect -1194 47822 -1187 47843
rect -1170 47822 -1166 47916
rect -1146 47822 -1142 47916
rect -1122 47822 -1118 47916
rect -1098 47822 -1094 47916
rect -1091 47915 -1077 47916
rect -1074 47915 -1067 47940
rect -1074 47822 -1070 47915
rect -1050 47822 -1046 47960
rect -1027 47895 -1019 47909
rect -1026 47891 -1019 47895
rect -1026 47822 -1022 47891
rect -1013 47822 -1005 47823
rect -1211 47820 -1005 47822
rect -1211 47819 -1197 47820
rect -1194 47795 -1187 47820
rect -1194 47726 -1190 47795
rect -1170 47726 -1166 47820
rect -1146 47726 -1142 47820
rect -1122 47726 -1118 47820
rect -1098 47726 -1094 47820
rect -1074 47726 -1070 47820
rect -1061 47741 -1056 47751
rect -1050 47741 -1046 47820
rect -1051 47727 -1046 47741
rect -1050 47726 -1046 47727
rect -1026 47726 -1022 47820
rect -1019 47819 -1005 47820
rect -1013 47813 -1008 47819
rect -1003 47799 -998 47813
rect -1002 47727 -998 47799
rect -1013 47726 -981 47727
rect -1523 47724 -981 47726
rect -1523 47723 -1509 47724
rect -1506 47699 -1499 47724
rect -1506 47630 -1502 47699
rect -1482 47630 -1478 47724
rect -1458 47630 -1454 47724
rect -1434 47630 -1430 47724
rect -1410 47630 -1406 47724
rect -1386 47630 -1382 47724
rect -1362 47655 -1358 47724
rect -1373 47654 -1339 47655
rect -1338 47654 -1334 47724
rect -1314 47654 -1310 47724
rect -1290 47654 -1286 47724
rect -1266 47654 -1262 47724
rect -1242 47654 -1238 47724
rect -1218 47654 -1214 47724
rect -1194 47654 -1190 47724
rect -1170 47654 -1166 47724
rect -1157 47693 -1152 47703
rect -1146 47693 -1142 47724
rect -1147 47679 -1142 47693
rect -1157 47669 -1152 47679
rect -1147 47655 -1142 47669
rect -1146 47654 -1142 47655
rect -1122 47654 -1118 47724
rect -1098 47654 -1094 47724
rect -1074 47654 -1070 47724
rect -1050 47654 -1046 47724
rect -1026 47675 -1022 47724
rect -1013 47717 -1008 47724
rect -1002 47717 -998 47724
rect -995 47723 -981 47724
rect -1003 47703 -998 47717
rect -1373 47652 -1029 47654
rect -1373 47645 -1368 47652
rect -1362 47645 -1358 47652
rect -1363 47631 -1358 47645
rect -1373 47630 -1339 47631
rect -2393 47628 -1339 47630
rect -2371 47534 -2366 47628
rect -2348 47534 -2343 47628
rect -2325 47626 -2320 47628
rect -2317 47626 -2309 47628
rect -2131 47626 -2129 47628
rect -2125 47626 -2095 47628
rect -2325 47614 -2317 47626
rect -2117 47621 -2095 47626
rect -2325 47594 -2320 47614
rect -2325 47586 -2317 47594
rect -2325 47534 -2320 47586
rect -2317 47578 -2309 47586
rect -2117 47577 -2095 47587
rect -2045 47584 -2037 47598
rect -2309 47538 -2301 47548
rect -2087 47544 -2076 47552
rect -2017 47548 -2015 47555
rect -2317 47534 -2309 47538
rect -2092 47536 -2087 47544
rect -2092 47534 -2077 47535
rect -2000 47534 -1992 47628
rect -1663 47626 -1655 47628
rect -1671 47614 -1663 47626
rect -1969 47577 -1929 47589
rect -1671 47586 -1663 47594
rect -1663 47578 -1655 47586
rect -1655 47538 -1647 47548
rect -1928 47534 -1924 47535
rect -1854 47534 -1680 47535
rect -1663 47534 -1655 47538
rect -1642 47534 -1637 47628
rect -1619 47534 -1614 47628
rect -1530 47534 -1526 47628
rect -1506 47535 -1502 47628
rect -1517 47534 -1483 47535
rect -2393 47532 -1483 47534
rect -2371 47510 -2366 47532
rect -2348 47510 -2343 47532
rect -2325 47510 -2320 47532
rect -2092 47527 -2037 47532
rect -2021 47527 -1969 47532
rect -1921 47527 -1913 47532
rect -1854 47528 -1680 47532
rect -2100 47525 -2092 47526
rect -2309 47510 -2301 47520
rect -2100 47519 -2087 47525
rect -2051 47512 -2026 47514
rect -2062 47510 -2012 47512
rect -2000 47510 -1992 47527
rect -1969 47519 -1921 47526
rect -1969 47510 -1964 47519
rect -1864 47510 -1796 47511
rect -1655 47510 -1647 47520
rect -1642 47510 -1637 47532
rect -1619 47510 -1614 47532
rect -1530 47510 -1526 47532
rect -1517 47525 -1512 47532
rect -1506 47525 -1502 47532
rect -1507 47511 -1502 47525
rect -1506 47510 -1502 47511
rect -1482 47510 -1478 47628
rect -1458 47510 -1454 47628
rect -1434 47510 -1430 47628
rect -1410 47510 -1406 47628
rect -1397 47597 -1392 47607
rect -1386 47597 -1382 47628
rect -1373 47621 -1368 47628
rect -1363 47607 -1358 47621
rect -1387 47583 -1382 47597
rect -1386 47510 -1382 47583
rect -1362 47531 -1358 47607
rect -1338 47579 -1334 47652
rect -1338 47558 -1331 47579
rect -1314 47558 -1310 47652
rect -1290 47583 -1286 47652
rect -1301 47582 -1267 47583
rect -1266 47582 -1262 47652
rect -1242 47582 -1238 47652
rect -1218 47582 -1214 47652
rect -1194 47582 -1190 47652
rect -1170 47582 -1166 47652
rect -1146 47582 -1142 47652
rect -1122 47627 -1118 47652
rect -1301 47580 -1125 47582
rect -1301 47573 -1296 47580
rect -1290 47573 -1286 47580
rect -1291 47559 -1286 47573
rect -1301 47558 -1267 47559
rect -1355 47556 -1267 47558
rect -1355 47555 -1341 47556
rect -1338 47531 -1331 47556
rect -2393 47508 -1365 47510
rect -2371 47462 -2366 47508
rect -2348 47462 -2343 47508
rect -2325 47462 -2320 47508
rect -2317 47504 -2309 47508
rect -2105 47501 -2092 47504
rect -2092 47478 -2062 47480
rect -2094 47474 -2062 47478
rect -2000 47462 -1992 47508
rect -1663 47504 -1655 47508
rect -1969 47501 -1921 47504
rect -1854 47478 -1806 47480
rect -1854 47474 -1680 47478
rect -1642 47462 -1637 47508
rect -1619 47462 -1614 47508
rect -1530 47462 -1526 47508
rect -1517 47477 -1512 47487
rect -1506 47477 -1502 47508
rect -1507 47463 -1502 47477
rect -1517 47462 -1483 47463
rect -2393 47460 -1483 47462
rect -2371 47438 -2366 47460
rect -2348 47438 -2343 47460
rect -2325 47438 -2320 47460
rect -2072 47458 -2036 47459
rect -2072 47452 -2054 47458
rect -2309 47444 -2301 47452
rect -2317 47438 -2309 47444
rect -2092 47443 -2062 47448
rect -2000 47439 -1992 47460
rect -1938 47459 -1906 47460
rect -1920 47458 -1906 47459
rect -1806 47452 -1680 47458
rect -1854 47443 -1806 47448
rect -1655 47444 -1647 47452
rect -1982 47439 -1966 47440
rect -2000 47438 -1966 47439
rect -1846 47438 -1806 47441
rect -1663 47438 -1655 47444
rect -1642 47438 -1637 47460
rect -1619 47438 -1614 47460
rect -1530 47438 -1526 47460
rect -1517 47453 -1512 47460
rect -1482 47459 -1478 47508
rect -1507 47439 -1502 47453
rect -1493 47449 -1485 47453
rect -1499 47439 -1493 47449
rect -1506 47438 -1502 47439
rect -2393 47436 -1485 47438
rect -2371 47414 -2366 47436
rect -2348 47414 -2343 47436
rect -2325 47414 -2320 47436
rect -2000 47434 -1966 47436
rect -2309 47416 -2301 47424
rect -2062 47423 -2054 47430
rect -2092 47416 -2084 47423
rect -2062 47416 -2026 47418
rect -2317 47414 -2309 47416
rect -2062 47414 -2012 47416
rect -2000 47414 -1992 47434
rect -1982 47433 -1966 47434
rect -1846 47432 -1806 47436
rect -1846 47425 -1798 47430
rect -1806 47423 -1798 47425
rect -1854 47421 -1846 47423
rect -1854 47416 -1806 47421
rect -1655 47416 -1647 47424
rect -1864 47414 -1796 47415
rect -1663 47414 -1655 47416
rect -1642 47414 -1637 47436
rect -1619 47414 -1614 47436
rect -1530 47414 -1526 47436
rect -1506 47414 -1502 47436
rect -1499 47435 -1485 47436
rect -1482 47435 -1475 47459
rect -1482 47414 -1478 47435
rect -1458 47414 -1454 47508
rect -1434 47414 -1430 47508
rect -1410 47414 -1406 47508
rect -1386 47414 -1382 47508
rect -1379 47507 -1365 47508
rect -1362 47507 -1355 47531
rect -1362 47414 -1358 47507
rect -1338 47414 -1334 47531
rect -1314 47414 -1310 47556
rect -1301 47549 -1296 47556
rect -1291 47535 -1286 47549
rect -1290 47414 -1286 47535
rect -1266 47507 -1262 47580
rect -1266 47486 -1259 47507
rect -1242 47486 -1238 47580
rect -1218 47486 -1214 47580
rect -1205 47501 -1200 47511
rect -1194 47501 -1190 47580
rect -1195 47487 -1190 47501
rect -1194 47486 -1190 47487
rect -1170 47486 -1166 47580
rect -1146 47486 -1142 47580
rect -1139 47579 -1125 47580
rect -1122 47579 -1115 47627
rect -1122 47486 -1118 47579
rect -1098 47486 -1094 47652
rect -1074 47486 -1070 47652
rect -1050 47486 -1046 47652
rect -1043 47651 -1029 47652
rect -1026 47651 -1019 47675
rect -1026 47486 -1022 47651
rect -1002 47486 -998 47703
rect -989 47693 -984 47703
rect -979 47679 -974 47693
rect -978 47651 -974 47679
rect -978 47627 -971 47651
rect -978 47486 -974 47627
rect -954 47603 -947 47627
rect -954 47486 -950 47603
rect -931 47559 -923 47573
rect -930 47555 -923 47559
rect -930 47486 -926 47555
rect -917 47486 -909 47487
rect -1283 47484 -909 47486
rect -1283 47483 -1269 47484
rect -1266 47459 -1259 47484
rect -1266 47414 -1262 47459
rect -1242 47414 -1238 47484
rect -1218 47414 -1214 47484
rect -1194 47414 -1190 47484
rect -1170 47435 -1166 47484
rect -2393 47412 -1173 47414
rect -2371 47366 -2366 47412
rect -2348 47366 -2343 47412
rect -2325 47366 -2320 47412
rect -2317 47408 -2309 47412
rect -2062 47408 -2054 47412
rect -2154 47404 -2138 47406
rect -2057 47404 -2054 47408
rect -2292 47398 -2054 47404
rect -2052 47398 -2044 47408
rect -2092 47382 -2062 47384
rect -2094 47378 -2062 47382
rect -2000 47366 -1992 47412
rect -1846 47405 -1806 47412
rect -1663 47408 -1655 47412
rect -1846 47398 -1680 47404
rect -1854 47382 -1806 47384
rect -1854 47378 -1680 47382
rect -1642 47366 -1637 47412
rect -1619 47366 -1614 47412
rect -1530 47366 -1526 47412
rect -1506 47366 -1502 47412
rect -1482 47411 -1478 47412
rect -2393 47364 -1485 47366
rect -2371 47342 -2366 47364
rect -2348 47342 -2343 47364
rect -2325 47342 -2320 47364
rect -2072 47362 -2036 47363
rect -2072 47356 -2054 47362
rect -2309 47348 -2301 47356
rect -2317 47342 -2309 47348
rect -2092 47347 -2062 47352
rect -2000 47343 -1992 47364
rect -1938 47363 -1906 47364
rect -1920 47362 -1906 47363
rect -1806 47356 -1680 47362
rect -1854 47347 -1806 47352
rect -1655 47348 -1647 47356
rect -1982 47343 -1966 47344
rect -2000 47342 -1966 47343
rect -1846 47342 -1806 47345
rect -1663 47342 -1655 47348
rect -1642 47342 -1637 47364
rect -1619 47342 -1614 47364
rect -1530 47342 -1526 47364
rect -1506 47342 -1502 47364
rect -1499 47363 -1485 47364
rect -1482 47363 -1475 47411
rect -1482 47342 -1478 47363
rect -1458 47342 -1454 47412
rect -1434 47342 -1430 47412
rect -1410 47342 -1406 47412
rect -1386 47342 -1382 47412
rect -1362 47342 -1358 47412
rect -1338 47342 -1334 47412
rect -1314 47391 -1310 47412
rect -1325 47390 -1291 47391
rect -1290 47390 -1286 47412
rect -1266 47390 -1262 47412
rect -1242 47390 -1238 47412
rect -1218 47390 -1214 47412
rect -1194 47390 -1190 47412
rect -1187 47411 -1173 47412
rect -1170 47411 -1163 47435
rect -1170 47390 -1166 47411
rect -1146 47390 -1142 47484
rect -1122 47390 -1118 47484
rect -1098 47390 -1094 47484
rect -1074 47390 -1070 47484
rect -1061 47405 -1056 47415
rect -1050 47405 -1046 47484
rect -1051 47391 -1046 47405
rect -1050 47390 -1046 47391
rect -1026 47390 -1022 47484
rect -1013 47429 -1008 47439
rect -1002 47429 -998 47484
rect -1003 47415 -998 47429
rect -1002 47390 -998 47415
rect -978 47390 -974 47484
rect -954 47390 -950 47484
rect -930 47390 -926 47484
rect -923 47483 -909 47484
rect -917 47477 -912 47483
rect -907 47463 -902 47477
rect -906 47390 -902 47463
rect -893 47390 -885 47391
rect -1325 47388 -885 47390
rect -1325 47381 -1320 47388
rect -1314 47381 -1310 47388
rect -1315 47367 -1310 47381
rect -1325 47357 -1320 47367
rect -1315 47343 -1310 47357
rect -1314 47342 -1310 47343
rect -1290 47342 -1286 47388
rect -1266 47342 -1262 47388
rect -1242 47342 -1238 47388
rect -1218 47342 -1214 47388
rect -1194 47343 -1190 47388
rect -1205 47342 -1171 47343
rect -2393 47340 -1171 47342
rect -2371 47318 -2366 47340
rect -2348 47318 -2343 47340
rect -2325 47318 -2320 47340
rect -2000 47338 -1966 47340
rect -2309 47320 -2301 47328
rect -2062 47327 -2054 47334
rect -2092 47320 -2084 47327
rect -2062 47320 -2026 47322
rect -2317 47318 -2309 47320
rect -2062 47318 -2012 47320
rect -2000 47318 -1992 47338
rect -1982 47337 -1966 47338
rect -1846 47336 -1806 47340
rect -1846 47329 -1798 47334
rect -1806 47327 -1798 47329
rect -1854 47325 -1846 47327
rect -1854 47320 -1806 47325
rect -1655 47320 -1647 47328
rect -1864 47318 -1796 47319
rect -1663 47318 -1655 47320
rect -1642 47318 -1637 47340
rect -1619 47318 -1614 47340
rect -1530 47318 -1526 47340
rect -1506 47318 -1502 47340
rect -1482 47318 -1478 47340
rect -1458 47318 -1454 47340
rect -1434 47318 -1430 47340
rect -1410 47318 -1406 47340
rect -1386 47318 -1382 47340
rect -1362 47318 -1358 47340
rect -1338 47318 -1334 47340
rect -1314 47318 -1310 47340
rect -1290 47318 -1286 47340
rect -1266 47318 -1262 47340
rect -1242 47318 -1238 47340
rect -1218 47318 -1214 47340
rect -1205 47333 -1200 47340
rect -1194 47333 -1190 47340
rect -1195 47319 -1190 47333
rect -1194 47318 -1190 47319
rect -1170 47318 -1166 47388
rect -1146 47318 -1142 47388
rect -1122 47318 -1118 47388
rect -1098 47318 -1094 47388
rect -1074 47318 -1070 47388
rect -1050 47318 -1046 47388
rect -1026 47339 -1022 47388
rect -2393 47316 -1029 47318
rect -2371 47270 -2366 47316
rect -2348 47270 -2343 47316
rect -2325 47270 -2320 47316
rect -2317 47312 -2309 47316
rect -2062 47312 -2054 47316
rect -2154 47308 -2138 47310
rect -2057 47308 -2054 47312
rect -2292 47302 -2054 47308
rect -2052 47302 -2044 47312
rect -2092 47286 -2062 47288
rect -2094 47282 -2062 47286
rect -2000 47270 -1992 47316
rect -1846 47309 -1806 47316
rect -1663 47312 -1655 47316
rect -1846 47302 -1680 47308
rect -1854 47286 -1806 47288
rect -1854 47282 -1680 47286
rect -1642 47270 -1637 47316
rect -1619 47270 -1614 47316
rect -1530 47270 -1526 47316
rect -1506 47270 -1502 47316
rect -1482 47270 -1478 47316
rect -1458 47270 -1454 47316
rect -1434 47270 -1430 47316
rect -1410 47270 -1406 47316
rect -1386 47270 -1382 47316
rect -1362 47270 -1358 47316
rect -1338 47270 -1334 47316
rect -1314 47270 -1310 47316
rect -1290 47315 -1286 47316
rect -2393 47268 -1293 47270
rect -2371 47246 -2366 47268
rect -2348 47246 -2343 47268
rect -2325 47246 -2320 47268
rect -2072 47266 -2036 47267
rect -2072 47260 -2054 47266
rect -2309 47252 -2301 47260
rect -2317 47246 -2309 47252
rect -2092 47251 -2062 47256
rect -2000 47247 -1992 47268
rect -1938 47267 -1906 47268
rect -1920 47266 -1906 47267
rect -1806 47260 -1680 47266
rect -1854 47251 -1806 47256
rect -1655 47252 -1647 47260
rect -1982 47247 -1966 47248
rect -2000 47246 -1966 47247
rect -1846 47246 -1806 47249
rect -1663 47246 -1655 47252
rect -1642 47246 -1637 47268
rect -1619 47246 -1614 47268
rect -1589 47246 -1555 47247
rect -2393 47244 -1555 47246
rect -2371 47222 -2366 47244
rect -2348 47222 -2343 47244
rect -2325 47222 -2320 47244
rect -2000 47242 -1966 47244
rect -2309 47224 -2301 47232
rect -2062 47231 -2054 47238
rect -2092 47224 -2084 47231
rect -2062 47224 -2026 47226
rect -2317 47222 -2309 47224
rect -2062 47222 -2012 47224
rect -2000 47222 -1992 47242
rect -1982 47241 -1966 47242
rect -1846 47240 -1806 47244
rect -1846 47233 -1798 47238
rect -1806 47231 -1798 47233
rect -1854 47229 -1846 47231
rect -1854 47224 -1806 47229
rect -1655 47224 -1647 47232
rect -1864 47222 -1796 47223
rect -1663 47222 -1655 47224
rect -1642 47222 -1637 47244
rect -1619 47222 -1614 47244
rect -1530 47222 -1526 47268
rect -1506 47222 -1502 47268
rect -1482 47222 -1478 47268
rect -1458 47222 -1454 47268
rect -1434 47222 -1430 47268
rect -1410 47222 -1406 47268
rect -1386 47222 -1382 47268
rect -1362 47222 -1358 47268
rect -1338 47222 -1334 47268
rect -1314 47222 -1310 47268
rect -1307 47267 -1293 47268
rect -1290 47267 -1283 47315
rect -1290 47222 -1286 47267
rect -1266 47222 -1262 47316
rect -1242 47222 -1238 47316
rect -1218 47222 -1214 47316
rect -1194 47222 -1190 47316
rect -1170 47267 -1166 47316
rect -1170 47243 -1163 47267
rect -1170 47222 -1166 47243
rect -1146 47222 -1142 47316
rect -1122 47222 -1118 47316
rect -1098 47222 -1094 47316
rect -1074 47222 -1070 47316
rect -1050 47223 -1046 47316
rect -1043 47315 -1029 47316
rect -1026 47315 -1019 47339
rect -1061 47222 -1027 47223
rect -2393 47220 -1027 47222
rect -2371 47174 -2366 47220
rect -2348 47174 -2343 47220
rect -2325 47174 -2320 47220
rect -2317 47216 -2309 47220
rect -2062 47216 -2054 47220
rect -2154 47212 -2138 47214
rect -2057 47212 -2054 47216
rect -2292 47206 -2054 47212
rect -2052 47206 -2044 47216
rect -2092 47190 -2062 47192
rect -2094 47186 -2062 47190
rect -2000 47174 -1992 47220
rect -1846 47213 -1806 47220
rect -1663 47216 -1655 47220
rect -1846 47206 -1680 47212
rect -1854 47190 -1806 47192
rect -1854 47186 -1680 47190
rect -1979 47174 -1945 47176
rect -1642 47174 -1637 47220
rect -1619 47174 -1614 47220
rect -1530 47174 -1526 47220
rect -1506 47174 -1502 47220
rect -1482 47174 -1478 47220
rect -1458 47174 -1454 47220
rect -1434 47174 -1430 47220
rect -1410 47174 -1406 47220
rect -1386 47174 -1382 47220
rect -1362 47174 -1358 47220
rect -1338 47174 -1334 47220
rect -1314 47174 -1310 47220
rect -1290 47174 -1286 47220
rect -1266 47174 -1262 47220
rect -1242 47174 -1238 47220
rect -1218 47174 -1214 47220
rect -1194 47174 -1190 47220
rect -1170 47174 -1166 47220
rect -1146 47174 -1142 47220
rect -1122 47174 -1118 47220
rect -1098 47174 -1094 47220
rect -1074 47174 -1070 47220
rect -1061 47213 -1056 47220
rect -1050 47213 -1046 47220
rect -1051 47199 -1046 47213
rect -1050 47174 -1046 47199
rect -1026 47174 -1022 47315
rect -1002 47174 -998 47388
rect -978 47363 -974 47388
rect -978 47339 -971 47363
rect -978 47174 -974 47339
rect -965 47189 -960 47199
rect -954 47189 -950 47388
rect -941 47309 -936 47319
rect -930 47309 -926 47388
rect -931 47295 -926 47309
rect -955 47175 -950 47189
rect -965 47174 -931 47175
rect -2393 47172 -931 47174
rect -2371 47126 -2366 47172
rect -2348 47126 -2343 47172
rect -2325 47126 -2320 47172
rect -2080 47171 -1906 47172
rect -2080 47170 -2036 47171
rect -2080 47164 -2054 47170
rect -2309 47156 -2301 47162
rect -2317 47146 -2309 47156
rect -2070 47155 -2040 47162
rect -2054 47147 -2040 47150
rect -2000 47145 -1992 47171
rect -1920 47170 -1906 47171
rect -1850 47164 -1846 47172
rect -1840 47164 -1792 47172
rect -1969 47152 -1966 47161
rect -1850 47157 -1802 47162
rect -1906 47155 -1802 47157
rect -1655 47156 -1647 47162
rect -1906 47154 -1850 47155
rect -1846 47147 -1802 47153
rect -1663 47146 -1655 47156
rect -1860 47145 -1798 47146
rect -2078 47138 -2070 47145
rect -2309 47128 -2301 47134
rect -2317 47126 -2309 47128
rect -2154 47126 -2145 47136
rect -2044 47135 -2040 47140
rect -2028 47138 -1945 47145
rect -1929 47138 -1794 47145
rect -2070 47128 -2040 47135
rect -2044 47126 -2028 47128
rect -2000 47126 -1992 47138
rect -1860 47137 -1798 47138
rect -1850 47128 -1802 47135
rect -1655 47128 -1647 47134
rect -1978 47126 -1942 47127
rect -1663 47126 -1655 47128
rect -1642 47126 -1637 47172
rect -1619 47126 -1614 47172
rect -1554 47158 -1547 47171
rect -1554 47147 -1547 47148
rect -1530 47126 -1526 47172
rect -1506 47126 -1502 47172
rect -1482 47126 -1478 47172
rect -1469 47141 -1464 47151
rect -1458 47141 -1454 47172
rect -1459 47127 -1454 47141
rect -1469 47126 -1435 47127
rect -2393 47124 -1435 47126
rect -2371 47006 -2366 47124
rect -2348 47006 -2343 47124
rect -2325 47086 -2320 47124
rect -2317 47118 -2309 47124
rect -2145 47120 -2138 47124
rect -2070 47120 -2054 47124
rect -2078 47111 -2054 47118
rect -2062 47086 -2032 47087
rect -2000 47086 -1992 47124
rect -1846 47120 -1802 47124
rect -1846 47110 -1792 47119
rect -1663 47118 -1655 47124
rect -1942 47088 -1937 47100
rect -1850 47097 -1822 47098
rect -1850 47093 -1802 47097
rect -2325 47078 -2317 47086
rect -2062 47084 -1961 47086
rect -2325 47058 -2320 47078
rect -2317 47070 -2309 47078
rect -2062 47071 -2040 47082
rect -2032 47077 -1961 47084
rect -1947 47078 -1942 47086
rect -1842 47084 -1794 47087
rect -2070 47066 -2022 47070
rect -2325 47046 -2317 47058
rect -2137 47049 -2121 47051
rect -2325 47030 -2320 47046
rect -2317 47042 -2309 47046
rect -2292 47044 -2085 47049
rect -2069 47044 -2032 47046
rect -2309 47030 -2301 47042
rect -2125 47038 -2121 47039
rect -2325 47018 -2317 47030
rect -2059 47022 -2045 47026
rect -2325 47006 -2320 47018
rect -2317 47014 -2309 47018
rect -2309 47006 -2301 47014
rect -2025 47010 -2022 47016
rect -2000 47010 -1992 47077
rect -1942 47076 -1937 47078
rect -1932 47068 -1927 47076
rect -1912 47073 -1896 47079
rect -1842 47071 -1802 47082
rect -1671 47078 -1663 47086
rect -1663 47070 -1655 47078
rect -1850 47066 -1680 47070
rect -1671 47046 -1663 47058
rect -1663 47042 -1655 47046
rect -1977 47035 -1929 47041
rect -1974 47026 -1944 47035
rect -1655 47030 -1647 47042
rect -1960 47025 -1944 47026
rect -1671 47018 -1663 47030
rect -1977 47013 -1929 47015
rect -1663 47014 -1655 47018
rect -2033 47008 -1992 47010
rect -2062 47006 -1992 47008
rect -1655 47006 -1647 47014
rect -1642 47006 -1637 47124
rect -1619 47006 -1614 47124
rect -1530 47006 -1526 47124
rect -1506 47006 -1502 47124
rect -1482 47006 -1478 47124
rect -1469 47117 -1464 47124
rect -1459 47103 -1454 47117
rect -1458 47006 -1454 47103
rect -1434 47075 -1430 47172
rect -1434 47054 -1427 47075
rect -1410 47054 -1406 47172
rect -1386 47054 -1382 47172
rect -1362 47054 -1358 47172
rect -1338 47054 -1334 47172
rect -1314 47054 -1310 47172
rect -1290 47054 -1286 47172
rect -1266 47079 -1262 47172
rect -1277 47078 -1243 47079
rect -1242 47078 -1238 47172
rect -1218 47127 -1214 47172
rect -1229 47126 -1195 47127
rect -1194 47126 -1190 47172
rect -1170 47126 -1166 47172
rect -1146 47126 -1142 47172
rect -1122 47126 -1118 47172
rect -1098 47126 -1094 47172
rect -1074 47126 -1070 47172
rect -1050 47126 -1046 47172
rect -1026 47147 -1022 47172
rect -1229 47124 -1029 47126
rect -1229 47117 -1224 47124
rect -1218 47117 -1214 47124
rect -1219 47103 -1214 47117
rect -1229 47093 -1224 47103
rect -1219 47079 -1214 47093
rect -1218 47078 -1214 47079
rect -1194 47078 -1190 47124
rect -1170 47078 -1166 47124
rect -1146 47078 -1142 47124
rect -1122 47078 -1118 47124
rect -1098 47078 -1094 47124
rect -1074 47078 -1070 47124
rect -1050 47078 -1046 47124
rect -1043 47123 -1029 47124
rect -1026 47123 -1019 47147
rect -1026 47078 -1022 47123
rect -1002 47078 -998 47172
rect -978 47078 -974 47172
rect -965 47165 -960 47172
rect -955 47151 -950 47165
rect -954 47078 -950 47151
rect -930 47123 -926 47295
rect -906 47243 -902 47388
rect -899 47387 -885 47388
rect -893 47381 -888 47387
rect -883 47367 -878 47381
rect -882 47272 -878 47367
rect -864 47291 -861 47292
rect -893 47261 -888 47271
rect -883 47247 -878 47261
rect -906 47219 -899 47243
rect -1277 47076 -933 47078
rect -1277 47069 -1272 47076
rect -1266 47069 -1262 47076
rect -1267 47055 -1262 47069
rect -1277 47054 -1243 47055
rect -1451 47052 -1243 47054
rect -1451 47051 -1437 47052
rect -1434 47027 -1427 47052
rect -1434 47006 -1430 47027
rect -1410 47006 -1406 47052
rect -1386 47006 -1382 47052
rect -1362 47006 -1358 47052
rect -1338 47006 -1334 47052
rect -1314 47006 -1310 47052
rect -1290 47006 -1286 47052
rect -1277 47045 -1272 47052
rect -1267 47031 -1262 47045
rect -1266 47006 -1262 47031
rect -1242 47006 -1238 47076
rect -1218 47006 -1214 47076
rect -1194 47051 -1190 47076
rect -2393 47004 -1197 47006
rect -2371 46910 -2366 47004
rect -2348 46910 -2343 47004
rect -2325 47002 -2320 47004
rect -2309 47002 -2301 47004
rect -2325 46990 -2317 47002
rect -2025 47000 -2022 47004
rect -2062 46990 -2032 46991
rect -2325 46970 -2320 46990
rect -2317 46986 -2309 46990
rect -2325 46962 -2317 46970
rect -2325 46910 -2320 46962
rect -2317 46954 -2309 46962
rect -2117 46953 -2095 46963
rect -2045 46960 -2037 46974
rect -2309 46914 -2301 46924
rect -2087 46920 -2076 46928
rect -2017 46924 -2015 46931
rect -2317 46910 -2309 46914
rect -2092 46912 -2087 46920
rect -2092 46910 -2077 46911
rect -2000 46910 -1992 47004
rect -1888 46997 -1874 47004
rect -1655 47002 -1647 47004
rect -1671 46990 -1663 47002
rect -1663 46986 -1655 46990
rect -1969 46953 -1929 46965
rect -1671 46962 -1663 46970
rect -1663 46954 -1655 46962
rect -1655 46914 -1647 46924
rect -1928 46910 -1924 46911
rect -1854 46910 -1680 46911
rect -1663 46910 -1655 46914
rect -1642 46910 -1637 47004
rect -1619 46910 -1614 47004
rect -1530 46910 -1526 47004
rect -1506 46910 -1502 47004
rect -1482 46910 -1478 47004
rect -1458 46910 -1454 47004
rect -1434 46910 -1430 47004
rect -1410 46910 -1406 47004
rect -1386 46910 -1382 47004
rect -1362 46911 -1358 47004
rect -1373 46910 -1339 46911
rect -2393 46908 -1339 46910
rect -2371 46886 -2366 46908
rect -2348 46886 -2343 46908
rect -2325 46886 -2320 46908
rect -2092 46903 -2037 46908
rect -2021 46903 -1969 46908
rect -1921 46903 -1913 46908
rect -1854 46904 -1680 46908
rect -2100 46901 -2092 46902
rect -2309 46886 -2301 46896
rect -2100 46895 -2087 46901
rect -2051 46888 -2026 46890
rect -2062 46886 -2012 46888
rect -2000 46886 -1992 46903
rect -1969 46895 -1921 46902
rect -1969 46886 -1964 46895
rect -1864 46886 -1796 46887
rect -1655 46886 -1647 46896
rect -1642 46886 -1637 46908
rect -1619 46886 -1614 46908
rect -1530 46886 -1526 46908
rect -1506 46886 -1502 46908
rect -1482 46886 -1478 46908
rect -1458 46886 -1454 46908
rect -1434 46886 -1430 46908
rect -1410 46886 -1406 46908
rect -1386 46887 -1382 46908
rect -1373 46901 -1368 46908
rect -1362 46901 -1358 46908
rect -1363 46887 -1358 46901
rect -1397 46886 -1363 46887
rect -2393 46884 -1363 46886
rect -2371 46838 -2366 46884
rect -2348 46838 -2343 46884
rect -2325 46838 -2320 46884
rect -2317 46880 -2309 46884
rect -2105 46877 -2092 46880
rect -2092 46854 -2062 46856
rect -2094 46850 -2062 46854
rect -2000 46838 -1992 46884
rect -1663 46880 -1655 46884
rect -1969 46877 -1921 46880
rect -1854 46854 -1806 46856
rect -1854 46850 -1680 46854
rect -1642 46838 -1637 46884
rect -1619 46838 -1614 46884
rect -1530 46838 -1526 46884
rect -1506 46838 -1502 46884
rect -1482 46838 -1478 46884
rect -1458 46838 -1454 46884
rect -1434 46838 -1430 46884
rect -1410 46838 -1406 46884
rect -1397 46877 -1392 46884
rect -1386 46877 -1382 46884
rect -1387 46863 -1382 46877
rect -1386 46838 -1382 46863
rect -1362 46838 -1358 46887
rect -1338 46838 -1334 47004
rect -1314 46838 -1310 47004
rect -1290 46838 -1286 47004
rect -1266 46838 -1262 47004
rect -1242 47003 -1238 47004
rect -1242 46982 -1235 47003
rect -1218 46982 -1214 47004
rect -1211 47003 -1197 47004
rect -1194 47003 -1187 47051
rect -1194 46982 -1190 47003
rect -1170 46982 -1166 47076
rect -1146 46982 -1142 47076
rect -1122 46982 -1118 47076
rect -1098 46982 -1094 47076
rect -1074 46982 -1070 47076
rect -1050 46982 -1046 47076
rect -1026 46982 -1022 47076
rect -1002 46982 -998 47076
rect -978 46982 -974 47076
rect -954 46982 -950 47076
rect -947 47075 -933 47076
rect -930 47075 -923 47123
rect -930 46982 -926 47075
rect -917 46997 -912 47007
rect -906 46997 -902 47219
rect -907 46983 -902 46997
rect -906 46982 -902 46983
rect -882 46982 -878 47247
rect -858 47206 -854 47272
rect -858 47171 -851 47195
rect -845 47189 -840 47199
rect -835 47175 -830 47189
rect -858 46983 -854 47171
rect -869 46982 -835 46983
rect -1259 46980 -835 46982
rect -1259 46979 -1245 46980
rect -1242 46955 -1235 46980
rect -1242 46838 -1238 46955
rect -1229 46949 -1224 46959
rect -1218 46949 -1214 46980
rect -1219 46935 -1214 46949
rect -1229 46925 -1224 46935
rect -1219 46911 -1214 46925
rect -1218 46838 -1214 46911
rect -1194 46883 -1190 46980
rect -2393 46836 -1197 46838
rect -2371 46790 -2366 46836
rect -2348 46790 -2343 46836
rect -2325 46790 -2320 46836
rect -2309 46820 -2301 46830
rect -2317 46814 -2309 46820
rect -2097 46814 -2095 46823
rect -2309 46792 -2301 46802
rect -2097 46800 -2095 46804
rect -2292 46799 -2095 46800
rect -2097 46797 -2095 46799
rect -2084 46792 -2083 46835
rect -2069 46828 -2054 46830
rect -2054 46812 -2018 46814
rect -2054 46810 -2004 46812
rect -2059 46806 -2045 46810
rect -2054 46804 -2049 46806
rect -2317 46790 -2309 46792
rect -2084 46790 -2054 46792
rect -2044 46790 -2039 46804
rect -2025 46794 -2014 46800
rect -2000 46794 -1992 46836
rect -1920 46834 -1906 46836
rect -1977 46819 -1929 46825
rect -1655 46820 -1647 46830
rect -1977 46809 -1966 46819
rect -1663 46814 -1655 46820
rect -1977 46797 -1929 46799
rect -2033 46790 -1992 46794
rect -1655 46792 -1647 46802
rect -1663 46790 -1655 46792
rect -1642 46790 -1637 46836
rect -1619 46790 -1614 46836
rect -1530 46790 -1526 46836
rect -1506 46790 -1502 46836
rect -1482 46790 -1478 46836
rect -1458 46791 -1454 46836
rect -1469 46790 -1435 46791
rect -2393 46788 -1435 46790
rect -2371 46694 -2366 46788
rect -2348 46694 -2343 46788
rect -2325 46754 -2320 46788
rect -2317 46786 -2309 46788
rect -2084 46775 -2083 46788
rect -2084 46774 -2054 46775
rect -2325 46746 -2317 46754
rect -2325 46694 -2320 46746
rect -2317 46738 -2309 46746
rect -2117 46737 -2095 46747
rect -2045 46744 -2037 46758
rect -2309 46698 -2301 46708
rect -2087 46704 -2076 46712
rect -2017 46708 -2015 46715
rect -2317 46694 -2309 46698
rect -2092 46696 -2087 46704
rect -2092 46694 -2077 46695
rect -2000 46694 -1992 46788
rect -1663 46786 -1655 46788
rect -1969 46737 -1929 46749
rect -1671 46746 -1663 46754
rect -1663 46738 -1655 46746
rect -1655 46698 -1647 46708
rect -1928 46694 -1924 46695
rect -1854 46694 -1680 46695
rect -1663 46694 -1655 46698
rect -1642 46694 -1637 46788
rect -1619 46694 -1614 46788
rect -1530 46694 -1526 46788
rect -1506 46694 -1502 46788
rect -1482 46694 -1478 46788
rect -1469 46781 -1464 46788
rect -1458 46781 -1454 46788
rect -1459 46767 -1454 46781
rect -1458 46694 -1454 46767
rect -1434 46715 -1430 46836
rect -2393 46692 -1437 46694
rect -2371 46670 -2366 46692
rect -2348 46670 -2343 46692
rect -2325 46670 -2320 46692
rect -2092 46687 -2037 46692
rect -2021 46687 -1969 46692
rect -1921 46687 -1913 46692
rect -1854 46688 -1680 46692
rect -2100 46685 -2092 46686
rect -2309 46670 -2301 46680
rect -2100 46679 -2087 46685
rect -2051 46672 -2026 46674
rect -2062 46670 -2012 46672
rect -2000 46670 -1992 46687
rect -1969 46679 -1921 46686
rect -1969 46670 -1964 46679
rect -1864 46670 -1796 46671
rect -1655 46670 -1647 46680
rect -1642 46670 -1637 46692
rect -1619 46670 -1614 46692
rect -1530 46670 -1526 46692
rect -1506 46670 -1502 46692
rect -1482 46670 -1478 46692
rect -1458 46670 -1454 46692
rect -1451 46691 -1437 46692
rect -1434 46691 -1427 46715
rect -1434 46670 -1430 46691
rect -1410 46670 -1406 46836
rect -1386 46670 -1382 46836
rect -1362 46811 -1358 46836
rect -1338 46835 -1334 46836
rect -1338 46811 -1331 46835
rect -1362 46787 -1355 46811
rect -1362 46670 -1358 46787
rect -1338 46670 -1334 46811
rect -1314 46670 -1310 46836
rect -1290 46670 -1286 46836
rect -1266 46670 -1262 46836
rect -1242 46670 -1238 46836
rect -1218 46670 -1214 46836
rect -1211 46835 -1197 46836
rect -1194 46835 -1187 46883
rect -1194 46670 -1190 46835
rect -1170 46670 -1166 46980
rect -1146 46670 -1142 46980
rect -1122 46670 -1118 46980
rect -1098 46670 -1094 46980
rect -1074 46670 -1070 46980
rect -1050 46671 -1046 46980
rect -1061 46670 -1027 46671
rect -2393 46668 -1027 46670
rect -2371 46622 -2366 46668
rect -2348 46622 -2343 46668
rect -2325 46622 -2320 46668
rect -2317 46664 -2309 46668
rect -2105 46661 -2092 46664
rect -2092 46638 -2062 46640
rect -2094 46634 -2062 46638
rect -2000 46622 -1992 46668
rect -1663 46664 -1655 46668
rect -1969 46661 -1921 46664
rect -1854 46638 -1806 46640
rect -1854 46634 -1680 46638
rect -1642 46622 -1637 46668
rect -1619 46622 -1614 46668
rect -1530 46622 -1526 46668
rect -1506 46622 -1502 46668
rect -1482 46622 -1478 46668
rect -1458 46622 -1454 46668
rect -1434 46622 -1430 46668
rect -1410 46622 -1406 46668
rect -1386 46622 -1382 46668
rect -1362 46622 -1358 46668
rect -1349 46637 -1344 46647
rect -1338 46637 -1334 46668
rect -1339 46623 -1334 46637
rect -1314 46622 -1310 46668
rect -1290 46622 -1286 46668
rect -1266 46622 -1262 46668
rect -1242 46622 -1238 46668
rect -1218 46622 -1214 46668
rect -1194 46622 -1190 46668
rect -1170 46622 -1166 46668
rect -1146 46622 -1142 46668
rect -1122 46622 -1118 46668
rect -1098 46622 -1094 46668
rect -1074 46622 -1070 46668
rect -1061 46661 -1056 46668
rect -1050 46661 -1046 46668
rect -1051 46647 -1046 46661
rect -1050 46622 -1046 46647
rect -1026 46622 -1022 46980
rect -1002 46622 -998 46980
rect -978 46743 -974 46980
rect -989 46742 -955 46743
rect -954 46742 -950 46980
rect -930 46742 -926 46980
rect -906 46742 -902 46980
rect -882 46931 -878 46980
rect -869 46973 -864 46980
rect -858 46973 -854 46980
rect -859 46959 -854 46973
rect -882 46907 -875 46931
rect -882 46742 -878 46907
rect -858 46742 -854 46959
rect -834 46907 -830 47175
rect -810 47099 -803 47123
rect -834 46883 -827 46907
rect -834 46742 -830 46883
rect -810 46742 -806 47099
rect -786 47051 -779 47075
rect -786 46863 -782 47051
rect -762 47027 -755 47051
rect -797 46862 -763 46863
rect -762 46862 -758 47027
rect -749 46949 -744 46959
rect -739 46935 -734 46949
rect -738 46862 -734 46935
rect -725 46862 -717 46863
rect -797 46860 -717 46862
rect -797 46853 -792 46860
rect -786 46853 -782 46860
rect -787 46839 -782 46853
rect -797 46829 -792 46839
rect -787 46815 -782 46829
rect -786 46742 -782 46815
rect -762 46787 -758 46860
rect -762 46766 -755 46787
rect -738 46767 -734 46860
rect -731 46859 -717 46860
rect -725 46853 -720 46859
rect -715 46839 -710 46853
rect -749 46766 -715 46767
rect -779 46764 -715 46766
rect -779 46763 -765 46764
rect -989 46740 -765 46742
rect -989 46733 -984 46740
rect -978 46733 -974 46740
rect -979 46719 -974 46733
rect -989 46709 -984 46719
rect -979 46695 -974 46709
rect -978 46671 -974 46695
rect -989 46670 -955 46671
rect -954 46670 -950 46740
rect -941 46685 -936 46695
rect -930 46685 -926 46740
rect -931 46671 -926 46685
rect -930 46670 -926 46671
rect -906 46670 -902 46740
rect -882 46670 -878 46740
rect -858 46670 -854 46740
rect -834 46670 -830 46740
rect -810 46670 -806 46740
rect -786 46670 -782 46740
rect -779 46739 -765 46740
rect -762 46739 -755 46764
rect -749 46757 -744 46764
rect -738 46757 -734 46764
rect -739 46743 -734 46757
rect -762 46670 -758 46739
rect -738 46670 -734 46743
rect -714 46691 -710 46839
rect -701 46733 -696 46743
rect -691 46719 -686 46733
rect -989 46668 -717 46670
rect -989 46661 -984 46668
rect -978 46661 -974 46668
rect -954 46667 -950 46668
rect -979 46647 -974 46661
rect -965 46657 -957 46661
rect -971 46647 -965 46657
rect -954 46646 -947 46667
rect -930 46646 -926 46668
rect -906 46646 -902 46668
rect -882 46646 -878 46668
rect -858 46646 -854 46668
rect -834 46646 -830 46668
rect -810 46646 -806 46668
rect -786 46646 -782 46668
rect -762 46646 -758 46668
rect -738 46646 -734 46668
rect -731 46667 -717 46668
rect -714 46667 -707 46691
rect -714 46646 -710 46667
rect -690 46646 -686 46719
rect -667 46647 -659 46661
rect -971 46644 -669 46646
rect -971 46643 -957 46644
rect -989 46622 -957 46623
rect -2393 46620 -957 46622
rect -2371 46598 -2366 46620
rect -2348 46598 -2343 46620
rect -2325 46598 -2320 46620
rect -2072 46618 -2036 46619
rect -2072 46612 -2054 46618
rect -2309 46604 -2301 46612
rect -2317 46598 -2309 46604
rect -2092 46603 -2062 46608
rect -2000 46599 -1992 46620
rect -1938 46619 -1906 46620
rect -1920 46618 -1906 46619
rect -1806 46612 -1680 46618
rect -1854 46603 -1806 46608
rect -1655 46604 -1647 46612
rect -1982 46599 -1966 46600
rect -2000 46598 -1966 46599
rect -1846 46598 -1806 46601
rect -1663 46598 -1655 46604
rect -1642 46598 -1637 46620
rect -1619 46598 -1614 46620
rect -1530 46598 -1526 46620
rect -1506 46598 -1502 46620
rect -1482 46598 -1478 46620
rect -1458 46598 -1454 46620
rect -1434 46598 -1430 46620
rect -1410 46598 -1406 46620
rect -1386 46599 -1382 46620
rect -1397 46598 -1363 46599
rect -1362 46598 -1358 46620
rect -1349 46598 -1315 46599
rect -2393 46596 -1315 46598
rect -2371 46574 -2366 46596
rect -2348 46574 -2343 46596
rect -2325 46574 -2320 46596
rect -2000 46594 -1966 46596
rect -2309 46576 -2301 46584
rect -2062 46583 -2054 46590
rect -2092 46576 -2084 46583
rect -2062 46576 -2026 46578
rect -2317 46574 -2309 46576
rect -2062 46574 -2012 46576
rect -2000 46574 -1992 46594
rect -1982 46593 -1966 46594
rect -1846 46592 -1806 46596
rect -1846 46585 -1798 46590
rect -1806 46583 -1798 46585
rect -1854 46581 -1846 46583
rect -1854 46576 -1806 46581
rect -1655 46576 -1647 46584
rect -1864 46574 -1796 46575
rect -1663 46574 -1655 46576
rect -1642 46574 -1637 46596
rect -1619 46574 -1614 46596
rect -1530 46574 -1526 46596
rect -1506 46574 -1502 46596
rect -1482 46574 -1478 46596
rect -1458 46574 -1454 46596
rect -1434 46574 -1430 46596
rect -1410 46574 -1406 46596
rect -1397 46589 -1392 46596
rect -1386 46589 -1382 46596
rect -1387 46575 -1382 46589
rect -1397 46574 -1363 46575
rect -2393 46572 -1363 46574
rect -2371 46526 -2366 46572
rect -2348 46526 -2343 46572
rect -2325 46526 -2320 46572
rect -2317 46568 -2309 46572
rect -2062 46568 -2054 46572
rect -2154 46564 -2138 46566
rect -2057 46564 -2054 46568
rect -2292 46558 -2054 46564
rect -2052 46558 -2044 46568
rect -2092 46542 -2062 46544
rect -2094 46538 -2062 46542
rect -2000 46526 -1992 46572
rect -1846 46565 -1806 46572
rect -1663 46568 -1655 46572
rect -1846 46558 -1680 46564
rect -1854 46542 -1806 46544
rect -1854 46538 -1680 46542
rect -1642 46526 -1637 46572
rect -1619 46526 -1614 46572
rect -1530 46526 -1526 46572
rect -1506 46526 -1502 46572
rect -1482 46526 -1478 46572
rect -1458 46526 -1454 46572
rect -1434 46526 -1430 46572
rect -1410 46526 -1406 46572
rect -1397 46565 -1392 46572
rect -1387 46551 -1382 46565
rect -1386 46526 -1382 46551
rect -1362 46526 -1358 46596
rect -1349 46589 -1344 46596
rect -1339 46575 -1334 46589
rect -1338 46526 -1334 46575
rect -1314 46571 -1310 46620
rect -1314 46547 -1307 46571
rect -1290 46526 -1286 46620
rect -1266 46526 -1262 46620
rect -1242 46526 -1238 46620
rect -1218 46526 -1214 46620
rect -1194 46526 -1190 46620
rect -1170 46526 -1166 46620
rect -1146 46526 -1142 46620
rect -1122 46526 -1118 46620
rect -1098 46551 -1094 46620
rect -1109 46550 -1075 46551
rect -1074 46550 -1070 46620
rect -1050 46550 -1046 46620
rect -1026 46595 -1022 46620
rect -1026 46571 -1019 46595
rect -1026 46550 -1022 46571
rect -1002 46550 -998 46620
rect -989 46613 -984 46620
rect -971 46619 -957 46620
rect -954 46619 -947 46644
rect -979 46599 -974 46613
rect -978 46550 -974 46599
rect -954 46595 -950 46619
rect -954 46571 -947 46595
rect -930 46550 -926 46644
rect -906 46619 -902 46644
rect -906 46595 -899 46619
rect -906 46550 -902 46595
rect -882 46550 -878 46644
rect -858 46550 -854 46644
rect -834 46550 -830 46644
rect -810 46550 -806 46644
rect -786 46550 -782 46644
rect -762 46550 -758 46644
rect -738 46550 -734 46644
rect -714 46550 -710 46644
rect -690 46550 -686 46644
rect -683 46643 -669 46644
rect -666 46643 -659 46647
rect -666 46550 -662 46643
rect -642 46571 -635 46595
rect -642 46550 -638 46571
rect -629 46550 -621 46551
rect -1109 46548 -621 46550
rect -1109 46541 -1104 46548
rect -1098 46541 -1094 46548
rect -1099 46527 -1094 46541
rect -1109 46526 -1075 46527
rect -2393 46524 -1075 46526
rect -2371 46502 -2366 46524
rect -2348 46502 -2343 46524
rect -2325 46502 -2320 46524
rect -2072 46522 -2036 46523
rect -2072 46516 -2054 46522
rect -2309 46508 -2301 46516
rect -2317 46502 -2309 46508
rect -2092 46507 -2062 46512
rect -2000 46503 -1992 46524
rect -1938 46523 -1906 46524
rect -1920 46522 -1906 46523
rect -1806 46516 -1680 46522
rect -1854 46507 -1806 46512
rect -1655 46508 -1647 46516
rect -1982 46503 -1966 46504
rect -2000 46502 -1966 46503
rect -1846 46502 -1806 46505
rect -1663 46502 -1655 46508
rect -1642 46502 -1637 46524
rect -1619 46502 -1614 46524
rect -1530 46502 -1526 46524
rect -1506 46502 -1502 46524
rect -1482 46502 -1478 46524
rect -1458 46502 -1454 46524
rect -1434 46502 -1430 46524
rect -1410 46503 -1406 46524
rect -1421 46502 -1387 46503
rect -2393 46500 -1387 46502
rect -2371 46478 -2366 46500
rect -2348 46478 -2343 46500
rect -2325 46478 -2320 46500
rect -2000 46498 -1966 46500
rect -2309 46480 -2301 46488
rect -2062 46487 -2054 46494
rect -2092 46480 -2084 46487
rect -2062 46480 -2026 46482
rect -2317 46478 -2309 46480
rect -2062 46478 -2012 46480
rect -2000 46478 -1992 46498
rect -1982 46497 -1966 46498
rect -1846 46496 -1806 46500
rect -1846 46489 -1798 46494
rect -1806 46487 -1798 46489
rect -1854 46485 -1846 46487
rect -1854 46480 -1806 46485
rect -1655 46480 -1647 46488
rect -1864 46478 -1796 46479
rect -1663 46478 -1655 46480
rect -1642 46478 -1637 46500
rect -1619 46478 -1614 46500
rect -1530 46478 -1526 46500
rect -1506 46478 -1502 46500
rect -1482 46478 -1478 46500
rect -1458 46478 -1454 46500
rect -1434 46478 -1430 46500
rect -1421 46493 -1416 46500
rect -1410 46493 -1406 46500
rect -1411 46479 -1406 46493
rect -1410 46478 -1406 46479
rect -1386 46478 -1382 46524
rect -1362 46523 -1358 46524
rect -2393 46476 -1365 46478
rect -2371 46430 -2366 46476
rect -2348 46430 -2343 46476
rect -2325 46430 -2320 46476
rect -2317 46472 -2309 46476
rect -2062 46472 -2054 46476
rect -2154 46468 -2138 46470
rect -2057 46468 -2054 46472
rect -2292 46462 -2054 46468
rect -2052 46462 -2044 46472
rect -2092 46446 -2062 46448
rect -2094 46442 -2062 46446
rect -2000 46430 -1992 46476
rect -1846 46469 -1806 46476
rect -1663 46472 -1655 46476
rect -1846 46462 -1680 46468
rect -1854 46446 -1806 46448
rect -1854 46442 -1680 46446
rect -1642 46430 -1637 46476
rect -1619 46430 -1614 46476
rect -1530 46430 -1526 46476
rect -1506 46430 -1502 46476
rect -1482 46430 -1478 46476
rect -1458 46430 -1454 46476
rect -1445 46445 -1440 46455
rect -1434 46445 -1430 46476
rect -1435 46431 -1430 46445
rect -1410 46430 -1406 46476
rect -1386 46430 -1382 46476
rect -1379 46475 -1365 46476
rect -1362 46475 -1355 46523
rect -1362 46430 -1358 46475
rect -1349 46469 -1344 46479
rect -1338 46469 -1334 46524
rect -1339 46455 -1334 46469
rect -1314 46499 -1307 46523
rect -1349 46430 -1315 46431
rect -2393 46428 -1315 46430
rect -2371 46406 -2366 46428
rect -2348 46406 -2343 46428
rect -2325 46406 -2320 46428
rect -2072 46426 -2036 46427
rect -2072 46420 -2054 46426
rect -2309 46412 -2301 46420
rect -2317 46406 -2309 46412
rect -2092 46411 -2062 46416
rect -2000 46407 -1992 46428
rect -1938 46427 -1906 46428
rect -1920 46426 -1906 46427
rect -1806 46420 -1680 46426
rect -1854 46411 -1806 46416
rect -1655 46412 -1647 46420
rect -1982 46407 -1966 46408
rect -2000 46406 -1966 46407
rect -1846 46406 -1806 46409
rect -1663 46406 -1655 46412
rect -1642 46406 -1637 46428
rect -1619 46406 -1614 46428
rect -1530 46406 -1526 46428
rect -1506 46406 -1502 46428
rect -1482 46406 -1478 46428
rect -1458 46406 -1454 46428
rect -1445 46406 -1411 46407
rect -2393 46404 -1411 46406
rect -2371 46382 -2366 46404
rect -2348 46382 -2343 46404
rect -2325 46382 -2320 46404
rect -2000 46402 -1966 46404
rect -2309 46384 -2301 46392
rect -2062 46391 -2054 46398
rect -2092 46384 -2084 46391
rect -2062 46384 -2026 46386
rect -2317 46382 -2309 46384
rect -2062 46382 -2012 46384
rect -2000 46382 -1992 46402
rect -1982 46401 -1966 46402
rect -1846 46400 -1806 46404
rect -1846 46393 -1798 46398
rect -1806 46391 -1798 46393
rect -1854 46389 -1846 46391
rect -1854 46384 -1806 46389
rect -1655 46384 -1647 46392
rect -1864 46382 -1796 46383
rect -1663 46382 -1655 46384
rect -1642 46382 -1637 46404
rect -1619 46382 -1614 46404
rect -1530 46382 -1526 46404
rect -1506 46382 -1502 46404
rect -1482 46383 -1478 46404
rect -1493 46382 -1459 46383
rect -2393 46380 -1459 46382
rect -2371 46334 -2366 46380
rect -2348 46334 -2343 46380
rect -2325 46334 -2320 46380
rect -2317 46376 -2309 46380
rect -2062 46376 -2054 46380
rect -2154 46372 -2138 46374
rect -2057 46372 -2054 46376
rect -2292 46366 -2054 46372
rect -2052 46366 -2044 46376
rect -2092 46350 -2062 46352
rect -2094 46346 -2062 46350
rect -2000 46334 -1992 46380
rect -1846 46373 -1806 46380
rect -1663 46376 -1655 46380
rect -1846 46366 -1680 46372
rect -1854 46350 -1806 46352
rect -1854 46346 -1680 46350
rect -1642 46334 -1637 46380
rect -1619 46334 -1614 46380
rect -1530 46334 -1526 46380
rect -1506 46334 -1502 46380
rect -1493 46373 -1488 46380
rect -1482 46373 -1478 46380
rect -1483 46359 -1478 46373
rect -1482 46334 -1478 46359
rect -1458 46334 -1454 46404
rect -1445 46397 -1440 46404
rect -1435 46383 -1430 46397
rect -1434 46334 -1430 46383
rect -1410 46379 -1406 46428
rect -1386 46427 -1382 46428
rect -1386 46403 -1379 46427
rect -1410 46355 -1403 46379
rect -1386 46334 -1382 46403
rect -1362 46334 -1358 46428
rect -1349 46421 -1344 46428
rect -1339 46407 -1334 46421
rect -1338 46334 -1334 46407
rect -1314 46403 -1310 46499
rect -1314 46379 -1307 46403
rect -2393 46332 -1317 46334
rect -2371 46310 -2366 46332
rect -2348 46310 -2343 46332
rect -2325 46310 -2320 46332
rect -2072 46330 -2036 46331
rect -2072 46324 -2054 46330
rect -2309 46316 -2301 46324
rect -2317 46310 -2309 46316
rect -2092 46315 -2062 46320
rect -2000 46311 -1992 46332
rect -1938 46331 -1906 46332
rect -1920 46330 -1906 46331
rect -1806 46324 -1680 46330
rect -1854 46315 -1806 46320
rect -1655 46316 -1647 46324
rect -1982 46311 -1966 46312
rect -2000 46310 -1966 46311
rect -1846 46310 -1806 46313
rect -1663 46310 -1655 46316
rect -1642 46310 -1637 46332
rect -1619 46310 -1614 46332
rect -1530 46310 -1526 46332
rect -1506 46310 -1502 46332
rect -1482 46310 -1478 46332
rect -1458 46310 -1454 46332
rect -1434 46310 -1430 46332
rect -2393 46308 -1413 46310
rect -2371 46286 -2366 46308
rect -2348 46286 -2343 46308
rect -2325 46286 -2320 46308
rect -2000 46306 -1966 46308
rect -2309 46288 -2301 46296
rect -2062 46295 -2054 46302
rect -2092 46288 -2084 46295
rect -2062 46288 -2026 46290
rect -2317 46286 -2309 46288
rect -2062 46286 -2012 46288
rect -2000 46286 -1992 46306
rect -1982 46305 -1966 46306
rect -1846 46304 -1806 46308
rect -1846 46297 -1798 46302
rect -1806 46295 -1798 46297
rect -1854 46293 -1846 46295
rect -1854 46288 -1806 46293
rect -1655 46288 -1647 46296
rect -1864 46286 -1796 46287
rect -1663 46286 -1655 46288
rect -1642 46286 -1637 46308
rect -1619 46286 -1614 46308
rect -1530 46286 -1526 46308
rect -1506 46286 -1502 46308
rect -1482 46286 -1478 46308
rect -1458 46307 -1454 46308
rect -2393 46284 -1461 46286
rect -2371 46214 -2366 46284
rect -2348 46214 -2343 46284
rect -2325 46214 -2320 46284
rect -2317 46280 -2309 46284
rect -2062 46280 -2054 46284
rect -2154 46276 -2138 46278
rect -2057 46276 -2054 46280
rect -2292 46270 -2054 46276
rect -2052 46270 -2044 46280
rect -2092 46254 -2062 46256
rect -2094 46250 -2062 46254
rect -2309 46220 -2301 46226
rect -2317 46214 -2309 46220
rect -2000 46214 -1992 46284
rect -1846 46277 -1806 46284
rect -1663 46280 -1655 46284
rect -1846 46270 -1680 46276
rect -1854 46254 -1806 46256
rect -1854 46250 -1680 46254
rect -1655 46220 -1647 46226
rect -1663 46214 -1655 46220
rect -1642 46214 -1637 46284
rect -1619 46214 -1614 46284
rect -1530 46214 -1526 46284
rect -1506 46214 -1502 46284
rect -1482 46214 -1478 46284
rect -1475 46283 -1461 46284
rect -1458 46283 -1451 46307
rect -1458 46214 -1454 46283
rect -1434 46214 -1430 46308
rect -1427 46307 -1413 46308
rect -1410 46307 -1403 46331
rect -1410 46214 -1406 46307
rect -1386 46214 -1382 46332
rect -1362 46214 -1358 46332
rect -1338 46214 -1334 46332
rect -1331 46331 -1317 46332
rect -1314 46331 -1307 46355
rect -1314 46214 -1310 46331
rect -1290 46214 -1286 46524
rect -1266 46214 -1262 46524
rect -1242 46239 -1238 46524
rect -1253 46238 -1219 46239
rect -1218 46238 -1214 46524
rect -1194 46238 -1190 46524
rect -1170 46238 -1166 46524
rect -1146 46238 -1142 46524
rect -1122 46238 -1118 46524
rect -1109 46517 -1104 46524
rect -1099 46503 -1094 46517
rect -1098 46238 -1094 46503
rect -1074 46475 -1070 46548
rect -1074 46454 -1067 46475
rect -1050 46454 -1046 46548
rect -1026 46454 -1022 46548
rect -1002 46454 -998 46548
rect -978 46454 -974 46548
rect -954 46523 -947 46547
rect -954 46454 -950 46523
rect -930 46454 -926 46548
rect -906 46454 -902 46548
rect -882 46454 -878 46548
rect -858 46454 -854 46548
rect -834 46454 -830 46548
rect -810 46454 -806 46548
rect -786 46454 -782 46548
rect -762 46454 -758 46548
rect -738 46454 -734 46548
rect -714 46454 -710 46548
rect -690 46454 -686 46548
rect -666 46454 -662 46548
rect -642 46454 -638 46548
rect -635 46547 -621 46548
rect -629 46541 -624 46547
rect -619 46527 -614 46541
rect -618 46480 -614 46527
rect -629 46469 -624 46479
rect -619 46455 -614 46469
rect -605 46465 -597 46469
rect -611 46455 -605 46465
rect -618 46454 -614 46455
rect -1091 46452 -597 46454
rect -1091 46451 -1077 46452
rect -1074 46427 -1067 46452
rect -1085 46277 -1080 46287
rect -1074 46277 -1070 46427
rect -1061 46301 -1056 46311
rect -1050 46301 -1046 46452
rect -1051 46287 -1046 46301
rect -1075 46263 -1070 46277
rect -1074 46238 -1070 46263
rect -1050 46238 -1046 46287
rect -1026 46238 -1022 46452
rect -1002 46359 -998 46452
rect -1013 46358 -979 46359
rect -978 46358 -974 46452
rect -954 46358 -950 46452
rect -930 46358 -926 46452
rect -906 46358 -902 46452
rect -882 46358 -878 46452
rect -858 46358 -854 46452
rect -834 46358 -830 46452
rect -810 46358 -806 46452
rect -786 46358 -782 46452
rect -762 46358 -758 46452
rect -738 46358 -734 46452
rect -714 46358 -710 46452
rect -690 46358 -686 46452
rect -666 46358 -662 46452
rect -642 46358 -638 46452
rect -618 46358 -614 46452
rect -611 46451 -597 46452
rect -594 46451 -587 46475
rect -594 46414 -590 46451
rect -594 46379 -587 46403
rect -594 46358 -590 46379
rect -570 46358 -566 46424
rect -557 46358 -549 46359
rect -1013 46356 -549 46358
rect -1013 46349 -1008 46356
rect -1002 46349 -998 46356
rect -1003 46335 -998 46349
rect -1013 46325 -1008 46335
rect -1003 46311 -998 46325
rect -1002 46238 -998 46311
rect -978 46283 -974 46356
rect -1253 46236 -981 46238
rect -1253 46229 -1248 46236
rect -1242 46229 -1238 46236
rect -1243 46215 -1238 46229
rect -1253 46214 -1219 46215
rect -2393 46212 -1219 46214
rect -2371 46118 -2366 46212
rect -2348 46118 -2343 46212
rect -2325 46150 -2320 46212
rect -2317 46210 -2309 46212
rect -2000 46211 -1966 46212
rect -2000 46210 -1982 46211
rect -1663 46210 -1655 46212
rect -2028 46202 -2018 46204
rect -2309 46192 -2301 46198
rect -2091 46192 -2061 46199
rect -2317 46182 -2309 46192
rect -2044 46190 -2028 46192
rect -2026 46190 -2014 46202
rect -2084 46184 -2061 46190
rect -2044 46188 -2014 46190
rect -2292 46174 -2054 46183
rect -2325 46142 -2317 46150
rect -2325 46122 -2320 46142
rect -2317 46134 -2309 46142
rect -2325 46118 -2317 46122
rect -2000 46118 -1992 46210
rect -1982 46209 -1966 46210
rect -1980 46192 -1932 46199
rect -1655 46192 -1647 46198
rect -1846 46174 -1680 46183
rect -1663 46182 -1655 46192
rect -1671 46142 -1663 46150
rect -1663 46134 -1655 46142
rect -1671 46118 -1663 46122
rect -1642 46118 -1637 46212
rect -1619 46118 -1614 46212
rect -1530 46118 -1526 46212
rect -1517 46157 -1512 46167
rect -1506 46157 -1502 46212
rect -1507 46143 -1502 46157
rect -1506 46118 -1502 46143
rect -1482 46118 -1478 46212
rect -1458 46118 -1454 46212
rect -1434 46118 -1430 46212
rect -1410 46118 -1406 46212
rect -1386 46118 -1382 46212
rect -1362 46118 -1358 46212
rect -1338 46118 -1334 46212
rect -1314 46118 -1310 46212
rect -1290 46118 -1286 46212
rect -1266 46118 -1262 46212
rect -1253 46205 -1248 46212
rect -1243 46191 -1238 46205
rect -1242 46118 -1238 46191
rect -1218 46163 -1214 46236
rect -2393 46116 -1221 46118
rect -2371 46070 -2366 46116
rect -2348 46070 -2343 46116
rect -2325 46108 -2317 46116
rect -2018 46115 -2004 46116
rect -2000 46115 -1992 46116
rect -2072 46114 -1928 46115
rect -2072 46108 -2053 46114
rect -2325 46092 -2320 46108
rect -2317 46106 -2309 46108
rect -2309 46094 -2301 46106
rect -2092 46099 -2062 46104
rect -2317 46092 -2309 46094
rect -2325 46080 -2317 46092
rect -2098 46086 -2096 46097
rect -2092 46086 -2084 46099
rect -2000 46098 -1992 46114
rect -1972 46108 -1928 46114
rect -1924 46108 -1918 46116
rect -1671 46108 -1663 46116
rect -1663 46106 -1655 46108
rect -2083 46088 -2062 46097
rect -2027 46096 -1992 46098
rect -2018 46088 -2002 46096
rect -2000 46088 -1992 46096
rect -2100 46081 -2096 46086
rect -2083 46081 -2053 46086
rect -2003 46084 -1990 46088
rect -1972 46086 -1964 46095
rect -1928 46094 -1924 46097
rect -1655 46094 -1647 46106
rect -1663 46092 -1655 46094
rect -2325 46070 -2320 46080
rect -2317 46078 -2309 46080
rect -2309 46070 -2301 46078
rect -2004 46074 -2003 46084
rect -2062 46070 -2012 46072
rect -2000 46070 -1992 46084
rect -1972 46081 -1924 46086
rect -1864 46081 -1796 46087
rect -1671 46080 -1663 46092
rect -1663 46078 -1655 46080
rect -1864 46070 -1796 46071
rect -1655 46070 -1647 46078
rect -1642 46070 -1637 46116
rect -1619 46070 -1614 46116
rect -1530 46070 -1526 46116
rect -1506 46070 -1502 46116
rect -1482 46091 -1478 46116
rect -2393 46068 -1485 46070
rect -2371 46022 -2366 46068
rect -2348 46022 -2343 46068
rect -2325 46064 -2320 46068
rect -2309 46066 -2301 46068
rect -2317 46064 -2309 46066
rect -2325 46052 -2317 46064
rect -2325 46022 -2320 46052
rect -2317 46050 -2309 46052
rect -2092 46038 -2062 46040
rect -2094 46034 -2062 46038
rect -2000 46022 -1992 46068
rect -1655 46066 -1647 46068
rect -1663 46064 -1655 46066
rect -1671 46052 -1663 46064
rect -1663 46050 -1655 46052
rect -1854 46038 -1806 46040
rect -1854 46034 -1680 46038
rect -1642 46022 -1637 46068
rect -1619 46022 -1614 46068
rect -1530 46022 -1526 46068
rect -1506 46022 -1502 46068
rect -1499 46067 -1485 46068
rect -1482 46067 -1475 46091
rect -1482 46022 -1478 46067
rect -1458 46022 -1454 46116
rect -1434 46022 -1430 46116
rect -1410 46022 -1406 46116
rect -1386 46022 -1382 46116
rect -1362 46022 -1358 46116
rect -1338 46022 -1334 46116
rect -1314 46022 -1310 46116
rect -1290 46022 -1286 46116
rect -1266 46022 -1262 46116
rect -1242 46022 -1238 46116
rect -1235 46115 -1221 46116
rect -1218 46115 -1211 46163
rect -1218 46022 -1214 46115
rect -1194 46022 -1190 46236
rect -1170 46022 -1166 46236
rect -1146 46022 -1142 46236
rect -1133 46061 -1128 46071
rect -1122 46061 -1118 46236
rect -1123 46047 -1118 46061
rect -1122 46022 -1118 46047
rect -1098 46022 -1094 46236
rect -1074 46022 -1070 46236
rect -1050 46211 -1046 46236
rect -1026 46235 -1022 46236
rect -1026 46211 -1019 46235
rect -1050 46187 -1043 46211
rect -1050 46022 -1046 46187
rect -1026 46022 -1022 46211
rect -1002 46022 -998 46236
rect -995 46235 -981 46236
rect -978 46235 -971 46283
rect -978 46022 -974 46235
rect -954 46022 -950 46356
rect -930 46022 -926 46356
rect -906 46022 -902 46356
rect -882 46022 -878 46356
rect -869 46085 -864 46095
rect -858 46085 -854 46356
rect -834 46143 -830 46356
rect -845 46142 -811 46143
rect -810 46142 -806 46356
rect -786 46142 -782 46356
rect -762 46142 -758 46356
rect -738 46142 -734 46356
rect -714 46142 -710 46356
rect -690 46142 -686 46356
rect -666 46142 -662 46356
rect -642 46142 -638 46356
rect -618 46142 -614 46356
rect -594 46142 -590 46356
rect -570 46142 -566 46356
rect -563 46355 -549 46356
rect -557 46349 -552 46355
rect -547 46335 -542 46349
rect -546 46142 -542 46335
rect -533 46229 -528 46239
rect -523 46215 -518 46229
rect -522 46142 -518 46215
rect -509 46142 -501 46143
rect -845 46140 -501 46142
rect -845 46133 -840 46140
rect -834 46133 -830 46140
rect -835 46119 -830 46133
rect -845 46109 -840 46119
rect -835 46095 -830 46109
rect -859 46071 -854 46085
rect -858 46022 -854 46071
rect -834 46022 -830 46095
rect -810 46067 -806 46140
rect -2393 46020 -813 46022
rect -2371 45998 -2366 46020
rect -2348 45998 -2343 46020
rect -2325 45998 -2320 46020
rect -2072 46018 -2036 46019
rect -2072 46012 -2054 46018
rect -2309 46004 -2301 46012
rect -2317 45998 -2309 46004
rect -2092 46003 -2062 46008
rect -2000 45999 -1992 46020
rect -1938 46019 -1906 46020
rect -1920 46018 -1906 46019
rect -1806 46012 -1680 46018
rect -1854 46003 -1806 46008
rect -1655 46004 -1647 46012
rect -1982 45999 -1966 46000
rect -2000 45998 -1966 45999
rect -1846 45998 -1806 46001
rect -1663 45998 -1655 46004
rect -1642 45998 -1637 46020
rect -1619 45998 -1614 46020
rect -1530 45998 -1526 46020
rect -1506 45998 -1502 46020
rect -1482 45998 -1478 46020
rect -1458 45998 -1454 46020
rect -1434 45998 -1430 46020
rect -1410 45998 -1406 46020
rect -1386 45998 -1382 46020
rect -1362 45998 -1358 46020
rect -1338 45998 -1334 46020
rect -1314 45998 -1310 46020
rect -1290 45998 -1286 46020
rect -1266 45998 -1262 46020
rect -1242 45998 -1238 46020
rect -1218 45998 -1214 46020
rect -1194 45998 -1190 46020
rect -1170 45998 -1166 46020
rect -1146 45998 -1142 46020
rect -1122 45998 -1118 46020
rect -1098 45998 -1094 46020
rect -1074 45998 -1070 46020
rect -1050 45998 -1046 46020
rect -1026 45998 -1022 46020
rect -1002 45998 -998 46020
rect -978 45998 -974 46020
rect -954 45998 -950 46020
rect -930 45998 -926 46020
rect -906 45998 -902 46020
rect -882 45998 -878 46020
rect -858 45999 -854 46020
rect -834 46019 -830 46020
rect -827 46019 -813 46020
rect -810 46019 -803 46067
rect -869 45998 -837 45999
rect -2393 45996 -837 45998
rect -2371 45974 -2366 45996
rect -2348 45974 -2343 45996
rect -2325 45974 -2320 45996
rect -2000 45994 -1966 45996
rect -2309 45976 -2301 45984
rect -2062 45983 -2054 45990
rect -2092 45976 -2084 45983
rect -2062 45976 -2026 45978
rect -2317 45974 -2309 45976
rect -2062 45974 -2012 45976
rect -2000 45974 -1992 45994
rect -1982 45993 -1966 45994
rect -1846 45992 -1806 45996
rect -1846 45985 -1798 45990
rect -1806 45983 -1798 45985
rect -1854 45981 -1846 45983
rect -1854 45976 -1806 45981
rect -1655 45976 -1647 45984
rect -1864 45974 -1796 45975
rect -1663 45974 -1655 45976
rect -1642 45974 -1637 45996
rect -1619 45974 -1614 45996
rect -1530 45974 -1526 45996
rect -1506 45974 -1502 45996
rect -1482 45974 -1478 45996
rect -1458 45974 -1454 45996
rect -1434 45974 -1430 45996
rect -1410 45974 -1406 45996
rect -1386 45974 -1382 45996
rect -1362 45974 -1358 45996
rect -1338 45974 -1334 45996
rect -1314 45974 -1310 45996
rect -1290 45974 -1286 45996
rect -1266 45974 -1262 45996
rect -1242 45974 -1238 45996
rect -1218 45974 -1214 45996
rect -1194 45974 -1190 45996
rect -1170 45974 -1166 45996
rect -1146 45974 -1142 45996
rect -1122 45974 -1118 45996
rect -1098 45995 -1094 45996
rect -2393 45972 -1101 45974
rect -2371 45926 -2366 45972
rect -2348 45926 -2343 45972
rect -2325 45926 -2320 45972
rect -2317 45968 -2309 45972
rect -2062 45968 -2054 45972
rect -2154 45964 -2138 45966
rect -2057 45964 -2054 45968
rect -2292 45958 -2054 45964
rect -2052 45958 -2044 45968
rect -2092 45942 -2062 45944
rect -2094 45938 -2062 45942
rect -2000 45926 -1992 45972
rect -1846 45965 -1806 45972
rect -1663 45968 -1655 45972
rect -1846 45958 -1680 45964
rect -1854 45942 -1806 45944
rect -1854 45938 -1680 45942
rect -1926 45926 -1892 45929
rect -1642 45926 -1637 45972
rect -1619 45926 -1614 45972
rect -1530 45926 -1526 45972
rect -1506 45926 -1502 45972
rect -1482 45926 -1478 45972
rect -1458 45926 -1454 45972
rect -1434 45926 -1430 45972
rect -1410 45926 -1406 45972
rect -1386 45926 -1382 45972
rect -1362 45926 -1358 45972
rect -1338 45926 -1334 45972
rect -1314 45926 -1310 45972
rect -1290 45926 -1286 45972
rect -1266 45926 -1262 45972
rect -1242 45926 -1238 45972
rect -1218 45926 -1214 45972
rect -1194 45926 -1190 45972
rect -1170 45926 -1166 45972
rect -1146 45926 -1142 45972
rect -1122 45926 -1118 45972
rect -1115 45971 -1101 45972
rect -1098 45971 -1091 45995
rect -1098 45926 -1094 45971
rect -1074 45926 -1070 45996
rect -1050 45926 -1046 45996
rect -1026 45926 -1022 45996
rect -1002 45926 -998 45996
rect -978 45926 -974 45996
rect -954 45926 -950 45996
rect -930 45926 -926 45996
rect -906 45926 -902 45996
rect -882 45926 -878 45996
rect -869 45989 -864 45996
rect -858 45989 -854 45996
rect -851 45995 -837 45996
rect -834 45995 -827 46019
rect -859 45975 -854 45989
rect -858 45926 -854 45975
rect -834 45926 -830 45995
rect -821 45941 -816 45951
rect -810 45941 -806 46019
rect -811 45927 -806 45941
rect -821 45926 -787 45927
rect -2393 45924 -787 45926
rect -2371 45902 -2366 45924
rect -2348 45902 -2343 45924
rect -2325 45902 -2320 45924
rect -2054 45923 -1906 45924
rect -2054 45922 -2036 45923
rect -2309 45908 -2301 45918
rect -2317 45902 -2309 45908
rect -2068 45907 -2038 45914
rect -2000 45906 -1992 45923
rect -1920 45922 -1906 45923
rect -1846 45916 -1794 45924
rect -1852 45909 -1804 45914
rect -1902 45907 -1804 45909
rect -1655 45908 -1647 45918
rect -2000 45904 -1975 45906
rect -1902 45905 -1852 45907
rect -2025 45902 -1975 45904
rect -1846 45902 -1804 45905
rect -1663 45902 -1655 45908
rect -1642 45902 -1637 45924
rect -1619 45902 -1614 45924
rect -1530 45902 -1526 45924
rect -1506 45902 -1502 45924
rect -1482 45902 -1478 45924
rect -1458 45902 -1454 45924
rect -1434 45902 -1430 45924
rect -1410 45902 -1406 45924
rect -1386 45902 -1382 45924
rect -1362 45902 -1358 45924
rect -1338 45902 -1334 45924
rect -1314 45902 -1310 45924
rect -1290 45902 -1286 45924
rect -1266 45902 -1262 45924
rect -1242 45902 -1238 45924
rect -1218 45902 -1214 45924
rect -1194 45902 -1190 45924
rect -1170 45902 -1166 45924
rect -1146 45902 -1142 45924
rect -1122 45902 -1118 45924
rect -1098 45902 -1094 45924
rect -1074 45902 -1070 45924
rect -1050 45902 -1046 45924
rect -1026 45902 -1022 45924
rect -1002 45902 -998 45924
rect -978 45902 -974 45924
rect -954 45902 -950 45924
rect -930 45902 -926 45924
rect -906 45902 -902 45924
rect -882 45902 -878 45924
rect -858 45903 -854 45924
rect -834 45923 -830 45924
rect -869 45902 -837 45903
rect -2393 45900 -837 45902
rect -2371 45878 -2366 45900
rect -2348 45878 -2343 45900
rect -2325 45878 -2320 45900
rect -2054 45899 -2038 45900
rect -2000 45899 -1966 45900
rect -1846 45899 -1804 45900
rect -2000 45898 -1975 45899
rect -2076 45890 -2054 45897
rect -2309 45880 -2301 45890
rect -2044 45887 -2038 45892
rect -2028 45890 -2001 45897
rect -2054 45880 -2038 45887
rect -2015 45889 -2001 45890
rect -2015 45880 -2014 45889
rect -2317 45878 -2309 45880
rect -2044 45878 -2028 45880
rect -2000 45878 -1992 45898
rect -1982 45897 -1975 45898
rect -1862 45897 -1798 45898
rect -1985 45890 -1796 45897
rect -1862 45889 -1798 45890
rect -1852 45880 -1804 45887
rect -1655 45880 -1647 45890
rect -1976 45878 -1940 45879
rect -1663 45878 -1655 45880
rect -1642 45878 -1637 45900
rect -1619 45878 -1614 45900
rect -1530 45878 -1526 45900
rect -1506 45878 -1502 45900
rect -1482 45878 -1478 45900
rect -1458 45878 -1454 45900
rect -1434 45878 -1430 45900
rect -1410 45878 -1406 45900
rect -1386 45878 -1382 45900
rect -1362 45878 -1358 45900
rect -1338 45878 -1334 45900
rect -1314 45878 -1310 45900
rect -1290 45878 -1286 45900
rect -1266 45878 -1262 45900
rect -1242 45878 -1238 45900
rect -1218 45878 -1214 45900
rect -1194 45878 -1190 45900
rect -1170 45878 -1166 45900
rect -1146 45878 -1142 45900
rect -1122 45878 -1118 45900
rect -1098 45878 -1094 45900
rect -1074 45878 -1070 45900
rect -1050 45878 -1046 45900
rect -1026 45878 -1022 45900
rect -1002 45878 -998 45900
rect -978 45878 -974 45900
rect -954 45878 -950 45900
rect -930 45878 -926 45900
rect -906 45878 -902 45900
rect -882 45878 -878 45900
rect -869 45893 -864 45900
rect -858 45893 -854 45900
rect -851 45899 -837 45900
rect -834 45899 -827 45923
rect -821 45917 -816 45924
rect -811 45903 -806 45917
rect -859 45879 -854 45893
rect -869 45878 -835 45879
rect -2393 45876 -835 45878
rect -2371 45435 -2366 45876
rect -2361 45455 -2353 45465
rect -2348 45455 -2343 45876
rect -2351 45439 -2343 45455
rect -2371 45409 -2363 45435
rect -2383 45237 -2376 45247
rect -2371 45237 -2366 45409
rect -2373 45226 -2366 45237
rect -2348 45226 -2343 45439
rect -2325 45842 -2320 45876
rect -2317 45874 -2309 45876
rect -2076 45863 -2054 45870
rect -2325 45834 -2317 45842
rect -2060 45836 -2030 45839
rect -2325 45814 -2320 45834
rect -2317 45826 -2309 45834
rect -2060 45823 -2038 45834
rect -2033 45827 -2030 45836
rect -2028 45832 -2027 45836
rect -2068 45818 -2038 45821
rect -2325 45798 -2317 45814
rect -2325 45721 -2320 45798
rect -2309 45786 -2301 45797
rect -2317 45781 -2309 45786
rect -2309 45758 -2301 45768
rect -2251 45762 -2093 45768
rect -2317 45752 -2309 45758
rect -2124 45755 -2108 45758
rect -2060 45755 -2030 45760
rect -2000 45759 -1992 45876
rect -1846 45872 -1804 45876
rect -1663 45874 -1655 45876
rect -1846 45862 -1794 45871
rect -1912 45851 -1884 45853
rect -1852 45845 -1804 45849
rect -1844 45836 -1796 45839
rect -1671 45834 -1663 45842
rect -1844 45823 -1804 45834
rect -1663 45826 -1655 45834
rect -1852 45818 -1680 45822
rect -1844 45796 -1837 45798
rect -1789 45796 -1680 45798
rect -1837 45787 -1789 45788
rect -1655 45786 -1647 45794
rect -1837 45772 -1796 45785
rect -1663 45778 -1655 45786
rect -1796 45762 -1789 45767
rect -1837 45760 -1796 45762
rect -2000 45756 -1990 45759
rect -1844 45758 -1837 45760
rect -1655 45758 -1647 45766
rect -2124 45742 -2113 45748
rect -2325 45711 -2317 45721
rect -2325 45692 -2320 45711
rect -2317 45705 -2309 45711
rect -2243 45694 -2221 45702
rect -2211 45694 -2201 45714
rect -2073 45694 -2065 45712
rect -2000 45694 -1992 45756
rect -1844 45755 -1796 45758
rect -1837 45742 -1796 45752
rect -1663 45750 -1655 45758
rect -1671 45710 -1663 45718
rect -1655 45710 -1647 45712
rect -1663 45702 -1647 45710
rect -1642 45702 -1637 45876
rect -1885 45694 -1877 45696
rect -1708 45694 -1672 45696
rect -2243 45693 -2213 45694
rect -2325 45683 -2317 45692
rect -2259 45687 -2211 45693
rect -2183 45687 -1877 45694
rect -1869 45687 -1758 45694
rect -1710 45688 -1672 45694
rect -1710 45687 -1692 45688
rect -2211 45683 -2201 45687
rect -2325 45663 -2320 45683
rect -2317 45676 -2309 45683
rect -2211 45676 -2198 45683
rect -2325 45655 -2317 45663
rect -2300 45656 -2292 45666
rect -2243 45657 -2228 45668
rect -2211 45660 -2181 45676
rect -2211 45657 -2201 45660
rect -2325 45635 -2320 45655
rect -2317 45647 -2309 45655
rect -2325 45627 -2317 45635
rect -2325 45607 -2320 45627
rect -2317 45619 -2309 45627
rect -2325 45598 -2317 45607
rect -2325 45579 -2320 45598
rect -2317 45591 -2309 45598
rect -2325 45570 -2317 45579
rect -2325 45550 -2320 45570
rect -2317 45563 -2309 45570
rect -2325 45542 -2317 45550
rect -2290 45543 -2282 45656
rect -2251 45646 -2240 45650
rect -2211 45646 -2181 45650
rect -2251 45643 -2181 45646
rect -2176 45636 -2173 45638
rect -2240 45629 -2173 45636
rect -2169 45631 -2163 45686
rect -2073 45650 -2065 45687
rect -2073 45646 -2043 45650
rect -2000 45646 -1992 45687
rect -1915 45656 -1907 45665
rect -1963 45650 -1955 45656
rect -1963 45646 -1915 45650
rect -1885 45646 -1877 45687
rect -1875 45682 -1869 45686
rect -1829 45664 -1781 45666
rect -1847 45660 -1781 45664
rect -1778 45660 -1771 45686
rect -1758 45679 -1710 45686
rect -1718 45672 -1710 45679
rect -1768 45662 -1760 45672
rect -1718 45670 -1700 45672
rect -2146 45643 -2135 45646
rect -2105 45643 -2043 45646
rect -2035 45643 -1989 45646
rect -1973 45643 -1915 45646
rect -1907 45643 -1854 45646
rect -2073 45641 -2043 45643
rect -2135 45629 -2105 45636
rect -2065 45634 -2043 45641
rect -2243 45618 -2240 45627
rect -2221 45621 -2213 45629
rect -2211 45621 -2208 45629
rect -2203 45622 -2173 45629
rect -2251 45611 -2240 45618
rect -2211 45618 -2203 45621
rect -2211 45611 -2181 45618
rect -2073 45611 -2043 45618
rect -2203 45588 -2173 45595
rect -2262 45570 -2240 45580
rect -2203 45579 -2176 45588
rect -2083 45577 -2075 45587
rect -2040 45577 -2035 45581
rect -2073 45565 -2043 45577
rect -2028 45565 -2023 45577
rect -2000 45570 -1992 45643
rect -1963 45640 -1955 45643
rect -1963 45639 -1915 45640
rect -1955 45629 -1907 45636
rect -1885 45632 -1877 45643
rect -1837 45638 -1828 45654
rect -1758 45647 -1750 45662
rect -1758 45646 -1692 45647
rect -1837 45636 -1833 45638
rect -1837 45634 -1835 45636
rect -1887 45629 -1851 45632
rect -1750 45629 -1702 45636
rect -1885 45624 -1877 45629
rect -1963 45611 -1915 45618
rect -1905 45579 -1897 45624
rect -1857 45606 -1851 45629
rect -1760 45621 -1758 45622
rect -1837 45611 -1789 45618
rect -1758 45612 -1750 45618
rect -1758 45611 -1710 45612
rect -1955 45576 -1915 45579
rect -1963 45570 -1962 45572
rect -2000 45567 -1981 45570
rect -1965 45567 -1962 45570
rect -1955 45570 -1907 45574
rect -1885 45570 -1877 45589
rect -1857 45576 -1851 45588
rect -1750 45584 -1702 45591
rect -1829 45576 -1789 45578
rect -1766 45574 -1760 45584
rect -1829 45570 -1781 45574
rect -1756 45570 -1740 45574
rect -1680 45570 -1672 45688
rect -1671 45682 -1663 45690
rect -1645 45686 -1637 45702
rect -1663 45674 -1655 45682
rect -1671 45654 -1663 45662
rect -1663 45646 -1655 45654
rect -1671 45626 -1663 45634
rect -1671 45610 -1669 45623
rect -1663 45618 -1655 45626
rect -1671 45598 -1663 45606
rect -1663 45590 -1655 45598
rect -1671 45570 -1663 45578
rect -1955 45567 -1837 45570
rect -1829 45567 -1740 45570
rect -2206 45557 -2176 45560
rect -2206 45554 -2203 45557
rect -2161 45555 -2145 45564
rect -2073 45562 -2065 45565
rect -2073 45561 -2043 45562
rect -2028 45561 -2012 45565
rect -2073 45554 -2065 45560
rect -2203 45553 -2176 45554
rect -2065 45553 -2043 45554
rect -2262 45547 -2232 45553
rect -2176 45547 -2173 45553
rect -2043 45547 -2035 45553
rect -2325 45522 -2320 45542
rect -2317 45534 -2309 45542
rect -2153 45541 -2146 45545
rect -2325 45514 -2317 45522
rect -2300 45518 -2292 45528
rect -2325 45494 -2320 45514
rect -2317 45506 -2309 45514
rect -2325 45486 -2317 45494
rect -2325 45466 -2320 45486
rect -2317 45478 -2309 45486
rect -2290 45485 -2282 45518
rect -2273 45514 -2264 45519
rect -2206 45514 -2176 45519
rect -2262 45507 -2232 45512
rect -2198 45503 -2176 45514
rect -2198 45489 -2176 45497
rect -2166 45481 -2158 45529
rect -2143 45525 -2136 45541
rect -2143 45514 -2113 45519
rect -2073 45514 -2065 45519
rect -2065 45512 -2043 45514
rect -2043 45507 -2035 45512
rect -2065 45486 -2043 45501
rect -2006 45485 -2004 45501
rect -2265 45471 -2260 45477
rect -2143 45471 -2113 45478
rect -2270 45470 -2240 45471
rect -2270 45467 -2265 45470
rect -2325 45458 -2317 45466
rect -2325 45438 -2320 45458
rect -2317 45450 -2309 45458
rect -2113 45455 -2105 45465
rect -2291 45443 -2270 45450
rect -2198 45448 -2168 45450
rect -2135 45449 -2105 45450
rect -2103 45449 -2095 45455
rect -2113 45448 -2105 45449
rect -2065 45448 -2035 45450
rect -2000 45448 -1992 45567
rect -1963 45560 -1960 45567
rect -1915 45563 -1905 45567
rect -1963 45559 -1955 45560
rect -1963 45553 -1915 45559
rect -1989 45526 -1973 45529
rect -1915 45526 -1907 45533
rect -1990 45491 -1989 45512
rect -1983 45448 -1981 45511
rect -1885 45502 -1877 45567
rect -1789 45562 -1778 45567
rect -1837 45559 -1829 45560
rect -1837 45553 -1789 45559
rect -1756 45558 -1740 45567
rect -1837 45543 -1829 45553
rect -1872 45524 -1867 45534
rect -1789 45526 -1781 45533
rect -1776 45526 -1769 45543
rect -1756 45536 -1750 45558
rect -1671 45554 -1669 45565
rect -1663 45562 -1655 45570
rect -1671 45542 -1663 45550
rect -1663 45534 -1655 45542
rect -1702 45524 -1696 45530
rect -1955 45500 -1915 45502
rect -1963 45498 -1955 45500
rect -1963 45491 -1915 45498
rect -1963 45483 -1955 45491
rect -1963 45482 -1915 45483
rect -1973 45476 -1965 45479
rect -1955 45476 -1907 45480
rect -1974 45473 -1907 45476
rect -1973 45469 -1965 45473
rect -1963 45469 -1960 45471
rect -1963 45465 -1915 45469
rect -1963 45457 -1955 45465
rect -1963 45453 -1915 45457
rect -1963 45450 -1955 45453
rect -2240 45443 -2206 45448
rect -2198 45443 -2143 45448
rect -2113 45443 -1981 45448
rect -1915 45443 -1907 45450
rect -2270 45438 -2266 45442
rect -2086 45439 -2070 45443
rect -2325 45430 -2317 45438
rect -2270 45431 -2240 45438
rect -2206 45431 -2176 45438
rect -2325 45410 -2320 45430
rect -2317 45422 -2309 45430
rect -2270 45426 -2266 45431
rect -2270 45422 -2266 45425
rect -2198 45422 -2176 45429
rect -2166 45422 -2158 45439
rect -2143 45431 -2113 45438
rect -2198 45413 -2168 45417
rect -2325 45402 -2317 45410
rect -2143 45408 -2136 45422
rect -2085 45417 -2060 45418
rect -2039 45417 -2035 45426
rect -2135 45410 -2105 45417
rect -2085 45410 -2035 45417
rect -2029 45410 -2025 45417
rect -2325 45389 -2320 45402
rect -2317 45394 -2309 45402
rect -2235 45392 -2232 45395
rect -2325 45363 -2317 45389
rect -2325 45354 -2320 45363
rect -2325 45346 -2317 45354
rect -2135 45346 -2119 45359
rect -2000 45351 -1992 45443
rect -1983 45425 -1981 45443
rect -1955 45425 -1915 45426
rect -1862 45422 -1857 45524
rect -1706 45520 -1702 45524
rect -1829 45508 -1789 45516
rect -1671 45514 -1663 45522
rect -1849 45500 -1842 45508
rect -1790 45500 -1781 45508
rect -1663 45506 -1655 45514
rect -1837 45491 -1829 45498
rect -1758 45491 -1732 45498
rect -1748 45482 -1732 45491
rect -1671 45486 -1663 45494
rect -1829 45473 -1781 45480
rect -1663 45478 -1655 45486
rect -1829 45467 -1789 45471
rect -1768 45468 -1760 45478
rect -1758 45467 -1750 45468
rect -1671 45458 -1663 45466
rect -1837 45455 -1780 45458
rect -1758 45452 -1748 45458
rect -1708 45452 -1690 45458
rect -1829 45443 -1781 45450
rect -1680 45441 -1672 45458
rect -1663 45450 -1655 45458
rect -1829 45432 -1791 45438
rect -1758 45432 -1710 45434
rect -1758 45425 -1692 45432
rect -1671 45430 -1663 45438
rect -1955 45414 -1907 45417
rect -1791 45414 -1781 45417
rect -1991 45410 -1839 45414
rect -1791 45410 -1780 45414
rect -1680 45407 -1672 45425
rect -1663 45422 -1655 45430
rect -1839 45397 -1791 45404
rect -1671 45402 -1663 45410
rect -1829 45391 -1791 45395
rect -1671 45392 -1669 45402
rect -1663 45394 -1655 45402
rect -1680 45376 -1672 45391
rect -1642 45376 -1637 45686
rect -1619 45636 -1614 45876
rect -1619 45610 -1611 45636
rect -1768 45360 -1760 45370
rect -1758 45353 -1710 45360
rect -2325 45326 -2320 45346
rect -2317 45338 -2306 45346
rect -2031 45343 -1992 45351
rect -1750 45349 -1710 45353
rect -1674 45348 -1663 45354
rect -2307 45330 -2306 45338
rect -2149 45341 -2135 45342
rect -2149 45337 -2119 45341
rect -2024 45332 -2021 45341
rect -2325 45318 -2317 45326
rect -2325 45270 -2320 45318
rect -2317 45310 -2306 45318
rect -2185 45316 -2169 45328
rect -2056 45325 -2040 45329
rect -2021 45325 -2008 45332
rect -2056 45314 -2054 45324
rect -2056 45313 -2048 45314
rect -2307 45274 -2306 45282
rect -2111 45281 -2054 45287
rect -2325 45262 -2314 45270
rect -2104 45263 -2101 45267
rect -2325 45242 -2320 45262
rect -2314 45254 -2306 45262
rect -2104 45260 -2101 45262
rect -2084 45260 -2054 45261
rect -2000 45260 -1992 45343
rect -1758 45342 -1750 45343
rect -1758 45341 -1749 45342
rect -1758 45340 -1710 45341
rect -1663 45338 -1658 45348
rect -1831 45330 -1783 45334
rect -1784 45317 -1783 45330
rect -1674 45320 -1663 45326
rect -1826 45315 -1796 45316
rect -1663 45310 -1658 45320
rect -1654 45316 -1647 45326
rect -1644 45302 -1637 45316
rect -1758 45284 -1750 45287
rect -1758 45281 -1710 45284
rect -1844 45269 -1828 45271
rect -1844 45268 -1792 45269
rect -1828 45267 -1792 45268
rect -1772 45267 -1758 45275
rect -1750 45272 -1702 45279
rect -1750 45264 -1710 45268
rect -1700 45264 -1692 45284
rect -1674 45276 -1665 45284
rect -1674 45264 -1666 45272
rect -1758 45260 -1710 45261
rect -2307 45246 -2306 45254
rect -2139 45250 -2123 45259
rect -2111 45254 -2016 45260
rect -2139 45243 -2111 45250
rect -2325 45234 -2314 45242
rect -2177 45236 -2161 45237
rect -2141 45236 -2119 45238
rect -2104 45236 -2101 45254
rect -2076 45243 -2046 45248
rect -2325 45226 -2320 45234
rect -2314 45226 -2306 45234
rect -2076 45232 -2054 45238
rect -2021 45235 -2016 45254
rect -2000 45254 -1818 45260
rect -1802 45254 -1776 45260
rect -1760 45254 -1710 45260
rect -1666 45256 -1658 45264
rect -2189 45226 -2175 45231
rect -2373 45224 -2175 45226
rect -2373 45223 -2359 45224
rect -2371 45086 -2366 45223
rect -2348 45171 -2343 45224
rect -2325 45214 -2320 45224
rect -2307 45218 -2306 45224
rect -2189 45223 -2175 45224
rect -2149 45222 -2119 45231
rect -2084 45230 -2036 45231
rect -2000 45230 -1992 45254
rect -1758 45252 -1710 45254
rect -1758 45250 -1755 45252
rect -1828 45243 -1792 45250
rect -1768 45241 -1760 45248
rect -1758 45243 -1757 45250
rect -1710 45249 -1702 45250
rect -1750 45243 -1702 45249
rect -1674 45248 -1665 45256
rect -1768 45238 -1764 45241
rect -1758 45238 -1755 45243
rect -1818 45230 -1789 45238
rect -1758 45231 -1754 45238
rect -1750 45233 -1710 45238
rect -1674 45236 -1666 45244
rect -1758 45230 -1692 45231
rect -2084 45228 -1692 45230
rect -1666 45228 -1658 45236
rect -2084 45225 -1690 45228
rect -2084 45222 -2054 45225
rect -2046 45223 -1710 45225
rect -2325 45206 -2314 45214
rect -2076 45213 -2046 45220
rect -2325 45186 -2320 45206
rect -2314 45198 -2306 45206
rect -2076 45205 -2054 45211
rect -2084 45201 -2054 45203
rect -2104 45198 -2054 45201
rect -2307 45190 -2306 45198
rect -2084 45195 -2054 45198
rect -2325 45172 -2314 45186
rect -2348 45147 -2341 45171
rect -2325 45156 -2320 45172
rect -2314 45170 -2309 45172
rect -2309 45158 -2298 45170
rect -2092 45167 -2060 45168
rect -2062 45162 -2060 45167
rect -2314 45156 -2309 45158
rect -2348 45086 -2343 45147
rect -2325 45144 -2314 45156
rect -2076 45152 -2062 45162
rect -2076 45146 -2046 45150
rect -2014 45149 -2003 45158
rect -2062 45144 -2046 45146
rect -2325 45128 -2320 45144
rect -2314 45142 -2309 45144
rect -2076 45143 -2062 45144
rect -2309 45130 -2298 45142
rect -2092 45137 -2076 45143
rect -2046 45137 -2026 45138
rect -2314 45128 -2309 45130
rect -2046 45128 -2042 45129
rect -2325 45116 -2314 45128
rect -2141 45124 -2134 45126
rect -2052 45124 -2046 45128
rect -2292 45119 -2111 45124
rect -2096 45122 -2046 45124
rect -2076 45119 -2046 45122
rect -2325 45086 -2320 45116
rect -2314 45114 -2309 45116
rect -2092 45102 -2062 45104
rect -2094 45098 -2062 45102
rect -2000 45086 -1992 45223
rect -1758 45222 -1710 45223
rect -1680 45220 -1665 45228
rect -1750 45213 -1702 45220
rect -1680 45216 -1672 45220
rect -1680 45211 -1666 45216
rect -1836 45207 -1820 45208
rect -1837 45203 -1820 45207
rect -1750 45205 -1710 45211
rect -1674 45208 -1666 45211
rect -1837 45196 -1789 45203
rect -1758 45202 -1710 45203
rect -1760 45199 -1692 45202
rect -1666 45200 -1658 45208
rect -1837 45195 -1820 45196
rect -1764 45195 -1692 45199
rect -1674 45195 -1665 45200
rect -1680 45192 -1665 45195
rect -1750 45176 -1702 45178
rect -1680 45168 -1672 45192
rect -1671 45172 -1666 45188
rect -1854 45167 -1806 45168
rect -1829 45152 -1806 45162
rect -1655 45160 -1650 45172
rect -1666 45156 -1655 45160
rect -1829 45146 -1798 45150
rect -1680 45149 -1672 45152
rect -1806 45144 -1798 45146
rect -1671 45144 -1666 45156
rect -1829 45143 -1806 45144
rect -1854 45141 -1829 45143
rect -1854 45137 -1806 45141
rect -1829 45125 -1806 45135
rect -1655 45132 -1650 45144
rect -1666 45128 -1655 45132
rect -1829 45119 -1680 45124
rect -1671 45116 -1666 45128
rect -1854 45102 -1806 45104
rect -1854 45098 -1680 45102
rect -1642 45086 -1637 45302
rect -1619 45300 -1614 45610
rect -1619 45226 -1612 45250
rect -1619 45086 -1614 45226
rect -1530 45086 -1526 45876
rect -1506 45086 -1502 45876
rect -1482 45086 -1478 45876
rect -1458 45086 -1454 45876
rect -1434 45086 -1430 45876
rect -1410 45207 -1406 45876
rect -1421 45206 -1387 45207
rect -1386 45206 -1382 45876
rect -1362 45206 -1358 45876
rect -1338 45206 -1334 45876
rect -1314 45206 -1310 45876
rect -1290 45206 -1286 45876
rect -1266 45206 -1262 45876
rect -1242 45206 -1238 45876
rect -1218 45206 -1214 45876
rect -1194 45206 -1190 45876
rect -1170 45206 -1166 45876
rect -1146 45206 -1142 45876
rect -1122 45206 -1118 45876
rect -1098 45206 -1094 45876
rect -1074 45206 -1070 45876
rect -1050 45206 -1046 45876
rect -1026 45206 -1022 45876
rect -1002 45206 -998 45876
rect -978 45206 -974 45876
rect -954 45206 -950 45876
rect -930 45206 -926 45876
rect -917 45845 -912 45855
rect -906 45845 -902 45876
rect -907 45831 -902 45845
rect -906 45206 -902 45831
rect -882 45779 -878 45876
rect -869 45869 -864 45876
rect -859 45855 -854 45869
rect -882 45755 -875 45779
rect -882 45206 -878 45755
rect -858 45206 -854 45855
rect -834 45827 -830 45899
rect -834 45779 -827 45827
rect -834 45206 -830 45779
rect -810 45206 -806 45903
rect -786 45875 -782 46140
rect -762 45927 -758 46140
rect -773 45926 -739 45927
rect -738 45926 -734 46140
rect -714 45926 -710 46140
rect -690 45926 -686 46140
rect -666 45926 -662 46140
rect -642 45926 -638 46140
rect -618 46047 -614 46140
rect -629 46046 -595 46047
rect -594 46046 -590 46140
rect -570 46046 -566 46140
rect -546 46046 -542 46140
rect -522 46046 -518 46140
rect -515 46139 -501 46140
rect -509 46133 -504 46139
rect -499 46119 -494 46133
rect -498 46046 -494 46119
rect -485 46046 -477 46047
rect -629 46044 -477 46046
rect -629 46037 -624 46044
rect -618 46037 -614 46044
rect -619 46023 -614 46037
rect -629 46013 -624 46023
rect -619 45999 -614 46013
rect -618 45926 -614 45999
rect -594 45971 -590 46044
rect -594 45950 -587 45971
rect -570 45950 -566 46044
rect -546 45950 -542 46044
rect -533 45965 -528 45975
rect -522 45965 -518 46044
rect -523 45951 -518 45965
rect -522 45950 -518 45951
rect -498 45950 -494 46044
rect -491 46043 -477 46044
rect -485 46037 -480 46043
rect -475 46023 -470 46037
rect -474 45950 -470 46023
rect -461 45950 -453 45951
rect -611 45948 -453 45950
rect -611 45947 -597 45948
rect -773 45924 -597 45926
rect -773 45917 -768 45924
rect -762 45917 -758 45924
rect -763 45903 -758 45917
rect -773 45893 -768 45903
rect -763 45879 -758 45893
rect -786 45827 -779 45875
rect -786 45206 -782 45827
rect -762 45206 -758 45879
rect -738 45851 -734 45924
rect -738 45803 -731 45851
rect -738 45206 -734 45803
rect -714 45206 -710 45924
rect -690 45206 -686 45924
rect -666 45206 -662 45924
rect -653 45725 -648 45735
rect -642 45725 -638 45924
rect -643 45711 -638 45725
rect -653 45701 -648 45711
rect -643 45687 -638 45701
rect -642 45206 -638 45687
rect -618 45659 -614 45924
rect -611 45923 -597 45924
rect -594 45923 -587 45948
rect -618 45611 -611 45659
rect -618 45206 -614 45611
rect -594 45206 -590 45923
rect -570 45206 -566 45948
rect -546 45206 -542 45948
rect -522 45206 -518 45948
rect -498 45899 -494 45948
rect -498 45875 -491 45899
rect -498 45206 -494 45875
rect -474 45206 -470 45948
rect -467 45947 -453 45948
rect -461 45941 -456 45947
rect -451 45927 -446 45941
rect -450 45206 -446 45927
rect -426 45851 -419 45875
rect -426 45206 -422 45851
rect -413 45725 -408 45735
rect -403 45711 -398 45725
rect -413 45293 -408 45303
rect -402 45293 -398 45711
rect -403 45279 -398 45293
rect -413 45206 -381 45207
rect -1421 45204 -381 45206
rect -1421 45197 -1416 45204
rect -1410 45197 -1406 45204
rect -1411 45183 -1406 45197
rect -1421 45173 -1416 45183
rect -1411 45159 -1406 45173
rect -1410 45086 -1406 45159
rect -1386 45131 -1382 45204
rect -2393 45084 -1389 45086
rect -2371 45062 -2366 45084
rect -2348 45062 -2343 45084
rect -2325 45062 -2320 45084
rect -2072 45082 -2036 45083
rect -2072 45076 -2054 45082
rect -2309 45068 -2301 45076
rect -2317 45062 -2309 45068
rect -2092 45067 -2062 45072
rect -2000 45063 -1992 45084
rect -1938 45083 -1906 45084
rect -1920 45082 -1906 45083
rect -1806 45076 -1680 45082
rect -1854 45067 -1806 45072
rect -1655 45068 -1647 45076
rect -1982 45063 -1966 45064
rect -2000 45062 -1966 45063
rect -1846 45062 -1806 45065
rect -1663 45062 -1655 45068
rect -1642 45062 -1637 45084
rect -1619 45062 -1614 45084
rect -1554 45070 -1547 45083
rect -1589 45062 -1555 45063
rect -2393 45060 -1555 45062
rect -2371 45038 -2366 45060
rect -2348 45038 -2343 45060
rect -2325 45038 -2320 45060
rect -2000 45058 -1966 45060
rect -2309 45040 -2301 45048
rect -2062 45047 -2054 45054
rect -2092 45040 -2084 45047
rect -2062 45040 -2026 45042
rect -2317 45038 -2309 45040
rect -2062 45038 -2012 45040
rect -2000 45038 -1992 45058
rect -1982 45057 -1966 45058
rect -1846 45056 -1806 45060
rect -1846 45049 -1798 45054
rect -1806 45047 -1798 45049
rect -1854 45045 -1846 45047
rect -1854 45040 -1806 45045
rect -1655 45040 -1647 45048
rect -1864 45038 -1796 45039
rect -1663 45038 -1655 45040
rect -1642 45038 -1637 45060
rect -1619 45038 -1614 45060
rect -1571 45059 -1557 45060
rect -1554 45059 -1547 45060
rect -1530 45038 -1526 45084
rect -1506 45038 -1502 45084
rect -1482 45038 -1478 45084
rect -1458 45038 -1454 45084
rect -1434 45038 -1430 45084
rect -1410 45038 -1406 45084
rect -1403 45083 -1389 45084
rect -1386 45083 -1379 45131
rect -1386 45038 -1382 45083
rect -1362 45038 -1358 45204
rect -1338 45038 -1334 45204
rect -1314 45111 -1310 45204
rect -1325 45110 -1291 45111
rect -1290 45110 -1286 45204
rect -1266 45110 -1262 45204
rect -1242 45110 -1238 45204
rect -1218 45110 -1214 45204
rect -1194 45110 -1190 45204
rect -1170 45110 -1166 45204
rect -1146 45110 -1142 45204
rect -1122 45110 -1118 45204
rect -1098 45110 -1094 45204
rect -1074 45110 -1070 45204
rect -1050 45110 -1046 45204
rect -1026 45110 -1022 45204
rect -1002 45110 -998 45204
rect -978 45110 -974 45204
rect -954 45110 -950 45204
rect -930 45110 -926 45204
rect -906 45110 -902 45204
rect -882 45110 -878 45204
rect -858 45110 -854 45204
rect -834 45110 -830 45204
rect -810 45110 -806 45204
rect -786 45110 -782 45204
rect -762 45110 -758 45204
rect -738 45110 -734 45204
rect -714 45110 -710 45204
rect -690 45110 -686 45204
rect -666 45110 -662 45204
rect -642 45110 -638 45204
rect -618 45110 -614 45204
rect -594 45110 -590 45204
rect -570 45110 -566 45204
rect -546 45110 -542 45204
rect -522 45110 -518 45204
rect -498 45110 -494 45204
rect -474 45110 -470 45204
rect -461 45125 -456 45135
rect -450 45125 -446 45204
rect -451 45111 -446 45125
rect -450 45110 -446 45111
rect -426 45110 -422 45204
rect -413 45197 -408 45204
rect -395 45203 -381 45204
rect -403 45183 -398 45197
rect -402 45110 -398 45183
rect -389 45110 -381 45111
rect -1325 45108 -381 45110
rect -1325 45101 -1320 45108
rect -1314 45101 -1310 45108
rect -1315 45087 -1310 45101
rect -1325 45077 -1320 45087
rect -1315 45063 -1310 45077
rect -1314 45038 -1310 45063
rect -1290 45038 -1286 45108
rect -1266 45038 -1262 45108
rect -1242 45038 -1238 45108
rect -1218 45038 -1214 45108
rect -1194 45038 -1190 45108
rect -1170 45038 -1166 45108
rect -1146 45038 -1142 45108
rect -1122 45038 -1118 45108
rect -1098 45038 -1094 45108
rect -1074 45038 -1070 45108
rect -1050 45038 -1046 45108
rect -1026 45038 -1022 45108
rect -1002 45038 -998 45108
rect -978 45038 -974 45108
rect -954 45038 -950 45108
rect -930 45038 -926 45108
rect -906 45038 -902 45108
rect -882 45038 -878 45108
rect -858 45038 -854 45108
rect -834 45038 -830 45108
rect -810 45038 -806 45108
rect -786 45038 -782 45108
rect -762 45038 -758 45108
rect -738 45038 -734 45108
rect -714 45038 -710 45108
rect -690 45038 -686 45108
rect -666 45038 -662 45108
rect -642 45038 -638 45108
rect -618 45038 -614 45108
rect -594 45038 -590 45108
rect -570 45038 -566 45108
rect -546 45038 -542 45108
rect -522 45038 -518 45108
rect -498 45038 -494 45108
rect -474 45038 -470 45108
rect -450 45038 -446 45108
rect -426 45059 -422 45108
rect -2393 45036 -429 45038
rect -2371 44990 -2366 45036
rect -2348 44990 -2343 45036
rect -2325 44990 -2320 45036
rect -2317 45032 -2309 45036
rect -2062 45032 -2054 45036
rect -2154 45028 -2138 45030
rect -2057 45028 -2054 45032
rect -2292 45022 -2054 45028
rect -2052 45022 -2044 45032
rect -2092 45006 -2062 45008
rect -2094 45002 -2062 45006
rect -2000 44990 -1992 45036
rect -1846 45029 -1806 45036
rect -1663 45032 -1655 45036
rect -1846 45022 -1680 45028
rect -1854 45006 -1806 45008
rect -1854 45002 -1680 45006
rect -1642 44990 -1637 45036
rect -1619 44990 -1614 45036
rect -1530 44990 -1526 45036
rect -1506 44990 -1502 45036
rect -1482 44990 -1478 45036
rect -1458 44990 -1454 45036
rect -1434 44990 -1430 45036
rect -1410 44990 -1406 45036
rect -1386 44990 -1382 45036
rect -1362 44990 -1358 45036
rect -1338 44990 -1334 45036
rect -1314 44990 -1310 45036
rect -1290 45035 -1286 45036
rect -2393 44988 -1293 44990
rect -2371 44966 -2366 44988
rect -2348 44966 -2343 44988
rect -2325 44966 -2320 44988
rect -2072 44986 -2036 44987
rect -2072 44980 -2054 44986
rect -2309 44972 -2301 44980
rect -2317 44966 -2309 44972
rect -2092 44971 -2062 44976
rect -2000 44967 -1992 44988
rect -1938 44987 -1906 44988
rect -1920 44986 -1906 44987
rect -1806 44980 -1680 44986
rect -1854 44971 -1806 44976
rect -1655 44972 -1647 44980
rect -1982 44967 -1966 44968
rect -2000 44966 -1966 44967
rect -1846 44966 -1806 44969
rect -1663 44966 -1655 44972
rect -1642 44966 -1637 44988
rect -1619 44966 -1614 44988
rect -1554 44974 -1547 44987
rect -2393 44964 -1557 44966
rect -2371 44942 -2366 44964
rect -2348 44942 -2343 44964
rect -2325 44942 -2320 44964
rect -2000 44962 -1966 44964
rect -2309 44944 -2301 44952
rect -2062 44951 -2054 44958
rect -2092 44944 -2084 44951
rect -2062 44944 -2026 44946
rect -2317 44942 -2309 44944
rect -2062 44942 -2012 44944
rect -2000 44942 -1992 44962
rect -1982 44961 -1966 44962
rect -1846 44960 -1806 44964
rect -1846 44953 -1798 44958
rect -1806 44951 -1798 44953
rect -1854 44949 -1846 44951
rect -1854 44944 -1806 44949
rect -1655 44944 -1647 44952
rect -1864 44942 -1796 44943
rect -1663 44942 -1655 44944
rect -1642 44942 -1637 44964
rect -1619 44942 -1614 44964
rect -1571 44963 -1557 44964
rect -1554 44963 -1547 44964
rect -1530 44942 -1526 44988
rect -1506 44942 -1502 44988
rect -1482 44942 -1478 44988
rect -1458 44942 -1454 44988
rect -1434 44942 -1430 44988
rect -1410 44942 -1406 44988
rect -1386 44942 -1382 44988
rect -1362 44942 -1358 44988
rect -1338 44942 -1334 44988
rect -1314 44942 -1310 44988
rect -1307 44987 -1293 44988
rect -1290 44987 -1283 45035
rect -1290 44942 -1286 44987
rect -1266 44942 -1262 45036
rect -1242 44942 -1238 45036
rect -1218 44942 -1214 45036
rect -1194 44942 -1190 45036
rect -1170 44942 -1166 45036
rect -1146 44942 -1142 45036
rect -1122 44942 -1118 45036
rect -1098 44942 -1094 45036
rect -1074 45015 -1070 45036
rect -1085 45014 -1051 45015
rect -1050 45014 -1046 45036
rect -1026 45014 -1022 45036
rect -1002 45014 -998 45036
rect -978 45014 -974 45036
rect -954 45014 -950 45036
rect -930 45014 -926 45036
rect -906 45014 -902 45036
rect -882 45014 -878 45036
rect -858 45014 -854 45036
rect -834 45014 -830 45036
rect -810 45014 -806 45036
rect -786 45014 -782 45036
rect -762 45014 -758 45036
rect -738 45014 -734 45036
rect -714 45014 -710 45036
rect -690 45014 -686 45036
rect -666 45014 -662 45036
rect -642 45014 -638 45036
rect -618 45014 -614 45036
rect -594 45014 -590 45036
rect -570 45014 -566 45036
rect -546 45014 -542 45036
rect -522 45014 -518 45036
rect -498 45014 -494 45036
rect -474 45014 -470 45036
rect -450 45014 -446 45036
rect -443 45035 -429 45036
rect -426 45035 -419 45059
rect -426 45014 -422 45035
rect -413 45029 -408 45039
rect -402 45029 -398 45108
rect -395 45107 -381 45108
rect -389 45101 -384 45107
rect -379 45087 -374 45101
rect -403 45015 -398 45029
rect -402 45014 -398 45015
rect -378 45014 -374 45087
rect -365 45014 -357 45015
rect -1085 45012 -357 45014
rect -1085 45005 -1080 45012
rect -1074 45005 -1070 45012
rect -1075 44991 -1070 45005
rect -1085 44981 -1080 44991
rect -1075 44967 -1070 44981
rect -1074 44942 -1070 44967
rect -1061 44957 -1056 44967
rect -1050 44957 -1046 45012
rect -1051 44943 -1046 44957
rect -1026 44943 -1022 45012
rect -1050 44942 -1046 44943
rect -1037 44942 -1003 44943
rect -2393 44940 -1003 44942
rect -2371 44870 -2366 44940
rect -2348 44870 -2343 44940
rect -2325 44870 -2320 44940
rect -2317 44936 -2309 44940
rect -2062 44936 -2054 44940
rect -2154 44932 -2138 44934
rect -2057 44932 -2054 44936
rect -2292 44926 -2054 44932
rect -2052 44926 -2044 44936
rect -2092 44910 -2062 44912
rect -2094 44906 -2062 44910
rect -2309 44876 -2301 44882
rect -2317 44870 -2309 44876
rect -2000 44870 -1992 44940
rect -1846 44933 -1806 44940
rect -1663 44936 -1655 44940
rect -1846 44926 -1680 44932
rect -1854 44910 -1806 44912
rect -1854 44906 -1680 44910
rect -1655 44876 -1647 44882
rect -1663 44870 -1655 44876
rect -1642 44870 -1637 44940
rect -1619 44870 -1614 44940
rect -1530 44870 -1526 44940
rect -1506 44870 -1502 44940
rect -1482 44870 -1478 44940
rect -1458 44870 -1454 44940
rect -1434 44870 -1430 44940
rect -1410 44870 -1406 44940
rect -1386 44870 -1382 44940
rect -1362 44870 -1358 44940
rect -1338 44870 -1334 44940
rect -1314 44870 -1310 44940
rect -1290 44870 -1286 44940
rect -1266 44870 -1262 44940
rect -1242 44870 -1238 44940
rect -1218 44870 -1214 44940
rect -1194 44895 -1190 44940
rect -1205 44894 -1171 44895
rect -1170 44894 -1166 44940
rect -1146 44894 -1142 44940
rect -1122 44894 -1118 44940
rect -1098 44894 -1094 44940
rect -1074 44894 -1070 44940
rect -1050 44939 -1046 44940
rect -1205 44892 -1053 44894
rect -1205 44885 -1200 44892
rect -1194 44885 -1190 44892
rect -1195 44871 -1190 44885
rect -1205 44870 -1171 44871
rect -2393 44868 -1171 44870
rect -2371 44774 -2366 44868
rect -2348 44774 -2343 44868
rect -2325 44806 -2320 44868
rect -2317 44866 -2309 44868
rect -2000 44867 -1966 44868
rect -2000 44866 -1982 44867
rect -1663 44866 -1655 44868
rect -2028 44858 -2018 44860
rect -2309 44848 -2301 44854
rect -2091 44848 -2061 44855
rect -2317 44838 -2309 44848
rect -2044 44846 -2028 44848
rect -2026 44846 -2014 44858
rect -2084 44840 -2061 44846
rect -2044 44844 -2014 44846
rect -2292 44830 -2054 44839
rect -2325 44798 -2317 44806
rect -2325 44778 -2320 44798
rect -2317 44790 -2309 44798
rect -2325 44774 -2317 44778
rect -2000 44774 -1992 44866
rect -1982 44865 -1966 44866
rect -1980 44848 -1932 44855
rect -1655 44848 -1647 44854
rect -1846 44830 -1680 44839
rect -1663 44838 -1655 44848
rect -1671 44798 -1663 44806
rect -1663 44790 -1655 44798
rect -1671 44774 -1663 44778
rect -1642 44774 -1637 44868
rect -1619 44774 -1614 44868
rect -1530 44774 -1526 44868
rect -1506 44774 -1502 44868
rect -1482 44774 -1478 44868
rect -1458 44774 -1454 44868
rect -1434 44774 -1430 44868
rect -1410 44774 -1406 44868
rect -1386 44774 -1382 44868
rect -1362 44774 -1358 44868
rect -1338 44774 -1334 44868
rect -1314 44774 -1310 44868
rect -1290 44774 -1286 44868
rect -1266 44774 -1262 44868
rect -1242 44774 -1238 44868
rect -1218 44774 -1214 44868
rect -1205 44861 -1200 44868
rect -1195 44847 -1190 44861
rect -1194 44774 -1190 44847
rect -1170 44819 -1166 44892
rect -2393 44772 -1173 44774
rect -2371 44726 -2366 44772
rect -2348 44726 -2343 44772
rect -2325 44766 -2317 44772
rect -2018 44770 -2004 44772
rect -2325 44750 -2320 44766
rect -2317 44762 -2309 44766
rect -2069 44764 -2053 44766
rect -2309 44750 -2301 44762
rect -2096 44753 -2095 44759
rect -2000 44754 -1992 44772
rect -1671 44766 -1663 44772
rect -1663 44762 -1655 44766
rect -1977 44755 -1929 44761
rect -2112 44750 -2095 44753
rect -2325 44738 -2317 44750
rect -2325 44726 -2320 44738
rect -2317 44734 -2309 44738
rect -2112 44737 -2096 44750
rect -2059 44746 -2053 44753
rect -2027 44752 -1992 44754
rect -2059 44742 -2045 44746
rect -2018 44744 -2017 44746
rect -2083 44737 -2053 44738
rect -2019 44736 -2017 44740
rect -2309 44726 -2301 44734
rect -2017 44730 -2009 44736
rect -2000 44730 -1992 44752
rect -1972 44738 -1929 44753
rect -1655 44750 -1647 44762
rect -1671 44738 -1663 44750
rect -1972 44737 -1924 44738
rect -1663 44734 -1655 44738
rect -2033 44726 -1992 44730
rect -1655 44726 -1647 44734
rect -1642 44726 -1637 44772
rect -1619 44726 -1614 44772
rect -1530 44726 -1526 44772
rect -1506 44726 -1502 44772
rect -1482 44726 -1478 44772
rect -1458 44726 -1454 44772
rect -1434 44726 -1430 44772
rect -1410 44726 -1406 44772
rect -1386 44726 -1382 44772
rect -1362 44726 -1358 44772
rect -1338 44726 -1334 44772
rect -1314 44726 -1310 44772
rect -1290 44726 -1286 44772
rect -1266 44726 -1262 44772
rect -1242 44726 -1238 44772
rect -1218 44726 -1214 44772
rect -1194 44726 -1190 44772
rect -1187 44771 -1173 44772
rect -1170 44771 -1163 44819
rect -1170 44726 -1166 44771
rect -1146 44726 -1142 44892
rect -1122 44726 -1118 44892
rect -1098 44726 -1094 44892
rect -1074 44726 -1070 44892
rect -1067 44891 -1053 44892
rect -1050 44891 -1043 44939
rect -1037 44933 -1032 44940
rect -1026 44933 -1022 44940
rect -1027 44919 -1022 44933
rect -1026 44891 -1022 44919
rect -1050 44726 -1046 44891
rect -1026 44867 -1019 44891
rect -1002 44867 -998 45012
rect -1026 44726 -1022 44867
rect -1002 44843 -995 44867
rect -1002 44726 -998 44843
rect -978 44726 -974 45012
rect -954 44726 -950 45012
rect -930 44726 -926 45012
rect -906 44726 -902 45012
rect -882 44799 -878 45012
rect -893 44798 -859 44799
rect -858 44798 -854 45012
rect -834 44798 -830 45012
rect -810 44798 -806 45012
rect -786 44798 -782 45012
rect -762 44798 -758 45012
rect -738 44798 -734 45012
rect -714 44798 -710 45012
rect -690 44798 -686 45012
rect -677 44813 -672 44823
rect -666 44813 -662 45012
rect -667 44799 -662 44813
rect -666 44798 -662 44799
rect -642 44798 -638 45012
rect -618 44798 -614 45012
rect -594 44798 -590 45012
rect -570 44798 -566 45012
rect -546 44798 -542 45012
rect -522 44798 -518 45012
rect -498 44798 -494 45012
rect -474 44798 -470 45012
rect -450 44798 -446 45012
rect -426 44798 -422 45012
rect -402 44798 -398 45012
rect -378 44963 -374 45012
rect -371 45011 -357 45012
rect -365 45005 -360 45011
rect -355 44991 -350 45005
rect -378 44939 -371 44963
rect -378 44798 -374 44939
rect -354 44798 -350 44991
rect -341 44885 -336 44895
rect -331 44871 -326 44885
rect -330 44798 -326 44871
rect -317 44798 -309 44799
rect -893 44796 -309 44798
rect -893 44789 -888 44796
rect -882 44789 -878 44796
rect -883 44775 -878 44789
rect -893 44765 -888 44775
rect -883 44751 -878 44765
rect -882 44726 -878 44751
rect -858 44726 -854 44796
rect -834 44726 -830 44796
rect -810 44726 -806 44796
rect -786 44726 -782 44796
rect -762 44726 -758 44796
rect -738 44726 -734 44796
rect -714 44726 -710 44796
rect -690 44726 -686 44796
rect -666 44726 -662 44796
rect -642 44747 -638 44796
rect -2393 44724 -645 44726
rect -2371 44606 -2366 44724
rect -2348 44606 -2343 44724
rect -2325 44722 -2320 44724
rect -2309 44722 -2301 44724
rect -2325 44710 -2317 44722
rect -2325 44690 -2320 44710
rect -2317 44706 -2309 44710
rect -2325 44682 -2317 44690
rect -2325 44662 -2320 44682
rect -2317 44674 -2309 44682
rect -2117 44673 -2095 44683
rect -2045 44680 -2037 44694
rect -2325 44646 -2317 44662
rect -2325 44630 -2320 44646
rect -2309 44634 -2301 44646
rect -2317 44630 -2309 44634
rect -2117 44632 -2095 44639
rect -2069 44638 -2041 44646
rect -2017 44644 -2015 44646
rect -2325 44618 -2317 44630
rect -2125 44623 -2095 44630
rect -2047 44628 -2011 44630
rect -2059 44626 -2011 44628
rect -2000 44626 -1992 44724
rect -1655 44722 -1647 44724
rect -1671 44710 -1663 44722
rect -1663 44706 -1655 44710
rect -1969 44673 -1929 44685
rect -1671 44682 -1663 44690
rect -1663 44674 -1655 44682
rect -1671 44646 -1663 44662
rect -1655 44634 -1647 44646
rect -1663 44630 -1655 44634
rect -2125 44621 -2117 44623
rect -2059 44622 -2045 44626
rect -2021 44623 -1992 44626
rect -1977 44623 -1929 44630
rect -2325 44606 -2320 44618
rect -2309 44606 -2301 44618
rect -2131 44613 -2129 44618
rect -2125 44615 -2095 44621
rect -2021 44616 -2009 44620
rect -2125 44613 -2117 44615
rect -2133 44606 -2129 44613
rect -2117 44606 -2087 44613
rect -2025 44610 -2021 44616
rect -2000 44610 -1992 44623
rect -1969 44615 -1929 44621
rect -1671 44618 -1663 44630
rect -2033 44606 -1992 44610
rect -1969 44606 -1921 44613
rect -1655 44606 -1647 44618
rect -1642 44606 -1637 44724
rect -1619 44606 -1614 44724
rect -1530 44606 -1526 44724
rect -1506 44606 -1502 44724
rect -1493 44693 -1488 44703
rect -1482 44693 -1478 44724
rect -1483 44679 -1478 44693
rect -1482 44606 -1478 44679
rect -1458 44627 -1454 44724
rect -2393 44604 -1461 44606
rect -2371 44510 -2366 44604
rect -2348 44510 -2343 44604
rect -2325 44602 -2320 44604
rect -2317 44602 -2309 44604
rect -2131 44602 -2129 44604
rect -2125 44602 -2095 44604
rect -2325 44590 -2317 44602
rect -2117 44597 -2095 44602
rect -2325 44570 -2320 44590
rect -2325 44562 -2317 44570
rect -2325 44510 -2320 44562
rect -2317 44554 -2309 44562
rect -2117 44553 -2095 44563
rect -2045 44560 -2037 44574
rect -2309 44514 -2301 44524
rect -2087 44520 -2076 44528
rect -2017 44524 -2015 44531
rect -2317 44510 -2309 44514
rect -2092 44512 -2087 44520
rect -2092 44510 -2077 44511
rect -2000 44510 -1992 44604
rect -1663 44602 -1655 44604
rect -1671 44590 -1663 44602
rect -1969 44553 -1929 44565
rect -1671 44562 -1663 44570
rect -1663 44554 -1655 44562
rect -1655 44514 -1647 44524
rect -1928 44510 -1924 44511
rect -1854 44510 -1680 44511
rect -1663 44510 -1655 44514
rect -1642 44510 -1637 44604
rect -1619 44510 -1614 44604
rect -1530 44510 -1526 44604
rect -1506 44510 -1502 44604
rect -1482 44510 -1478 44604
rect -1475 44603 -1461 44604
rect -1458 44603 -1451 44627
rect -1458 44510 -1454 44603
rect -1445 44573 -1440 44583
rect -1434 44573 -1430 44724
rect -1435 44559 -1430 44573
rect -1434 44511 -1430 44559
rect -1445 44510 -1411 44511
rect -2393 44508 -1411 44510
rect -2371 44486 -2366 44508
rect -2348 44486 -2343 44508
rect -2325 44486 -2320 44508
rect -2092 44503 -2037 44508
rect -2021 44503 -1969 44508
rect -1921 44503 -1913 44508
rect -1854 44504 -1680 44508
rect -2100 44501 -2092 44502
rect -2309 44486 -2301 44496
rect -2100 44495 -2087 44501
rect -2051 44488 -2026 44490
rect -2062 44486 -2012 44488
rect -2000 44486 -1992 44503
rect -1969 44495 -1921 44502
rect -1969 44486 -1964 44495
rect -1864 44486 -1796 44487
rect -1655 44486 -1647 44496
rect -1642 44486 -1637 44508
rect -1619 44486 -1614 44508
rect -1530 44486 -1526 44508
rect -1506 44486 -1502 44508
rect -1482 44486 -1478 44508
rect -1458 44486 -1454 44508
rect -1445 44501 -1440 44508
rect -1434 44501 -1430 44508
rect -1410 44507 -1406 44724
rect -1435 44487 -1430 44501
rect -1421 44497 -1413 44501
rect -1427 44487 -1421 44497
rect -1434 44486 -1430 44487
rect -2393 44484 -1413 44486
rect -2371 44414 -2366 44484
rect -2348 44414 -2343 44484
rect -2325 44414 -2320 44484
rect -2317 44480 -2309 44484
rect -2105 44477 -2092 44480
rect -2092 44454 -2062 44456
rect -2094 44450 -2062 44454
rect -2309 44420 -2301 44426
rect -2317 44414 -2309 44420
rect -2000 44414 -1992 44484
rect -1663 44480 -1655 44484
rect -1969 44477 -1921 44480
rect -1854 44454 -1806 44456
rect -1854 44450 -1680 44454
rect -1655 44420 -1647 44426
rect -1663 44414 -1655 44420
rect -1642 44414 -1637 44484
rect -1619 44414 -1614 44484
rect -1530 44414 -1526 44484
rect -1506 44414 -1502 44484
rect -1482 44414 -1478 44484
rect -1458 44414 -1454 44484
rect -1434 44414 -1430 44484
rect -1427 44483 -1413 44484
rect -1410 44483 -1403 44507
rect -1410 44435 -1406 44483
rect -1397 44477 -1392 44487
rect -1386 44477 -1382 44724
rect -1387 44463 -1382 44477
rect -2393 44412 -1413 44414
rect -2371 44318 -2366 44412
rect -2348 44318 -2343 44412
rect -2325 44350 -2320 44412
rect -2317 44410 -2309 44412
rect -2000 44411 -1966 44412
rect -2000 44410 -1982 44411
rect -1663 44410 -1655 44412
rect -2028 44402 -2018 44404
rect -2309 44392 -2301 44398
rect -2091 44392 -2061 44399
rect -2317 44382 -2309 44392
rect -2044 44390 -2028 44392
rect -2026 44390 -2014 44402
rect -2084 44384 -2061 44390
rect -2044 44388 -2014 44390
rect -2292 44374 -2054 44383
rect -2325 44342 -2317 44350
rect -2325 44322 -2320 44342
rect -2317 44334 -2309 44342
rect -2325 44318 -2317 44322
rect -2000 44318 -1992 44410
rect -1982 44409 -1966 44410
rect -1980 44392 -1932 44399
rect -1655 44392 -1647 44398
rect -1846 44374 -1680 44383
rect -1663 44382 -1655 44392
rect -1671 44342 -1663 44350
rect -1663 44334 -1655 44342
rect -1671 44318 -1663 44322
rect -1642 44318 -1637 44412
rect -1619 44318 -1614 44412
rect -1530 44318 -1526 44412
rect -1506 44318 -1502 44412
rect -1482 44318 -1478 44412
rect -1458 44318 -1454 44412
rect -1434 44318 -1430 44412
rect -1427 44411 -1413 44412
rect -1410 44411 -1403 44435
rect -1410 44318 -1406 44411
rect -1386 44318 -1382 44463
rect -1362 44411 -1358 44724
rect -1362 44387 -1355 44411
rect -1362 44318 -1358 44387
rect -1338 44318 -1334 44724
rect -1314 44318 -1310 44724
rect -1290 44318 -1286 44724
rect -1266 44318 -1262 44724
rect -1242 44318 -1238 44724
rect -1218 44318 -1214 44724
rect -1194 44318 -1190 44724
rect -1170 44318 -1166 44724
rect -1146 44318 -1142 44724
rect -1122 44318 -1118 44724
rect -1098 44318 -1094 44724
rect -1074 44318 -1070 44724
rect -1050 44318 -1046 44724
rect -1026 44318 -1022 44724
rect -1002 44318 -998 44724
rect -978 44318 -974 44724
rect -954 44318 -950 44724
rect -930 44318 -926 44724
rect -906 44318 -902 44724
rect -882 44318 -878 44724
rect -858 44723 -854 44724
rect -858 44675 -851 44723
rect -858 44318 -854 44675
rect -834 44318 -830 44724
rect -810 44318 -806 44724
rect -786 44318 -782 44724
rect -762 44318 -758 44724
rect -738 44318 -734 44724
rect -714 44318 -710 44724
rect -690 44318 -686 44724
rect -666 44318 -662 44724
rect -659 44723 -645 44724
rect -642 44723 -635 44747
rect -642 44318 -638 44723
rect -618 44318 -614 44796
rect -594 44318 -590 44796
rect -570 44318 -566 44796
rect -546 44318 -542 44796
rect -522 44318 -518 44796
rect -498 44318 -494 44796
rect -474 44318 -470 44796
rect -461 44717 -456 44727
rect -450 44717 -446 44796
rect -451 44703 -446 44717
rect -450 44559 -446 44703
rect -426 44651 -422 44796
rect -426 44627 -419 44651
rect -461 44558 -427 44559
rect -426 44558 -422 44627
rect -402 44558 -398 44796
rect -378 44558 -374 44796
rect -365 44597 -360 44607
rect -354 44597 -350 44796
rect -355 44583 -350 44597
rect -354 44558 -350 44583
rect -330 44558 -326 44796
rect -323 44795 -309 44796
rect -317 44789 -312 44795
rect -307 44775 -302 44789
rect -306 44558 -302 44775
rect -293 44645 -288 44655
rect -283 44631 -278 44645
rect -282 44558 -278 44631
rect -269 44558 -261 44559
rect -461 44556 -261 44558
rect -461 44549 -456 44556
rect -450 44549 -446 44556
rect -451 44535 -446 44549
rect -461 44525 -456 44535
rect -451 44511 -446 44525
rect -450 44318 -446 44511
rect -426 44483 -422 44556
rect -426 44435 -419 44483
rect -426 44318 -422 44435
rect -402 44318 -398 44556
rect -389 44357 -384 44367
rect -378 44357 -374 44556
rect -379 44343 -374 44357
rect -389 44333 -384 44343
rect -378 44333 -374 44343
rect -379 44319 -374 44333
rect -389 44318 -355 44319
rect -2393 44316 -355 44318
rect -2371 44270 -2366 44316
rect -2348 44270 -2343 44316
rect -2325 44308 -2317 44316
rect -2018 44315 -2004 44316
rect -2000 44315 -1992 44316
rect -2072 44314 -1928 44315
rect -2072 44308 -2053 44314
rect -2325 44292 -2320 44308
rect -2317 44306 -2309 44308
rect -2309 44294 -2301 44306
rect -2092 44299 -2062 44304
rect -2317 44292 -2309 44294
rect -2325 44280 -2317 44292
rect -2098 44286 -2096 44297
rect -2092 44286 -2084 44299
rect -2000 44298 -1992 44314
rect -1972 44308 -1928 44314
rect -1924 44308 -1918 44316
rect -1671 44308 -1663 44316
rect -1663 44306 -1655 44308
rect -2083 44288 -2062 44297
rect -2027 44296 -1992 44298
rect -2018 44288 -2002 44296
rect -2000 44288 -1992 44296
rect -2100 44281 -2096 44286
rect -2083 44281 -2053 44286
rect -2003 44284 -1990 44288
rect -1972 44286 -1964 44295
rect -1928 44294 -1924 44297
rect -1655 44294 -1647 44306
rect -1663 44292 -1655 44294
rect -2325 44270 -2320 44280
rect -2317 44278 -2309 44280
rect -2309 44270 -2301 44278
rect -2004 44274 -2003 44284
rect -2062 44270 -2012 44272
rect -2000 44270 -1992 44284
rect -1972 44281 -1924 44286
rect -1864 44281 -1796 44287
rect -1671 44280 -1663 44292
rect -1663 44278 -1655 44280
rect -1864 44270 -1796 44271
rect -1655 44270 -1647 44278
rect -1642 44270 -1637 44316
rect -1619 44270 -1614 44316
rect -1530 44270 -1526 44316
rect -1506 44270 -1502 44316
rect -1482 44270 -1478 44316
rect -1458 44270 -1454 44316
rect -1434 44270 -1430 44316
rect -1410 44270 -1406 44316
rect -1386 44270 -1382 44316
rect -1362 44270 -1358 44316
rect -1338 44270 -1334 44316
rect -1314 44270 -1310 44316
rect -1290 44270 -1286 44316
rect -1266 44270 -1262 44316
rect -1242 44270 -1238 44316
rect -1218 44270 -1214 44316
rect -1194 44270 -1190 44316
rect -1170 44270 -1166 44316
rect -1146 44270 -1142 44316
rect -1122 44270 -1118 44316
rect -1098 44270 -1094 44316
rect -1074 44270 -1070 44316
rect -1050 44270 -1046 44316
rect -1026 44270 -1022 44316
rect -1002 44270 -998 44316
rect -978 44270 -974 44316
rect -954 44270 -950 44316
rect -930 44270 -926 44316
rect -906 44270 -902 44316
rect -882 44270 -878 44316
rect -858 44270 -854 44316
rect -834 44270 -830 44316
rect -810 44270 -806 44316
rect -786 44270 -782 44316
rect -762 44270 -758 44316
rect -738 44270 -734 44316
rect -714 44270 -710 44316
rect -690 44270 -686 44316
rect -666 44270 -662 44316
rect -642 44270 -638 44316
rect -618 44270 -614 44316
rect -594 44270 -590 44316
rect -570 44270 -566 44316
rect -546 44270 -542 44316
rect -522 44270 -518 44316
rect -498 44270 -494 44316
rect -474 44270 -470 44316
rect -450 44270 -446 44316
rect -426 44270 -422 44316
rect -402 44270 -398 44316
rect -389 44309 -384 44316
rect -379 44295 -374 44309
rect -378 44270 -374 44295
rect -354 44291 -350 44556
rect -330 44531 -326 44556
rect -330 44507 -323 44531
rect -365 44270 -357 44271
rect -2393 44268 -357 44270
rect -2371 44222 -2366 44268
rect -2348 44222 -2343 44268
rect -2325 44264 -2320 44268
rect -2309 44266 -2301 44268
rect -2317 44264 -2309 44266
rect -2325 44252 -2317 44264
rect -2325 44222 -2320 44252
rect -2317 44250 -2309 44252
rect -2092 44238 -2062 44240
rect -2094 44234 -2062 44238
rect -2000 44222 -1992 44268
rect -1655 44266 -1647 44268
rect -1663 44264 -1655 44266
rect -1671 44252 -1663 44264
rect -1663 44250 -1655 44252
rect -1854 44238 -1806 44240
rect -1854 44234 -1680 44238
rect -1642 44222 -1637 44268
rect -1619 44222 -1614 44268
rect -1530 44222 -1526 44268
rect -1506 44222 -1502 44268
rect -1482 44222 -1478 44268
rect -1458 44222 -1454 44268
rect -1434 44222 -1430 44268
rect -1410 44222 -1406 44268
rect -1386 44222 -1382 44268
rect -1362 44222 -1358 44268
rect -1338 44222 -1334 44268
rect -1314 44222 -1310 44268
rect -1290 44222 -1286 44268
rect -1266 44222 -1262 44268
rect -1242 44222 -1238 44268
rect -1218 44222 -1214 44268
rect -1194 44222 -1190 44268
rect -1170 44222 -1166 44268
rect -1146 44222 -1142 44268
rect -1122 44222 -1118 44268
rect -1098 44222 -1094 44268
rect -1085 44237 -1080 44247
rect -1074 44237 -1070 44268
rect -1075 44223 -1070 44237
rect -1085 44222 -1051 44223
rect -2393 44220 -1051 44222
rect -2371 44198 -2366 44220
rect -2348 44198 -2343 44220
rect -2325 44198 -2320 44220
rect -2072 44218 -2036 44219
rect -2072 44212 -2054 44218
rect -2309 44204 -2301 44212
rect -2317 44198 -2309 44204
rect -2092 44203 -2062 44208
rect -2000 44199 -1992 44220
rect -1938 44219 -1906 44220
rect -1920 44218 -1906 44219
rect -1806 44212 -1680 44218
rect -1854 44203 -1806 44208
rect -1655 44204 -1647 44212
rect -1982 44199 -1966 44200
rect -2000 44198 -1966 44199
rect -1846 44198 -1806 44201
rect -1663 44198 -1655 44204
rect -1642 44198 -1637 44220
rect -1619 44198 -1614 44220
rect -1554 44206 -1547 44219
rect -2393 44196 -1557 44198
rect -2371 44174 -2366 44196
rect -2348 44174 -2343 44196
rect -2325 44174 -2320 44196
rect -2000 44194 -1966 44196
rect -2309 44176 -2301 44184
rect -2062 44183 -2054 44190
rect -2092 44176 -2084 44183
rect -2062 44176 -2026 44178
rect -2317 44174 -2309 44176
rect -2062 44174 -2012 44176
rect -2000 44174 -1992 44194
rect -1982 44193 -1966 44194
rect -1846 44192 -1806 44196
rect -1846 44185 -1798 44190
rect -1806 44183 -1798 44185
rect -1854 44181 -1846 44183
rect -1854 44176 -1806 44181
rect -1655 44176 -1647 44184
rect -1864 44174 -1796 44175
rect -1663 44174 -1655 44176
rect -1642 44174 -1637 44196
rect -1619 44174 -1614 44196
rect -1571 44195 -1557 44196
rect -1554 44195 -1547 44196
rect -1530 44174 -1526 44220
rect -1506 44174 -1502 44220
rect -1482 44174 -1478 44220
rect -1458 44174 -1454 44220
rect -1434 44174 -1430 44220
rect -1410 44174 -1406 44220
rect -1386 44174 -1382 44220
rect -1362 44174 -1358 44220
rect -1338 44174 -1334 44220
rect -1314 44174 -1310 44220
rect -1290 44174 -1286 44220
rect -1266 44174 -1262 44220
rect -1242 44174 -1238 44220
rect -1218 44174 -1214 44220
rect -1194 44174 -1190 44220
rect -1181 44189 -1176 44199
rect -1170 44189 -1166 44220
rect -1171 44175 -1166 44189
rect -1170 44174 -1166 44175
rect -1146 44174 -1142 44220
rect -1122 44174 -1118 44220
rect -1098 44174 -1094 44220
rect -1085 44213 -1080 44220
rect -1075 44199 -1070 44213
rect -1074 44174 -1070 44199
rect -1050 44174 -1046 44268
rect -1026 44174 -1022 44268
rect -1002 44174 -998 44268
rect -978 44174 -974 44268
rect -954 44174 -950 44268
rect -930 44174 -926 44268
rect -906 44174 -902 44268
rect -882 44174 -878 44268
rect -858 44174 -854 44268
rect -834 44174 -830 44268
rect -810 44174 -806 44268
rect -786 44174 -782 44268
rect -762 44174 -758 44268
rect -738 44174 -734 44268
rect -714 44174 -710 44268
rect -690 44174 -686 44268
rect -666 44174 -662 44268
rect -642 44174 -638 44268
rect -618 44174 -614 44268
rect -594 44174 -590 44268
rect -570 44174 -566 44268
rect -546 44174 -542 44268
rect -522 44174 -518 44268
rect -498 44174 -494 44268
rect -474 44174 -470 44268
rect -450 44174 -446 44268
rect -426 44174 -422 44268
rect -402 44174 -398 44268
rect -378 44174 -374 44268
rect -371 44267 -357 44268
rect -365 44261 -360 44267
rect -354 44261 -347 44291
rect -355 44247 -347 44261
rect -354 44246 -347 44247
rect -330 44246 -326 44507
rect -306 44246 -302 44556
rect -282 44246 -278 44556
rect -275 44555 -261 44556
rect -269 44549 -264 44555
rect -259 44535 -254 44549
rect -258 44246 -254 44535
rect -245 44405 -240 44415
rect -235 44391 -230 44405
rect -234 44246 -230 44391
rect -211 44319 -203 44333
rect -210 44315 -203 44319
rect -210 44246 -206 44315
rect -197 44246 -189 44247
rect -371 44244 -189 44246
rect -371 44243 -357 44244
rect -354 44219 -347 44244
rect -354 44174 -350 44219
rect -330 44195 -326 44244
rect -2393 44172 -333 44174
rect -2371 44126 -2366 44172
rect -2348 44126 -2343 44172
rect -2325 44126 -2320 44172
rect -2317 44168 -2309 44172
rect -2062 44168 -2054 44172
rect -2154 44164 -2138 44166
rect -2057 44164 -2054 44168
rect -2292 44158 -2054 44164
rect -2052 44158 -2044 44168
rect -2092 44142 -2062 44144
rect -2094 44138 -2062 44142
rect -2000 44126 -1992 44172
rect -1846 44165 -1806 44172
rect -1663 44168 -1655 44172
rect -1846 44158 -1680 44164
rect -1854 44142 -1806 44144
rect -1854 44138 -1680 44142
rect -1642 44126 -1637 44172
rect -1619 44126 -1614 44172
rect -1530 44126 -1526 44172
rect -1506 44126 -1502 44172
rect -1482 44126 -1478 44172
rect -1458 44126 -1454 44172
rect -1434 44126 -1430 44172
rect -1410 44126 -1406 44172
rect -1386 44126 -1382 44172
rect -1362 44126 -1358 44172
rect -1338 44126 -1334 44172
rect -1314 44126 -1310 44172
rect -1290 44126 -1286 44172
rect -1266 44126 -1262 44172
rect -1242 44126 -1238 44172
rect -1218 44126 -1214 44172
rect -1194 44126 -1190 44172
rect -1170 44126 -1166 44172
rect -1157 44141 -1152 44151
rect -1146 44141 -1142 44172
rect -1147 44127 -1142 44141
rect -1157 44126 -1123 44127
rect -2393 44124 -1123 44126
rect -2371 44102 -2366 44124
rect -2348 44102 -2343 44124
rect -2325 44102 -2320 44124
rect -2072 44122 -2036 44123
rect -2072 44116 -2054 44122
rect -2309 44108 -2301 44116
rect -2317 44102 -2309 44108
rect -2092 44107 -2062 44112
rect -2000 44103 -1992 44124
rect -1938 44123 -1906 44124
rect -1920 44122 -1906 44123
rect -1806 44116 -1680 44122
rect -1854 44107 -1806 44112
rect -1655 44108 -1647 44116
rect -1982 44103 -1966 44104
rect -2000 44102 -1966 44103
rect -1846 44102 -1806 44105
rect -1663 44102 -1655 44108
rect -1642 44102 -1637 44124
rect -1619 44102 -1614 44124
rect -1530 44102 -1526 44124
rect -1506 44102 -1502 44124
rect -1482 44102 -1478 44124
rect -1458 44102 -1454 44124
rect -1434 44102 -1430 44124
rect -1410 44102 -1406 44124
rect -1386 44102 -1382 44124
rect -1362 44102 -1358 44124
rect -1338 44102 -1334 44124
rect -1314 44102 -1310 44124
rect -1290 44102 -1286 44124
rect -1266 44102 -1262 44124
rect -1242 44102 -1238 44124
rect -1218 44102 -1214 44124
rect -1194 44102 -1190 44124
rect -1170 44102 -1166 44124
rect -1157 44117 -1152 44124
rect -1147 44103 -1139 44117
rect -2393 44100 -1149 44102
rect -2371 44078 -2366 44100
rect -2348 44078 -2343 44100
rect -2325 44078 -2320 44100
rect -2000 44098 -1966 44100
rect -2309 44080 -2301 44088
rect -2062 44087 -2054 44094
rect -2092 44080 -2084 44087
rect -2062 44080 -2026 44082
rect -2317 44078 -2309 44080
rect -2062 44078 -2012 44080
rect -2000 44078 -1992 44098
rect -1982 44097 -1966 44098
rect -1846 44096 -1806 44100
rect -1846 44089 -1798 44094
rect -1806 44087 -1798 44089
rect -1854 44085 -1846 44087
rect -1854 44080 -1806 44085
rect -1655 44080 -1647 44088
rect -1864 44078 -1796 44079
rect -1663 44078 -1655 44080
rect -1642 44078 -1637 44100
rect -1619 44078 -1614 44100
rect -1530 44078 -1526 44100
rect -1506 44078 -1502 44100
rect -1482 44078 -1478 44100
rect -1458 44078 -1454 44100
rect -1434 44078 -1430 44100
rect -1410 44078 -1406 44100
rect -1386 44078 -1382 44100
rect -1362 44078 -1358 44100
rect -1338 44078 -1334 44100
rect -1314 44078 -1310 44100
rect -1290 44078 -1286 44100
rect -1266 44078 -1262 44100
rect -1242 44078 -1238 44100
rect -1218 44078 -1214 44100
rect -1194 44078 -1190 44100
rect -1170 44078 -1166 44100
rect -1163 44099 -1149 44100
rect -1146 44099 -1139 44103
rect -1146 44078 -1142 44099
rect -1122 44078 -1118 44172
rect -1098 44078 -1094 44172
rect -1074 44078 -1070 44172
rect -1050 44171 -1046 44172
rect -1050 44150 -1043 44171
rect -1026 44150 -1022 44172
rect -1002 44150 -998 44172
rect -978 44150 -974 44172
rect -954 44150 -950 44172
rect -930 44150 -926 44172
rect -906 44150 -902 44172
rect -882 44150 -878 44172
rect -858 44150 -854 44172
rect -834 44150 -830 44172
rect -810 44150 -806 44172
rect -786 44150 -782 44172
rect -762 44150 -758 44172
rect -738 44150 -734 44172
rect -714 44150 -710 44172
rect -690 44150 -686 44172
rect -666 44150 -662 44172
rect -642 44150 -638 44172
rect -618 44150 -614 44172
rect -594 44150 -590 44172
rect -570 44150 -566 44172
rect -546 44150 -542 44172
rect -522 44150 -518 44172
rect -498 44150 -494 44172
rect -474 44150 -470 44172
rect -450 44150 -446 44172
rect -426 44150 -422 44172
rect -402 44150 -398 44172
rect -378 44150 -374 44172
rect -354 44150 -350 44172
rect -347 44171 -333 44172
rect -330 44171 -323 44195
rect -330 44150 -326 44171
rect -306 44150 -302 44244
rect -282 44150 -278 44244
rect -269 44165 -264 44175
rect -258 44165 -254 44244
rect -259 44151 -254 44165
rect -258 44150 -254 44151
rect -234 44150 -230 44244
rect -210 44150 -206 44244
rect -203 44243 -189 44244
rect -197 44237 -192 44243
rect -187 44223 -182 44237
rect -186 44150 -182 44223
rect -173 44150 -165 44151
rect -1067 44148 -165 44150
rect -1067 44147 -1053 44148
rect -1050 44123 -1043 44148
rect -1050 44078 -1046 44123
rect -1026 44078 -1022 44148
rect -1002 44078 -998 44148
rect -978 44078 -974 44148
rect -954 44078 -950 44148
rect -941 44093 -936 44103
rect -930 44093 -926 44148
rect -931 44079 -926 44093
rect -930 44078 -926 44079
rect -906 44078 -902 44148
rect -882 44078 -878 44148
rect -858 44078 -854 44148
rect -834 44078 -830 44148
rect -810 44078 -806 44148
rect -786 44078 -782 44148
rect -762 44078 -758 44148
rect -738 44078 -734 44148
rect -714 44078 -710 44148
rect -690 44078 -686 44148
rect -666 44078 -662 44148
rect -642 44078 -638 44148
rect -618 44078 -614 44148
rect -594 44078 -590 44148
rect -570 44078 -566 44148
rect -546 44078 -542 44148
rect -522 44078 -518 44148
rect -498 44078 -494 44148
rect -474 44078 -470 44148
rect -450 44078 -446 44148
rect -426 44078 -422 44148
rect -402 44078 -398 44148
rect -378 44078 -374 44148
rect -354 44078 -350 44148
rect -330 44078 -326 44148
rect -306 44078 -302 44148
rect -282 44078 -278 44148
rect -258 44079 -254 44148
rect -234 44099 -230 44148
rect -269 44078 -237 44079
rect -2393 44076 -237 44078
rect -2371 44030 -2366 44076
rect -2348 44030 -2343 44076
rect -2325 44030 -2320 44076
rect -2317 44072 -2309 44076
rect -2062 44072 -2054 44076
rect -2154 44068 -2138 44070
rect -2057 44068 -2054 44072
rect -2292 44062 -2054 44068
rect -2052 44062 -2044 44072
rect -2092 44046 -2062 44048
rect -2094 44042 -2062 44046
rect -2000 44030 -1992 44076
rect -1846 44069 -1806 44076
rect -1663 44072 -1655 44076
rect -1846 44062 -1680 44068
rect -1854 44046 -1806 44048
rect -1854 44042 -1680 44046
rect -1979 44030 -1945 44032
rect -1642 44030 -1637 44076
rect -1619 44030 -1614 44076
rect -1530 44030 -1526 44076
rect -1506 44030 -1502 44076
rect -1482 44030 -1478 44076
rect -1458 44030 -1454 44076
rect -1434 44030 -1430 44076
rect -1410 44030 -1406 44076
rect -1386 44030 -1382 44076
rect -1362 44030 -1358 44076
rect -1338 44030 -1334 44076
rect -1314 44030 -1310 44076
rect -1290 44030 -1286 44076
rect -1266 44030 -1262 44076
rect -1242 44030 -1238 44076
rect -1218 44030 -1214 44076
rect -1194 44030 -1190 44076
rect -1170 44030 -1166 44076
rect -1146 44030 -1142 44076
rect -1122 44075 -1118 44076
rect -2393 44028 -1125 44030
rect -2371 43982 -2366 44028
rect -2348 43982 -2343 44028
rect -2325 43982 -2320 44028
rect -2080 44027 -1906 44028
rect -2080 44026 -2036 44027
rect -2080 44020 -2054 44026
rect -2309 44012 -2301 44018
rect -2317 44002 -2309 44012
rect -2070 44011 -2040 44018
rect -2054 44003 -2040 44006
rect -2000 44001 -1992 44027
rect -1920 44026 -1906 44027
rect -1850 44020 -1846 44028
rect -1840 44020 -1792 44028
rect -1969 44008 -1966 44017
rect -1850 44013 -1802 44018
rect -1906 44011 -1802 44013
rect -1655 44012 -1647 44018
rect -1906 44010 -1850 44011
rect -1846 44003 -1802 44009
rect -1663 44002 -1655 44012
rect -1860 44001 -1798 44002
rect -2078 43994 -2070 44001
rect -2309 43984 -2301 43990
rect -2317 43982 -2309 43984
rect -2154 43982 -2145 43992
rect -2044 43991 -2040 43996
rect -2028 43994 -1945 44001
rect -1929 43994 -1794 44001
rect -2070 43984 -2040 43991
rect -2044 43982 -2028 43984
rect -2000 43982 -1992 43994
rect -1860 43993 -1798 43994
rect -1850 43984 -1802 43991
rect -1655 43984 -1647 43990
rect -1978 43982 -1942 43983
rect -1663 43982 -1655 43984
rect -1642 43982 -1637 44028
rect -1619 43982 -1614 44028
rect -1589 43982 -1555 43983
rect -2393 43980 -1555 43982
rect -2371 43862 -2366 43980
rect -2348 43862 -2343 43980
rect -2325 43942 -2320 43980
rect -2317 43974 -2309 43980
rect -2145 43976 -2138 43980
rect -2070 43976 -2054 43980
rect -2078 43967 -2054 43974
rect -2062 43942 -2032 43943
rect -2000 43942 -1992 43980
rect -1846 43976 -1802 43980
rect -1846 43966 -1792 43975
rect -1663 43974 -1655 43980
rect -1942 43944 -1937 43956
rect -1850 43953 -1822 43954
rect -1850 43949 -1802 43953
rect -2325 43934 -2317 43942
rect -2062 43940 -1961 43942
rect -2325 43914 -2320 43934
rect -2317 43926 -2309 43934
rect -2062 43927 -2040 43938
rect -2032 43933 -1961 43940
rect -1947 43934 -1942 43942
rect -1842 43940 -1794 43943
rect -2070 43922 -2022 43926
rect -2325 43902 -2317 43914
rect -2137 43905 -2121 43907
rect -2325 43886 -2320 43902
rect -2317 43898 -2309 43902
rect -2292 43900 -2085 43905
rect -2069 43900 -2032 43902
rect -2309 43886 -2301 43898
rect -2125 43894 -2121 43895
rect -2325 43874 -2317 43886
rect -2059 43878 -2045 43882
rect -2325 43862 -2320 43874
rect -2317 43870 -2309 43874
rect -2309 43862 -2301 43870
rect -2025 43866 -2022 43872
rect -2000 43866 -1992 43933
rect -1942 43932 -1937 43934
rect -1932 43924 -1927 43932
rect -1912 43929 -1896 43935
rect -1842 43927 -1802 43938
rect -1671 43934 -1663 43942
rect -1663 43926 -1655 43934
rect -1850 43922 -1680 43926
rect -1671 43902 -1663 43914
rect -1663 43898 -1655 43902
rect -1977 43891 -1929 43897
rect -1974 43882 -1944 43891
rect -1655 43886 -1647 43898
rect -1960 43881 -1944 43882
rect -1671 43874 -1663 43886
rect -1977 43869 -1929 43871
rect -1663 43870 -1655 43874
rect -2033 43864 -1992 43866
rect -2062 43862 -1992 43864
rect -1655 43862 -1647 43870
rect -1642 43862 -1637 43980
rect -1619 43862 -1614 43980
rect -1554 43894 -1547 43907
rect -1554 43883 -1547 43884
rect -1530 43862 -1526 44028
rect -1506 43862 -1502 44028
rect -1482 43862 -1478 44028
rect -1458 43862 -1454 44028
rect -1434 43863 -1430 44028
rect -1445 43862 -1411 43863
rect -2393 43860 -1411 43862
rect -2371 43742 -2366 43860
rect -2348 43742 -2343 43860
rect -2325 43858 -2320 43860
rect -2309 43858 -2301 43860
rect -2325 43846 -2317 43858
rect -2025 43856 -2022 43860
rect -2062 43846 -2032 43847
rect -2325 43826 -2320 43846
rect -2317 43842 -2309 43846
rect -2325 43818 -2317 43826
rect -2325 43798 -2320 43818
rect -2317 43810 -2309 43818
rect -2117 43809 -2095 43819
rect -2045 43816 -2037 43830
rect -2325 43782 -2317 43798
rect -2325 43766 -2320 43782
rect -2309 43770 -2301 43782
rect -2317 43766 -2309 43770
rect -2117 43768 -2095 43775
rect -2069 43774 -2041 43782
rect -2017 43780 -2015 43782
rect -2325 43754 -2317 43766
rect -2125 43759 -2095 43766
rect -2047 43764 -2011 43766
rect -2059 43762 -2011 43764
rect -2000 43762 -1992 43860
rect -1888 43853 -1874 43860
rect -1655 43858 -1647 43860
rect -1671 43846 -1663 43858
rect -1663 43842 -1655 43846
rect -1969 43809 -1929 43821
rect -1671 43818 -1663 43826
rect -1663 43810 -1655 43818
rect -1671 43782 -1663 43798
rect -1655 43770 -1647 43782
rect -1663 43766 -1655 43770
rect -2125 43757 -2117 43759
rect -2059 43758 -2045 43762
rect -2021 43759 -1992 43762
rect -1977 43759 -1929 43766
rect -2325 43742 -2320 43754
rect -2309 43742 -2301 43754
rect -2131 43749 -2129 43754
rect -2125 43751 -2095 43757
rect -2021 43752 -2009 43756
rect -2125 43749 -2117 43751
rect -2133 43742 -2129 43749
rect -2117 43742 -2087 43749
rect -2025 43746 -2021 43752
rect -2000 43746 -1992 43759
rect -1969 43751 -1929 43757
rect -1671 43754 -1663 43766
rect -2033 43742 -1992 43746
rect -1969 43742 -1921 43749
rect -1655 43742 -1647 43754
rect -1642 43742 -1637 43860
rect -1619 43742 -1614 43860
rect -1530 43742 -1526 43860
rect -1506 43742 -1502 43860
rect -1482 43742 -1478 43860
rect -1458 43742 -1454 43860
rect -1445 43853 -1440 43860
rect -1434 43853 -1430 43860
rect -1435 43839 -1430 43853
rect -1434 43742 -1430 43839
rect -1410 43787 -1406 44028
rect -1410 43763 -1403 43787
rect -1410 43742 -1406 43763
rect -1386 43742 -1382 44028
rect -1373 43829 -1368 43839
rect -1362 43829 -1358 44028
rect -1363 43815 -1358 43829
rect -1362 43743 -1358 43815
rect -1338 43763 -1334 44028
rect -1373 43742 -1341 43743
rect -2393 43740 -1341 43742
rect -2371 43646 -2366 43740
rect -2348 43646 -2343 43740
rect -2325 43738 -2320 43740
rect -2317 43738 -2309 43740
rect -2131 43738 -2129 43740
rect -2125 43738 -2095 43740
rect -2325 43726 -2317 43738
rect -2117 43733 -2095 43738
rect -2325 43706 -2320 43726
rect -2325 43698 -2317 43706
rect -2325 43646 -2320 43698
rect -2317 43690 -2309 43698
rect -2117 43689 -2095 43699
rect -2045 43696 -2037 43710
rect -2309 43650 -2301 43658
rect -2317 43646 -2309 43650
rect -2000 43646 -1992 43740
rect -1663 43738 -1655 43740
rect -1671 43726 -1663 43738
rect -1969 43689 -1929 43701
rect -1671 43698 -1663 43706
rect -1663 43690 -1655 43698
rect -1655 43650 -1647 43658
rect -1663 43646 -1655 43650
rect -1642 43646 -1637 43740
rect -1619 43646 -1614 43740
rect -1530 43646 -1526 43740
rect -1506 43646 -1502 43740
rect -1482 43646 -1478 43740
rect -1458 43646 -1454 43740
rect -1434 43646 -1430 43740
rect -1410 43646 -1406 43740
rect -1397 43709 -1392 43719
rect -1386 43709 -1382 43740
rect -1373 43733 -1368 43740
rect -1362 43733 -1358 43740
rect -1355 43739 -1341 43740
rect -1338 43739 -1331 43763
rect -1363 43719 -1358 43733
rect -1387 43695 -1382 43709
rect -1386 43646 -1382 43695
rect -1362 43646 -1358 43719
rect -1338 43667 -1334 43739
rect -2393 43644 -2026 43646
rect -2021 43644 -1341 43646
rect -2371 43550 -2366 43644
rect -2348 43550 -2343 43644
rect -2325 43582 -2320 43644
rect -2317 43642 -2309 43644
rect -2309 43622 -2301 43630
rect -2317 43614 -2309 43622
rect -2123 43617 -2116 43622
rect -2123 43615 -2092 43617
rect -2091 43616 -2087 43632
rect -2026 43624 -2021 43636
rect -2037 43620 -2021 43624
rect -2292 43613 -2087 43615
rect -2123 43611 -2116 43613
rect -2325 43574 -2317 43582
rect -2325 43554 -2320 43574
rect -2317 43566 -2309 43574
rect -2325 43550 -2317 43554
rect -2000 43550 -1992 43644
rect -1663 43642 -1655 43644
rect -1969 43616 -1932 43632
rect -1655 43622 -1647 43630
rect -1969 43613 -1680 43615
rect -1663 43614 -1655 43622
rect -1671 43574 -1663 43582
rect -1663 43566 -1655 43574
rect -1671 43550 -1663 43554
rect -1642 43550 -1637 43644
rect -1619 43550 -1614 43644
rect -1530 43550 -1526 43644
rect -1506 43550 -1502 43644
rect -1493 43565 -1488 43575
rect -1482 43565 -1478 43644
rect -1483 43551 -1478 43565
rect -1493 43550 -1459 43551
rect -2393 43548 -1459 43550
rect -2371 43502 -2366 43548
rect -2348 43502 -2343 43548
rect -2325 43540 -2317 43548
rect -2018 43547 -2004 43548
rect -2000 43547 -1992 43548
rect -2072 43546 -1928 43547
rect -2072 43540 -2053 43546
rect -2325 43524 -2320 43540
rect -2317 43538 -2309 43540
rect -2309 43526 -2301 43538
rect -2092 43531 -2062 43536
rect -2317 43524 -2309 43526
rect -2325 43512 -2317 43524
rect -2098 43518 -2096 43529
rect -2092 43518 -2084 43531
rect -2000 43530 -1992 43546
rect -1972 43540 -1928 43546
rect -1924 43540 -1918 43548
rect -1671 43540 -1663 43548
rect -1663 43538 -1655 43540
rect -2083 43520 -2062 43529
rect -2027 43528 -1992 43530
rect -2018 43520 -2002 43528
rect -2000 43520 -1992 43528
rect -2100 43513 -2096 43518
rect -2083 43513 -2053 43518
rect -2003 43516 -1990 43520
rect -1972 43518 -1964 43527
rect -1928 43526 -1924 43529
rect -1655 43526 -1647 43538
rect -1663 43524 -1655 43526
rect -2325 43502 -2320 43512
rect -2317 43510 -2309 43512
rect -2309 43502 -2301 43510
rect -2004 43506 -2003 43516
rect -2062 43502 -2012 43504
rect -2000 43502 -1992 43516
rect -1972 43513 -1924 43518
rect -1864 43513 -1796 43519
rect -1671 43512 -1663 43524
rect -1663 43510 -1655 43512
rect -1864 43502 -1796 43503
rect -1655 43502 -1647 43510
rect -1642 43502 -1637 43548
rect -1619 43502 -1614 43548
rect -1530 43502 -1526 43548
rect -1506 43502 -1502 43548
rect -1493 43541 -1488 43548
rect -1483 43527 -1478 43541
rect -1482 43502 -1478 43527
rect -1458 43502 -1454 43644
rect -1434 43502 -1430 43644
rect -1410 43502 -1406 43644
rect -1386 43502 -1382 43644
rect -1362 43643 -1358 43644
rect -1355 43643 -1341 43644
rect -1338 43643 -1331 43667
rect -1362 43619 -1355 43643
rect -1362 43502 -1358 43619
rect -1338 43502 -1334 43643
rect -1314 43502 -1310 44028
rect -1301 43661 -1296 43671
rect -1290 43661 -1286 44028
rect -1291 43647 -1286 43661
rect -1301 43637 -1296 43647
rect -1291 43623 -1286 43637
rect -1290 43502 -1286 43623
rect -1266 43595 -1262 44028
rect -1266 43574 -1259 43595
rect -1242 43574 -1238 44028
rect -1218 43574 -1214 44028
rect -1194 43574 -1190 44028
rect -1170 43574 -1166 44028
rect -1146 43574 -1142 44028
rect -1139 44027 -1125 44028
rect -1122 44027 -1115 44075
rect -1122 43815 -1118 44027
rect -1133 43814 -1099 43815
rect -1098 43814 -1094 44076
rect -1074 43814 -1070 44076
rect -1050 43814 -1046 44076
rect -1026 43814 -1022 44076
rect -1002 43814 -998 44076
rect -978 43814 -974 44076
rect -954 43814 -950 44076
rect -930 43814 -926 44076
rect -906 44027 -902 44076
rect -906 44003 -899 44027
rect -906 43814 -902 44003
rect -882 43814 -878 44076
rect -858 43814 -854 44076
rect -834 43814 -830 44076
rect -810 43814 -806 44076
rect -786 43814 -782 44076
rect -762 43814 -758 44076
rect -738 43814 -734 44076
rect -714 43814 -710 44076
rect -690 43814 -686 44076
rect -666 43814 -662 44076
rect -642 43814 -638 44076
rect -618 43814 -614 44076
rect -594 43814 -590 44076
rect -581 43949 -576 43959
rect -570 43949 -566 44076
rect -571 43935 -566 43949
rect -570 43814 -566 43935
rect -546 43883 -542 44076
rect -546 43859 -539 43883
rect -546 43814 -542 43859
rect -522 43814 -518 44076
rect -498 43814 -494 44076
rect -474 43814 -470 44076
rect -450 43814 -446 44076
rect -426 43814 -422 44076
rect -402 44055 -398 44076
rect -413 44054 -379 44055
rect -378 44054 -374 44076
rect -354 44054 -350 44076
rect -330 44054 -326 44076
rect -306 44054 -302 44076
rect -282 44054 -278 44076
rect -269 44069 -264 44076
rect -258 44069 -254 44076
rect -251 44075 -237 44076
rect -234 44075 -227 44099
rect -259 44055 -254 44069
rect -258 44054 -254 44055
rect -234 44054 -230 44075
rect -210 44054 -206 44148
rect -186 44054 -182 44148
rect -179 44147 -165 44148
rect -173 44141 -168 44147
rect -163 44127 -158 44141
rect -162 44054 -158 44127
rect -149 44054 -141 44055
rect -413 44052 -141 44054
rect -413 44045 -408 44052
rect -402 44045 -398 44052
rect -403 44031 -398 44045
rect -413 44021 -408 44031
rect -403 44007 -398 44021
rect -402 43814 -398 44007
rect -378 43979 -374 44052
rect -378 43931 -371 43979
rect -378 43814 -374 43931
rect -354 43814 -350 44052
rect -330 43814 -326 44052
rect -306 43814 -302 44052
rect -282 43814 -278 44052
rect -269 43925 -264 43935
rect -258 43925 -254 44052
rect -259 43911 -254 43925
rect -234 44003 -230 44052
rect -234 43979 -227 44003
rect -269 43901 -264 43911
rect -259 43887 -254 43901
rect -258 43814 -254 43887
rect -234 43859 -230 43979
rect -1133 43812 -237 43814
rect -1133 43805 -1128 43812
rect -1122 43805 -1118 43812
rect -1123 43791 -1118 43805
rect -1133 43781 -1128 43791
rect -1123 43767 -1118 43781
rect -1122 43574 -1118 43767
rect -1098 43739 -1094 43812
rect -1098 43691 -1091 43739
rect -1098 43574 -1094 43691
rect -1074 43574 -1070 43812
rect -1050 43574 -1046 43812
rect -1026 43574 -1022 43812
rect -1002 43574 -998 43812
rect -978 43574 -974 43812
rect -954 43574 -950 43812
rect -930 43574 -926 43812
rect -906 43574 -902 43812
rect -882 43574 -878 43812
rect -858 43574 -854 43812
rect -834 43574 -830 43812
rect -810 43574 -806 43812
rect -786 43574 -782 43812
rect -762 43574 -758 43812
rect -738 43574 -734 43812
rect -714 43574 -710 43812
rect -690 43574 -686 43812
rect -666 43574 -662 43812
rect -642 43574 -638 43812
rect -618 43574 -614 43812
rect -594 43574 -590 43812
rect -570 43574 -566 43812
rect -546 43574 -542 43812
rect -522 43574 -518 43812
rect -498 43574 -494 43812
rect -474 43574 -470 43812
rect -450 43574 -446 43812
rect -426 43574 -422 43812
rect -402 43574 -398 43812
rect -378 43574 -374 43812
rect -354 43574 -350 43812
rect -330 43574 -326 43812
rect -306 43574 -302 43812
rect -282 43574 -278 43812
rect -258 43574 -254 43812
rect -251 43811 -237 43812
rect -234 43811 -227 43859
rect -234 43574 -230 43811
rect -210 43574 -206 44052
rect -186 43574 -182 44052
rect -173 43589 -168 43599
rect -162 43589 -158 44052
rect -155 44051 -141 44052
rect -149 44045 -144 44051
rect -139 44031 -134 44045
rect -163 43575 -158 43589
rect -162 43574 -158 43575
rect -138 43574 -134 44031
rect -125 43925 -120 43935
rect -115 43911 -110 43925
rect -114 43574 -110 43911
rect -101 43805 -96 43815
rect -91 43791 -86 43805
rect -90 43574 -86 43791
rect -77 43661 -72 43671
rect -67 43647 -62 43661
rect -66 43574 -62 43647
rect -53 43574 -45 43575
rect -1283 43572 -45 43574
rect -1283 43571 -1269 43572
rect -1266 43547 -1259 43572
rect -1266 43502 -1262 43547
rect -1242 43502 -1238 43572
rect -1218 43502 -1214 43572
rect -1194 43502 -1190 43572
rect -1170 43502 -1166 43572
rect -1146 43502 -1142 43572
rect -1122 43502 -1118 43572
rect -1098 43502 -1094 43572
rect -1074 43502 -1070 43572
rect -1050 43502 -1046 43572
rect -1026 43502 -1022 43572
rect -1013 43541 -1008 43551
rect -1002 43541 -998 43572
rect -1003 43527 -998 43541
rect -1013 43517 -1008 43527
rect -1003 43503 -998 43517
rect -1002 43502 -998 43503
rect -978 43502 -974 43572
rect -954 43502 -950 43572
rect -930 43502 -926 43572
rect -906 43502 -902 43572
rect -882 43502 -878 43572
rect -858 43502 -854 43572
rect -834 43502 -830 43572
rect -810 43502 -806 43572
rect -786 43502 -782 43572
rect -762 43502 -758 43572
rect -738 43502 -734 43572
rect -714 43502 -710 43572
rect -690 43502 -686 43572
rect -666 43502 -662 43572
rect -642 43502 -638 43572
rect -618 43502 -614 43572
rect -594 43502 -590 43572
rect -570 43502 -566 43572
rect -546 43502 -542 43572
rect -522 43502 -518 43572
rect -498 43502 -494 43572
rect -474 43502 -470 43572
rect -450 43502 -446 43572
rect -426 43502 -422 43572
rect -402 43502 -398 43572
rect -378 43502 -374 43572
rect -354 43502 -350 43572
rect -330 43502 -326 43572
rect -306 43502 -302 43572
rect -282 43502 -278 43572
rect -258 43502 -254 43572
rect -234 43502 -230 43572
rect -210 43502 -206 43572
rect -186 43502 -182 43572
rect -173 43517 -168 43527
rect -162 43517 -158 43572
rect -138 43523 -134 43572
rect -163 43503 -158 43517
rect -149 43513 -141 43517
rect -155 43503 -149 43513
rect -173 43502 -141 43503
rect -2393 43500 -141 43502
rect -2371 43454 -2366 43500
rect -2348 43454 -2343 43500
rect -2325 43496 -2320 43500
rect -2309 43498 -2301 43500
rect -2317 43496 -2309 43498
rect -2325 43484 -2317 43496
rect -2325 43454 -2320 43484
rect -2317 43482 -2309 43484
rect -2092 43470 -2062 43472
rect -2094 43466 -2062 43470
rect -2000 43454 -1992 43500
rect -1655 43498 -1647 43500
rect -1663 43496 -1655 43498
rect -1671 43484 -1663 43496
rect -1663 43482 -1655 43484
rect -1854 43470 -1806 43472
rect -1854 43466 -1680 43470
rect -1642 43454 -1637 43500
rect -1619 43454 -1614 43500
rect -1530 43454 -1526 43500
rect -1506 43454 -1502 43500
rect -1482 43454 -1478 43500
rect -1458 43499 -1454 43500
rect -2393 43452 -1461 43454
rect -2371 43430 -2366 43452
rect -2348 43430 -2343 43452
rect -2325 43430 -2320 43452
rect -2072 43450 -2036 43451
rect -2072 43444 -2054 43450
rect -2309 43436 -2301 43444
rect -2317 43430 -2309 43436
rect -2092 43435 -2062 43440
rect -2000 43431 -1992 43452
rect -1938 43451 -1906 43452
rect -1920 43450 -1906 43451
rect -1806 43444 -1680 43450
rect -1854 43435 -1806 43440
rect -1655 43436 -1647 43444
rect -1982 43431 -1966 43432
rect -2000 43430 -1966 43431
rect -1846 43430 -1806 43433
rect -1663 43430 -1655 43436
rect -1642 43430 -1637 43452
rect -1619 43430 -1614 43452
rect -1530 43430 -1526 43452
rect -1506 43430 -1502 43452
rect -1482 43430 -1478 43452
rect -1475 43451 -1461 43452
rect -1458 43451 -1451 43499
rect -1458 43430 -1454 43451
rect -1434 43430 -1430 43500
rect -1410 43430 -1406 43500
rect -1386 43430 -1382 43500
rect -1362 43430 -1358 43500
rect -1338 43430 -1334 43500
rect -1314 43430 -1310 43500
rect -1290 43430 -1286 43500
rect -1266 43430 -1262 43500
rect -1242 43430 -1238 43500
rect -1218 43430 -1214 43500
rect -1194 43430 -1190 43500
rect -1170 43430 -1166 43500
rect -1146 43430 -1142 43500
rect -1122 43430 -1118 43500
rect -1098 43430 -1094 43500
rect -1074 43430 -1070 43500
rect -1050 43430 -1046 43500
rect -1026 43430 -1022 43500
rect -1002 43430 -998 43500
rect -978 43475 -974 43500
rect -978 43454 -971 43475
rect -954 43454 -950 43500
rect -930 43454 -926 43500
rect -906 43454 -902 43500
rect -882 43454 -878 43500
rect -858 43454 -854 43500
rect -834 43454 -830 43500
rect -810 43454 -806 43500
rect -786 43454 -782 43500
rect -762 43454 -758 43500
rect -738 43454 -734 43500
rect -714 43454 -710 43500
rect -690 43454 -686 43500
rect -666 43454 -662 43500
rect -642 43454 -638 43500
rect -618 43454 -614 43500
rect -594 43479 -590 43500
rect -605 43478 -571 43479
rect -570 43478 -566 43500
rect -546 43478 -542 43500
rect -522 43478 -518 43500
rect -498 43478 -494 43500
rect -474 43478 -470 43500
rect -450 43478 -446 43500
rect -426 43478 -422 43500
rect -402 43478 -398 43500
rect -378 43478 -374 43500
rect -354 43478 -350 43500
rect -330 43478 -326 43500
rect -306 43478 -302 43500
rect -282 43478 -278 43500
rect -258 43478 -254 43500
rect -234 43478 -230 43500
rect -210 43478 -206 43500
rect -186 43478 -182 43500
rect -173 43493 -168 43500
rect -155 43499 -141 43500
rect -138 43499 -131 43523
rect -163 43479 -158 43493
rect -162 43478 -158 43479
rect -138 43478 -134 43499
rect -114 43478 -110 43572
rect -90 43478 -86 43572
rect -66 43478 -62 43572
rect -59 43571 -45 43572
rect -53 43565 -48 43571
rect -43 43551 -38 43565
rect -42 43478 -38 43551
rect -605 43476 -21 43478
rect -605 43469 -600 43476
rect -594 43469 -590 43476
rect -595 43455 -590 43469
rect -605 43454 -571 43455
rect -995 43452 -571 43454
rect -995 43451 -981 43452
rect -2393 43428 -981 43430
rect -2371 43406 -2366 43428
rect -2348 43406 -2343 43428
rect -2325 43406 -2320 43428
rect -2000 43426 -1966 43428
rect -2309 43408 -2301 43416
rect -2062 43415 -2054 43422
rect -2092 43408 -2084 43415
rect -2062 43408 -2026 43410
rect -2317 43406 -2309 43408
rect -2062 43406 -2012 43408
rect -2000 43406 -1992 43426
rect -1982 43425 -1966 43426
rect -1846 43424 -1806 43428
rect -1846 43417 -1798 43422
rect -1806 43415 -1798 43417
rect -1854 43413 -1846 43415
rect -1854 43408 -1806 43413
rect -1655 43408 -1647 43416
rect -1864 43406 -1796 43407
rect -1663 43406 -1655 43408
rect -1642 43406 -1637 43428
rect -1619 43406 -1614 43428
rect -1530 43406 -1526 43428
rect -1506 43406 -1502 43428
rect -1482 43406 -1478 43428
rect -1458 43406 -1454 43428
rect -1434 43406 -1430 43428
rect -1410 43406 -1406 43428
rect -1386 43406 -1382 43428
rect -1362 43406 -1358 43428
rect -1338 43406 -1334 43428
rect -1314 43406 -1310 43428
rect -1290 43406 -1286 43428
rect -1266 43406 -1262 43428
rect -1242 43406 -1238 43428
rect -1218 43406 -1214 43428
rect -1194 43406 -1190 43428
rect -1170 43406 -1166 43428
rect -1146 43406 -1142 43428
rect -1122 43406 -1118 43428
rect -1098 43406 -1094 43428
rect -1074 43406 -1070 43428
rect -1050 43406 -1046 43428
rect -1026 43406 -1022 43428
rect -1002 43406 -998 43428
rect -995 43427 -981 43428
rect -978 43427 -971 43452
rect -978 43406 -974 43427
rect -954 43406 -950 43452
rect -930 43406 -926 43452
rect -917 43421 -912 43431
rect -906 43421 -902 43452
rect -907 43407 -902 43421
rect -906 43406 -902 43407
rect -882 43406 -878 43452
rect -858 43406 -854 43452
rect -834 43406 -830 43452
rect -810 43406 -806 43452
rect -786 43406 -782 43452
rect -762 43406 -758 43452
rect -738 43406 -734 43452
rect -714 43406 -710 43452
rect -690 43406 -686 43452
rect -666 43406 -662 43452
rect -642 43406 -638 43452
rect -618 43406 -614 43452
rect -605 43445 -600 43452
rect -595 43431 -590 43445
rect -594 43406 -590 43431
rect -570 43406 -566 43476
rect -546 43406 -542 43476
rect -522 43406 -518 43476
rect -498 43406 -494 43476
rect -474 43406 -470 43476
rect -450 43406 -446 43476
rect -426 43407 -422 43476
rect -437 43406 -403 43407
rect -2393 43404 -403 43406
rect -2371 43358 -2366 43404
rect -2348 43358 -2343 43404
rect -2325 43358 -2320 43404
rect -2317 43400 -2309 43404
rect -2062 43400 -2054 43404
rect -2154 43396 -2138 43398
rect -2057 43396 -2054 43400
rect -2292 43390 -2054 43396
rect -2052 43390 -2044 43400
rect -2092 43374 -2062 43376
rect -2094 43370 -2062 43374
rect -2000 43358 -1992 43404
rect -1846 43397 -1806 43404
rect -1663 43400 -1655 43404
rect -1846 43390 -1680 43396
rect -1854 43374 -1806 43376
rect -1854 43370 -1680 43374
rect -1642 43358 -1637 43404
rect -1619 43358 -1614 43404
rect -1530 43358 -1526 43404
rect -1506 43358 -1502 43404
rect -1482 43358 -1478 43404
rect -1458 43358 -1454 43404
rect -1434 43358 -1430 43404
rect -1410 43358 -1406 43404
rect -1386 43358 -1382 43404
rect -1362 43358 -1358 43404
rect -1338 43358 -1334 43404
rect -1325 43373 -1320 43383
rect -1314 43373 -1310 43404
rect -1315 43359 -1310 43373
rect -1325 43358 -1291 43359
rect -2393 43356 -1291 43358
rect -2371 43334 -2366 43356
rect -2348 43334 -2343 43356
rect -2325 43334 -2320 43356
rect -2072 43354 -2036 43355
rect -2072 43348 -2054 43354
rect -2309 43340 -2301 43348
rect -2317 43334 -2309 43340
rect -2092 43339 -2062 43344
rect -2000 43335 -1992 43356
rect -1938 43355 -1906 43356
rect -1920 43354 -1906 43355
rect -1806 43348 -1680 43354
rect -1854 43339 -1806 43344
rect -1655 43340 -1647 43348
rect -1982 43335 -1966 43336
rect -2000 43334 -1966 43335
rect -1846 43334 -1806 43337
rect -1663 43334 -1655 43340
rect -1642 43334 -1637 43356
rect -1619 43334 -1614 43356
rect -1530 43334 -1526 43356
rect -1506 43334 -1502 43356
rect -1482 43334 -1478 43356
rect -1458 43335 -1454 43356
rect -1469 43334 -1435 43335
rect -1434 43334 -1430 43356
rect -1410 43334 -1406 43356
rect -1386 43334 -1382 43356
rect -1362 43334 -1358 43356
rect -1338 43334 -1334 43356
rect -1325 43349 -1320 43356
rect -1315 43335 -1310 43349
rect -1314 43334 -1310 43335
rect -1290 43334 -1286 43404
rect -1266 43334 -1262 43404
rect -1242 43334 -1238 43404
rect -1218 43334 -1214 43404
rect -1194 43334 -1190 43404
rect -1170 43334 -1166 43404
rect -1146 43334 -1142 43404
rect -1122 43334 -1118 43404
rect -1098 43359 -1094 43404
rect -1109 43358 -1075 43359
rect -1074 43358 -1070 43404
rect -1050 43358 -1046 43404
rect -1026 43358 -1022 43404
rect -1002 43358 -998 43404
rect -978 43358 -974 43404
rect -954 43358 -950 43404
rect -930 43358 -926 43404
rect -906 43358 -902 43404
rect -882 43358 -878 43404
rect -858 43358 -854 43404
rect -834 43358 -830 43404
rect -810 43358 -806 43404
rect -786 43358 -782 43404
rect -762 43358 -758 43404
rect -738 43358 -734 43404
rect -714 43358 -710 43404
rect -690 43358 -686 43404
rect -666 43358 -662 43404
rect -642 43358 -638 43404
rect -618 43358 -614 43404
rect -594 43358 -590 43404
rect -570 43403 -566 43404
rect -570 43382 -563 43403
rect -546 43382 -542 43404
rect -522 43382 -518 43404
rect -498 43382 -494 43404
rect -474 43382 -470 43404
rect -450 43382 -446 43404
rect -437 43397 -432 43404
rect -426 43397 -422 43404
rect -427 43383 -422 43397
rect -426 43382 -422 43383
rect -402 43382 -398 43476
rect -378 43382 -374 43476
rect -354 43382 -350 43476
rect -330 43382 -326 43476
rect -306 43382 -302 43476
rect -282 43382 -278 43476
rect -258 43382 -254 43476
rect -234 43382 -230 43476
rect -210 43382 -206 43476
rect -186 43382 -182 43476
rect -162 43382 -158 43476
rect -138 43451 -134 43476
rect -138 43403 -131 43451
rect -138 43382 -134 43403
rect -114 43382 -110 43476
rect -90 43382 -86 43476
rect -66 43382 -62 43476
rect -42 43382 -38 43476
rect -35 43475 -21 43476
rect -18 43475 -11 43499
rect -18 43382 -14 43475
rect 6 43451 13 43475
rect 6 43382 10 43451
rect 30 43427 37 43451
rect 30 43382 34 43427
rect 43 43382 51 43383
rect -587 43380 51 43382
rect -587 43379 -573 43380
rect -1109 43356 -573 43358
rect -1109 43349 -1104 43356
rect -1098 43349 -1094 43356
rect -1099 43335 -1094 43349
rect -1109 43334 -1075 43335
rect -2393 43332 -1075 43334
rect -2371 43310 -2366 43332
rect -2348 43310 -2343 43332
rect -2325 43310 -2320 43332
rect -2000 43330 -1966 43332
rect -2309 43312 -2301 43320
rect -2062 43319 -2054 43326
rect -2092 43312 -2084 43319
rect -2062 43312 -2026 43314
rect -2317 43310 -2309 43312
rect -2062 43310 -2012 43312
rect -2000 43310 -1992 43330
rect -1982 43329 -1966 43330
rect -1846 43328 -1806 43332
rect -1846 43321 -1798 43326
rect -1806 43319 -1798 43321
rect -1854 43317 -1846 43319
rect -1854 43312 -1806 43317
rect -1655 43312 -1647 43320
rect -1864 43310 -1796 43311
rect -1663 43310 -1655 43312
rect -1642 43310 -1637 43332
rect -1619 43310 -1614 43332
rect -1530 43310 -1526 43332
rect -1506 43310 -1502 43332
rect -1482 43310 -1478 43332
rect -1469 43325 -1464 43332
rect -1458 43325 -1454 43332
rect -1459 43311 -1454 43325
rect -1469 43310 -1435 43311
rect -2393 43308 -1435 43310
rect -2371 43238 -2366 43308
rect -2348 43238 -2343 43308
rect -2325 43238 -2320 43308
rect -2317 43304 -2309 43308
rect -2062 43304 -2054 43308
rect -2154 43300 -2138 43302
rect -2057 43300 -2054 43304
rect -2292 43294 -2054 43300
rect -2052 43294 -2044 43304
rect -2092 43278 -2062 43280
rect -2094 43274 -2062 43278
rect -2309 43244 -2301 43250
rect -2317 43238 -2309 43244
rect -2000 43238 -1992 43308
rect -1846 43301 -1806 43308
rect -1663 43304 -1655 43308
rect -1846 43294 -1680 43300
rect -1854 43278 -1806 43280
rect -1854 43274 -1680 43278
rect -1655 43244 -1647 43250
rect -1663 43238 -1655 43244
rect -1642 43238 -1637 43308
rect -1619 43238 -1614 43308
rect -1530 43238 -1526 43308
rect -1506 43238 -1502 43308
rect -1482 43238 -1478 43308
rect -1469 43301 -1464 43308
rect -1459 43287 -1454 43301
rect -1458 43238 -1454 43287
rect -1434 43259 -1430 43332
rect -1410 43263 -1406 43332
rect -1421 43262 -1387 43263
rect -1386 43262 -1382 43332
rect -1362 43262 -1358 43332
rect -1338 43262 -1334 43332
rect -1314 43262 -1310 43332
rect -1290 43307 -1286 43332
rect -1421 43260 -1293 43262
rect -1434 43238 -1427 43259
rect -1421 43253 -1416 43260
rect -1410 43253 -1406 43260
rect -1411 43239 -1406 43253
rect -1421 43238 -1387 43239
rect -2393 43236 -1387 43238
rect -2371 43142 -2366 43236
rect -2348 43142 -2343 43236
rect -2325 43174 -2320 43236
rect -2317 43234 -2309 43236
rect -2000 43235 -1966 43236
rect -2000 43234 -1982 43235
rect -1663 43234 -1655 43236
rect -2028 43226 -2018 43228
rect -2309 43216 -2301 43222
rect -2091 43216 -2061 43223
rect -2317 43206 -2309 43216
rect -2044 43214 -2028 43216
rect -2026 43214 -2014 43226
rect -2084 43208 -2061 43214
rect -2044 43212 -2014 43214
rect -2292 43198 -2054 43207
rect -2325 43166 -2317 43174
rect -2325 43146 -2320 43166
rect -2317 43158 -2309 43166
rect -2325 43142 -2317 43146
rect -2000 43142 -1992 43234
rect -1982 43233 -1966 43234
rect -1980 43216 -1932 43223
rect -1655 43216 -1647 43222
rect -1846 43198 -1680 43207
rect -1663 43206 -1655 43216
rect -1671 43166 -1663 43174
rect -1663 43158 -1655 43166
rect -1671 43142 -1663 43146
rect -1642 43142 -1637 43236
rect -1619 43142 -1614 43236
rect -1530 43142 -1526 43236
rect -1506 43142 -1502 43236
rect -1482 43142 -1478 43236
rect -1458 43142 -1454 43236
rect -1451 43235 -1437 43236
rect -1434 43211 -1427 43236
rect -1421 43229 -1416 43236
rect -1411 43215 -1406 43229
rect -1434 43142 -1430 43211
rect -1410 43142 -1406 43215
rect -1386 43187 -1382 43260
rect -1386 43167 -1379 43187
rect -1397 43166 -1363 43167
rect -1362 43166 -1358 43260
rect -1338 43166 -1334 43260
rect -1314 43166 -1310 43260
rect -1307 43259 -1293 43260
rect -1290 43259 -1283 43307
rect -1290 43166 -1286 43259
rect -1266 43166 -1262 43332
rect -1242 43166 -1238 43332
rect -1229 43181 -1224 43191
rect -1218 43181 -1214 43332
rect -1219 43167 -1214 43181
rect -1218 43166 -1214 43167
rect -1194 43166 -1190 43332
rect -1170 43166 -1166 43332
rect -1146 43166 -1142 43332
rect -1122 43166 -1118 43332
rect -1109 43325 -1104 43332
rect -1099 43311 -1094 43325
rect -1098 43166 -1094 43311
rect -1074 43283 -1070 43356
rect -1074 43262 -1067 43283
rect -1050 43262 -1046 43356
rect -1026 43262 -1022 43356
rect -1002 43262 -998 43356
rect -978 43262 -974 43356
rect -954 43262 -950 43356
rect -930 43262 -926 43356
rect -906 43262 -902 43356
rect -882 43355 -878 43356
rect -882 43331 -875 43355
rect -882 43262 -878 43331
rect -858 43262 -854 43356
rect -834 43262 -830 43356
rect -810 43262 -806 43356
rect -786 43262 -782 43356
rect -762 43262 -758 43356
rect -738 43262 -734 43356
rect -714 43262 -710 43356
rect -690 43262 -686 43356
rect -666 43262 -662 43356
rect -642 43262 -638 43356
rect -618 43262 -614 43356
rect -594 43262 -590 43356
rect -587 43355 -573 43356
rect -570 43355 -563 43380
rect -570 43262 -566 43355
rect -546 43262 -542 43380
rect -522 43262 -518 43380
rect -498 43262 -494 43380
rect -474 43262 -470 43380
rect -450 43262 -446 43380
rect -426 43262 -422 43380
rect -402 43331 -398 43380
rect -402 43307 -395 43331
rect -402 43262 -398 43307
rect -378 43262 -374 43380
rect -354 43262 -350 43380
rect -330 43262 -326 43380
rect -306 43262 -302 43380
rect -282 43262 -278 43380
rect -258 43262 -254 43380
rect -234 43262 -230 43380
rect -210 43262 -206 43380
rect -186 43262 -182 43380
rect -162 43262 -158 43380
rect -138 43262 -134 43380
rect -114 43262 -110 43380
rect -90 43262 -86 43380
rect -66 43262 -62 43380
rect -42 43262 -38 43380
rect -18 43262 -14 43380
rect 6 43262 10 43380
rect 30 43262 34 43380
rect 37 43379 51 43380
rect 43 43373 48 43379
rect 53 43359 58 43373
rect 54 43262 58 43359
rect 78 43283 85 43307
rect 78 43262 82 43283
rect 91 43262 99 43263
rect -1091 43260 99 43262
rect -1091 43259 -1077 43260
rect -1074 43235 -1067 43260
rect -1074 43166 -1070 43235
rect -1050 43166 -1046 43260
rect -1026 43166 -1022 43260
rect -1002 43166 -998 43260
rect -978 43166 -974 43260
rect -954 43166 -950 43260
rect -930 43166 -926 43260
rect -906 43166 -902 43260
rect -882 43166 -878 43260
rect -858 43166 -854 43260
rect -834 43166 -830 43260
rect -810 43166 -806 43260
rect -786 43166 -782 43260
rect -762 43166 -758 43260
rect -738 43166 -734 43260
rect -714 43166 -710 43260
rect -690 43166 -686 43260
rect -666 43166 -662 43260
rect -642 43166 -638 43260
rect -618 43166 -614 43260
rect -594 43166 -590 43260
rect -570 43166 -566 43260
rect -546 43166 -542 43260
rect -522 43166 -518 43260
rect -498 43166 -494 43260
rect -474 43166 -470 43260
rect -450 43166 -446 43260
rect -426 43166 -422 43260
rect -402 43166 -398 43260
rect -378 43166 -374 43260
rect -354 43166 -350 43260
rect -330 43166 -326 43260
rect -306 43166 -302 43260
rect -282 43166 -278 43260
rect -258 43166 -254 43260
rect -234 43166 -230 43260
rect -210 43166 -206 43260
rect -186 43166 -182 43260
rect -162 43166 -158 43260
rect -138 43166 -134 43260
rect -114 43166 -110 43260
rect -90 43166 -86 43260
rect -66 43166 -62 43260
rect -42 43166 -38 43260
rect -18 43166 -14 43260
rect 6 43166 10 43260
rect 30 43166 34 43260
rect 54 43166 58 43260
rect 78 43166 82 43260
rect 85 43259 99 43260
rect 91 43253 96 43259
rect 101 43239 106 43253
rect 102 43166 106 43239
rect 115 43166 123 43167
rect -1397 43164 123 43166
rect -1397 43163 -1389 43164
rect -1386 43157 -1379 43164
rect -1387 43143 -1379 43157
rect -1397 43142 -1389 43143
rect -2393 43140 -1389 43142
rect -2371 43094 -2366 43140
rect -2348 43094 -2343 43140
rect -2325 43132 -2317 43140
rect -2018 43139 -2004 43140
rect -2000 43139 -1992 43140
rect -2072 43138 -1928 43139
rect -2072 43132 -2053 43138
rect -2325 43116 -2320 43132
rect -2317 43130 -2309 43132
rect -2309 43118 -2301 43130
rect -2092 43123 -2062 43128
rect -2317 43116 -2309 43118
rect -2325 43104 -2317 43116
rect -2098 43110 -2096 43121
rect -2092 43110 -2084 43123
rect -2000 43122 -1992 43138
rect -1972 43132 -1928 43138
rect -1924 43132 -1918 43140
rect -1671 43132 -1663 43140
rect -1663 43130 -1655 43132
rect -2083 43112 -2062 43121
rect -2027 43120 -1992 43122
rect -2018 43112 -2002 43120
rect -2000 43112 -1992 43120
rect -2100 43105 -2096 43110
rect -2083 43105 -2053 43110
rect -2003 43108 -1990 43112
rect -1972 43110 -1964 43119
rect -1928 43118 -1924 43121
rect -1655 43118 -1647 43130
rect -1663 43116 -1655 43118
rect -2325 43094 -2320 43104
rect -2317 43102 -2309 43104
rect -2309 43094 -2301 43102
rect -2004 43098 -2003 43108
rect -2062 43094 -2012 43096
rect -2000 43094 -1992 43108
rect -1972 43105 -1924 43110
rect -1864 43105 -1796 43111
rect -1671 43104 -1663 43116
rect -1663 43102 -1655 43104
rect -1864 43094 -1796 43095
rect -1655 43094 -1647 43102
rect -1642 43094 -1637 43140
rect -1619 43094 -1614 43140
rect -1530 43094 -1526 43140
rect -1506 43094 -1502 43140
rect -1482 43094 -1478 43140
rect -1458 43094 -1454 43140
rect -1434 43094 -1430 43140
rect -1410 43094 -1406 43140
rect -1403 43139 -1389 43140
rect -1397 43133 -1392 43139
rect -1387 43119 -1382 43133
rect -1386 43094 -1382 43119
rect -1362 43094 -1358 43164
rect -1338 43094 -1334 43164
rect -1314 43094 -1310 43164
rect -1290 43094 -1286 43164
rect -1266 43094 -1262 43164
rect -1242 43094 -1238 43164
rect -1218 43094 -1214 43164
rect -1194 43115 -1190 43164
rect -2393 43092 -1197 43094
rect -2371 43022 -2366 43092
rect -2348 43022 -2343 43092
rect -2325 43088 -2320 43092
rect -2309 43090 -2301 43092
rect -2317 43088 -2309 43090
rect -2325 43076 -2317 43088
rect -2325 43022 -2320 43076
rect -2317 43074 -2309 43076
rect -2092 43062 -2062 43064
rect -2094 43058 -2062 43062
rect -2309 43028 -2301 43034
rect -2317 43022 -2309 43028
rect -2000 43022 -1992 43092
rect -1655 43090 -1647 43092
rect -1663 43088 -1655 43090
rect -1671 43076 -1663 43088
rect -1663 43074 -1655 43076
rect -1854 43062 -1806 43064
rect -1854 43058 -1680 43062
rect -1655 43028 -1647 43034
rect -1663 43022 -1655 43028
rect -1642 43022 -1637 43092
rect -1619 43022 -1614 43092
rect -1530 43022 -1526 43092
rect -1506 43022 -1502 43092
rect -1482 43022 -1478 43092
rect -1458 43022 -1454 43092
rect -1434 43022 -1430 43092
rect -1410 43022 -1406 43092
rect -1386 43022 -1382 43092
rect -1362 43091 -1358 43092
rect -1362 43043 -1355 43091
rect -1362 43022 -1358 43043
rect -1338 43022 -1334 43092
rect -1314 43022 -1310 43092
rect -1290 43022 -1286 43092
rect -1266 43022 -1262 43092
rect -1242 43022 -1238 43092
rect -1218 43022 -1214 43092
rect -1211 43091 -1197 43092
rect -1194 43091 -1187 43115
rect -1194 43022 -1190 43091
rect -1170 43022 -1166 43164
rect -1146 43022 -1142 43164
rect -1122 43022 -1118 43164
rect -1098 43022 -1094 43164
rect -1074 43022 -1070 43164
rect -1050 43022 -1046 43164
rect -1037 43085 -1032 43095
rect -1026 43085 -1022 43164
rect -1027 43071 -1022 43085
rect -1026 43022 -1022 43071
rect -1002 43022 -998 43164
rect -978 43022 -974 43164
rect -954 43022 -950 43164
rect -930 43022 -926 43164
rect -906 43022 -902 43164
rect -893 43037 -888 43047
rect -882 43037 -878 43164
rect -883 43023 -878 43037
rect -893 43022 -859 43023
rect -2393 43020 -859 43022
rect -2371 42926 -2366 43020
rect -2348 42926 -2343 43020
rect -2325 42958 -2320 43020
rect -2317 43018 -2309 43020
rect -2000 43019 -1966 43020
rect -2000 43018 -1982 43019
rect -1663 43018 -1655 43020
rect -2028 43010 -2018 43012
rect -2309 43000 -2301 43006
rect -2091 43000 -2061 43007
rect -2317 42990 -2309 43000
rect -2044 42998 -2028 43000
rect -2026 42998 -2014 43010
rect -2084 42992 -2061 42998
rect -2044 42996 -2014 42998
rect -2292 42982 -2054 42991
rect -2325 42950 -2317 42958
rect -2325 42930 -2320 42950
rect -2317 42942 -2309 42950
rect -2325 42926 -2317 42930
rect -2000 42926 -1992 43018
rect -1982 43017 -1966 43018
rect -1980 43000 -1932 43007
rect -1655 43000 -1647 43006
rect -1846 42982 -1680 42991
rect -1663 42990 -1655 43000
rect -1671 42950 -1663 42958
rect -1663 42942 -1655 42950
rect -1671 42926 -1663 42930
rect -1642 42926 -1637 43020
rect -1619 42926 -1614 43020
rect -1530 42926 -1526 43020
rect -1506 42926 -1502 43020
rect -1482 42926 -1478 43020
rect -1458 42926 -1454 43020
rect -1434 42926 -1430 43020
rect -1410 42926 -1406 43020
rect -1386 42926 -1382 43020
rect -1362 42926 -1358 43020
rect -1338 42926 -1334 43020
rect -1314 42926 -1310 43020
rect -1290 42926 -1286 43020
rect -1266 42926 -1262 43020
rect -1242 42926 -1238 43020
rect -1218 42926 -1214 43020
rect -1194 42926 -1190 43020
rect -1170 42926 -1166 43020
rect -1146 42926 -1142 43020
rect -1122 42926 -1118 43020
rect -1098 42926 -1094 43020
rect -1074 42926 -1070 43020
rect -1050 42926 -1046 43020
rect -1026 42926 -1022 43020
rect -1002 43019 -998 43020
rect -1002 42995 -995 43019
rect -1002 42926 -998 42995
rect -978 42926 -974 43020
rect -954 42926 -950 43020
rect -930 42926 -926 43020
rect -906 42926 -902 43020
rect -893 43013 -888 43020
rect -883 42999 -878 43013
rect -882 42926 -878 42999
rect -858 42971 -854 43164
rect -2393 42924 -861 42926
rect -2371 42878 -2366 42924
rect -2348 42878 -2343 42924
rect -2325 42916 -2317 42924
rect -2018 42923 -2004 42924
rect -2000 42923 -1992 42924
rect -2072 42922 -1928 42923
rect -2072 42916 -2053 42922
rect -2325 42900 -2320 42916
rect -2317 42914 -2309 42916
rect -2309 42902 -2301 42914
rect -2092 42907 -2062 42912
rect -2317 42900 -2309 42902
rect -2325 42888 -2317 42900
rect -2098 42894 -2096 42905
rect -2092 42894 -2084 42907
rect -2000 42906 -1992 42922
rect -1972 42916 -1928 42922
rect -1924 42916 -1918 42924
rect -1671 42916 -1663 42924
rect -1663 42914 -1655 42916
rect -2083 42896 -2062 42905
rect -2027 42904 -1992 42906
rect -2018 42896 -2002 42904
rect -2000 42896 -1992 42904
rect -2100 42889 -2096 42894
rect -2083 42889 -2053 42894
rect -2003 42892 -1990 42896
rect -1972 42894 -1964 42903
rect -1928 42902 -1924 42905
rect -1655 42902 -1647 42914
rect -1663 42900 -1655 42902
rect -2325 42878 -2320 42888
rect -2317 42886 -2309 42888
rect -2309 42878 -2301 42886
rect -2004 42882 -2003 42892
rect -2062 42878 -2012 42880
rect -2000 42878 -1992 42892
rect -1972 42889 -1924 42894
rect -1864 42889 -1796 42895
rect -1671 42888 -1663 42900
rect -1663 42886 -1655 42888
rect -1864 42878 -1796 42879
rect -1655 42878 -1647 42886
rect -1642 42878 -1637 42924
rect -1619 42878 -1614 42924
rect -1530 42878 -1526 42924
rect -1506 42878 -1502 42924
rect -1482 42878 -1478 42924
rect -1458 42878 -1454 42924
rect -1434 42878 -1430 42924
rect -1410 42878 -1406 42924
rect -1386 42878 -1382 42924
rect -1362 42878 -1358 42924
rect -1338 42878 -1334 42924
rect -1314 42878 -1310 42924
rect -1290 42878 -1286 42924
rect -1266 42878 -1262 42924
rect -1242 42878 -1238 42924
rect -1218 42878 -1214 42924
rect -1194 42878 -1190 42924
rect -1170 42878 -1166 42924
rect -1146 42878 -1142 42924
rect -1122 42878 -1118 42924
rect -1098 42878 -1094 42924
rect -1074 42878 -1070 42924
rect -1050 42878 -1046 42924
rect -1026 42878 -1022 42924
rect -1002 42878 -998 42924
rect -978 42878 -974 42924
rect -954 42878 -950 42924
rect -930 42878 -926 42924
rect -906 42878 -902 42924
rect -882 42878 -878 42924
rect -875 42923 -861 42924
rect -858 42923 -851 42971
rect -858 42878 -854 42923
rect -834 42878 -830 43164
rect -810 42878 -806 43164
rect -786 42878 -782 43164
rect -762 42878 -758 43164
rect -738 42878 -734 43164
rect -725 42965 -720 42975
rect -714 42965 -710 43164
rect -715 42951 -710 42965
rect -714 42878 -710 42951
rect -690 42899 -686 43164
rect -666 42951 -662 43164
rect -677 42950 -643 42951
rect -642 42950 -638 43164
rect -618 42950 -614 43164
rect -594 42950 -590 43164
rect -581 43109 -576 43119
rect -570 43109 -566 43164
rect -571 43095 -566 43109
rect -570 42950 -566 43095
rect -546 43043 -542 43164
rect -546 43019 -539 43043
rect -546 42950 -542 43019
rect -522 42950 -518 43164
rect -498 42950 -494 43164
rect -474 42950 -470 43164
rect -450 42950 -446 43164
rect -426 42950 -422 43164
rect -413 42965 -408 42975
rect -402 42965 -398 43164
rect -403 42951 -398 42965
rect -378 42950 -374 43164
rect -354 42950 -350 43164
rect -330 42950 -326 43164
rect -306 42950 -302 43164
rect -282 42950 -278 43164
rect -258 42950 -254 43164
rect -234 42950 -230 43164
rect -210 42950 -206 43164
rect -186 42950 -182 43164
rect -162 42950 -158 43164
rect -138 42950 -134 43164
rect -114 42950 -110 43164
rect -90 42950 -86 43164
rect -66 42950 -62 43164
rect -42 42950 -38 43164
rect -18 42950 -14 43164
rect 6 42950 10 43164
rect 30 42950 34 43164
rect 54 42950 58 43164
rect 78 42950 82 43164
rect 102 42950 106 43164
rect 109 43163 123 43164
rect 115 43157 120 43163
rect 125 43143 130 43157
rect 126 42950 130 43143
rect 139 43037 144 43047
rect 149 43023 154 43037
rect 150 42950 154 43023
rect 173 42951 181 42965
rect -677 42948 171 42950
rect -677 42941 -672 42948
rect -666 42941 -662 42948
rect -667 42927 -662 42941
rect -2393 42876 -693 42878
rect -2371 42830 -2366 42876
rect -2348 42830 -2343 42876
rect -2325 42872 -2320 42876
rect -2309 42874 -2301 42876
rect -2317 42872 -2309 42874
rect -2325 42860 -2317 42872
rect -2325 42830 -2320 42860
rect -2317 42858 -2309 42860
rect -2092 42846 -2062 42848
rect -2094 42842 -2062 42846
rect -2000 42830 -1992 42876
rect -1655 42874 -1647 42876
rect -1663 42872 -1655 42874
rect -1671 42860 -1663 42872
rect -1663 42858 -1655 42860
rect -1854 42846 -1806 42848
rect -1854 42842 -1680 42846
rect -1642 42830 -1637 42876
rect -1619 42830 -1614 42876
rect -1530 42830 -1526 42876
rect -1506 42830 -1502 42876
rect -1482 42830 -1478 42876
rect -1458 42830 -1454 42876
rect -1434 42830 -1430 42876
rect -1410 42830 -1406 42876
rect -1386 42830 -1382 42876
rect -1362 42830 -1358 42876
rect -1338 42830 -1334 42876
rect -1314 42830 -1310 42876
rect -1290 42830 -1286 42876
rect -1266 42830 -1262 42876
rect -1242 42830 -1238 42876
rect -1218 42830 -1214 42876
rect -1194 42830 -1190 42876
rect -1170 42830 -1166 42876
rect -1146 42830 -1142 42876
rect -1122 42830 -1118 42876
rect -1098 42830 -1094 42876
rect -1074 42830 -1070 42876
rect -1050 42830 -1046 42876
rect -1026 42830 -1022 42876
rect -1002 42830 -998 42876
rect -978 42830 -974 42876
rect -954 42830 -950 42876
rect -930 42830 -926 42876
rect -906 42830 -902 42876
rect -882 42830 -878 42876
rect -858 42830 -854 42876
rect -834 42830 -830 42876
rect -810 42830 -806 42876
rect -786 42830 -782 42876
rect -762 42830 -758 42876
rect -738 42830 -734 42876
rect -714 42830 -710 42876
rect -707 42875 -693 42876
rect -690 42875 -683 42899
rect -677 42893 -672 42903
rect -667 42879 -662 42893
rect -690 42830 -686 42875
rect -666 42830 -662 42879
rect -642 42875 -638 42948
rect -642 42851 -635 42875
rect -618 42830 -614 42948
rect -594 42830 -590 42948
rect -570 42830 -566 42948
rect -546 42830 -542 42948
rect -522 42832 -518 42948
rect -509 42893 -504 42903
rect -498 42893 -494 42948
rect -499 42879 -494 42893
rect -509 42854 -475 42855
rect -474 42854 -470 42948
rect -450 42854 -446 42948
rect -426 42854 -422 42948
rect -413 42917 -408 42927
rect -403 42903 -398 42917
rect -402 42854 -398 42903
rect -378 42899 -374 42948
rect -378 42878 -371 42899
rect -354 42878 -350 42948
rect -330 42878 -326 42948
rect -306 42878 -302 42948
rect -282 42878 -278 42948
rect -258 42878 -254 42948
rect -234 42878 -230 42948
rect -210 42878 -206 42948
rect -186 42878 -182 42948
rect -162 42878 -158 42948
rect -138 42878 -134 42948
rect -114 42878 -110 42948
rect -90 42878 -86 42948
rect -66 42878 -62 42948
rect -42 42878 -38 42948
rect -18 42878 -14 42948
rect -5 42917 0 42927
rect 6 42917 10 42948
rect 5 42903 10 42917
rect -5 42878 29 42879
rect -395 42876 29 42878
rect -395 42875 -381 42876
rect -378 42875 -371 42876
rect -354 42854 -350 42876
rect -330 42854 -326 42876
rect -306 42854 -302 42876
rect -282 42854 -278 42876
rect -258 42854 -254 42876
rect -234 42854 -230 42876
rect -210 42854 -206 42876
rect -186 42854 -182 42876
rect -162 42854 -158 42876
rect -138 42854 -134 42876
rect -114 42854 -110 42876
rect -90 42854 -86 42876
rect -66 42854 -62 42876
rect -42 42854 -38 42876
rect -18 42854 -14 42876
rect -5 42869 0 42876
rect 5 42855 10 42869
rect 6 42854 10 42855
rect 30 42854 34 42948
rect 54 42854 58 42948
rect 78 42854 82 42948
rect 102 42854 106 42948
rect 126 42854 130 42948
rect 150 42854 154 42948
rect 157 42947 171 42948
rect 174 42947 181 42951
rect 174 42854 178 42947
rect 198 42875 205 42899
rect 198 42854 202 42875
rect -509 42852 219 42854
rect -509 42845 -504 42852
rect -499 42842 -494 42845
rect -499 42831 -494 42832
rect -533 42830 -499 42831
rect -2393 42828 -499 42830
rect -2371 42806 -2366 42828
rect -2348 42806 -2343 42828
rect -2325 42806 -2320 42828
rect -2072 42826 -2036 42827
rect -2072 42820 -2054 42826
rect -2309 42812 -2301 42820
rect -2317 42806 -2309 42812
rect -2092 42811 -2062 42816
rect -2000 42807 -1992 42828
rect -1938 42827 -1906 42828
rect -1920 42826 -1906 42827
rect -1806 42820 -1680 42826
rect -1854 42811 -1806 42816
rect -1655 42812 -1647 42820
rect -1982 42807 -1966 42808
rect -2000 42806 -1966 42807
rect -1846 42806 -1806 42809
rect -1663 42806 -1655 42812
rect -1642 42806 -1637 42828
rect -1619 42806 -1614 42828
rect -1530 42806 -1526 42828
rect -1506 42806 -1502 42828
rect -1482 42806 -1478 42828
rect -1458 42806 -1454 42828
rect -1434 42806 -1430 42828
rect -1410 42806 -1406 42828
rect -1386 42806 -1382 42828
rect -1362 42806 -1358 42828
rect -1338 42806 -1334 42828
rect -1314 42806 -1310 42828
rect -1290 42806 -1286 42828
rect -1266 42806 -1262 42828
rect -1242 42806 -1238 42828
rect -1218 42806 -1214 42828
rect -1194 42806 -1190 42828
rect -1170 42806 -1166 42828
rect -1146 42806 -1142 42828
rect -1122 42806 -1118 42828
rect -1098 42806 -1094 42828
rect -1074 42806 -1070 42828
rect -1050 42806 -1046 42828
rect -1026 42806 -1022 42828
rect -1002 42806 -998 42828
rect -978 42806 -974 42828
rect -954 42806 -950 42828
rect -930 42806 -926 42828
rect -906 42806 -902 42828
rect -882 42806 -878 42828
rect -858 42806 -854 42828
rect -834 42806 -830 42828
rect -810 42806 -806 42828
rect -786 42806 -782 42828
rect -762 42806 -758 42828
rect -738 42807 -734 42828
rect -749 42806 -715 42807
rect -714 42806 -710 42828
rect -690 42806 -686 42828
rect -666 42806 -662 42828
rect -2393 42804 -645 42806
rect -2371 42782 -2366 42804
rect -2348 42782 -2343 42804
rect -2325 42782 -2320 42804
rect -2000 42802 -1966 42804
rect -2309 42784 -2301 42792
rect -2062 42791 -2054 42798
rect -2092 42784 -2084 42791
rect -2062 42784 -2026 42786
rect -2317 42782 -2309 42784
rect -2062 42782 -2012 42784
rect -2000 42782 -1992 42802
rect -1982 42801 -1966 42802
rect -1846 42800 -1806 42804
rect -1846 42793 -1798 42798
rect -1806 42791 -1798 42793
rect -1854 42789 -1846 42791
rect -1854 42784 -1806 42789
rect -1655 42784 -1647 42792
rect -1864 42782 -1796 42783
rect -1663 42782 -1655 42784
rect -1642 42782 -1637 42804
rect -1619 42782 -1614 42804
rect -1530 42782 -1526 42804
rect -1506 42782 -1502 42804
rect -1482 42782 -1478 42804
rect -1458 42782 -1454 42804
rect -1434 42782 -1430 42804
rect -1410 42782 -1406 42804
rect -1386 42782 -1382 42804
rect -1362 42782 -1358 42804
rect -1338 42782 -1334 42804
rect -1314 42782 -1310 42804
rect -1290 42782 -1286 42804
rect -1266 42782 -1262 42804
rect -1242 42782 -1238 42804
rect -1218 42782 -1214 42804
rect -1194 42782 -1190 42804
rect -1170 42782 -1166 42804
rect -1146 42782 -1142 42804
rect -1122 42782 -1118 42804
rect -1098 42782 -1094 42804
rect -1074 42782 -1070 42804
rect -1050 42782 -1046 42804
rect -1026 42782 -1022 42804
rect -1002 42782 -998 42804
rect -978 42782 -974 42804
rect -954 42782 -950 42804
rect -930 42782 -926 42804
rect -906 42782 -902 42804
rect -882 42782 -878 42804
rect -858 42782 -854 42804
rect -834 42782 -830 42804
rect -810 42782 -806 42804
rect -786 42782 -782 42804
rect -762 42782 -758 42804
rect -749 42797 -744 42804
rect -738 42797 -734 42804
rect -739 42783 -734 42797
rect -749 42782 -715 42783
rect -2393 42780 -715 42782
rect -2371 42710 -2366 42780
rect -2348 42710 -2343 42780
rect -2325 42710 -2320 42780
rect -2317 42776 -2309 42780
rect -2062 42776 -2054 42780
rect -2154 42772 -2138 42774
rect -2057 42772 -2054 42776
rect -2292 42766 -2054 42772
rect -2052 42766 -2044 42776
rect -2092 42750 -2062 42752
rect -2094 42746 -2062 42750
rect -2309 42716 -2301 42722
rect -2317 42710 -2309 42716
rect -2000 42710 -1992 42780
rect -1846 42773 -1806 42780
rect -1663 42776 -1655 42780
rect -1846 42766 -1680 42772
rect -1854 42750 -1806 42752
rect -1854 42746 -1680 42750
rect -1655 42716 -1647 42722
rect -1663 42710 -1655 42716
rect -1642 42710 -1637 42780
rect -1619 42710 -1614 42780
rect -1530 42710 -1526 42780
rect -1506 42710 -1502 42780
rect -1482 42710 -1478 42780
rect -1458 42710 -1454 42780
rect -1434 42710 -1430 42780
rect -1410 42710 -1406 42780
rect -1386 42710 -1382 42780
rect -1362 42710 -1358 42780
rect -1338 42710 -1334 42780
rect -1314 42710 -1310 42780
rect -1290 42710 -1286 42780
rect -1266 42710 -1262 42780
rect -1242 42710 -1238 42780
rect -1218 42710 -1214 42780
rect -1194 42710 -1190 42780
rect -1170 42710 -1166 42780
rect -1146 42710 -1142 42780
rect -1122 42710 -1118 42780
rect -1098 42710 -1094 42780
rect -1074 42710 -1070 42780
rect -1050 42710 -1046 42780
rect -1026 42710 -1022 42780
rect -1002 42710 -998 42780
rect -978 42710 -974 42780
rect -954 42710 -950 42780
rect -930 42710 -926 42780
rect -906 42710 -902 42780
rect -882 42710 -878 42780
rect -858 42710 -854 42780
rect -834 42710 -830 42780
rect -810 42710 -806 42780
rect -786 42710 -782 42780
rect -762 42710 -758 42780
rect -749 42773 -744 42780
rect -739 42759 -734 42773
rect -738 42710 -734 42759
rect -714 42731 -710 42804
rect -714 42710 -707 42731
rect -690 42710 -686 42804
rect -666 42710 -662 42804
rect -659 42803 -645 42804
rect -642 42803 -635 42827
rect -642 42710 -638 42803
rect -618 42710 -614 42828
rect -594 42710 -590 42828
rect -570 42710 -566 42828
rect -546 42710 -542 42828
rect -533 42821 -528 42828
rect -474 42827 -470 42852
rect -523 42807 -518 42821
rect -533 42797 -528 42807
rect -523 42783 -518 42797
rect -522 42710 -518 42783
rect -498 42766 -494 42808
rect -474 42803 -467 42827
rect -474 42755 -467 42779
rect -498 42742 -491 42755
rect -2393 42708 -501 42710
rect -2371 42614 -2366 42708
rect -2348 42614 -2343 42708
rect -2325 42646 -2320 42708
rect -2317 42706 -2309 42708
rect -2000 42707 -1966 42708
rect -2000 42706 -1982 42707
rect -1663 42706 -1655 42708
rect -2028 42698 -2018 42700
rect -2309 42688 -2301 42694
rect -2091 42688 -2061 42695
rect -2317 42678 -2309 42688
rect -2044 42686 -2028 42688
rect -2026 42686 -2014 42698
rect -2084 42680 -2061 42686
rect -2044 42684 -2014 42686
rect -2292 42670 -2054 42679
rect -2325 42638 -2317 42646
rect -2325 42618 -2320 42638
rect -2317 42630 -2309 42638
rect -2325 42614 -2317 42618
rect -2000 42614 -1992 42706
rect -1982 42705 -1966 42706
rect -1980 42688 -1932 42695
rect -1655 42688 -1647 42694
rect -1846 42670 -1680 42679
rect -1663 42678 -1655 42688
rect -1671 42638 -1663 42646
rect -1663 42630 -1655 42638
rect -1926 42614 -1892 42617
rect -1671 42614 -1663 42618
rect -1642 42614 -1637 42708
rect -1619 42614 -1614 42708
rect -1530 42614 -1526 42708
rect -1506 42614 -1502 42708
rect -1482 42614 -1478 42708
rect -1458 42614 -1454 42708
rect -1434 42614 -1430 42708
rect -1410 42614 -1406 42708
rect -1386 42614 -1382 42708
rect -1362 42614 -1358 42708
rect -1338 42614 -1334 42708
rect -1314 42614 -1310 42708
rect -1290 42614 -1286 42708
rect -1266 42614 -1262 42708
rect -1242 42614 -1238 42708
rect -1218 42614 -1214 42708
rect -1194 42614 -1190 42708
rect -1170 42614 -1166 42708
rect -1146 42614 -1142 42708
rect -1133 42653 -1128 42663
rect -1122 42653 -1118 42708
rect -1123 42639 -1118 42653
rect -1122 42614 -1118 42639
rect -1109 42629 -1104 42639
rect -1098 42629 -1094 42708
rect -1099 42615 -1094 42629
rect -1109 42614 -1075 42615
rect -2393 42612 -1075 42614
rect -2371 42566 -2366 42612
rect -2348 42566 -2343 42612
rect -2325 42606 -2317 42612
rect -2053 42610 -1972 42612
rect -2325 42590 -2320 42606
rect -2317 42602 -2309 42606
rect -2069 42602 -2068 42603
rect -2309 42590 -2301 42602
rect -2069 42595 -2038 42602
rect -2069 42593 -2068 42595
rect -2000 42594 -1992 42610
rect -1926 42607 -1924 42612
rect -1916 42604 -1914 42607
rect -1671 42606 -1663 42612
rect -1982 42594 -1916 42603
rect -1663 42602 -1655 42606
rect -2325 42578 -2317 42590
rect -2068 42587 -2053 42593
rect -2027 42592 -1992 42594
rect -2076 42578 -2053 42585
rect -2011 42584 -2002 42592
rect -2000 42584 -1992 42592
rect -1655 42590 -1647 42602
rect -2003 42582 -1992 42584
rect -2325 42566 -2320 42578
rect -2317 42574 -2309 42578
rect -2309 42566 -2301 42574
rect -2015 42570 -2003 42582
rect -2000 42566 -1992 42582
rect -1972 42578 -1924 42585
rect -1862 42577 -1680 42586
rect -1671 42578 -1663 42590
rect -1663 42574 -1655 42578
rect -1976 42566 -1940 42567
rect -1655 42566 -1647 42574
rect -1642 42566 -1637 42612
rect -1619 42566 -1614 42612
rect -1530 42566 -1526 42612
rect -1506 42566 -1502 42612
rect -1482 42566 -1478 42612
rect -1458 42566 -1454 42612
rect -1434 42566 -1430 42612
rect -1410 42566 -1406 42612
rect -1386 42566 -1382 42612
rect -1362 42566 -1358 42612
rect -1338 42566 -1334 42612
rect -1314 42566 -1310 42612
rect -1290 42566 -1286 42612
rect -1266 42566 -1262 42612
rect -1242 42566 -1238 42612
rect -1218 42566 -1214 42612
rect -1194 42566 -1190 42612
rect -1170 42566 -1166 42612
rect -1146 42566 -1142 42612
rect -1122 42566 -1118 42612
rect -1109 42605 -1104 42612
rect -1099 42591 -1094 42605
rect -1098 42587 -1094 42591
rect -2393 42564 -1101 42566
rect -2371 42470 -2366 42564
rect -2348 42470 -2343 42564
rect -2325 42562 -2320 42564
rect -2309 42562 -2301 42564
rect -2325 42550 -2317 42562
rect -2325 42530 -2320 42550
rect -2317 42546 -2309 42550
rect -2325 42522 -2317 42530
rect -2060 42524 -2030 42527
rect -2325 42470 -2320 42522
rect -2317 42514 -2309 42522
rect -2060 42511 -2038 42522
rect -2033 42515 -2030 42524
rect -2028 42520 -2027 42524
rect -2068 42506 -2038 42509
rect -2309 42474 -2301 42482
rect -2317 42470 -2309 42474
rect -2000 42470 -1992 42564
rect -1655 42562 -1647 42564
rect -1671 42550 -1663 42562
rect -1663 42546 -1655 42550
rect -1912 42539 -1884 42541
rect -1852 42533 -1804 42537
rect -1844 42524 -1796 42527
rect -1671 42522 -1663 42530
rect -1844 42511 -1804 42522
rect -1663 42514 -1655 42522
rect -1852 42506 -1680 42510
rect -1655 42474 -1647 42482
rect -1663 42470 -1655 42474
rect -1642 42470 -1637 42564
rect -1619 42470 -1614 42564
rect -1530 42470 -1526 42564
rect -1506 42470 -1502 42564
rect -1482 42470 -1478 42564
rect -1458 42470 -1454 42564
rect -1434 42470 -1430 42564
rect -1410 42495 -1406 42564
rect -1421 42494 -1387 42495
rect -1386 42494 -1382 42564
rect -1362 42494 -1358 42564
rect -1338 42494 -1334 42564
rect -1314 42494 -1310 42564
rect -1290 42494 -1286 42564
rect -1266 42494 -1262 42564
rect -1242 42494 -1238 42564
rect -1218 42494 -1214 42564
rect -1194 42494 -1190 42564
rect -1181 42533 -1176 42543
rect -1170 42533 -1166 42564
rect -1171 42519 -1166 42533
rect -1170 42494 -1166 42519
rect -1146 42494 -1142 42564
rect -1122 42494 -1118 42564
rect -1115 42563 -1101 42564
rect -1098 42563 -1091 42587
rect -1074 42563 -1070 42708
rect -1098 42494 -1094 42563
rect -1074 42515 -1067 42563
rect -1074 42494 -1070 42515
rect -1050 42494 -1046 42708
rect -1026 42494 -1022 42708
rect -1002 42494 -998 42708
rect -978 42494 -974 42708
rect -954 42494 -950 42708
rect -930 42494 -926 42708
rect -906 42494 -902 42708
rect -882 42494 -878 42708
rect -858 42494 -854 42708
rect -834 42494 -830 42708
rect -810 42494 -806 42708
rect -786 42494 -782 42708
rect -762 42494 -758 42708
rect -738 42494 -734 42708
rect -731 42707 -717 42708
rect -714 42683 -707 42708
rect -714 42494 -710 42683
rect -690 42494 -686 42708
rect -666 42494 -662 42708
rect -642 42494 -638 42708
rect -618 42494 -614 42708
rect -594 42494 -590 42708
rect -581 42557 -576 42567
rect -570 42557 -566 42708
rect -557 42581 -552 42591
rect -546 42581 -542 42708
rect -547 42567 -542 42581
rect -571 42543 -566 42557
rect -570 42494 -566 42543
rect -546 42494 -542 42567
rect -522 42515 -518 42708
rect -515 42707 -501 42708
rect -498 42707 -491 42732
rect -1421 42492 -525 42494
rect -1421 42485 -1416 42492
rect -1410 42485 -1406 42492
rect -1411 42471 -1406 42485
rect -1421 42470 -1387 42471
rect -2393 42468 -2020 42470
rect -2012 42468 -1387 42470
rect -2371 42374 -2366 42468
rect -2348 42374 -2343 42468
rect -2325 42406 -2320 42468
rect -2317 42466 -2309 42468
rect -2062 42455 -2061 42456
rect -2060 42455 -2049 42468
rect -2309 42446 -2301 42454
rect -2068 42448 -2061 42455
rect -2020 42448 -2012 42460
rect -2317 42438 -2309 42446
rect -2124 42439 -2108 42441
rect -2060 42439 -2049 42448
rect -2020 42446 -2004 42448
rect -2000 42446 -1992 42468
rect -1972 42466 -1958 42468
rect -1663 42466 -1655 42468
rect -1958 42465 -1942 42466
rect -1980 42448 -1932 42455
rect -1655 42446 -1647 42454
rect -2292 42438 -2049 42439
rect -2036 42438 -2030 42446
rect -2020 42444 -1992 42446
rect -2292 42431 -2030 42438
rect -2292 42430 -2049 42431
rect -2031 42430 -2030 42431
rect -2026 42430 -2020 42436
rect -2325 42398 -2317 42406
rect -2325 42378 -2320 42398
rect -2317 42390 -2309 42398
rect -2325 42374 -2317 42378
rect -2000 42374 -1992 42444
rect -1844 42430 -1680 42439
rect -1663 42438 -1655 42446
rect -1671 42398 -1663 42406
rect -1663 42390 -1655 42398
rect -1671 42374 -1663 42378
rect -1642 42374 -1637 42468
rect -1619 42374 -1614 42468
rect -1530 42374 -1526 42468
rect -1506 42374 -1502 42468
rect -1482 42374 -1478 42468
rect -1458 42374 -1454 42468
rect -1434 42374 -1430 42468
rect -1421 42461 -1416 42468
rect -1411 42447 -1406 42461
rect -1410 42374 -1406 42447
rect -1386 42419 -1382 42492
rect -2393 42372 -1389 42374
rect -2371 42326 -2366 42372
rect -2348 42326 -2343 42372
rect -2325 42364 -2317 42372
rect -2018 42371 -2004 42372
rect -2000 42371 -1992 42372
rect -2072 42370 -1928 42371
rect -2072 42364 -2053 42370
rect -2325 42348 -2320 42364
rect -2317 42362 -2309 42364
rect -2309 42350 -2301 42362
rect -2092 42355 -2062 42360
rect -2317 42348 -2309 42350
rect -2325 42336 -2317 42348
rect -2098 42342 -2096 42353
rect -2092 42342 -2084 42355
rect -2000 42354 -1992 42370
rect -1972 42364 -1928 42370
rect -1924 42364 -1918 42372
rect -1671 42364 -1663 42372
rect -1663 42362 -1655 42364
rect -2083 42344 -2062 42353
rect -2027 42352 -1992 42354
rect -2018 42344 -2002 42352
rect -2000 42344 -1992 42352
rect -2100 42337 -2096 42342
rect -2083 42337 -2053 42342
rect -2003 42340 -1990 42344
rect -1972 42342 -1964 42351
rect -1928 42350 -1924 42353
rect -1655 42350 -1647 42362
rect -1663 42348 -1655 42350
rect -2325 42326 -2320 42336
rect -2317 42334 -2309 42336
rect -2309 42326 -2301 42334
rect -2004 42330 -2003 42340
rect -2062 42326 -2012 42328
rect -2000 42326 -1992 42340
rect -1972 42337 -1924 42342
rect -1864 42337 -1796 42343
rect -1671 42336 -1663 42348
rect -1663 42334 -1655 42336
rect -1864 42326 -1796 42327
rect -1655 42326 -1647 42334
rect -1642 42326 -1637 42372
rect -1619 42326 -1614 42372
rect -1530 42327 -1526 42372
rect -1541 42326 -1507 42327
rect -2393 42324 -1507 42326
rect -2371 42254 -2366 42324
rect -2348 42254 -2343 42324
rect -2325 42320 -2320 42324
rect -2309 42322 -2301 42324
rect -2317 42320 -2309 42322
rect -2325 42308 -2317 42320
rect -2325 42254 -2320 42308
rect -2317 42306 -2309 42308
rect -2092 42294 -2062 42296
rect -2094 42290 -2062 42294
rect -2309 42260 -2301 42266
rect -2317 42254 -2309 42260
rect -2000 42254 -1992 42324
rect -1655 42322 -1647 42324
rect -1663 42320 -1655 42322
rect -1671 42308 -1663 42320
rect -1663 42306 -1655 42308
rect -1854 42294 -1806 42296
rect -1854 42290 -1680 42294
rect -1655 42260 -1647 42266
rect -1663 42254 -1655 42260
rect -1642 42254 -1637 42324
rect -1619 42254 -1614 42324
rect -1541 42317 -1536 42324
rect -1530 42317 -1526 42324
rect -1531 42303 -1526 42317
rect -1530 42254 -1526 42303
rect -1506 42254 -1502 42372
rect -1482 42254 -1478 42372
rect -1458 42254 -1454 42372
rect -1434 42254 -1430 42372
rect -1410 42254 -1406 42372
rect -1403 42371 -1389 42372
rect -1386 42371 -1379 42419
rect -1386 42254 -1382 42371
rect -1362 42254 -1358 42492
rect -1338 42254 -1334 42492
rect -1314 42254 -1310 42492
rect -1290 42254 -1286 42492
rect -1266 42254 -1262 42492
rect -1242 42254 -1238 42492
rect -1218 42254 -1214 42492
rect -1194 42254 -1190 42492
rect -1181 42341 -1176 42351
rect -1170 42341 -1166 42492
rect -1171 42327 -1166 42341
rect -1170 42254 -1166 42327
rect -1146 42467 -1142 42492
rect -1146 42443 -1139 42467
rect -1146 42275 -1142 42443
rect -2393 42252 -1149 42254
rect -2371 42038 -2366 42252
rect -2348 42038 -2343 42252
rect -2325 42190 -2320 42252
rect -2317 42250 -2309 42252
rect -2000 42251 -1966 42252
rect -2000 42250 -1982 42251
rect -1663 42250 -1655 42252
rect -2028 42242 -2018 42244
rect -2309 42232 -2301 42238
rect -2091 42232 -2061 42239
rect -2317 42222 -2309 42232
rect -2044 42230 -2028 42232
rect -2026 42230 -2014 42242
rect -2084 42224 -2061 42230
rect -2044 42228 -2014 42230
rect -2292 42214 -2054 42223
rect -2325 42182 -2317 42190
rect -2325 42162 -2320 42182
rect -2317 42174 -2309 42182
rect -2325 42146 -2317 42162
rect -2325 42130 -2320 42146
rect -2309 42134 -2301 42146
rect -2317 42130 -2309 42134
rect -2103 42130 -2096 42132
rect -2083 42130 -2053 42132
rect -2325 42118 -2317 42130
rect -2103 42121 -2053 42130
rect -2018 42128 -2017 42134
rect -2003 42128 -2002 42130
rect -2026 42124 -2017 42128
rect -2325 42102 -2320 42118
rect -2309 42106 -2301 42118
rect -2017 42114 -2012 42124
rect -2317 42102 -2309 42106
rect -2325 42090 -2317 42102
rect -2325 42070 -2320 42090
rect -2325 42062 -2317 42070
rect -2325 42042 -2320 42062
rect -2317 42054 -2309 42062
rect -2325 42038 -2317 42042
rect -2000 42038 -1992 42250
rect -1982 42249 -1966 42250
rect -1980 42232 -1932 42239
rect -1655 42232 -1647 42238
rect -1846 42214 -1680 42223
rect -1663 42222 -1655 42232
rect -1671 42182 -1663 42190
rect -1663 42174 -1655 42182
rect -1671 42146 -1663 42162
rect -1655 42134 -1647 42146
rect -1972 42130 -1924 42132
rect -1663 42130 -1655 42134
rect -1972 42121 -1922 42130
rect -1671 42118 -1663 42130
rect -1655 42106 -1647 42118
rect -1663 42102 -1655 42106
rect -1671 42090 -1663 42102
rect -1671 42062 -1663 42070
rect -1663 42054 -1655 42062
rect -1671 42038 -1663 42042
rect -1642 42038 -1637 42252
rect -1619 42038 -1614 42252
rect -1530 42038 -1526 42252
rect -1506 42251 -1502 42252
rect -1506 42227 -1499 42251
rect -1506 42038 -1502 42227
rect -1482 42038 -1478 42252
rect -1458 42038 -1454 42252
rect -1434 42038 -1430 42252
rect -1410 42038 -1406 42252
rect -1386 42038 -1382 42252
rect -1362 42038 -1358 42252
rect -1338 42038 -1334 42252
rect -1314 42038 -1310 42252
rect -1290 42038 -1286 42252
rect -1266 42038 -1262 42252
rect -1242 42038 -1238 42252
rect -1218 42038 -1214 42252
rect -1194 42038 -1190 42252
rect -1170 42038 -1166 42252
rect -1163 42251 -1149 42252
rect -1146 42251 -1139 42275
rect -1146 42038 -1142 42251
rect -1122 42038 -1118 42492
rect -1098 42038 -1094 42492
rect -1074 42038 -1070 42492
rect -1050 42038 -1046 42492
rect -1037 42053 -1032 42063
rect -1026 42053 -1022 42492
rect -1027 42039 -1022 42053
rect -1037 42038 -1003 42039
rect -2393 42036 -1003 42038
rect -2371 41990 -2366 42036
rect -2348 41990 -2343 42036
rect -2325 42030 -2317 42036
rect -2018 42034 -2004 42036
rect -2325 42014 -2320 42030
rect -2317 42026 -2309 42030
rect -2069 42028 -2053 42030
rect -2309 42014 -2301 42026
rect -2096 42017 -2095 42023
rect -2000 42018 -1992 42036
rect -1671 42030 -1663 42036
rect -1663 42026 -1655 42030
rect -1977 42019 -1929 42025
rect -2112 42014 -2095 42017
rect -2325 42002 -2317 42014
rect -2325 41990 -2320 42002
rect -2317 41998 -2309 42002
rect -2112 42001 -2096 42014
rect -2059 42010 -2053 42017
rect -2027 42016 -1992 42018
rect -2059 42006 -2045 42010
rect -2018 42008 -2017 42010
rect -2083 42001 -2053 42002
rect -2019 42000 -2017 42004
rect -2309 41990 -2301 41998
rect -2017 41994 -2009 42000
rect -2000 41994 -1992 42016
rect -1972 42002 -1929 42017
rect -1655 42014 -1647 42026
rect -1671 42002 -1663 42014
rect -1972 42001 -1924 42002
rect -1663 41998 -1655 42002
rect -2033 41990 -1992 41994
rect -1655 41990 -1647 41998
rect -1642 41990 -1637 42036
rect -1619 41990 -1614 42036
rect -1530 41990 -1526 42036
rect -1506 41990 -1502 42036
rect -1482 41990 -1478 42036
rect -1458 41990 -1454 42036
rect -1434 41990 -1430 42036
rect -1410 41990 -1406 42036
rect -1386 41990 -1382 42036
rect -1362 41990 -1358 42036
rect -1338 41990 -1334 42036
rect -1314 41990 -1310 42036
rect -1290 41990 -1286 42036
rect -1266 41990 -1262 42036
rect -1242 41990 -1238 42036
rect -1218 41990 -1214 42036
rect -1194 41990 -1190 42036
rect -1170 41990 -1166 42036
rect -1146 41990 -1142 42036
rect -1122 41990 -1118 42036
rect -1098 41990 -1094 42036
rect -1074 41990 -1070 42036
rect -1050 41990 -1046 42036
rect -1037 42029 -1032 42036
rect -1027 42015 -1022 42029
rect -1026 41990 -1022 42015
rect -1002 41990 -998 42492
rect -978 41990 -974 42492
rect -954 41990 -950 42492
rect -930 41990 -926 42492
rect -906 41990 -902 42492
rect -882 41990 -878 42492
rect -858 41990 -854 42492
rect -834 41990 -830 42492
rect -810 41990 -806 42492
rect -786 41991 -782 42492
rect -797 41990 -763 41991
rect -2393 41988 -763 41990
rect -2371 41894 -2366 41988
rect -2348 41894 -2343 41988
rect -2325 41986 -2320 41988
rect -2309 41986 -2301 41988
rect -2325 41974 -2317 41986
rect -2325 41954 -2320 41974
rect -2317 41970 -2309 41974
rect -2325 41946 -2317 41954
rect -2325 41894 -2320 41946
rect -2317 41938 -2309 41946
rect -2117 41937 -2095 41947
rect -2045 41944 -2037 41958
rect -2309 41898 -2301 41908
rect -2087 41904 -2076 41912
rect -2017 41908 -2015 41915
rect -2317 41894 -2309 41898
rect -2092 41896 -2087 41904
rect -2092 41894 -2077 41895
rect -2000 41894 -1992 41988
rect -1655 41986 -1647 41988
rect -1671 41974 -1663 41986
rect -1663 41970 -1655 41974
rect -1969 41937 -1929 41949
rect -1671 41946 -1663 41954
rect -1663 41938 -1655 41946
rect -1655 41898 -1647 41908
rect -1928 41894 -1924 41895
rect -1854 41894 -1680 41895
rect -1663 41894 -1655 41898
rect -1642 41894 -1637 41988
rect -1619 41894 -1614 41988
rect -1530 41894 -1526 41988
rect -1506 41894 -1502 41988
rect -1482 41894 -1478 41988
rect -1458 41943 -1454 41988
rect -1469 41942 -1435 41943
rect -1434 41942 -1430 41988
rect -1410 41942 -1406 41988
rect -1386 41942 -1382 41988
rect -1362 41942 -1358 41988
rect -1338 41942 -1334 41988
rect -1314 41942 -1310 41988
rect -1290 41942 -1286 41988
rect -1266 41942 -1262 41988
rect -1242 41942 -1238 41988
rect -1218 41942 -1214 41988
rect -1194 41942 -1190 41988
rect -1170 41942 -1166 41988
rect -1146 41942 -1142 41988
rect -1122 41942 -1118 41988
rect -1098 41942 -1094 41988
rect -1074 41942 -1070 41988
rect -1050 41942 -1046 41988
rect -1026 41942 -1022 41988
rect -1002 41987 -998 41988
rect -1002 41966 -995 41987
rect -978 41966 -974 41988
rect -954 41967 -950 41988
rect -965 41966 -931 41967
rect -1019 41964 -931 41966
rect -1019 41963 -1005 41964
rect -1469 41940 -1005 41942
rect -1469 41933 -1464 41940
rect -1458 41933 -1454 41940
rect -1459 41919 -1454 41933
rect -1469 41909 -1464 41919
rect -1459 41895 -1454 41909
rect -1458 41894 -1454 41895
rect -1434 41894 -1430 41940
rect -1410 41894 -1406 41940
rect -1386 41894 -1382 41940
rect -1362 41894 -1358 41940
rect -1338 41894 -1334 41940
rect -1314 41894 -1310 41940
rect -1290 41894 -1286 41940
rect -1266 41894 -1262 41940
rect -1242 41894 -1238 41940
rect -1218 41894 -1214 41940
rect -1194 41894 -1190 41940
rect -1170 41894 -1166 41940
rect -1146 41894 -1142 41940
rect -1122 41894 -1118 41940
rect -1098 41894 -1094 41940
rect -1074 41894 -1070 41940
rect -1050 41894 -1046 41940
rect -1026 41894 -1022 41940
rect -1019 41939 -1005 41940
rect -1002 41939 -995 41964
rect -1002 41894 -998 41939
rect -978 41894 -974 41964
rect -965 41957 -960 41964
rect -954 41957 -950 41964
rect -955 41943 -950 41957
rect -954 41894 -950 41943
rect -930 41894 -926 41988
rect -906 41894 -902 41988
rect -882 41894 -878 41988
rect -858 41894 -854 41988
rect -834 41894 -830 41988
rect -810 41894 -806 41988
rect -797 41981 -792 41988
rect -786 41981 -782 41988
rect -787 41967 -782 41981
rect -786 41894 -782 41967
rect -762 41915 -758 42492
rect -2393 41892 -765 41894
rect -2371 41870 -2366 41892
rect -2348 41870 -2343 41892
rect -2325 41870 -2320 41892
rect -2092 41887 -2037 41892
rect -2021 41887 -1969 41892
rect -1921 41887 -1913 41892
rect -1854 41888 -1680 41892
rect -2100 41885 -2092 41886
rect -2309 41870 -2301 41880
rect -2100 41879 -2087 41885
rect -2051 41872 -2026 41874
rect -2062 41870 -2012 41872
rect -2000 41870 -1992 41887
rect -1969 41879 -1921 41886
rect -1969 41870 -1964 41879
rect -1864 41870 -1796 41871
rect -1655 41870 -1647 41880
rect -1642 41870 -1637 41892
rect -1619 41870 -1614 41892
rect -1530 41870 -1526 41892
rect -1506 41870 -1502 41892
rect -1482 41870 -1478 41892
rect -1458 41870 -1454 41892
rect -1434 41870 -1430 41892
rect -1410 41870 -1406 41892
rect -1386 41870 -1382 41892
rect -1362 41870 -1358 41892
rect -1338 41870 -1334 41892
rect -1314 41870 -1310 41892
rect -1290 41870 -1286 41892
rect -1266 41870 -1262 41892
rect -1242 41870 -1238 41892
rect -1218 41870 -1214 41892
rect -1194 41870 -1190 41892
rect -1170 41870 -1166 41892
rect -1146 41870 -1142 41892
rect -1122 41870 -1118 41892
rect -1098 41870 -1094 41892
rect -1074 41870 -1070 41892
rect -1050 41870 -1046 41892
rect -1026 41870 -1022 41892
rect -1002 41870 -998 41892
rect -978 41870 -974 41892
rect -954 41870 -950 41892
rect -930 41891 -926 41892
rect -2393 41868 -933 41870
rect -2371 41798 -2366 41868
rect -2348 41798 -2343 41868
rect -2325 41798 -2320 41868
rect -2317 41864 -2309 41868
rect -2105 41861 -2092 41864
rect -2092 41838 -2062 41840
rect -2094 41834 -2062 41838
rect -2309 41804 -2301 41810
rect -2317 41798 -2309 41804
rect -2000 41798 -1992 41868
rect -1663 41864 -1655 41868
rect -1969 41861 -1921 41864
rect -1854 41838 -1806 41840
rect -1854 41834 -1680 41838
rect -1655 41804 -1647 41810
rect -1663 41798 -1655 41804
rect -1642 41798 -1637 41868
rect -1619 41798 -1614 41868
rect -1530 41798 -1526 41868
rect -1506 41798 -1502 41868
rect -1482 41798 -1478 41868
rect -1458 41798 -1454 41868
rect -1434 41867 -1430 41868
rect -1434 41819 -1427 41867
rect -1434 41798 -1430 41819
rect -1410 41798 -1406 41868
rect -1386 41798 -1382 41868
rect -1362 41798 -1358 41868
rect -1338 41798 -1334 41868
rect -1314 41798 -1310 41868
rect -1290 41798 -1286 41868
rect -1277 41813 -1272 41823
rect -1266 41813 -1262 41868
rect -1267 41799 -1262 41813
rect -1277 41798 -1243 41799
rect -2393 41796 -1243 41798
rect -2371 41342 -2366 41796
rect -2348 41342 -2343 41796
rect -2325 41734 -2320 41796
rect -2317 41794 -2309 41796
rect -2000 41795 -1966 41796
rect -2000 41794 -1982 41795
rect -1663 41794 -1655 41796
rect -2028 41786 -2018 41788
rect -2309 41776 -2301 41782
rect -2091 41776 -2061 41783
rect -2317 41766 -2309 41776
rect -2044 41774 -2028 41776
rect -2026 41774 -2014 41786
rect -2084 41768 -2061 41774
rect -2044 41772 -2014 41774
rect -2292 41758 -2054 41767
rect -2325 41726 -2317 41734
rect -2325 41706 -2320 41726
rect -2317 41718 -2309 41726
rect -2325 41690 -2317 41706
rect -2325 41674 -2320 41690
rect -2309 41678 -2301 41690
rect -2317 41674 -2309 41678
rect -2103 41674 -2096 41676
rect -2083 41674 -2053 41676
rect -2325 41662 -2317 41674
rect -2103 41665 -2053 41674
rect -2018 41672 -2017 41678
rect -2003 41672 -2002 41674
rect -2026 41668 -2017 41672
rect -2325 41646 -2320 41662
rect -2309 41650 -2301 41662
rect -2017 41658 -2012 41668
rect -2317 41646 -2309 41650
rect -2325 41634 -2317 41646
rect -2325 41614 -2320 41634
rect -2325 41606 -2317 41614
rect -2325 41586 -2320 41606
rect -2317 41598 -2309 41606
rect -2325 41570 -2317 41586
rect -2325 41554 -2320 41570
rect -2309 41558 -2301 41570
rect -2317 41554 -2309 41558
rect -2103 41554 -2096 41556
rect -2083 41554 -2053 41556
rect -2325 41542 -2317 41554
rect -2103 41545 -2053 41554
rect -2018 41552 -2017 41558
rect -2003 41552 -2002 41554
rect -2026 41548 -2017 41552
rect -2325 41526 -2320 41542
rect -2309 41530 -2301 41542
rect -2017 41538 -2012 41548
rect -2317 41526 -2309 41530
rect -2325 41514 -2317 41526
rect -2325 41494 -2320 41514
rect -2325 41486 -2317 41494
rect -2325 41466 -2320 41486
rect -2317 41478 -2309 41486
rect -2325 41450 -2317 41466
rect -2325 41434 -2320 41450
rect -2309 41438 -2301 41450
rect -2317 41434 -2309 41438
rect -2103 41434 -2096 41436
rect -2083 41434 -2053 41436
rect -2325 41422 -2317 41434
rect -2103 41425 -2053 41434
rect -2018 41432 -2017 41438
rect -2003 41432 -2002 41434
rect -2026 41428 -2017 41432
rect -2325 41406 -2320 41422
rect -2309 41410 -2301 41422
rect -2017 41418 -2012 41428
rect -2317 41406 -2309 41410
rect -2325 41394 -2317 41406
rect -2325 41374 -2320 41394
rect -2325 41366 -2317 41374
rect -2325 41346 -2320 41366
rect -2317 41358 -2309 41366
rect -2325 41342 -2317 41346
rect -2000 41342 -1992 41794
rect -1982 41793 -1966 41794
rect -1980 41776 -1932 41783
rect -1655 41776 -1647 41782
rect -1846 41758 -1680 41767
rect -1663 41766 -1655 41776
rect -1671 41726 -1663 41734
rect -1663 41718 -1655 41726
rect -1671 41690 -1663 41706
rect -1655 41678 -1647 41690
rect -1972 41674 -1924 41676
rect -1663 41674 -1655 41678
rect -1972 41665 -1922 41674
rect -1671 41662 -1663 41674
rect -1655 41650 -1647 41662
rect -1663 41646 -1655 41650
rect -1671 41634 -1663 41646
rect -1671 41606 -1663 41614
rect -1663 41598 -1655 41606
rect -1671 41570 -1663 41586
rect -1655 41558 -1647 41570
rect -1972 41554 -1924 41556
rect -1663 41554 -1655 41558
rect -1972 41545 -1922 41554
rect -1671 41542 -1663 41554
rect -1655 41530 -1647 41542
rect -1663 41526 -1655 41530
rect -1671 41514 -1663 41526
rect -1671 41486 -1663 41494
rect -1663 41478 -1655 41486
rect -1671 41450 -1663 41466
rect -1655 41438 -1647 41450
rect -1972 41434 -1924 41436
rect -1663 41434 -1655 41438
rect -1972 41425 -1922 41434
rect -1671 41422 -1663 41434
rect -1655 41410 -1647 41422
rect -1663 41406 -1655 41410
rect -1671 41394 -1663 41406
rect -1671 41366 -1663 41374
rect -1663 41358 -1655 41366
rect -1926 41342 -1892 41345
rect -1671 41342 -1663 41346
rect -1642 41342 -1637 41796
rect -1619 41342 -1614 41796
rect -1530 41342 -1526 41796
rect -1517 41357 -1512 41367
rect -1506 41357 -1502 41796
rect -1507 41343 -1502 41357
rect -1517 41342 -1483 41343
rect -2393 41340 -1483 41342
rect -2371 41294 -2366 41340
rect -2348 41294 -2343 41340
rect -2325 41334 -2317 41340
rect -2053 41338 -1972 41340
rect -2325 41318 -2320 41334
rect -2317 41330 -2309 41334
rect -2069 41330 -2068 41331
rect -2309 41318 -2301 41330
rect -2069 41323 -2038 41330
rect -2069 41321 -2068 41323
rect -2000 41322 -1992 41338
rect -1926 41335 -1924 41340
rect -1916 41332 -1914 41335
rect -1671 41334 -1663 41340
rect -1982 41322 -1916 41331
rect -1663 41330 -1655 41334
rect -2325 41306 -2317 41318
rect -2068 41315 -2053 41321
rect -2027 41320 -1992 41322
rect -2076 41306 -2053 41313
rect -2011 41312 -2002 41320
rect -2000 41312 -1992 41320
rect -1655 41318 -1647 41330
rect -2003 41310 -1992 41312
rect -2325 41294 -2320 41306
rect -2317 41302 -2309 41306
rect -2309 41294 -2301 41302
rect -2015 41298 -2003 41310
rect -2000 41294 -1992 41310
rect -1972 41306 -1924 41313
rect -1862 41305 -1680 41314
rect -1671 41306 -1663 41318
rect -1663 41302 -1655 41306
rect -1976 41294 -1940 41295
rect -1655 41294 -1647 41302
rect -1642 41294 -1637 41340
rect -1619 41294 -1614 41340
rect -1530 41294 -1526 41340
rect -1517 41333 -1512 41340
rect -1507 41319 -1502 41333
rect -1506 41294 -1502 41319
rect -1482 41294 -1478 41796
rect -1458 41294 -1454 41796
rect -1434 41294 -1430 41796
rect -1410 41294 -1406 41796
rect -1397 41381 -1392 41391
rect -1386 41381 -1382 41796
rect -1387 41367 -1382 41381
rect -1386 41294 -1382 41367
rect -1362 41315 -1358 41796
rect -1349 41501 -1344 41511
rect -1338 41501 -1334 41796
rect -1339 41487 -1334 41501
rect -2393 41292 -1365 41294
rect -2371 41222 -2366 41292
rect -2348 41222 -2343 41292
rect -2325 41290 -2320 41292
rect -2309 41290 -2301 41292
rect -2325 41278 -2317 41290
rect -2325 41258 -2320 41278
rect -2317 41274 -2309 41278
rect -2325 41250 -2317 41258
rect -2060 41252 -2030 41255
rect -2325 41222 -2320 41250
rect -2317 41242 -2309 41250
rect -2060 41239 -2038 41250
rect -2033 41243 -2030 41252
rect -2028 41248 -2027 41252
rect -2068 41234 -2038 41237
rect -2000 41222 -1992 41292
rect -1655 41290 -1647 41292
rect -1671 41278 -1663 41290
rect -1663 41274 -1655 41278
rect -1912 41267 -1884 41269
rect -1852 41261 -1804 41265
rect -1844 41252 -1796 41255
rect -1671 41250 -1663 41258
rect -1844 41239 -1804 41250
rect -1663 41242 -1655 41250
rect -1852 41234 -1680 41238
rect -1979 41222 -1945 41224
rect -1642 41222 -1637 41292
rect -1619 41222 -1614 41292
rect -1530 41222 -1526 41292
rect -1506 41222 -1502 41292
rect -1482 41291 -1478 41292
rect -1482 41270 -1475 41291
rect -1458 41270 -1454 41292
rect -1434 41270 -1430 41292
rect -1410 41270 -1406 41292
rect -1386 41270 -1382 41292
rect -1379 41291 -1365 41292
rect -1362 41291 -1355 41315
rect -1362 41270 -1358 41291
rect -1338 41270 -1334 41487
rect -1314 41435 -1310 41796
rect -1314 41411 -1307 41435
rect -1314 41270 -1310 41411
rect -1290 41270 -1286 41796
rect -1277 41789 -1272 41796
rect -1267 41775 -1262 41789
rect -1266 41270 -1262 41775
rect -1242 41747 -1238 41868
rect -1242 41699 -1235 41747
rect -1242 41270 -1238 41699
rect -1218 41270 -1214 41868
rect -1194 41270 -1190 41868
rect -1170 41270 -1166 41868
rect -1157 41741 -1152 41751
rect -1146 41741 -1142 41868
rect -1147 41727 -1142 41741
rect -1146 41270 -1142 41727
rect -1122 41675 -1118 41868
rect -1122 41651 -1115 41675
rect -1122 41270 -1118 41651
rect -1098 41270 -1094 41868
rect -1074 41270 -1070 41868
rect -1050 41463 -1046 41868
rect -1061 41462 -1027 41463
rect -1026 41462 -1022 41868
rect -1002 41462 -998 41868
rect -978 41462 -974 41868
rect -954 41462 -950 41868
rect -947 41867 -933 41868
rect -930 41867 -923 41891
rect -930 41462 -926 41867
rect -906 41462 -902 41892
rect -882 41462 -878 41892
rect -858 41462 -854 41892
rect -845 41621 -840 41631
rect -834 41621 -830 41892
rect -835 41607 -830 41621
rect -834 41462 -830 41607
rect -810 41555 -806 41892
rect -797 41861 -792 41871
rect -786 41861 -782 41892
rect -779 41891 -765 41892
rect -762 41891 -755 41915
rect -787 41847 -782 41861
rect -810 41531 -803 41555
rect -810 41462 -806 41531
rect -786 41462 -782 41847
rect -762 41795 -758 41891
rect -762 41771 -755 41795
rect -762 41462 -758 41771
rect -738 41462 -734 42492
rect -714 41462 -710 42492
rect -690 41462 -686 42492
rect -666 41462 -662 42492
rect -642 41462 -638 42492
rect -618 41583 -614 42492
rect -629 41582 -595 41583
rect -594 41582 -590 42492
rect -570 41582 -566 42492
rect -546 42491 -542 42492
rect -539 42491 -525 42492
rect -522 42491 -515 42515
rect -546 42467 -539 42491
rect -546 41582 -542 42467
rect -522 41582 -518 42491
rect -509 42077 -504 42087
rect -498 42077 -494 42707
rect -499 42063 -494 42077
rect -498 41582 -494 42063
rect -474 42011 -470 42752
rect -474 41987 -467 42011
rect -474 41582 -470 41987
rect -450 41582 -446 42852
rect -426 41582 -422 42852
rect -402 41582 -398 42852
rect -378 42827 -371 42851
rect -378 41582 -374 42827
rect -365 42725 -360 42735
rect -354 42725 -350 42852
rect -355 42711 -350 42725
rect -365 42701 -360 42711
rect -355 42687 -350 42701
rect -354 41582 -350 42687
rect -330 42659 -326 42852
rect -330 42638 -323 42659
rect -306 42638 -302 42852
rect -282 42638 -278 42852
rect -258 42638 -254 42852
rect -234 42638 -230 42852
rect -210 42638 -206 42852
rect -186 42638 -182 42852
rect -162 42638 -158 42852
rect -138 42638 -134 42852
rect -114 42638 -110 42852
rect -90 42638 -86 42852
rect -66 42638 -62 42852
rect -42 42638 -38 42852
rect -18 42638 -14 42852
rect 6 42638 10 42852
rect 30 42851 34 42852
rect 30 42827 37 42851
rect 30 42779 37 42803
rect 30 42638 34 42779
rect 54 42638 58 42852
rect 78 42638 82 42852
rect 102 42638 106 42852
rect 126 42638 130 42852
rect 150 42638 154 42852
rect 174 42638 178 42852
rect 198 42638 202 42852
rect 205 42851 219 42852
rect 222 42851 229 42875
rect 222 42638 226 42851
rect 246 42827 253 42851
rect 246 42638 250 42827
rect 270 42803 277 42827
rect 270 42638 274 42803
rect 283 42725 288 42735
rect 293 42711 298 42725
rect 294 42638 298 42711
rect 307 42638 315 42639
rect -347 42636 315 42638
rect -347 42635 -333 42636
rect -330 42611 -323 42636
rect -330 41582 -326 42611
rect -306 41582 -302 42636
rect -282 41582 -278 42636
rect -258 41582 -254 42636
rect -234 41582 -230 42636
rect -210 41582 -206 42636
rect -197 42413 -192 42423
rect -186 42413 -182 42636
rect -187 42399 -182 42413
rect -186 41582 -182 42399
rect -162 42347 -158 42636
rect -162 42323 -155 42347
rect -162 42159 -158 42323
rect -138 42279 -134 42636
rect -149 42278 -115 42279
rect -114 42278 -110 42636
rect -90 42278 -86 42636
rect -66 42278 -62 42636
rect -42 42278 -38 42636
rect -18 42399 -14 42636
rect -29 42398 5 42399
rect 6 42398 10 42636
rect 30 42398 34 42636
rect 54 42398 58 42636
rect 78 42398 82 42636
rect 102 42398 106 42636
rect 126 42398 130 42636
rect 150 42398 154 42636
rect 174 42398 178 42636
rect 198 42398 202 42636
rect 222 42398 226 42636
rect 246 42398 250 42636
rect 270 42398 274 42636
rect 294 42398 298 42636
rect 301 42635 315 42636
rect 307 42629 312 42635
rect 317 42615 322 42629
rect 318 42398 322 42615
rect 331 42485 336 42495
rect 341 42471 346 42485
rect 342 42398 346 42471
rect 355 42398 363 42399
rect -29 42396 363 42398
rect -29 42389 -24 42396
rect -18 42389 -14 42396
rect -19 42375 -14 42389
rect -29 42365 -24 42375
rect -19 42351 -14 42365
rect -18 42278 -14 42351
rect 6 42323 10 42396
rect -149 42276 3 42278
rect -149 42269 -144 42276
rect -138 42269 -134 42276
rect -139 42255 -134 42269
rect -149 42245 -144 42255
rect -139 42231 -134 42245
rect -173 42158 -139 42159
rect -138 42158 -134 42231
rect -114 42203 -110 42276
rect -173 42156 -117 42158
rect -173 42149 -168 42156
rect -162 42149 -158 42156
rect -163 42135 -158 42149
rect -173 42125 -168 42135
rect -163 42111 -158 42125
rect -162 41582 -158 42111
rect -138 42083 -134 42156
rect -131 42155 -117 42156
rect -114 42155 -107 42203
rect -138 42062 -131 42083
rect -114 42062 -110 42155
rect -90 42062 -86 42276
rect -66 42062 -62 42276
rect -42 42062 -38 42276
rect -18 42062 -14 42276
rect -11 42275 3 42276
rect 6 42275 13 42323
rect 6 42062 10 42275
rect 30 42062 34 42396
rect 43 42197 48 42207
rect 54 42197 58 42396
rect 53 42183 58 42197
rect 54 42062 58 42183
rect 78 42131 82 42396
rect 78 42107 85 42131
rect 78 42062 82 42107
rect 102 42062 106 42396
rect 126 42062 130 42396
rect 150 42062 154 42396
rect 174 42062 178 42396
rect 198 42062 202 42396
rect 222 42062 226 42396
rect 246 42062 250 42396
rect 270 42062 274 42396
rect 294 42062 298 42396
rect 318 42062 322 42396
rect 342 42062 346 42396
rect 349 42395 363 42396
rect 355 42389 360 42395
rect 365 42375 370 42389
rect 366 42062 370 42375
rect 379 42269 384 42279
rect 389 42255 394 42269
rect 390 42062 394 42255
rect 403 42149 408 42159
rect 413 42135 418 42149
rect 414 42062 418 42135
rect 427 42062 435 42063
rect -155 42060 435 42062
rect -155 42059 -141 42060
rect -138 42035 -131 42060
rect -138 41582 -134 42035
rect -114 41582 -110 42060
rect -90 41582 -86 42060
rect -66 41582 -62 42060
rect -53 41885 -48 41895
rect -42 41885 -38 42060
rect -43 41871 -38 41885
rect -42 41582 -38 41871
rect -18 41819 -14 42060
rect -18 41795 -11 41819
rect -18 41582 -14 41795
rect 6 41582 10 42060
rect 30 41582 34 42060
rect 43 41693 48 41703
rect 54 41693 58 42060
rect 53 41679 58 41693
rect 43 41669 48 41679
rect 53 41655 58 41669
rect 54 41582 58 41655
rect 78 41627 82 42060
rect -629 41580 75 41582
rect -629 41573 -624 41580
rect -618 41573 -614 41580
rect -619 41559 -614 41573
rect -629 41549 -624 41559
rect -619 41535 -614 41549
rect -618 41462 -614 41535
rect -594 41507 -590 41580
rect -1061 41460 -597 41462
rect -1061 41453 -1056 41460
rect -1050 41453 -1046 41460
rect -1051 41439 -1046 41453
rect -1061 41429 -1056 41439
rect -1051 41415 -1046 41429
rect -1050 41270 -1046 41415
rect -1026 41387 -1022 41460
rect -1026 41366 -1019 41387
rect -1002 41366 -998 41460
rect -978 41366 -974 41460
rect -954 41366 -950 41460
rect -930 41366 -926 41460
rect -906 41366 -902 41460
rect -882 41366 -878 41460
rect -858 41366 -854 41460
rect -834 41366 -830 41460
rect -810 41366 -806 41460
rect -786 41366 -782 41460
rect -762 41366 -758 41460
rect -738 41366 -734 41460
rect -714 41366 -710 41460
rect -690 41366 -686 41460
rect -666 41366 -662 41460
rect -642 41366 -638 41460
rect -618 41366 -614 41460
rect -611 41459 -597 41460
rect -594 41459 -587 41507
rect -594 41366 -590 41459
rect -570 41366 -566 41580
rect -546 41366 -542 41580
rect -522 41366 -518 41580
rect -498 41366 -494 41580
rect -474 41366 -470 41580
rect -450 41366 -446 41580
rect -426 41366 -422 41580
rect -402 41366 -398 41580
rect -378 41366 -374 41580
rect -354 41366 -350 41580
rect -330 41366 -326 41580
rect -306 41366 -302 41580
rect -282 41366 -278 41580
rect -258 41366 -254 41580
rect -234 41366 -230 41580
rect -210 41366 -206 41580
rect -186 41366 -182 41580
rect -162 41366 -158 41580
rect -138 41366 -134 41580
rect -114 41366 -110 41580
rect -90 41366 -86 41580
rect -66 41366 -62 41580
rect -42 41366 -38 41580
rect -18 41366 -14 41580
rect 6 41366 10 41580
rect 30 41366 34 41580
rect 54 41366 58 41580
rect 61 41579 75 41580
rect 78 41579 85 41627
rect 78 41366 82 41579
rect 102 41366 106 42060
rect 126 41366 130 42060
rect 150 41366 154 42060
rect 174 41366 178 42060
rect 198 41366 202 42060
rect 222 41366 226 42060
rect 246 41366 250 42060
rect 270 41366 274 42060
rect 294 41366 298 42060
rect 318 41366 322 42060
rect 342 41366 346 42060
rect 366 41366 370 42060
rect 390 41366 394 42060
rect 414 41366 418 42060
rect 421 42059 435 42060
rect 427 42053 432 42059
rect 437 42039 442 42053
rect 438 41366 442 42039
rect 451 41933 456 41943
rect 461 41919 466 41933
rect 462 41366 466 41919
rect 475 41813 480 41823
rect 485 41799 490 41813
rect 486 41366 490 41799
rect 499 41693 504 41703
rect 509 41679 514 41693
rect 510 41366 514 41679
rect 523 41573 528 41583
rect 533 41559 538 41573
rect 534 41366 538 41559
rect 547 41453 552 41463
rect 557 41439 562 41453
rect 558 41366 562 41439
rect 571 41366 579 41367
rect -1043 41364 579 41366
rect -1043 41363 -1029 41364
rect -1026 41339 -1019 41364
rect -1026 41270 -1022 41339
rect -1002 41270 -998 41364
rect -978 41270 -974 41364
rect -954 41270 -950 41364
rect -930 41270 -926 41364
rect -906 41270 -902 41364
rect -882 41270 -878 41364
rect -858 41270 -854 41364
rect -834 41270 -830 41364
rect -810 41270 -806 41364
rect -786 41270 -782 41364
rect -762 41270 -758 41364
rect -738 41270 -734 41364
rect -714 41270 -710 41364
rect -690 41270 -686 41364
rect -666 41270 -662 41364
rect -642 41270 -638 41364
rect -618 41270 -614 41364
rect -594 41270 -590 41364
rect -570 41270 -566 41364
rect -546 41270 -542 41364
rect -522 41270 -518 41364
rect -498 41270 -494 41364
rect -474 41270 -470 41364
rect -450 41270 -446 41364
rect -426 41270 -422 41364
rect -402 41270 -398 41364
rect -378 41270 -374 41364
rect -354 41270 -350 41364
rect -341 41309 -336 41319
rect -330 41309 -326 41364
rect -331 41295 -326 41309
rect -330 41270 -326 41295
rect -306 41270 -302 41364
rect -282 41270 -278 41364
rect -258 41270 -254 41364
rect -234 41270 -230 41364
rect -210 41270 -206 41364
rect -186 41270 -182 41364
rect -162 41270 -158 41364
rect -138 41270 -134 41364
rect -114 41271 -110 41364
rect -125 41270 -91 41271
rect -1499 41268 -91 41270
rect -1499 41267 -1485 41268
rect -1482 41243 -1475 41268
rect -1482 41222 -1478 41243
rect -1458 41222 -1454 41268
rect -1434 41222 -1430 41268
rect -1410 41222 -1406 41268
rect -1386 41222 -1382 41268
rect -1362 41222 -1358 41268
rect -1338 41222 -1334 41268
rect -1314 41222 -1310 41268
rect -1290 41222 -1286 41268
rect -1266 41222 -1262 41268
rect -1242 41222 -1238 41268
rect -1218 41222 -1214 41268
rect -1194 41222 -1190 41268
rect -1170 41222 -1166 41268
rect -1146 41222 -1142 41268
rect -1122 41222 -1118 41268
rect -1098 41222 -1094 41268
rect -1074 41222 -1070 41268
rect -1050 41222 -1046 41268
rect -1026 41222 -1022 41268
rect -1002 41222 -998 41268
rect -978 41222 -974 41268
rect -954 41222 -950 41268
rect -930 41222 -926 41268
rect -906 41222 -902 41268
rect -882 41222 -878 41268
rect -858 41222 -854 41268
rect -834 41222 -830 41268
rect -810 41222 -806 41268
rect -786 41222 -782 41268
rect -762 41222 -758 41268
rect -738 41222 -734 41268
rect -725 41237 -720 41247
rect -714 41237 -710 41268
rect -715 41223 -710 41237
rect -725 41222 -691 41223
rect -2393 41220 -691 41222
rect -2371 41174 -2366 41220
rect -2348 41174 -2343 41220
rect -2325 41174 -2320 41220
rect -2309 41202 -2301 41210
rect -2068 41203 -2040 41210
rect -2317 41194 -2309 41202
rect -2000 41193 -1992 41220
rect -1850 41212 -1844 41220
rect -1840 41212 -1792 41220
rect -1894 41210 -1850 41211
rect -1958 41208 -1955 41209
rect -1969 41202 -1955 41208
rect -1894 41203 -1802 41210
rect -1894 41202 -1850 41203
rect -1655 41202 -1647 41210
rect -1969 41200 -1942 41202
rect -1955 41193 -1942 41200
rect -1844 41195 -1802 41201
rect -1663 41194 -1655 41202
rect -1860 41193 -1796 41194
rect -2040 41186 -2020 41193
rect -2004 41186 -1945 41193
rect -1929 41191 -1794 41193
rect -1929 41186 -1850 41191
rect -1844 41186 -1794 41191
rect -2309 41174 -2301 41182
rect -2136 41174 -2129 41184
rect -2068 41176 -2040 41183
rect -2020 41174 -2004 41176
rect -2000 41174 -1992 41186
rect -1844 41185 -1796 41186
rect -1850 41176 -1802 41183
rect -1978 41174 -1942 41175
rect -1655 41174 -1647 41182
rect -1642 41174 -1637 41220
rect -1619 41174 -1614 41220
rect -1530 41174 -1526 41220
rect -1506 41174 -1502 41220
rect -1482 41174 -1478 41220
rect -1458 41174 -1454 41220
rect -1434 41174 -1430 41220
rect -1410 41174 -1406 41220
rect -1386 41174 -1382 41220
rect -1362 41174 -1358 41220
rect -1338 41174 -1334 41220
rect -1314 41174 -1310 41220
rect -1290 41174 -1286 41220
rect -1266 41174 -1262 41220
rect -1242 41174 -1238 41220
rect -1218 41174 -1214 41220
rect -1194 41174 -1190 41220
rect -1170 41174 -1166 41220
rect -1146 41174 -1142 41220
rect -1122 41174 -1118 41220
rect -1098 41174 -1094 41220
rect -1074 41174 -1070 41220
rect -1050 41174 -1046 41220
rect -1026 41174 -1022 41220
rect -1002 41174 -998 41220
rect -978 41174 -974 41220
rect -954 41174 -950 41220
rect -930 41174 -926 41220
rect -906 41174 -902 41220
rect -882 41174 -878 41220
rect -858 41174 -854 41220
rect -834 41174 -830 41220
rect -810 41174 -806 41220
rect -786 41174 -782 41220
rect -762 41174 -758 41220
rect -738 41174 -734 41220
rect -725 41213 -720 41220
rect -715 41199 -710 41213
rect -714 41174 -710 41199
rect -690 41174 -686 41268
rect -666 41174 -662 41268
rect -642 41174 -638 41268
rect -618 41174 -614 41268
rect -594 41174 -590 41268
rect -570 41174 -566 41268
rect -546 41174 -542 41268
rect -522 41174 -518 41268
rect -498 41174 -494 41268
rect -474 41174 -470 41268
rect -450 41174 -446 41268
rect -426 41174 -422 41268
rect -402 41174 -398 41268
rect -378 41174 -374 41268
rect -354 41174 -350 41268
rect -330 41174 -326 41268
rect -306 41243 -302 41268
rect -306 41219 -299 41243
rect -306 41174 -302 41219
rect -282 41174 -278 41268
rect -258 41174 -254 41268
rect -234 41174 -230 41268
rect -210 41174 -206 41268
rect -186 41174 -182 41268
rect -162 41174 -158 41268
rect -138 41174 -134 41268
rect -125 41261 -120 41268
rect -114 41261 -110 41268
rect -115 41247 -110 41261
rect -114 41174 -110 41247
rect -90 41195 -86 41364
rect -2393 41172 -93 41174
rect -2371 41078 -2366 41172
rect -2348 41078 -2343 41172
rect -2325 41134 -2320 41172
rect -2317 41166 -2309 41172
rect -2124 41168 -2117 41172
rect -2060 41168 -2040 41172
rect -2060 41159 -2030 41166
rect -2062 41134 -2032 41135
rect -2000 41134 -1992 41172
rect -1844 41168 -1802 41172
rect -1844 41158 -1792 41167
rect -1663 41166 -1655 41172
rect -1942 41136 -1937 41148
rect -1850 41145 -1822 41146
rect -1850 41141 -1802 41145
rect -2325 41126 -2317 41134
rect -2062 41132 -1961 41134
rect -2325 41106 -2320 41126
rect -2317 41118 -2309 41126
rect -2062 41119 -2040 41130
rect -2032 41125 -1961 41132
rect -1947 41126 -1942 41134
rect -1842 41132 -1794 41135
rect -2070 41114 -2022 41118
rect -2325 41096 -2317 41106
rect -2325 41078 -2320 41096
rect -2317 41090 -2309 41096
rect -2000 41086 -1992 41125
rect -1942 41124 -1937 41126
rect -1932 41116 -1927 41124
rect -1912 41121 -1896 41127
rect -1842 41119 -1802 41130
rect -1671 41126 -1663 41134
rect -1663 41118 -1655 41126
rect -1850 41114 -1680 41118
rect -1937 41100 -1934 41105
rect -1924 41100 -1921 41105
rect -1671 41096 -1663 41106
rect -1842 41092 -1806 41094
rect -1924 41086 -1916 41091
rect -1663 41090 -1655 41096
rect -1854 41086 -1806 41090
rect -2070 41083 -2062 41086
rect -2032 41083 -1960 41086
rect -1944 41083 -1806 41086
rect -2000 41080 -1992 41083
rect -1916 41081 -1914 41083
rect -2033 41078 -1992 41080
rect -1842 41079 -1806 41081
rect -1864 41078 -1796 41079
rect -1642 41078 -1637 41172
rect -1619 41078 -1614 41172
rect -1530 41078 -1526 41172
rect -1506 41078 -1502 41172
rect -1482 41078 -1478 41172
rect -1458 41078 -1454 41172
rect -1434 41078 -1430 41172
rect -1410 41078 -1406 41172
rect -1386 41078 -1382 41172
rect -1362 41078 -1358 41172
rect -1338 41078 -1334 41172
rect -1314 41078 -1310 41172
rect -1290 41078 -1286 41172
rect -1266 41078 -1262 41172
rect -1242 41078 -1238 41172
rect -1218 41078 -1214 41172
rect -1194 41078 -1190 41172
rect -1170 41078 -1166 41172
rect -1146 41078 -1142 41172
rect -1122 41078 -1118 41172
rect -1098 41078 -1094 41172
rect -1074 41078 -1070 41172
rect -1050 41078 -1046 41172
rect -1026 41078 -1022 41172
rect -1002 41078 -998 41172
rect -978 41078 -974 41172
rect -954 41078 -950 41172
rect -930 41078 -926 41172
rect -906 41078 -902 41172
rect -882 41078 -878 41172
rect -858 41078 -854 41172
rect -834 41078 -830 41172
rect -810 41078 -806 41172
rect -786 41078 -782 41172
rect -762 41078 -758 41172
rect -738 41078 -734 41172
rect -714 41078 -710 41172
rect -690 41171 -686 41172
rect -690 41150 -683 41171
rect -666 41150 -662 41172
rect -642 41150 -638 41172
rect -618 41150 -614 41172
rect -594 41150 -590 41172
rect -570 41150 -566 41172
rect -546 41150 -542 41172
rect -522 41150 -518 41172
rect -498 41150 -494 41172
rect -474 41150 -470 41172
rect -450 41150 -446 41172
rect -426 41150 -422 41172
rect -402 41150 -398 41172
rect -378 41150 -374 41172
rect -354 41150 -350 41172
rect -330 41150 -326 41172
rect -306 41150 -302 41172
rect -282 41150 -278 41172
rect -258 41150 -254 41172
rect -234 41150 -230 41172
rect -210 41150 -206 41172
rect -186 41150 -182 41172
rect -162 41150 -158 41172
rect -138 41150 -134 41172
rect -114 41150 -110 41172
rect -107 41171 -93 41172
rect -90 41171 -83 41195
rect -90 41150 -86 41171
rect -66 41150 -62 41364
rect -42 41150 -38 41364
rect -18 41150 -14 41364
rect 6 41150 10 41364
rect 30 41150 34 41364
rect 54 41150 58 41364
rect 78 41150 82 41364
rect 102 41150 106 41364
rect 115 41285 120 41295
rect 126 41285 130 41364
rect 125 41271 130 41285
rect 126 41151 130 41271
rect 150 41219 154 41364
rect 150 41195 157 41219
rect 115 41150 149 41151
rect -707 41148 149 41150
rect -707 41147 -693 41148
rect -690 41123 -683 41148
rect -690 41078 -686 41123
rect -666 41078 -662 41148
rect -642 41078 -638 41148
rect -618 41078 -614 41148
rect -594 41078 -590 41148
rect -570 41079 -566 41148
rect -581 41078 -547 41079
rect -2393 41076 -547 41078
rect -2371 41054 -2366 41076
rect -2348 41054 -2343 41076
rect -2325 41068 -2317 41076
rect -2062 41073 -2032 41076
rect -2000 41073 -1992 41076
rect -1974 41074 -1960 41076
rect -1904 41073 -1798 41076
rect -2080 41069 -2009 41073
rect -2023 41068 -2009 41069
rect -2000 41071 -1798 41073
rect -2000 41069 -1854 41071
rect -1842 41069 -1798 41071
rect -2325 41054 -2320 41068
rect -2317 41062 -2309 41068
rect -2023 41059 -2022 41064
rect -2000 41059 -1992 41069
rect -1671 41068 -1663 41076
rect -1842 41065 -1806 41067
rect -1854 41059 -1806 41063
rect -1663 41062 -1655 41068
rect -2070 41056 -2062 41059
rect -2032 41056 -1904 41059
rect -1888 41056 -1806 41059
rect -2074 41054 -2062 41056
rect -2000 41054 -1992 41056
rect -1642 41054 -1637 41076
rect -1619 41054 -1614 41076
rect -1530 41054 -1526 41076
rect -1506 41054 -1502 41076
rect -1482 41054 -1478 41076
rect -1458 41054 -1454 41076
rect -1434 41054 -1430 41076
rect -1410 41054 -1406 41076
rect -1386 41054 -1382 41076
rect -1362 41054 -1358 41076
rect -1338 41054 -1334 41076
rect -1314 41054 -1310 41076
rect -1290 41054 -1286 41076
rect -1266 41054 -1262 41076
rect -1242 41054 -1238 41076
rect -1218 41054 -1214 41076
rect -1194 41054 -1190 41076
rect -1170 41054 -1166 41076
rect -1146 41054 -1142 41076
rect -1122 41054 -1118 41076
rect -1098 41054 -1094 41076
rect -1074 41054 -1070 41076
rect -1050 41054 -1046 41076
rect -1026 41054 -1022 41076
rect -1002 41054 -998 41076
rect -978 41054 -974 41076
rect -954 41054 -950 41076
rect -930 41054 -926 41076
rect -906 41054 -902 41076
rect -882 41054 -878 41076
rect -858 41054 -854 41076
rect -834 41054 -830 41076
rect -810 41054 -806 41076
rect -786 41054 -782 41076
rect -762 41054 -758 41076
rect -738 41054 -734 41076
rect -714 41054 -710 41076
rect -690 41054 -686 41076
rect -666 41054 -662 41076
rect -642 41054 -638 41076
rect -618 41054 -614 41076
rect -594 41054 -590 41076
rect -581 41069 -576 41076
rect -570 41069 -566 41076
rect -571 41055 -566 41069
rect -570 41054 -566 41055
rect -546 41054 -542 41148
rect -522 41054 -518 41148
rect -498 41054 -494 41148
rect -485 41117 -480 41127
rect -474 41117 -470 41148
rect -475 41103 -470 41117
rect -485 41093 -480 41103
rect -475 41079 -470 41093
rect -474 41054 -470 41079
rect -450 41054 -446 41148
rect -426 41054 -422 41148
rect -402 41054 -398 41148
rect -378 41054 -374 41148
rect -354 41054 -350 41148
rect -330 41054 -326 41148
rect -306 41054 -302 41148
rect -282 41054 -278 41148
rect -258 41054 -254 41148
rect -234 41054 -230 41148
rect -210 41054 -206 41148
rect -186 41054 -182 41148
rect -162 41054 -158 41148
rect -138 41054 -134 41148
rect -114 41054 -110 41148
rect -90 41054 -86 41148
rect -66 41054 -62 41148
rect -42 41054 -38 41148
rect -18 41054 -14 41148
rect 6 41054 10 41148
rect 30 41054 34 41148
rect 54 41054 58 41148
rect 78 41054 82 41148
rect 102 41054 106 41148
rect 115 41141 120 41148
rect 126 41141 130 41148
rect 125 41127 130 41141
rect 126 41054 130 41127
rect 150 41075 154 41195
rect -2393 41052 -2062 41054
rect -2050 41052 147 41054
rect -2371 41006 -2366 41052
rect -2348 41006 -2343 41052
rect -2325 41050 -2320 41052
rect -2325 41040 -2317 41050
rect -2062 41042 -2032 41049
rect -2325 41020 -2320 41040
rect -2317 41034 -2309 41040
rect -2062 41038 -2034 41042
rect -2325 41012 -2317 41020
rect -2101 41015 -2071 41018
rect -2325 41006 -2320 41012
rect -2317 41006 -2309 41012
rect -2000 41010 -1992 41052
rect -1888 41045 -1874 41052
rect -1842 41051 -1806 41052
rect -1842 41042 -1798 41049
rect -1671 41040 -1663 41050
rect -1842 41038 -1806 41040
rect -1663 41034 -1655 41040
rect -1854 41024 -1680 41028
rect -1846 41015 -1798 41018
rect -2079 41009 -2043 41010
rect -2007 41009 -1991 41010
rect -2079 41008 -2071 41009
rect -2079 41006 -2029 41008
rect -2011 41006 -1991 41009
rect -1846 41007 -1806 41013
rect -1671 41012 -1663 41020
rect -1864 41006 -1796 41007
rect -1663 41006 -1655 41012
rect -1642 41006 -1637 41052
rect -1619 41006 -1614 41052
rect -1530 41006 -1526 41052
rect -1506 41006 -1502 41052
rect -1482 41006 -1478 41052
rect -1458 41006 -1454 41052
rect -1434 41006 -1430 41052
rect -1410 41006 -1406 41052
rect -1386 41006 -1382 41052
rect -1362 41006 -1358 41052
rect -1338 41006 -1334 41052
rect -1314 41006 -1310 41052
rect -1290 41006 -1286 41052
rect -1266 41006 -1262 41052
rect -1242 41006 -1238 41052
rect -1218 41006 -1214 41052
rect -1194 41006 -1190 41052
rect -1170 41006 -1166 41052
rect -1146 41006 -1142 41052
rect -1122 41006 -1118 41052
rect -1098 41006 -1094 41052
rect -1074 41006 -1070 41052
rect -1050 41006 -1046 41052
rect -1026 41006 -1022 41052
rect -1002 41006 -998 41052
rect -978 41006 -974 41052
rect -954 41006 -950 41052
rect -930 41006 -926 41052
rect -906 41006 -902 41052
rect -882 41006 -878 41052
rect -858 41006 -854 41052
rect -834 41006 -830 41052
rect -810 41006 -806 41052
rect -786 41006 -782 41052
rect -762 41006 -758 41052
rect -738 41006 -734 41052
rect -714 41006 -710 41052
rect -690 41006 -686 41052
rect -666 41006 -662 41052
rect -642 41006 -638 41052
rect -618 41006 -614 41052
rect -594 41006 -590 41052
rect -570 41006 -566 41052
rect -546 41006 -542 41052
rect -522 41006 -518 41052
rect -498 41006 -494 41052
rect -474 41006 -470 41052
rect -450 41051 -446 41052
rect -450 41030 -443 41051
rect -426 41030 -422 41052
rect -402 41030 -398 41052
rect -378 41030 -374 41052
rect -354 41030 -350 41052
rect -330 41030 -326 41052
rect -306 41030 -302 41052
rect -282 41030 -278 41052
rect -258 41030 -254 41052
rect -234 41030 -230 41052
rect -210 41030 -206 41052
rect -186 41030 -182 41052
rect -162 41030 -158 41052
rect -138 41030 -134 41052
rect -114 41030 -110 41052
rect -90 41030 -86 41052
rect -66 41030 -62 41052
rect -42 41030 -38 41052
rect -18 41030 -14 41052
rect 6 41030 10 41052
rect 30 41030 34 41052
rect 54 41030 58 41052
rect 78 41030 82 41052
rect 102 41030 106 41052
rect 126 41030 130 41052
rect 133 41051 147 41052
rect 150 41051 157 41075
rect 150 41030 154 41051
rect 174 41030 178 41364
rect 198 41030 202 41364
rect 222 41030 226 41364
rect 246 41030 250 41364
rect 270 41030 274 41364
rect 294 41030 298 41364
rect 318 41031 322 41364
rect 307 41030 341 41031
rect -467 41028 341 41030
rect -467 41027 -453 41028
rect -2393 41004 -453 41006
rect -2371 40958 -2366 41004
rect -2348 40958 -2343 41004
rect -2325 40992 -2320 41004
rect -2079 41002 -2071 41004
rect -2072 41000 -2071 41002
rect -2109 40995 -2101 41000
rect -2101 40993 -2079 40995
rect -2069 40993 -2068 41000
rect -2325 40984 -2317 40992
rect -2079 40988 -2071 40993
rect -2325 40964 -2320 40984
rect -2317 40976 -2309 40984
rect -2074 40979 -2071 40988
rect -2069 40984 -2068 40988
rect -2109 40970 -2079 40973
rect -2325 40958 -2317 40964
rect -2000 40958 -1992 41004
rect -1846 41002 -1806 41004
rect -1854 40997 -1806 41001
rect -1854 40995 -1846 40997
rect -1846 40993 -1806 40995
rect -1806 40991 -1798 40993
rect -1846 40988 -1798 40991
rect -1846 40975 -1806 40986
rect -1671 40984 -1663 40992
rect -1663 40976 -1655 40984
rect -1854 40970 -1680 40974
rect -1671 40958 -1663 40964
rect -1642 40958 -1637 41004
rect -1619 40958 -1614 41004
rect -1530 40958 -1526 41004
rect -1506 40958 -1502 41004
rect -1482 40958 -1478 41004
rect -1458 40958 -1454 41004
rect -1434 40958 -1430 41004
rect -1410 40958 -1406 41004
rect -1386 40958 -1382 41004
rect -1362 40958 -1358 41004
rect -1338 40958 -1334 41004
rect -1314 40958 -1310 41004
rect -1290 40958 -1286 41004
rect -1266 40958 -1262 41004
rect -1242 40958 -1238 41004
rect -1218 40958 -1214 41004
rect -1194 40958 -1190 41004
rect -1170 40958 -1166 41004
rect -1146 40958 -1142 41004
rect -1122 40958 -1118 41004
rect -1098 40958 -1094 41004
rect -1074 40958 -1070 41004
rect -1050 40958 -1046 41004
rect -1026 40958 -1022 41004
rect -1002 40958 -998 41004
rect -978 40958 -974 41004
rect -954 40958 -950 41004
rect -930 40958 -926 41004
rect -906 40958 -902 41004
rect -882 40958 -878 41004
rect -858 40958 -854 41004
rect -834 40958 -830 41004
rect -810 40958 -806 41004
rect -786 40958 -782 41004
rect -762 40958 -758 41004
rect -738 40958 -734 41004
rect -714 40958 -710 41004
rect -690 40958 -686 41004
rect -666 40958 -662 41004
rect -642 40958 -638 41004
rect -618 40958 -614 41004
rect -594 40958 -590 41004
rect -570 40958 -566 41004
rect -546 41003 -542 41004
rect -546 40979 -539 41003
rect -546 40958 -542 40979
rect -522 40958 -518 41004
rect -498 40958 -494 41004
rect -474 40958 -470 41004
rect -467 41003 -453 41004
rect -450 41003 -443 41028
rect -450 40958 -446 41003
rect -426 40958 -422 41028
rect -402 40958 -398 41028
rect -378 40958 -374 41028
rect -354 40958 -350 41028
rect -330 40958 -326 41028
rect -306 40958 -302 41028
rect -282 40958 -278 41028
rect -258 40958 -254 41028
rect -234 40958 -230 41028
rect -210 40958 -206 41028
rect -186 40958 -182 41028
rect -162 40958 -158 41028
rect -138 40958 -134 41028
rect -114 40958 -110 41028
rect -90 40958 -86 41028
rect -66 40958 -62 41028
rect -42 40958 -38 41028
rect -18 40958 -14 41028
rect 6 40958 10 41028
rect 30 40958 34 41028
rect 54 40958 58 41028
rect 78 40958 82 41028
rect 102 40958 106 41028
rect 126 40958 130 41028
rect 150 40958 154 41028
rect 174 40958 178 41028
rect 187 40973 192 40983
rect 198 40973 202 41028
rect 197 40959 202 40973
rect 187 40958 221 40959
rect -2393 40956 221 40958
rect -2371 40934 -2366 40956
rect -2348 40934 -2343 40956
rect -2325 40948 -2317 40956
rect -2325 40934 -2320 40948
rect -2309 40936 -2301 40948
rect -2092 40939 -2062 40944
rect -2000 40936 -1992 40956
rect -2317 40934 -2309 40936
rect -2000 40934 -1983 40936
rect -1906 40934 -1904 40956
rect -1806 40948 -1680 40954
rect -1671 40948 -1663 40956
rect -1854 40939 -1806 40944
rect -1846 40934 -1806 40937
rect -1655 40936 -1647 40948
rect -1663 40934 -1655 40936
rect -1642 40934 -1637 40956
rect -1619 40934 -1614 40956
rect -1530 40934 -1526 40956
rect -1506 40934 -1502 40956
rect -1482 40934 -1478 40956
rect -1458 40934 -1454 40956
rect -1434 40934 -1430 40956
rect -1410 40934 -1406 40956
rect -1386 40934 -1382 40956
rect -1362 40934 -1358 40956
rect -1338 40934 -1334 40956
rect -1314 40934 -1310 40956
rect -1290 40934 -1286 40956
rect -1266 40934 -1262 40956
rect -1242 40934 -1238 40956
rect -1218 40934 -1214 40956
rect -1194 40934 -1190 40956
rect -1170 40934 -1166 40956
rect -1146 40934 -1142 40956
rect -1122 40934 -1118 40956
rect -1098 40934 -1094 40956
rect -1074 40934 -1070 40956
rect -1050 40934 -1046 40956
rect -1026 40934 -1022 40956
rect -1002 40934 -998 40956
rect -978 40934 -974 40956
rect -954 40934 -950 40956
rect -930 40934 -926 40956
rect -906 40934 -902 40956
rect -882 40934 -878 40956
rect -858 40934 -854 40956
rect -834 40934 -830 40956
rect -810 40934 -806 40956
rect -786 40934 -782 40956
rect -762 40934 -758 40956
rect -738 40934 -734 40956
rect -714 40934 -710 40956
rect -690 40934 -686 40956
rect -666 40934 -662 40956
rect -642 40934 -638 40956
rect -618 40934 -614 40956
rect -594 40934 -590 40956
rect -570 40934 -566 40956
rect -546 40934 -542 40956
rect -522 40934 -518 40956
rect -498 40934 -494 40956
rect -474 40934 -470 40956
rect -450 40934 -446 40956
rect -426 40934 -422 40956
rect -402 40934 -398 40956
rect -378 40934 -374 40956
rect -354 40934 -350 40956
rect -330 40934 -326 40956
rect -306 40934 -302 40956
rect -282 40934 -278 40956
rect -258 40934 -254 40956
rect -234 40934 -230 40956
rect -210 40934 -206 40956
rect -186 40934 -182 40956
rect -162 40934 -158 40956
rect -138 40934 -134 40956
rect -114 40934 -110 40956
rect -90 40934 -86 40956
rect -66 40934 -62 40956
rect -42 40934 -38 40956
rect -18 40934 -14 40956
rect 6 40934 10 40956
rect 30 40934 34 40956
rect 54 40934 58 40956
rect 78 40934 82 40956
rect 102 40934 106 40956
rect 126 40934 130 40956
rect 150 40934 154 40956
rect 174 40934 178 40956
rect 187 40949 192 40956
rect 197 40935 202 40949
rect 198 40934 202 40935
rect 222 40934 226 41028
rect 246 40934 250 41028
rect 270 40934 274 41028
rect 294 40934 298 41028
rect 307 41021 312 41028
rect 318 41021 322 41028
rect 317 41007 322 41021
rect 318 40934 322 41007
rect 342 40955 346 41364
rect -2393 40932 339 40934
rect -2371 40910 -2366 40932
rect -2348 40910 -2343 40932
rect -2325 40920 -2317 40932
rect -2071 40928 -2062 40932
rect -2013 40930 -1983 40932
rect -2000 40929 -1983 40930
rect -2325 40910 -2320 40920
rect -2309 40910 -2301 40920
rect -2100 40919 -2092 40926
rect -2064 40924 -2062 40927
rect -2061 40919 -2059 40924
rect -2071 40914 -2062 40919
rect -2071 40912 -2026 40914
rect -2066 40910 -2012 40912
rect -2000 40910 -1992 40929
rect -1906 40927 -1904 40932
rect -1846 40928 -1806 40932
rect -1846 40921 -1798 40926
rect -1806 40919 -1798 40921
rect -1671 40920 -1663 40932
rect -1854 40917 -1846 40919
rect -1854 40912 -1806 40917
rect -1864 40910 -1796 40911
rect -1655 40910 -1647 40920
rect -1642 40910 -1637 40932
rect -1619 40910 -1614 40932
rect -1530 40910 -1526 40932
rect -1506 40910 -1502 40932
rect -1482 40910 -1478 40932
rect -1458 40910 -1454 40932
rect -1434 40910 -1430 40932
rect -1410 40910 -1406 40932
rect -1386 40910 -1382 40932
rect -1362 40910 -1358 40932
rect -1338 40910 -1334 40932
rect -1314 40910 -1310 40932
rect -1290 40910 -1286 40932
rect -1266 40910 -1262 40932
rect -1242 40910 -1238 40932
rect -1218 40910 -1214 40932
rect -1194 40910 -1190 40932
rect -1170 40910 -1166 40932
rect -1146 40910 -1142 40932
rect -1122 40910 -1118 40932
rect -1098 40910 -1094 40932
rect -1074 40910 -1070 40932
rect -1050 40910 -1046 40932
rect -1026 40910 -1022 40932
rect -1002 40910 -998 40932
rect -978 40910 -974 40932
rect -954 40910 -950 40932
rect -930 40910 -926 40932
rect -906 40910 -902 40932
rect -882 40910 -878 40932
rect -858 40910 -854 40932
rect -834 40910 -830 40932
rect -810 40910 -806 40932
rect -786 40910 -782 40932
rect -762 40910 -758 40932
rect -738 40910 -734 40932
rect -714 40910 -710 40932
rect -690 40910 -686 40932
rect -666 40910 -662 40932
rect -642 40910 -638 40932
rect -618 40910 -614 40932
rect -594 40910 -590 40932
rect -570 40910 -566 40932
rect -546 40910 -542 40932
rect -522 40910 -518 40932
rect -498 40910 -494 40932
rect -474 40910 -470 40932
rect -450 40910 -446 40932
rect -426 40910 -422 40932
rect -402 40910 -398 40932
rect -378 40910 -374 40932
rect -354 40910 -350 40932
rect -330 40910 -326 40932
rect -306 40910 -302 40932
rect -282 40910 -278 40932
rect -258 40910 -254 40932
rect -234 40910 -230 40932
rect -210 40910 -206 40932
rect -186 40910 -182 40932
rect -162 40910 -158 40932
rect -138 40910 -134 40932
rect -114 40910 -110 40932
rect -90 40910 -86 40932
rect -66 40910 -62 40932
rect -42 40910 -38 40932
rect -18 40910 -14 40932
rect 6 40910 10 40932
rect 30 40910 34 40932
rect 54 40910 58 40932
rect 78 40910 82 40932
rect 102 40910 106 40932
rect 126 40910 130 40932
rect 150 40910 154 40932
rect 174 40910 178 40932
rect 198 40910 202 40932
rect 222 40910 226 40932
rect 246 40910 250 40932
rect 270 40910 274 40932
rect 294 40911 298 40932
rect 283 40910 317 40911
rect -2393 40908 317 40910
rect -2371 40838 -2366 40908
rect -2348 40838 -2343 40908
rect -2325 40904 -2320 40908
rect -2317 40904 -2309 40908
rect -2325 40892 -2317 40904
rect -2066 40903 -2062 40908
rect -2147 40900 -2134 40902
rect -2292 40894 -2071 40900
rect -2325 40838 -2320 40892
rect -2092 40878 -2062 40880
rect -2094 40874 -2062 40878
rect -2309 40844 -2301 40850
rect -2317 40838 -2309 40844
rect -2000 40838 -1992 40908
rect -1846 40901 -1806 40908
rect -1663 40904 -1655 40908
rect -1846 40894 -1680 40900
rect -1671 40892 -1663 40904
rect -1854 40878 -1806 40880
rect -1854 40874 -1680 40878
rect -1655 40844 -1647 40850
rect -1663 40838 -1655 40844
rect -1642 40838 -1637 40908
rect -1619 40838 -1614 40908
rect -1530 40838 -1526 40908
rect -1506 40838 -1502 40908
rect -1482 40838 -1478 40908
rect -1458 40838 -1454 40908
rect -1434 40838 -1430 40908
rect -1410 40838 -1406 40908
rect -1386 40838 -1382 40908
rect -1362 40838 -1358 40908
rect -1338 40838 -1334 40908
rect -1314 40838 -1310 40908
rect -1290 40838 -1286 40908
rect -1266 40838 -1262 40908
rect -1242 40838 -1238 40908
rect -1218 40838 -1214 40908
rect -1194 40838 -1190 40908
rect -1170 40838 -1166 40908
rect -1146 40838 -1142 40908
rect -1122 40838 -1118 40908
rect -1098 40838 -1094 40908
rect -1074 40838 -1070 40908
rect -1050 40838 -1046 40908
rect -1026 40838 -1022 40908
rect -1002 40838 -998 40908
rect -978 40838 -974 40908
rect -954 40838 -950 40908
rect -930 40838 -926 40908
rect -906 40838 -902 40908
rect -882 40838 -878 40908
rect -858 40838 -854 40908
rect -834 40838 -830 40908
rect -810 40838 -806 40908
rect -786 40838 -782 40908
rect -762 40838 -758 40908
rect -738 40838 -734 40908
rect -714 40838 -710 40908
rect -690 40838 -686 40908
rect -666 40838 -662 40908
rect -642 40838 -638 40908
rect -618 40838 -614 40908
rect -594 40838 -590 40908
rect -570 40838 -566 40908
rect -546 40838 -542 40908
rect -522 40838 -518 40908
rect -498 40838 -494 40908
rect -474 40838 -470 40908
rect -450 40863 -446 40908
rect -461 40862 -427 40863
rect -426 40862 -422 40908
rect -402 40862 -398 40908
rect -378 40862 -374 40908
rect -354 40862 -350 40908
rect -330 40862 -326 40908
rect -306 40862 -302 40908
rect -282 40862 -278 40908
rect -258 40862 -254 40908
rect -234 40862 -230 40908
rect -210 40862 -206 40908
rect -186 40862 -182 40908
rect -162 40862 -158 40908
rect -138 40862 -134 40908
rect -114 40862 -110 40908
rect -90 40862 -86 40908
rect -66 40862 -62 40908
rect -42 40862 -38 40908
rect -18 40862 -14 40908
rect 6 40862 10 40908
rect 30 40862 34 40908
rect 54 40862 58 40908
rect 78 40862 82 40908
rect 102 40862 106 40908
rect 126 40862 130 40908
rect 150 40862 154 40908
rect 174 40862 178 40908
rect 198 40862 202 40908
rect 222 40907 226 40908
rect -461 40860 219 40862
rect -461 40853 -456 40860
rect -450 40853 -446 40860
rect -451 40839 -446 40853
rect -461 40838 -427 40839
rect -2393 40836 -427 40838
rect -2371 40742 -2366 40836
rect -2348 40742 -2343 40836
rect -2325 40774 -2320 40836
rect -2317 40834 -2309 40836
rect -2000 40835 -1966 40836
rect -2000 40834 -1982 40835
rect -1663 40834 -1655 40836
rect -2028 40826 -2018 40828
rect -2309 40816 -2301 40822
rect -2091 40816 -2061 40823
rect -2317 40806 -2309 40816
rect -2044 40814 -2028 40816
rect -2026 40814 -2014 40826
rect -2084 40808 -2061 40814
rect -2044 40812 -2014 40814
rect -2292 40798 -2054 40807
rect -2325 40766 -2317 40774
rect -2325 40746 -2320 40766
rect -2317 40758 -2309 40766
rect -2325 40742 -2317 40746
rect -2000 40742 -1992 40834
rect -1982 40833 -1966 40834
rect -1980 40816 -1932 40823
rect -1655 40816 -1647 40822
rect -1846 40798 -1680 40807
rect -1663 40806 -1655 40816
rect -1671 40766 -1663 40774
rect -1663 40758 -1655 40766
rect -1671 40742 -1663 40746
rect -1642 40742 -1637 40836
rect -1619 40742 -1614 40836
rect -1530 40742 -1526 40836
rect -1506 40742 -1502 40836
rect -1482 40742 -1478 40836
rect -1458 40742 -1454 40836
rect -1434 40742 -1430 40836
rect -1410 40742 -1406 40836
rect -1386 40742 -1382 40836
rect -1362 40742 -1358 40836
rect -1338 40742 -1334 40836
rect -1325 40781 -1320 40791
rect -1314 40781 -1310 40836
rect -1315 40767 -1310 40781
rect -1314 40742 -1310 40767
rect -1290 40742 -1286 40836
rect -1266 40742 -1262 40836
rect -1242 40742 -1238 40836
rect -1218 40742 -1214 40836
rect -1194 40742 -1190 40836
rect -1170 40742 -1166 40836
rect -1146 40742 -1142 40836
rect -1122 40742 -1118 40836
rect -1098 40742 -1094 40836
rect -1074 40742 -1070 40836
rect -1050 40742 -1046 40836
rect -1026 40742 -1022 40836
rect -1002 40742 -998 40836
rect -978 40742 -974 40836
rect -954 40742 -950 40836
rect -930 40742 -926 40836
rect -906 40742 -902 40836
rect -882 40742 -878 40836
rect -858 40742 -854 40836
rect -834 40742 -830 40836
rect -810 40742 -806 40836
rect -786 40742 -782 40836
rect -762 40742 -758 40836
rect -738 40742 -734 40836
rect -714 40742 -710 40836
rect -690 40742 -686 40836
rect -666 40742 -662 40836
rect -642 40742 -638 40836
rect -618 40742 -614 40836
rect -605 40757 -600 40767
rect -594 40757 -590 40836
rect -595 40743 -590 40757
rect -605 40742 -571 40743
rect -2393 40740 -1969 40742
rect -1955 40740 -571 40742
rect -2371 40694 -2366 40740
rect -2348 40694 -2343 40740
rect -2325 40730 -2317 40740
rect -2080 40738 -1969 40740
rect -2080 40732 -2053 40738
rect -2325 40714 -2320 40730
rect -2309 40718 -2301 40730
rect -2070 40723 -2040 40730
rect -2000 40722 -1992 40738
rect -1972 40734 -1969 40738
rect -1972 40732 -1955 40734
rect -1955 40722 -1850 40731
rect -1671 40730 -1663 40740
rect -2317 40714 -2309 40718
rect -2070 40715 -2053 40721
rect -2027 40720 -1992 40722
rect -1969 40720 -1955 40721
rect -2325 40702 -2317 40714
rect -2292 40705 -2053 40714
rect -2325 40694 -2320 40702
rect -2309 40694 -2301 40702
rect -2000 40694 -1992 40720
rect -1655 40718 -1647 40730
rect -1663 40714 -1655 40718
rect -1972 40706 -1924 40713
rect -1945 40705 -1929 40706
rect -1860 40705 -1680 40714
rect -1671 40702 -1663 40714
rect -1978 40694 -1942 40695
rect -1655 40694 -1647 40702
rect -1642 40694 -1637 40740
rect -1619 40694 -1614 40740
rect -1530 40694 -1526 40740
rect -1506 40694 -1502 40740
rect -1482 40694 -1478 40740
rect -1458 40694 -1454 40740
rect -1434 40694 -1430 40740
rect -1410 40694 -1406 40740
rect -1386 40694 -1382 40740
rect -1362 40694 -1358 40740
rect -1338 40694 -1334 40740
rect -1314 40694 -1310 40740
rect -1290 40715 -1286 40740
rect -2393 40692 -1293 40694
rect -2371 40598 -2366 40692
rect -2348 40598 -2343 40692
rect -2325 40686 -2320 40692
rect -2309 40690 -2301 40692
rect -2317 40686 -2309 40690
rect -2325 40674 -2317 40686
rect -2325 40654 -2320 40674
rect -2062 40654 -2032 40655
rect -2000 40654 -1992 40692
rect -1655 40690 -1647 40692
rect -1663 40686 -1655 40690
rect -1671 40674 -1663 40686
rect -1942 40656 -1937 40668
rect -1850 40665 -1822 40666
rect -1850 40661 -1802 40665
rect -2325 40646 -2317 40654
rect -2062 40652 -1961 40654
rect -2325 40626 -2320 40646
rect -2317 40638 -2309 40646
rect -2062 40639 -2040 40650
rect -2032 40645 -1961 40652
rect -1947 40646 -1942 40654
rect -1842 40652 -1794 40655
rect -2070 40634 -2022 40638
rect -2325 40614 -2317 40626
rect -2325 40598 -2320 40614
rect -2317 40610 -2309 40614
rect -2309 40598 -2301 40610
rect -2068 40603 -2038 40610
rect -2000 40600 -1992 40645
rect -1942 40644 -1937 40646
rect -1932 40636 -1927 40644
rect -1912 40641 -1896 40647
rect -1842 40639 -1802 40650
rect -1671 40646 -1663 40654
rect -1663 40638 -1655 40646
rect -1850 40634 -1680 40638
rect -1937 40620 -1934 40622
rect -1926 40620 -1921 40625
rect -1926 40615 -1924 40620
rect -1916 40612 -1914 40615
rect -1842 40612 -1794 40621
rect -1671 40614 -1663 40626
rect -1924 40602 -1916 40611
rect -1663 40610 -1655 40614
rect -1852 40603 -1804 40610
rect -1916 40601 -1914 40602
rect -2025 40599 -1991 40600
rect -2025 40598 -1975 40599
rect -1842 40598 -1804 40601
rect -1655 40598 -1647 40610
rect -1642 40598 -1637 40692
rect -1619 40598 -1614 40692
rect -1530 40598 -1526 40692
rect -1506 40598 -1502 40692
rect -1482 40647 -1478 40692
rect -1493 40646 -1459 40647
rect -1458 40646 -1454 40692
rect -1434 40646 -1430 40692
rect -1410 40646 -1406 40692
rect -1386 40646 -1382 40692
rect -1362 40646 -1358 40692
rect -1338 40646 -1334 40692
rect -1314 40646 -1310 40692
rect -1307 40691 -1293 40692
rect -1290 40691 -1283 40715
rect -1290 40646 -1286 40691
rect -1266 40646 -1262 40740
rect -1242 40646 -1238 40740
rect -1218 40646 -1214 40740
rect -1194 40646 -1190 40740
rect -1170 40646 -1166 40740
rect -1146 40646 -1142 40740
rect -1122 40646 -1118 40740
rect -1098 40646 -1094 40740
rect -1074 40646 -1070 40740
rect -1050 40646 -1046 40740
rect -1026 40646 -1022 40740
rect -1002 40646 -998 40740
rect -978 40646 -974 40740
rect -954 40646 -950 40740
rect -930 40646 -926 40740
rect -906 40646 -902 40740
rect -882 40646 -878 40740
rect -858 40646 -854 40740
rect -834 40646 -830 40740
rect -810 40646 -806 40740
rect -786 40646 -782 40740
rect -762 40646 -758 40740
rect -738 40646 -734 40740
rect -714 40646 -710 40740
rect -690 40646 -686 40740
rect -666 40646 -662 40740
rect -642 40646 -638 40740
rect -618 40646 -614 40740
rect -605 40733 -600 40740
rect -595 40719 -590 40733
rect -594 40646 -590 40719
rect -570 40691 -566 40836
rect -570 40670 -563 40691
rect -546 40670 -542 40836
rect -522 40670 -518 40836
rect -498 40670 -494 40836
rect -474 40670 -470 40836
rect -461 40829 -456 40836
rect -451 40815 -446 40829
rect -450 40670 -446 40815
rect -426 40787 -422 40860
rect -426 40766 -419 40787
rect -402 40766 -398 40860
rect -378 40766 -374 40860
rect -354 40766 -350 40860
rect -330 40766 -326 40860
rect -306 40766 -302 40860
rect -282 40766 -278 40860
rect -258 40766 -254 40860
rect -234 40766 -230 40860
rect -210 40766 -206 40860
rect -186 40766 -182 40860
rect -162 40766 -158 40860
rect -138 40766 -134 40860
rect -114 40766 -110 40860
rect -90 40766 -86 40860
rect -66 40766 -62 40860
rect -42 40766 -38 40860
rect -18 40766 -14 40860
rect 6 40766 10 40860
rect 30 40766 34 40860
rect 54 40766 58 40860
rect 78 40766 82 40860
rect 102 40766 106 40860
rect 126 40766 130 40860
rect 150 40766 154 40860
rect 174 40766 178 40860
rect 198 40766 202 40860
rect 205 40859 219 40860
rect 222 40859 229 40907
rect 222 40766 226 40859
rect 246 40766 250 40908
rect 270 40766 274 40908
rect 283 40901 288 40908
rect 294 40901 298 40908
rect 293 40887 298 40901
rect 294 40766 298 40887
rect 318 40835 322 40932
rect 325 40931 339 40932
rect 342 40931 349 40955
rect 318 40811 325 40835
rect 318 40766 322 40811
rect 342 40766 346 40931
rect 366 40766 370 41364
rect 379 40997 384 41007
rect 390 40997 394 41364
rect 389 40983 394 40997
rect 390 40766 394 40983
rect 414 40931 418 41364
rect 414 40907 421 40931
rect 414 40766 418 40907
rect 438 40766 442 41364
rect 462 40766 466 41364
rect 475 41165 480 41175
rect 486 41165 490 41364
rect 485 41151 490 41165
rect 486 40766 490 41151
rect 510 41099 514 41364
rect 510 41075 517 41099
rect 510 40766 514 41075
rect 534 40766 538 41364
rect 558 40766 562 41364
rect 565 41363 579 41364
rect 571 41357 576 41363
rect 581 41343 586 41357
rect 582 40766 586 41343
rect 595 41237 600 41247
rect 605 41223 610 41237
rect 606 40766 610 41223
rect 619 41117 624 41127
rect 629 41103 634 41117
rect 619 41045 624 41055
rect 630 41045 634 41103
rect 629 41031 634 41045
rect 643 41041 651 41045
rect 637 41031 643 41041
rect 630 40766 634 41031
rect 643 40973 648 40983
rect 653 40959 661 40973
rect 654 40955 661 40959
rect 643 40925 648 40935
rect 654 40925 658 40955
rect 653 40911 658 40925
rect 643 40853 648 40863
rect 653 40839 658 40853
rect 667 40849 675 40853
rect 661 40839 667 40849
rect 654 40766 658 40839
rect 667 40766 675 40767
rect -443 40764 675 40766
rect -443 40763 -429 40764
rect -426 40739 -419 40764
rect -426 40670 -422 40739
rect -402 40670 -398 40764
rect -378 40670 -374 40764
rect -354 40670 -350 40764
rect -330 40670 -326 40764
rect -306 40670 -302 40764
rect -282 40670 -278 40764
rect -258 40670 -254 40764
rect -234 40670 -230 40764
rect -210 40670 -206 40764
rect -186 40670 -182 40764
rect -162 40670 -158 40764
rect -138 40670 -134 40764
rect -125 40685 -120 40695
rect -114 40685 -110 40764
rect -115 40671 -110 40685
rect -114 40670 -110 40671
rect -90 40670 -86 40764
rect -66 40670 -62 40764
rect -42 40670 -38 40764
rect -18 40670 -14 40764
rect 6 40670 10 40764
rect 30 40671 34 40764
rect 19 40670 53 40671
rect -587 40668 53 40670
rect -587 40667 -573 40668
rect -1493 40644 -573 40646
rect -1493 40637 -1488 40644
rect -1482 40637 -1478 40644
rect -1483 40623 -1478 40637
rect -1493 40613 -1488 40623
rect -1483 40599 -1478 40613
rect -1482 40598 -1478 40599
rect -1458 40598 -1454 40644
rect -1434 40598 -1430 40644
rect -1410 40598 -1406 40644
rect -1386 40598 -1382 40644
rect -1362 40598 -1358 40644
rect -1338 40598 -1334 40644
rect -1314 40598 -1310 40644
rect -1290 40598 -1286 40644
rect -1266 40598 -1262 40644
rect -1242 40598 -1238 40644
rect -1218 40598 -1214 40644
rect -1194 40598 -1190 40644
rect -1170 40599 -1166 40644
rect -1181 40598 -1147 40599
rect -2393 40596 -1147 40598
rect -2371 40574 -2366 40596
rect -2348 40574 -2343 40596
rect -2325 40586 -2317 40596
rect -2076 40586 -2068 40593
rect -2062 40586 -2001 40593
rect -2325 40574 -2320 40586
rect -2317 40582 -2309 40586
rect -2015 40585 -2001 40586
rect -2309 40574 -2301 40582
rect -2068 40576 -2062 40583
rect -2000 40578 -1992 40596
rect -1974 40594 -1960 40596
rect -1842 40595 -1804 40596
rect -1862 40593 -1794 40594
rect -1985 40591 -1794 40593
rect -1985 40586 -1852 40591
rect -1842 40585 -1794 40591
rect -1671 40586 -1663 40596
rect -2015 40576 -1985 40578
rect -1852 40576 -1804 40583
rect -1663 40582 -1655 40586
rect -2000 40574 -1992 40576
rect -1976 40574 -1940 40575
rect -1655 40574 -1647 40582
rect -1642 40574 -1637 40596
rect -1619 40574 -1614 40596
rect -1530 40574 -1526 40596
rect -1506 40574 -1502 40596
rect -1482 40574 -1478 40596
rect -1458 40574 -1454 40596
rect -1434 40574 -1430 40596
rect -1410 40574 -1406 40596
rect -1386 40574 -1382 40596
rect -1362 40574 -1358 40596
rect -1338 40574 -1334 40596
rect -1314 40574 -1310 40596
rect -1290 40574 -1286 40596
rect -1266 40574 -1262 40596
rect -1242 40574 -1238 40596
rect -1218 40574 -1214 40596
rect -1194 40574 -1190 40596
rect -1181 40589 -1176 40596
rect -1170 40589 -1166 40596
rect -1171 40575 -1166 40589
rect -1170 40574 -1166 40575
rect -1146 40574 -1142 40644
rect -1122 40574 -1118 40644
rect -1098 40574 -1094 40644
rect -1074 40574 -1070 40644
rect -1050 40574 -1046 40644
rect -1026 40574 -1022 40644
rect -1002 40574 -998 40644
rect -978 40574 -974 40644
rect -954 40574 -950 40644
rect -930 40574 -926 40644
rect -906 40574 -902 40644
rect -882 40574 -878 40644
rect -858 40574 -854 40644
rect -834 40574 -830 40644
rect -810 40574 -806 40644
rect -786 40574 -782 40644
rect -762 40574 -758 40644
rect -738 40574 -734 40644
rect -714 40574 -710 40644
rect -690 40574 -686 40644
rect -666 40574 -662 40644
rect -642 40574 -638 40644
rect -618 40574 -614 40644
rect -594 40574 -590 40644
rect -587 40643 -573 40644
rect -570 40643 -563 40668
rect -570 40574 -566 40643
rect -546 40574 -542 40668
rect -522 40574 -518 40668
rect -498 40574 -494 40668
rect -474 40574 -470 40668
rect -450 40574 -446 40668
rect -426 40574 -422 40668
rect -402 40574 -398 40668
rect -378 40574 -374 40668
rect -354 40574 -350 40668
rect -330 40574 -326 40668
rect -306 40574 -302 40668
rect -282 40574 -278 40668
rect -258 40574 -254 40668
rect -234 40574 -230 40668
rect -210 40574 -206 40668
rect -186 40574 -182 40668
rect -162 40574 -158 40668
rect -138 40574 -134 40668
rect -114 40574 -110 40668
rect -90 40619 -86 40668
rect -90 40595 -83 40619
rect -90 40574 -86 40595
rect -66 40574 -62 40668
rect -42 40574 -38 40668
rect -18 40574 -14 40668
rect 6 40574 10 40668
rect 19 40661 24 40668
rect 30 40661 34 40668
rect 29 40647 34 40661
rect 30 40574 34 40647
rect 54 40595 58 40764
rect -2393 40572 51 40574
rect -2371 40502 -2366 40572
rect -2348 40502 -2343 40572
rect -2325 40570 -2320 40572
rect -2309 40570 -2301 40572
rect -2325 40558 -2317 40570
rect -2062 40559 -2032 40566
rect -2325 40538 -2320 40558
rect -2317 40554 -2309 40558
rect -2325 40530 -2317 40538
rect -2060 40532 -2030 40535
rect -2325 40502 -2320 40530
rect -2317 40522 -2309 40530
rect -2060 40519 -2038 40530
rect -2033 40523 -2030 40532
rect -2028 40528 -2027 40532
rect -2068 40514 -2038 40517
rect -2000 40502 -1992 40572
rect -1888 40567 -1874 40572
rect -1842 40568 -1804 40572
rect -1655 40570 -1647 40572
rect -1902 40565 -1874 40567
rect -1842 40558 -1794 40567
rect -1671 40558 -1663 40570
rect -1663 40554 -1655 40558
rect -1912 40547 -1884 40549
rect -1852 40541 -1804 40545
rect -1844 40532 -1796 40535
rect -1671 40530 -1663 40538
rect -1844 40519 -1804 40530
rect -1663 40522 -1655 40530
rect -1852 40514 -1680 40518
rect -1642 40502 -1637 40572
rect -1619 40502 -1614 40572
rect -1530 40502 -1526 40572
rect -1506 40502 -1502 40572
rect -1482 40502 -1478 40572
rect -1458 40571 -1454 40572
rect -1458 40550 -1451 40571
rect -1434 40550 -1430 40572
rect -1410 40550 -1406 40572
rect -1386 40550 -1382 40572
rect -1362 40550 -1358 40572
rect -1338 40550 -1334 40572
rect -1314 40550 -1310 40572
rect -1290 40550 -1286 40572
rect -1266 40550 -1262 40572
rect -1242 40550 -1238 40572
rect -1218 40550 -1214 40572
rect -1194 40550 -1190 40572
rect -1170 40550 -1166 40572
rect -1146 40550 -1142 40572
rect -1122 40550 -1118 40572
rect -1098 40550 -1094 40572
rect -1074 40550 -1070 40572
rect -1050 40550 -1046 40572
rect -1026 40550 -1022 40572
rect -1002 40550 -998 40572
rect -978 40550 -974 40572
rect -954 40550 -950 40572
rect -930 40550 -926 40572
rect -906 40550 -902 40572
rect -882 40550 -878 40572
rect -858 40550 -854 40572
rect -834 40550 -830 40572
rect -810 40550 -806 40572
rect -786 40550 -782 40572
rect -762 40550 -758 40572
rect -738 40550 -734 40572
rect -714 40550 -710 40572
rect -690 40550 -686 40572
rect -666 40550 -662 40572
rect -642 40550 -638 40572
rect -618 40550 -614 40572
rect -594 40550 -590 40572
rect -570 40550 -566 40572
rect -546 40550 -542 40572
rect -522 40550 -518 40572
rect -498 40550 -494 40572
rect -474 40550 -470 40572
rect -450 40550 -446 40572
rect -426 40550 -422 40572
rect -402 40550 -398 40572
rect -378 40550 -374 40572
rect -354 40550 -350 40572
rect -330 40550 -326 40572
rect -306 40550 -302 40572
rect -282 40550 -278 40572
rect -258 40550 -254 40572
rect -234 40550 -230 40572
rect -210 40550 -206 40572
rect -186 40550 -182 40572
rect -162 40550 -158 40572
rect -138 40550 -134 40572
rect -114 40551 -110 40572
rect -125 40550 -91 40551
rect -1475 40548 -91 40550
rect -1475 40547 -1461 40548
rect -1458 40523 -1451 40548
rect -1458 40502 -1454 40523
rect -1434 40502 -1430 40548
rect -1410 40502 -1406 40548
rect -1386 40502 -1382 40548
rect -1362 40502 -1358 40548
rect -1338 40502 -1334 40548
rect -1314 40502 -1310 40548
rect -1290 40502 -1286 40548
rect -1266 40502 -1262 40548
rect -1242 40502 -1238 40548
rect -1218 40502 -1214 40548
rect -1194 40502 -1190 40548
rect -1170 40502 -1166 40548
rect -1146 40523 -1142 40548
rect -2393 40500 -1149 40502
rect -2371 40478 -2366 40500
rect -2348 40478 -2343 40500
rect -2325 40478 -2320 40500
rect -2309 40482 -2301 40492
rect -2068 40483 -2062 40488
rect -2317 40478 -2309 40482
rect -2060 40478 -2050 40483
rect -2000 40478 -1992 40500
rect -1806 40492 -1680 40498
rect -1854 40483 -1806 40488
rect -1655 40482 -1647 40492
rect -1972 40478 -1964 40479
rect -1958 40478 -1942 40480
rect -1844 40478 -1806 40481
rect -1663 40478 -1655 40482
rect -1642 40478 -1637 40500
rect -1619 40478 -1614 40500
rect -1530 40478 -1526 40500
rect -1506 40478 -1502 40500
rect -1482 40478 -1478 40500
rect -1458 40478 -1454 40500
rect -1434 40478 -1430 40500
rect -1410 40478 -1406 40500
rect -1386 40478 -1382 40500
rect -1362 40478 -1358 40500
rect -1338 40478 -1334 40500
rect -1314 40478 -1310 40500
rect -1290 40478 -1286 40500
rect -1266 40478 -1262 40500
rect -1242 40478 -1238 40500
rect -1218 40478 -1214 40500
rect -1194 40478 -1190 40500
rect -1170 40478 -1166 40500
rect -1163 40499 -1149 40500
rect -1146 40499 -1139 40523
rect -1146 40478 -1142 40499
rect -1122 40478 -1118 40548
rect -1098 40478 -1094 40548
rect -1074 40478 -1070 40548
rect -1050 40478 -1046 40548
rect -1026 40478 -1022 40548
rect -1002 40478 -998 40548
rect -978 40478 -974 40548
rect -954 40478 -950 40548
rect -930 40478 -926 40548
rect -906 40478 -902 40548
rect -882 40478 -878 40548
rect -858 40478 -854 40548
rect -834 40478 -830 40548
rect -810 40478 -806 40548
rect -786 40478 -782 40548
rect -762 40478 -758 40548
rect -738 40478 -734 40548
rect -714 40478 -710 40548
rect -690 40478 -686 40548
rect -666 40478 -662 40548
rect -642 40478 -638 40548
rect -618 40478 -614 40548
rect -594 40478 -590 40548
rect -570 40478 -566 40548
rect -546 40478 -542 40548
rect -522 40478 -518 40548
rect -498 40478 -494 40548
rect -474 40478 -470 40548
rect -450 40478 -446 40548
rect -426 40478 -422 40548
rect -402 40478 -398 40548
rect -378 40478 -374 40548
rect -354 40478 -350 40548
rect -330 40478 -326 40548
rect -306 40478 -302 40548
rect -282 40478 -278 40548
rect -258 40478 -254 40548
rect -234 40478 -230 40548
rect -210 40478 -206 40548
rect -186 40478 -182 40548
rect -162 40478 -158 40548
rect -138 40478 -134 40548
rect -125 40541 -120 40548
rect -114 40541 -110 40548
rect -115 40527 -110 40541
rect -114 40478 -110 40527
rect -90 40478 -86 40572
rect -66 40478 -62 40572
rect -42 40478 -38 40572
rect -18 40478 -14 40572
rect 6 40478 10 40572
rect 30 40478 34 40572
rect 37 40571 51 40572
rect 54 40571 61 40595
rect 54 40478 58 40571
rect 78 40478 82 40764
rect 102 40478 106 40764
rect 115 40565 120 40575
rect 126 40565 130 40764
rect 125 40551 130 40565
rect 126 40478 130 40551
rect 150 40499 154 40764
rect -2393 40476 147 40478
rect -2371 40454 -2366 40476
rect -2348 40454 -2343 40476
rect -2325 40454 -2320 40476
rect -2060 40470 -2050 40476
rect -2309 40454 -2301 40464
rect -2060 40463 -2030 40470
rect -2000 40466 -1992 40476
rect -1972 40474 -1942 40476
rect -1958 40473 -1942 40474
rect -1844 40472 -1806 40476
rect -2068 40456 -2062 40463
rect -2062 40454 -2036 40456
rect -2393 40452 -2036 40454
rect -2030 40454 -2012 40456
rect -2004 40454 -1990 40466
rect -1844 40465 -1798 40470
rect -1806 40463 -1798 40465
rect -1854 40461 -1844 40463
rect -1854 40456 -1806 40461
rect -1864 40454 -1796 40455
rect -1655 40454 -1647 40464
rect -1642 40454 -1637 40476
rect -1619 40454 -1614 40476
rect -1530 40454 -1526 40476
rect -1506 40454 -1502 40476
rect -1482 40454 -1478 40476
rect -1458 40454 -1454 40476
rect -1434 40454 -1430 40476
rect -1410 40454 -1406 40476
rect -1386 40454 -1382 40476
rect -1362 40454 -1358 40476
rect -1338 40454 -1334 40476
rect -1314 40454 -1310 40476
rect -1290 40454 -1286 40476
rect -1266 40454 -1262 40476
rect -1242 40454 -1238 40476
rect -1218 40454 -1214 40476
rect -1194 40454 -1190 40476
rect -1170 40454 -1166 40476
rect -1146 40454 -1142 40476
rect -1122 40454 -1118 40476
rect -1098 40454 -1094 40476
rect -1074 40454 -1070 40476
rect -1050 40454 -1046 40476
rect -1026 40454 -1022 40476
rect -1002 40454 -998 40476
rect -978 40454 -974 40476
rect -954 40454 -950 40476
rect -930 40454 -926 40476
rect -906 40454 -902 40476
rect -882 40454 -878 40476
rect -858 40454 -854 40476
rect -834 40454 -830 40476
rect -810 40454 -806 40476
rect -786 40454 -782 40476
rect -762 40454 -758 40476
rect -738 40454 -734 40476
rect -714 40454 -710 40476
rect -690 40454 -686 40476
rect -666 40454 -662 40476
rect -642 40454 -638 40476
rect -618 40454 -614 40476
rect -594 40454 -590 40476
rect -570 40454 -566 40476
rect -546 40454 -542 40476
rect -522 40454 -518 40476
rect -498 40454 -494 40476
rect -474 40454 -470 40476
rect -450 40454 -446 40476
rect -426 40454 -422 40476
rect -402 40454 -398 40476
rect -378 40454 -374 40476
rect -354 40454 -350 40476
rect -330 40454 -326 40476
rect -306 40454 -302 40476
rect -282 40454 -278 40476
rect -258 40454 -254 40476
rect -234 40454 -230 40476
rect -210 40454 -206 40476
rect -186 40454 -182 40476
rect -162 40454 -158 40476
rect -138 40454 -134 40476
rect -114 40454 -110 40476
rect -90 40475 -86 40476
rect -2030 40452 -93 40454
rect -2371 40406 -2366 40452
rect -2348 40406 -2343 40452
rect -2325 40406 -2320 40452
rect -2317 40448 -2309 40452
rect -2060 40448 -2050 40452
rect -2060 40446 -2036 40448
rect -2060 40444 -2030 40446
rect -2292 40438 -2030 40444
rect -2092 40422 -2062 40424
rect -2094 40418 -2062 40422
rect -2000 40406 -1992 40452
rect -1844 40445 -1806 40452
rect -1663 40448 -1655 40452
rect -1844 40438 -1680 40444
rect -1854 40422 -1806 40424
rect -1854 40418 -1680 40422
rect -1642 40406 -1637 40452
rect -1619 40406 -1614 40452
rect -1530 40406 -1526 40452
rect -1506 40406 -1502 40452
rect -1482 40406 -1478 40452
rect -1458 40406 -1454 40452
rect -1434 40406 -1430 40452
rect -1410 40406 -1406 40452
rect -1386 40406 -1382 40452
rect -1362 40406 -1358 40452
rect -1338 40406 -1334 40452
rect -1314 40406 -1310 40452
rect -1290 40406 -1286 40452
rect -1266 40406 -1262 40452
rect -1242 40406 -1238 40452
rect -1218 40406 -1214 40452
rect -1194 40406 -1190 40452
rect -1170 40406 -1166 40452
rect -1146 40406 -1142 40452
rect -1122 40406 -1118 40452
rect -1098 40406 -1094 40452
rect -1074 40406 -1070 40452
rect -1050 40406 -1046 40452
rect -1026 40406 -1022 40452
rect -1002 40406 -998 40452
rect -978 40406 -974 40452
rect -954 40406 -950 40452
rect -930 40406 -926 40452
rect -906 40406 -902 40452
rect -882 40406 -878 40452
rect -858 40406 -854 40452
rect -834 40406 -830 40452
rect -810 40406 -806 40452
rect -786 40406 -782 40452
rect -762 40406 -758 40452
rect -738 40406 -734 40452
rect -714 40406 -710 40452
rect -690 40406 -686 40452
rect -666 40406 -662 40452
rect -642 40406 -638 40452
rect -618 40406 -614 40452
rect -594 40406 -590 40452
rect -570 40406 -566 40452
rect -546 40406 -542 40452
rect -522 40406 -518 40452
rect -498 40406 -494 40452
rect -474 40406 -470 40452
rect -450 40406 -446 40452
rect -426 40406 -422 40452
rect -402 40406 -398 40452
rect -378 40406 -374 40452
rect -354 40406 -350 40452
rect -330 40406 -326 40452
rect -306 40406 -302 40452
rect -282 40406 -278 40452
rect -258 40406 -254 40452
rect -234 40406 -230 40452
rect -210 40406 -206 40452
rect -186 40406 -182 40452
rect -162 40406 -158 40452
rect -138 40406 -134 40452
rect -114 40406 -110 40452
rect -107 40451 -93 40452
rect -90 40451 -83 40475
rect -90 40406 -86 40451
rect -66 40406 -62 40476
rect -42 40406 -38 40476
rect -18 40406 -14 40476
rect 6 40406 10 40476
rect 19 40445 24 40455
rect 30 40445 34 40476
rect 29 40431 34 40445
rect 30 40406 34 40431
rect 54 40406 58 40476
rect 78 40406 82 40476
rect 102 40406 106 40476
rect 126 40406 130 40476
rect 133 40475 147 40476
rect 150 40475 157 40499
rect 150 40406 154 40475
rect 174 40406 178 40764
rect 198 40406 202 40764
rect 222 40406 226 40764
rect 235 40517 240 40527
rect 246 40517 250 40764
rect 245 40503 250 40517
rect 235 40493 240 40503
rect 245 40479 250 40493
rect 246 40406 250 40479
rect 270 40451 274 40764
rect -2393 40404 267 40406
rect -2371 40382 -2366 40404
rect -2348 40382 -2343 40404
rect -2325 40382 -2320 40404
rect -2072 40402 -2036 40403
rect -2072 40396 -2054 40402
rect -2309 40388 -2301 40396
rect -2317 40382 -2309 40388
rect -2092 40387 -2062 40392
rect -2000 40383 -1992 40404
rect -1938 40403 -1906 40404
rect -1920 40402 -1906 40403
rect -1806 40396 -1680 40402
rect -1854 40387 -1806 40392
rect -1655 40388 -1647 40396
rect -1982 40383 -1966 40384
rect -2000 40382 -1966 40383
rect -1846 40382 -1806 40385
rect -1663 40382 -1655 40388
rect -1642 40382 -1637 40404
rect -1619 40382 -1614 40404
rect -1530 40382 -1526 40404
rect -1506 40382 -1502 40404
rect -1482 40382 -1478 40404
rect -1458 40382 -1454 40404
rect -1434 40382 -1430 40404
rect -1410 40382 -1406 40404
rect -1386 40382 -1382 40404
rect -1362 40382 -1358 40404
rect -1338 40382 -1334 40404
rect -1314 40382 -1310 40404
rect -1290 40382 -1286 40404
rect -1266 40382 -1262 40404
rect -1242 40382 -1238 40404
rect -1218 40382 -1214 40404
rect -1194 40382 -1190 40404
rect -1170 40382 -1166 40404
rect -1146 40382 -1142 40404
rect -1122 40382 -1118 40404
rect -1098 40382 -1094 40404
rect -1074 40382 -1070 40404
rect -1050 40382 -1046 40404
rect -1026 40382 -1022 40404
rect -1002 40382 -998 40404
rect -978 40382 -974 40404
rect -954 40382 -950 40404
rect -930 40382 -926 40404
rect -906 40382 -902 40404
rect -882 40382 -878 40404
rect -858 40382 -854 40404
rect -834 40382 -830 40404
rect -810 40382 -806 40404
rect -786 40382 -782 40404
rect -762 40382 -758 40404
rect -738 40383 -734 40404
rect -749 40382 -715 40383
rect -2393 40380 -715 40382
rect -2371 40358 -2366 40380
rect -2348 40358 -2343 40380
rect -2325 40358 -2320 40380
rect -2000 40378 -1966 40380
rect -2309 40360 -2301 40368
rect -2062 40367 -2054 40374
rect -2092 40360 -2084 40367
rect -2062 40360 -2026 40362
rect -2317 40358 -2309 40360
rect -2062 40358 -2012 40360
rect -2000 40358 -1992 40378
rect -1982 40377 -1966 40378
rect -1846 40376 -1806 40380
rect -1846 40369 -1798 40374
rect -1806 40367 -1798 40369
rect -1854 40365 -1846 40367
rect -1854 40360 -1806 40365
rect -1655 40360 -1647 40368
rect -1864 40358 -1796 40359
rect -1663 40358 -1655 40360
rect -1642 40358 -1637 40380
rect -1619 40358 -1614 40380
rect -1530 40358 -1526 40380
rect -1506 40358 -1502 40380
rect -1482 40358 -1478 40380
rect -1458 40358 -1454 40380
rect -1434 40358 -1430 40380
rect -1410 40358 -1406 40380
rect -1386 40358 -1382 40380
rect -1362 40358 -1358 40380
rect -1338 40358 -1334 40380
rect -1314 40358 -1310 40380
rect -1290 40358 -1286 40380
rect -1266 40358 -1262 40380
rect -1242 40358 -1238 40380
rect -1218 40358 -1214 40380
rect -1194 40358 -1190 40380
rect -1170 40358 -1166 40380
rect -1146 40358 -1142 40380
rect -1122 40359 -1118 40380
rect -1133 40358 -1099 40359
rect -2393 40356 -1099 40358
rect -2371 40310 -2366 40356
rect -2348 40310 -2343 40356
rect -2325 40310 -2320 40356
rect -2317 40352 -2309 40356
rect -2062 40352 -2054 40356
rect -2154 40348 -2138 40350
rect -2057 40348 -2054 40352
rect -2292 40342 -2054 40348
rect -2052 40342 -2044 40352
rect -2092 40326 -2062 40328
rect -2094 40322 -2062 40326
rect -2000 40310 -1992 40356
rect -1846 40349 -1806 40356
rect -1663 40352 -1655 40356
rect -1846 40342 -1680 40348
rect -1854 40326 -1806 40328
rect -1854 40322 -1680 40326
rect -1642 40310 -1637 40356
rect -1619 40310 -1614 40356
rect -1530 40310 -1526 40356
rect -1506 40310 -1502 40356
rect -1482 40310 -1478 40356
rect -1458 40310 -1454 40356
rect -1434 40310 -1430 40356
rect -1410 40310 -1406 40356
rect -1386 40310 -1382 40356
rect -1362 40310 -1358 40356
rect -1338 40310 -1334 40356
rect -1314 40310 -1310 40356
rect -1290 40310 -1286 40356
rect -1266 40310 -1262 40356
rect -1242 40310 -1238 40356
rect -1218 40310 -1214 40356
rect -1194 40310 -1190 40356
rect -1170 40310 -1166 40356
rect -1146 40310 -1142 40356
rect -1133 40349 -1128 40356
rect -1122 40349 -1118 40356
rect -1123 40335 -1118 40349
rect -1122 40310 -1118 40335
rect -1098 40310 -1094 40380
rect -1074 40310 -1070 40380
rect -1050 40310 -1046 40380
rect -1026 40310 -1022 40380
rect -1002 40310 -998 40380
rect -978 40310 -974 40380
rect -954 40310 -950 40380
rect -930 40310 -926 40380
rect -906 40310 -902 40380
rect -882 40310 -878 40380
rect -858 40310 -854 40380
rect -834 40310 -830 40380
rect -810 40310 -806 40380
rect -786 40310 -782 40380
rect -762 40310 -758 40380
rect -749 40373 -744 40380
rect -738 40373 -734 40380
rect -739 40359 -734 40373
rect -738 40310 -734 40359
rect -714 40310 -710 40404
rect -690 40310 -686 40404
rect -666 40310 -662 40404
rect -642 40310 -638 40404
rect -618 40310 -614 40404
rect -594 40310 -590 40404
rect -570 40310 -566 40404
rect -546 40310 -542 40404
rect -522 40310 -518 40404
rect -498 40310 -494 40404
rect -474 40310 -470 40404
rect -450 40310 -446 40404
rect -426 40310 -422 40404
rect -402 40310 -398 40404
rect -378 40310 -374 40404
rect -354 40310 -350 40404
rect -330 40310 -326 40404
rect -317 40325 -312 40335
rect -306 40325 -302 40404
rect -307 40311 -302 40325
rect -317 40310 -283 40311
rect -2393 40308 -283 40310
rect -2371 40286 -2366 40308
rect -2348 40286 -2343 40308
rect -2325 40286 -2320 40308
rect -2072 40306 -2036 40307
rect -2072 40300 -2054 40306
rect -2309 40292 -2301 40300
rect -2317 40286 -2309 40292
rect -2092 40291 -2062 40296
rect -2000 40287 -1992 40308
rect -1938 40307 -1906 40308
rect -1920 40306 -1906 40307
rect -1806 40300 -1680 40306
rect -1854 40291 -1806 40296
rect -1655 40292 -1647 40300
rect -1982 40287 -1966 40288
rect -2000 40286 -1966 40287
rect -1846 40286 -1806 40289
rect -1663 40286 -1655 40292
rect -1642 40286 -1637 40308
rect -1619 40286 -1614 40308
rect -1530 40286 -1526 40308
rect -1506 40286 -1502 40308
rect -1482 40286 -1478 40308
rect -1458 40286 -1454 40308
rect -1434 40286 -1430 40308
rect -1410 40286 -1406 40308
rect -1386 40286 -1382 40308
rect -1362 40286 -1358 40308
rect -1338 40286 -1334 40308
rect -1314 40286 -1310 40308
rect -1290 40286 -1286 40308
rect -1266 40286 -1262 40308
rect -1242 40286 -1238 40308
rect -1218 40286 -1214 40308
rect -1194 40286 -1190 40308
rect -1170 40286 -1166 40308
rect -1146 40286 -1142 40308
rect -1122 40286 -1118 40308
rect -1098 40286 -1094 40308
rect -1074 40286 -1070 40308
rect -1050 40286 -1046 40308
rect -1026 40286 -1022 40308
rect -1002 40286 -998 40308
rect -978 40286 -974 40308
rect -954 40286 -950 40308
rect -930 40286 -926 40308
rect -906 40286 -902 40308
rect -882 40286 -878 40308
rect -858 40286 -854 40308
rect -834 40286 -830 40308
rect -810 40286 -806 40308
rect -786 40286 -782 40308
rect -762 40286 -758 40308
rect -738 40286 -734 40308
rect -714 40307 -710 40308
rect -2393 40284 -717 40286
rect -2371 40262 -2366 40284
rect -2348 40262 -2343 40284
rect -2325 40262 -2320 40284
rect -2000 40282 -1966 40284
rect -2309 40264 -2301 40272
rect -2062 40271 -2054 40278
rect -2092 40264 -2084 40271
rect -2062 40264 -2026 40266
rect -2317 40262 -2309 40264
rect -2062 40262 -2012 40264
rect -2000 40262 -1992 40282
rect -1982 40281 -1966 40282
rect -1846 40280 -1806 40284
rect -1846 40273 -1798 40278
rect -1806 40271 -1798 40273
rect -1854 40269 -1846 40271
rect -1854 40264 -1806 40269
rect -1655 40264 -1647 40272
rect -1864 40262 -1796 40263
rect -1663 40262 -1655 40264
rect -1642 40262 -1637 40284
rect -1619 40262 -1614 40284
rect -1530 40262 -1526 40284
rect -1506 40262 -1502 40284
rect -1482 40262 -1478 40284
rect -1458 40262 -1454 40284
rect -1434 40262 -1430 40284
rect -1410 40262 -1406 40284
rect -1386 40263 -1382 40284
rect -1397 40262 -1363 40263
rect -2393 40260 -1363 40262
rect -2371 39843 -2366 40260
rect -2361 39863 -2353 39873
rect -2348 39863 -2343 40260
rect -2351 39847 -2343 39863
rect -2371 39817 -2363 39843
rect -2383 39645 -2376 39655
rect -2371 39645 -2366 39817
rect -2373 39634 -2366 39645
rect -2348 39634 -2343 39847
rect -2325 40129 -2320 40260
rect -2317 40256 -2309 40260
rect -2062 40256 -2054 40260
rect -2154 40252 -2138 40254
rect -2057 40252 -2054 40256
rect -2292 40246 -2054 40252
rect -2052 40246 -2044 40256
rect -2092 40230 -2062 40232
rect -2094 40226 -2062 40230
rect -2309 40196 -2301 40205
rect -2317 40189 -2309 40196
rect -2309 40168 -2301 40176
rect -2251 40170 -2093 40176
rect -2317 40160 -2309 40168
rect -2154 40163 -2138 40166
rect -2084 40163 -2054 40168
rect -2143 40150 -2138 40156
rect -2325 40119 -2317 40129
rect -2325 40100 -2320 40119
rect -2317 40113 -2309 40119
rect -2243 40102 -2221 40110
rect -2211 40102 -2201 40122
rect -2073 40102 -2065 40120
rect -2000 40102 -1992 40260
rect -1846 40253 -1806 40260
rect -1663 40256 -1655 40260
rect -1846 40246 -1680 40252
rect -1854 40230 -1806 40232
rect -1854 40226 -1680 40230
rect -1915 40196 -1906 40206
rect -1846 40204 -1837 40206
rect -1790 40204 -1680 40206
rect -1655 40196 -1647 40202
rect -1905 40187 -1896 40196
rect -1837 40195 -1790 40196
rect -1837 40180 -1798 40193
rect -1663 40186 -1655 40196
rect -1798 40170 -1790 40175
rect -1837 40168 -1798 40170
rect -1655 40168 -1647 40174
rect -1846 40166 -1837 40168
rect -1846 40163 -1798 40166
rect -1837 40150 -1798 40160
rect -1663 40158 -1655 40168
rect -1671 40118 -1663 40126
rect -1655 40118 -1647 40120
rect -1663 40110 -1647 40118
rect -1642 40110 -1637 40260
rect -1885 40102 -1877 40104
rect -1708 40102 -1672 40104
rect -2243 40101 -2213 40102
rect -2325 40091 -2317 40100
rect -2259 40095 -2211 40101
rect -2183 40095 -1877 40102
rect -1869 40095 -1758 40102
rect -1710 40096 -1672 40102
rect -1710 40095 -1692 40096
rect -2211 40091 -2201 40095
rect -2325 40071 -2320 40091
rect -2317 40084 -2309 40091
rect -2211 40084 -2198 40091
rect -2325 40063 -2317 40071
rect -2300 40064 -2292 40074
rect -2243 40065 -2228 40076
rect -2211 40068 -2181 40084
rect -2211 40065 -2201 40068
rect -2325 40043 -2320 40063
rect -2317 40055 -2309 40063
rect -2325 40035 -2317 40043
rect -2325 40015 -2320 40035
rect -2317 40027 -2309 40035
rect -2325 40006 -2317 40015
rect -2325 39987 -2320 40006
rect -2317 39999 -2309 40006
rect -2325 39978 -2317 39987
rect -2325 39958 -2320 39978
rect -2317 39971 -2309 39978
rect -2325 39950 -2317 39958
rect -2290 39951 -2282 40064
rect -2251 40054 -2240 40058
rect -2211 40054 -2181 40058
rect -2251 40051 -2181 40054
rect -2176 40044 -2173 40046
rect -2240 40037 -2173 40044
rect -2169 40039 -2163 40094
rect -2073 40058 -2065 40095
rect -2073 40054 -2043 40058
rect -2000 40054 -1992 40095
rect -1915 40064 -1907 40073
rect -1963 40058 -1955 40064
rect -1963 40054 -1915 40058
rect -1885 40054 -1877 40095
rect -1875 40090 -1869 40094
rect -1829 40072 -1781 40074
rect -1847 40068 -1781 40072
rect -1778 40068 -1771 40094
rect -1758 40087 -1710 40094
rect -1718 40080 -1710 40087
rect -1768 40070 -1760 40080
rect -1718 40078 -1700 40080
rect -2146 40051 -2135 40054
rect -2105 40051 -2043 40054
rect -2035 40051 -1989 40054
rect -1973 40051 -1915 40054
rect -1907 40051 -1854 40054
rect -2073 40049 -2043 40051
rect -2135 40037 -2105 40044
rect -2065 40042 -2043 40049
rect -2243 40026 -2240 40035
rect -2221 40029 -2213 40037
rect -2211 40029 -2208 40037
rect -2203 40030 -2173 40037
rect -2251 40019 -2240 40026
rect -2211 40026 -2203 40029
rect -2211 40019 -2181 40026
rect -2073 40019 -2043 40026
rect -2203 39996 -2173 40003
rect -2262 39978 -2240 39988
rect -2203 39987 -2176 39996
rect -2083 39985 -2075 39995
rect -2040 39985 -2035 39989
rect -2073 39973 -2043 39985
rect -2028 39973 -2023 39985
rect -2000 39978 -1992 40051
rect -1963 40048 -1955 40051
rect -1963 40047 -1915 40048
rect -1955 40037 -1907 40044
rect -1885 40040 -1877 40051
rect -1837 40046 -1828 40062
rect -1758 40055 -1750 40070
rect -1758 40054 -1692 40055
rect -1837 40044 -1833 40046
rect -1837 40042 -1835 40044
rect -1887 40037 -1851 40040
rect -1750 40037 -1702 40044
rect -1885 40032 -1877 40037
rect -1963 40019 -1915 40026
rect -1905 39987 -1897 40032
rect -1857 40014 -1851 40037
rect -1760 40029 -1758 40030
rect -1837 40019 -1789 40026
rect -1758 40020 -1750 40026
rect -1758 40019 -1710 40020
rect -1955 39984 -1915 39987
rect -1963 39978 -1962 39980
rect -2000 39975 -1981 39978
rect -1965 39975 -1962 39978
rect -1955 39978 -1907 39982
rect -1885 39978 -1877 39997
rect -1857 39984 -1851 39996
rect -1750 39992 -1702 39999
rect -1829 39984 -1789 39986
rect -1766 39982 -1760 39992
rect -1829 39978 -1781 39982
rect -1756 39978 -1740 39982
rect -1680 39978 -1672 40096
rect -1671 40090 -1663 40098
rect -1645 40094 -1637 40110
rect -1663 40082 -1655 40090
rect -1671 40062 -1663 40070
rect -1663 40054 -1655 40062
rect -1671 40034 -1663 40042
rect -1671 40018 -1669 40031
rect -1663 40026 -1655 40034
rect -1671 40006 -1663 40014
rect -1663 39998 -1655 40006
rect -1671 39978 -1663 39986
rect -1955 39975 -1837 39978
rect -1829 39975 -1740 39978
rect -2206 39965 -2176 39968
rect -2206 39962 -2203 39965
rect -2161 39963 -2145 39972
rect -2073 39970 -2065 39973
rect -2073 39969 -2043 39970
rect -2028 39969 -2012 39973
rect -2073 39962 -2065 39968
rect -2203 39961 -2176 39962
rect -2065 39961 -2043 39962
rect -2262 39955 -2232 39961
rect -2176 39955 -2173 39961
rect -2043 39955 -2035 39961
rect -2325 39930 -2320 39950
rect -2317 39942 -2309 39950
rect -2153 39949 -2146 39953
rect -2325 39922 -2317 39930
rect -2300 39926 -2292 39936
rect -2325 39902 -2320 39922
rect -2317 39914 -2309 39922
rect -2325 39894 -2317 39902
rect -2325 39874 -2320 39894
rect -2317 39886 -2309 39894
rect -2290 39893 -2282 39926
rect -2273 39922 -2264 39927
rect -2206 39922 -2176 39927
rect -2262 39915 -2232 39920
rect -2198 39911 -2176 39922
rect -2198 39897 -2176 39905
rect -2166 39889 -2158 39937
rect -2143 39933 -2136 39949
rect -2143 39922 -2113 39927
rect -2073 39922 -2065 39927
rect -2065 39920 -2043 39922
rect -2043 39915 -2035 39920
rect -2065 39894 -2043 39909
rect -2006 39893 -2004 39909
rect -2265 39879 -2260 39885
rect -2143 39879 -2113 39886
rect -2270 39878 -2240 39879
rect -2270 39875 -2265 39878
rect -2325 39866 -2317 39874
rect -2325 39846 -2320 39866
rect -2317 39858 -2309 39866
rect -2113 39863 -2105 39873
rect -2291 39851 -2270 39858
rect -2198 39856 -2168 39858
rect -2135 39857 -2105 39858
rect -2103 39857 -2095 39863
rect -2113 39856 -2105 39857
rect -2065 39856 -2035 39858
rect -2000 39856 -1992 39975
rect -1963 39968 -1960 39975
rect -1915 39971 -1905 39975
rect -1963 39967 -1955 39968
rect -1963 39961 -1915 39967
rect -1989 39934 -1973 39937
rect -1915 39934 -1907 39941
rect -1990 39899 -1989 39920
rect -1983 39856 -1981 39919
rect -1885 39910 -1877 39975
rect -1789 39970 -1778 39975
rect -1837 39967 -1829 39968
rect -1837 39961 -1789 39967
rect -1756 39966 -1740 39975
rect -1837 39951 -1829 39961
rect -1872 39932 -1867 39942
rect -1789 39934 -1781 39941
rect -1776 39934 -1769 39951
rect -1756 39944 -1750 39966
rect -1671 39962 -1669 39973
rect -1663 39970 -1655 39978
rect -1671 39950 -1663 39958
rect -1663 39942 -1655 39950
rect -1702 39932 -1696 39938
rect -1955 39908 -1915 39910
rect -1963 39906 -1955 39908
rect -1963 39899 -1915 39906
rect -1963 39891 -1955 39899
rect -1963 39890 -1915 39891
rect -1973 39884 -1965 39887
rect -1955 39884 -1907 39888
rect -1974 39881 -1907 39884
rect -1973 39877 -1965 39881
rect -1963 39877 -1960 39879
rect -1963 39873 -1915 39877
rect -1963 39865 -1955 39873
rect -1963 39861 -1915 39865
rect -1963 39858 -1955 39861
rect -2240 39851 -2206 39856
rect -2198 39851 -2143 39856
rect -2113 39851 -1981 39856
rect -1915 39851 -1907 39858
rect -2270 39846 -2266 39850
rect -2086 39847 -2070 39851
rect -2325 39838 -2317 39846
rect -2270 39839 -2240 39846
rect -2206 39839 -2176 39846
rect -2325 39818 -2320 39838
rect -2317 39830 -2309 39838
rect -2270 39834 -2266 39839
rect -2270 39830 -2266 39833
rect -2198 39830 -2176 39837
rect -2166 39830 -2158 39847
rect -2143 39839 -2113 39846
rect -2198 39821 -2168 39825
rect -2325 39810 -2317 39818
rect -2143 39816 -2136 39830
rect -2085 39825 -2060 39826
rect -2039 39825 -2035 39834
rect -2135 39818 -2105 39825
rect -2085 39818 -2035 39825
rect -2029 39818 -2025 39825
rect -2325 39797 -2320 39810
rect -2317 39802 -2309 39810
rect -2235 39800 -2232 39803
rect -2325 39771 -2317 39797
rect -2325 39762 -2320 39771
rect -2325 39754 -2317 39762
rect -2135 39754 -2119 39767
rect -2000 39759 -1992 39851
rect -1983 39833 -1981 39851
rect -1955 39833 -1915 39834
rect -1862 39830 -1857 39932
rect -1706 39928 -1702 39932
rect -1829 39916 -1789 39924
rect -1671 39922 -1663 39930
rect -1849 39908 -1842 39916
rect -1790 39908 -1781 39916
rect -1663 39914 -1655 39922
rect -1837 39899 -1829 39906
rect -1758 39899 -1732 39906
rect -1748 39890 -1732 39899
rect -1671 39894 -1663 39902
rect -1829 39881 -1781 39888
rect -1663 39886 -1655 39894
rect -1829 39875 -1789 39879
rect -1768 39876 -1760 39886
rect -1758 39875 -1750 39876
rect -1671 39866 -1663 39874
rect -1837 39863 -1780 39866
rect -1758 39860 -1748 39866
rect -1708 39860 -1690 39866
rect -1829 39851 -1781 39858
rect -1680 39849 -1672 39866
rect -1663 39858 -1655 39866
rect -1829 39840 -1791 39846
rect -1758 39840 -1710 39842
rect -1758 39833 -1692 39840
rect -1671 39838 -1663 39846
rect -1955 39822 -1907 39825
rect -1791 39822 -1781 39825
rect -1991 39818 -1839 39822
rect -1791 39818 -1780 39822
rect -1680 39815 -1672 39833
rect -1663 39830 -1655 39838
rect -1839 39805 -1791 39812
rect -1671 39810 -1663 39818
rect -1829 39799 -1791 39803
rect -1671 39800 -1669 39810
rect -1663 39802 -1655 39810
rect -1680 39784 -1672 39799
rect -1642 39784 -1637 40094
rect -1619 40044 -1614 40260
rect -1619 40018 -1611 40044
rect -1768 39768 -1760 39778
rect -1758 39761 -1710 39768
rect -2325 39734 -2320 39754
rect -2317 39746 -2306 39754
rect -2031 39751 -1992 39759
rect -1750 39757 -1710 39761
rect -1674 39756 -1663 39762
rect -2307 39738 -2306 39746
rect -2149 39749 -2135 39750
rect -2149 39745 -2119 39749
rect -2024 39740 -2021 39749
rect -2325 39726 -2317 39734
rect -2325 39678 -2320 39726
rect -2317 39718 -2306 39726
rect -2185 39724 -2169 39736
rect -2056 39733 -2040 39737
rect -2021 39733 -2008 39740
rect -2056 39722 -2054 39732
rect -2056 39721 -2048 39722
rect -2307 39682 -2306 39690
rect -2111 39689 -2054 39695
rect -2325 39670 -2314 39678
rect -2104 39671 -2101 39675
rect -2325 39650 -2320 39670
rect -2314 39662 -2306 39670
rect -2104 39668 -2101 39670
rect -2084 39668 -2054 39669
rect -2000 39668 -1992 39751
rect -1758 39750 -1750 39751
rect -1758 39749 -1749 39750
rect -1758 39748 -1710 39749
rect -1663 39746 -1658 39756
rect -1831 39738 -1783 39742
rect -1784 39725 -1783 39738
rect -1674 39728 -1663 39734
rect -1826 39723 -1796 39724
rect -1663 39718 -1658 39728
rect -1654 39724 -1647 39734
rect -1644 39710 -1637 39724
rect -1758 39692 -1750 39695
rect -1758 39689 -1710 39692
rect -1844 39677 -1828 39679
rect -1844 39676 -1792 39677
rect -1828 39675 -1792 39676
rect -1772 39675 -1758 39683
rect -1750 39680 -1702 39687
rect -1750 39672 -1710 39676
rect -1700 39672 -1692 39692
rect -1674 39684 -1665 39692
rect -1674 39672 -1666 39680
rect -1758 39668 -1710 39669
rect -2307 39654 -2306 39662
rect -2139 39658 -2123 39667
rect -2111 39662 -2016 39668
rect -2139 39651 -2111 39658
rect -2325 39642 -2314 39650
rect -2177 39644 -2161 39645
rect -2141 39644 -2119 39646
rect -2104 39644 -2101 39662
rect -2076 39651 -2046 39656
rect -2325 39634 -2320 39642
rect -2314 39634 -2306 39642
rect -2076 39640 -2054 39646
rect -2021 39643 -2016 39662
rect -2000 39662 -1818 39668
rect -1802 39662 -1776 39668
rect -1760 39662 -1710 39668
rect -1666 39664 -1658 39672
rect -2189 39634 -2175 39639
rect -2373 39632 -2175 39634
rect -2373 39631 -2359 39632
rect -2371 39494 -2366 39631
rect -2348 39579 -2343 39632
rect -2325 39622 -2320 39632
rect -2307 39626 -2306 39632
rect -2189 39631 -2175 39632
rect -2149 39630 -2119 39639
rect -2084 39638 -2036 39639
rect -2000 39638 -1992 39662
rect -1758 39660 -1710 39662
rect -1758 39658 -1755 39660
rect -1828 39651 -1792 39658
rect -1768 39649 -1760 39656
rect -1758 39651 -1757 39658
rect -1710 39657 -1702 39658
rect -1750 39651 -1702 39657
rect -1674 39656 -1665 39664
rect -1768 39646 -1764 39649
rect -1758 39646 -1755 39651
rect -1818 39638 -1789 39646
rect -1758 39639 -1754 39646
rect -1750 39641 -1710 39646
rect -1674 39644 -1666 39652
rect -1758 39638 -1692 39639
rect -2084 39636 -1692 39638
rect -1666 39636 -1658 39644
rect -2084 39633 -1690 39636
rect -2084 39630 -2054 39633
rect -2046 39631 -1710 39633
rect -2325 39614 -2314 39622
rect -2076 39621 -2046 39628
rect -2325 39594 -2320 39614
rect -2314 39606 -2306 39614
rect -2076 39613 -2054 39619
rect -2084 39609 -2054 39611
rect -2104 39606 -2054 39609
rect -2307 39598 -2306 39606
rect -2084 39603 -2054 39606
rect -2325 39580 -2314 39594
rect -2348 39555 -2341 39579
rect -2325 39564 -2320 39580
rect -2314 39578 -2309 39580
rect -2309 39566 -2298 39578
rect -2092 39575 -2060 39576
rect -2062 39570 -2060 39575
rect -2314 39564 -2309 39566
rect -2348 39494 -2343 39555
rect -2325 39552 -2314 39564
rect -2076 39560 -2062 39570
rect -2076 39554 -2046 39558
rect -2014 39557 -2003 39566
rect -2062 39552 -2046 39554
rect -2325 39536 -2320 39552
rect -2314 39550 -2309 39552
rect -2076 39551 -2062 39552
rect -2309 39538 -2298 39550
rect -2092 39545 -2076 39551
rect -2046 39545 -2026 39546
rect -2314 39536 -2309 39538
rect -2046 39536 -2042 39537
rect -2325 39524 -2314 39536
rect -2141 39532 -2134 39534
rect -2052 39532 -2046 39536
rect -2292 39527 -2111 39532
rect -2096 39530 -2046 39532
rect -2076 39527 -2046 39530
rect -2325 39494 -2320 39524
rect -2314 39522 -2309 39524
rect -2092 39510 -2062 39512
rect -2094 39506 -2062 39510
rect -2000 39494 -1992 39631
rect -1758 39630 -1710 39631
rect -1680 39628 -1665 39636
rect -1750 39621 -1702 39628
rect -1680 39624 -1672 39628
rect -1680 39619 -1666 39624
rect -1836 39615 -1820 39616
rect -1837 39611 -1820 39615
rect -1750 39613 -1710 39619
rect -1674 39616 -1666 39619
rect -1837 39604 -1789 39611
rect -1758 39610 -1710 39611
rect -1760 39607 -1692 39610
rect -1666 39608 -1658 39616
rect -1837 39603 -1820 39604
rect -1764 39603 -1692 39607
rect -1674 39603 -1665 39608
rect -1680 39600 -1665 39603
rect -1750 39584 -1702 39586
rect -1680 39576 -1672 39600
rect -1671 39580 -1666 39596
rect -1854 39575 -1806 39576
rect -1829 39560 -1806 39570
rect -1655 39568 -1650 39580
rect -1666 39564 -1655 39568
rect -1829 39554 -1798 39558
rect -1680 39557 -1672 39560
rect -1806 39552 -1798 39554
rect -1671 39552 -1666 39564
rect -1829 39551 -1806 39552
rect -1854 39549 -1829 39551
rect -1854 39545 -1806 39549
rect -1829 39533 -1806 39543
rect -1655 39540 -1650 39552
rect -1666 39536 -1655 39540
rect -1829 39527 -1680 39532
rect -1671 39524 -1666 39536
rect -1854 39510 -1806 39512
rect -1854 39506 -1680 39510
rect -1642 39494 -1637 39710
rect -1619 39708 -1614 40018
rect -1619 39634 -1612 39658
rect -1619 39494 -1614 39634
rect -1530 39494 -1526 40260
rect -1506 39494 -1502 40260
rect -1482 39494 -1478 40260
rect -1458 39494 -1454 40260
rect -1434 39494 -1430 40260
rect -1410 39494 -1406 40260
rect -1397 40253 -1392 40260
rect -1386 40253 -1382 40260
rect -1387 40239 -1382 40253
rect -1386 39494 -1382 40239
rect -1362 40187 -1358 40284
rect -1362 40163 -1355 40187
rect -1362 39494 -1358 40163
rect -1338 39494 -1334 40284
rect -1314 39494 -1310 40284
rect -1301 39533 -1296 39543
rect -1290 39533 -1286 40284
rect -1291 39519 -1286 39533
rect -1290 39494 -1286 39519
rect -1266 39494 -1262 40284
rect -1242 39494 -1238 40284
rect -1218 39494 -1214 40284
rect -1194 39494 -1190 40284
rect -1181 39509 -1176 39519
rect -1170 39509 -1166 40284
rect -1171 39495 -1166 39509
rect -1181 39494 -1147 39495
rect -2393 39492 -1147 39494
rect -2371 39470 -2366 39492
rect -2348 39470 -2343 39492
rect -2325 39470 -2320 39492
rect -2072 39490 -2036 39491
rect -2072 39484 -2054 39490
rect -2309 39476 -2301 39484
rect -2317 39470 -2309 39476
rect -2092 39475 -2062 39480
rect -2000 39471 -1992 39492
rect -1938 39491 -1906 39492
rect -1920 39490 -1906 39491
rect -1806 39484 -1680 39490
rect -1854 39475 -1806 39480
rect -1655 39476 -1647 39484
rect -1982 39471 -1966 39472
rect -2000 39470 -1966 39471
rect -1846 39470 -1806 39473
rect -1663 39470 -1655 39476
rect -1642 39470 -1637 39492
rect -1619 39470 -1614 39492
rect -1530 39470 -1526 39492
rect -1506 39470 -1502 39492
rect -1482 39470 -1478 39492
rect -1458 39470 -1454 39492
rect -1434 39470 -1430 39492
rect -1410 39470 -1406 39492
rect -1386 39470 -1382 39492
rect -1362 39470 -1358 39492
rect -1338 39470 -1334 39492
rect -1314 39470 -1310 39492
rect -1290 39470 -1286 39492
rect -1266 39470 -1262 39492
rect -1242 39470 -1238 39492
rect -1218 39470 -1214 39492
rect -1194 39470 -1190 39492
rect -1181 39485 -1176 39492
rect -1171 39471 -1166 39485
rect -1170 39470 -1166 39471
rect -1146 39470 -1142 40284
rect -1122 39470 -1118 40284
rect -1098 40283 -1094 40284
rect -1098 40259 -1091 40283
rect -1098 39470 -1094 40259
rect -1074 39470 -1070 40284
rect -1050 39470 -1046 40284
rect -1026 39470 -1022 40284
rect -1002 39470 -998 40284
rect -989 40085 -984 40095
rect -978 40085 -974 40284
rect -979 40071 -974 40085
rect -989 40061 -984 40071
rect -979 40047 -974 40061
rect -978 39470 -974 40047
rect -954 40019 -950 40284
rect -954 39971 -947 40019
rect -954 39470 -950 39971
rect -930 39470 -926 40284
rect -906 39471 -902 40284
rect -917 39470 -883 39471
rect -2393 39468 -883 39470
rect -2371 39446 -2366 39468
rect -2348 39446 -2343 39468
rect -2325 39446 -2320 39468
rect -2000 39466 -1966 39468
rect -2309 39448 -2301 39456
rect -2062 39455 -2054 39462
rect -2092 39448 -2084 39455
rect -2062 39448 -2026 39450
rect -2317 39446 -2309 39448
rect -2062 39446 -2012 39448
rect -2000 39446 -1992 39466
rect -1982 39465 -1966 39466
rect -1846 39464 -1806 39468
rect -1846 39457 -1798 39462
rect -1806 39455 -1798 39457
rect -1854 39453 -1846 39455
rect -1854 39448 -1806 39453
rect -1655 39448 -1647 39456
rect -1864 39446 -1796 39447
rect -1663 39446 -1655 39448
rect -1642 39446 -1637 39468
rect -1619 39446 -1614 39468
rect -1530 39446 -1526 39468
rect -1506 39446 -1502 39468
rect -1482 39446 -1478 39468
rect -1458 39446 -1454 39468
rect -1434 39446 -1430 39468
rect -1410 39446 -1406 39468
rect -1386 39446 -1382 39468
rect -1362 39446 -1358 39468
rect -1338 39446 -1334 39468
rect -1314 39446 -1310 39468
rect -1290 39446 -1286 39468
rect -1266 39467 -1262 39468
rect -2393 39444 -1269 39446
rect -2371 39398 -2366 39444
rect -2348 39398 -2343 39444
rect -2325 39398 -2320 39444
rect -2317 39440 -2309 39444
rect -2062 39440 -2054 39444
rect -2154 39436 -2138 39438
rect -2057 39436 -2054 39440
rect -2292 39430 -2054 39436
rect -2052 39430 -2044 39440
rect -2092 39414 -2062 39416
rect -2094 39410 -2062 39414
rect -2000 39398 -1992 39444
rect -1846 39437 -1806 39444
rect -1663 39440 -1655 39444
rect -1846 39430 -1680 39436
rect -1854 39414 -1806 39416
rect -1854 39410 -1680 39414
rect -1642 39398 -1637 39444
rect -1619 39398 -1614 39444
rect -1530 39398 -1526 39444
rect -1506 39398 -1502 39444
rect -1482 39398 -1478 39444
rect -1458 39398 -1454 39444
rect -1434 39398 -1430 39444
rect -1410 39398 -1406 39444
rect -1386 39398 -1382 39444
rect -1362 39398 -1358 39444
rect -1338 39398 -1334 39444
rect -1314 39398 -1310 39444
rect -1290 39398 -1286 39444
rect -1283 39443 -1269 39444
rect -1266 39443 -1259 39467
rect -1266 39398 -1262 39443
rect -1242 39398 -1238 39468
rect -1218 39398 -1214 39468
rect -1194 39398 -1190 39468
rect -1170 39398 -1166 39468
rect -1146 39443 -1142 39468
rect -2393 39396 -1149 39398
rect -2371 39374 -2366 39396
rect -2348 39374 -2343 39396
rect -2325 39374 -2320 39396
rect -2072 39394 -2036 39395
rect -2072 39388 -2054 39394
rect -2309 39380 -2301 39388
rect -2317 39374 -2309 39380
rect -2092 39379 -2062 39384
rect -2000 39375 -1992 39396
rect -1938 39395 -1906 39396
rect -1920 39394 -1906 39395
rect -1806 39388 -1680 39394
rect -1854 39379 -1806 39384
rect -1655 39380 -1647 39388
rect -1982 39375 -1966 39376
rect -2000 39374 -1966 39375
rect -1846 39374 -1806 39377
rect -1663 39374 -1655 39380
rect -1642 39374 -1637 39396
rect -1619 39374 -1614 39396
rect -1530 39374 -1526 39396
rect -1506 39374 -1502 39396
rect -1482 39374 -1478 39396
rect -1458 39374 -1454 39396
rect -1434 39374 -1430 39396
rect -1410 39374 -1406 39396
rect -1386 39374 -1382 39396
rect -1362 39374 -1358 39396
rect -1338 39374 -1334 39396
rect -1314 39374 -1310 39396
rect -1290 39374 -1286 39396
rect -1266 39374 -1262 39396
rect -1242 39374 -1238 39396
rect -1218 39374 -1214 39396
rect -1194 39374 -1190 39396
rect -1170 39374 -1166 39396
rect -1163 39395 -1149 39396
rect -1146 39395 -1139 39443
rect -1146 39374 -1142 39395
rect -1122 39374 -1118 39468
rect -1098 39374 -1094 39468
rect -1074 39374 -1070 39468
rect -1050 39374 -1046 39468
rect -1026 39374 -1022 39468
rect -1002 39374 -998 39468
rect -978 39374 -974 39468
rect -954 39374 -950 39468
rect -930 39374 -926 39468
rect -917 39461 -912 39468
rect -906 39461 -902 39468
rect -907 39447 -902 39461
rect -906 39374 -902 39447
rect -882 39395 -878 40284
rect -2393 39372 -885 39374
rect -2371 39350 -2366 39372
rect -2348 39350 -2343 39372
rect -2325 39350 -2320 39372
rect -2000 39370 -1966 39372
rect -2309 39352 -2301 39360
rect -2062 39359 -2054 39366
rect -2092 39352 -2084 39359
rect -2062 39352 -2026 39354
rect -2317 39350 -2309 39352
rect -2062 39350 -2012 39352
rect -2000 39350 -1992 39370
rect -1982 39369 -1966 39370
rect -1846 39368 -1806 39372
rect -1846 39361 -1798 39366
rect -1806 39359 -1798 39361
rect -1854 39357 -1846 39359
rect -1854 39352 -1806 39357
rect -1655 39352 -1647 39360
rect -1864 39350 -1796 39351
rect -1663 39350 -1655 39352
rect -1642 39350 -1637 39372
rect -1619 39350 -1614 39372
rect -1530 39350 -1526 39372
rect -1506 39350 -1502 39372
rect -1482 39350 -1478 39372
rect -1458 39350 -1454 39372
rect -1434 39350 -1430 39372
rect -1410 39350 -1406 39372
rect -1386 39350 -1382 39372
rect -1362 39350 -1358 39372
rect -1338 39350 -1334 39372
rect -1314 39350 -1310 39372
rect -1290 39350 -1286 39372
rect -1266 39350 -1262 39372
rect -1242 39350 -1238 39372
rect -1218 39350 -1214 39372
rect -1194 39350 -1190 39372
rect -1170 39350 -1166 39372
rect -1146 39350 -1142 39372
rect -1122 39350 -1118 39372
rect -1098 39350 -1094 39372
rect -1074 39350 -1070 39372
rect -1050 39350 -1046 39372
rect -1026 39350 -1022 39372
rect -1002 39350 -998 39372
rect -978 39350 -974 39372
rect -954 39350 -950 39372
rect -930 39350 -926 39372
rect -906 39350 -902 39372
rect -899 39371 -885 39372
rect -882 39371 -875 39395
rect -882 39350 -878 39371
rect -858 39350 -854 40284
rect -834 39350 -830 40284
rect -810 39350 -806 40284
rect -786 39350 -782 40284
rect -762 39350 -758 40284
rect -738 39350 -734 40284
rect -731 40283 -717 40284
rect -714 40283 -707 40307
rect -714 39350 -710 40283
rect -690 39350 -686 40308
rect -666 39350 -662 40308
rect -653 39701 -648 39711
rect -642 39701 -638 40308
rect -643 39687 -638 39701
rect -642 39350 -638 39687
rect -618 39635 -614 40308
rect -618 39611 -611 39635
rect -618 39350 -614 39611
rect -594 39350 -590 40308
rect -570 39350 -566 40308
rect -546 39350 -542 40308
rect -522 39350 -518 40308
rect -498 39350 -494 40308
rect -474 39350 -470 40308
rect -450 39350 -446 40308
rect -426 39350 -422 40308
rect -413 39365 -408 39375
rect -402 39365 -398 40308
rect -403 39351 -398 39365
rect -402 39350 -398 39351
rect -378 39350 -374 40308
rect -354 39350 -350 40308
rect -330 39350 -326 40308
rect -317 40301 -312 40308
rect -307 40287 -302 40301
rect -306 39350 -302 40287
rect -282 40259 -278 40404
rect -282 40211 -275 40259
rect -282 39350 -278 40211
rect -258 39350 -254 40404
rect -234 39350 -230 40404
rect -210 39350 -206 40404
rect -186 39350 -182 40404
rect -162 39350 -158 40404
rect -138 39350 -134 40404
rect -114 39350 -110 40404
rect -90 39350 -86 40404
rect -66 39350 -62 40404
rect -42 39350 -38 40404
rect -18 39350 -14 40404
rect 6 39350 10 40404
rect 30 39350 34 40404
rect 54 40379 58 40404
rect 54 40355 61 40379
rect 54 39350 58 40355
rect 78 39350 82 40404
rect 102 39350 106 40404
rect 126 39350 130 40404
rect 139 39437 144 39447
rect 150 39437 154 40404
rect 163 40133 168 40143
rect 174 40133 178 40404
rect 173 40119 178 40133
rect 163 40109 168 40119
rect 173 40095 178 40109
rect 149 39423 154 39437
rect 150 39350 154 39423
rect 174 39371 178 40095
rect 198 40067 202 40404
rect 198 40019 205 40067
rect -2393 39348 171 39350
rect -2371 39302 -2366 39348
rect -2348 39302 -2343 39348
rect -2325 39302 -2320 39348
rect -2317 39344 -2309 39348
rect -2062 39344 -2054 39348
rect -2154 39340 -2138 39342
rect -2057 39340 -2054 39344
rect -2292 39334 -2054 39340
rect -2052 39334 -2044 39344
rect -2092 39318 -2062 39320
rect -2094 39314 -2062 39318
rect -2000 39302 -1992 39348
rect -1846 39341 -1806 39348
rect -1663 39344 -1655 39348
rect -1846 39334 -1680 39340
rect -1854 39318 -1806 39320
rect -1854 39314 -1680 39318
rect -1642 39302 -1637 39348
rect -1619 39302 -1614 39348
rect -1530 39302 -1526 39348
rect -1506 39302 -1502 39348
rect -1482 39302 -1478 39348
rect -1458 39302 -1454 39348
rect -1434 39302 -1430 39348
rect -1410 39302 -1406 39348
rect -1386 39302 -1382 39348
rect -1362 39302 -1358 39348
rect -1338 39302 -1334 39348
rect -1314 39302 -1310 39348
rect -1290 39302 -1286 39348
rect -1266 39302 -1262 39348
rect -1242 39302 -1238 39348
rect -1218 39302 -1214 39348
rect -1194 39302 -1190 39348
rect -1170 39302 -1166 39348
rect -1146 39302 -1142 39348
rect -1122 39302 -1118 39348
rect -1098 39302 -1094 39348
rect -1074 39302 -1070 39348
rect -1050 39302 -1046 39348
rect -1026 39302 -1022 39348
rect -1002 39302 -998 39348
rect -978 39302 -974 39348
rect -954 39302 -950 39348
rect -930 39302 -926 39348
rect -906 39302 -902 39348
rect -882 39302 -878 39348
rect -858 39302 -854 39348
rect -834 39302 -830 39348
rect -810 39302 -806 39348
rect -786 39302 -782 39348
rect -762 39302 -758 39348
rect -738 39302 -734 39348
rect -714 39302 -710 39348
rect -690 39302 -686 39348
rect -666 39302 -662 39348
rect -642 39302 -638 39348
rect -618 39302 -614 39348
rect -594 39302 -590 39348
rect -570 39302 -566 39348
rect -546 39302 -542 39348
rect -522 39302 -518 39348
rect -498 39302 -494 39348
rect -474 39302 -470 39348
rect -450 39302 -446 39348
rect -426 39302 -422 39348
rect -402 39302 -398 39348
rect -378 39302 -374 39348
rect -354 39302 -350 39348
rect -330 39302 -326 39348
rect -306 39302 -302 39348
rect -282 39302 -278 39348
rect -258 39302 -254 39348
rect -234 39302 -230 39348
rect -210 39302 -206 39348
rect -186 39302 -182 39348
rect -162 39302 -158 39348
rect -138 39302 -134 39348
rect -114 39302 -110 39348
rect -90 39302 -86 39348
rect -66 39302 -62 39348
rect -42 39302 -38 39348
rect -18 39302 -14 39348
rect 6 39302 10 39348
rect 30 39302 34 39348
rect 54 39302 58 39348
rect 78 39302 82 39348
rect 102 39302 106 39348
rect 126 39302 130 39348
rect 150 39302 154 39348
rect 157 39347 171 39348
rect 174 39347 181 39371
rect 174 39302 178 39347
rect 198 39302 202 40019
rect 222 39302 226 40404
rect 235 39605 240 39615
rect 246 39605 250 40404
rect 253 40403 267 40404
rect 270 40403 277 40451
rect 245 39591 250 39605
rect 235 39581 240 39591
rect 245 39567 250 39581
rect 246 39302 250 39567
rect 270 39539 274 40403
rect 270 39518 277 39539
rect 294 39518 298 40764
rect 307 39557 312 39567
rect 318 39557 322 40764
rect 317 39543 322 39557
rect 318 39518 322 39543
rect 342 39518 346 40764
rect 366 39518 370 40764
rect 390 39518 394 40764
rect 414 40431 418 40764
rect 403 40430 437 40431
rect 438 40430 442 40764
rect 462 40430 466 40764
rect 486 40430 490 40764
rect 510 40430 514 40764
rect 534 40430 538 40764
rect 558 40430 562 40764
rect 582 40430 586 40764
rect 606 40430 610 40764
rect 630 40430 634 40764
rect 654 40430 658 40764
rect 661 40763 675 40764
rect 667 40757 672 40763
rect 677 40743 682 40757
rect 678 40430 682 40743
rect 691 40637 696 40647
rect 701 40623 706 40637
rect 702 40430 706 40623
rect 715 40517 720 40527
rect 725 40503 730 40517
rect 715 40469 720 40479
rect 726 40469 730 40503
rect 725 40455 730 40469
rect 715 40430 747 40431
rect 403 40428 747 40430
rect 403 40421 408 40428
rect 414 40421 418 40428
rect 413 40407 418 40421
rect 403 40397 408 40407
rect 413 40383 418 40397
rect 414 39518 418 40383
rect 438 40355 442 40428
rect 438 40334 445 40355
rect 462 40334 466 40428
rect 486 40334 490 40428
rect 510 40334 514 40428
rect 534 40334 538 40428
rect 558 40334 562 40428
rect 582 40334 586 40428
rect 606 40334 610 40428
rect 630 40334 634 40428
rect 654 40334 658 40428
rect 678 40334 682 40428
rect 702 40334 706 40428
rect 715 40421 720 40428
rect 733 40427 747 40428
rect 725 40407 730 40421
rect 726 40334 730 40407
rect 739 40334 747 40335
rect 421 40332 747 40334
rect 421 40331 435 40332
rect 438 40307 445 40332
rect 438 39518 442 40307
rect 462 39518 466 40332
rect 486 39518 490 40332
rect 510 39518 514 40332
rect 534 39518 538 40332
rect 558 39518 562 40332
rect 582 39518 586 40332
rect 606 39518 610 40332
rect 630 39518 634 40332
rect 654 39518 658 40332
rect 678 39518 682 40332
rect 702 39518 706 40332
rect 726 39518 730 40332
rect 733 40331 747 40332
rect 739 40325 744 40331
rect 749 40311 754 40325
rect 739 40277 744 40287
rect 750 40277 754 40311
rect 749 40263 754 40277
rect 739 40133 744 40143
rect 749 40119 754 40133
rect 750 39518 754 40119
rect 774 40043 781 40067
rect 774 39518 778 40043
rect 787 39605 792 39615
rect 797 39591 802 39605
rect 798 39518 802 39591
rect 811 39518 819 39519
rect 253 39516 819 39518
rect 253 39515 267 39516
rect 270 39491 277 39516
rect 270 39302 274 39491
rect 294 39302 298 39516
rect 318 39302 322 39516
rect 342 39491 346 39516
rect 342 39467 349 39491
rect 342 39302 346 39467
rect 366 39423 370 39516
rect 355 39422 389 39423
rect 390 39422 394 39516
rect 414 39422 418 39516
rect 438 39422 442 39516
rect 462 39422 466 39516
rect 486 39422 490 39516
rect 510 39422 514 39516
rect 534 39422 538 39516
rect 558 39422 562 39516
rect 582 39422 586 39516
rect 606 39422 610 39516
rect 630 39422 634 39516
rect 654 39422 658 39516
rect 678 39422 682 39516
rect 702 39422 706 39516
rect 726 39422 730 39516
rect 750 39422 754 39516
rect 774 39422 778 39516
rect 798 39422 802 39516
rect 805 39515 819 39516
rect 811 39509 816 39515
rect 821 39495 826 39509
rect 822 39422 826 39495
rect 835 39422 843 39423
rect 355 39420 843 39422
rect 355 39413 360 39420
rect 366 39413 370 39420
rect 365 39399 370 39413
rect 355 39389 360 39399
rect 365 39375 370 39389
rect 366 39302 370 39375
rect 390 39347 394 39420
rect -2393 39300 387 39302
rect -2371 39278 -2366 39300
rect -2348 39278 -2343 39300
rect -2325 39278 -2320 39300
rect -2072 39298 -2036 39299
rect -2072 39292 -2054 39298
rect -2309 39284 -2301 39292
rect -2317 39278 -2309 39284
rect -2092 39283 -2062 39288
rect -2000 39279 -1992 39300
rect -1938 39299 -1906 39300
rect -1920 39298 -1906 39299
rect -1806 39292 -1680 39298
rect -1854 39283 -1806 39288
rect -1655 39284 -1647 39292
rect -1982 39279 -1966 39280
rect -2000 39278 -1966 39279
rect -1846 39278 -1806 39281
rect -1663 39278 -1655 39284
rect -1642 39278 -1637 39300
rect -1619 39278 -1614 39300
rect -1530 39278 -1526 39300
rect -1506 39278 -1502 39300
rect -1482 39278 -1478 39300
rect -1458 39278 -1454 39300
rect -1434 39278 -1430 39300
rect -1410 39278 -1406 39300
rect -1386 39278 -1382 39300
rect -1362 39278 -1358 39300
rect -1338 39278 -1334 39300
rect -1314 39278 -1310 39300
rect -1290 39278 -1286 39300
rect -1266 39278 -1262 39300
rect -1242 39278 -1238 39300
rect -1218 39278 -1214 39300
rect -1194 39278 -1190 39300
rect -1170 39278 -1166 39300
rect -1146 39278 -1142 39300
rect -1122 39278 -1118 39300
rect -1098 39278 -1094 39300
rect -1074 39278 -1070 39300
rect -1050 39278 -1046 39300
rect -1026 39278 -1022 39300
rect -1002 39278 -998 39300
rect -978 39278 -974 39300
rect -954 39278 -950 39300
rect -930 39278 -926 39300
rect -906 39278 -902 39300
rect -882 39278 -878 39300
rect -858 39278 -854 39300
rect -834 39278 -830 39300
rect -810 39278 -806 39300
rect -786 39278 -782 39300
rect -762 39278 -758 39300
rect -738 39278 -734 39300
rect -714 39278 -710 39300
rect -690 39278 -686 39300
rect -666 39278 -662 39300
rect -642 39278 -638 39300
rect -618 39278 -614 39300
rect -594 39278 -590 39300
rect -570 39278 -566 39300
rect -546 39278 -542 39300
rect -522 39278 -518 39300
rect -498 39278 -494 39300
rect -474 39278 -470 39300
rect -450 39278 -446 39300
rect -426 39278 -422 39300
rect -402 39278 -398 39300
rect -378 39299 -374 39300
rect -2393 39276 -381 39278
rect -2371 39254 -2366 39276
rect -2348 39254 -2343 39276
rect -2325 39254 -2320 39276
rect -2000 39274 -1966 39276
rect -2309 39256 -2301 39264
rect -2062 39263 -2054 39270
rect -2092 39256 -2084 39263
rect -2062 39256 -2026 39258
rect -2317 39254 -2309 39256
rect -2062 39254 -2012 39256
rect -2000 39254 -1992 39274
rect -1982 39273 -1966 39274
rect -1846 39272 -1806 39276
rect -1846 39265 -1798 39270
rect -1806 39263 -1798 39265
rect -1854 39261 -1846 39263
rect -1854 39256 -1806 39261
rect -1655 39256 -1647 39264
rect -1864 39254 -1796 39255
rect -1663 39254 -1655 39256
rect -1642 39254 -1637 39276
rect -1619 39254 -1614 39276
rect -1530 39254 -1526 39276
rect -1506 39254 -1502 39276
rect -1482 39254 -1478 39276
rect -1458 39254 -1454 39276
rect -1434 39254 -1430 39276
rect -1410 39254 -1406 39276
rect -1386 39254 -1382 39276
rect -1362 39254 -1358 39276
rect -1338 39254 -1334 39276
rect -1314 39254 -1310 39276
rect -1290 39254 -1286 39276
rect -1266 39254 -1262 39276
rect -1242 39254 -1238 39276
rect -1218 39254 -1214 39276
rect -1194 39254 -1190 39276
rect -1170 39254 -1166 39276
rect -1146 39254 -1142 39276
rect -1122 39254 -1118 39276
rect -1098 39254 -1094 39276
rect -1074 39254 -1070 39276
rect -1050 39254 -1046 39276
rect -1026 39254 -1022 39276
rect -1002 39254 -998 39276
rect -978 39254 -974 39276
rect -954 39254 -950 39276
rect -930 39254 -926 39276
rect -906 39254 -902 39276
rect -882 39254 -878 39276
rect -858 39254 -854 39276
rect -834 39254 -830 39276
rect -810 39254 -806 39276
rect -786 39254 -782 39276
rect -762 39254 -758 39276
rect -738 39254 -734 39276
rect -714 39254 -710 39276
rect -690 39254 -686 39276
rect -666 39254 -662 39276
rect -642 39254 -638 39276
rect -618 39254 -614 39276
rect -594 39254 -590 39276
rect -570 39254 -566 39276
rect -546 39254 -542 39276
rect -522 39254 -518 39276
rect -498 39254 -494 39276
rect -474 39254 -470 39276
rect -450 39254 -446 39276
rect -426 39254 -422 39276
rect -402 39254 -398 39276
rect -395 39275 -381 39276
rect -378 39275 -371 39299
rect -378 39254 -374 39275
rect -354 39254 -350 39300
rect -330 39254 -326 39300
rect -306 39254 -302 39300
rect -282 39254 -278 39300
rect -258 39254 -254 39300
rect -234 39254 -230 39300
rect -210 39254 -206 39300
rect -186 39254 -182 39300
rect -162 39254 -158 39300
rect -138 39254 -134 39300
rect -114 39254 -110 39300
rect -90 39254 -86 39300
rect -66 39254 -62 39300
rect -42 39254 -38 39300
rect -18 39254 -14 39300
rect 6 39254 10 39300
rect 30 39254 34 39300
rect 54 39254 58 39300
rect 78 39254 82 39300
rect 102 39254 106 39300
rect 126 39254 130 39300
rect 150 39254 154 39300
rect 174 39254 178 39300
rect 198 39254 202 39300
rect 222 39254 226 39300
rect 246 39254 250 39300
rect 270 39254 274 39300
rect 294 39254 298 39300
rect 318 39254 322 39300
rect 342 39254 346 39300
rect 366 39254 370 39300
rect 373 39299 387 39300
rect 390 39299 397 39347
rect 390 39254 394 39299
rect 414 39254 418 39420
rect 438 39254 442 39420
rect 462 39254 466 39420
rect 486 39254 490 39420
rect 510 39254 514 39420
rect 534 39254 538 39420
rect 558 39254 562 39420
rect 582 39327 586 39420
rect 571 39326 605 39327
rect 606 39326 610 39420
rect 630 39326 634 39420
rect 654 39326 658 39420
rect 678 39326 682 39420
rect 691 39341 696 39351
rect 702 39341 706 39420
rect 701 39327 706 39341
rect 702 39326 706 39327
rect 726 39326 730 39420
rect 750 39326 754 39420
rect 774 39326 778 39420
rect 798 39326 802 39420
rect 822 39326 826 39420
rect 829 39419 843 39420
rect 835 39413 840 39419
rect 845 39399 850 39413
rect 846 39326 850 39399
rect 859 39326 867 39327
rect 571 39324 867 39326
rect 571 39317 576 39324
rect 582 39317 586 39324
rect 581 39303 586 39317
rect 571 39293 576 39303
rect 581 39279 586 39293
rect 582 39254 586 39279
rect 606 39254 610 39324
rect 630 39254 634 39324
rect 654 39254 658 39324
rect 678 39254 682 39324
rect 702 39254 706 39324
rect 726 39275 730 39324
rect -2393 39252 723 39254
rect -2371 39206 -2366 39252
rect -2348 39206 -2343 39252
rect -2325 39206 -2320 39252
rect -2317 39248 -2309 39252
rect -2062 39248 -2054 39252
rect -2154 39244 -2138 39246
rect -2057 39244 -2054 39248
rect -2292 39238 -2054 39244
rect -2052 39238 -2044 39248
rect -2092 39222 -2062 39224
rect -2094 39218 -2062 39222
rect -2000 39206 -1992 39252
rect -1846 39245 -1806 39252
rect -1663 39248 -1655 39252
rect -1846 39238 -1680 39244
rect -1854 39222 -1806 39224
rect -1854 39218 -1680 39222
rect -1979 39206 -1945 39208
rect -1642 39206 -1637 39252
rect -1619 39206 -1614 39252
rect -1530 39206 -1526 39252
rect -1506 39206 -1502 39252
rect -1482 39206 -1478 39252
rect -1458 39206 -1454 39252
rect -1434 39206 -1430 39252
rect -1410 39206 -1406 39252
rect -1386 39206 -1382 39252
rect -1362 39206 -1358 39252
rect -1338 39206 -1334 39252
rect -1314 39206 -1310 39252
rect -1290 39206 -1286 39252
rect -1266 39206 -1262 39252
rect -1242 39206 -1238 39252
rect -1218 39206 -1214 39252
rect -1194 39206 -1190 39252
rect -1170 39206 -1166 39252
rect -1146 39206 -1142 39252
rect -1122 39206 -1118 39252
rect -1098 39206 -1094 39252
rect -1074 39206 -1070 39252
rect -1050 39206 -1046 39252
rect -1026 39206 -1022 39252
rect -1002 39206 -998 39252
rect -978 39206 -974 39252
rect -954 39206 -950 39252
rect -930 39206 -926 39252
rect -906 39206 -902 39252
rect -882 39206 -878 39252
rect -858 39206 -854 39252
rect -834 39206 -830 39252
rect -810 39206 -806 39252
rect -786 39206 -782 39252
rect -762 39206 -758 39252
rect -738 39206 -734 39252
rect -714 39206 -710 39252
rect -690 39206 -686 39252
rect -666 39206 -662 39252
rect -653 39221 -648 39231
rect -642 39221 -638 39252
rect -643 39207 -638 39221
rect -653 39206 -619 39207
rect -2393 39204 -619 39206
rect -2371 39158 -2366 39204
rect -2348 39158 -2343 39204
rect -2325 39158 -2320 39204
rect -2080 39203 -1906 39204
rect -2080 39202 -2036 39203
rect -2080 39196 -2054 39202
rect -2309 39188 -2301 39194
rect -2317 39178 -2309 39188
rect -2070 39187 -2040 39194
rect -2054 39179 -2040 39182
rect -2000 39177 -1992 39203
rect -1920 39202 -1906 39203
rect -1850 39196 -1846 39204
rect -1840 39196 -1792 39204
rect -1969 39184 -1966 39193
rect -1850 39189 -1802 39194
rect -1906 39187 -1802 39189
rect -1655 39188 -1647 39194
rect -1906 39186 -1850 39187
rect -1846 39179 -1802 39185
rect -1663 39178 -1655 39188
rect -1860 39177 -1798 39178
rect -2078 39170 -2070 39177
rect -2309 39160 -2301 39166
rect -2317 39158 -2309 39160
rect -2154 39158 -2145 39168
rect -2044 39167 -2040 39172
rect -2028 39170 -1945 39177
rect -1929 39170 -1794 39177
rect -2070 39160 -2040 39167
rect -2044 39158 -2028 39160
rect -2000 39158 -1992 39170
rect -1860 39169 -1798 39170
rect -1850 39160 -1802 39167
rect -1655 39160 -1647 39166
rect -1978 39158 -1942 39159
rect -1663 39158 -1655 39160
rect -1642 39158 -1637 39204
rect -1619 39158 -1614 39204
rect -1530 39158 -1526 39204
rect -1506 39158 -1502 39204
rect -1482 39158 -1478 39204
rect -1458 39158 -1454 39204
rect -1434 39158 -1430 39204
rect -1410 39158 -1406 39204
rect -1386 39158 -1382 39204
rect -1362 39158 -1358 39204
rect -1338 39158 -1334 39204
rect -1314 39158 -1310 39204
rect -1290 39158 -1286 39204
rect -1266 39158 -1262 39204
rect -1242 39158 -1238 39204
rect -1218 39158 -1214 39204
rect -1194 39158 -1190 39204
rect -1170 39158 -1166 39204
rect -1146 39158 -1142 39204
rect -1122 39158 -1118 39204
rect -1098 39158 -1094 39204
rect -1074 39158 -1070 39204
rect -1050 39158 -1046 39204
rect -1026 39158 -1022 39204
rect -1002 39158 -998 39204
rect -978 39158 -974 39204
rect -954 39158 -950 39204
rect -930 39158 -926 39204
rect -906 39158 -902 39204
rect -882 39158 -878 39204
rect -858 39158 -854 39204
rect -834 39158 -830 39204
rect -810 39158 -806 39204
rect -786 39158 -782 39204
rect -762 39158 -758 39204
rect -738 39158 -734 39204
rect -714 39158 -710 39204
rect -690 39158 -686 39204
rect -666 39158 -662 39204
rect -653 39197 -648 39204
rect -643 39183 -638 39197
rect -642 39158 -638 39183
rect -618 39158 -614 39252
rect -594 39158 -590 39252
rect -570 39158 -566 39252
rect -546 39158 -542 39252
rect -522 39158 -518 39252
rect -498 39158 -494 39252
rect -474 39158 -470 39252
rect -450 39158 -446 39252
rect -426 39158 -422 39252
rect -402 39158 -398 39252
rect -378 39158 -374 39252
rect -354 39158 -350 39252
rect -330 39158 -326 39252
rect -306 39158 -302 39252
rect -282 39158 -278 39252
rect -258 39158 -254 39252
rect -234 39158 -230 39252
rect -210 39158 -206 39252
rect -186 39158 -182 39252
rect -162 39158 -158 39252
rect -138 39158 -134 39252
rect -114 39158 -110 39252
rect -90 39158 -86 39252
rect -66 39158 -62 39252
rect -42 39158 -38 39252
rect -18 39158 -14 39252
rect 6 39158 10 39252
rect 30 39158 34 39252
rect 54 39158 58 39252
rect 78 39158 82 39252
rect 102 39158 106 39252
rect 126 39158 130 39252
rect 150 39158 154 39252
rect 174 39158 178 39252
rect 198 39158 202 39252
rect 222 39158 226 39252
rect 246 39158 250 39252
rect 270 39158 274 39252
rect 294 39158 298 39252
rect 318 39158 322 39252
rect 342 39158 346 39252
rect 366 39158 370 39252
rect 390 39158 394 39252
rect 414 39158 418 39252
rect 438 39158 442 39252
rect 462 39158 466 39252
rect 486 39158 490 39252
rect 510 39159 514 39252
rect 499 39158 533 39159
rect -2393 39156 533 39158
rect -2371 39038 -2366 39156
rect -2348 39038 -2343 39156
rect -2325 39118 -2320 39156
rect -2317 39150 -2309 39156
rect -2145 39152 -2138 39156
rect -2070 39152 -2054 39156
rect -2078 39143 -2054 39150
rect -2062 39118 -2032 39119
rect -2000 39118 -1992 39156
rect -1846 39152 -1802 39156
rect -1846 39142 -1792 39151
rect -1663 39150 -1655 39156
rect -1942 39120 -1937 39132
rect -1850 39129 -1822 39130
rect -1850 39125 -1802 39129
rect -2325 39110 -2317 39118
rect -2062 39116 -1961 39118
rect -2325 39090 -2320 39110
rect -2317 39102 -2309 39110
rect -2062 39103 -2040 39114
rect -2032 39109 -1961 39116
rect -1947 39110 -1942 39118
rect -1842 39116 -1794 39119
rect -2070 39098 -2022 39102
rect -2325 39078 -2317 39090
rect -2137 39081 -2121 39083
rect -2325 39062 -2320 39078
rect -2317 39074 -2309 39078
rect -2292 39076 -2085 39081
rect -2069 39076 -2032 39078
rect -2309 39062 -2301 39074
rect -2125 39070 -2121 39071
rect -2325 39050 -2317 39062
rect -2059 39054 -2045 39058
rect -2325 39038 -2320 39050
rect -2317 39046 -2309 39050
rect -2309 39038 -2301 39046
rect -2025 39042 -2022 39048
rect -2000 39042 -1992 39109
rect -1942 39108 -1937 39110
rect -1932 39100 -1927 39108
rect -1912 39105 -1896 39111
rect -1842 39103 -1802 39114
rect -1671 39110 -1663 39118
rect -1663 39102 -1655 39110
rect -1850 39098 -1680 39102
rect -1671 39078 -1663 39090
rect -1663 39074 -1655 39078
rect -1977 39067 -1929 39073
rect -1974 39058 -1944 39067
rect -1655 39062 -1647 39074
rect -1960 39057 -1944 39058
rect -1671 39050 -1663 39062
rect -1977 39045 -1929 39047
rect -1663 39046 -1655 39050
rect -2033 39040 -1992 39042
rect -2062 39038 -1992 39040
rect -1655 39038 -1647 39046
rect -1642 39038 -1637 39156
rect -1619 39038 -1614 39156
rect -1530 39038 -1526 39156
rect -1506 39038 -1502 39156
rect -1482 39038 -1478 39156
rect -1458 39038 -1454 39156
rect -1434 39038 -1430 39156
rect -1410 39038 -1406 39156
rect -1386 39038 -1382 39156
rect -1362 39038 -1358 39156
rect -1338 39038 -1334 39156
rect -1314 39039 -1310 39156
rect -1325 39038 -1291 39039
rect -2393 39036 -1291 39038
rect -2371 38942 -2366 39036
rect -2348 38942 -2343 39036
rect -2325 39034 -2320 39036
rect -2309 39034 -2301 39036
rect -2325 39022 -2317 39034
rect -2025 39032 -2022 39036
rect -2062 39022 -2032 39023
rect -2325 39002 -2320 39022
rect -2317 39018 -2309 39022
rect -2325 38994 -2317 39002
rect -2325 38942 -2320 38994
rect -2317 38986 -2309 38994
rect -2117 38985 -2095 38995
rect -2045 38992 -2037 39006
rect -2309 38946 -2301 38956
rect -2087 38952 -2076 38960
rect -2017 38956 -2015 38963
rect -2317 38942 -2309 38946
rect -2092 38944 -2087 38952
rect -2092 38942 -2077 38943
rect -2000 38942 -1992 39036
rect -1888 39029 -1874 39036
rect -1655 39034 -1647 39036
rect -1671 39022 -1663 39034
rect -1663 39018 -1655 39022
rect -1969 38985 -1929 38997
rect -1671 38994 -1663 39002
rect -1663 38986 -1655 38994
rect -1655 38946 -1647 38956
rect -1928 38942 -1924 38943
rect -1854 38942 -1680 38943
rect -1663 38942 -1655 38946
rect -1642 38942 -1637 39036
rect -1619 38942 -1614 39036
rect -1530 38943 -1526 39036
rect -1541 38942 -1507 38943
rect -2393 38940 -1507 38942
rect -2371 38918 -2366 38940
rect -2348 38918 -2343 38940
rect -2325 38918 -2320 38940
rect -2092 38935 -2037 38940
rect -2021 38935 -1969 38940
rect -1921 38935 -1913 38940
rect -1854 38936 -1680 38940
rect -2100 38933 -2092 38934
rect -2309 38918 -2301 38928
rect -2100 38927 -2087 38933
rect -2051 38920 -2026 38922
rect -2062 38918 -2012 38920
rect -2000 38918 -1992 38935
rect -1969 38927 -1921 38934
rect -1969 38918 -1964 38927
rect -1864 38918 -1796 38919
rect -1655 38918 -1647 38928
rect -1642 38918 -1637 38940
rect -1619 38918 -1614 38940
rect -1541 38933 -1536 38940
rect -1530 38933 -1526 38940
rect -1531 38919 -1526 38933
rect -1530 38918 -1526 38919
rect -1506 38918 -1502 39036
rect -1482 38918 -1478 39036
rect -1458 38918 -1454 39036
rect -1434 38918 -1430 39036
rect -1410 38918 -1406 39036
rect -1386 38918 -1382 39036
rect -1362 38918 -1358 39036
rect -1338 38918 -1334 39036
rect -1325 39029 -1320 39036
rect -1314 39029 -1310 39036
rect -1315 39015 -1310 39029
rect -1314 38918 -1310 39015
rect -1290 38963 -1286 39156
rect -1290 38939 -1283 38963
rect -1290 38918 -1286 38939
rect -1266 38918 -1262 39156
rect -1242 38918 -1238 39156
rect -1218 38918 -1214 39156
rect -1194 38918 -1190 39156
rect -1170 38918 -1166 39156
rect -1146 38918 -1142 39156
rect -1122 38918 -1118 39156
rect -1098 38918 -1094 39156
rect -1074 38918 -1070 39156
rect -1050 38918 -1046 39156
rect -1026 38918 -1022 39156
rect -1002 38918 -998 39156
rect -978 38918 -974 39156
rect -954 38918 -950 39156
rect -930 38918 -926 39156
rect -906 38918 -902 39156
rect -882 38918 -878 39156
rect -858 38918 -854 39156
rect -834 38918 -830 39156
rect -810 39111 -806 39156
rect -821 39110 -787 39111
rect -786 39110 -782 39156
rect -762 39110 -758 39156
rect -738 39110 -734 39156
rect -714 39110 -710 39156
rect -690 39110 -686 39156
rect -666 39110 -662 39156
rect -642 39110 -638 39156
rect -618 39155 -614 39156
rect -618 39134 -611 39155
rect -594 39134 -590 39156
rect -570 39134 -566 39156
rect -546 39134 -542 39156
rect -522 39134 -518 39156
rect -498 39134 -494 39156
rect -474 39134 -470 39156
rect -450 39134 -446 39156
rect -426 39134 -422 39156
rect -402 39134 -398 39156
rect -378 39135 -374 39156
rect -389 39134 -355 39135
rect -635 39132 -355 39134
rect -635 39131 -621 39132
rect -821 39108 -621 39110
rect -821 39101 -816 39108
rect -810 39101 -806 39108
rect -811 39087 -806 39101
rect -821 39077 -816 39087
rect -811 39063 -806 39077
rect -810 38918 -806 39063
rect -786 39035 -782 39108
rect -786 39014 -779 39035
rect -762 39014 -758 39108
rect -738 39014 -734 39108
rect -714 39014 -710 39108
rect -690 39014 -686 39108
rect -666 39014 -662 39108
rect -642 39014 -638 39108
rect -635 39107 -621 39108
rect -618 39107 -611 39132
rect -618 39014 -614 39107
rect -594 39014 -590 39132
rect -570 39014 -566 39132
rect -546 39014 -542 39132
rect -522 39014 -518 39132
rect -498 39014 -494 39132
rect -474 39014 -470 39132
rect -450 39014 -446 39132
rect -426 39014 -422 39132
rect -402 39014 -398 39132
rect -389 39125 -384 39132
rect -378 39125 -374 39132
rect -379 39111 -374 39125
rect -378 39014 -374 39111
rect -354 39059 -350 39156
rect -354 39035 -347 39059
rect -354 39014 -350 39035
rect -330 39014 -326 39156
rect -306 39014 -302 39156
rect -282 39014 -278 39156
rect -258 39014 -254 39156
rect -234 39014 -230 39156
rect -210 39014 -206 39156
rect -186 39014 -182 39156
rect -162 39014 -158 39156
rect -138 39014 -134 39156
rect -114 39014 -110 39156
rect -90 39014 -86 39156
rect -66 39014 -62 39156
rect -42 39014 -38 39156
rect -18 39014 -14 39156
rect 6 39014 10 39156
rect 30 39014 34 39156
rect 54 39014 58 39156
rect 78 39014 82 39156
rect 102 39014 106 39156
rect 126 39014 130 39156
rect 150 39014 154 39156
rect 174 39014 178 39156
rect 198 39014 202 39156
rect 222 39014 226 39156
rect 246 39014 250 39156
rect 270 39014 274 39156
rect 294 39014 298 39156
rect 318 39014 322 39156
rect 342 39014 346 39156
rect 366 39014 370 39156
rect 390 39014 394 39156
rect 414 39014 418 39156
rect 438 39014 442 39156
rect 462 39014 466 39156
rect 486 39014 490 39156
rect 499 39149 504 39156
rect 510 39149 514 39156
rect 509 39135 514 39149
rect 510 39014 514 39135
rect 534 39083 538 39252
rect 534 39059 541 39083
rect 534 39014 538 39059
rect 558 39014 562 39252
rect 582 39014 586 39252
rect 606 39251 610 39252
rect 606 39230 613 39251
rect 630 39230 634 39252
rect 654 39230 658 39252
rect 678 39230 682 39252
rect 702 39230 706 39252
rect 709 39251 723 39252
rect 726 39251 733 39275
rect 726 39230 730 39251
rect 750 39230 754 39324
rect 774 39230 778 39324
rect 798 39230 802 39324
rect 822 39230 826 39324
rect 835 39245 840 39255
rect 846 39245 850 39324
rect 853 39323 867 39324
rect 859 39317 864 39323
rect 869 39303 874 39317
rect 859 39269 864 39279
rect 870 39269 874 39303
rect 869 39255 874 39269
rect 845 39231 850 39245
rect 835 39230 869 39231
rect 589 39228 869 39230
rect 589 39227 603 39228
rect 606 39203 613 39228
rect 606 39014 610 39203
rect 630 39014 634 39228
rect 654 39015 658 39228
rect 643 39014 677 39015
rect -803 39012 677 39014
rect -803 39011 -789 39012
rect -786 38987 -779 39012
rect -786 38918 -782 38987
rect -762 38918 -758 39012
rect -738 38918 -734 39012
rect -714 38918 -710 39012
rect -690 38918 -686 39012
rect -666 38918 -662 39012
rect -642 38918 -638 39012
rect -618 38918 -614 39012
rect -594 38918 -590 39012
rect -570 38918 -566 39012
rect -546 38918 -542 39012
rect -522 38918 -518 39012
rect -498 38918 -494 39012
rect -474 38918 -470 39012
rect -450 38918 -446 39012
rect -426 38918 -422 39012
rect -402 38918 -398 39012
rect -378 38918 -374 39012
rect -354 38918 -350 39012
rect -330 38918 -326 39012
rect -306 38918 -302 39012
rect -282 38919 -278 39012
rect -293 38918 -259 38919
rect -2393 38916 -259 38918
rect -2371 38870 -2366 38916
rect -2348 38870 -2343 38916
rect -2325 38870 -2320 38916
rect -2317 38912 -2309 38916
rect -2105 38909 -2092 38912
rect -2092 38886 -2062 38888
rect -2094 38882 -2062 38886
rect -2000 38870 -1992 38916
rect -1663 38912 -1655 38916
rect -1969 38909 -1921 38912
rect -1854 38886 -1806 38888
rect -1854 38882 -1680 38886
rect -1642 38870 -1637 38916
rect -1619 38870 -1614 38916
rect -1530 38870 -1526 38916
rect -1506 38870 -1502 38916
rect -1482 38870 -1478 38916
rect -1458 38870 -1454 38916
rect -1434 38870 -1430 38916
rect -1410 38870 -1406 38916
rect -1386 38870 -1382 38916
rect -1362 38870 -1358 38916
rect -1338 38870 -1334 38916
rect -1314 38870 -1310 38916
rect -1290 38870 -1286 38916
rect -1266 38870 -1262 38916
rect -1242 38870 -1238 38916
rect -1218 38870 -1214 38916
rect -1194 38870 -1190 38916
rect -1170 38870 -1166 38916
rect -1146 38870 -1142 38916
rect -1122 38870 -1118 38916
rect -1098 38870 -1094 38916
rect -1074 38870 -1070 38916
rect -1050 38870 -1046 38916
rect -1026 38870 -1022 38916
rect -1002 38870 -998 38916
rect -978 38870 -974 38916
rect -954 38870 -950 38916
rect -930 38870 -926 38916
rect -906 38870 -902 38916
rect -882 38870 -878 38916
rect -858 38870 -854 38916
rect -834 38870 -830 38916
rect -810 38870 -806 38916
rect -786 38870 -782 38916
rect -762 38870 -758 38916
rect -738 38870 -734 38916
rect -714 38870 -710 38916
rect -690 38870 -686 38916
rect -666 38870 -662 38916
rect -642 38870 -638 38916
rect -618 38870 -614 38916
rect -594 38870 -590 38916
rect -570 38870 -566 38916
rect -546 38870 -542 38916
rect -522 38870 -518 38916
rect -498 38870 -494 38916
rect -474 38870 -470 38916
rect -450 38870 -446 38916
rect -426 38870 -422 38916
rect -402 38870 -398 38916
rect -378 38870 -374 38916
rect -365 38885 -360 38895
rect -354 38885 -350 38916
rect -355 38871 -350 38885
rect -365 38870 -331 38871
rect -2393 38868 -331 38870
rect -2371 38846 -2366 38868
rect -2348 38846 -2343 38868
rect -2325 38846 -2320 38868
rect -2072 38866 -2036 38867
rect -2072 38860 -2054 38866
rect -2309 38852 -2301 38860
rect -2317 38846 -2309 38852
rect -2092 38851 -2062 38856
rect -2000 38847 -1992 38868
rect -1938 38867 -1906 38868
rect -1920 38866 -1906 38867
rect -1806 38860 -1680 38866
rect -1854 38851 -1806 38856
rect -1655 38852 -1647 38860
rect -1982 38847 -1966 38848
rect -2000 38846 -1966 38847
rect -1846 38846 -1806 38849
rect -1663 38846 -1655 38852
rect -1642 38846 -1637 38868
rect -1619 38846 -1614 38868
rect -1589 38846 -1555 38847
rect -2393 38844 -1555 38846
rect -2371 38822 -2366 38844
rect -2348 38822 -2343 38844
rect -2325 38822 -2320 38844
rect -2000 38842 -1966 38844
rect -2309 38824 -2301 38832
rect -2062 38831 -2054 38838
rect -2092 38824 -2084 38831
rect -2062 38824 -2026 38826
rect -2317 38822 -2309 38824
rect -2062 38822 -2012 38824
rect -2000 38822 -1992 38842
rect -1982 38841 -1966 38842
rect -1846 38840 -1806 38844
rect -1846 38833 -1798 38838
rect -1806 38831 -1798 38833
rect -1854 38829 -1846 38831
rect -1854 38824 -1806 38829
rect -1655 38824 -1647 38832
rect -1864 38822 -1796 38823
rect -1663 38822 -1655 38824
rect -1642 38822 -1637 38844
rect -1619 38822 -1614 38844
rect -1530 38822 -1526 38868
rect -1506 38867 -1502 38868
rect -1506 38843 -1499 38867
rect -1506 38822 -1502 38843
rect -1482 38822 -1478 38868
rect -1458 38822 -1454 38868
rect -1434 38822 -1430 38868
rect -1410 38822 -1406 38868
rect -1386 38822 -1382 38868
rect -1362 38822 -1358 38868
rect -1338 38822 -1334 38868
rect -1314 38822 -1310 38868
rect -1290 38822 -1286 38868
rect -1266 38822 -1262 38868
rect -1242 38822 -1238 38868
rect -1218 38822 -1214 38868
rect -1194 38822 -1190 38868
rect -1170 38822 -1166 38868
rect -1146 38822 -1142 38868
rect -1122 38822 -1118 38868
rect -1098 38822 -1094 38868
rect -1074 38822 -1070 38868
rect -1050 38822 -1046 38868
rect -1026 38822 -1022 38868
rect -1002 38822 -998 38868
rect -978 38822 -974 38868
rect -954 38822 -950 38868
rect -930 38822 -926 38868
rect -906 38822 -902 38868
rect -882 38822 -878 38868
rect -858 38822 -854 38868
rect -834 38822 -830 38868
rect -810 38822 -806 38868
rect -786 38822 -782 38868
rect -762 38822 -758 38868
rect -738 38822 -734 38868
rect -714 38822 -710 38868
rect -690 38822 -686 38868
rect -666 38822 -662 38868
rect -642 38822 -638 38868
rect -618 38822 -614 38868
rect -594 38822 -590 38868
rect -570 38822 -566 38868
rect -546 38822 -542 38868
rect -522 38822 -518 38868
rect -498 38822 -494 38868
rect -474 38822 -470 38868
rect -450 38822 -446 38868
rect -426 38822 -422 38868
rect -402 38822 -398 38868
rect -378 38822 -374 38868
rect -365 38861 -360 38868
rect -355 38847 -350 38861
rect -354 38822 -350 38847
rect -330 38822 -326 38916
rect -306 38822 -302 38916
rect -293 38909 -288 38916
rect -282 38909 -278 38916
rect -283 38895 -278 38909
rect -282 38823 -278 38895
rect -258 38843 -254 39012
rect -293 38822 -261 38823
rect -2393 38820 -261 38822
rect -2371 38774 -2366 38820
rect -2348 38774 -2343 38820
rect -2325 38774 -2320 38820
rect -2317 38816 -2309 38820
rect -2062 38816 -2054 38820
rect -2154 38812 -2138 38814
rect -2057 38812 -2054 38816
rect -2292 38806 -2054 38812
rect -2052 38806 -2044 38816
rect -2092 38790 -2062 38792
rect -2094 38786 -2062 38790
rect -2000 38774 -1992 38820
rect -1846 38813 -1806 38820
rect -1663 38816 -1655 38820
rect -1846 38806 -1680 38812
rect -1854 38790 -1806 38792
rect -1854 38786 -1680 38790
rect -1642 38774 -1637 38820
rect -1619 38774 -1614 38820
rect -1530 38774 -1526 38820
rect -1506 38774 -1502 38820
rect -1482 38774 -1478 38820
rect -1458 38774 -1454 38820
rect -1434 38774 -1430 38820
rect -1410 38774 -1406 38820
rect -1386 38774 -1382 38820
rect -1362 38774 -1358 38820
rect -1338 38774 -1334 38820
rect -1314 38774 -1310 38820
rect -1290 38774 -1286 38820
rect -1266 38774 -1262 38820
rect -1242 38774 -1238 38820
rect -1218 38774 -1214 38820
rect -1194 38774 -1190 38820
rect -1170 38774 -1166 38820
rect -1146 38774 -1142 38820
rect -1122 38774 -1118 38820
rect -1098 38774 -1094 38820
rect -1074 38774 -1070 38820
rect -1050 38774 -1046 38820
rect -1026 38774 -1022 38820
rect -1002 38774 -998 38820
rect -978 38774 -974 38820
rect -954 38774 -950 38820
rect -930 38774 -926 38820
rect -906 38774 -902 38820
rect -882 38774 -878 38820
rect -858 38774 -854 38820
rect -834 38774 -830 38820
rect -810 38774 -806 38820
rect -786 38774 -782 38820
rect -762 38774 -758 38820
rect -738 38774 -734 38820
rect -714 38774 -710 38820
rect -690 38774 -686 38820
rect -666 38774 -662 38820
rect -642 38774 -638 38820
rect -618 38774 -614 38820
rect -594 38774 -590 38820
rect -570 38774 -566 38820
rect -546 38774 -542 38820
rect -522 38774 -518 38820
rect -498 38774 -494 38820
rect -474 38774 -470 38820
rect -450 38774 -446 38820
rect -426 38774 -422 38820
rect -402 38774 -398 38820
rect -378 38774 -374 38820
rect -354 38774 -350 38820
rect -330 38819 -326 38820
rect -2393 38772 -333 38774
rect -2371 38750 -2366 38772
rect -2348 38750 -2343 38772
rect -2325 38750 -2320 38772
rect -2072 38770 -2036 38771
rect -2072 38764 -2054 38770
rect -2309 38756 -2301 38764
rect -2317 38750 -2309 38756
rect -2092 38755 -2062 38760
rect -2000 38751 -1992 38772
rect -1938 38771 -1906 38772
rect -1920 38770 -1906 38771
rect -1806 38764 -1680 38770
rect -1854 38755 -1806 38760
rect -1655 38756 -1647 38764
rect -1982 38751 -1966 38752
rect -2000 38750 -1966 38751
rect -1846 38750 -1806 38753
rect -1663 38750 -1655 38756
rect -1642 38750 -1637 38772
rect -1619 38750 -1614 38772
rect -1554 38758 -1547 38771
rect -2393 38748 -1557 38750
rect -2371 38726 -2366 38748
rect -2348 38726 -2343 38748
rect -2325 38726 -2320 38748
rect -2000 38746 -1966 38748
rect -2309 38728 -2301 38736
rect -2062 38735 -2054 38742
rect -2092 38728 -2084 38735
rect -2062 38728 -2026 38730
rect -2317 38726 -2309 38728
rect -2062 38726 -2012 38728
rect -2000 38726 -1992 38746
rect -1982 38745 -1966 38746
rect -1846 38744 -1806 38748
rect -1846 38737 -1798 38742
rect -1806 38735 -1798 38737
rect -1854 38733 -1846 38735
rect -1854 38728 -1806 38733
rect -1655 38728 -1647 38736
rect -1864 38726 -1796 38727
rect -1663 38726 -1655 38728
rect -1642 38726 -1637 38748
rect -1619 38726 -1614 38748
rect -1571 38747 -1557 38748
rect -1554 38747 -1547 38748
rect -1530 38726 -1526 38772
rect -1506 38726 -1502 38772
rect -1482 38726 -1478 38772
rect -1458 38726 -1454 38772
rect -1434 38726 -1430 38772
rect -1410 38726 -1406 38772
rect -1386 38726 -1382 38772
rect -1362 38726 -1358 38772
rect -1338 38726 -1334 38772
rect -1314 38726 -1310 38772
rect -1290 38726 -1286 38772
rect -1266 38726 -1262 38772
rect -1253 38741 -1248 38751
rect -1242 38741 -1238 38772
rect -1243 38727 -1238 38741
rect -1242 38726 -1238 38727
rect -1218 38726 -1214 38772
rect -1194 38726 -1190 38772
rect -1170 38726 -1166 38772
rect -1146 38726 -1142 38772
rect -1122 38726 -1118 38772
rect -1098 38726 -1094 38772
rect -1074 38726 -1070 38772
rect -1050 38726 -1046 38772
rect -1026 38726 -1022 38772
rect -1002 38726 -998 38772
rect -978 38726 -974 38772
rect -954 38726 -950 38772
rect -930 38726 -926 38772
rect -906 38726 -902 38772
rect -882 38726 -878 38772
rect -858 38726 -854 38772
rect -834 38726 -830 38772
rect -810 38726 -806 38772
rect -786 38726 -782 38772
rect -762 38726 -758 38772
rect -738 38726 -734 38772
rect -714 38726 -710 38772
rect -690 38726 -686 38772
rect -666 38726 -662 38772
rect -642 38726 -638 38772
rect -618 38726 -614 38772
rect -594 38726 -590 38772
rect -570 38726 -566 38772
rect -546 38726 -542 38772
rect -522 38726 -518 38772
rect -498 38726 -494 38772
rect -474 38726 -470 38772
rect -450 38726 -446 38772
rect -426 38726 -422 38772
rect -402 38726 -398 38772
rect -378 38726 -374 38772
rect -354 38726 -350 38772
rect -347 38771 -333 38772
rect -330 38771 -323 38819
rect -330 38726 -326 38771
rect -306 38726 -302 38820
rect -293 38813 -288 38820
rect -282 38813 -278 38820
rect -275 38819 -261 38820
rect -258 38819 -251 38843
rect -283 38799 -278 38813
rect -282 38726 -278 38799
rect -258 38747 -254 38819
rect -2393 38724 -261 38726
rect -2371 38678 -2366 38724
rect -2348 38678 -2343 38724
rect -2325 38678 -2320 38724
rect -2317 38720 -2309 38724
rect -2062 38720 -2054 38724
rect -2154 38716 -2138 38718
rect -2057 38716 -2054 38720
rect -2292 38710 -2054 38716
rect -2052 38710 -2044 38720
rect -2092 38694 -2062 38696
rect -2094 38690 -2062 38694
rect -2000 38678 -1992 38724
rect -1846 38717 -1806 38724
rect -1663 38720 -1655 38724
rect -1846 38710 -1680 38716
rect -1854 38694 -1806 38696
rect -1854 38690 -1680 38694
rect -1642 38678 -1637 38724
rect -1619 38678 -1614 38724
rect -1530 38678 -1526 38724
rect -1506 38678 -1502 38724
rect -1482 38678 -1478 38724
rect -1458 38678 -1454 38724
rect -1434 38678 -1430 38724
rect -1410 38678 -1406 38724
rect -1386 38678 -1382 38724
rect -1362 38678 -1358 38724
rect -1338 38678 -1334 38724
rect -1314 38678 -1310 38724
rect -1290 38678 -1286 38724
rect -1266 38678 -1262 38724
rect -1242 38678 -1238 38724
rect -1218 38678 -1214 38724
rect -1194 38678 -1190 38724
rect -1170 38678 -1166 38724
rect -1146 38678 -1142 38724
rect -1122 38678 -1118 38724
rect -1098 38678 -1094 38724
rect -1074 38678 -1070 38724
rect -1050 38678 -1046 38724
rect -1026 38678 -1022 38724
rect -1002 38678 -998 38724
rect -978 38678 -974 38724
rect -954 38678 -950 38724
rect -930 38678 -926 38724
rect -906 38678 -902 38724
rect -882 38678 -878 38724
rect -858 38678 -854 38724
rect -834 38678 -830 38724
rect -810 38678 -806 38724
rect -786 38678 -782 38724
rect -762 38678 -758 38724
rect -738 38678 -734 38724
rect -714 38678 -710 38724
rect -690 38678 -686 38724
rect -666 38678 -662 38724
rect -642 38678 -638 38724
rect -618 38678 -614 38724
rect -594 38678 -590 38724
rect -570 38678 -566 38724
rect -546 38678 -542 38724
rect -522 38678 -518 38724
rect -498 38678 -494 38724
rect -474 38678 -470 38724
rect -450 38678 -446 38724
rect -426 38678 -422 38724
rect -402 38678 -398 38724
rect -378 38678 -374 38724
rect -354 38678 -350 38724
rect -330 38678 -326 38724
rect -306 38678 -302 38724
rect -282 38678 -278 38724
rect -275 38723 -261 38724
rect -258 38723 -251 38747
rect -258 38678 -254 38723
rect -234 38678 -230 39012
rect -210 38799 -206 39012
rect -221 38798 -187 38799
rect -186 38798 -182 39012
rect -162 38798 -158 39012
rect -138 38798 -134 39012
rect -114 38798 -110 39012
rect -90 38798 -86 39012
rect -66 38798 -62 39012
rect -42 38798 -38 39012
rect -18 38798 -14 39012
rect 6 38798 10 39012
rect 30 38798 34 39012
rect 54 38798 58 39012
rect 78 38798 82 39012
rect 91 38981 96 38991
rect 102 38981 106 39012
rect 101 38967 106 38981
rect 91 38957 96 38967
rect 101 38943 106 38957
rect 102 38798 106 38943
rect 126 38915 130 39012
rect 126 38894 133 38915
rect 150 38894 154 39012
rect 174 38894 178 39012
rect 198 38894 202 39012
rect 222 38894 226 39012
rect 246 38894 250 39012
rect 270 38894 274 39012
rect 294 38894 298 39012
rect 318 38894 322 39012
rect 342 38894 346 39012
rect 366 38894 370 39012
rect 390 38894 394 39012
rect 414 38894 418 39012
rect 438 38894 442 39012
rect 462 38894 466 39012
rect 486 38894 490 39012
rect 510 38894 514 39012
rect 534 38894 538 39012
rect 558 38894 562 39012
rect 582 38894 586 39012
rect 606 38894 610 39012
rect 630 38894 634 39012
rect 643 39005 648 39012
rect 654 39005 658 39012
rect 653 38991 658 39005
rect 654 38894 658 38991
rect 678 38939 682 39228
rect 678 38915 685 38939
rect 678 38894 682 38915
rect 702 38894 706 39228
rect 726 38894 730 39228
rect 750 38894 754 39228
rect 774 38894 778 39228
rect 798 38894 802 39228
rect 822 38894 826 39228
rect 835 39221 840 39228
rect 845 39207 850 39221
rect 846 38894 850 39207
rect 859 39101 864 39111
rect 869 39087 874 39101
rect 870 38894 874 39087
rect 883 38981 888 38991
rect 893 38967 898 38981
rect 894 38894 898 38967
rect 907 38894 915 38895
rect 109 38892 915 38894
rect 109 38891 123 38892
rect 126 38867 133 38892
rect 126 38798 130 38867
rect 150 38798 154 38892
rect 174 38798 178 38892
rect 198 38798 202 38892
rect 222 38798 226 38892
rect 246 38798 250 38892
rect 270 38798 274 38892
rect 294 38798 298 38892
rect 318 38798 322 38892
rect 342 38798 346 38892
rect 366 38798 370 38892
rect 390 38798 394 38892
rect 414 38798 418 38892
rect 438 38798 442 38892
rect 462 38798 466 38892
rect 486 38798 490 38892
rect 510 38798 514 38892
rect 534 38798 538 38892
rect 558 38798 562 38892
rect 582 38798 586 38892
rect 606 38798 610 38892
rect 630 38798 634 38892
rect 654 38798 658 38892
rect 678 38798 682 38892
rect 702 38798 706 38892
rect 726 38798 730 38892
rect 750 38798 754 38892
rect 774 38798 778 38892
rect 798 38798 802 38892
rect 822 38798 826 38892
rect 846 38798 850 38892
rect 870 38798 874 38892
rect 894 38798 898 38892
rect 901 38891 915 38892
rect 907 38885 912 38891
rect 917 38871 922 38885
rect 918 38798 922 38871
rect 931 38798 939 38799
rect -221 38796 939 38798
rect -221 38789 -216 38796
rect -210 38789 -206 38796
rect -211 38775 -206 38789
rect -221 38765 -216 38775
rect -211 38751 -206 38765
rect -210 38678 -206 38751
rect -186 38723 -182 38796
rect -2393 38676 -189 38678
rect -2371 38654 -2366 38676
rect -2348 38654 -2343 38676
rect -2325 38654 -2320 38676
rect -2072 38674 -2036 38675
rect -2072 38668 -2054 38674
rect -2309 38660 -2301 38668
rect -2317 38654 -2309 38660
rect -2092 38659 -2062 38664
rect -2000 38655 -1992 38676
rect -1938 38675 -1906 38676
rect -1920 38674 -1906 38675
rect -1806 38668 -1680 38674
rect -1854 38659 -1806 38664
rect -1655 38660 -1647 38668
rect -1982 38655 -1966 38656
rect -2000 38654 -1966 38655
rect -1846 38654 -1806 38657
rect -1663 38654 -1655 38660
rect -1642 38654 -1637 38676
rect -1619 38654 -1614 38676
rect -1530 38654 -1526 38676
rect -1506 38654 -1502 38676
rect -1482 38654 -1478 38676
rect -1458 38654 -1454 38676
rect -1434 38654 -1430 38676
rect -1410 38654 -1406 38676
rect -1386 38654 -1382 38676
rect -1362 38654 -1358 38676
rect -1338 38654 -1334 38676
rect -1314 38654 -1310 38676
rect -1290 38654 -1286 38676
rect -1266 38654 -1262 38676
rect -1242 38654 -1238 38676
rect -1218 38675 -1214 38676
rect -2393 38652 -1221 38654
rect -2371 38630 -2366 38652
rect -2348 38630 -2343 38652
rect -2325 38630 -2320 38652
rect -2000 38650 -1966 38652
rect -2309 38632 -2301 38640
rect -2062 38639 -2054 38646
rect -2092 38632 -2084 38639
rect -2062 38632 -2026 38634
rect -2317 38630 -2309 38632
rect -2062 38630 -2012 38632
rect -2000 38630 -1992 38650
rect -1982 38649 -1966 38650
rect -1846 38648 -1806 38652
rect -1846 38641 -1798 38646
rect -1806 38639 -1798 38641
rect -1854 38637 -1846 38639
rect -1854 38632 -1806 38637
rect -1655 38632 -1647 38640
rect -1864 38630 -1796 38631
rect -1663 38630 -1655 38632
rect -1642 38630 -1637 38652
rect -1619 38630 -1614 38652
rect -1530 38630 -1526 38652
rect -1506 38630 -1502 38652
rect -1482 38630 -1478 38652
rect -1458 38630 -1454 38652
rect -1434 38630 -1430 38652
rect -1410 38630 -1406 38652
rect -1386 38630 -1382 38652
rect -1362 38630 -1358 38652
rect -1338 38630 -1334 38652
rect -1314 38630 -1310 38652
rect -1290 38630 -1286 38652
rect -1266 38630 -1262 38652
rect -1242 38630 -1238 38652
rect -1235 38651 -1221 38652
rect -1218 38651 -1211 38675
rect -1218 38630 -1214 38651
rect -1194 38630 -1190 38676
rect -1170 38630 -1166 38676
rect -1146 38630 -1142 38676
rect -1122 38630 -1118 38676
rect -1098 38630 -1094 38676
rect -1074 38630 -1070 38676
rect -1050 38630 -1046 38676
rect -1026 38630 -1022 38676
rect -1002 38630 -998 38676
rect -978 38630 -974 38676
rect -954 38630 -950 38676
rect -930 38630 -926 38676
rect -906 38630 -902 38676
rect -882 38630 -878 38676
rect -858 38630 -854 38676
rect -834 38630 -830 38676
rect -810 38630 -806 38676
rect -786 38630 -782 38676
rect -762 38630 -758 38676
rect -738 38630 -734 38676
rect -714 38630 -710 38676
rect -690 38630 -686 38676
rect -666 38630 -662 38676
rect -642 38630 -638 38676
rect -618 38630 -614 38676
rect -594 38630 -590 38676
rect -570 38630 -566 38676
rect -546 38630 -542 38676
rect -522 38630 -518 38676
rect -498 38630 -494 38676
rect -474 38630 -470 38676
rect -450 38630 -446 38676
rect -426 38630 -422 38676
rect -402 38630 -398 38676
rect -378 38630 -374 38676
rect -354 38630 -350 38676
rect -330 38630 -326 38676
rect -306 38630 -302 38676
rect -282 38630 -278 38676
rect -258 38630 -254 38676
rect -234 38630 -230 38676
rect -210 38630 -206 38676
rect -203 38675 -189 38676
rect -186 38675 -179 38723
rect -186 38630 -182 38675
rect -162 38630 -158 38796
rect -138 38630 -134 38796
rect -114 38703 -110 38796
rect -125 38702 -91 38703
rect -90 38702 -86 38796
rect -66 38702 -62 38796
rect -42 38702 -38 38796
rect -18 38702 -14 38796
rect 6 38702 10 38796
rect 30 38702 34 38796
rect 54 38702 58 38796
rect 78 38702 82 38796
rect 102 38702 106 38796
rect 126 38702 130 38796
rect 150 38702 154 38796
rect 174 38702 178 38796
rect 198 38702 202 38796
rect 222 38702 226 38796
rect 246 38702 250 38796
rect 270 38702 274 38796
rect 294 38702 298 38796
rect 318 38702 322 38796
rect 342 38702 346 38796
rect 366 38702 370 38796
rect 390 38702 394 38796
rect 414 38702 418 38796
rect 438 38702 442 38796
rect 462 38702 466 38796
rect 486 38702 490 38796
rect 499 38717 504 38727
rect 510 38717 514 38796
rect 509 38703 514 38717
rect 510 38702 514 38703
rect 534 38702 538 38796
rect 558 38702 562 38796
rect 582 38702 586 38796
rect 606 38702 610 38796
rect 630 38702 634 38796
rect 654 38702 658 38796
rect 678 38702 682 38796
rect 702 38702 706 38796
rect 726 38702 730 38796
rect 750 38702 754 38796
rect 774 38702 778 38796
rect 798 38702 802 38796
rect 822 38702 826 38796
rect 846 38702 850 38796
rect 870 38702 874 38796
rect 894 38702 898 38796
rect 918 38702 922 38796
rect 925 38795 939 38796
rect 931 38789 936 38795
rect 941 38775 946 38789
rect 942 38702 946 38775
rect 955 38702 963 38703
rect -125 38700 963 38702
rect -125 38693 -120 38700
rect -114 38693 -110 38700
rect -115 38679 -110 38693
rect -125 38669 -120 38679
rect -115 38655 -110 38669
rect -114 38630 -110 38655
rect -90 38630 -86 38700
rect -66 38630 -62 38700
rect -42 38630 -38 38700
rect -18 38630 -14 38700
rect 6 38630 10 38700
rect 30 38630 34 38700
rect 54 38630 58 38700
rect 78 38630 82 38700
rect 102 38630 106 38700
rect 126 38630 130 38700
rect 150 38630 154 38700
rect 174 38630 178 38700
rect 198 38630 202 38700
rect 222 38630 226 38700
rect 246 38630 250 38700
rect 270 38630 274 38700
rect 294 38630 298 38700
rect 318 38630 322 38700
rect 342 38630 346 38700
rect 366 38630 370 38700
rect 390 38630 394 38700
rect 414 38630 418 38700
rect 438 38630 442 38700
rect 462 38630 466 38700
rect 486 38630 490 38700
rect 510 38630 514 38700
rect 523 38645 528 38655
rect 534 38651 538 38700
rect 534 38645 541 38651
rect 533 38631 541 38645
rect -2393 38628 531 38630
rect -2371 38582 -2366 38628
rect -2348 38582 -2343 38628
rect -2325 38582 -2320 38628
rect -2317 38624 -2309 38628
rect -2062 38624 -2054 38628
rect -2154 38620 -2138 38622
rect -2057 38620 -2054 38624
rect -2292 38614 -2054 38620
rect -2052 38614 -2044 38624
rect -2092 38598 -2062 38600
rect -2094 38594 -2062 38598
rect -2000 38582 -1992 38628
rect -1846 38621 -1806 38628
rect -1663 38624 -1655 38628
rect -1846 38614 -1680 38620
rect -1854 38598 -1806 38600
rect -1854 38594 -1680 38598
rect -1642 38582 -1637 38628
rect -1619 38582 -1614 38628
rect -1530 38582 -1526 38628
rect -1506 38582 -1502 38628
rect -1482 38582 -1478 38628
rect -1458 38582 -1454 38628
rect -1434 38582 -1430 38628
rect -1410 38582 -1406 38628
rect -1386 38582 -1382 38628
rect -1362 38582 -1358 38628
rect -1338 38582 -1334 38628
rect -1314 38582 -1310 38628
rect -1290 38582 -1286 38628
rect -1266 38582 -1262 38628
rect -1242 38582 -1238 38628
rect -1218 38582 -1214 38628
rect -1194 38582 -1190 38628
rect -1170 38582 -1166 38628
rect -1146 38582 -1142 38628
rect -1122 38582 -1118 38628
rect -1098 38582 -1094 38628
rect -1074 38582 -1070 38628
rect -1050 38582 -1046 38628
rect -1026 38582 -1022 38628
rect -1002 38582 -998 38628
rect -978 38582 -974 38628
rect -954 38582 -950 38628
rect -930 38582 -926 38628
rect -906 38582 -902 38628
rect -882 38582 -878 38628
rect -858 38582 -854 38628
rect -834 38582 -830 38628
rect -810 38582 -806 38628
rect -786 38582 -782 38628
rect -762 38582 -758 38628
rect -738 38582 -734 38628
rect -725 38597 -720 38607
rect -714 38597 -710 38628
rect -715 38583 -710 38597
rect -725 38582 -691 38583
rect -2393 38580 -691 38582
rect -2371 38558 -2366 38580
rect -2348 38558 -2343 38580
rect -2325 38558 -2320 38580
rect -2072 38578 -2036 38579
rect -2072 38572 -2054 38578
rect -2309 38564 -2301 38572
rect -2317 38558 -2309 38564
rect -2092 38563 -2062 38568
rect -2000 38559 -1992 38580
rect -1938 38579 -1906 38580
rect -1920 38578 -1906 38579
rect -1806 38572 -1680 38578
rect -1854 38563 -1806 38568
rect -1655 38564 -1647 38572
rect -1982 38559 -1966 38560
rect -2000 38558 -1966 38559
rect -1846 38558 -1806 38561
rect -1663 38558 -1655 38564
rect -1642 38558 -1637 38580
rect -1619 38558 -1614 38580
rect -1530 38558 -1526 38580
rect -1506 38558 -1502 38580
rect -1482 38558 -1478 38580
rect -1458 38558 -1454 38580
rect -1434 38558 -1430 38580
rect -1410 38558 -1406 38580
rect -1386 38558 -1382 38580
rect -1362 38558 -1358 38580
rect -1338 38558 -1334 38580
rect -1314 38558 -1310 38580
rect -1290 38558 -1286 38580
rect -1266 38558 -1262 38580
rect -1242 38558 -1238 38580
rect -1218 38558 -1214 38580
rect -1194 38558 -1190 38580
rect -1170 38558 -1166 38580
rect -1146 38558 -1142 38580
rect -1122 38558 -1118 38580
rect -1098 38558 -1094 38580
rect -1074 38558 -1070 38580
rect -1050 38558 -1046 38580
rect -1026 38558 -1022 38580
rect -1002 38558 -998 38580
rect -978 38558 -974 38580
rect -954 38558 -950 38580
rect -930 38559 -926 38580
rect -941 38558 -907 38559
rect -2393 38556 -907 38558
rect -2371 38534 -2366 38556
rect -2348 38534 -2343 38556
rect -2325 38534 -2320 38556
rect -2000 38554 -1966 38556
rect -2309 38536 -2301 38544
rect -2062 38543 -2054 38550
rect -2092 38536 -2084 38543
rect -2062 38536 -2026 38538
rect -2317 38534 -2309 38536
rect -2062 38534 -2012 38536
rect -2000 38534 -1992 38554
rect -1982 38553 -1966 38554
rect -1846 38552 -1806 38556
rect -1846 38545 -1798 38550
rect -1806 38543 -1798 38545
rect -1854 38541 -1846 38543
rect -1854 38536 -1806 38541
rect -1655 38536 -1647 38544
rect -1864 38534 -1796 38535
rect -1663 38534 -1655 38536
rect -1642 38534 -1637 38556
rect -1619 38534 -1614 38556
rect -1530 38534 -1526 38556
rect -1506 38534 -1502 38556
rect -1482 38534 -1478 38556
rect -1458 38534 -1454 38556
rect -1434 38534 -1430 38556
rect -1410 38534 -1406 38556
rect -1386 38534 -1382 38556
rect -1362 38534 -1358 38556
rect -1338 38534 -1334 38556
rect -1314 38534 -1310 38556
rect -1290 38534 -1286 38556
rect -1266 38534 -1262 38556
rect -1242 38534 -1238 38556
rect -1218 38534 -1214 38556
rect -1194 38534 -1190 38556
rect -1170 38534 -1166 38556
rect -1146 38534 -1142 38556
rect -1122 38534 -1118 38556
rect -1098 38534 -1094 38556
rect -1074 38534 -1070 38556
rect -1050 38534 -1046 38556
rect -1026 38534 -1022 38556
rect -1002 38534 -998 38556
rect -978 38534 -974 38556
rect -954 38534 -950 38556
rect -941 38549 -936 38556
rect -930 38549 -926 38556
rect -931 38535 -926 38549
rect -930 38534 -926 38535
rect -906 38534 -902 38580
rect -882 38534 -878 38580
rect -858 38534 -854 38580
rect -834 38534 -830 38580
rect -810 38534 -806 38580
rect -786 38534 -782 38580
rect -762 38534 -758 38580
rect -738 38534 -734 38580
rect -725 38573 -720 38580
rect -715 38559 -710 38573
rect -714 38534 -710 38559
rect -690 38534 -686 38628
rect -666 38534 -662 38628
rect -642 38534 -638 38628
rect -618 38534 -614 38628
rect -594 38534 -590 38628
rect -570 38534 -566 38628
rect -546 38534 -542 38628
rect -522 38534 -518 38628
rect -498 38534 -494 38628
rect -474 38534 -470 38628
rect -450 38534 -446 38628
rect -426 38534 -422 38628
rect -402 38534 -398 38628
rect -378 38534 -374 38628
rect -354 38534 -350 38628
rect -330 38534 -326 38628
rect -306 38534 -302 38628
rect -282 38534 -278 38628
rect -258 38534 -254 38628
rect -234 38534 -230 38628
rect -210 38534 -206 38628
rect -186 38534 -182 38628
rect -162 38534 -158 38628
rect -138 38534 -134 38628
rect -114 38534 -110 38628
rect -90 38627 -86 38628
rect -90 38606 -83 38627
rect -66 38606 -62 38628
rect -42 38606 -38 38628
rect -18 38606 -14 38628
rect 6 38606 10 38628
rect 30 38606 34 38628
rect 54 38606 58 38628
rect 78 38606 82 38628
rect 102 38606 106 38628
rect 126 38606 130 38628
rect 150 38606 154 38628
rect 174 38606 178 38628
rect 198 38606 202 38628
rect 222 38606 226 38628
rect 246 38606 250 38628
rect 270 38606 274 38628
rect 294 38606 298 38628
rect 318 38606 322 38628
rect 342 38606 346 38628
rect 366 38606 370 38628
rect 390 38606 394 38628
rect 414 38606 418 38628
rect 438 38606 442 38628
rect 462 38606 466 38628
rect 486 38606 490 38628
rect 510 38606 514 38628
rect 517 38627 531 38628
rect 534 38627 541 38631
rect 534 38606 538 38627
rect 558 38606 562 38700
rect 582 38606 586 38700
rect 606 38606 610 38700
rect 630 38606 634 38700
rect 654 38606 658 38700
rect 667 38621 672 38631
rect 678 38621 682 38700
rect 677 38607 682 38621
rect 678 38606 682 38607
rect 702 38606 706 38700
rect 726 38606 730 38700
rect 750 38606 754 38700
rect 774 38606 778 38700
rect 798 38606 802 38700
rect 822 38606 826 38700
rect 846 38606 850 38700
rect 870 38606 874 38700
rect 894 38606 898 38700
rect 918 38606 922 38700
rect 942 38606 946 38700
rect 949 38699 963 38700
rect 955 38693 960 38699
rect 965 38679 970 38693
rect 966 38606 970 38679
rect 979 38606 987 38607
rect -107 38604 987 38606
rect -107 38603 -93 38604
rect -90 38579 -83 38604
rect -90 38534 -86 38579
rect -66 38534 -62 38604
rect -42 38534 -38 38604
rect -18 38534 -14 38604
rect 6 38534 10 38604
rect 30 38534 34 38604
rect 54 38534 58 38604
rect 78 38534 82 38604
rect 102 38534 106 38604
rect 126 38534 130 38604
rect 150 38534 154 38604
rect 174 38534 178 38604
rect 198 38534 202 38604
rect 222 38534 226 38604
rect 246 38534 250 38604
rect 270 38534 274 38604
rect 294 38534 298 38604
rect 318 38534 322 38604
rect 342 38534 346 38604
rect 366 38534 370 38604
rect 390 38534 394 38604
rect 414 38534 418 38604
rect 438 38534 442 38604
rect 462 38534 466 38604
rect 486 38534 490 38604
rect 510 38534 514 38604
rect 534 38534 538 38604
rect 558 38579 562 38604
rect 558 38555 565 38579
rect 558 38534 562 38555
rect 582 38534 586 38604
rect 606 38534 610 38604
rect 630 38534 634 38604
rect 654 38534 658 38604
rect 678 38534 682 38604
rect 702 38555 706 38604
rect -2393 38532 699 38534
rect -2371 38486 -2366 38532
rect -2348 38486 -2343 38532
rect -2325 38486 -2320 38532
rect -2317 38528 -2309 38532
rect -2062 38528 -2054 38532
rect -2154 38524 -2138 38526
rect -2057 38524 -2054 38528
rect -2292 38518 -2054 38524
rect -2052 38518 -2044 38528
rect -2092 38502 -2062 38504
rect -2094 38498 -2062 38502
rect -2000 38486 -1992 38532
rect -1846 38525 -1806 38532
rect -1663 38528 -1655 38532
rect -1846 38518 -1680 38524
rect -1854 38502 -1806 38504
rect -1854 38498 -1680 38502
rect -1642 38486 -1637 38532
rect -1619 38486 -1614 38532
rect -1530 38486 -1526 38532
rect -1506 38486 -1502 38532
rect -1482 38486 -1478 38532
rect -1458 38486 -1454 38532
rect -1434 38486 -1430 38532
rect -1410 38486 -1406 38532
rect -1386 38486 -1382 38532
rect -1362 38486 -1358 38532
rect -1338 38486 -1334 38532
rect -1314 38486 -1310 38532
rect -1290 38486 -1286 38532
rect -1266 38486 -1262 38532
rect -1242 38486 -1238 38532
rect -1218 38486 -1214 38532
rect -1194 38486 -1190 38532
rect -1170 38486 -1166 38532
rect -1146 38486 -1142 38532
rect -1122 38486 -1118 38532
rect -1098 38486 -1094 38532
rect -1074 38486 -1070 38532
rect -1050 38486 -1046 38532
rect -1026 38486 -1022 38532
rect -1002 38486 -998 38532
rect -978 38486 -974 38532
rect -954 38486 -950 38532
rect -930 38486 -926 38532
rect -906 38486 -902 38532
rect -882 38486 -878 38532
rect -858 38486 -854 38532
rect -834 38486 -830 38532
rect -810 38486 -806 38532
rect -786 38486 -782 38532
rect -762 38486 -758 38532
rect -738 38486 -734 38532
rect -714 38486 -710 38532
rect -690 38531 -686 38532
rect -2393 38484 -693 38486
rect -2371 38462 -2366 38484
rect -2348 38462 -2343 38484
rect -2325 38462 -2320 38484
rect -2072 38482 -2036 38483
rect -2072 38476 -2054 38482
rect -2309 38468 -2301 38476
rect -2317 38462 -2309 38468
rect -2092 38467 -2062 38472
rect -2000 38463 -1992 38484
rect -1938 38483 -1906 38484
rect -1920 38482 -1906 38483
rect -1806 38476 -1680 38482
rect -1854 38467 -1806 38472
rect -1655 38468 -1647 38476
rect -1982 38463 -1966 38464
rect -2000 38462 -1966 38463
rect -1846 38462 -1806 38465
rect -1663 38462 -1655 38468
rect -1642 38462 -1637 38484
rect -1619 38462 -1614 38484
rect -1530 38462 -1526 38484
rect -1506 38462 -1502 38484
rect -1482 38462 -1478 38484
rect -1458 38462 -1454 38484
rect -1434 38462 -1430 38484
rect -1410 38462 -1406 38484
rect -1386 38462 -1382 38484
rect -1362 38462 -1358 38484
rect -1338 38462 -1334 38484
rect -1314 38462 -1310 38484
rect -1290 38462 -1286 38484
rect -1266 38462 -1262 38484
rect -1242 38462 -1238 38484
rect -1218 38462 -1214 38484
rect -1194 38462 -1190 38484
rect -1170 38462 -1166 38484
rect -1146 38462 -1142 38484
rect -1122 38462 -1118 38484
rect -1098 38462 -1094 38484
rect -1074 38462 -1070 38484
rect -1050 38462 -1046 38484
rect -1026 38462 -1022 38484
rect -1002 38462 -998 38484
rect -978 38462 -974 38484
rect -954 38462 -950 38484
rect -930 38462 -926 38484
rect -906 38483 -902 38484
rect -2393 38460 -909 38462
rect -2371 38438 -2366 38460
rect -2348 38438 -2343 38460
rect -2325 38438 -2320 38460
rect -2000 38458 -1966 38460
rect -2309 38440 -2301 38448
rect -2062 38447 -2054 38454
rect -2092 38440 -2084 38447
rect -2062 38440 -2026 38442
rect -2317 38438 -2309 38440
rect -2062 38438 -2012 38440
rect -2000 38438 -1992 38458
rect -1982 38457 -1966 38458
rect -1846 38456 -1806 38460
rect -1846 38449 -1798 38454
rect -1806 38447 -1798 38449
rect -1854 38445 -1846 38447
rect -1854 38440 -1806 38445
rect -1655 38440 -1647 38448
rect -1864 38438 -1796 38439
rect -1663 38438 -1655 38440
rect -1642 38438 -1637 38460
rect -1619 38438 -1614 38460
rect -1530 38438 -1526 38460
rect -1506 38438 -1502 38460
rect -1482 38438 -1478 38460
rect -1458 38438 -1454 38460
rect -1434 38438 -1430 38460
rect -1410 38438 -1406 38460
rect -1386 38438 -1382 38460
rect -1362 38438 -1358 38460
rect -1338 38438 -1334 38460
rect -1314 38438 -1310 38460
rect -1290 38438 -1286 38460
rect -1266 38438 -1262 38460
rect -1242 38438 -1238 38460
rect -1218 38438 -1214 38460
rect -1194 38438 -1190 38460
rect -1170 38438 -1166 38460
rect -1146 38438 -1142 38460
rect -1122 38438 -1118 38460
rect -1098 38438 -1094 38460
rect -1074 38438 -1070 38460
rect -1050 38438 -1046 38460
rect -1026 38438 -1022 38460
rect -1002 38438 -998 38460
rect -978 38438 -974 38460
rect -954 38438 -950 38460
rect -930 38438 -926 38460
rect -923 38459 -909 38460
rect -906 38459 -899 38483
rect -906 38438 -902 38459
rect -882 38438 -878 38484
rect -858 38438 -854 38484
rect -834 38438 -830 38484
rect -810 38438 -806 38484
rect -786 38438 -782 38484
rect -773 38453 -768 38463
rect -762 38453 -758 38484
rect -763 38439 -758 38453
rect -762 38438 -758 38439
rect -738 38438 -734 38484
rect -714 38438 -710 38484
rect -707 38483 -693 38484
rect -690 38483 -683 38531
rect -690 38438 -686 38483
rect -666 38438 -662 38532
rect -642 38438 -638 38532
rect -618 38438 -614 38532
rect -594 38438 -590 38532
rect -570 38438 -566 38532
rect -546 38438 -542 38532
rect -522 38438 -518 38532
rect -498 38438 -494 38532
rect -474 38438 -470 38532
rect -450 38438 -446 38532
rect -426 38438 -422 38532
rect -402 38438 -398 38532
rect -378 38438 -374 38532
rect -354 38438 -350 38532
rect -330 38438 -326 38532
rect -306 38438 -302 38532
rect -282 38438 -278 38532
rect -258 38438 -254 38532
rect -234 38438 -230 38532
rect -210 38438 -206 38532
rect -186 38438 -182 38532
rect -162 38438 -158 38532
rect -138 38438 -134 38532
rect -114 38438 -110 38532
rect -90 38438 -86 38532
rect -66 38438 -62 38532
rect -42 38438 -38 38532
rect -18 38438 -14 38532
rect 6 38438 10 38532
rect 30 38438 34 38532
rect 54 38438 58 38532
rect 78 38438 82 38532
rect 102 38438 106 38532
rect 126 38438 130 38532
rect 150 38439 154 38532
rect 139 38438 173 38439
rect -2393 38436 173 38438
rect -2371 38390 -2366 38436
rect -2348 38390 -2343 38436
rect -2325 38390 -2320 38436
rect -2317 38432 -2309 38436
rect -2062 38432 -2054 38436
rect -2154 38428 -2138 38430
rect -2057 38428 -2054 38432
rect -2292 38422 -2054 38428
rect -2052 38422 -2044 38432
rect -2092 38406 -2062 38408
rect -2094 38402 -2062 38406
rect -2000 38390 -1992 38436
rect -1846 38429 -1806 38436
rect -1663 38432 -1655 38436
rect -1846 38422 -1680 38428
rect -1854 38406 -1806 38408
rect -1854 38402 -1680 38406
rect -1642 38390 -1637 38436
rect -1619 38390 -1614 38436
rect -1530 38390 -1526 38436
rect -1506 38390 -1502 38436
rect -1482 38390 -1478 38436
rect -1458 38390 -1454 38436
rect -1434 38390 -1430 38436
rect -1410 38390 -1406 38436
rect -1386 38390 -1382 38436
rect -1362 38390 -1358 38436
rect -1338 38390 -1334 38436
rect -1314 38390 -1310 38436
rect -1290 38390 -1286 38436
rect -1266 38390 -1262 38436
rect -1242 38390 -1238 38436
rect -1218 38390 -1214 38436
rect -1194 38390 -1190 38436
rect -1170 38390 -1166 38436
rect -1146 38390 -1142 38436
rect -1122 38390 -1118 38436
rect -1098 38390 -1094 38436
rect -1074 38390 -1070 38436
rect -1050 38390 -1046 38436
rect -1026 38390 -1022 38436
rect -1002 38390 -998 38436
rect -978 38390 -974 38436
rect -954 38390 -950 38436
rect -930 38390 -926 38436
rect -906 38390 -902 38436
rect -882 38390 -878 38436
rect -858 38390 -854 38436
rect -834 38390 -830 38436
rect -810 38390 -806 38436
rect -786 38390 -782 38436
rect -762 38390 -758 38436
rect -738 38390 -734 38436
rect -714 38390 -710 38436
rect -690 38390 -686 38436
rect -666 38390 -662 38436
rect -642 38390 -638 38436
rect -618 38390 -614 38436
rect -594 38390 -590 38436
rect -570 38390 -566 38436
rect -546 38390 -542 38436
rect -522 38390 -518 38436
rect -498 38390 -494 38436
rect -474 38390 -470 38436
rect -450 38390 -446 38436
rect -426 38390 -422 38436
rect -402 38390 -398 38436
rect -378 38390 -374 38436
rect -354 38390 -350 38436
rect -330 38390 -326 38436
rect -306 38390 -302 38436
rect -282 38390 -278 38436
rect -258 38390 -254 38436
rect -234 38390 -230 38436
rect -210 38390 -206 38436
rect -186 38390 -182 38436
rect -162 38390 -158 38436
rect -138 38390 -134 38436
rect -114 38390 -110 38436
rect -90 38390 -86 38436
rect -66 38390 -62 38436
rect -42 38390 -38 38436
rect -18 38390 -14 38436
rect 6 38390 10 38436
rect 30 38390 34 38436
rect 54 38390 58 38436
rect 78 38390 82 38436
rect 102 38390 106 38436
rect 126 38390 130 38436
rect 139 38429 144 38436
rect 150 38429 154 38436
rect 149 38415 154 38429
rect 150 38390 154 38415
rect 174 38390 178 38532
rect 198 38390 202 38532
rect 222 38390 226 38532
rect 246 38390 250 38532
rect 270 38390 274 38532
rect 294 38390 298 38532
rect 318 38390 322 38532
rect 331 38405 336 38415
rect 342 38405 346 38532
rect 341 38391 346 38405
rect 331 38390 365 38391
rect -2393 38388 365 38390
rect -2371 38366 -2366 38388
rect -2348 38366 -2343 38388
rect -2325 38366 -2320 38388
rect -2072 38386 -2036 38387
rect -2072 38380 -2054 38386
rect -2309 38372 -2301 38380
rect -2317 38366 -2309 38372
rect -2092 38371 -2062 38376
rect -2000 38367 -1992 38388
rect -1938 38387 -1906 38388
rect -1920 38386 -1906 38387
rect -1806 38380 -1680 38386
rect -1854 38371 -1806 38376
rect -1655 38372 -1647 38380
rect -1982 38367 -1966 38368
rect -2000 38366 -1966 38367
rect -1846 38366 -1806 38369
rect -1663 38366 -1655 38372
rect -1642 38366 -1637 38388
rect -1619 38366 -1614 38388
rect -1530 38366 -1526 38388
rect -1506 38366 -1502 38388
rect -1482 38366 -1478 38388
rect -1458 38366 -1454 38388
rect -1434 38366 -1430 38388
rect -1410 38366 -1406 38388
rect -1386 38366 -1382 38388
rect -1362 38366 -1358 38388
rect -1338 38366 -1334 38388
rect -1314 38366 -1310 38388
rect -1290 38366 -1286 38388
rect -1266 38366 -1262 38388
rect -1242 38366 -1238 38388
rect -1218 38366 -1214 38388
rect -1194 38366 -1190 38388
rect -1170 38366 -1166 38388
rect -1146 38366 -1142 38388
rect -1122 38366 -1118 38388
rect -1098 38366 -1094 38388
rect -1074 38366 -1070 38388
rect -1050 38366 -1046 38388
rect -1026 38366 -1022 38388
rect -1002 38366 -998 38388
rect -978 38366 -974 38388
rect -954 38366 -950 38388
rect -930 38366 -926 38388
rect -906 38366 -902 38388
rect -882 38366 -878 38388
rect -858 38366 -854 38388
rect -834 38366 -830 38388
rect -810 38366 -806 38388
rect -786 38366 -782 38388
rect -762 38366 -758 38388
rect -738 38387 -734 38388
rect -2393 38364 -741 38366
rect -2371 38342 -2366 38364
rect -2348 38342 -2343 38364
rect -2325 38342 -2320 38364
rect -2000 38362 -1966 38364
rect -2309 38344 -2301 38352
rect -2062 38351 -2054 38358
rect -2092 38344 -2084 38351
rect -2062 38344 -2026 38346
rect -2317 38342 -2309 38344
rect -2062 38342 -2012 38344
rect -2000 38342 -1992 38362
rect -1982 38361 -1966 38362
rect -1846 38360 -1806 38364
rect -1846 38353 -1798 38358
rect -1806 38351 -1798 38353
rect -1854 38349 -1846 38351
rect -1854 38344 -1806 38349
rect -1655 38344 -1647 38352
rect -1864 38342 -1796 38343
rect -1663 38342 -1655 38344
rect -1642 38342 -1637 38364
rect -1619 38342 -1614 38364
rect -1530 38342 -1526 38364
rect -1506 38342 -1502 38364
rect -1482 38342 -1478 38364
rect -1458 38342 -1454 38364
rect -1434 38342 -1430 38364
rect -1410 38342 -1406 38364
rect -1386 38342 -1382 38364
rect -1362 38342 -1358 38364
rect -1338 38342 -1334 38364
rect -1314 38342 -1310 38364
rect -1290 38342 -1286 38364
rect -1266 38342 -1262 38364
rect -1242 38342 -1238 38364
rect -1218 38342 -1214 38364
rect -1194 38342 -1190 38364
rect -1170 38342 -1166 38364
rect -1146 38342 -1142 38364
rect -1122 38342 -1118 38364
rect -1098 38342 -1094 38364
rect -1074 38342 -1070 38364
rect -1050 38342 -1046 38364
rect -1026 38342 -1022 38364
rect -1002 38342 -998 38364
rect -978 38342 -974 38364
rect -954 38342 -950 38364
rect -930 38342 -926 38364
rect -906 38342 -902 38364
rect -882 38342 -878 38364
rect -858 38342 -854 38364
rect -834 38342 -830 38364
rect -810 38342 -806 38364
rect -786 38342 -782 38364
rect -762 38342 -758 38364
rect -755 38363 -741 38364
rect -738 38363 -731 38387
rect -738 38342 -734 38363
rect -714 38342 -710 38388
rect -690 38342 -686 38388
rect -666 38342 -662 38388
rect -642 38342 -638 38388
rect -618 38342 -614 38388
rect -594 38342 -590 38388
rect -570 38342 -566 38388
rect -546 38342 -542 38388
rect -522 38342 -518 38388
rect -498 38342 -494 38388
rect -474 38342 -470 38388
rect -450 38342 -446 38388
rect -426 38342 -422 38388
rect -402 38342 -398 38388
rect -378 38342 -374 38388
rect -354 38342 -350 38388
rect -330 38342 -326 38388
rect -306 38342 -302 38388
rect -282 38342 -278 38388
rect -258 38342 -254 38388
rect -234 38342 -230 38388
rect -210 38342 -206 38388
rect -186 38342 -182 38388
rect -162 38342 -158 38388
rect -138 38342 -134 38388
rect -114 38342 -110 38388
rect -90 38342 -86 38388
rect -66 38342 -62 38388
rect -42 38342 -38 38388
rect -18 38342 -14 38388
rect 6 38342 10 38388
rect 30 38342 34 38388
rect 54 38342 58 38388
rect 78 38342 82 38388
rect 102 38342 106 38388
rect 115 38357 120 38367
rect 126 38357 130 38388
rect 125 38343 130 38357
rect 126 38342 130 38343
rect 150 38342 154 38388
rect 174 38363 178 38388
rect -2393 38340 171 38342
rect -2371 38294 -2366 38340
rect -2348 38294 -2343 38340
rect -2325 38294 -2320 38340
rect -2317 38336 -2309 38340
rect -2062 38336 -2054 38340
rect -2154 38332 -2138 38334
rect -2057 38332 -2054 38336
rect -2292 38326 -2054 38332
rect -2052 38326 -2044 38336
rect -2092 38310 -2062 38312
rect -2094 38306 -2062 38310
rect -2000 38294 -1992 38340
rect -1846 38333 -1806 38340
rect -1663 38336 -1655 38340
rect -1846 38326 -1680 38332
rect -1854 38310 -1806 38312
rect -1854 38306 -1680 38310
rect -1642 38294 -1637 38340
rect -1619 38294 -1614 38340
rect -1530 38294 -1526 38340
rect -1506 38294 -1502 38340
rect -1482 38294 -1478 38340
rect -1458 38294 -1454 38340
rect -1434 38294 -1430 38340
rect -1410 38294 -1406 38340
rect -1386 38294 -1382 38340
rect -1362 38294 -1358 38340
rect -1338 38294 -1334 38340
rect -1314 38294 -1310 38340
rect -1290 38294 -1286 38340
rect -1266 38294 -1262 38340
rect -1242 38294 -1238 38340
rect -1218 38294 -1214 38340
rect -1194 38294 -1190 38340
rect -1170 38294 -1166 38340
rect -1146 38294 -1142 38340
rect -1122 38294 -1118 38340
rect -1098 38294 -1094 38340
rect -1074 38294 -1070 38340
rect -1050 38294 -1046 38340
rect -1026 38294 -1022 38340
rect -1002 38294 -998 38340
rect -978 38294 -974 38340
rect -954 38294 -950 38340
rect -930 38294 -926 38340
rect -906 38294 -902 38340
rect -882 38294 -878 38340
rect -869 38309 -864 38319
rect -858 38309 -854 38340
rect -859 38295 -854 38309
rect -869 38294 -835 38295
rect -2393 38292 -835 38294
rect -2371 38270 -2366 38292
rect -2348 38270 -2343 38292
rect -2325 38270 -2320 38292
rect -2072 38290 -2036 38291
rect -2072 38284 -2054 38290
rect -2309 38276 -2301 38284
rect -2317 38270 -2309 38276
rect -2092 38275 -2062 38280
rect -2000 38271 -1992 38292
rect -1938 38291 -1906 38292
rect -1920 38290 -1906 38291
rect -1806 38284 -1680 38290
rect -1854 38275 -1806 38280
rect -1655 38276 -1647 38284
rect -1982 38271 -1966 38272
rect -2000 38270 -1966 38271
rect -1846 38270 -1806 38273
rect -1663 38270 -1655 38276
rect -1642 38270 -1637 38292
rect -1619 38270 -1614 38292
rect -1530 38270 -1526 38292
rect -1506 38270 -1502 38292
rect -1482 38270 -1478 38292
rect -1458 38270 -1454 38292
rect -1434 38270 -1430 38292
rect -1410 38270 -1406 38292
rect -1386 38270 -1382 38292
rect -1362 38270 -1358 38292
rect -1338 38270 -1334 38292
rect -1314 38270 -1310 38292
rect -1290 38270 -1286 38292
rect -1266 38270 -1262 38292
rect -1242 38270 -1238 38292
rect -1218 38270 -1214 38292
rect -1194 38270 -1190 38292
rect -1170 38270 -1166 38292
rect -1146 38270 -1142 38292
rect -1122 38270 -1118 38292
rect -1098 38270 -1094 38292
rect -1074 38270 -1070 38292
rect -1050 38270 -1046 38292
rect -1026 38270 -1022 38292
rect -1002 38270 -998 38292
rect -978 38270 -974 38292
rect -954 38270 -950 38292
rect -930 38270 -926 38292
rect -906 38270 -902 38292
rect -882 38270 -878 38292
rect -869 38285 -864 38292
rect -859 38271 -854 38285
rect -858 38270 -854 38271
rect -834 38270 -830 38340
rect -810 38270 -806 38340
rect -786 38270 -782 38340
rect -762 38270 -758 38340
rect -738 38270 -734 38340
rect -714 38270 -710 38340
rect -690 38270 -686 38340
rect -666 38270 -662 38340
rect -642 38270 -638 38340
rect -618 38270 -614 38340
rect -594 38270 -590 38340
rect -570 38270 -566 38340
rect -546 38270 -542 38340
rect -522 38270 -518 38340
rect -498 38270 -494 38340
rect -474 38270 -470 38340
rect -450 38270 -446 38340
rect -426 38270 -422 38340
rect -402 38270 -398 38340
rect -378 38270 -374 38340
rect -354 38270 -350 38340
rect -330 38270 -326 38340
rect -306 38270 -302 38340
rect -282 38270 -278 38340
rect -258 38270 -254 38340
rect -234 38270 -230 38340
rect -210 38270 -206 38340
rect -186 38270 -182 38340
rect -162 38270 -158 38340
rect -138 38270 -134 38340
rect -114 38270 -110 38340
rect -90 38270 -86 38340
rect -66 38270 -62 38340
rect -42 38270 -38 38340
rect -18 38270 -14 38340
rect 6 38270 10 38340
rect 30 38270 34 38340
rect 54 38270 58 38340
rect 78 38270 82 38340
rect 102 38270 106 38340
rect 126 38271 130 38340
rect 150 38291 154 38340
rect 157 38339 171 38340
rect 174 38339 181 38363
rect 115 38270 147 38271
rect -2393 38268 147 38270
rect -2371 38246 -2366 38268
rect -2348 38246 -2343 38268
rect -2325 38246 -2320 38268
rect -2000 38266 -1966 38268
rect -2309 38248 -2301 38256
rect -2062 38255 -2054 38262
rect -2092 38248 -2084 38255
rect -2062 38248 -2026 38250
rect -2317 38246 -2309 38248
rect -2062 38246 -2012 38248
rect -2000 38246 -1992 38266
rect -1982 38265 -1966 38266
rect -1846 38264 -1806 38268
rect -1846 38257 -1798 38262
rect -1806 38255 -1798 38257
rect -1854 38253 -1846 38255
rect -1854 38248 -1806 38253
rect -1655 38248 -1647 38256
rect -1864 38246 -1796 38247
rect -1663 38246 -1655 38248
rect -1642 38246 -1637 38268
rect -1619 38246 -1614 38268
rect -1530 38246 -1526 38268
rect -1506 38246 -1502 38268
rect -1482 38246 -1478 38268
rect -1458 38246 -1454 38268
rect -1434 38246 -1430 38268
rect -1410 38246 -1406 38268
rect -1386 38246 -1382 38268
rect -1362 38246 -1358 38268
rect -1338 38246 -1334 38268
rect -1314 38247 -1310 38268
rect -1325 38246 -1291 38247
rect -2393 38244 -1291 38246
rect -2371 38198 -2366 38244
rect -2348 38198 -2343 38244
rect -2325 38198 -2320 38244
rect -2317 38240 -2309 38244
rect -2062 38240 -2054 38244
rect -2154 38236 -2138 38238
rect -2057 38236 -2054 38240
rect -2292 38230 -2054 38236
rect -2052 38230 -2044 38240
rect -2092 38214 -2062 38216
rect -2094 38210 -2062 38214
rect -2000 38198 -1992 38244
rect -1846 38237 -1806 38244
rect -1663 38240 -1655 38244
rect -1846 38230 -1680 38236
rect -1854 38214 -1806 38216
rect -1854 38210 -1680 38214
rect -1642 38198 -1637 38244
rect -1619 38198 -1614 38244
rect -1530 38198 -1526 38244
rect -1506 38198 -1502 38244
rect -1482 38198 -1478 38244
rect -1458 38198 -1454 38244
rect -1434 38198 -1430 38244
rect -1410 38198 -1406 38244
rect -1386 38198 -1382 38244
rect -1362 38198 -1358 38244
rect -1338 38198 -1334 38244
rect -1325 38237 -1320 38244
rect -1314 38237 -1310 38244
rect -1315 38223 -1310 38237
rect -1314 38198 -1310 38223
rect -1290 38198 -1286 38268
rect -1266 38198 -1262 38268
rect -1242 38198 -1238 38268
rect -1218 38198 -1214 38268
rect -1194 38198 -1190 38268
rect -1170 38198 -1166 38268
rect -1146 38198 -1142 38268
rect -1122 38198 -1118 38268
rect -1098 38198 -1094 38268
rect -1074 38198 -1070 38268
rect -1050 38198 -1046 38268
rect -1026 38198 -1022 38268
rect -1002 38198 -998 38268
rect -978 38198 -974 38268
rect -954 38198 -950 38268
rect -930 38198 -926 38268
rect -906 38198 -902 38268
rect -882 38198 -878 38268
rect -858 38198 -854 38268
rect -834 38243 -830 38268
rect -2393 38196 -837 38198
rect -2371 38174 -2366 38196
rect -2348 38174 -2343 38196
rect -2325 38174 -2320 38196
rect -2072 38194 -2036 38195
rect -2072 38188 -2054 38194
rect -2309 38180 -2301 38188
rect -2317 38174 -2309 38180
rect -2092 38179 -2062 38184
rect -2000 38175 -1992 38196
rect -1938 38195 -1906 38196
rect -1920 38194 -1906 38195
rect -1806 38188 -1680 38194
rect -1854 38179 -1806 38184
rect -1655 38180 -1647 38188
rect -1982 38175 -1966 38176
rect -2000 38174 -1966 38175
rect -1846 38174 -1806 38177
rect -1663 38174 -1655 38180
rect -1642 38174 -1637 38196
rect -1619 38174 -1614 38196
rect -1530 38174 -1526 38196
rect -1506 38174 -1502 38196
rect -1482 38174 -1478 38196
rect -1458 38174 -1454 38196
rect -1434 38174 -1430 38196
rect -1410 38174 -1406 38196
rect -1386 38174 -1382 38196
rect -1362 38174 -1358 38196
rect -1338 38174 -1334 38196
rect -1314 38174 -1310 38196
rect -1290 38174 -1286 38196
rect -1266 38174 -1262 38196
rect -1242 38174 -1238 38196
rect -1218 38174 -1214 38196
rect -1194 38174 -1190 38196
rect -1170 38174 -1166 38196
rect -1146 38174 -1142 38196
rect -1122 38174 -1118 38196
rect -1098 38174 -1094 38196
rect -1074 38174 -1070 38196
rect -1050 38174 -1046 38196
rect -1026 38174 -1022 38196
rect -1002 38174 -998 38196
rect -978 38174 -974 38196
rect -954 38174 -950 38196
rect -930 38174 -926 38196
rect -906 38174 -902 38196
rect -882 38174 -878 38196
rect -858 38174 -854 38196
rect -851 38195 -837 38196
rect -834 38195 -827 38243
rect -834 38174 -830 38195
rect -810 38174 -806 38268
rect -786 38174 -782 38268
rect -762 38174 -758 38268
rect -738 38174 -734 38268
rect -714 38174 -710 38268
rect -690 38174 -686 38268
rect -666 38174 -662 38268
rect -642 38174 -638 38268
rect -618 38174 -614 38268
rect -594 38174 -590 38268
rect -570 38174 -566 38268
rect -546 38174 -542 38268
rect -522 38174 -518 38268
rect -498 38174 -494 38268
rect -474 38174 -470 38268
rect -450 38174 -446 38268
rect -426 38174 -422 38268
rect -402 38174 -398 38268
rect -378 38174 -374 38268
rect -354 38174 -350 38268
rect -330 38174 -326 38268
rect -306 38174 -302 38268
rect -282 38223 -278 38268
rect -293 38222 -259 38223
rect -258 38222 -254 38268
rect -234 38222 -230 38268
rect -210 38222 -206 38268
rect -186 38222 -182 38268
rect -162 38222 -158 38268
rect -138 38222 -134 38268
rect -114 38222 -110 38268
rect -90 38222 -86 38268
rect -66 38222 -62 38268
rect -42 38222 -38 38268
rect -18 38222 -14 38268
rect 6 38222 10 38268
rect 30 38222 34 38268
rect 54 38222 58 38268
rect 78 38222 82 38268
rect 102 38222 106 38268
rect 115 38261 120 38268
rect 126 38261 130 38268
rect 133 38267 147 38268
rect 150 38267 157 38291
rect 125 38247 130 38261
rect 126 38222 130 38247
rect 150 38222 154 38267
rect 174 38222 178 38339
rect 198 38222 202 38388
rect 222 38222 226 38388
rect 246 38222 250 38388
rect 270 38222 274 38388
rect 294 38222 298 38388
rect 318 38222 322 38388
rect 331 38381 336 38388
rect 341 38367 346 38381
rect 342 38222 346 38367
rect 366 38339 370 38532
rect 366 38318 373 38339
rect 390 38318 394 38532
rect 414 38318 418 38532
rect 438 38318 442 38532
rect 462 38318 466 38532
rect 486 38318 490 38532
rect 510 38318 514 38532
rect 534 38318 538 38532
rect 558 38318 562 38532
rect 582 38318 586 38532
rect 606 38511 610 38532
rect 595 38510 629 38511
rect 630 38510 634 38532
rect 654 38510 658 38532
rect 678 38510 682 38532
rect 685 38531 699 38532
rect 702 38531 709 38555
rect 702 38510 706 38531
rect 726 38510 730 38604
rect 739 38525 744 38535
rect 750 38525 754 38604
rect 749 38511 754 38525
rect 750 38510 754 38511
rect 774 38510 778 38604
rect 798 38510 802 38604
rect 822 38510 826 38604
rect 846 38510 850 38604
rect 870 38510 874 38604
rect 894 38510 898 38604
rect 918 38510 922 38604
rect 942 38510 946 38604
rect 966 38510 970 38604
rect 973 38603 987 38604
rect 979 38597 984 38603
rect 989 38583 994 38597
rect 990 38510 994 38583
rect 1003 38510 1011 38511
rect 595 38508 1011 38510
rect 595 38501 600 38508
rect 606 38501 610 38508
rect 605 38487 610 38501
rect 595 38477 600 38487
rect 605 38463 610 38477
rect 606 38318 610 38463
rect 630 38435 634 38508
rect 630 38414 637 38435
rect 654 38414 658 38508
rect 678 38414 682 38508
rect 702 38414 706 38508
rect 726 38414 730 38508
rect 750 38414 754 38508
rect 774 38459 778 38508
rect 774 38435 781 38459
rect 774 38414 778 38435
rect 798 38414 802 38508
rect 822 38414 826 38508
rect 846 38414 850 38508
rect 870 38414 874 38508
rect 894 38414 898 38508
rect 918 38414 922 38508
rect 942 38414 946 38508
rect 966 38414 970 38508
rect 990 38414 994 38508
rect 997 38507 1011 38508
rect 1003 38501 1008 38507
rect 1013 38487 1018 38501
rect 1014 38414 1018 38487
rect 1027 38414 1035 38415
rect 613 38412 1035 38414
rect 613 38411 627 38412
rect 630 38387 637 38412
rect 630 38318 634 38387
rect 654 38318 658 38412
rect 678 38318 682 38412
rect 702 38318 706 38412
rect 726 38318 730 38412
rect 750 38318 754 38412
rect 774 38318 778 38412
rect 798 38318 802 38412
rect 822 38318 826 38412
rect 846 38318 850 38412
rect 870 38318 874 38412
rect 894 38318 898 38412
rect 918 38318 922 38412
rect 942 38318 946 38412
rect 966 38318 970 38412
rect 990 38318 994 38412
rect 1014 38318 1018 38412
rect 1021 38411 1035 38412
rect 1027 38405 1032 38411
rect 1037 38391 1042 38405
rect 1027 38333 1032 38343
rect 1038 38333 1042 38391
rect 1037 38319 1042 38333
rect 1051 38329 1059 38333
rect 1045 38319 1051 38329
rect 1027 38318 1059 38319
rect 349 38316 1059 38318
rect 349 38315 363 38316
rect 366 38291 373 38316
rect 366 38222 370 38291
rect 390 38222 394 38316
rect 414 38222 418 38316
rect 438 38222 442 38316
rect 462 38222 466 38316
rect 486 38222 490 38316
rect 510 38222 514 38316
rect 534 38222 538 38316
rect 558 38222 562 38316
rect 582 38222 586 38316
rect 606 38222 610 38316
rect 630 38222 634 38316
rect 654 38222 658 38316
rect 678 38222 682 38316
rect 702 38222 706 38316
rect 726 38222 730 38316
rect 750 38222 754 38316
rect 774 38222 778 38316
rect 798 38222 802 38316
rect 822 38222 826 38316
rect 846 38222 850 38316
rect 870 38222 874 38316
rect 894 38222 898 38316
rect 918 38222 922 38316
rect 942 38222 946 38316
rect 966 38222 970 38316
rect 990 38222 994 38316
rect 1014 38222 1018 38316
rect 1027 38309 1032 38316
rect 1045 38315 1059 38316
rect 1037 38295 1042 38309
rect 1038 38222 1042 38295
rect 1051 38222 1059 38223
rect -293 38220 1059 38222
rect -293 38213 -288 38220
rect -282 38213 -278 38220
rect -283 38199 -278 38213
rect -293 38189 -288 38199
rect -283 38175 -278 38189
rect -282 38174 -278 38175
rect -258 38174 -254 38220
rect -234 38174 -230 38220
rect -210 38174 -206 38220
rect -186 38174 -182 38220
rect -162 38174 -158 38220
rect -138 38174 -134 38220
rect -114 38174 -110 38220
rect -90 38174 -86 38220
rect -66 38174 -62 38220
rect -42 38175 -38 38220
rect -53 38174 -19 38175
rect -2393 38172 -19 38174
rect -2371 38150 -2366 38172
rect -2348 38150 -2343 38172
rect -2325 38150 -2320 38172
rect -2000 38170 -1966 38172
rect -2309 38152 -2301 38160
rect -2062 38159 -2054 38166
rect -2092 38152 -2084 38159
rect -2062 38152 -2026 38154
rect -2317 38150 -2309 38152
rect -2062 38150 -2012 38152
rect -2000 38150 -1992 38170
rect -1982 38169 -1966 38170
rect -1846 38168 -1806 38172
rect -1846 38161 -1798 38166
rect -1806 38159 -1798 38161
rect -1854 38157 -1846 38159
rect -1854 38152 -1806 38157
rect -1655 38152 -1647 38160
rect -1864 38150 -1796 38151
rect -1663 38150 -1655 38152
rect -1642 38150 -1637 38172
rect -1619 38150 -1614 38172
rect -1530 38150 -1526 38172
rect -1506 38150 -1502 38172
rect -1482 38150 -1478 38172
rect -1458 38150 -1454 38172
rect -1434 38150 -1430 38172
rect -1410 38150 -1406 38172
rect -1386 38150 -1382 38172
rect -1362 38150 -1358 38172
rect -1338 38150 -1334 38172
rect -1314 38150 -1310 38172
rect -1290 38171 -1286 38172
rect -2393 38148 -1293 38150
rect -2371 38102 -2366 38148
rect -2348 38102 -2343 38148
rect -2325 38102 -2320 38148
rect -2317 38144 -2309 38148
rect -2062 38144 -2054 38148
rect -2154 38140 -2138 38142
rect -2057 38140 -2054 38144
rect -2292 38134 -2054 38140
rect -2052 38134 -2044 38144
rect -2092 38118 -2062 38120
rect -2094 38114 -2062 38118
rect -2000 38102 -1992 38148
rect -1846 38141 -1806 38148
rect -1663 38144 -1655 38148
rect -1846 38134 -1680 38140
rect -1854 38118 -1806 38120
rect -1854 38114 -1680 38118
rect -1642 38102 -1637 38148
rect -1619 38102 -1614 38148
rect -1530 38102 -1526 38148
rect -1506 38102 -1502 38148
rect -1482 38102 -1478 38148
rect -1458 38102 -1454 38148
rect -1434 38102 -1430 38148
rect -1410 38102 -1406 38148
rect -1386 38102 -1382 38148
rect -1362 38102 -1358 38148
rect -1338 38102 -1334 38148
rect -1314 38102 -1310 38148
rect -1307 38147 -1293 38148
rect -1290 38147 -1283 38171
rect -1290 38102 -1286 38147
rect -1266 38102 -1262 38172
rect -1242 38102 -1238 38172
rect -1218 38102 -1214 38172
rect -1194 38102 -1190 38172
rect -1170 38102 -1166 38172
rect -1146 38102 -1142 38172
rect -1122 38102 -1118 38172
rect -1098 38102 -1094 38172
rect -1074 38102 -1070 38172
rect -1050 38102 -1046 38172
rect -1026 38102 -1022 38172
rect -1002 38102 -998 38172
rect -978 38102 -974 38172
rect -954 38102 -950 38172
rect -930 38102 -926 38172
rect -906 38102 -902 38172
rect -882 38102 -878 38172
rect -858 38102 -854 38172
rect -834 38102 -830 38172
rect -810 38102 -806 38172
rect -786 38102 -782 38172
rect -762 38102 -758 38172
rect -738 38102 -734 38172
rect -714 38102 -710 38172
rect -690 38102 -686 38172
rect -666 38102 -662 38172
rect -642 38102 -638 38172
rect -618 38102 -614 38172
rect -594 38102 -590 38172
rect -570 38102 -566 38172
rect -546 38102 -542 38172
rect -522 38102 -518 38172
rect -498 38102 -494 38172
rect -474 38102 -470 38172
rect -450 38102 -446 38172
rect -426 38102 -422 38172
rect -402 38102 -398 38172
rect -378 38102 -374 38172
rect -354 38102 -350 38172
rect -330 38102 -326 38172
rect -306 38102 -302 38172
rect -282 38102 -278 38172
rect -269 38141 -264 38151
rect -258 38147 -254 38172
rect -258 38141 -251 38147
rect -259 38127 -251 38141
rect -2393 38100 -261 38102
rect -2371 38078 -2366 38100
rect -2348 38078 -2343 38100
rect -2325 38078 -2320 38100
rect -2072 38098 -2036 38099
rect -2072 38092 -2054 38098
rect -2309 38084 -2301 38092
rect -2317 38078 -2309 38084
rect -2092 38083 -2062 38088
rect -2000 38079 -1992 38100
rect -1938 38099 -1906 38100
rect -1920 38098 -1906 38099
rect -1806 38092 -1680 38098
rect -1854 38083 -1806 38088
rect -1655 38084 -1647 38092
rect -1982 38079 -1966 38080
rect -2000 38078 -1966 38079
rect -1846 38078 -1806 38081
rect -1663 38078 -1655 38084
rect -1642 38078 -1637 38100
rect -1619 38078 -1614 38100
rect -1530 38078 -1526 38100
rect -1506 38078 -1502 38100
rect -1482 38078 -1478 38100
rect -1458 38078 -1454 38100
rect -1434 38078 -1430 38100
rect -1410 38078 -1406 38100
rect -1386 38079 -1382 38100
rect -1397 38078 -1363 38079
rect -2393 38076 -1363 38078
rect -2371 38054 -2366 38076
rect -2348 38054 -2343 38076
rect -2325 38054 -2320 38076
rect -2000 38074 -1966 38076
rect -2309 38056 -2301 38064
rect -2062 38063 -2054 38070
rect -2092 38056 -2084 38063
rect -2062 38056 -2026 38058
rect -2317 38054 -2309 38056
rect -2062 38054 -2012 38056
rect -2000 38054 -1992 38074
rect -1982 38073 -1966 38074
rect -1846 38072 -1806 38076
rect -1846 38065 -1798 38070
rect -1806 38063 -1798 38065
rect -1854 38061 -1846 38063
rect -1854 38056 -1806 38061
rect -1655 38056 -1647 38064
rect -1864 38054 -1796 38055
rect -1663 38054 -1655 38056
rect -1642 38054 -1637 38076
rect -1619 38054 -1614 38076
rect -1530 38054 -1526 38076
rect -1506 38054 -1502 38076
rect -1482 38054 -1478 38076
rect -1458 38054 -1454 38076
rect -1434 38054 -1430 38076
rect -1410 38054 -1406 38076
rect -1397 38069 -1392 38076
rect -1386 38069 -1382 38076
rect -1387 38055 -1382 38069
rect -1386 38054 -1382 38055
rect -1362 38054 -1358 38100
rect -1338 38054 -1334 38100
rect -1314 38054 -1310 38100
rect -1290 38054 -1286 38100
rect -1266 38054 -1262 38100
rect -1242 38054 -1238 38100
rect -1218 38054 -1214 38100
rect -1194 38054 -1190 38100
rect -1170 38054 -1166 38100
rect -1146 38054 -1142 38100
rect -1122 38054 -1118 38100
rect -1098 38054 -1094 38100
rect -1074 38054 -1070 38100
rect -1050 38054 -1046 38100
rect -1026 38054 -1022 38100
rect -1002 38054 -998 38100
rect -978 38054 -974 38100
rect -954 38054 -950 38100
rect -930 38054 -926 38100
rect -906 38054 -902 38100
rect -882 38054 -878 38100
rect -858 38054 -854 38100
rect -834 38054 -830 38100
rect -810 38054 -806 38100
rect -786 38054 -782 38100
rect -762 38054 -758 38100
rect -738 38054 -734 38100
rect -714 38054 -710 38100
rect -690 38054 -686 38100
rect -666 38054 -662 38100
rect -642 38054 -638 38100
rect -618 38054 -614 38100
rect -594 38054 -590 38100
rect -570 38054 -566 38100
rect -546 38054 -542 38100
rect -522 38054 -518 38100
rect -498 38054 -494 38100
rect -474 38054 -470 38100
rect -450 38054 -446 38100
rect -426 38054 -422 38100
rect -402 38054 -398 38100
rect -378 38054 -374 38100
rect -354 38054 -350 38100
rect -330 38054 -326 38100
rect -306 38054 -302 38100
rect -282 38054 -278 38100
rect -275 38099 -261 38100
rect -258 38099 -251 38127
rect -258 38054 -254 38099
rect -234 38075 -230 38172
rect -2393 38052 -237 38054
rect -2371 38006 -2366 38052
rect -2348 38006 -2343 38052
rect -2325 38006 -2320 38052
rect -2317 38048 -2309 38052
rect -2062 38048 -2054 38052
rect -2154 38044 -2138 38046
rect -2057 38044 -2054 38048
rect -2292 38038 -2054 38044
rect -2052 38038 -2044 38048
rect -2092 38022 -2062 38024
rect -2094 38018 -2062 38022
rect -2000 38006 -1992 38052
rect -1846 38045 -1806 38052
rect -1663 38048 -1655 38052
rect -1846 38038 -1680 38044
rect -1854 38022 -1806 38024
rect -1854 38018 -1680 38022
rect -1642 38006 -1637 38052
rect -1619 38006 -1614 38052
rect -1530 38006 -1526 38052
rect -1506 38006 -1502 38052
rect -1482 38006 -1478 38052
rect -1458 38006 -1454 38052
rect -1434 38006 -1430 38052
rect -1410 38006 -1406 38052
rect -1397 38021 -1392 38031
rect -1386 38021 -1382 38052
rect -1387 38007 -1382 38021
rect -1397 38006 -1363 38007
rect -2393 38004 -1363 38006
rect -2371 37982 -2366 38004
rect -2348 37982 -2343 38004
rect -2325 37982 -2320 38004
rect -2072 38002 -2036 38003
rect -2072 37996 -2054 38002
rect -2309 37988 -2301 37996
rect -2317 37982 -2309 37988
rect -2092 37987 -2062 37992
rect -2000 37983 -1992 38004
rect -1938 38003 -1906 38004
rect -1920 38002 -1906 38003
rect -1806 37996 -1680 38002
rect -1854 37987 -1806 37992
rect -1655 37988 -1647 37996
rect -1982 37983 -1966 37984
rect -2000 37982 -1966 37983
rect -1846 37982 -1806 37985
rect -1663 37982 -1655 37988
rect -1642 37982 -1637 38004
rect -1619 37982 -1614 38004
rect -1530 37982 -1526 38004
rect -1506 37982 -1502 38004
rect -1482 37982 -1478 38004
rect -1458 37982 -1454 38004
rect -1434 37982 -1430 38004
rect -1410 37982 -1406 38004
rect -1397 37997 -1392 38004
rect -1362 38003 -1358 38052
rect -1387 37983 -1382 37997
rect -1373 37993 -1365 37997
rect -1379 37983 -1373 37993
rect -1386 37982 -1382 37983
rect -2393 37980 -1365 37982
rect -2371 37958 -2366 37980
rect -2348 37958 -2343 37980
rect -2325 37958 -2320 37980
rect -2000 37978 -1966 37980
rect -2309 37960 -2301 37968
rect -2062 37967 -2054 37974
rect -2092 37960 -2084 37967
rect -2062 37960 -2026 37962
rect -2317 37958 -2309 37960
rect -2062 37958 -2012 37960
rect -2000 37958 -1992 37978
rect -1982 37977 -1966 37978
rect -1846 37976 -1806 37980
rect -1846 37969 -1798 37974
rect -1806 37967 -1798 37969
rect -1854 37965 -1846 37967
rect -1854 37960 -1806 37965
rect -1655 37960 -1647 37968
rect -1864 37958 -1796 37959
rect -1663 37958 -1655 37960
rect -1642 37958 -1637 37980
rect -1619 37958 -1614 37980
rect -1530 37958 -1526 37980
rect -1506 37958 -1502 37980
rect -1482 37958 -1478 37980
rect -1458 37958 -1454 37980
rect -1434 37958 -1430 37980
rect -1410 37958 -1406 37980
rect -1386 37958 -1382 37980
rect -1379 37979 -1365 37980
rect -1362 37979 -1355 38003
rect -1362 37958 -1358 37979
rect -1338 37958 -1334 38052
rect -1314 37958 -1310 38052
rect -1290 37958 -1286 38052
rect -1266 37958 -1262 38052
rect -1242 37958 -1238 38052
rect -1218 37958 -1214 38052
rect -1194 37958 -1190 38052
rect -1170 37958 -1166 38052
rect -1146 37958 -1142 38052
rect -1122 37958 -1118 38052
rect -1098 37958 -1094 38052
rect -1074 37958 -1070 38052
rect -1050 37958 -1046 38052
rect -1026 37958 -1022 38052
rect -1002 37958 -998 38052
rect -978 37958 -974 38052
rect -954 37958 -950 38052
rect -930 37958 -926 38052
rect -906 37958 -902 38052
rect -882 37958 -878 38052
rect -858 37958 -854 38052
rect -834 37958 -830 38052
rect -810 37958 -806 38052
rect -786 37958 -782 38052
rect -762 37958 -758 38052
rect -738 37959 -734 38052
rect -749 37958 -715 37959
rect -2393 37956 -715 37958
rect -2371 37910 -2366 37956
rect -2348 37910 -2343 37956
rect -2325 37910 -2320 37956
rect -2317 37952 -2309 37956
rect -2062 37952 -2054 37956
rect -2154 37948 -2138 37950
rect -2057 37948 -2054 37952
rect -2292 37942 -2054 37948
rect -2052 37942 -2044 37952
rect -2092 37926 -2062 37928
rect -2094 37922 -2062 37926
rect -2000 37910 -1992 37956
rect -1846 37949 -1806 37956
rect -1663 37952 -1655 37956
rect -1846 37942 -1680 37948
rect -1854 37926 -1806 37928
rect -1854 37922 -1680 37926
rect -1642 37910 -1637 37956
rect -1619 37910 -1614 37956
rect -1530 37910 -1526 37956
rect -1506 37910 -1502 37956
rect -1482 37910 -1478 37956
rect -1458 37910 -1454 37956
rect -1434 37910 -1430 37956
rect -1410 37910 -1406 37956
rect -1386 37910 -1382 37956
rect -1362 37955 -1358 37956
rect -2393 37908 -1365 37910
rect -2371 37886 -2366 37908
rect -2348 37886 -2343 37908
rect -2325 37886 -2320 37908
rect -2072 37906 -2036 37907
rect -2072 37900 -2054 37906
rect -2309 37892 -2301 37900
rect -2317 37886 -2309 37892
rect -2092 37891 -2062 37896
rect -2000 37887 -1992 37908
rect -1938 37907 -1906 37908
rect -1920 37906 -1906 37907
rect -1806 37900 -1680 37906
rect -1854 37891 -1806 37896
rect -1655 37892 -1647 37900
rect -1982 37887 -1966 37888
rect -2000 37886 -1966 37887
rect -1846 37886 -1806 37889
rect -1663 37886 -1655 37892
rect -1642 37886 -1637 37908
rect -1619 37886 -1614 37908
rect -1530 37886 -1526 37908
rect -1506 37886 -1502 37908
rect -1482 37886 -1478 37908
rect -1458 37886 -1454 37908
rect -1434 37886 -1430 37908
rect -1410 37886 -1406 37908
rect -1386 37886 -1382 37908
rect -1379 37907 -1365 37908
rect -1362 37907 -1355 37955
rect -1362 37886 -1358 37907
rect -1338 37886 -1334 37956
rect -1314 37886 -1310 37956
rect -1290 37886 -1286 37956
rect -1266 37886 -1262 37956
rect -1242 37886 -1238 37956
rect -1218 37886 -1214 37956
rect -1194 37886 -1190 37956
rect -1170 37886 -1166 37956
rect -1146 37886 -1142 37956
rect -1122 37886 -1118 37956
rect -1098 37886 -1094 37956
rect -1074 37886 -1070 37956
rect -1050 37886 -1046 37956
rect -1026 37886 -1022 37956
rect -1002 37886 -998 37956
rect -978 37886 -974 37956
rect -954 37886 -950 37956
rect -930 37886 -926 37956
rect -906 37886 -902 37956
rect -882 37886 -878 37956
rect -858 37886 -854 37956
rect -834 37886 -830 37956
rect -810 37886 -806 37956
rect -786 37886 -782 37956
rect -762 37886 -758 37956
rect -749 37949 -744 37956
rect -738 37949 -734 37956
rect -739 37935 -734 37949
rect -738 37886 -734 37935
rect -714 37886 -710 38052
rect -690 37935 -686 38052
rect -701 37934 -667 37935
rect -666 37934 -662 38052
rect -642 37934 -638 38052
rect -618 37934 -614 38052
rect -594 37934 -590 38052
rect -570 37934 -566 38052
rect -546 37934 -542 38052
rect -522 37934 -518 38052
rect -498 37934 -494 38052
rect -474 37934 -470 38052
rect -450 37934 -446 38052
rect -426 37934 -422 38052
rect -402 37934 -398 38052
rect -378 37934 -374 38052
rect -354 37934 -350 38052
rect -330 37934 -326 38052
rect -306 37934 -302 38052
rect -282 37934 -278 38052
rect -258 37934 -254 38052
rect -251 38051 -237 38052
rect -234 38051 -227 38075
rect -234 37934 -230 38051
rect -210 37934 -206 38172
rect -186 37934 -182 38172
rect -162 37934 -158 38172
rect -138 37934 -134 38172
rect -114 37934 -110 38172
rect -90 37934 -86 38172
rect -66 37934 -62 38172
rect -53 38165 -48 38172
rect -42 38165 -38 38172
rect -43 38151 -38 38165
rect -42 37934 -38 38151
rect -18 38099 -14 38220
rect -18 38075 -11 38099
rect -18 37934 -14 38075
rect 6 37934 10 38220
rect 30 37934 34 38220
rect 54 37934 58 38220
rect 78 37934 82 38220
rect 102 37934 106 38220
rect 115 38045 120 38055
rect 126 38045 130 38220
rect 125 38031 130 38045
rect 126 37934 130 38031
rect 150 38195 154 38220
rect 150 38171 157 38195
rect 150 37979 154 38171
rect 150 37955 157 37979
rect 150 37934 154 37955
rect 174 37934 178 38220
rect 198 37934 202 38220
rect 222 37934 226 38220
rect 246 37934 250 38220
rect 270 37934 274 38220
rect 294 37934 298 38220
rect 318 37934 322 38220
rect 342 37934 346 38220
rect 366 37934 370 38220
rect 390 37934 394 38220
rect 414 37934 418 38220
rect 438 37934 442 38220
rect 462 37934 466 38220
rect 486 37934 490 38220
rect 510 37934 514 38220
rect 534 37934 538 38220
rect 558 37934 562 38220
rect 582 37934 586 38220
rect 606 37934 610 38220
rect 630 37934 634 38220
rect 654 37934 658 38220
rect 678 37934 682 38220
rect 702 37934 706 38220
rect 726 37934 730 38220
rect 750 37934 754 38220
rect 774 37934 778 38220
rect 798 38127 802 38220
rect 787 38126 821 38127
rect 822 38126 826 38220
rect 846 38126 850 38220
rect 870 38126 874 38220
rect 894 38126 898 38220
rect 918 38126 922 38220
rect 942 38126 946 38220
rect 966 38126 970 38220
rect 990 38126 994 38220
rect 1014 38126 1018 38220
rect 1038 38126 1042 38220
rect 1045 38219 1059 38220
rect 1051 38213 1056 38219
rect 1061 38199 1066 38213
rect 1062 38126 1066 38199
rect 1075 38126 1083 38127
rect 787 38124 1083 38126
rect 787 38117 792 38124
rect 798 38117 802 38124
rect 797 38103 802 38117
rect 787 38093 792 38103
rect 797 38079 802 38093
rect 798 37934 802 38079
rect 822 38051 826 38124
rect 822 38030 829 38051
rect 846 38030 850 38124
rect 870 38030 874 38124
rect 894 38030 898 38124
rect 918 38030 922 38124
rect 942 38030 946 38124
rect 966 38030 970 38124
rect 990 38030 994 38124
rect 1014 38030 1018 38124
rect 1038 38030 1042 38124
rect 1062 38030 1066 38124
rect 1069 38123 1083 38124
rect 1075 38117 1080 38123
rect 1085 38103 1090 38117
rect 1086 38030 1090 38103
rect 1099 38030 1107 38031
rect 805 38028 1107 38030
rect 805 38027 819 38028
rect 822 38003 829 38028
rect 822 37934 826 38003
rect 846 37934 850 38028
rect 870 37934 874 38028
rect 894 37934 898 38028
rect 918 37934 922 38028
rect 942 37934 946 38028
rect 966 37934 970 38028
rect 990 37934 994 38028
rect 1014 37934 1018 38028
rect 1038 37934 1042 38028
rect 1062 37934 1066 38028
rect 1086 37934 1090 38028
rect 1093 38027 1107 38028
rect 1099 38021 1104 38027
rect 1109 38007 1114 38021
rect 1099 37973 1104 37983
rect 1110 37973 1114 38007
rect 1109 37959 1114 37973
rect 1099 37934 1131 37935
rect -701 37932 1131 37934
rect -701 37925 -696 37932
rect -690 37925 -686 37932
rect -691 37911 -686 37925
rect -701 37901 -696 37911
rect -691 37887 -686 37901
rect -690 37886 -686 37887
rect -666 37886 -662 37932
rect -642 37886 -638 37932
rect -618 37886 -614 37932
rect -594 37886 -590 37932
rect -570 37886 -566 37932
rect -546 37886 -542 37932
rect -522 37886 -518 37932
rect -498 37886 -494 37932
rect -474 37886 -470 37932
rect -450 37886 -446 37932
rect -426 37886 -422 37932
rect -402 37886 -398 37932
rect -378 37886 -374 37932
rect -354 37886 -350 37932
rect -330 37886 -326 37932
rect -306 37886 -302 37932
rect -282 37886 -278 37932
rect -258 37886 -254 37932
rect -234 37886 -230 37932
rect -210 37886 -206 37932
rect -186 37886 -182 37932
rect -162 37886 -158 37932
rect -138 37886 -134 37932
rect -114 37886 -110 37932
rect -90 37886 -86 37932
rect -66 37886 -62 37932
rect -42 37886 -38 37932
rect -18 37886 -14 37932
rect 6 37886 10 37932
rect 30 37886 34 37932
rect 54 37886 58 37932
rect 78 37886 82 37932
rect 102 37886 106 37932
rect 126 37886 130 37932
rect 150 37886 154 37932
rect 174 37886 178 37932
rect 198 37886 202 37932
rect 222 37886 226 37932
rect 246 37886 250 37932
rect 270 37886 274 37932
rect 294 37886 298 37932
rect 318 37886 322 37932
rect 342 37886 346 37932
rect 366 37886 370 37932
rect 390 37886 394 37932
rect 414 37886 418 37932
rect 438 37886 442 37932
rect 462 37886 466 37932
rect 486 37886 490 37932
rect 510 37886 514 37932
rect 534 37886 538 37932
rect 558 37886 562 37932
rect 582 37886 586 37932
rect 606 37886 610 37932
rect 630 37886 634 37932
rect 654 37886 658 37932
rect 678 37886 682 37932
rect 702 37886 706 37932
rect 726 37886 730 37932
rect 750 37886 754 37932
rect 774 37886 778 37932
rect 798 37886 802 37932
rect 822 37886 826 37932
rect 846 37886 850 37932
rect 870 37886 874 37932
rect 894 37886 898 37932
rect 918 37886 922 37932
rect 942 37886 946 37932
rect 966 37887 970 37932
rect 955 37886 989 37887
rect -2393 37884 989 37886
rect -2371 37862 -2366 37884
rect -2348 37862 -2343 37884
rect -2325 37862 -2320 37884
rect -2000 37882 -1966 37884
rect -2309 37864 -2301 37872
rect -2062 37871 -2054 37878
rect -2092 37864 -2084 37871
rect -2062 37864 -2026 37866
rect -2317 37862 -2309 37864
rect -2062 37862 -2012 37864
rect -2000 37862 -1992 37882
rect -1982 37881 -1966 37882
rect -1846 37880 -1806 37884
rect -1846 37873 -1798 37878
rect -1806 37871 -1798 37873
rect -1854 37869 -1846 37871
rect -1854 37864 -1806 37869
rect -1655 37864 -1647 37872
rect -1864 37862 -1796 37863
rect -1663 37862 -1655 37864
rect -1642 37862 -1637 37884
rect -1619 37862 -1614 37884
rect -1530 37862 -1526 37884
rect -1506 37862 -1502 37884
rect -1482 37862 -1478 37884
rect -1458 37862 -1454 37884
rect -1434 37862 -1430 37884
rect -1410 37862 -1406 37884
rect -1386 37862 -1382 37884
rect -1362 37862 -1358 37884
rect -1338 37862 -1334 37884
rect -1314 37862 -1310 37884
rect -1290 37862 -1286 37884
rect -1266 37862 -1262 37884
rect -1242 37862 -1238 37884
rect -1218 37862 -1214 37884
rect -1194 37862 -1190 37884
rect -1170 37862 -1166 37884
rect -1146 37862 -1142 37884
rect -1122 37862 -1118 37884
rect -1098 37862 -1094 37884
rect -1074 37862 -1070 37884
rect -1050 37862 -1046 37884
rect -1026 37862 -1022 37884
rect -1002 37862 -998 37884
rect -978 37862 -974 37884
rect -954 37862 -950 37884
rect -930 37862 -926 37884
rect -906 37862 -902 37884
rect -882 37862 -878 37884
rect -858 37862 -854 37884
rect -834 37862 -830 37884
rect -810 37862 -806 37884
rect -786 37862 -782 37884
rect -762 37862 -758 37884
rect -738 37862 -734 37884
rect -714 37883 -710 37884
rect -2393 37860 -717 37862
rect -2371 37814 -2366 37860
rect -2348 37814 -2343 37860
rect -2325 37814 -2320 37860
rect -2317 37856 -2309 37860
rect -2062 37856 -2054 37860
rect -2154 37852 -2138 37854
rect -2057 37852 -2054 37856
rect -2292 37846 -2054 37852
rect -2052 37846 -2044 37856
rect -2092 37830 -2062 37832
rect -2094 37826 -2062 37830
rect -2000 37814 -1992 37860
rect -1846 37853 -1806 37860
rect -1663 37856 -1655 37860
rect -1846 37846 -1680 37852
rect -1854 37830 -1806 37832
rect -1854 37826 -1680 37830
rect -1642 37814 -1637 37860
rect -1619 37814 -1614 37860
rect -1530 37814 -1526 37860
rect -1506 37814 -1502 37860
rect -1482 37814 -1478 37860
rect -1458 37814 -1454 37860
rect -1434 37814 -1430 37860
rect -1410 37814 -1406 37860
rect -1397 37829 -1392 37839
rect -1386 37829 -1382 37860
rect -1387 37815 -1382 37829
rect -1397 37814 -1363 37815
rect -2393 37812 -1363 37814
rect -2371 37790 -2366 37812
rect -2348 37790 -2343 37812
rect -2325 37790 -2320 37812
rect -2072 37810 -2036 37811
rect -2072 37804 -2054 37810
rect -2309 37796 -2301 37804
rect -2317 37790 -2309 37796
rect -2092 37795 -2062 37800
rect -2000 37791 -1992 37812
rect -1938 37811 -1906 37812
rect -1920 37810 -1906 37811
rect -1806 37804 -1680 37810
rect -1854 37795 -1806 37800
rect -1655 37796 -1647 37804
rect -1982 37791 -1966 37792
rect -2000 37790 -1966 37791
rect -1846 37790 -1806 37793
rect -1663 37790 -1655 37796
rect -1642 37790 -1637 37812
rect -1619 37790 -1614 37812
rect -1530 37790 -1526 37812
rect -1506 37790 -1502 37812
rect -1482 37790 -1478 37812
rect -1458 37790 -1454 37812
rect -1434 37790 -1430 37812
rect -1410 37790 -1406 37812
rect -1397 37805 -1392 37812
rect -1387 37791 -1382 37805
rect -1362 37791 -1358 37860
rect -1386 37790 -1382 37791
rect -1373 37790 -1339 37791
rect -2393 37788 -1339 37790
rect -2371 37766 -2366 37788
rect -2348 37766 -2343 37788
rect -2325 37766 -2320 37788
rect -2000 37786 -1966 37788
rect -2309 37768 -2301 37776
rect -2062 37775 -2054 37782
rect -2092 37768 -2084 37775
rect -2062 37768 -2026 37770
rect -2317 37766 -2309 37768
rect -2062 37766 -2012 37768
rect -2000 37766 -1992 37786
rect -1982 37785 -1966 37786
rect -1846 37784 -1806 37788
rect -1846 37777 -1798 37782
rect -1806 37775 -1798 37777
rect -1854 37773 -1846 37775
rect -1854 37768 -1806 37773
rect -1655 37768 -1647 37776
rect -1864 37766 -1796 37767
rect -1663 37766 -1655 37768
rect -1642 37766 -1637 37788
rect -1619 37766 -1614 37788
rect -1530 37766 -1526 37788
rect -1506 37766 -1502 37788
rect -1482 37766 -1478 37788
rect -1458 37766 -1454 37788
rect -1434 37766 -1430 37788
rect -1410 37766 -1406 37788
rect -1386 37766 -1382 37788
rect -1373 37781 -1368 37788
rect -1362 37781 -1358 37788
rect -1363 37767 -1358 37781
rect -1338 37767 -1334 37860
rect -1362 37766 -1358 37767
rect -1349 37766 -1315 37767
rect -2393 37764 -1315 37766
rect -2371 37718 -2366 37764
rect -2348 37718 -2343 37764
rect -2325 37718 -2320 37764
rect -2317 37760 -2309 37764
rect -2062 37760 -2054 37764
rect -2154 37756 -2138 37758
rect -2057 37756 -2054 37760
rect -2292 37750 -2054 37756
rect -2052 37750 -2044 37760
rect -2092 37734 -2062 37736
rect -2094 37730 -2062 37734
rect -2000 37718 -1992 37764
rect -1846 37757 -1806 37764
rect -1663 37760 -1655 37764
rect -1846 37750 -1680 37756
rect -1854 37734 -1806 37736
rect -1854 37730 -1680 37734
rect -1642 37718 -1637 37764
rect -1619 37718 -1614 37764
rect -1530 37718 -1526 37764
rect -1506 37718 -1502 37764
rect -1482 37718 -1478 37764
rect -1458 37718 -1454 37764
rect -1434 37718 -1430 37764
rect -1410 37718 -1406 37764
rect -1386 37718 -1382 37764
rect -1362 37763 -1358 37764
rect -2393 37716 -1365 37718
rect -2371 37694 -2366 37716
rect -2348 37694 -2343 37716
rect -2325 37694 -2320 37716
rect -2072 37714 -2036 37715
rect -2072 37708 -2054 37714
rect -2309 37700 -2301 37708
rect -2317 37694 -2309 37700
rect -2092 37699 -2062 37704
rect -2000 37695 -1992 37716
rect -1938 37715 -1906 37716
rect -1920 37714 -1906 37715
rect -1806 37708 -1680 37714
rect -1854 37699 -1806 37704
rect -1655 37700 -1647 37708
rect -1982 37695 -1966 37696
rect -2000 37694 -1966 37695
rect -1846 37694 -1806 37697
rect -1663 37694 -1655 37700
rect -1642 37694 -1637 37716
rect -1619 37694 -1614 37716
rect -1530 37694 -1526 37716
rect -1506 37694 -1502 37716
rect -1482 37694 -1478 37716
rect -1458 37694 -1454 37716
rect -1434 37694 -1430 37716
rect -1410 37694 -1406 37716
rect -1386 37694 -1382 37716
rect -1379 37715 -1365 37716
rect -1362 37715 -1355 37763
rect -1349 37757 -1344 37764
rect -1338 37757 -1334 37764
rect -1339 37743 -1334 37757
rect -1338 37715 -1334 37743
rect -1362 37694 -1358 37715
rect -2393 37692 -1341 37694
rect -2371 37670 -2366 37692
rect -2348 37670 -2343 37692
rect -2325 37670 -2320 37692
rect -2000 37690 -1966 37692
rect -2309 37672 -2301 37680
rect -2062 37679 -2054 37686
rect -2092 37672 -2084 37679
rect -2062 37672 -2026 37674
rect -2317 37670 -2309 37672
rect -2062 37670 -2012 37672
rect -2000 37670 -1992 37690
rect -1982 37689 -1966 37690
rect -1846 37688 -1806 37692
rect -1846 37681 -1798 37686
rect -1806 37679 -1798 37681
rect -1854 37677 -1846 37679
rect -1854 37672 -1806 37677
rect -1655 37672 -1647 37680
rect -1864 37670 -1796 37671
rect -1663 37670 -1655 37672
rect -1642 37670 -1637 37692
rect -1619 37670 -1614 37692
rect -1530 37670 -1526 37692
rect -1506 37670 -1502 37692
rect -1482 37670 -1478 37692
rect -1458 37670 -1454 37692
rect -1434 37670 -1430 37692
rect -1410 37670 -1406 37692
rect -1386 37670 -1382 37692
rect -1362 37670 -1358 37692
rect -1355 37691 -1341 37692
rect -1338 37691 -1331 37715
rect -1314 37691 -1310 37860
rect -1338 37670 -1334 37691
rect -2393 37668 -1317 37670
rect -2371 37622 -2366 37668
rect -2348 37622 -2343 37668
rect -2325 37622 -2320 37668
rect -2317 37664 -2309 37668
rect -2062 37664 -2054 37668
rect -2154 37660 -2138 37662
rect -2057 37660 -2054 37664
rect -2292 37654 -2054 37660
rect -2052 37654 -2044 37664
rect -2092 37638 -2062 37640
rect -2094 37634 -2062 37638
rect -2000 37622 -1992 37668
rect -1846 37661 -1806 37668
rect -1663 37664 -1655 37668
rect -1846 37654 -1680 37660
rect -1854 37638 -1806 37640
rect -1854 37634 -1680 37638
rect -1642 37622 -1637 37668
rect -1619 37622 -1614 37668
rect -1530 37622 -1526 37668
rect -1506 37622 -1502 37668
rect -1482 37622 -1478 37668
rect -1458 37622 -1454 37668
rect -1434 37622 -1430 37668
rect -1410 37622 -1406 37668
rect -1386 37622 -1382 37668
rect -1362 37622 -1358 37668
rect -1338 37622 -1334 37668
rect -1331 37667 -1317 37668
rect -1314 37667 -1307 37691
rect -1314 37622 -1310 37667
rect -1290 37622 -1286 37860
rect -1266 37622 -1262 37860
rect -1242 37622 -1238 37860
rect -1218 37622 -1214 37860
rect -1194 37622 -1190 37860
rect -1170 37622 -1166 37860
rect -1146 37622 -1142 37860
rect -1122 37622 -1118 37860
rect -1098 37622 -1094 37860
rect -1074 37622 -1070 37860
rect -1050 37622 -1046 37860
rect -1026 37622 -1022 37860
rect -1002 37622 -998 37860
rect -978 37622 -974 37860
rect -954 37622 -950 37860
rect -930 37622 -926 37860
rect -906 37622 -902 37860
rect -882 37622 -878 37860
rect -858 37622 -854 37860
rect -834 37622 -830 37860
rect -810 37622 -806 37860
rect -786 37622 -782 37860
rect -762 37622 -758 37860
rect -738 37622 -734 37860
rect -731 37859 -717 37860
rect -714 37859 -707 37883
rect -714 37622 -710 37859
rect -690 37622 -686 37884
rect -666 37859 -662 37884
rect -666 37838 -659 37859
rect -642 37838 -638 37884
rect -618 37838 -614 37884
rect -594 37838 -590 37884
rect -570 37838 -566 37884
rect -546 37838 -542 37884
rect -522 37838 -518 37884
rect -498 37838 -494 37884
rect -474 37838 -470 37884
rect -450 37838 -446 37884
rect -426 37838 -422 37884
rect -402 37838 -398 37884
rect -378 37838 -374 37884
rect -354 37838 -350 37884
rect -330 37838 -326 37884
rect -306 37838 -302 37884
rect -282 37838 -278 37884
rect -258 37838 -254 37884
rect -234 37838 -230 37884
rect -210 37838 -206 37884
rect -186 37838 -182 37884
rect -162 37838 -158 37884
rect -138 37838 -134 37884
rect -114 37838 -110 37884
rect -90 37838 -86 37884
rect -66 37838 -62 37884
rect -42 37838 -38 37884
rect -18 37838 -14 37884
rect 6 37838 10 37884
rect 30 37838 34 37884
rect 54 37838 58 37884
rect 78 37838 82 37884
rect 102 37838 106 37884
rect 126 37838 130 37884
rect 150 37838 154 37884
rect 174 37838 178 37884
rect 198 37838 202 37884
rect 222 37838 226 37884
rect 246 37838 250 37884
rect 270 37838 274 37884
rect 294 37838 298 37884
rect 318 37838 322 37884
rect 342 37838 346 37884
rect 366 37838 370 37884
rect 390 37838 394 37884
rect 414 37838 418 37884
rect 438 37838 442 37884
rect 462 37838 466 37884
rect 486 37838 490 37884
rect 510 37838 514 37884
rect 534 37838 538 37884
rect 558 37838 562 37884
rect 582 37838 586 37884
rect 606 37838 610 37884
rect 630 37838 634 37884
rect 654 37838 658 37884
rect 678 37838 682 37884
rect 702 37838 706 37884
rect 726 37838 730 37884
rect 750 37838 754 37884
rect 774 37838 778 37884
rect 798 37838 802 37884
rect 822 37838 826 37884
rect 846 37838 850 37884
rect 870 37838 874 37884
rect 894 37838 898 37884
rect 918 37838 922 37884
rect 942 37838 946 37884
rect 955 37877 960 37884
rect 966 37877 970 37884
rect 965 37863 970 37877
rect 966 37838 970 37863
rect 990 37838 994 37932
rect 1014 37838 1018 37932
rect 1038 37838 1042 37932
rect 1051 37853 1056 37863
rect 1062 37853 1066 37932
rect 1061 37839 1066 37853
rect 1062 37838 1066 37839
rect 1086 37838 1090 37932
rect 1099 37925 1104 37932
rect 1117 37931 1131 37932
rect 1109 37911 1114 37925
rect 1110 37838 1114 37911
rect 1123 37838 1131 37839
rect -683 37836 1131 37838
rect -683 37835 -669 37836
rect -666 37811 -659 37836
rect -666 37622 -662 37811
rect -642 37622 -638 37836
rect -618 37622 -614 37836
rect -594 37622 -590 37836
rect -570 37622 -566 37836
rect -546 37622 -542 37836
rect -522 37622 -518 37836
rect -498 37622 -494 37836
rect -474 37622 -470 37836
rect -450 37622 -446 37836
rect -426 37622 -422 37836
rect -402 37622 -398 37836
rect -378 37622 -374 37836
rect -354 37622 -350 37836
rect -330 37622 -326 37836
rect -306 37622 -302 37836
rect -282 37622 -278 37836
rect -258 37622 -254 37836
rect -234 37622 -230 37836
rect -210 37622 -206 37836
rect -186 37622 -182 37836
rect -162 37622 -158 37836
rect -138 37622 -134 37836
rect -114 37622 -110 37836
rect -90 37622 -86 37836
rect -66 37622 -62 37836
rect -42 37622 -38 37836
rect -18 37622 -14 37836
rect 6 37622 10 37836
rect 30 37622 34 37836
rect 54 37622 58 37836
rect 78 37622 82 37836
rect 102 37622 106 37836
rect 126 37622 130 37836
rect 150 37743 154 37836
rect 139 37742 173 37743
rect 174 37742 178 37836
rect 198 37742 202 37836
rect 222 37742 226 37836
rect 246 37742 250 37836
rect 270 37742 274 37836
rect 294 37742 298 37836
rect 318 37742 322 37836
rect 342 37742 346 37836
rect 366 37742 370 37836
rect 390 37742 394 37836
rect 414 37742 418 37836
rect 438 37742 442 37836
rect 462 37742 466 37836
rect 486 37742 490 37836
rect 510 37742 514 37836
rect 534 37742 538 37836
rect 558 37742 562 37836
rect 582 37742 586 37836
rect 606 37742 610 37836
rect 630 37742 634 37836
rect 654 37742 658 37836
rect 678 37742 682 37836
rect 702 37742 706 37836
rect 726 37742 730 37836
rect 750 37742 754 37836
rect 774 37742 778 37836
rect 798 37742 802 37836
rect 822 37742 826 37836
rect 846 37742 850 37836
rect 870 37742 874 37836
rect 894 37742 898 37836
rect 918 37742 922 37836
rect 942 37742 946 37836
rect 966 37742 970 37836
rect 990 37811 994 37836
rect 990 37787 997 37811
rect 990 37742 994 37787
rect 1014 37742 1018 37836
rect 1038 37742 1042 37836
rect 1062 37742 1066 37836
rect 1086 37787 1090 37836
rect 1086 37763 1093 37787
rect 1086 37742 1090 37763
rect 1110 37742 1114 37836
rect 1117 37835 1131 37836
rect 1123 37829 1128 37835
rect 1133 37815 1138 37829
rect 1134 37742 1138 37815
rect 1147 37742 1155 37743
rect 139 37740 1155 37742
rect 139 37733 144 37740
rect 150 37733 154 37740
rect 149 37719 154 37733
rect 139 37709 144 37719
rect 149 37695 154 37709
rect 150 37622 154 37695
rect 174 37667 178 37740
rect -2393 37620 171 37622
rect -2371 37574 -2366 37620
rect -2348 37574 -2343 37620
rect -2325 37574 -2320 37620
rect -2309 37604 -2301 37614
rect -2317 37598 -2309 37604
rect -2097 37598 -2095 37607
rect -2309 37576 -2301 37586
rect -2097 37584 -2095 37588
rect -2292 37583 -2095 37584
rect -2097 37581 -2095 37583
rect -2084 37576 -2083 37619
rect -2069 37612 -2054 37614
rect -2054 37596 -2018 37598
rect -2054 37594 -2004 37596
rect -2059 37590 -2045 37594
rect -2054 37588 -2049 37590
rect -2317 37574 -2309 37576
rect -2084 37574 -2054 37576
rect -2044 37574 -2039 37588
rect -2025 37578 -2014 37584
rect -2000 37578 -1992 37620
rect -1920 37618 -1906 37620
rect -1977 37603 -1929 37609
rect -1655 37604 -1647 37614
rect -1977 37593 -1966 37603
rect -1663 37598 -1655 37604
rect -1977 37581 -1929 37583
rect -2033 37574 -1992 37578
rect -1655 37576 -1647 37586
rect -1663 37574 -1655 37576
rect -1642 37574 -1637 37620
rect -1619 37574 -1614 37620
rect -1530 37574 -1526 37620
rect -1506 37574 -1502 37620
rect -1482 37574 -1478 37620
rect -1458 37574 -1454 37620
rect -1434 37574 -1430 37620
rect -1410 37574 -1406 37620
rect -1386 37574 -1382 37620
rect -1362 37575 -1358 37620
rect -1373 37574 -1339 37575
rect -2393 37572 -1339 37574
rect -2371 37454 -2366 37572
rect -2348 37454 -2343 37572
rect -2325 37538 -2320 37572
rect -2317 37570 -2309 37572
rect -2084 37559 -2083 37572
rect -2084 37558 -2054 37559
rect -2325 37530 -2317 37538
rect -2325 37510 -2320 37530
rect -2317 37522 -2309 37530
rect -2117 37521 -2095 37531
rect -2045 37528 -2037 37542
rect -2325 37494 -2317 37510
rect -2325 37478 -2320 37494
rect -2309 37482 -2301 37494
rect -2317 37478 -2309 37482
rect -2117 37480 -2095 37487
rect -2069 37486 -2041 37494
rect -2017 37492 -2015 37494
rect -2325 37466 -2317 37478
rect -2125 37471 -2095 37478
rect -2047 37476 -2011 37478
rect -2059 37474 -2011 37476
rect -2000 37474 -1992 37572
rect -1663 37570 -1655 37572
rect -1969 37521 -1929 37533
rect -1671 37530 -1663 37538
rect -1663 37522 -1655 37530
rect -1671 37494 -1663 37510
rect -1655 37482 -1647 37494
rect -1663 37478 -1655 37482
rect -2125 37469 -2117 37471
rect -2059 37470 -2045 37474
rect -2021 37471 -1992 37474
rect -1977 37471 -1929 37478
rect -2325 37454 -2320 37466
rect -2309 37454 -2301 37466
rect -2131 37461 -2129 37466
rect -2125 37463 -2095 37469
rect -2021 37464 -2009 37468
rect -2125 37461 -2117 37463
rect -2133 37454 -2129 37461
rect -2117 37454 -2087 37461
rect -2025 37458 -2021 37464
rect -2000 37458 -1992 37471
rect -1969 37463 -1929 37469
rect -1671 37466 -1663 37478
rect -2033 37454 -1992 37458
rect -1969 37454 -1921 37461
rect -1655 37454 -1647 37466
rect -1642 37454 -1637 37572
rect -1619 37454 -1614 37572
rect -1530 37454 -1526 37572
rect -1506 37454 -1502 37572
rect -1482 37454 -1478 37572
rect -1458 37454 -1454 37572
rect -1434 37454 -1430 37572
rect -1410 37454 -1406 37572
rect -1386 37454 -1382 37572
rect -1373 37565 -1368 37572
rect -1362 37565 -1358 37572
rect -1363 37551 -1358 37565
rect -1362 37455 -1358 37551
rect -1349 37541 -1344 37551
rect -1338 37541 -1334 37620
rect -1339 37527 -1334 37541
rect -1338 37499 -1334 37527
rect -1338 37475 -1331 37499
rect -1314 37475 -1310 37620
rect -1373 37454 -1339 37455
rect -2393 37452 -1339 37454
rect -2371 37358 -2366 37452
rect -2348 37358 -2343 37452
rect -2325 37450 -2320 37452
rect -2317 37450 -2309 37452
rect -2131 37450 -2129 37452
rect -2125 37450 -2095 37452
rect -2325 37438 -2317 37450
rect -2117 37445 -2095 37450
rect -2325 37418 -2320 37438
rect -2325 37410 -2317 37418
rect -2325 37358 -2320 37410
rect -2317 37402 -2309 37410
rect -2117 37401 -2095 37411
rect -2045 37408 -2037 37422
rect -2309 37362 -2301 37370
rect -2317 37358 -2309 37362
rect -2000 37358 -1992 37452
rect -1663 37450 -1655 37452
rect -1671 37438 -1663 37450
rect -1969 37401 -1929 37413
rect -1671 37410 -1663 37418
rect -1663 37402 -1655 37410
rect -1655 37362 -1647 37370
rect -1663 37358 -1655 37362
rect -1642 37358 -1637 37452
rect -1619 37358 -1614 37452
rect -1530 37358 -1526 37452
rect -1506 37358 -1502 37452
rect -1482 37358 -1478 37452
rect -1458 37358 -1454 37452
rect -1434 37358 -1430 37452
rect -1410 37358 -1406 37452
rect -1386 37358 -1382 37452
rect -1373 37445 -1368 37452
rect -1362 37445 -1358 37452
rect -1363 37431 -1358 37445
rect -1362 37358 -1358 37431
rect -1338 37379 -1334 37475
rect -1314 37451 -1307 37475
rect -2393 37356 -2026 37358
rect -2021 37356 -1341 37358
rect -2371 37214 -2366 37356
rect -2348 37214 -2343 37356
rect -2325 37294 -2320 37356
rect -2317 37354 -2309 37356
rect -2309 37334 -2301 37342
rect -2317 37326 -2309 37334
rect -2123 37329 -2116 37334
rect -2123 37327 -2092 37329
rect -2091 37328 -2087 37344
rect -2026 37336 -2021 37348
rect -2037 37332 -2021 37336
rect -2292 37325 -2087 37327
rect -2123 37323 -2116 37325
rect -2325 37286 -2317 37294
rect -2325 37238 -2320 37286
rect -2317 37278 -2309 37286
rect -2083 37252 -2053 37254
rect -2124 37241 -2119 37246
rect -2325 37234 -2317 37238
rect -2325 37214 -2320 37234
rect -2317 37222 -2306 37234
rect -2112 37229 -2107 37241
rect -2018 37232 -2002 37238
rect -2159 37228 -2107 37229
rect -2159 37225 -2096 37228
rect -2083 37225 -2053 37228
rect -2018 37223 -2017 37228
rect -2307 37218 -2306 37222
rect -2017 37218 -2008 37223
rect -2000 37214 -1992 37356
rect -1663 37354 -1655 37356
rect -1969 37328 -1932 37344
rect -1655 37334 -1647 37342
rect -1969 37325 -1680 37327
rect -1663 37326 -1655 37334
rect -1671 37286 -1663 37294
rect -1663 37278 -1655 37286
rect -1972 37252 -1924 37254
rect -1674 37237 -1663 37238
rect -1946 37228 -1932 37237
rect -1972 37225 -1924 37228
rect -1794 37226 -1758 37234
rect -1794 37225 -1680 37226
rect -1663 37222 -1658 37237
rect -1923 37214 -1889 37215
rect -1642 37214 -1637 37356
rect -1619 37214 -1614 37356
rect -1530 37214 -1526 37356
rect -1506 37214 -1502 37356
rect -1482 37214 -1478 37356
rect -1458 37214 -1454 37356
rect -1434 37214 -1430 37356
rect -1410 37214 -1406 37356
rect -1386 37214 -1382 37356
rect -1362 37214 -1358 37356
rect -1355 37355 -1341 37356
rect -1338 37355 -1331 37379
rect -1338 37214 -1334 37355
rect -1314 37214 -1310 37451
rect -1290 37214 -1286 37620
rect -1266 37214 -1262 37620
rect -1242 37214 -1238 37620
rect -1218 37214 -1214 37620
rect -1194 37214 -1190 37620
rect -1170 37214 -1166 37620
rect -1146 37214 -1142 37620
rect -1122 37214 -1118 37620
rect -1098 37214 -1094 37620
rect -1074 37214 -1070 37620
rect -1050 37214 -1046 37620
rect -1037 37301 -1032 37311
rect -1026 37301 -1022 37620
rect -1027 37287 -1022 37301
rect -1026 37214 -1022 37287
rect -1002 37235 -998 37620
rect -2393 37212 -1005 37214
rect -2371 37142 -2366 37212
rect -2348 37142 -2343 37212
rect -2325 37210 -2320 37212
rect -2325 37206 -2317 37210
rect -2325 37158 -2320 37206
rect -2317 37194 -2306 37206
rect -2153 37180 -2147 37182
rect -2153 37178 -2101 37180
rect -2153 37172 -2054 37178
rect -2307 37162 -2306 37170
rect -2325 37150 -2314 37158
rect -2104 37154 -2101 37158
rect -2104 37152 -2101 37153
rect -2000 37152 -1992 37212
rect -1674 37209 -1663 37210
rect -1663 37194 -1658 37209
rect -1758 37175 -1692 37181
rect -1758 37172 -1710 37175
rect -1750 37163 -1702 37170
rect -1917 37156 -1901 37162
rect -1828 37158 -1792 37162
rect -1916 37152 -1914 37156
rect -1750 37155 -1710 37161
rect -1700 37155 -1692 37175
rect -1674 37164 -1665 37173
rect -1674 37152 -1666 37161
rect -2325 37142 -2320 37150
rect -2314 37142 -2306 37150
rect -2139 37143 -2123 37152
rect -2111 37145 -2016 37152
rect -2139 37142 -2111 37143
rect -2104 37142 -2101 37145
rect -2021 37142 -2016 37145
rect -2000 37145 -1818 37152
rect -1802 37145 -1776 37152
rect -1760 37145 -1710 37152
rect -1666 37145 -1658 37152
rect -2000 37142 -1992 37145
rect -1758 37143 -1755 37145
rect -1758 37142 -1757 37143
rect -1710 37142 -1702 37143
rect -1674 37142 -1665 37145
rect -1642 37142 -1637 37212
rect -1619 37142 -1614 37212
rect -1530 37142 -1526 37212
rect -1506 37142 -1502 37212
rect -1482 37142 -1478 37212
rect -1458 37142 -1454 37212
rect -1434 37142 -1430 37212
rect -1410 37142 -1406 37212
rect -1386 37142 -1382 37212
rect -1362 37142 -1358 37212
rect -1338 37142 -1334 37212
rect -1314 37142 -1310 37212
rect -1290 37142 -1286 37212
rect -1266 37142 -1262 37212
rect -1242 37142 -1238 37212
rect -1218 37142 -1214 37212
rect -1194 37142 -1190 37212
rect -1170 37142 -1166 37212
rect -1146 37142 -1142 37212
rect -1122 37142 -1118 37212
rect -1098 37142 -1094 37212
rect -1074 37142 -1070 37212
rect -1050 37142 -1046 37212
rect -1026 37142 -1022 37212
rect -1019 37211 -1005 37212
rect -1002 37211 -995 37235
rect -1002 37142 -998 37211
rect -978 37142 -974 37620
rect -954 37142 -950 37620
rect -941 37157 -936 37167
rect -930 37157 -926 37620
rect -931 37143 -926 37157
rect -930 37142 -926 37143
rect -906 37142 -902 37620
rect -882 37142 -878 37620
rect -858 37142 -854 37620
rect -834 37142 -830 37620
rect -810 37142 -806 37620
rect -786 37142 -782 37620
rect -762 37142 -758 37620
rect -738 37142 -734 37620
rect -714 37142 -710 37620
rect -690 37142 -686 37620
rect -666 37142 -662 37620
rect -642 37142 -638 37620
rect -618 37142 -614 37620
rect -594 37142 -590 37620
rect -570 37142 -566 37620
rect -546 37142 -542 37620
rect -522 37142 -518 37620
rect -498 37142 -494 37620
rect -474 37142 -470 37620
rect -450 37142 -446 37620
rect -426 37142 -422 37620
rect -402 37142 -398 37620
rect -378 37142 -374 37620
rect -354 37142 -350 37620
rect -330 37142 -326 37620
rect -306 37142 -302 37620
rect -282 37142 -278 37620
rect -258 37142 -254 37620
rect -234 37142 -230 37620
rect -210 37142 -206 37620
rect -186 37142 -182 37620
rect -162 37142 -158 37620
rect -138 37142 -134 37620
rect -114 37142 -110 37620
rect -90 37142 -86 37620
rect -66 37142 -62 37620
rect -42 37142 -38 37620
rect -18 37142 -14 37620
rect 6 37142 10 37620
rect 30 37142 34 37620
rect 54 37142 58 37620
rect 78 37142 82 37620
rect 102 37142 106 37620
rect 126 37142 130 37620
rect 150 37142 154 37620
rect 157 37619 171 37620
rect 174 37619 181 37667
rect 174 37142 178 37619
rect 198 37142 202 37740
rect 222 37142 226 37740
rect 246 37142 250 37740
rect 270 37142 274 37740
rect 283 37685 288 37695
rect 294 37685 298 37740
rect 293 37671 298 37685
rect 294 37143 298 37671
rect 318 37619 322 37740
rect 318 37595 325 37619
rect 283 37142 317 37143
rect -2393 37140 317 37142
rect -2371 37070 -2366 37140
rect -2348 37070 -2343 37140
rect -2325 37130 -2320 37140
rect -2307 37134 -2306 37140
rect -2139 37136 -2111 37140
rect -2325 37122 -2314 37130
rect -2141 37127 -2119 37131
rect -2325 37102 -2320 37122
rect -2314 37114 -2306 37122
rect -2149 37115 -2141 37122
rect -2307 37106 -2306 37114
rect -2104 37112 -2101 37140
rect -2076 37136 -2046 37139
rect -2076 37123 -2054 37131
rect -2021 37128 -2016 37140
rect -2084 37121 -2036 37122
rect -2000 37121 -1992 37140
rect -1931 37136 -1895 37140
rect -1768 37132 -1760 37140
rect -1758 37136 -1757 37140
rect -1750 37136 -1702 37140
rect -1674 37136 -1665 37140
rect -1768 37131 -1764 37132
rect -1758 37131 -1755 37136
rect -1932 37121 -1917 37130
rect -2084 37118 -1917 37121
rect -1916 37121 -1905 37123
rect -1758 37122 -1754 37131
rect -1750 37124 -1710 37131
rect -1674 37124 -1666 37133
rect -1758 37121 -1692 37122
rect -1916 37119 -1692 37121
rect -1916 37118 -1690 37119
rect -2084 37114 -2054 37118
rect -2046 37114 -1932 37118
rect -1921 37114 -1710 37118
rect -1680 37116 -1672 37119
rect -1666 37117 -1658 37124
rect -2054 37112 -2046 37113
rect -2155 37106 -2139 37112
rect -2076 37106 -2046 37112
rect -2325 37094 -2314 37102
rect -2149 37096 -2139 37106
rect -2076 37096 -2054 37104
rect -2325 37074 -2320 37094
rect -2314 37086 -2306 37094
rect -2104 37091 -2054 37094
rect -2084 37088 -2054 37091
rect -2307 37078 -2306 37086
rect -2325 37070 -2314 37074
rect -2000 37070 -1992 37114
rect -1710 37112 -1702 37113
rect -1750 37106 -1702 37112
rect -1680 37108 -1665 37116
rect -1919 37104 -1916 37106
rect -1680 37104 -1672 37108
rect -1932 37102 -1916 37104
rect -1750 37096 -1710 37104
rect -1674 37096 -1666 37104
rect -1837 37088 -1789 37094
rect -1760 37092 -1692 37095
rect -1764 37088 -1692 37092
rect -1666 37088 -1658 37096
rect -1680 37080 -1665 37088
rect -1979 37070 -1945 37072
rect -1680 37070 -1672 37080
rect -1642 37070 -1637 37140
rect -1619 37070 -1614 37140
rect -1530 37070 -1526 37140
rect -1506 37070 -1502 37140
rect -1482 37070 -1478 37140
rect -1458 37070 -1454 37140
rect -1434 37070 -1430 37140
rect -1410 37070 -1406 37140
rect -1386 37070 -1382 37140
rect -1362 37070 -1358 37140
rect -1338 37070 -1334 37140
rect -1314 37070 -1310 37140
rect -1290 37070 -1286 37140
rect -1266 37070 -1262 37140
rect -1242 37070 -1238 37140
rect -1218 37070 -1214 37140
rect -1194 37070 -1190 37140
rect -1170 37070 -1166 37140
rect -1146 37070 -1142 37140
rect -1122 37070 -1118 37140
rect -1098 37070 -1094 37140
rect -1074 37070 -1070 37140
rect -1050 37070 -1046 37140
rect -1026 37070 -1022 37140
rect -1002 37070 -998 37140
rect -978 37070 -974 37140
rect -954 37070 -950 37140
rect -930 37070 -926 37140
rect -906 37091 -902 37140
rect -2393 37068 -909 37070
rect -2371 36926 -2366 37068
rect -2348 36926 -2343 37068
rect -2325 37058 -2314 37068
rect -2072 37060 -2046 37061
rect -2325 37042 -2320 37058
rect -2309 37046 -2298 37058
rect -2046 37055 -2040 37059
rect -2314 37042 -2309 37046
rect -2070 37043 -2046 37055
rect -2325 37030 -2314 37042
rect -2129 37039 -2111 37042
rect -2076 37041 -2070 37042
rect -2076 37039 -2046 37041
rect -2076 37037 -2070 37039
rect -2070 37034 -2046 37037
rect -2046 37032 -2040 37034
rect -2145 37030 -2129 37032
rect -2070 37030 -2040 37032
rect -2325 37014 -2320 37030
rect -2309 37018 -2298 37030
rect -2314 37014 -2309 37018
rect -2141 37016 -2129 37030
rect -2070 37016 -2046 37028
rect -2325 37002 -2314 37014
rect -2076 37012 -2046 37014
rect -2325 36982 -2320 37002
rect -2062 36982 -2032 36983
rect -2000 36982 -1992 37068
rect -1908 37066 -1894 37068
rect -1810 37060 -1799 37062
rect -1850 37055 -1802 37059
rect -1934 37050 -1923 37052
rect -1909 37050 -1898 37052
rect -1923 37042 -1919 37050
rect -1829 37043 -1802 37055
rect -1680 37042 -1672 37068
rect -1666 37060 -1665 37068
rect -1655 37048 -1650 37058
rect -1666 37042 -1655 37048
rect -1924 37026 -1919 37042
rect -1802 37041 -1781 37042
rect -1829 37039 -1781 37041
rect -1750 37039 -1702 37042
rect -1802 37037 -1794 37039
rect -1829 37034 -1802 37037
rect -1850 37032 -1829 37034
rect -1666 37032 -1665 37042
rect -1850 37030 -1802 37032
rect -1829 37016 -1802 37028
rect -1655 37020 -1650 37030
rect -1829 37012 -1792 37015
rect -1666 37014 -1655 37020
rect -1666 37004 -1665 37014
rect -1942 36984 -1937 36996
rect -1850 36993 -1822 36994
rect -1850 36989 -1802 36993
rect -2325 36974 -2317 36982
rect -2062 36980 -1961 36982
rect -2325 36954 -2320 36974
rect -2317 36966 -2309 36974
rect -2062 36967 -2040 36978
rect -2032 36973 -1961 36980
rect -1947 36974 -1942 36982
rect -1842 36980 -1794 36983
rect -2070 36962 -2022 36966
rect -2325 36942 -2317 36954
rect -2325 36926 -2320 36942
rect -2317 36938 -2309 36942
rect -2309 36926 -2301 36938
rect -2068 36931 -2038 36938
rect -2000 36928 -1992 36973
rect -1942 36972 -1937 36974
rect -1932 36964 -1927 36972
rect -1912 36969 -1896 36975
rect -1842 36967 -1802 36978
rect -1671 36974 -1663 36982
rect -1663 36966 -1655 36974
rect -1850 36962 -1680 36966
rect -1937 36948 -1934 36950
rect -1926 36948 -1921 36953
rect -1926 36943 -1924 36948
rect -1916 36940 -1914 36943
rect -1842 36940 -1794 36949
rect -1671 36942 -1663 36954
rect -1924 36930 -1916 36939
rect -1663 36938 -1655 36942
rect -1852 36931 -1804 36938
rect -1916 36929 -1914 36930
rect -2025 36927 -1991 36928
rect -2025 36926 -1975 36927
rect -1842 36926 -1804 36929
rect -1655 36926 -1647 36938
rect -1642 36926 -1637 37068
rect -1619 36926 -1614 37068
rect -1530 36926 -1526 37068
rect -1506 36926 -1502 37068
rect -1482 36926 -1478 37068
rect -1458 36926 -1454 37068
rect -1434 36926 -1430 37068
rect -1410 36926 -1406 37068
rect -1386 36926 -1382 37068
rect -1362 36926 -1358 37068
rect -1338 36926 -1334 37068
rect -1314 36926 -1310 37068
rect -1290 36926 -1286 37068
rect -1266 36926 -1262 37068
rect -1242 36926 -1238 37068
rect -1218 36926 -1214 37068
rect -1194 36926 -1190 37068
rect -1170 36926 -1166 37068
rect -1146 36926 -1142 37068
rect -1122 36926 -1118 37068
rect -1098 36926 -1094 37068
rect -1074 36926 -1070 37068
rect -1050 36926 -1046 37068
rect -1026 36926 -1022 37068
rect -1002 36926 -998 37068
rect -978 36926 -974 37068
rect -954 36926 -950 37068
rect -930 36926 -926 37068
rect -923 37067 -909 37068
rect -906 37067 -899 37091
rect -906 36926 -902 37067
rect -882 36926 -878 37140
rect -858 36926 -854 37140
rect -834 36926 -830 37140
rect -810 36926 -806 37140
rect -786 36926 -782 37140
rect -762 36926 -758 37140
rect -738 36926 -734 37140
rect -714 36926 -710 37140
rect -690 36926 -686 37140
rect -666 36926 -662 37140
rect -642 36926 -638 37140
rect -618 36926 -614 37140
rect -594 36926 -590 37140
rect -570 36926 -566 37140
rect -557 37013 -552 37023
rect -546 37013 -542 37140
rect -547 36999 -542 37013
rect -546 36926 -542 36999
rect -522 36947 -518 37140
rect -533 36926 -525 36927
rect -2393 36924 -525 36926
rect -2371 36902 -2366 36924
rect -2348 36902 -2343 36924
rect -2325 36914 -2317 36924
rect -2076 36914 -2068 36921
rect -2062 36914 -2001 36921
rect -2325 36902 -2320 36914
rect -2317 36910 -2309 36914
rect -2015 36913 -2001 36914
rect -2309 36902 -2301 36910
rect -2068 36904 -2062 36911
rect -2000 36906 -1992 36924
rect -1974 36922 -1960 36924
rect -1842 36923 -1804 36924
rect -1862 36921 -1794 36922
rect -1985 36919 -1794 36921
rect -1985 36914 -1852 36919
rect -1842 36913 -1794 36919
rect -1671 36914 -1663 36924
rect -2015 36904 -1985 36906
rect -1852 36904 -1804 36911
rect -1663 36910 -1655 36914
rect -2000 36902 -1992 36904
rect -1976 36902 -1940 36903
rect -1655 36902 -1647 36910
rect -1642 36902 -1637 36924
rect -1619 36902 -1614 36924
rect -1530 36902 -1526 36924
rect -1506 36902 -1502 36924
rect -1482 36902 -1478 36924
rect -1458 36902 -1454 36924
rect -1434 36902 -1430 36924
rect -1410 36902 -1406 36924
rect -1386 36902 -1382 36924
rect -1362 36902 -1358 36924
rect -1338 36903 -1334 36924
rect -1349 36902 -1315 36903
rect -2393 36900 -1315 36902
rect -2371 36830 -2366 36900
rect -2348 36830 -2343 36900
rect -2325 36898 -2320 36900
rect -2309 36898 -2301 36900
rect -2325 36886 -2317 36898
rect -2062 36887 -2032 36894
rect -2325 36866 -2320 36886
rect -2317 36882 -2309 36886
rect -2325 36858 -2317 36866
rect -2060 36860 -2030 36863
rect -2325 36838 -2320 36858
rect -2317 36850 -2309 36858
rect -2060 36847 -2038 36858
rect -2033 36851 -2030 36860
rect -2028 36856 -2027 36860
rect -2068 36842 -2038 36845
rect -2325 36830 -2317 36838
rect -2000 36830 -1992 36900
rect -1888 36895 -1874 36900
rect -1842 36896 -1804 36900
rect -1655 36898 -1647 36900
rect -1902 36893 -1874 36895
rect -1842 36886 -1794 36895
rect -1671 36886 -1663 36898
rect -1663 36882 -1655 36886
rect -1912 36875 -1884 36877
rect -1852 36869 -1804 36873
rect -1844 36860 -1796 36863
rect -1671 36858 -1663 36866
rect -1844 36847 -1804 36858
rect -1663 36850 -1655 36858
rect -1852 36842 -1680 36846
rect -1926 36830 -1892 36833
rect -1671 36830 -1663 36838
rect -1642 36830 -1637 36900
rect -1619 36830 -1614 36900
rect -1530 36830 -1526 36900
rect -1506 36830 -1502 36900
rect -1482 36830 -1478 36900
rect -1458 36830 -1454 36900
rect -1434 36830 -1430 36900
rect -1410 36830 -1406 36900
rect -1386 36830 -1382 36900
rect -1373 36869 -1368 36879
rect -1362 36869 -1358 36900
rect -1349 36893 -1344 36900
rect -1338 36893 -1334 36900
rect -1339 36879 -1334 36893
rect -1363 36855 -1358 36869
rect -1362 36830 -1358 36855
rect -1338 36830 -1334 36879
rect -1314 36830 -1310 36924
rect -1290 36830 -1286 36924
rect -1266 36830 -1262 36924
rect -1242 36830 -1238 36924
rect -1218 36830 -1214 36924
rect -1194 36830 -1190 36924
rect -1170 36830 -1166 36924
rect -1146 36830 -1142 36924
rect -1122 36830 -1118 36924
rect -1098 36830 -1094 36924
rect -1074 36830 -1070 36924
rect -1050 36830 -1046 36924
rect -1026 36830 -1022 36924
rect -1002 36830 -998 36924
rect -978 36830 -974 36924
rect -954 36830 -950 36924
rect -930 36830 -926 36924
rect -906 36830 -902 36924
rect -882 36830 -878 36924
rect -858 36830 -854 36924
rect -834 36830 -830 36924
rect -810 36830 -806 36924
rect -786 36830 -782 36924
rect -762 36830 -758 36924
rect -738 36830 -734 36924
rect -714 36830 -710 36924
rect -690 36830 -686 36924
rect -666 36830 -662 36924
rect -642 36830 -638 36924
rect -618 36830 -614 36924
rect -594 36830 -590 36924
rect -570 36830 -566 36924
rect -546 36830 -542 36924
rect -539 36923 -525 36924
rect -522 36923 -515 36947
rect -533 36917 -528 36923
rect -522 36917 -518 36923
rect -523 36903 -518 36917
rect -522 36830 -518 36903
rect -498 36851 -494 37140
rect -2393 36828 -501 36830
rect -2371 36806 -2366 36828
rect -2348 36806 -2343 36828
rect -2325 36822 -2317 36828
rect -2325 36806 -2320 36822
rect -2309 36810 -2301 36822
rect -2068 36811 -2038 36818
rect -2317 36806 -2309 36810
rect -2000 36808 -1992 36828
rect -1844 36820 -1794 36828
rect -1671 36822 -1663 36828
rect -1852 36811 -1804 36818
rect -1655 36810 -1647 36822
rect -2025 36807 -1991 36808
rect -2025 36806 -1975 36807
rect -1844 36806 -1804 36809
rect -1663 36806 -1655 36810
rect -1642 36806 -1637 36828
rect -1619 36806 -1614 36828
rect -1530 36806 -1526 36828
rect -1506 36806 -1502 36828
rect -1482 36806 -1478 36828
rect -1458 36806 -1454 36828
rect -1434 36806 -1430 36828
rect -1410 36806 -1406 36828
rect -1386 36806 -1382 36828
rect -1362 36806 -1358 36828
rect -1338 36806 -1334 36828
rect -1314 36827 -1310 36828
rect -2393 36804 -1317 36806
rect -2371 36782 -2366 36804
rect -2348 36782 -2343 36804
rect -2325 36794 -2317 36804
rect -2060 36794 -2020 36801
rect -2004 36796 -2001 36801
rect -2015 36794 -2001 36796
rect -2000 36794 -1992 36804
rect -1972 36802 -1958 36804
rect -1844 36803 -1804 36804
rect -1862 36801 -1796 36802
rect -1985 36799 -1796 36801
rect -1985 36794 -1852 36799
rect -2325 36782 -2320 36794
rect -2309 36782 -2301 36794
rect -2068 36784 -2060 36791
rect -2015 36784 -1990 36794
rect -1844 36793 -1796 36799
rect -1671 36794 -1663 36804
rect -1852 36784 -1804 36791
rect -2020 36782 -2004 36784
rect -2000 36782 -1992 36784
rect -1976 36782 -1940 36783
rect -1655 36782 -1647 36794
rect -1642 36782 -1637 36804
rect -1619 36782 -1614 36804
rect -1530 36782 -1526 36804
rect -1506 36782 -1502 36804
rect -1482 36782 -1478 36804
rect -1458 36782 -1454 36804
rect -1434 36782 -1430 36804
rect -1410 36782 -1406 36804
rect -1386 36782 -1382 36804
rect -1362 36782 -1358 36804
rect -1338 36803 -1334 36804
rect -1331 36803 -1317 36804
rect -1314 36803 -1307 36827
rect -2393 36780 -1341 36782
rect -2371 36710 -2366 36780
rect -2348 36710 -2343 36780
rect -2325 36778 -2320 36780
rect -2317 36778 -2309 36780
rect -2325 36766 -2317 36778
rect -2060 36767 -2030 36774
rect -2325 36746 -2320 36766
rect -2325 36738 -2317 36746
rect -2060 36740 -2030 36743
rect -2325 36710 -2320 36738
rect -2317 36730 -2309 36738
rect -2060 36727 -2038 36738
rect -2033 36731 -2030 36740
rect -2028 36736 -2027 36740
rect -2068 36722 -2038 36725
rect -2000 36710 -1992 36780
rect -1844 36776 -1804 36780
rect -1663 36778 -1655 36780
rect -1844 36766 -1794 36775
rect -1671 36766 -1663 36778
rect -1912 36755 -1884 36757
rect -1852 36749 -1804 36753
rect -1844 36740 -1796 36743
rect -1671 36738 -1663 36746
rect -1844 36727 -1804 36738
rect -1663 36730 -1655 36738
rect -1852 36722 -1680 36726
rect -1642 36710 -1637 36780
rect -1619 36710 -1614 36780
rect -1530 36710 -1526 36780
rect -1506 36710 -1502 36780
rect -1482 36710 -1478 36780
rect -1458 36710 -1454 36780
rect -1434 36710 -1430 36780
rect -1410 36710 -1406 36780
rect -1386 36710 -1382 36780
rect -1362 36710 -1358 36780
rect -1355 36779 -1341 36780
rect -1338 36779 -1331 36803
rect -1338 36710 -1334 36779
rect -1314 36710 -1310 36803
rect -1290 36710 -1286 36828
rect -1266 36710 -1262 36828
rect -1242 36710 -1238 36828
rect -1218 36710 -1214 36828
rect -1194 36710 -1190 36828
rect -1170 36710 -1166 36828
rect -1146 36710 -1142 36828
rect -1122 36710 -1118 36828
rect -1098 36710 -1094 36828
rect -1074 36710 -1070 36828
rect -1050 36710 -1046 36828
rect -1026 36710 -1022 36828
rect -1002 36710 -998 36828
rect -978 36710 -974 36828
rect -954 36710 -950 36828
rect -930 36710 -926 36828
rect -906 36710 -902 36828
rect -882 36710 -878 36828
rect -858 36710 -854 36828
rect -834 36710 -830 36828
rect -810 36710 -806 36828
rect -786 36710 -782 36828
rect -762 36710 -758 36828
rect -738 36710 -734 36828
rect -714 36710 -710 36828
rect -690 36710 -686 36828
rect -666 36710 -662 36828
rect -642 36710 -638 36828
rect -618 36710 -614 36828
rect -594 36710 -590 36828
rect -570 36710 -566 36828
rect -546 36710 -542 36828
rect -522 36710 -518 36828
rect -515 36827 -501 36828
rect -498 36827 -491 36851
rect -498 36735 -494 36827
rect -509 36734 -475 36735
rect -474 36734 -470 37140
rect -450 36734 -446 37140
rect -426 36734 -422 37140
rect -402 36734 -398 37140
rect -389 37085 -384 37095
rect -378 37085 -374 37140
rect -379 37071 -374 37085
rect -389 37061 -384 37071
rect -379 37047 -374 37061
rect -378 36734 -374 37047
rect -354 37019 -350 37140
rect -354 36998 -347 37019
rect -330 36998 -326 37140
rect -306 36998 -302 37140
rect -282 36998 -278 37140
rect -258 36998 -254 37140
rect -234 36998 -230 37140
rect -210 36998 -206 37140
rect -186 36998 -182 37140
rect -162 36998 -158 37140
rect -138 36998 -134 37140
rect -114 36998 -110 37140
rect -90 36998 -86 37140
rect -66 36998 -62 37140
rect -42 36998 -38 37140
rect -18 36998 -14 37140
rect 6 36998 10 37140
rect 30 36998 34 37140
rect 54 36998 58 37140
rect 78 36998 82 37140
rect 102 36998 106 37140
rect 126 36998 130 37140
rect 150 36998 154 37140
rect 174 36998 178 37140
rect 198 36998 202 37140
rect 222 36998 226 37140
rect 246 36998 250 37140
rect 270 36998 274 37140
rect 283 37133 288 37140
rect 294 37133 298 37140
rect 293 37119 298 37133
rect 294 36998 298 37119
rect 318 37067 322 37595
rect 318 37043 325 37067
rect 318 36998 322 37043
rect 342 36998 346 37740
rect 366 37527 370 37740
rect 355 37526 389 37527
rect 390 37526 394 37740
rect 414 37526 418 37740
rect 438 37526 442 37740
rect 462 37526 466 37740
rect 486 37526 490 37740
rect 510 37526 514 37740
rect 534 37526 538 37740
rect 558 37526 562 37740
rect 582 37526 586 37740
rect 606 37526 610 37740
rect 630 37526 634 37740
rect 654 37526 658 37740
rect 678 37526 682 37740
rect 702 37526 706 37740
rect 726 37526 730 37740
rect 750 37526 754 37740
rect 774 37526 778 37740
rect 798 37526 802 37740
rect 822 37526 826 37740
rect 846 37526 850 37740
rect 870 37526 874 37740
rect 894 37526 898 37740
rect 918 37526 922 37740
rect 942 37526 946 37740
rect 966 37526 970 37740
rect 990 37526 994 37740
rect 1014 37526 1018 37740
rect 1038 37647 1042 37740
rect 1027 37646 1061 37647
rect 1062 37646 1066 37740
rect 1086 37646 1090 37740
rect 1110 37646 1114 37740
rect 1134 37646 1138 37740
rect 1141 37739 1155 37740
rect 1147 37733 1152 37739
rect 1157 37719 1162 37733
rect 1147 37661 1152 37671
rect 1158 37661 1162 37719
rect 1157 37647 1162 37661
rect 1171 37657 1179 37661
rect 1165 37647 1171 37657
rect 1147 37646 1179 37647
rect 1027 37644 1179 37646
rect 1027 37637 1032 37644
rect 1038 37637 1042 37644
rect 1037 37623 1042 37637
rect 1027 37613 1032 37623
rect 1037 37599 1042 37613
rect 1038 37526 1042 37599
rect 1062 37571 1066 37644
rect 355 37524 1059 37526
rect 355 37517 360 37524
rect 366 37517 370 37524
rect 365 37503 370 37517
rect 355 37493 360 37503
rect 365 37479 370 37493
rect 366 36998 370 37479
rect 390 37451 394 37524
rect 390 37430 397 37451
rect 414 37430 418 37524
rect 438 37430 442 37524
rect 462 37430 466 37524
rect 486 37430 490 37524
rect 510 37430 514 37524
rect 534 37430 538 37524
rect 558 37430 562 37524
rect 582 37430 586 37524
rect 606 37430 610 37524
rect 630 37430 634 37524
rect 654 37431 658 37524
rect 643 37430 677 37431
rect 373 37428 677 37430
rect 373 37427 387 37428
rect 390 37403 397 37428
rect 390 36998 394 37403
rect 414 36998 418 37428
rect 438 36998 442 37428
rect 462 36998 466 37428
rect 486 36998 490 37428
rect 510 36998 514 37428
rect 523 37373 528 37383
rect 534 37373 538 37428
rect 533 37359 538 37373
rect 523 37349 528 37359
rect 533 37335 538 37349
rect 534 36998 538 37335
rect 558 37307 562 37428
rect 558 37259 565 37307
rect 558 36998 562 37259
rect 582 36998 586 37428
rect 606 36998 610 37428
rect 630 36998 634 37428
rect 643 37421 648 37428
rect 654 37421 658 37428
rect 653 37407 658 37421
rect 654 36998 658 37407
rect 678 37355 682 37524
rect 678 37331 685 37355
rect 678 36998 682 37331
rect 702 36998 706 37524
rect 726 36998 730 37524
rect 750 36998 754 37524
rect 774 36998 778 37524
rect 798 36998 802 37524
rect 822 36998 826 37524
rect 846 36998 850 37524
rect 870 36998 874 37524
rect 894 36998 898 37524
rect 918 36998 922 37524
rect 942 36998 946 37524
rect 966 36998 970 37524
rect 990 36998 994 37524
rect 1003 37253 1008 37263
rect 1014 37253 1018 37524
rect 1013 37239 1018 37253
rect 1003 37229 1008 37239
rect 1013 37215 1018 37229
rect 1014 36998 1018 37215
rect 1038 37187 1042 37524
rect 1045 37523 1059 37524
rect 1062 37523 1069 37571
rect 1038 37139 1045 37187
rect 1038 36998 1042 37139
rect 1062 36998 1066 37523
rect 1086 36998 1090 37644
rect 1110 36998 1114 37644
rect 1134 36998 1138 37644
rect 1147 37637 1152 37644
rect 1165 37643 1179 37644
rect 1157 37623 1162 37637
rect 1158 36998 1162 37623
rect 1171 37517 1176 37527
rect 1181 37503 1186 37517
rect 1182 36998 1186 37503
rect 1195 37373 1200 37383
rect 1205 37359 1210 37373
rect 1206 36998 1210 37359
rect 1219 37253 1224 37263
rect 1229 37239 1234 37253
rect 1219 37205 1224 37215
rect 1230 37205 1234 37239
rect 1229 37191 1234 37205
rect 1219 37085 1224 37095
rect 1229 37071 1234 37085
rect 1230 36999 1234 37071
rect 1219 36998 1251 36999
rect -371 36996 1251 36998
rect -371 36995 -357 36996
rect -354 36971 -347 36996
rect -354 36734 -350 36971
rect -330 36734 -326 36996
rect -306 36734 -302 36996
rect -282 36734 -278 36996
rect -258 36734 -254 36996
rect -234 36734 -230 36996
rect -210 36734 -206 36996
rect -186 36734 -182 36996
rect -162 36734 -158 36996
rect -138 36734 -134 36996
rect -114 36734 -110 36996
rect -90 36734 -86 36996
rect -66 36855 -62 36996
rect -77 36854 -43 36855
rect -42 36854 -38 36996
rect -18 36854 -14 36996
rect 6 36854 10 36996
rect 30 36854 34 36996
rect 54 36854 58 36996
rect 78 36854 82 36996
rect 102 36854 106 36996
rect 126 36854 130 36996
rect 150 36854 154 36996
rect 174 36854 178 36996
rect 198 36854 202 36996
rect 222 36854 226 36996
rect 246 36854 250 36996
rect 270 36854 274 36996
rect 294 36854 298 36996
rect 318 36854 322 36996
rect 342 36854 346 36996
rect 366 36854 370 36996
rect 390 36854 394 36996
rect 414 36854 418 36996
rect 438 36854 442 36996
rect 462 36854 466 36996
rect 486 36854 490 36996
rect 510 36854 514 36996
rect 534 36854 538 36996
rect 558 36854 562 36996
rect 582 36854 586 36996
rect 606 36854 610 36996
rect 630 36854 634 36996
rect 654 36854 658 36996
rect 667 36965 672 36975
rect 678 36965 682 36996
rect 677 36951 682 36965
rect 667 36941 672 36951
rect 677 36927 682 36941
rect 678 36854 682 36927
rect 702 36899 706 36996
rect -77 36852 699 36854
rect -77 36845 -72 36852
rect -66 36845 -62 36852
rect -67 36831 -62 36845
rect -77 36821 -72 36831
rect -67 36807 -62 36821
rect -66 36734 -62 36807
rect -42 36779 -38 36852
rect -42 36758 -35 36779
rect -18 36758 -14 36852
rect 6 36758 10 36852
rect 30 36758 34 36852
rect 54 36758 58 36852
rect 78 36758 82 36852
rect 102 36758 106 36852
rect 126 36758 130 36852
rect 150 36758 154 36852
rect 174 36758 178 36852
rect 198 36758 202 36852
rect 222 36758 226 36852
rect 246 36758 250 36852
rect 270 36758 274 36852
rect 294 36758 298 36852
rect 318 36758 322 36852
rect 342 36758 346 36852
rect 366 36758 370 36852
rect 390 36758 394 36852
rect 414 36758 418 36852
rect 438 36758 442 36852
rect 462 36758 466 36852
rect 486 36758 490 36852
rect 510 36758 514 36852
rect 534 36758 538 36852
rect 558 36758 562 36852
rect 582 36758 586 36852
rect 606 36758 610 36852
rect 630 36758 634 36852
rect 654 36758 658 36852
rect 678 36758 682 36852
rect 685 36851 699 36852
rect 702 36851 709 36899
rect 702 36758 706 36851
rect 726 36758 730 36996
rect 750 36758 754 36996
rect 774 36758 778 36996
rect 798 36758 802 36996
rect 822 36758 826 36996
rect 846 36758 850 36996
rect 870 36758 874 36996
rect 894 36758 898 36996
rect 918 36758 922 36996
rect 942 36758 946 36996
rect 966 36758 970 36996
rect 990 36758 994 36996
rect 1014 36758 1018 36996
rect 1038 36758 1042 36996
rect 1062 36758 1066 36996
rect 1086 36758 1090 36996
rect 1110 36758 1114 36996
rect 1134 36758 1138 36996
rect 1158 36758 1162 36996
rect 1182 36758 1186 36996
rect 1206 36759 1210 36996
rect 1219 36989 1224 36996
rect 1230 36989 1234 36996
rect 1237 36995 1251 36996
rect 1229 36975 1234 36989
rect 1219 36965 1224 36975
rect 1229 36951 1234 36965
rect 1219 36773 1224 36783
rect 1230 36773 1234 36951
rect 1243 36845 1248 36855
rect 1253 36831 1258 36845
rect 1243 36797 1248 36807
rect 1254 36797 1258 36831
rect 1253 36783 1258 36797
rect 1229 36759 1234 36773
rect 1195 36758 1229 36759
rect -59 36756 1229 36758
rect -59 36755 -45 36756
rect -509 36732 -45 36734
rect -509 36725 -504 36732
rect -498 36725 -494 36732
rect -499 36711 -494 36725
rect -509 36710 -475 36711
rect -2393 36708 -475 36710
rect -2371 36686 -2366 36708
rect -2348 36686 -2343 36708
rect -2325 36686 -2320 36708
rect -2309 36690 -2301 36700
rect -2068 36691 -2062 36696
rect -2317 36686 -2309 36690
rect -2060 36686 -2050 36691
rect -2000 36686 -1992 36708
rect -1806 36700 -1680 36706
rect -1854 36691 -1806 36696
rect -1655 36690 -1647 36700
rect -1972 36686 -1964 36687
rect -1958 36686 -1942 36688
rect -1844 36686 -1806 36689
rect -1663 36686 -1655 36690
rect -1642 36686 -1637 36708
rect -1619 36686 -1614 36708
rect -1530 36686 -1526 36708
rect -1506 36686 -1502 36708
rect -1482 36686 -1478 36708
rect -1458 36686 -1454 36708
rect -1434 36686 -1430 36708
rect -1410 36686 -1406 36708
rect -1386 36686 -1382 36708
rect -1362 36686 -1358 36708
rect -1338 36686 -1334 36708
rect -1314 36686 -1310 36708
rect -1290 36686 -1286 36708
rect -1266 36686 -1262 36708
rect -1242 36686 -1238 36708
rect -1218 36686 -1214 36708
rect -1194 36686 -1190 36708
rect -1170 36686 -1166 36708
rect -1146 36686 -1142 36708
rect -1122 36686 -1118 36708
rect -1098 36686 -1094 36708
rect -1074 36686 -1070 36708
rect -1050 36686 -1046 36708
rect -1026 36686 -1022 36708
rect -1002 36686 -998 36708
rect -978 36686 -974 36708
rect -954 36686 -950 36708
rect -930 36686 -926 36708
rect -906 36686 -902 36708
rect -882 36686 -878 36708
rect -858 36686 -854 36708
rect -834 36686 -830 36708
rect -810 36686 -806 36708
rect -786 36686 -782 36708
rect -762 36686 -758 36708
rect -738 36686 -734 36708
rect -714 36686 -710 36708
rect -690 36686 -686 36708
rect -666 36686 -662 36708
rect -642 36686 -638 36708
rect -618 36686 -614 36708
rect -594 36686 -590 36708
rect -570 36686 -566 36708
rect -546 36687 -542 36708
rect -557 36686 -523 36687
rect -2393 36684 -523 36686
rect -2371 36662 -2366 36684
rect -2348 36662 -2343 36684
rect -2325 36662 -2320 36684
rect -2060 36678 -2050 36684
rect -2309 36662 -2301 36672
rect -2060 36671 -2030 36678
rect -2000 36674 -1992 36684
rect -1972 36682 -1942 36684
rect -1958 36681 -1942 36682
rect -1844 36680 -1806 36684
rect -2068 36664 -2062 36671
rect -2062 36662 -2036 36664
rect -2393 36660 -2036 36662
rect -2030 36662 -2012 36664
rect -2004 36662 -1990 36674
rect -1844 36673 -1798 36678
rect -1806 36671 -1798 36673
rect -1854 36669 -1844 36671
rect -1854 36664 -1806 36669
rect -1864 36662 -1796 36663
rect -1655 36662 -1647 36672
rect -1642 36662 -1637 36684
rect -1619 36662 -1614 36684
rect -1530 36662 -1526 36684
rect -1506 36662 -1502 36684
rect -1482 36662 -1478 36684
rect -1458 36662 -1454 36684
rect -1434 36662 -1430 36684
rect -1410 36662 -1406 36684
rect -1386 36662 -1382 36684
rect -1362 36662 -1358 36684
rect -1338 36662 -1334 36684
rect -1314 36662 -1310 36684
rect -1290 36662 -1286 36684
rect -1266 36662 -1262 36684
rect -1242 36662 -1238 36684
rect -1218 36662 -1214 36684
rect -1194 36662 -1190 36684
rect -1170 36662 -1166 36684
rect -1146 36662 -1142 36684
rect -1122 36662 -1118 36684
rect -1098 36662 -1094 36684
rect -1074 36662 -1070 36684
rect -1050 36663 -1046 36684
rect -1061 36662 -1027 36663
rect -2030 36660 -1027 36662
rect -2371 36614 -2366 36660
rect -2348 36614 -2343 36660
rect -2325 36614 -2320 36660
rect -2317 36656 -2309 36660
rect -2060 36656 -2050 36660
rect -2060 36654 -2036 36656
rect -2060 36652 -2030 36654
rect -2292 36646 -2030 36652
rect -2092 36630 -2062 36632
rect -2094 36626 -2062 36630
rect -2000 36614 -1992 36660
rect -1844 36653 -1806 36660
rect -1663 36656 -1655 36660
rect -1844 36646 -1680 36652
rect -1854 36630 -1806 36632
rect -1854 36626 -1680 36630
rect -1926 36614 -1892 36617
rect -1642 36614 -1637 36660
rect -1619 36614 -1614 36660
rect -1530 36614 -1526 36660
rect -1506 36614 -1502 36660
rect -1482 36614 -1478 36660
rect -1458 36614 -1454 36660
rect -1434 36614 -1430 36660
rect -1410 36614 -1406 36660
rect -1386 36614 -1382 36660
rect -1362 36614 -1358 36660
rect -1338 36614 -1334 36660
rect -1314 36614 -1310 36660
rect -1290 36614 -1286 36660
rect -1266 36614 -1262 36660
rect -1242 36614 -1238 36660
rect -1218 36614 -1214 36660
rect -1194 36614 -1190 36660
rect -1170 36614 -1166 36660
rect -1146 36614 -1142 36660
rect -1122 36614 -1118 36660
rect -1098 36614 -1094 36660
rect -1074 36614 -1070 36660
rect -1061 36653 -1056 36660
rect -1050 36653 -1046 36660
rect -1051 36639 -1046 36653
rect -1061 36629 -1056 36639
rect -1050 36629 -1046 36639
rect -1051 36615 -1046 36629
rect -1061 36614 -1027 36615
rect -2393 36612 -1027 36614
rect -2371 36590 -2366 36612
rect -2348 36590 -2343 36612
rect -2325 36590 -2320 36612
rect -2054 36611 -1906 36612
rect -2054 36610 -2036 36611
rect -2309 36596 -2301 36606
rect -2317 36590 -2309 36596
rect -2068 36595 -2038 36602
rect -2000 36594 -1992 36611
rect -1920 36610 -1906 36611
rect -1846 36604 -1794 36612
rect -1852 36597 -1804 36602
rect -1902 36595 -1804 36597
rect -1655 36596 -1647 36606
rect -2000 36592 -1975 36594
rect -1902 36593 -1852 36595
rect -2025 36590 -1975 36592
rect -1846 36590 -1804 36593
rect -1663 36590 -1655 36596
rect -1642 36590 -1637 36612
rect -1619 36590 -1614 36612
rect -1530 36590 -1526 36612
rect -1506 36590 -1502 36612
rect -1482 36590 -1478 36612
rect -1458 36590 -1454 36612
rect -1434 36590 -1430 36612
rect -1410 36590 -1406 36612
rect -1386 36590 -1382 36612
rect -1362 36590 -1358 36612
rect -1338 36590 -1334 36612
rect -1314 36590 -1310 36612
rect -1290 36590 -1286 36612
rect -1266 36590 -1262 36612
rect -1242 36591 -1238 36612
rect -1253 36590 -1219 36591
rect -2393 36588 -1219 36590
rect -2371 36566 -2366 36588
rect -2348 36566 -2343 36588
rect -2325 36566 -2320 36588
rect -2054 36587 -2038 36588
rect -2000 36587 -1966 36588
rect -1846 36587 -1804 36588
rect -2000 36586 -1975 36587
rect -2076 36578 -2054 36585
rect -2309 36568 -2301 36578
rect -2044 36575 -2038 36580
rect -2028 36578 -2001 36585
rect -2054 36568 -2038 36575
rect -2015 36577 -2001 36578
rect -2015 36568 -2014 36577
rect -2317 36566 -2309 36568
rect -2044 36566 -2028 36568
rect -2000 36566 -1992 36586
rect -1982 36585 -1975 36586
rect -1862 36585 -1798 36586
rect -1985 36578 -1796 36585
rect -1862 36577 -1798 36578
rect -1852 36568 -1804 36575
rect -1655 36568 -1647 36578
rect -1976 36566 -1940 36567
rect -1663 36566 -1655 36568
rect -1642 36566 -1637 36588
rect -1619 36566 -1614 36588
rect -1530 36566 -1526 36588
rect -1506 36566 -1502 36588
rect -1482 36566 -1478 36588
rect -1458 36566 -1454 36588
rect -1434 36566 -1430 36588
rect -1410 36566 -1406 36588
rect -1386 36566 -1382 36588
rect -1362 36566 -1358 36588
rect -1338 36566 -1334 36588
rect -1314 36566 -1310 36588
rect -1290 36566 -1286 36588
rect -1266 36566 -1262 36588
rect -1253 36581 -1248 36588
rect -1242 36581 -1238 36588
rect -1243 36567 -1238 36581
rect -1242 36566 -1238 36567
rect -1218 36566 -1214 36612
rect -1194 36566 -1190 36612
rect -1170 36566 -1166 36612
rect -1146 36566 -1142 36612
rect -1122 36566 -1118 36612
rect -1098 36566 -1094 36612
rect -1074 36566 -1070 36612
rect -1061 36605 -1056 36612
rect -1051 36591 -1046 36605
rect -1050 36566 -1046 36591
rect -1026 36587 -1022 36684
rect -2393 36564 -1029 36566
rect -2371 36494 -2366 36564
rect -2348 36494 -2343 36564
rect -2325 36530 -2320 36564
rect -2317 36562 -2309 36564
rect -2076 36551 -2054 36558
rect -2325 36522 -2317 36530
rect -2060 36524 -2030 36527
rect -2325 36494 -2320 36522
rect -2317 36514 -2309 36522
rect -2060 36511 -2038 36522
rect -2033 36515 -2030 36524
rect -2028 36520 -2027 36524
rect -2068 36506 -2038 36509
rect -2000 36494 -1992 36564
rect -1846 36560 -1804 36564
rect -1663 36562 -1655 36564
rect -1846 36550 -1794 36559
rect -1912 36539 -1884 36541
rect -1852 36533 -1804 36537
rect -1844 36524 -1796 36527
rect -1671 36522 -1663 36530
rect -1844 36511 -1804 36522
rect -1663 36514 -1655 36522
rect -1852 36506 -1680 36510
rect -1642 36494 -1637 36564
rect -1619 36494 -1614 36564
rect -1530 36494 -1526 36564
rect -1506 36494 -1502 36564
rect -1482 36494 -1478 36564
rect -1458 36494 -1454 36564
rect -1434 36494 -1430 36564
rect -1410 36494 -1406 36564
rect -1386 36494 -1382 36564
rect -1362 36494 -1358 36564
rect -1338 36494 -1334 36564
rect -1314 36494 -1310 36564
rect -1290 36494 -1286 36564
rect -1266 36494 -1262 36564
rect -1242 36494 -1238 36564
rect -1218 36515 -1214 36564
rect -2393 36492 -1221 36494
rect -2371 36470 -2366 36492
rect -2348 36470 -2343 36492
rect -2325 36470 -2320 36492
rect -2309 36474 -2301 36484
rect -2068 36475 -2062 36480
rect -2317 36470 -2309 36474
rect -2060 36470 -2050 36475
rect -2000 36470 -1992 36492
rect -1806 36484 -1680 36490
rect -1854 36475 -1806 36480
rect -1655 36474 -1647 36484
rect -1972 36470 -1964 36471
rect -1958 36470 -1942 36472
rect -1844 36470 -1806 36473
rect -1663 36470 -1655 36474
rect -1642 36470 -1637 36492
rect -1619 36470 -1614 36492
rect -1530 36470 -1526 36492
rect -1506 36470 -1502 36492
rect -1482 36470 -1478 36492
rect -1458 36470 -1454 36492
rect -1434 36470 -1430 36492
rect -1410 36470 -1406 36492
rect -1386 36470 -1382 36492
rect -1362 36470 -1358 36492
rect -1338 36470 -1334 36492
rect -1314 36470 -1310 36492
rect -1290 36470 -1286 36492
rect -1266 36470 -1262 36492
rect -1242 36470 -1238 36492
rect -1235 36491 -1221 36492
rect -1218 36491 -1211 36515
rect -1218 36470 -1214 36491
rect -1194 36470 -1190 36564
rect -1170 36470 -1166 36564
rect -1146 36470 -1142 36564
rect -1122 36470 -1118 36564
rect -1098 36470 -1094 36564
rect -1074 36470 -1070 36564
rect -1050 36470 -1046 36564
rect -1043 36563 -1029 36564
rect -1026 36542 -1019 36587
rect -1002 36542 -998 36684
rect -978 36542 -974 36684
rect -954 36542 -950 36684
rect -930 36542 -926 36684
rect -906 36542 -902 36684
rect -882 36542 -878 36684
rect -858 36542 -854 36684
rect -834 36542 -830 36684
rect -810 36542 -806 36684
rect -786 36542 -782 36684
rect -762 36542 -758 36684
rect -738 36542 -734 36684
rect -714 36542 -710 36684
rect -690 36542 -686 36684
rect -666 36542 -662 36684
rect -642 36542 -638 36684
rect -618 36542 -614 36684
rect -594 36542 -590 36684
rect -570 36542 -566 36684
rect -557 36677 -552 36684
rect -546 36677 -542 36684
rect -547 36663 -542 36677
rect -546 36542 -542 36663
rect -522 36611 -518 36708
rect -509 36701 -504 36708
rect -499 36687 -494 36701
rect -522 36587 -515 36611
rect -522 36542 -518 36587
rect -498 36542 -494 36687
rect -474 36659 -470 36732
rect -474 36638 -467 36659
rect -450 36638 -446 36732
rect -426 36638 -422 36732
rect -402 36638 -398 36732
rect -378 36638 -374 36732
rect -354 36638 -350 36732
rect -330 36638 -326 36732
rect -306 36638 -302 36732
rect -282 36638 -278 36732
rect -258 36638 -254 36732
rect -234 36638 -230 36732
rect -210 36638 -206 36732
rect -186 36638 -182 36732
rect -162 36638 -158 36732
rect -138 36638 -134 36732
rect -114 36638 -110 36732
rect -90 36638 -86 36732
rect -66 36638 -62 36732
rect -59 36731 -45 36732
rect -42 36731 -35 36756
rect -42 36638 -38 36731
rect -18 36638 -14 36756
rect 6 36638 10 36756
rect 30 36638 34 36756
rect 54 36638 58 36756
rect 78 36638 82 36756
rect 102 36638 106 36756
rect 126 36638 130 36756
rect 150 36638 154 36756
rect 174 36638 178 36756
rect 198 36638 202 36756
rect 222 36638 226 36756
rect 246 36638 250 36756
rect 270 36638 274 36756
rect 294 36638 298 36756
rect 318 36638 322 36756
rect 342 36638 346 36756
rect 366 36638 370 36756
rect 390 36638 394 36756
rect 414 36638 418 36756
rect 438 36638 442 36756
rect 462 36638 466 36756
rect 486 36638 490 36756
rect 510 36638 514 36756
rect 534 36638 538 36756
rect 558 36638 562 36756
rect 582 36638 586 36756
rect 606 36638 610 36756
rect 630 36638 634 36756
rect 654 36638 658 36756
rect 678 36638 682 36756
rect 702 36638 706 36756
rect 726 36638 730 36756
rect 750 36638 754 36756
rect 774 36638 778 36756
rect 798 36638 802 36756
rect 822 36638 826 36756
rect 846 36638 850 36756
rect 870 36638 874 36756
rect 894 36638 898 36756
rect 918 36638 922 36756
rect 942 36638 946 36756
rect 966 36638 970 36756
rect 990 36638 994 36756
rect 1014 36638 1018 36756
rect 1038 36638 1042 36756
rect 1062 36638 1066 36756
rect 1086 36638 1090 36756
rect 1110 36638 1114 36756
rect 1134 36638 1138 36756
rect 1158 36638 1162 36756
rect 1182 36638 1186 36756
rect 1195 36749 1200 36756
rect 1206 36749 1210 36756
rect 1205 36735 1210 36749
rect 1195 36725 1200 36735
rect 1205 36711 1210 36725
rect 1206 36638 1210 36711
rect 1219 36638 1227 36639
rect -491 36636 1227 36638
rect -491 36635 -477 36636
rect -474 36611 -467 36636
rect -474 36542 -470 36611
rect -450 36542 -446 36636
rect -426 36542 -422 36636
rect -402 36542 -398 36636
rect -378 36542 -374 36636
rect -354 36542 -350 36636
rect -330 36542 -326 36636
rect -306 36542 -302 36636
rect -282 36542 -278 36636
rect -258 36542 -254 36636
rect -234 36542 -230 36636
rect -210 36542 -206 36636
rect -186 36542 -182 36636
rect -162 36542 -158 36636
rect -138 36542 -134 36636
rect -114 36542 -110 36636
rect -90 36542 -86 36636
rect -66 36542 -62 36636
rect -42 36542 -38 36636
rect -18 36542 -14 36636
rect 6 36542 10 36636
rect 30 36542 34 36636
rect 54 36542 58 36636
rect 78 36542 82 36636
rect 102 36542 106 36636
rect 126 36542 130 36636
rect 150 36542 154 36636
rect 174 36542 178 36636
rect 198 36542 202 36636
rect 222 36542 226 36636
rect 246 36542 250 36636
rect 270 36542 274 36636
rect 294 36542 298 36636
rect 318 36542 322 36636
rect 342 36542 346 36636
rect 366 36542 370 36636
rect 379 36557 384 36567
rect 390 36557 394 36636
rect 389 36543 394 36557
rect 390 36542 394 36543
rect 414 36542 418 36636
rect 438 36543 442 36636
rect 427 36542 461 36543
rect -1043 36540 461 36542
rect -1043 36539 -1029 36540
rect -1026 36515 -1019 36540
rect -1026 36470 -1022 36515
rect -1002 36470 -998 36540
rect -978 36470 -974 36540
rect -954 36470 -950 36540
rect -930 36470 -926 36540
rect -906 36470 -902 36540
rect -882 36470 -878 36540
rect -858 36470 -854 36540
rect -834 36470 -830 36540
rect -810 36470 -806 36540
rect -786 36470 -782 36540
rect -762 36470 -758 36540
rect -738 36470 -734 36540
rect -714 36470 -710 36540
rect -690 36470 -686 36540
rect -666 36470 -662 36540
rect -642 36470 -638 36540
rect -618 36470 -614 36540
rect -594 36470 -590 36540
rect -570 36470 -566 36540
rect -546 36470 -542 36540
rect -522 36470 -518 36540
rect -498 36470 -494 36540
rect -474 36470 -470 36540
rect -450 36470 -446 36540
rect -426 36470 -422 36540
rect -413 36509 -408 36519
rect -402 36509 -398 36540
rect -403 36495 -398 36509
rect -413 36485 -408 36495
rect -403 36471 -398 36485
rect -402 36470 -398 36471
rect -378 36470 -374 36540
rect -354 36470 -350 36540
rect -330 36470 -326 36540
rect -306 36470 -302 36540
rect -282 36470 -278 36540
rect -258 36470 -254 36540
rect -234 36470 -230 36540
rect -210 36470 -206 36540
rect -186 36470 -182 36540
rect -162 36470 -158 36540
rect -138 36470 -134 36540
rect -114 36470 -110 36540
rect -90 36470 -86 36540
rect -66 36470 -62 36540
rect -42 36470 -38 36540
rect -18 36470 -14 36540
rect 6 36470 10 36540
rect 30 36470 34 36540
rect 54 36470 58 36540
rect 78 36470 82 36540
rect 102 36470 106 36540
rect 126 36470 130 36540
rect 150 36470 154 36540
rect 174 36470 178 36540
rect 198 36470 202 36540
rect 222 36470 226 36540
rect 246 36470 250 36540
rect 270 36470 274 36540
rect 294 36471 298 36540
rect 283 36470 317 36471
rect -2393 36468 317 36470
rect -2371 36446 -2366 36468
rect -2348 36446 -2343 36468
rect -2325 36446 -2320 36468
rect -2060 36462 -2050 36468
rect -2309 36446 -2301 36456
rect -2060 36455 -2030 36462
rect -2000 36458 -1992 36468
rect -1972 36466 -1942 36468
rect -1958 36465 -1942 36466
rect -1844 36464 -1806 36468
rect -2068 36448 -2062 36455
rect -2062 36446 -2036 36448
rect -2393 36444 -2036 36446
rect -2030 36446 -2012 36448
rect -2004 36446 -1990 36458
rect -1844 36457 -1798 36462
rect -1806 36455 -1798 36457
rect -1854 36453 -1844 36455
rect -1854 36448 -1806 36453
rect -1864 36446 -1796 36447
rect -1655 36446 -1647 36456
rect -1642 36446 -1637 36468
rect -1619 36446 -1614 36468
rect -1530 36446 -1526 36468
rect -1506 36446 -1502 36468
rect -1482 36446 -1478 36468
rect -1458 36446 -1454 36468
rect -1434 36446 -1430 36468
rect -1410 36446 -1406 36468
rect -1386 36446 -1382 36468
rect -1362 36446 -1358 36468
rect -1338 36446 -1334 36468
rect -1314 36446 -1310 36468
rect -1290 36446 -1286 36468
rect -1266 36446 -1262 36468
rect -1242 36446 -1238 36468
rect -1218 36446 -1214 36468
rect -1194 36446 -1190 36468
rect -1170 36446 -1166 36468
rect -1146 36446 -1142 36468
rect -1122 36446 -1118 36468
rect -1098 36446 -1094 36468
rect -1074 36446 -1070 36468
rect -1050 36446 -1046 36468
rect -1026 36446 -1022 36468
rect -1002 36446 -998 36468
rect -978 36446 -974 36468
rect -954 36446 -950 36468
rect -930 36446 -926 36468
rect -906 36446 -902 36468
rect -882 36446 -878 36468
rect -858 36446 -854 36468
rect -834 36446 -830 36468
rect -810 36446 -806 36468
rect -786 36446 -782 36468
rect -762 36446 -758 36468
rect -738 36446 -734 36468
rect -714 36446 -710 36468
rect -690 36446 -686 36468
rect -666 36446 -662 36468
rect -642 36446 -638 36468
rect -618 36446 -614 36468
rect -594 36447 -590 36468
rect -605 36446 -571 36447
rect -2030 36444 -571 36446
rect -2371 36398 -2366 36444
rect -2348 36398 -2343 36444
rect -2325 36398 -2320 36444
rect -2317 36440 -2309 36444
rect -2060 36440 -2050 36444
rect -2060 36438 -2036 36440
rect -2060 36436 -2030 36438
rect -2292 36430 -2030 36436
rect -2092 36414 -2062 36416
rect -2094 36410 -2062 36414
rect -2000 36398 -1992 36444
rect -1844 36437 -1806 36444
rect -1663 36440 -1655 36444
rect -1844 36430 -1680 36436
rect -1854 36414 -1806 36416
rect -1854 36410 -1680 36414
rect -1642 36398 -1637 36444
rect -1619 36398 -1614 36444
rect -1530 36398 -1526 36444
rect -1506 36398 -1502 36444
rect -1482 36398 -1478 36444
rect -1458 36398 -1454 36444
rect -1434 36398 -1430 36444
rect -1410 36398 -1406 36444
rect -1386 36398 -1382 36444
rect -1362 36398 -1358 36444
rect -1338 36398 -1334 36444
rect -1314 36398 -1310 36444
rect -1290 36398 -1286 36444
rect -1266 36398 -1262 36444
rect -1242 36398 -1238 36444
rect -1218 36398 -1214 36444
rect -1194 36398 -1190 36444
rect -1170 36398 -1166 36444
rect -1146 36398 -1142 36444
rect -1122 36398 -1118 36444
rect -1098 36398 -1094 36444
rect -1074 36398 -1070 36444
rect -1050 36398 -1046 36444
rect -1026 36398 -1022 36444
rect -1002 36398 -998 36444
rect -978 36398 -974 36444
rect -954 36398 -950 36444
rect -930 36398 -926 36444
rect -906 36398 -902 36444
rect -882 36398 -878 36444
rect -858 36398 -854 36444
rect -834 36398 -830 36444
rect -810 36398 -806 36444
rect -786 36398 -782 36444
rect -762 36398 -758 36444
rect -738 36398 -734 36444
rect -714 36398 -710 36444
rect -690 36398 -686 36444
rect -666 36398 -662 36444
rect -642 36398 -638 36444
rect -618 36398 -614 36444
rect -605 36437 -600 36444
rect -594 36437 -590 36444
rect -595 36423 -590 36437
rect -605 36413 -600 36423
rect -594 36413 -590 36423
rect -595 36399 -590 36413
rect -605 36398 -571 36399
rect -2393 36396 -571 36398
rect -2371 36374 -2366 36396
rect -2348 36374 -2343 36396
rect -2325 36374 -2320 36396
rect -2072 36394 -2036 36395
rect -2072 36388 -2054 36394
rect -2309 36380 -2301 36388
rect -2317 36374 -2309 36380
rect -2092 36379 -2062 36384
rect -2000 36375 -1992 36396
rect -1938 36395 -1906 36396
rect -1920 36394 -1906 36395
rect -1806 36388 -1680 36394
rect -1854 36379 -1806 36384
rect -1655 36380 -1647 36388
rect -1982 36375 -1966 36376
rect -2000 36374 -1966 36375
rect -1846 36374 -1806 36377
rect -1663 36374 -1655 36380
rect -1642 36374 -1637 36396
rect -1619 36374 -1614 36396
rect -1530 36374 -1526 36396
rect -1506 36374 -1502 36396
rect -1482 36374 -1478 36396
rect -1458 36374 -1454 36396
rect -1434 36374 -1430 36396
rect -1410 36374 -1406 36396
rect -1386 36374 -1382 36396
rect -1362 36374 -1358 36396
rect -1338 36374 -1334 36396
rect -1314 36374 -1310 36396
rect -1290 36374 -1286 36396
rect -1266 36374 -1262 36396
rect -1242 36374 -1238 36396
rect -1218 36374 -1214 36396
rect -1194 36374 -1190 36396
rect -1170 36374 -1166 36396
rect -1146 36374 -1142 36396
rect -1122 36374 -1118 36396
rect -1098 36374 -1094 36396
rect -1074 36374 -1070 36396
rect -1050 36374 -1046 36396
rect -1026 36374 -1022 36396
rect -1002 36374 -998 36396
rect -978 36374 -974 36396
rect -954 36374 -950 36396
rect -930 36374 -926 36396
rect -906 36374 -902 36396
rect -882 36374 -878 36396
rect -858 36374 -854 36396
rect -834 36374 -830 36396
rect -810 36374 -806 36396
rect -786 36374 -782 36396
rect -762 36374 -758 36396
rect -738 36374 -734 36396
rect -714 36374 -710 36396
rect -690 36374 -686 36396
rect -666 36374 -662 36396
rect -642 36374 -638 36396
rect -618 36374 -614 36396
rect -605 36389 -600 36396
rect -595 36375 -590 36389
rect -594 36374 -590 36375
rect -570 36374 -566 36468
rect -546 36374 -542 36468
rect -522 36374 -518 36468
rect -498 36374 -494 36468
rect -474 36374 -470 36468
rect -450 36374 -446 36468
rect -426 36374 -422 36468
rect -402 36374 -398 36468
rect -378 36443 -374 36468
rect -378 36422 -371 36443
rect -354 36422 -350 36468
rect -330 36422 -326 36468
rect -306 36422 -302 36468
rect -282 36422 -278 36468
rect -258 36422 -254 36468
rect -234 36422 -230 36468
rect -210 36422 -206 36468
rect -186 36422 -182 36468
rect -162 36422 -158 36468
rect -138 36422 -134 36468
rect -114 36422 -110 36468
rect -90 36422 -86 36468
rect -66 36422 -62 36468
rect -42 36422 -38 36468
rect -18 36422 -14 36468
rect 6 36422 10 36468
rect 30 36422 34 36468
rect 54 36422 58 36468
rect 78 36422 82 36468
rect 102 36422 106 36468
rect 126 36422 130 36468
rect 150 36422 154 36468
rect 174 36422 178 36468
rect 198 36422 202 36468
rect 222 36422 226 36468
rect 246 36422 250 36468
rect 270 36422 274 36468
rect 283 36461 288 36468
rect 294 36461 298 36468
rect 293 36447 298 36461
rect 294 36422 298 36447
rect 318 36422 322 36540
rect 342 36422 346 36540
rect 366 36422 370 36540
rect 390 36422 394 36540
rect 414 36491 418 36540
rect 427 36533 432 36540
rect 438 36533 442 36540
rect 437 36519 442 36533
rect 414 36467 421 36491
rect 414 36422 418 36467
rect 438 36422 442 36519
rect 462 36467 466 36636
rect 462 36443 469 36467
rect 462 36422 466 36443
rect 486 36422 490 36636
rect 510 36422 514 36636
rect 534 36422 538 36636
rect 558 36422 562 36636
rect 582 36422 586 36636
rect 606 36422 610 36636
rect 630 36422 634 36636
rect 654 36422 658 36636
rect 678 36422 682 36636
rect 702 36422 706 36636
rect 726 36422 730 36636
rect 750 36422 754 36636
rect 774 36422 778 36636
rect 798 36422 802 36636
rect 822 36422 826 36636
rect 846 36422 850 36636
rect 870 36422 874 36636
rect 894 36422 898 36636
rect 918 36422 922 36636
rect 942 36422 946 36636
rect 966 36422 970 36636
rect 990 36422 994 36636
rect 1014 36422 1018 36636
rect 1038 36422 1042 36636
rect 1062 36422 1066 36636
rect 1086 36422 1090 36636
rect 1110 36422 1114 36636
rect 1134 36422 1138 36636
rect 1158 36422 1162 36636
rect 1182 36422 1186 36636
rect 1206 36422 1210 36636
rect 1213 36635 1227 36636
rect 1219 36629 1224 36635
rect 1229 36615 1234 36629
rect 1230 36422 1234 36615
rect 1243 36509 1248 36519
rect 1253 36495 1258 36509
rect 1254 36422 1258 36495
rect 1267 36422 1275 36423
rect -395 36420 1275 36422
rect -395 36419 -381 36420
rect -378 36395 -371 36420
rect -378 36374 -374 36395
rect -354 36374 -350 36420
rect -330 36374 -326 36420
rect -306 36374 -302 36420
rect -282 36374 -278 36420
rect -258 36374 -254 36420
rect -234 36374 -230 36420
rect -210 36374 -206 36420
rect -186 36374 -182 36420
rect -162 36374 -158 36420
rect -138 36374 -134 36420
rect -114 36374 -110 36420
rect -90 36374 -86 36420
rect -66 36374 -62 36420
rect -42 36374 -38 36420
rect -18 36374 -14 36420
rect 6 36374 10 36420
rect 30 36374 34 36420
rect 54 36374 58 36420
rect 78 36374 82 36420
rect 102 36374 106 36420
rect 126 36374 130 36420
rect 150 36374 154 36420
rect 174 36374 178 36420
rect 198 36374 202 36420
rect 222 36374 226 36420
rect 246 36374 250 36420
rect 270 36374 274 36420
rect 294 36374 298 36420
rect 318 36395 322 36420
rect 307 36374 315 36375
rect -2393 36372 315 36374
rect -2371 36350 -2366 36372
rect -2348 36350 -2343 36372
rect -2325 36350 -2320 36372
rect -2000 36370 -1966 36372
rect -2309 36352 -2301 36360
rect -2062 36359 -2054 36366
rect -2092 36352 -2084 36359
rect -2062 36352 -2026 36354
rect -2317 36350 -2309 36352
rect -2062 36350 -2012 36352
rect -2000 36350 -1992 36370
rect -1982 36369 -1966 36370
rect -1846 36368 -1806 36372
rect -1846 36361 -1798 36366
rect -1806 36359 -1798 36361
rect -1854 36357 -1846 36359
rect -1854 36352 -1806 36357
rect -1655 36352 -1647 36360
rect -1864 36350 -1796 36351
rect -1663 36350 -1655 36352
rect -1642 36350 -1637 36372
rect -1619 36350 -1614 36372
rect -1530 36350 -1526 36372
rect -1506 36350 -1502 36372
rect -1482 36350 -1478 36372
rect -1458 36350 -1454 36372
rect -1434 36350 -1430 36372
rect -1410 36350 -1406 36372
rect -1386 36350 -1382 36372
rect -1362 36350 -1358 36372
rect -1338 36350 -1334 36372
rect -1314 36350 -1310 36372
rect -1290 36350 -1286 36372
rect -1266 36350 -1262 36372
rect -1242 36350 -1238 36372
rect -1218 36350 -1214 36372
rect -1194 36350 -1190 36372
rect -1170 36350 -1166 36372
rect -1146 36350 -1142 36372
rect -1122 36350 -1118 36372
rect -1098 36350 -1094 36372
rect -1074 36350 -1070 36372
rect -1050 36350 -1046 36372
rect -1026 36350 -1022 36372
rect -1002 36350 -998 36372
rect -978 36350 -974 36372
rect -954 36350 -950 36372
rect -930 36350 -926 36372
rect -906 36350 -902 36372
rect -882 36350 -878 36372
rect -858 36350 -854 36372
rect -834 36350 -830 36372
rect -810 36350 -806 36372
rect -786 36350 -782 36372
rect -762 36350 -758 36372
rect -738 36350 -734 36372
rect -714 36350 -710 36372
rect -690 36350 -686 36372
rect -666 36350 -662 36372
rect -642 36350 -638 36372
rect -618 36350 -614 36372
rect -594 36350 -590 36372
rect -570 36371 -566 36372
rect -2393 36348 -573 36350
rect -2371 36302 -2366 36348
rect -2348 36302 -2343 36348
rect -2325 36302 -2320 36348
rect -2317 36344 -2309 36348
rect -2062 36344 -2054 36348
rect -2154 36340 -2138 36342
rect -2057 36340 -2054 36344
rect -2292 36334 -2054 36340
rect -2052 36334 -2044 36344
rect -2092 36318 -2062 36320
rect -2094 36314 -2062 36318
rect -2000 36302 -1992 36348
rect -1846 36341 -1806 36348
rect -1663 36344 -1655 36348
rect -1846 36334 -1680 36340
rect -1854 36318 -1806 36320
rect -1854 36314 -1680 36318
rect -1979 36302 -1945 36304
rect -1642 36302 -1637 36348
rect -1619 36302 -1614 36348
rect -1530 36302 -1526 36348
rect -1506 36302 -1502 36348
rect -1482 36302 -1478 36348
rect -1458 36302 -1454 36348
rect -1434 36302 -1430 36348
rect -1410 36302 -1406 36348
rect -1386 36302 -1382 36348
rect -1362 36302 -1358 36348
rect -1338 36302 -1334 36348
rect -1314 36302 -1310 36348
rect -1290 36302 -1286 36348
rect -1266 36302 -1262 36348
rect -1242 36302 -1238 36348
rect -1218 36302 -1214 36348
rect -1194 36302 -1190 36348
rect -1170 36302 -1166 36348
rect -1146 36302 -1142 36348
rect -1122 36302 -1118 36348
rect -1098 36302 -1094 36348
rect -1074 36302 -1070 36348
rect -1050 36302 -1046 36348
rect -1026 36302 -1022 36348
rect -1002 36302 -998 36348
rect -978 36302 -974 36348
rect -954 36302 -950 36348
rect -930 36302 -926 36348
rect -906 36302 -902 36348
rect -882 36302 -878 36348
rect -858 36302 -854 36348
rect -834 36302 -830 36348
rect -810 36302 -806 36348
rect -786 36302 -782 36348
rect -762 36302 -758 36348
rect -738 36302 -734 36348
rect -714 36302 -710 36348
rect -690 36302 -686 36348
rect -666 36302 -662 36348
rect -642 36302 -638 36348
rect -618 36302 -614 36348
rect -594 36302 -590 36348
rect -587 36347 -573 36348
rect -2393 36300 -573 36302
rect -2371 36254 -2366 36300
rect -2348 36254 -2343 36300
rect -2325 36254 -2320 36300
rect -2080 36299 -1906 36300
rect -2080 36298 -2036 36299
rect -2080 36292 -2054 36298
rect -2309 36284 -2301 36290
rect -2317 36274 -2309 36284
rect -2070 36283 -2040 36290
rect -2054 36275 -2040 36278
rect -2000 36273 -1992 36299
rect -1920 36298 -1906 36299
rect -1850 36292 -1846 36300
rect -1840 36292 -1792 36300
rect -1969 36280 -1966 36289
rect -1850 36285 -1802 36290
rect -1906 36283 -1802 36285
rect -1655 36284 -1647 36290
rect -1906 36282 -1850 36283
rect -1846 36275 -1802 36281
rect -1663 36274 -1655 36284
rect -1860 36273 -1798 36274
rect -2078 36266 -2070 36273
rect -2309 36256 -2301 36262
rect -2317 36254 -2309 36256
rect -2154 36254 -2145 36264
rect -2044 36263 -2040 36268
rect -2028 36266 -1945 36273
rect -1929 36266 -1794 36273
rect -2070 36256 -2040 36263
rect -2044 36254 -2028 36256
rect -2000 36254 -1992 36266
rect -1860 36265 -1798 36266
rect -1850 36256 -1802 36263
rect -1655 36256 -1647 36262
rect -1978 36254 -1942 36255
rect -1663 36254 -1655 36256
rect -1642 36254 -1637 36300
rect -1619 36254 -1614 36300
rect -1530 36254 -1526 36300
rect -1506 36254 -1502 36300
rect -1482 36254 -1478 36300
rect -1458 36254 -1454 36300
rect -1434 36254 -1430 36300
rect -1410 36254 -1406 36300
rect -1386 36254 -1382 36300
rect -1362 36254 -1358 36300
rect -1338 36254 -1334 36300
rect -1314 36254 -1310 36300
rect -1290 36254 -1286 36300
rect -1266 36254 -1262 36300
rect -1242 36254 -1238 36300
rect -1218 36254 -1214 36300
rect -1194 36254 -1190 36300
rect -1170 36254 -1166 36300
rect -1146 36254 -1142 36300
rect -1122 36254 -1118 36300
rect -1098 36254 -1094 36300
rect -1074 36254 -1070 36300
rect -1050 36254 -1046 36300
rect -1026 36254 -1022 36300
rect -1002 36254 -998 36300
rect -978 36254 -974 36300
rect -954 36254 -950 36300
rect -930 36254 -926 36300
rect -906 36254 -902 36300
rect -882 36254 -878 36300
rect -858 36254 -854 36300
rect -834 36254 -830 36300
rect -810 36254 -806 36300
rect -786 36254 -782 36300
rect -762 36254 -758 36300
rect -738 36254 -734 36300
rect -714 36254 -710 36300
rect -690 36254 -686 36300
rect -666 36254 -662 36300
rect -642 36254 -638 36300
rect -618 36254 -614 36300
rect -594 36254 -590 36300
rect -587 36299 -573 36300
rect -570 36299 -563 36371
rect -570 36254 -566 36299
rect -546 36254 -542 36372
rect -522 36254 -518 36372
rect -498 36254 -494 36372
rect -474 36254 -470 36372
rect -450 36254 -446 36372
rect -426 36254 -422 36372
rect -402 36254 -398 36372
rect -378 36254 -374 36372
rect -354 36254 -350 36372
rect -330 36254 -326 36372
rect -306 36254 -302 36372
rect -282 36254 -278 36372
rect -258 36254 -254 36372
rect -234 36254 -230 36372
rect -210 36254 -206 36372
rect -186 36254 -182 36372
rect -162 36254 -158 36372
rect -138 36254 -134 36372
rect -114 36254 -110 36372
rect -90 36254 -86 36372
rect -66 36254 -62 36372
rect -42 36254 -38 36372
rect -18 36254 -14 36372
rect 6 36254 10 36372
rect 30 36254 34 36372
rect 54 36254 58 36372
rect 78 36254 82 36372
rect 102 36254 106 36372
rect 126 36254 130 36372
rect 150 36254 154 36372
rect 174 36254 178 36372
rect 198 36254 202 36372
rect 222 36254 226 36372
rect 246 36254 250 36372
rect 270 36254 274 36372
rect 294 36254 298 36372
rect 301 36371 315 36372
rect 318 36371 325 36395
rect 307 36365 312 36371
rect 318 36365 322 36371
rect 317 36351 322 36365
rect 318 36254 322 36351
rect 342 36299 346 36420
rect 342 36275 349 36299
rect 342 36254 346 36275
rect 366 36254 370 36420
rect 390 36254 394 36420
rect 414 36254 418 36420
rect 438 36255 442 36420
rect 427 36254 461 36255
rect -2393 36252 461 36254
rect -2371 36158 -2366 36252
rect -2348 36158 -2343 36252
rect -2325 36214 -2320 36252
rect -2317 36246 -2309 36252
rect -2145 36248 -2138 36252
rect -2070 36248 -2054 36252
rect -2078 36239 -2054 36246
rect -2062 36214 -2032 36215
rect -2000 36214 -1992 36252
rect -1846 36248 -1802 36252
rect -1846 36238 -1792 36247
rect -1663 36246 -1655 36252
rect -1942 36216 -1937 36228
rect -1850 36225 -1822 36226
rect -1850 36221 -1802 36225
rect -2325 36206 -2317 36214
rect -2062 36212 -1961 36214
rect -2325 36186 -2320 36206
rect -2317 36198 -2309 36206
rect -2062 36199 -2040 36210
rect -2032 36205 -1961 36212
rect -1947 36206 -1942 36214
rect -1842 36212 -1794 36215
rect -2070 36194 -2022 36198
rect -2325 36174 -2317 36186
rect -2325 36158 -2320 36174
rect -2317 36170 -2309 36174
rect -2309 36158 -2301 36170
rect -2068 36163 -2038 36170
rect -2000 36160 -1992 36205
rect -1942 36204 -1937 36206
rect -1932 36196 -1927 36204
rect -1912 36201 -1896 36207
rect -1842 36199 -1802 36210
rect -1671 36206 -1663 36214
rect -1663 36198 -1655 36206
rect -1850 36194 -1680 36198
rect -1937 36180 -1934 36182
rect -1926 36180 -1921 36185
rect -1926 36175 -1924 36180
rect -1916 36172 -1914 36175
rect -1842 36172 -1794 36181
rect -1671 36174 -1663 36186
rect -1924 36162 -1916 36171
rect -1663 36170 -1655 36174
rect -1852 36163 -1804 36170
rect -1916 36161 -1914 36162
rect -2025 36159 -1991 36160
rect -2025 36158 -1975 36159
rect -1842 36158 -1804 36161
rect -1655 36158 -1647 36170
rect -1642 36158 -1637 36252
rect -1619 36158 -1614 36252
rect -1530 36158 -1526 36252
rect -1506 36158 -1502 36252
rect -1482 36158 -1478 36252
rect -1458 36158 -1454 36252
rect -1434 36158 -1430 36252
rect -1410 36158 -1406 36252
rect -1386 36158 -1382 36252
rect -1362 36158 -1358 36252
rect -1338 36158 -1334 36252
rect -1314 36158 -1310 36252
rect -1290 36158 -1286 36252
rect -1266 36158 -1262 36252
rect -1242 36158 -1238 36252
rect -1218 36158 -1214 36252
rect -1194 36158 -1190 36252
rect -1170 36158 -1166 36252
rect -1146 36158 -1142 36252
rect -1122 36158 -1118 36252
rect -1098 36158 -1094 36252
rect -1074 36158 -1070 36252
rect -1050 36158 -1046 36252
rect -1026 36158 -1022 36252
rect -1002 36158 -998 36252
rect -978 36158 -974 36252
rect -954 36158 -950 36252
rect -930 36158 -926 36252
rect -906 36158 -902 36252
rect -882 36158 -878 36252
rect -858 36158 -854 36252
rect -834 36158 -830 36252
rect -810 36158 -806 36252
rect -786 36158 -782 36252
rect -762 36207 -758 36252
rect -773 36206 -739 36207
rect -738 36206 -734 36252
rect -714 36206 -710 36252
rect -690 36206 -686 36252
rect -666 36206 -662 36252
rect -642 36206 -638 36252
rect -618 36206 -614 36252
rect -594 36206 -590 36252
rect -570 36206 -566 36252
rect -546 36206 -542 36252
rect -522 36206 -518 36252
rect -498 36206 -494 36252
rect -474 36206 -470 36252
rect -450 36206 -446 36252
rect -426 36206 -422 36252
rect -402 36206 -398 36252
rect -378 36206 -374 36252
rect -354 36206 -350 36252
rect -330 36206 -326 36252
rect -306 36206 -302 36252
rect -282 36206 -278 36252
rect -258 36206 -254 36252
rect -234 36206 -230 36252
rect -210 36206 -206 36252
rect -186 36206 -182 36252
rect -162 36206 -158 36252
rect -138 36206 -134 36252
rect -114 36206 -110 36252
rect -90 36206 -86 36252
rect -66 36206 -62 36252
rect -42 36206 -38 36252
rect -18 36206 -14 36252
rect 6 36206 10 36252
rect 30 36206 34 36252
rect 54 36206 58 36252
rect 78 36206 82 36252
rect 102 36206 106 36252
rect 126 36206 130 36252
rect 150 36206 154 36252
rect 174 36206 178 36252
rect 198 36206 202 36252
rect 222 36206 226 36252
rect 246 36206 250 36252
rect 270 36206 274 36252
rect 294 36206 298 36252
rect 318 36206 322 36252
rect 342 36206 346 36252
rect 366 36206 370 36252
rect 390 36206 394 36252
rect 414 36206 418 36252
rect 427 36245 432 36252
rect 438 36245 442 36252
rect 437 36231 442 36245
rect 438 36206 442 36231
rect 462 36206 466 36420
rect 486 36206 490 36420
rect 510 36206 514 36420
rect 534 36206 538 36420
rect 558 36206 562 36420
rect 582 36206 586 36420
rect 606 36206 610 36420
rect 630 36206 634 36420
rect 654 36206 658 36420
rect 678 36206 682 36420
rect 702 36327 706 36420
rect 691 36326 725 36327
rect 726 36326 730 36420
rect 750 36326 754 36420
rect 774 36326 778 36420
rect 798 36326 802 36420
rect 822 36326 826 36420
rect 846 36326 850 36420
rect 870 36326 874 36420
rect 894 36326 898 36420
rect 918 36326 922 36420
rect 942 36326 946 36420
rect 966 36326 970 36420
rect 990 36326 994 36420
rect 1014 36326 1018 36420
rect 1038 36326 1042 36420
rect 1062 36326 1066 36420
rect 1086 36326 1090 36420
rect 1110 36326 1114 36420
rect 1134 36326 1138 36420
rect 1158 36326 1162 36420
rect 1182 36326 1186 36420
rect 1206 36326 1210 36420
rect 1230 36326 1234 36420
rect 1254 36326 1258 36420
rect 1261 36419 1275 36420
rect 1267 36413 1272 36419
rect 1277 36399 1282 36413
rect 1267 36341 1272 36351
rect 1278 36341 1282 36399
rect 1277 36327 1282 36341
rect 1291 36337 1299 36341
rect 1285 36327 1291 36337
rect 1267 36326 1299 36327
rect 691 36324 1299 36326
rect 691 36317 696 36324
rect 702 36317 706 36324
rect 701 36303 706 36317
rect 691 36293 696 36303
rect 701 36279 706 36293
rect 702 36206 706 36279
rect 726 36251 730 36324
rect 726 36230 733 36251
rect 750 36230 754 36324
rect 774 36230 778 36324
rect 798 36230 802 36324
rect 822 36230 826 36324
rect 846 36230 850 36324
rect 870 36230 874 36324
rect 894 36230 898 36324
rect 918 36230 922 36324
rect 942 36230 946 36324
rect 966 36230 970 36324
rect 990 36231 994 36324
rect 979 36230 1013 36231
rect 709 36228 1013 36230
rect 709 36227 723 36228
rect -773 36204 723 36206
rect -773 36197 -768 36204
rect -762 36197 -758 36204
rect -763 36183 -758 36197
rect -773 36173 -768 36183
rect -763 36159 -758 36173
rect -762 36158 -758 36159
rect -738 36158 -734 36204
rect -714 36158 -710 36204
rect -690 36158 -686 36204
rect -666 36158 -662 36204
rect -642 36158 -638 36204
rect -618 36158 -614 36204
rect -594 36158 -590 36204
rect -570 36158 -566 36204
rect -546 36158 -542 36204
rect -522 36158 -518 36204
rect -498 36158 -494 36204
rect -474 36158 -470 36204
rect -450 36158 -446 36204
rect -426 36158 -422 36204
rect -402 36158 -398 36204
rect -378 36158 -374 36204
rect -354 36158 -350 36204
rect -330 36158 -326 36204
rect -306 36158 -302 36204
rect -282 36158 -278 36204
rect -258 36158 -254 36204
rect -234 36158 -230 36204
rect -210 36158 -206 36204
rect -186 36158 -182 36204
rect -162 36158 -158 36204
rect -138 36158 -134 36204
rect -114 36158 -110 36204
rect -90 36158 -86 36204
rect -66 36158 -62 36204
rect -42 36158 -38 36204
rect -18 36158 -14 36204
rect 6 36158 10 36204
rect 30 36158 34 36204
rect 54 36158 58 36204
rect 78 36158 82 36204
rect 102 36158 106 36204
rect 126 36158 130 36204
rect 150 36158 154 36204
rect 174 36158 178 36204
rect 198 36158 202 36204
rect 222 36158 226 36204
rect 246 36158 250 36204
rect 270 36158 274 36204
rect 294 36158 298 36204
rect 318 36158 322 36204
rect 342 36158 346 36204
rect 366 36158 370 36204
rect 390 36158 394 36204
rect 414 36158 418 36204
rect 438 36158 442 36204
rect 462 36179 466 36204
rect -2393 36156 459 36158
rect -2371 36134 -2366 36156
rect -2348 36134 -2343 36156
rect -2325 36146 -2317 36156
rect -2076 36146 -2068 36153
rect -2062 36146 -2001 36153
rect -2325 36134 -2320 36146
rect -2317 36142 -2309 36146
rect -2015 36145 -2001 36146
rect -2309 36134 -2301 36142
rect -2068 36136 -2062 36143
rect -2000 36138 -1992 36156
rect -1974 36154 -1960 36156
rect -1842 36155 -1804 36156
rect -1862 36153 -1794 36154
rect -1985 36151 -1794 36153
rect -1985 36146 -1852 36151
rect -1842 36145 -1794 36151
rect -1671 36146 -1663 36156
rect -2015 36136 -1985 36138
rect -1852 36136 -1804 36143
rect -1663 36142 -1655 36146
rect -2000 36134 -1992 36136
rect -1976 36134 -1940 36135
rect -1655 36134 -1647 36142
rect -1642 36134 -1637 36156
rect -1619 36134 -1614 36156
rect -1530 36134 -1526 36156
rect -1506 36134 -1502 36156
rect -1482 36134 -1478 36156
rect -1458 36134 -1454 36156
rect -1434 36134 -1430 36156
rect -1410 36134 -1406 36156
rect -1386 36134 -1382 36156
rect -1362 36134 -1358 36156
rect -1338 36134 -1334 36156
rect -1314 36134 -1310 36156
rect -1290 36134 -1286 36156
rect -1266 36134 -1262 36156
rect -1242 36134 -1238 36156
rect -1218 36134 -1214 36156
rect -1194 36134 -1190 36156
rect -1170 36134 -1166 36156
rect -1146 36134 -1142 36156
rect -1122 36134 -1118 36156
rect -1098 36134 -1094 36156
rect -1074 36134 -1070 36156
rect -1050 36134 -1046 36156
rect -1026 36134 -1022 36156
rect -1002 36134 -998 36156
rect -978 36134 -974 36156
rect -954 36134 -950 36156
rect -930 36134 -926 36156
rect -906 36134 -902 36156
rect -882 36134 -878 36156
rect -858 36134 -854 36156
rect -834 36134 -830 36156
rect -810 36134 -806 36156
rect -786 36134 -782 36156
rect -762 36134 -758 36156
rect -738 36134 -734 36156
rect -714 36134 -710 36156
rect -690 36134 -686 36156
rect -666 36134 -662 36156
rect -642 36134 -638 36156
rect -618 36134 -614 36156
rect -594 36134 -590 36156
rect -570 36134 -566 36156
rect -546 36134 -542 36156
rect -522 36134 -518 36156
rect -498 36134 -494 36156
rect -474 36134 -470 36156
rect -450 36134 -446 36156
rect -426 36134 -422 36156
rect -402 36134 -398 36156
rect -378 36134 -374 36156
rect -354 36134 -350 36156
rect -330 36134 -326 36156
rect -306 36134 -302 36156
rect -282 36134 -278 36156
rect -258 36134 -254 36156
rect -234 36134 -230 36156
rect -210 36134 -206 36156
rect -186 36134 -182 36156
rect -162 36134 -158 36156
rect -138 36134 -134 36156
rect -114 36134 -110 36156
rect -90 36134 -86 36156
rect -66 36134 -62 36156
rect -42 36134 -38 36156
rect -18 36134 -14 36156
rect 6 36134 10 36156
rect 30 36134 34 36156
rect 54 36134 58 36156
rect 78 36134 82 36156
rect 102 36134 106 36156
rect 126 36134 130 36156
rect 150 36134 154 36156
rect 174 36134 178 36156
rect 198 36134 202 36156
rect 222 36134 226 36156
rect 246 36134 250 36156
rect 270 36134 274 36156
rect 294 36134 298 36156
rect 318 36134 322 36156
rect 342 36134 346 36156
rect 366 36134 370 36156
rect 390 36134 394 36156
rect 414 36134 418 36156
rect 438 36134 442 36156
rect 445 36155 459 36156
rect 462 36155 469 36179
rect 462 36134 466 36155
rect 486 36134 490 36204
rect 510 36134 514 36204
rect 534 36134 538 36204
rect 558 36134 562 36204
rect 582 36134 586 36204
rect 606 36134 610 36204
rect 630 36134 634 36204
rect 654 36134 658 36204
rect 678 36134 682 36204
rect 702 36134 706 36204
rect 709 36203 723 36204
rect 726 36203 733 36228
rect 726 36134 730 36203
rect 750 36134 754 36228
rect 774 36134 778 36228
rect 798 36134 802 36228
rect 822 36134 826 36228
rect 846 36134 850 36228
rect 870 36134 874 36228
rect 894 36134 898 36228
rect 918 36134 922 36228
rect 942 36134 946 36228
rect 966 36134 970 36228
rect 979 36221 984 36228
rect 990 36221 994 36228
rect 989 36207 994 36221
rect 990 36134 994 36207
rect 1014 36155 1018 36324
rect -2393 36132 1011 36134
rect -2371 36062 -2366 36132
rect -2348 36062 -2343 36132
rect -2325 36130 -2320 36132
rect -2309 36130 -2301 36132
rect -2325 36118 -2317 36130
rect -2062 36119 -2032 36126
rect -2325 36098 -2320 36118
rect -2317 36114 -2309 36118
rect -2325 36090 -2317 36098
rect -2060 36092 -2030 36095
rect -2325 36070 -2320 36090
rect -2317 36082 -2309 36090
rect -2060 36079 -2038 36090
rect -2033 36083 -2030 36092
rect -2028 36088 -2027 36092
rect -2068 36074 -2038 36077
rect -2325 36062 -2317 36070
rect -2000 36065 -1992 36132
rect -1888 36127 -1874 36132
rect -1842 36128 -1804 36132
rect -1655 36130 -1647 36132
rect -1902 36125 -1874 36127
rect -1842 36118 -1794 36127
rect -1671 36118 -1663 36130
rect -1663 36114 -1655 36118
rect -1912 36107 -1884 36109
rect -1852 36101 -1804 36105
rect -1844 36092 -1796 36095
rect -1671 36090 -1663 36098
rect -1844 36079 -1804 36090
rect -1663 36082 -1655 36090
rect -1852 36074 -1680 36078
rect -2119 36062 -2069 36064
rect -2007 36062 -1977 36065
rect -1926 36062 -1892 36065
rect -1671 36062 -1663 36070
rect -1642 36062 -1637 36132
rect -1619 36062 -1614 36132
rect -1530 36062 -1526 36132
rect -1506 36062 -1502 36132
rect -1482 36062 -1478 36132
rect -1458 36062 -1454 36132
rect -1434 36062 -1430 36132
rect -1410 36062 -1406 36132
rect -1386 36062 -1382 36132
rect -1362 36062 -1358 36132
rect -1338 36062 -1334 36132
rect -1314 36062 -1310 36132
rect -1290 36062 -1286 36132
rect -1266 36062 -1262 36132
rect -1242 36062 -1238 36132
rect -1218 36062 -1214 36132
rect -1194 36062 -1190 36132
rect -1170 36062 -1166 36132
rect -1146 36062 -1142 36132
rect -1122 36062 -1118 36132
rect -1098 36062 -1094 36132
rect -1074 36062 -1070 36132
rect -1050 36062 -1046 36132
rect -1026 36062 -1022 36132
rect -1002 36062 -998 36132
rect -978 36062 -974 36132
rect -954 36062 -950 36132
rect -930 36062 -926 36132
rect -906 36062 -902 36132
rect -882 36062 -878 36132
rect -858 36062 -854 36132
rect -834 36062 -830 36132
rect -810 36062 -806 36132
rect -786 36062 -782 36132
rect -762 36062 -758 36132
rect -738 36131 -734 36132
rect -738 36110 -731 36131
rect -714 36110 -710 36132
rect -690 36110 -686 36132
rect -666 36110 -662 36132
rect -642 36110 -638 36132
rect -618 36110 -614 36132
rect -594 36110 -590 36132
rect -570 36110 -566 36132
rect -546 36110 -542 36132
rect -522 36110 -518 36132
rect -498 36110 -494 36132
rect -474 36110 -470 36132
rect -450 36110 -446 36132
rect -426 36110 -422 36132
rect -402 36110 -398 36132
rect -378 36110 -374 36132
rect -354 36110 -350 36132
rect -330 36110 -326 36132
rect -306 36110 -302 36132
rect -282 36110 -278 36132
rect -258 36110 -254 36132
rect -234 36110 -230 36132
rect -210 36110 -206 36132
rect -186 36110 -182 36132
rect -162 36110 -158 36132
rect -138 36110 -134 36132
rect -114 36110 -110 36132
rect -90 36110 -86 36132
rect -66 36110 -62 36132
rect -42 36110 -38 36132
rect -18 36110 -14 36132
rect 6 36110 10 36132
rect 30 36110 34 36132
rect 54 36110 58 36132
rect 78 36110 82 36132
rect 102 36110 106 36132
rect 126 36110 130 36132
rect 150 36110 154 36132
rect 174 36110 178 36132
rect 198 36110 202 36132
rect 222 36110 226 36132
rect 246 36110 250 36132
rect 270 36110 274 36132
rect 294 36110 298 36132
rect 318 36110 322 36132
rect 342 36110 346 36132
rect 366 36110 370 36132
rect 390 36110 394 36132
rect 414 36110 418 36132
rect 438 36110 442 36132
rect 462 36110 466 36132
rect 486 36110 490 36132
rect 510 36110 514 36132
rect 534 36110 538 36132
rect 558 36110 562 36132
rect 582 36110 586 36132
rect 606 36110 610 36132
rect 630 36110 634 36132
rect 654 36110 658 36132
rect 678 36110 682 36132
rect 702 36110 706 36132
rect 726 36110 730 36132
rect 750 36110 754 36132
rect 774 36110 778 36132
rect 798 36110 802 36132
rect 822 36110 826 36132
rect 846 36110 850 36132
rect 870 36110 874 36132
rect 894 36110 898 36132
rect 918 36110 922 36132
rect 942 36110 946 36132
rect 966 36110 970 36132
rect 990 36110 994 36132
rect 997 36131 1011 36132
rect 1014 36131 1021 36155
rect 1014 36110 1018 36131
rect 1038 36110 1042 36324
rect 1062 36110 1066 36324
rect 1086 36110 1090 36324
rect 1110 36110 1114 36324
rect 1134 36110 1138 36324
rect 1158 36110 1162 36324
rect 1182 36110 1186 36324
rect 1206 36110 1210 36324
rect 1230 36110 1234 36324
rect 1254 36111 1258 36324
rect 1267 36317 1272 36324
rect 1285 36323 1299 36324
rect 1277 36303 1282 36317
rect 1267 36125 1272 36135
rect 1278 36125 1282 36303
rect 1291 36197 1296 36207
rect 1301 36183 1306 36197
rect 1291 36149 1296 36159
rect 1302 36149 1306 36183
rect 1301 36135 1306 36149
rect 1277 36111 1282 36125
rect 1243 36110 1277 36111
rect -755 36108 1277 36110
rect -755 36107 -741 36108
rect -738 36083 -731 36108
rect -738 36062 -734 36083
rect -714 36062 -710 36108
rect -690 36062 -686 36108
rect -666 36062 -662 36108
rect -642 36062 -638 36108
rect -618 36062 -614 36108
rect -594 36062 -590 36108
rect -570 36062 -566 36108
rect -546 36062 -542 36108
rect -522 36062 -518 36108
rect -498 36062 -494 36108
rect -474 36062 -470 36108
rect -450 36062 -446 36108
rect -426 36062 -422 36108
rect -402 36062 -398 36108
rect -378 36062 -374 36108
rect -354 36062 -350 36108
rect -330 36062 -326 36108
rect -306 36062 -302 36108
rect -282 36062 -278 36108
rect -258 36062 -254 36108
rect -234 36062 -230 36108
rect -210 36062 -206 36108
rect -186 36062 -182 36108
rect -162 36062 -158 36108
rect -138 36062 -134 36108
rect -114 36062 -110 36108
rect -90 36062 -86 36108
rect -66 36062 -62 36108
rect -42 36062 -38 36108
rect -18 36062 -14 36108
rect 6 36062 10 36108
rect 30 36062 34 36108
rect 54 36062 58 36108
rect 78 36062 82 36108
rect 102 36062 106 36108
rect 126 36062 130 36108
rect 150 36062 154 36108
rect 174 36062 178 36108
rect 198 36062 202 36108
rect 222 36062 226 36108
rect 246 36062 250 36108
rect 270 36062 274 36108
rect 294 36062 298 36108
rect 318 36062 322 36108
rect 342 36062 346 36108
rect 366 36062 370 36108
rect 390 36062 394 36108
rect 414 36062 418 36108
rect 438 36062 442 36108
rect 462 36062 466 36108
rect 486 36062 490 36108
rect 510 36062 514 36108
rect 534 36062 538 36108
rect 558 36062 562 36108
rect 582 36062 586 36108
rect 606 36062 610 36108
rect 630 36062 634 36108
rect 654 36062 658 36108
rect 678 36062 682 36108
rect 702 36062 706 36108
rect 726 36062 730 36108
rect 739 36077 744 36087
rect 750 36077 754 36108
rect 749 36063 754 36077
rect 739 36062 773 36063
rect -2393 36060 773 36062
rect -2371 36038 -2366 36060
rect -2348 36038 -2343 36060
rect -2325 36056 -2317 36060
rect -2325 36040 -2320 36056
rect -2317 36054 -2309 36056
rect -2309 36042 -2301 36054
rect -2000 36046 -1992 36060
rect -1671 36056 -1663 36060
rect -1663 36054 -1655 36056
rect -1844 36052 -1806 36054
rect -1854 36046 -1806 36050
rect -2068 36043 -2060 36046
rect -2030 36043 -1958 36046
rect -1942 36043 -1806 36046
rect -2317 36040 -2309 36042
rect -2000 36040 -1992 36043
rect -1655 36042 -1647 36054
rect -2325 36038 -2317 36040
rect -2033 36038 -1992 36040
rect -1844 36039 -1806 36041
rect -1663 36040 -1655 36042
rect -1864 36038 -1796 36039
rect -1671 36038 -1663 36040
rect -1642 36038 -1637 36060
rect -1619 36038 -1614 36060
rect -1530 36038 -1526 36060
rect -1506 36038 -1502 36060
rect -1482 36038 -1478 36060
rect -1458 36038 -1454 36060
rect -1434 36038 -1430 36060
rect -1410 36038 -1406 36060
rect -1386 36038 -1382 36060
rect -1362 36038 -1358 36060
rect -1338 36038 -1334 36060
rect -1314 36038 -1310 36060
rect -1290 36038 -1286 36060
rect -1266 36038 -1262 36060
rect -1242 36038 -1238 36060
rect -1218 36038 -1214 36060
rect -1194 36038 -1190 36060
rect -1170 36038 -1166 36060
rect -1146 36038 -1142 36060
rect -1122 36038 -1118 36060
rect -1098 36038 -1094 36060
rect -1074 36038 -1070 36060
rect -1050 36038 -1046 36060
rect -1026 36038 -1022 36060
rect -1002 36038 -998 36060
rect -978 36038 -974 36060
rect -954 36038 -950 36060
rect -930 36038 -926 36060
rect -906 36038 -902 36060
rect -882 36039 -878 36060
rect -893 36038 -859 36039
rect -2393 36036 -859 36038
rect -2371 36014 -2366 36036
rect -2348 36014 -2343 36036
rect -2325 36028 -2317 36036
rect -2060 36033 -2030 36036
rect -2000 36033 -1992 36036
rect -1972 36034 -1958 36036
rect -1904 36033 -1798 36036
rect -2078 36029 -2020 36033
rect -2023 36028 -2020 36029
rect -2000 36031 -1798 36033
rect -2000 36029 -1854 36031
rect -1844 36029 -1798 36031
rect -2325 36014 -2320 36028
rect -2317 36026 -2309 36028
rect -2020 36026 -2004 36028
rect -2000 36026 -1992 36029
rect -1671 36028 -1663 36036
rect -2309 36014 -2301 36026
rect -2020 36024 -1992 36026
rect -1844 36025 -1806 36027
rect -1663 36026 -1655 36028
rect -2023 36019 -1992 36024
rect -1854 36019 -1806 36023
rect -2068 36016 -2060 36019
rect -2030 36016 -1806 36019
rect -2074 36014 -2060 36016
rect -2020 36014 -2004 36016
rect -2000 36014 -1992 36016
rect -1655 36014 -1647 36026
rect -1642 36014 -1637 36036
rect -1619 36014 -1614 36036
rect -1530 36014 -1526 36036
rect -1506 36014 -1502 36036
rect -1482 36014 -1478 36036
rect -1458 36014 -1454 36036
rect -1434 36014 -1430 36036
rect -1410 36014 -1406 36036
rect -1386 36014 -1382 36036
rect -1362 36014 -1358 36036
rect -1338 36014 -1334 36036
rect -1314 36014 -1310 36036
rect -1290 36014 -1286 36036
rect -1266 36014 -1262 36036
rect -1242 36014 -1238 36036
rect -1218 36014 -1214 36036
rect -1194 36014 -1190 36036
rect -1170 36014 -1166 36036
rect -1146 36014 -1142 36036
rect -1122 36014 -1118 36036
rect -1098 36014 -1094 36036
rect -1074 36014 -1070 36036
rect -1050 36014 -1046 36036
rect -1026 36014 -1022 36036
rect -1002 36014 -998 36036
rect -978 36014 -974 36036
rect -954 36014 -950 36036
rect -930 36014 -926 36036
rect -906 36014 -902 36036
rect -893 36029 -888 36036
rect -882 36029 -878 36036
rect -883 36015 -878 36029
rect -882 36014 -878 36015
rect -858 36014 -854 36060
rect -834 36014 -830 36060
rect -810 36014 -806 36060
rect -786 36014 -782 36060
rect -762 36014 -758 36060
rect -738 36014 -734 36060
rect -714 36014 -710 36060
rect -690 36014 -686 36060
rect -666 36014 -662 36060
rect -642 36014 -638 36060
rect -618 36014 -614 36060
rect -594 36014 -590 36060
rect -570 36014 -566 36060
rect -546 36014 -542 36060
rect -522 36014 -518 36060
rect -498 36014 -494 36060
rect -474 36014 -470 36060
rect -450 36014 -446 36060
rect -426 36014 -422 36060
rect -402 36014 -398 36060
rect -378 36014 -374 36060
rect -354 36014 -350 36060
rect -330 36014 -326 36060
rect -306 36014 -302 36060
rect -282 36014 -278 36060
rect -258 36014 -254 36060
rect -234 36014 -230 36060
rect -210 36014 -206 36060
rect -186 36014 -182 36060
rect -162 36014 -158 36060
rect -138 36014 -134 36060
rect -114 36014 -110 36060
rect -90 36014 -86 36060
rect -66 36014 -62 36060
rect -42 36014 -38 36060
rect -18 36014 -14 36060
rect 6 36014 10 36060
rect 30 36014 34 36060
rect 54 36014 58 36060
rect 78 36014 82 36060
rect 102 36014 106 36060
rect 126 36014 130 36060
rect 150 36014 154 36060
rect 174 36014 178 36060
rect 198 36014 202 36060
rect 222 36014 226 36060
rect 246 36014 250 36060
rect 270 36014 274 36060
rect 294 36014 298 36060
rect 318 36014 322 36060
rect 342 36014 346 36060
rect 366 36014 370 36060
rect 390 36014 394 36060
rect 414 36014 418 36060
rect 438 36014 442 36060
rect 462 36014 466 36060
rect 486 36014 490 36060
rect 510 36014 514 36060
rect 534 36014 538 36060
rect 558 36014 562 36060
rect 582 36014 586 36060
rect 606 36014 610 36060
rect 630 36014 634 36060
rect 654 36014 658 36060
rect 678 36014 682 36060
rect 702 36014 706 36060
rect 726 36014 730 36060
rect 739 36053 744 36060
rect 749 36039 754 36053
rect 750 36014 754 36039
rect 774 36014 778 36108
rect 798 36014 802 36108
rect 822 36014 826 36108
rect 846 36014 850 36108
rect 870 36014 874 36108
rect 894 36014 898 36108
rect 918 36014 922 36108
rect 942 36014 946 36108
rect 966 36014 970 36108
rect 990 36014 994 36108
rect 1014 36014 1018 36108
rect 1038 36014 1042 36108
rect 1062 36015 1066 36108
rect 1051 36014 1085 36015
rect -2393 36012 -2060 36014
rect -2050 36012 1085 36014
rect -2371 35966 -2366 36012
rect -2348 35966 -2343 36012
rect -2325 36000 -2317 36012
rect -2109 36009 -2108 36012
rect -2117 36002 -2108 36009
rect -2325 35980 -2320 36000
rect -2317 35998 -2309 36000
rect -2109 35998 -2108 36002
rect -2060 36002 -2030 36009
rect -2060 35998 -2034 36002
rect -2325 35972 -2317 35980
rect -2101 35975 -2071 35978
rect -2325 35966 -2320 35972
rect -2317 35966 -2309 35972
rect -2000 35970 -1992 36012
rect -1844 36011 -1806 36012
rect -1844 36002 -1798 36009
rect -1671 36000 -1663 36012
rect -1844 35998 -1806 36000
rect -1663 35998 -1655 36000
rect -1854 35984 -1680 35988
rect -1846 35975 -1798 35978
rect -2079 35969 -2043 35970
rect -2007 35969 -1991 35970
rect -2079 35968 -2071 35969
rect -2079 35966 -2029 35968
rect -2011 35966 -1991 35969
rect -1846 35967 -1806 35973
rect -1671 35972 -1663 35980
rect -1864 35966 -1796 35967
rect -1663 35966 -1655 35972
rect -1642 35966 -1637 36012
rect -1619 35966 -1614 36012
rect -1530 35966 -1526 36012
rect -1506 35966 -1502 36012
rect -1482 35966 -1478 36012
rect -1458 35966 -1454 36012
rect -1434 35966 -1430 36012
rect -1410 35966 -1406 36012
rect -1386 35966 -1382 36012
rect -1362 35966 -1358 36012
rect -1338 35966 -1334 36012
rect -1314 35966 -1310 36012
rect -1290 35966 -1286 36012
rect -1266 35966 -1262 36012
rect -1242 35966 -1238 36012
rect -1218 35966 -1214 36012
rect -1194 35966 -1190 36012
rect -1170 35966 -1166 36012
rect -1146 35966 -1142 36012
rect -1122 35966 -1118 36012
rect -1098 35966 -1094 36012
rect -1074 35966 -1070 36012
rect -1050 35966 -1046 36012
rect -1026 35966 -1022 36012
rect -1002 35966 -998 36012
rect -978 35966 -974 36012
rect -954 35966 -950 36012
rect -930 35966 -926 36012
rect -906 35966 -902 36012
rect -882 35966 -878 36012
rect -858 35966 -854 36012
rect -834 35966 -830 36012
rect -810 35966 -806 36012
rect -786 35966 -782 36012
rect -762 35966 -758 36012
rect -738 35966 -734 36012
rect -714 35966 -710 36012
rect -690 35966 -686 36012
rect -666 35966 -662 36012
rect -642 35966 -638 36012
rect -618 35966 -614 36012
rect -594 35966 -590 36012
rect -570 35966 -566 36012
rect -546 35966 -542 36012
rect -522 35966 -518 36012
rect -498 35966 -494 36012
rect -474 35966 -470 36012
rect -450 35966 -446 36012
rect -426 35966 -422 36012
rect -402 35966 -398 36012
rect -378 35966 -374 36012
rect -354 35966 -350 36012
rect -330 35966 -326 36012
rect -306 35966 -302 36012
rect -282 35966 -278 36012
rect -258 35966 -254 36012
rect -234 35966 -230 36012
rect -210 35966 -206 36012
rect -186 35966 -182 36012
rect -162 35966 -158 36012
rect -138 35966 -134 36012
rect -114 35966 -110 36012
rect -90 35966 -86 36012
rect -66 35966 -62 36012
rect -53 35981 -48 35991
rect -42 35981 -38 36012
rect -43 35967 -38 35981
rect -42 35966 -38 35967
rect -18 35966 -14 36012
rect 6 35966 10 36012
rect 30 35966 34 36012
rect 54 35966 58 36012
rect 78 35966 82 36012
rect 102 35966 106 36012
rect 126 35966 130 36012
rect 150 35966 154 36012
rect 174 35966 178 36012
rect 198 35966 202 36012
rect 222 35966 226 36012
rect 246 35966 250 36012
rect 270 35966 274 36012
rect 294 35966 298 36012
rect 318 35966 322 36012
rect 342 35966 346 36012
rect 366 35966 370 36012
rect 390 35966 394 36012
rect 414 35966 418 36012
rect 438 35966 442 36012
rect 462 35966 466 36012
rect 486 35966 490 36012
rect 510 35966 514 36012
rect 534 35966 538 36012
rect 558 35966 562 36012
rect 582 35966 586 36012
rect 606 35966 610 36012
rect 630 35966 634 36012
rect 654 35966 658 36012
rect 678 35966 682 36012
rect 702 35966 706 36012
rect 726 35966 730 36012
rect 750 35966 754 36012
rect 774 36011 778 36012
rect -2393 35964 771 35966
rect -2371 35918 -2366 35964
rect -2348 35918 -2343 35964
rect -2325 35952 -2320 35964
rect -2079 35962 -2071 35964
rect -2072 35960 -2071 35962
rect -2109 35955 -2101 35960
rect -2101 35953 -2079 35955
rect -2069 35953 -2068 35960
rect -2325 35944 -2317 35952
rect -2079 35948 -2071 35953
rect -2325 35918 -2320 35944
rect -2317 35936 -2309 35944
rect -2074 35939 -2071 35948
rect -2069 35944 -2068 35948
rect -2109 35930 -2079 35933
rect -2082 35918 -2071 35919
rect -2000 35918 -1992 35964
rect -1846 35962 -1806 35964
rect -1854 35957 -1806 35961
rect -1854 35955 -1846 35957
rect -1846 35953 -1806 35955
rect -1806 35951 -1798 35953
rect -1846 35948 -1798 35951
rect -1846 35935 -1806 35946
rect -1671 35944 -1663 35952
rect -1663 35936 -1655 35944
rect -1854 35930 -1680 35934
rect -1979 35918 -1945 35920
rect -1642 35918 -1637 35964
rect -1619 35918 -1614 35964
rect -1530 35918 -1526 35964
rect -1506 35918 -1502 35964
rect -1482 35918 -1478 35964
rect -1458 35918 -1454 35964
rect -1434 35918 -1430 35964
rect -1410 35918 -1406 35964
rect -1386 35943 -1382 35964
rect -1397 35942 -1363 35943
rect -1362 35942 -1358 35964
rect -1338 35942 -1334 35964
rect -1314 35942 -1310 35964
rect -1290 35942 -1286 35964
rect -1266 35942 -1262 35964
rect -1242 35942 -1238 35964
rect -1218 35942 -1214 35964
rect -1194 35942 -1190 35964
rect -1170 35942 -1166 35964
rect -1146 35942 -1142 35964
rect -1122 35942 -1118 35964
rect -1098 35942 -1094 35964
rect -1074 35942 -1070 35964
rect -1050 35942 -1046 35964
rect -1026 35942 -1022 35964
rect -1002 35942 -998 35964
rect -978 35942 -974 35964
rect -954 35942 -950 35964
rect -930 35942 -926 35964
rect -906 35942 -902 35964
rect -882 35942 -878 35964
rect -858 35963 -854 35964
rect -1397 35940 -861 35942
rect -1397 35933 -1392 35940
rect -1386 35933 -1382 35940
rect -1387 35919 -1382 35933
rect -1397 35918 -1363 35919
rect -2393 35916 -1363 35918
rect -2371 35870 -2366 35916
rect -2348 35870 -2343 35916
rect -2325 35870 -2320 35916
rect -2082 35907 -2071 35916
rect -2070 35906 -2059 35907
rect -2309 35896 -2301 35906
rect -2070 35899 -2040 35906
rect -2317 35890 -2309 35896
rect -2070 35894 -2059 35899
rect -2070 35891 -2040 35894
rect -2070 35889 -2059 35891
rect -2000 35889 -1992 35916
rect -1850 35908 -1846 35916
rect -1840 35908 -1792 35916
rect -1896 35906 -1850 35907
rect -1896 35899 -1802 35906
rect -1896 35898 -1850 35899
rect -1846 35891 -1802 35897
rect -1655 35896 -1647 35906
rect -1663 35890 -1655 35896
rect -1860 35889 -1798 35890
rect -2078 35882 -2070 35889
rect -2061 35882 -2045 35884
rect -2040 35882 -1945 35889
rect -1929 35887 -1794 35889
rect -1929 35882 -1850 35887
rect -1846 35882 -1794 35887
rect -2070 35880 -2045 35882
rect -2309 35870 -2301 35878
rect -2147 35870 -2145 35880
rect -2070 35870 -2040 35880
rect -2000 35870 -1992 35882
rect -1846 35881 -1798 35882
rect -1850 35872 -1802 35879
rect -1978 35870 -1942 35871
rect -1655 35870 -1647 35878
rect -1642 35870 -1637 35916
rect -1619 35870 -1614 35916
rect -1530 35870 -1526 35916
rect -1506 35870 -1502 35916
rect -1482 35870 -1478 35916
rect -1458 35870 -1454 35916
rect -1434 35870 -1430 35916
rect -1410 35870 -1406 35916
rect -1397 35909 -1392 35916
rect -1387 35895 -1382 35909
rect -1386 35870 -1382 35895
rect -1362 35870 -1358 35940
rect -1338 35870 -1334 35940
rect -1314 35870 -1310 35940
rect -1290 35870 -1286 35940
rect -1266 35870 -1262 35940
rect -1242 35870 -1238 35940
rect -1218 35870 -1214 35940
rect -1194 35870 -1190 35940
rect -1170 35870 -1166 35940
rect -1146 35870 -1142 35940
rect -1122 35870 -1118 35940
rect -1098 35870 -1094 35940
rect -1074 35870 -1070 35940
rect -1050 35870 -1046 35940
rect -1026 35870 -1022 35940
rect -1002 35870 -998 35940
rect -978 35870 -974 35940
rect -954 35870 -950 35940
rect -930 35870 -926 35940
rect -906 35871 -902 35940
rect -917 35870 -883 35871
rect -2393 35868 -883 35870
rect -2371 35774 -2366 35868
rect -2348 35774 -2343 35868
rect -2325 35830 -2320 35868
rect -2317 35862 -2309 35868
rect -2145 35864 -2131 35868
rect -2072 35862 -2071 35864
rect -2070 35862 -2059 35868
rect -2078 35855 -2071 35862
rect -2070 35854 -2059 35855
rect -2062 35830 -2032 35831
rect -2000 35830 -1992 35868
rect -1846 35864 -1802 35868
rect -1846 35854 -1792 35863
rect -1663 35862 -1655 35868
rect -1942 35832 -1937 35844
rect -1850 35841 -1822 35842
rect -1850 35837 -1802 35841
rect -2325 35822 -2317 35830
rect -2062 35828 -1961 35830
rect -2325 35802 -2320 35822
rect -2317 35814 -2309 35822
rect -2062 35815 -2040 35826
rect -2032 35821 -1961 35828
rect -1947 35822 -1942 35830
rect -1842 35828 -1794 35831
rect -2070 35810 -2022 35814
rect -2325 35788 -2317 35802
rect -2072 35794 -2032 35795
rect -2102 35788 -2032 35794
rect -2325 35774 -2320 35788
rect -2317 35786 -2309 35788
rect -2309 35774 -2301 35786
rect -2070 35779 -2062 35784
rect -2000 35774 -1992 35821
rect -1942 35820 -1937 35822
rect -1932 35812 -1927 35820
rect -1912 35817 -1896 35823
rect -1842 35815 -1802 35826
rect -1671 35822 -1663 35830
rect -1663 35814 -1655 35822
rect -1850 35810 -1680 35814
rect -1924 35796 -1921 35798
rect -1806 35788 -1680 35794
rect -1671 35788 -1663 35802
rect -1663 35786 -1655 35788
rect -1854 35779 -1806 35784
rect -1974 35774 -1964 35775
rect -1960 35774 -1944 35776
rect -1842 35774 -1806 35777
rect -1655 35774 -1647 35786
rect -1642 35774 -1637 35868
rect -1619 35774 -1614 35868
rect -1530 35774 -1526 35868
rect -1506 35774 -1502 35868
rect -1482 35774 -1478 35868
rect -1458 35774 -1454 35868
rect -1434 35774 -1430 35868
rect -1410 35774 -1406 35868
rect -1386 35774 -1382 35868
rect -1362 35867 -1358 35868
rect -1362 35846 -1355 35867
rect -1338 35846 -1334 35868
rect -1314 35846 -1310 35868
rect -1290 35846 -1286 35868
rect -1266 35846 -1262 35868
rect -1242 35846 -1238 35868
rect -1218 35846 -1214 35868
rect -1194 35846 -1190 35868
rect -1170 35846 -1166 35868
rect -1146 35846 -1142 35868
rect -1122 35846 -1118 35868
rect -1098 35846 -1094 35868
rect -1074 35846 -1070 35868
rect -1050 35846 -1046 35868
rect -1026 35846 -1022 35868
rect -1002 35846 -998 35868
rect -978 35846 -974 35868
rect -954 35846 -950 35868
rect -930 35846 -926 35868
rect -917 35861 -912 35868
rect -906 35861 -902 35868
rect -907 35847 -902 35861
rect -906 35846 -902 35847
rect -882 35846 -878 35940
rect -875 35939 -861 35940
rect -858 35939 -851 35963
rect -858 35846 -854 35939
rect -834 35846 -830 35964
rect -810 35846 -806 35964
rect -786 35846 -782 35964
rect -762 35846 -758 35964
rect -738 35846 -734 35964
rect -714 35846 -710 35964
rect -690 35846 -686 35964
rect -666 35846 -662 35964
rect -642 35846 -638 35964
rect -618 35846 -614 35964
rect -594 35846 -590 35964
rect -570 35846 -566 35964
rect -546 35846 -542 35964
rect -522 35846 -518 35964
rect -498 35846 -494 35964
rect -474 35846 -470 35964
rect -450 35846 -446 35964
rect -426 35846 -422 35964
rect -402 35846 -398 35964
rect -378 35846 -374 35964
rect -354 35846 -350 35964
rect -330 35846 -326 35964
rect -306 35846 -302 35964
rect -282 35846 -278 35964
rect -258 35846 -254 35964
rect -234 35846 -230 35964
rect -210 35846 -206 35964
rect -186 35846 -182 35964
rect -162 35846 -158 35964
rect -138 35846 -134 35964
rect -114 35846 -110 35964
rect -90 35846 -86 35964
rect -66 35846 -62 35964
rect -42 35846 -38 35964
rect -18 35915 -14 35964
rect -18 35891 -11 35915
rect -18 35846 -14 35891
rect 6 35846 10 35964
rect 30 35846 34 35964
rect 54 35847 58 35964
rect 43 35846 77 35847
rect -1379 35844 77 35846
rect -1379 35843 -1365 35844
rect -1362 35819 -1355 35844
rect -1362 35774 -1358 35819
rect -1338 35775 -1334 35844
rect -1349 35774 -1315 35775
rect -2393 35772 -1315 35774
rect -2371 35750 -2366 35772
rect -2348 35750 -2343 35772
rect -2325 35760 -2317 35772
rect -2325 35750 -2320 35760
rect -2317 35758 -2309 35760
rect -2062 35759 -2032 35766
rect -2309 35750 -2301 35758
rect -2070 35752 -2062 35759
rect -2000 35754 -1992 35772
rect -1974 35770 -1944 35772
rect -1960 35769 -1944 35770
rect -1842 35768 -1806 35772
rect -1842 35761 -1798 35766
rect -1806 35759 -1798 35761
rect -1671 35760 -1663 35772
rect -1854 35757 -1842 35759
rect -1663 35758 -1655 35760
rect -2062 35750 -2036 35752
rect -2393 35748 -2036 35750
rect -2032 35750 -2012 35752
rect -2004 35750 -1974 35754
rect -1854 35752 -1806 35757
rect -1864 35750 -1796 35751
rect -1655 35750 -1647 35758
rect -1642 35750 -1637 35772
rect -1619 35750 -1614 35772
rect -1530 35750 -1526 35772
rect -1506 35750 -1502 35772
rect -1482 35750 -1478 35772
rect -1458 35750 -1454 35772
rect -1434 35750 -1430 35772
rect -1410 35750 -1406 35772
rect -1386 35750 -1382 35772
rect -1362 35750 -1358 35772
rect -1349 35765 -1344 35772
rect -1338 35765 -1334 35772
rect -1339 35751 -1334 35765
rect -1338 35750 -1334 35751
rect -1314 35750 -1310 35844
rect -1290 35750 -1286 35844
rect -1266 35750 -1262 35844
rect -1242 35750 -1238 35844
rect -1218 35750 -1214 35844
rect -1194 35750 -1190 35844
rect -1170 35750 -1166 35844
rect -1146 35750 -1142 35844
rect -1122 35750 -1118 35844
rect -1098 35750 -1094 35844
rect -1074 35750 -1070 35844
rect -1050 35750 -1046 35844
rect -1026 35750 -1022 35844
rect -1002 35750 -998 35844
rect -978 35750 -974 35844
rect -954 35750 -950 35844
rect -930 35750 -926 35844
rect -906 35750 -902 35844
rect -882 35795 -878 35844
rect -882 35771 -875 35795
rect -882 35750 -878 35771
rect -858 35750 -854 35844
rect -834 35750 -830 35844
rect -810 35750 -806 35844
rect -786 35750 -782 35844
rect -762 35750 -758 35844
rect -738 35750 -734 35844
rect -714 35750 -710 35844
rect -690 35750 -686 35844
rect -666 35750 -662 35844
rect -642 35750 -638 35844
rect -618 35750 -614 35844
rect -594 35750 -590 35844
rect -570 35750 -566 35844
rect -546 35750 -542 35844
rect -522 35750 -518 35844
rect -498 35750 -494 35844
rect -474 35750 -470 35844
rect -450 35750 -446 35844
rect -426 35750 -422 35844
rect -402 35750 -398 35844
rect -378 35750 -374 35844
rect -354 35750 -350 35844
rect -330 35750 -326 35844
rect -306 35750 -302 35844
rect -282 35750 -278 35844
rect -258 35750 -254 35844
rect -234 35750 -230 35844
rect -210 35750 -206 35844
rect -186 35750 -182 35844
rect -162 35750 -158 35844
rect -138 35750 -134 35844
rect -114 35750 -110 35844
rect -90 35750 -86 35844
rect -66 35750 -62 35844
rect -42 35750 -38 35844
rect -18 35750 -14 35844
rect 6 35750 10 35844
rect 30 35750 34 35844
rect 43 35837 48 35844
rect 54 35837 58 35844
rect 53 35823 58 35837
rect 54 35750 58 35823
rect 78 35771 82 35964
rect -2032 35748 75 35750
rect -2371 35702 -2366 35748
rect -2348 35702 -2343 35748
rect -2325 35744 -2320 35748
rect -2309 35746 -2301 35748
rect -2317 35744 -2309 35746
rect -2325 35732 -2317 35744
rect -2052 35742 -2036 35744
rect -2052 35740 -2032 35742
rect -2062 35734 -2032 35740
rect -2325 35702 -2320 35732
rect -2317 35730 -2309 35732
rect -2092 35718 -2062 35720
rect -2094 35714 -2062 35718
rect -2000 35702 -1992 35748
rect -1904 35741 -1874 35748
rect -1842 35741 -1806 35748
rect -1655 35746 -1647 35748
rect -1663 35744 -1655 35746
rect -1842 35734 -1680 35740
rect -1671 35732 -1663 35744
rect -1663 35730 -1655 35732
rect -1854 35718 -1806 35720
rect -1854 35714 -1680 35718
rect -1642 35702 -1637 35748
rect -1619 35702 -1614 35748
rect -1530 35702 -1526 35748
rect -1506 35702 -1502 35748
rect -1482 35702 -1478 35748
rect -1458 35702 -1454 35748
rect -1434 35702 -1430 35748
rect -1410 35702 -1406 35748
rect -1386 35702 -1382 35748
rect -1362 35702 -1358 35748
rect -1338 35702 -1334 35748
rect -1314 35702 -1310 35748
rect -1290 35702 -1286 35748
rect -1266 35702 -1262 35748
rect -1242 35702 -1238 35748
rect -1218 35702 -1214 35748
rect -1194 35702 -1190 35748
rect -1170 35702 -1166 35748
rect -1146 35702 -1142 35748
rect -1122 35702 -1118 35748
rect -1098 35702 -1094 35748
rect -1074 35702 -1070 35748
rect -1050 35702 -1046 35748
rect -1026 35702 -1022 35748
rect -1002 35702 -998 35748
rect -978 35702 -974 35748
rect -954 35702 -950 35748
rect -930 35702 -926 35748
rect -906 35702 -902 35748
rect -882 35702 -878 35748
rect -858 35702 -854 35748
rect -834 35702 -830 35748
rect -810 35702 -806 35748
rect -786 35702 -782 35748
rect -773 35717 -768 35727
rect -762 35717 -758 35748
rect -763 35703 -758 35717
rect -773 35702 -739 35703
rect -2393 35700 -739 35702
rect -2371 35678 -2366 35700
rect -2348 35678 -2343 35700
rect -2325 35678 -2320 35700
rect -2072 35698 -2036 35699
rect -2072 35692 -2054 35698
rect -2309 35684 -2301 35692
rect -2317 35678 -2309 35684
rect -2092 35683 -2062 35688
rect -2000 35679 -1992 35700
rect -1938 35699 -1906 35700
rect -1920 35698 -1906 35699
rect -1806 35692 -1680 35698
rect -1854 35683 -1806 35688
rect -1655 35684 -1647 35692
rect -1982 35679 -1966 35680
rect -2000 35678 -1966 35679
rect -1846 35678 -1806 35681
rect -1663 35678 -1655 35684
rect -1642 35678 -1637 35700
rect -1619 35678 -1614 35700
rect -1530 35678 -1526 35700
rect -1506 35678 -1502 35700
rect -1482 35678 -1478 35700
rect -1458 35678 -1454 35700
rect -1434 35678 -1430 35700
rect -1410 35679 -1406 35700
rect -1421 35678 -1387 35679
rect -2393 35676 -1387 35678
rect -2371 35654 -2366 35676
rect -2348 35654 -2343 35676
rect -2325 35654 -2320 35676
rect -2000 35674 -1966 35676
rect -2309 35656 -2301 35664
rect -2062 35663 -2054 35670
rect -2092 35656 -2084 35663
rect -2062 35656 -2026 35658
rect -2317 35654 -2309 35656
rect -2062 35654 -2012 35656
rect -2000 35654 -1992 35674
rect -1982 35673 -1966 35674
rect -1846 35672 -1806 35676
rect -1846 35665 -1798 35670
rect -1806 35663 -1798 35665
rect -1854 35661 -1846 35663
rect -1854 35656 -1806 35661
rect -1655 35656 -1647 35664
rect -1864 35654 -1796 35655
rect -1663 35654 -1655 35656
rect -1642 35654 -1637 35676
rect -1619 35654 -1614 35676
rect -1530 35654 -1526 35676
rect -1506 35654 -1502 35676
rect -1482 35654 -1478 35676
rect -1458 35654 -1454 35676
rect -1434 35654 -1430 35676
rect -1421 35669 -1416 35676
rect -1410 35669 -1406 35676
rect -1411 35655 -1406 35669
rect -1410 35654 -1406 35655
rect -1386 35654 -1382 35700
rect -1362 35654 -1358 35700
rect -1338 35654 -1334 35700
rect -1314 35699 -1310 35700
rect -1314 35675 -1307 35699
rect -1314 35654 -1310 35675
rect -1290 35654 -1286 35700
rect -1266 35655 -1262 35700
rect -1277 35654 -1243 35655
rect -2393 35652 -1243 35654
rect -2371 35606 -2366 35652
rect -2348 35606 -2343 35652
rect -2325 35606 -2320 35652
rect -2317 35648 -2309 35652
rect -2062 35648 -2054 35652
rect -2154 35644 -2138 35646
rect -2057 35644 -2054 35648
rect -2292 35638 -2054 35644
rect -2052 35638 -2044 35648
rect -2092 35622 -2062 35624
rect -2094 35618 -2062 35622
rect -2000 35606 -1992 35652
rect -1846 35645 -1806 35652
rect -1663 35648 -1655 35652
rect -1846 35638 -1680 35644
rect -1854 35622 -1806 35624
rect -1854 35618 -1680 35622
rect -1979 35606 -1945 35608
rect -1642 35606 -1637 35652
rect -1619 35606 -1614 35652
rect -1530 35606 -1526 35652
rect -1506 35606 -1502 35652
rect -1493 35621 -1488 35631
rect -1482 35621 -1478 35652
rect -1483 35607 -1478 35621
rect -1493 35606 -1459 35607
rect -2393 35604 -1459 35606
rect -2371 35558 -2366 35604
rect -2348 35558 -2343 35604
rect -2325 35558 -2320 35604
rect -2080 35603 -1906 35604
rect -2080 35602 -2036 35603
rect -2080 35596 -2054 35602
rect -2309 35588 -2301 35594
rect -2317 35578 -2309 35588
rect -2070 35587 -2040 35594
rect -2054 35579 -2040 35582
rect -2000 35577 -1992 35603
rect -1920 35602 -1906 35603
rect -1850 35596 -1846 35604
rect -1840 35596 -1792 35604
rect -1969 35584 -1966 35593
rect -1850 35589 -1802 35594
rect -1906 35587 -1802 35589
rect -1655 35588 -1647 35594
rect -1906 35586 -1850 35587
rect -1846 35579 -1802 35585
rect -1663 35578 -1655 35588
rect -1860 35577 -1798 35578
rect -2078 35570 -2070 35577
rect -2309 35560 -2301 35566
rect -2317 35558 -2309 35560
rect -2154 35558 -2145 35568
rect -2044 35567 -2040 35572
rect -2028 35570 -1945 35577
rect -1929 35570 -1794 35577
rect -2070 35560 -2040 35567
rect -2044 35558 -2028 35560
rect -2000 35558 -1992 35570
rect -1860 35569 -1798 35570
rect -1850 35560 -1802 35567
rect -1655 35560 -1647 35566
rect -1978 35558 -1942 35559
rect -1663 35558 -1655 35560
rect -1642 35558 -1637 35604
rect -1619 35558 -1614 35604
rect -1530 35558 -1526 35604
rect -1506 35558 -1502 35604
rect -1493 35597 -1488 35604
rect -1483 35583 -1478 35597
rect -1482 35558 -1478 35583
rect -1458 35558 -1454 35652
rect -1434 35558 -1430 35652
rect -1410 35558 -1406 35652
rect -1386 35603 -1382 35652
rect -1386 35579 -1379 35603
rect -1386 35558 -1382 35579
rect -1362 35558 -1358 35652
rect -1338 35558 -1334 35652
rect -1314 35558 -1310 35652
rect -1290 35558 -1286 35652
rect -1277 35645 -1272 35652
rect -1266 35645 -1262 35652
rect -1267 35631 -1262 35645
rect -1266 35558 -1262 35631
rect -1242 35579 -1238 35700
rect -2393 35556 -1245 35558
rect -2371 35462 -2366 35556
rect -2348 35462 -2343 35556
rect -2325 35518 -2320 35556
rect -2317 35550 -2309 35556
rect -2145 35552 -2138 35556
rect -2070 35552 -2054 35556
rect -2078 35543 -2054 35550
rect -2062 35518 -2032 35519
rect -2000 35518 -1992 35556
rect -1846 35552 -1802 35556
rect -1846 35542 -1792 35551
rect -1663 35550 -1655 35556
rect -1942 35520 -1937 35532
rect -1850 35529 -1822 35530
rect -1850 35525 -1802 35529
rect -2325 35510 -2317 35518
rect -2062 35516 -1961 35518
rect -2325 35490 -2320 35510
rect -2317 35502 -2309 35510
rect -2062 35503 -2040 35514
rect -2032 35509 -1961 35516
rect -1947 35510 -1942 35518
rect -1842 35516 -1794 35519
rect -2070 35498 -2022 35502
rect -2325 35476 -2317 35490
rect -2072 35482 -2032 35483
rect -2102 35476 -2032 35482
rect -2325 35462 -2320 35476
rect -2317 35474 -2309 35476
rect -2309 35462 -2301 35474
rect -2070 35467 -2062 35472
rect -2000 35462 -1992 35509
rect -1942 35508 -1937 35510
rect -1932 35500 -1927 35508
rect -1912 35505 -1896 35511
rect -1842 35503 -1802 35514
rect -1671 35510 -1663 35518
rect -1663 35502 -1655 35510
rect -1850 35498 -1680 35502
rect -1924 35484 -1921 35486
rect -1806 35476 -1680 35482
rect -1671 35476 -1663 35490
rect -1663 35474 -1655 35476
rect -1854 35467 -1806 35472
rect -1974 35462 -1964 35463
rect -1960 35462 -1944 35464
rect -1842 35462 -1806 35465
rect -1655 35462 -1647 35474
rect -1642 35462 -1637 35556
rect -1619 35462 -1614 35556
rect -1530 35462 -1526 35556
rect -1506 35462 -1502 35556
rect -1482 35462 -1478 35556
rect -1458 35555 -1454 35556
rect -1458 35534 -1451 35555
rect -1434 35534 -1430 35556
rect -1410 35534 -1406 35556
rect -1386 35534 -1382 35556
rect -1362 35534 -1358 35556
rect -1338 35534 -1334 35556
rect -1314 35534 -1310 35556
rect -1290 35534 -1286 35556
rect -1266 35534 -1262 35556
rect -1259 35555 -1245 35556
rect -1242 35555 -1235 35579
rect -1242 35534 -1238 35555
rect -1218 35534 -1214 35700
rect -1194 35534 -1190 35700
rect -1170 35534 -1166 35700
rect -1146 35534 -1142 35700
rect -1122 35535 -1118 35700
rect -1133 35534 -1099 35535
rect -1475 35532 -1099 35534
rect -1475 35531 -1461 35532
rect -1458 35507 -1451 35532
rect -1458 35462 -1454 35507
rect -1434 35462 -1430 35532
rect -1410 35462 -1406 35532
rect -1386 35462 -1382 35532
rect -1362 35463 -1358 35532
rect -1373 35462 -1339 35463
rect -2393 35460 -1339 35462
rect -2371 35438 -2366 35460
rect -2348 35438 -2343 35460
rect -2325 35448 -2317 35460
rect -2325 35438 -2320 35448
rect -2317 35446 -2309 35448
rect -2062 35447 -2032 35454
rect -2309 35438 -2301 35446
rect -2070 35440 -2062 35447
rect -2000 35442 -1992 35460
rect -1974 35458 -1944 35460
rect -1960 35457 -1944 35458
rect -1842 35456 -1806 35460
rect -1842 35449 -1798 35454
rect -1806 35447 -1798 35449
rect -1671 35448 -1663 35460
rect -1854 35445 -1842 35447
rect -1663 35446 -1655 35448
rect -2062 35438 -2036 35440
rect -2393 35436 -2036 35438
rect -2032 35438 -2012 35440
rect -2004 35438 -1974 35442
rect -1854 35440 -1806 35445
rect -1864 35438 -1796 35439
rect -1655 35438 -1647 35446
rect -1642 35438 -1637 35460
rect -1619 35438 -1614 35460
rect -1530 35438 -1526 35460
rect -1506 35438 -1502 35460
rect -1482 35438 -1478 35460
rect -1458 35438 -1454 35460
rect -1434 35438 -1430 35460
rect -1410 35438 -1406 35460
rect -1386 35438 -1382 35460
rect -1373 35453 -1368 35460
rect -1362 35453 -1358 35460
rect -1363 35439 -1358 35453
rect -1362 35438 -1358 35439
rect -1338 35438 -1334 35532
rect -1314 35438 -1310 35532
rect -1290 35438 -1286 35532
rect -1266 35438 -1262 35532
rect -1242 35438 -1238 35532
rect -1218 35438 -1214 35532
rect -1194 35438 -1190 35532
rect -1170 35438 -1166 35532
rect -1146 35438 -1142 35532
rect -1133 35525 -1128 35532
rect -1122 35525 -1118 35532
rect -1123 35511 -1118 35525
rect -1122 35438 -1118 35511
rect -1098 35459 -1094 35700
rect -2032 35436 -1101 35438
rect -2371 35390 -2366 35436
rect -2348 35390 -2343 35436
rect -2325 35432 -2320 35436
rect -2309 35434 -2301 35436
rect -2317 35432 -2309 35434
rect -2325 35420 -2317 35432
rect -2052 35430 -2036 35432
rect -2052 35428 -2032 35430
rect -2062 35422 -2032 35428
rect -2325 35390 -2320 35420
rect -2317 35418 -2309 35420
rect -2092 35406 -2062 35408
rect -2094 35402 -2062 35406
rect -2000 35390 -1992 35436
rect -1904 35429 -1874 35436
rect -1842 35429 -1806 35436
rect -1655 35434 -1647 35436
rect -1663 35432 -1655 35434
rect -1842 35422 -1680 35428
rect -1671 35420 -1663 35432
rect -1663 35418 -1655 35420
rect -1854 35406 -1806 35408
rect -1854 35402 -1680 35406
rect -1642 35390 -1637 35436
rect -1619 35390 -1614 35436
rect -1530 35390 -1526 35436
rect -1506 35390 -1502 35436
rect -1482 35390 -1478 35436
rect -1458 35390 -1454 35436
rect -1434 35390 -1430 35436
rect -1410 35390 -1406 35436
rect -1386 35390 -1382 35436
rect -1362 35390 -1358 35436
rect -1338 35390 -1334 35436
rect -1314 35390 -1310 35436
rect -1290 35390 -1286 35436
rect -1266 35390 -1262 35436
rect -1242 35390 -1238 35436
rect -1218 35390 -1214 35436
rect -1194 35390 -1190 35436
rect -1170 35390 -1166 35436
rect -1146 35390 -1142 35436
rect -1122 35390 -1118 35436
rect -1115 35435 -1101 35436
rect -1098 35435 -1091 35459
rect -1098 35390 -1094 35435
rect -1074 35390 -1070 35700
rect -1050 35390 -1046 35700
rect -1026 35390 -1022 35700
rect -1002 35390 -998 35700
rect -978 35390 -974 35700
rect -954 35390 -950 35700
rect -930 35390 -926 35700
rect -906 35390 -902 35700
rect -882 35390 -878 35700
rect -858 35390 -854 35700
rect -834 35390 -830 35700
rect -810 35390 -806 35700
rect -786 35390 -782 35700
rect -773 35693 -768 35700
rect -763 35679 -758 35693
rect -762 35390 -758 35679
rect -738 35651 -734 35748
rect -738 35630 -731 35651
rect -714 35630 -710 35748
rect -690 35630 -686 35748
rect -666 35630 -662 35748
rect -642 35630 -638 35748
rect -618 35630 -614 35748
rect -594 35630 -590 35748
rect -570 35630 -566 35748
rect -546 35630 -542 35748
rect -522 35630 -518 35748
rect -498 35630 -494 35748
rect -474 35630 -470 35748
rect -450 35630 -446 35748
rect -426 35630 -422 35748
rect -402 35630 -398 35748
rect -378 35630 -374 35748
rect -354 35630 -350 35748
rect -330 35630 -326 35748
rect -306 35630 -302 35748
rect -282 35630 -278 35748
rect -258 35630 -254 35748
rect -234 35630 -230 35748
rect -210 35630 -206 35748
rect -186 35630 -182 35748
rect -162 35630 -158 35748
rect -138 35630 -134 35748
rect -114 35630 -110 35748
rect -90 35630 -86 35748
rect -66 35630 -62 35748
rect -42 35630 -38 35748
rect -18 35630 -14 35748
rect 6 35630 10 35748
rect 30 35630 34 35748
rect 54 35630 58 35748
rect 61 35747 75 35748
rect 78 35747 85 35771
rect 78 35630 82 35747
rect 102 35630 106 35964
rect 126 35630 130 35964
rect 150 35630 154 35964
rect 174 35630 178 35964
rect 198 35630 202 35964
rect 222 35630 226 35964
rect 246 35630 250 35964
rect 270 35630 274 35964
rect 294 35630 298 35964
rect 318 35630 322 35964
rect 342 35630 346 35964
rect 366 35630 370 35964
rect 390 35630 394 35964
rect 414 35630 418 35964
rect 438 35630 442 35964
rect 462 35630 466 35964
rect 486 35630 490 35964
rect 510 35630 514 35964
rect 534 35630 538 35964
rect 558 35630 562 35964
rect 582 35630 586 35964
rect 606 35630 610 35964
rect 630 35630 634 35964
rect 654 35630 658 35964
rect 678 35630 682 35964
rect 702 35630 706 35964
rect 726 35630 730 35964
rect 750 35630 754 35964
rect 757 35963 771 35964
rect 774 35963 781 36011
rect 774 35630 778 35963
rect 798 35630 802 36012
rect 822 35630 826 36012
rect 846 35630 850 36012
rect 870 35630 874 36012
rect 894 35630 898 36012
rect 907 35813 912 35823
rect 918 35813 922 36012
rect 917 35799 922 35813
rect 907 35789 912 35799
rect 917 35775 922 35789
rect 918 35630 922 35775
rect 942 35747 946 36012
rect 942 35726 949 35747
rect 966 35726 970 36012
rect 990 35726 994 36012
rect 1014 35726 1018 36012
rect 1038 35726 1042 36012
rect 1051 36005 1056 36012
rect 1062 36005 1066 36012
rect 1061 35991 1066 36005
rect 1062 35726 1066 35991
rect 1086 35939 1090 36108
rect 1086 35915 1093 35939
rect 1086 35726 1090 35915
rect 1110 35726 1114 36108
rect 1134 35726 1138 36108
rect 1158 35726 1162 36108
rect 1182 35726 1186 36108
rect 1206 35726 1210 36108
rect 1230 35726 1234 36108
rect 1243 36101 1248 36108
rect 1254 36101 1258 36108
rect 1253 36087 1258 36101
rect 1243 36077 1248 36087
rect 1253 36063 1258 36077
rect 1243 35957 1248 35967
rect 1254 35957 1258 36063
rect 1253 35943 1258 35957
rect 1243 35933 1248 35943
rect 1253 35919 1258 35933
rect 1254 35726 1258 35919
rect 1267 35813 1272 35823
rect 1277 35799 1282 35813
rect 1267 35741 1272 35751
rect 1278 35741 1282 35799
rect 1277 35727 1282 35741
rect 1291 35737 1299 35741
rect 1285 35727 1291 35737
rect 1267 35726 1299 35727
rect 925 35724 1299 35726
rect 925 35723 939 35724
rect 942 35699 949 35724
rect 942 35630 946 35699
rect 966 35630 970 35724
rect 990 35630 994 35724
rect 1014 35630 1018 35724
rect 1038 35630 1042 35724
rect 1062 35630 1066 35724
rect 1086 35630 1090 35724
rect 1110 35630 1114 35724
rect 1134 35630 1138 35724
rect 1158 35630 1162 35724
rect 1182 35630 1186 35724
rect 1206 35630 1210 35724
rect 1230 35630 1234 35724
rect 1254 35630 1258 35724
rect 1267 35717 1272 35724
rect 1285 35723 1299 35724
rect 1277 35703 1282 35717
rect 1278 35630 1282 35703
rect 1291 35630 1299 35631
rect -755 35628 1299 35630
rect -755 35627 -741 35628
rect -738 35603 -731 35628
rect -738 35390 -734 35603
rect -714 35390 -710 35628
rect -690 35390 -686 35628
rect -666 35390 -662 35628
rect -642 35390 -638 35628
rect -629 35429 -624 35439
rect -618 35429 -614 35628
rect -619 35415 -614 35429
rect -629 35405 -624 35415
rect -618 35405 -614 35415
rect -619 35391 -614 35405
rect -629 35390 -595 35391
rect -2393 35388 -595 35390
rect -2371 35366 -2366 35388
rect -2348 35366 -2343 35388
rect -2325 35366 -2320 35388
rect -2072 35386 -2036 35387
rect -2072 35380 -2054 35386
rect -2309 35372 -2301 35380
rect -2317 35366 -2309 35372
rect -2092 35371 -2062 35376
rect -2000 35367 -1992 35388
rect -1938 35387 -1906 35388
rect -1920 35386 -1906 35387
rect -1806 35380 -1680 35386
rect -1854 35371 -1806 35376
rect -1655 35372 -1647 35380
rect -1982 35367 -1966 35368
rect -2000 35366 -1966 35367
rect -1846 35366 -1806 35369
rect -1663 35366 -1655 35372
rect -1642 35366 -1637 35388
rect -1619 35366 -1614 35388
rect -1530 35366 -1526 35388
rect -1506 35366 -1502 35388
rect -1482 35366 -1478 35388
rect -1458 35366 -1454 35388
rect -1434 35366 -1430 35388
rect -1410 35366 -1406 35388
rect -1386 35366 -1382 35388
rect -1362 35366 -1358 35388
rect -1338 35387 -1334 35388
rect -2393 35364 -1341 35366
rect -2371 35342 -2366 35364
rect -2348 35342 -2343 35364
rect -2325 35342 -2320 35364
rect -2000 35362 -1966 35364
rect -2309 35344 -2301 35352
rect -2062 35351 -2054 35358
rect -2092 35344 -2084 35351
rect -2062 35344 -2026 35346
rect -2317 35342 -2309 35344
rect -2062 35342 -2012 35344
rect -2000 35342 -1992 35362
rect -1982 35361 -1966 35362
rect -1846 35360 -1806 35364
rect -1846 35353 -1798 35358
rect -1806 35351 -1798 35353
rect -1854 35349 -1846 35351
rect -1854 35344 -1806 35349
rect -1655 35344 -1647 35352
rect -1864 35342 -1796 35343
rect -1663 35342 -1655 35344
rect -1642 35342 -1637 35364
rect -1619 35342 -1614 35364
rect -1530 35342 -1526 35364
rect -1506 35342 -1502 35364
rect -1482 35342 -1478 35364
rect -1458 35342 -1454 35364
rect -1434 35342 -1430 35364
rect -1410 35342 -1406 35364
rect -1386 35342 -1382 35364
rect -1362 35342 -1358 35364
rect -1355 35363 -1341 35364
rect -1338 35363 -1331 35387
rect -1338 35342 -1334 35363
rect -1314 35342 -1310 35388
rect -1290 35342 -1286 35388
rect -1266 35342 -1262 35388
rect -1242 35342 -1238 35388
rect -1218 35342 -1214 35388
rect -1194 35342 -1190 35388
rect -1170 35342 -1166 35388
rect -1146 35342 -1142 35388
rect -1122 35342 -1118 35388
rect -1098 35342 -1094 35388
rect -1074 35342 -1070 35388
rect -1050 35342 -1046 35388
rect -1026 35342 -1022 35388
rect -1002 35342 -998 35388
rect -978 35342 -974 35388
rect -954 35342 -950 35388
rect -930 35342 -926 35388
rect -906 35342 -902 35388
rect -882 35342 -878 35388
rect -858 35342 -854 35388
rect -834 35342 -830 35388
rect -810 35342 -806 35388
rect -786 35342 -782 35388
rect -762 35342 -758 35388
rect -738 35342 -734 35388
rect -714 35342 -710 35388
rect -690 35342 -686 35388
rect -666 35342 -662 35388
rect -642 35342 -638 35388
rect -629 35381 -624 35388
rect -619 35367 -614 35381
rect -618 35342 -614 35367
rect -594 35363 -590 35628
rect -2393 35340 -597 35342
rect -2371 35294 -2366 35340
rect -2348 35294 -2343 35340
rect -2325 35294 -2320 35340
rect -2317 35336 -2309 35340
rect -2062 35336 -2054 35340
rect -2154 35332 -2138 35334
rect -2057 35332 -2054 35336
rect -2292 35326 -2054 35332
rect -2052 35326 -2044 35336
rect -2092 35310 -2062 35312
rect -2094 35306 -2062 35310
rect -2000 35294 -1992 35340
rect -1846 35333 -1806 35340
rect -1663 35336 -1655 35340
rect -1846 35326 -1680 35332
rect -1854 35310 -1806 35312
rect -1854 35306 -1680 35310
rect -1642 35294 -1637 35340
rect -1619 35294 -1614 35340
rect -1530 35294 -1526 35340
rect -1506 35294 -1502 35340
rect -1482 35294 -1478 35340
rect -1458 35294 -1454 35340
rect -1434 35294 -1430 35340
rect -1410 35294 -1406 35340
rect -1386 35294 -1382 35340
rect -1362 35294 -1358 35340
rect -1338 35294 -1334 35340
rect -1314 35294 -1310 35340
rect -1290 35294 -1286 35340
rect -1266 35294 -1262 35340
rect -1242 35294 -1238 35340
rect -1218 35294 -1214 35340
rect -1194 35294 -1190 35340
rect -1170 35294 -1166 35340
rect -1146 35294 -1142 35340
rect -1122 35294 -1118 35340
rect -1098 35294 -1094 35340
rect -1074 35294 -1070 35340
rect -1050 35294 -1046 35340
rect -1026 35294 -1022 35340
rect -1002 35294 -998 35340
rect -978 35294 -974 35340
rect -954 35294 -950 35340
rect -930 35294 -926 35340
rect -906 35294 -902 35340
rect -882 35294 -878 35340
rect -858 35294 -854 35340
rect -834 35294 -830 35340
rect -810 35294 -806 35340
rect -786 35294 -782 35340
rect -762 35294 -758 35340
rect -738 35294 -734 35340
rect -714 35294 -710 35340
rect -690 35294 -686 35340
rect -666 35294 -662 35340
rect -642 35294 -638 35340
rect -618 35294 -614 35340
rect -611 35339 -597 35340
rect -2393 35292 -597 35294
rect -2371 35270 -2366 35292
rect -2348 35270 -2343 35292
rect -2325 35270 -2320 35292
rect -2072 35290 -2036 35291
rect -2072 35284 -2054 35290
rect -2309 35276 -2301 35284
rect -2317 35270 -2309 35276
rect -2092 35275 -2062 35280
rect -2000 35271 -1992 35292
rect -1938 35291 -1906 35292
rect -1920 35290 -1906 35291
rect -1806 35284 -1680 35290
rect -1854 35275 -1806 35280
rect -1655 35276 -1647 35284
rect -1982 35271 -1966 35272
rect -2000 35270 -1966 35271
rect -1846 35270 -1806 35273
rect -1663 35270 -1655 35276
rect -1642 35270 -1637 35292
rect -1619 35270 -1614 35292
rect -1530 35270 -1526 35292
rect -1506 35270 -1502 35292
rect -1482 35270 -1478 35292
rect -1458 35270 -1454 35292
rect -1434 35270 -1430 35292
rect -1410 35270 -1406 35292
rect -1386 35270 -1382 35292
rect -1362 35270 -1358 35292
rect -1338 35270 -1334 35292
rect -1314 35270 -1310 35292
rect -1290 35270 -1286 35292
rect -1266 35270 -1262 35292
rect -1242 35270 -1238 35292
rect -1218 35270 -1214 35292
rect -1194 35270 -1190 35292
rect -1170 35270 -1166 35292
rect -1146 35270 -1142 35292
rect -1122 35270 -1118 35292
rect -1098 35270 -1094 35292
rect -1074 35270 -1070 35292
rect -1050 35270 -1046 35292
rect -1026 35270 -1022 35292
rect -1002 35270 -998 35292
rect -978 35270 -974 35292
rect -954 35270 -950 35292
rect -930 35270 -926 35292
rect -906 35270 -902 35292
rect -882 35270 -878 35292
rect -858 35270 -854 35292
rect -834 35270 -830 35292
rect -810 35270 -806 35292
rect -786 35270 -782 35292
rect -762 35270 -758 35292
rect -738 35270 -734 35292
rect -714 35270 -710 35292
rect -690 35270 -686 35292
rect -666 35270 -662 35292
rect -642 35270 -638 35292
rect -618 35270 -614 35292
rect -611 35291 -597 35292
rect -594 35291 -587 35363
rect -594 35270 -590 35291
rect -570 35270 -566 35628
rect -546 35270 -542 35628
rect -522 35270 -518 35628
rect -498 35270 -494 35628
rect -474 35270 -470 35628
rect -461 35549 -456 35559
rect -450 35549 -446 35628
rect -451 35535 -446 35549
rect -461 35357 -456 35367
rect -450 35357 -446 35535
rect -451 35343 -446 35357
rect -450 35271 -446 35343
rect -426 35483 -422 35628
rect -426 35459 -419 35483
rect -426 35291 -422 35459
rect -461 35270 -429 35271
rect -2393 35268 -429 35270
rect -2371 35246 -2366 35268
rect -2348 35246 -2343 35268
rect -2325 35246 -2320 35268
rect -2000 35266 -1966 35268
rect -2309 35248 -2301 35256
rect -2062 35255 -2054 35262
rect -2092 35248 -2084 35255
rect -2062 35248 -2026 35250
rect -2317 35246 -2309 35248
rect -2062 35246 -2012 35248
rect -2000 35246 -1992 35266
rect -1982 35265 -1966 35266
rect -1846 35264 -1806 35268
rect -1846 35257 -1798 35262
rect -1806 35255 -1798 35257
rect -1854 35253 -1846 35255
rect -1854 35248 -1806 35253
rect -1655 35248 -1647 35256
rect -1864 35246 -1796 35247
rect -1663 35246 -1655 35248
rect -1642 35246 -1637 35268
rect -1619 35246 -1614 35268
rect -1530 35246 -1526 35268
rect -1506 35246 -1502 35268
rect -1482 35246 -1478 35268
rect -1458 35246 -1454 35268
rect -1434 35246 -1430 35268
rect -1410 35246 -1406 35268
rect -1386 35246 -1382 35268
rect -1362 35246 -1358 35268
rect -1338 35246 -1334 35268
rect -1314 35246 -1310 35268
rect -1290 35246 -1286 35268
rect -1266 35246 -1262 35268
rect -1242 35246 -1238 35268
rect -1218 35246 -1214 35268
rect -1194 35246 -1190 35268
rect -1170 35246 -1166 35268
rect -1146 35246 -1142 35268
rect -1122 35246 -1118 35268
rect -1098 35246 -1094 35268
rect -1074 35246 -1070 35268
rect -1050 35246 -1046 35268
rect -1026 35246 -1022 35268
rect -1002 35246 -998 35268
rect -978 35246 -974 35268
rect -954 35246 -950 35268
rect -930 35246 -926 35268
rect -906 35246 -902 35268
rect -882 35246 -878 35268
rect -858 35246 -854 35268
rect -834 35246 -830 35268
rect -810 35246 -806 35268
rect -786 35246 -782 35268
rect -762 35246 -758 35268
rect -738 35246 -734 35268
rect -714 35246 -710 35268
rect -690 35246 -686 35268
rect -666 35246 -662 35268
rect -642 35246 -638 35268
rect -618 35246 -614 35268
rect -594 35246 -590 35268
rect -570 35246 -566 35268
rect -546 35246 -542 35268
rect -522 35246 -518 35268
rect -498 35246 -494 35268
rect -474 35246 -470 35268
rect -461 35261 -456 35268
rect -450 35261 -446 35268
rect -443 35267 -429 35268
rect -426 35267 -419 35291
rect -451 35247 -446 35261
rect -450 35246 -446 35247
rect -426 35246 -422 35267
rect -402 35246 -398 35628
rect -378 35246 -374 35628
rect -354 35246 -350 35628
rect -330 35246 -326 35628
rect -306 35246 -302 35628
rect -282 35246 -278 35628
rect -258 35247 -254 35628
rect -269 35246 -235 35247
rect -2393 35244 -235 35246
rect -2371 35198 -2366 35244
rect -2348 35198 -2343 35244
rect -2325 35198 -2320 35244
rect -2317 35240 -2309 35244
rect -2062 35240 -2054 35244
rect -2154 35236 -2138 35238
rect -2057 35236 -2054 35240
rect -2292 35230 -2054 35236
rect -2052 35230 -2044 35240
rect -2092 35214 -2062 35216
rect -2094 35210 -2062 35214
rect -2000 35198 -1992 35244
rect -1846 35237 -1806 35244
rect -1663 35240 -1655 35244
rect -1846 35230 -1680 35236
rect -1854 35214 -1806 35216
rect -1854 35210 -1680 35214
rect -1642 35198 -1637 35244
rect -1619 35198 -1614 35244
rect -1530 35198 -1526 35244
rect -1506 35198 -1502 35244
rect -1482 35198 -1478 35244
rect -1458 35198 -1454 35244
rect -1434 35198 -1430 35244
rect -1410 35198 -1406 35244
rect -1386 35198 -1382 35244
rect -1362 35198 -1358 35244
rect -1338 35198 -1334 35244
rect -1314 35198 -1310 35244
rect -1290 35198 -1286 35244
rect -1266 35198 -1262 35244
rect -1242 35198 -1238 35244
rect -1218 35198 -1214 35244
rect -1194 35198 -1190 35244
rect -1170 35198 -1166 35244
rect -1146 35198 -1142 35244
rect -1122 35198 -1118 35244
rect -1098 35198 -1094 35244
rect -1074 35198 -1070 35244
rect -1050 35198 -1046 35244
rect -1026 35198 -1022 35244
rect -1002 35198 -998 35244
rect -978 35198 -974 35244
rect -954 35198 -950 35244
rect -930 35198 -926 35244
rect -906 35198 -902 35244
rect -882 35198 -878 35244
rect -858 35198 -854 35244
rect -834 35198 -830 35244
rect -810 35198 -806 35244
rect -786 35198 -782 35244
rect -762 35198 -758 35244
rect -738 35198 -734 35244
rect -714 35198 -710 35244
rect -690 35198 -686 35244
rect -666 35198 -662 35244
rect -642 35198 -638 35244
rect -618 35198 -614 35244
rect -594 35198 -590 35244
rect -570 35198 -566 35244
rect -546 35198 -542 35244
rect -522 35198 -518 35244
rect -498 35198 -494 35244
rect -474 35198 -470 35244
rect -450 35198 -446 35244
rect -426 35198 -422 35244
rect -402 35198 -398 35244
rect -378 35198 -374 35244
rect -354 35198 -350 35244
rect -330 35198 -326 35244
rect -306 35198 -302 35244
rect -282 35198 -278 35244
rect -269 35237 -264 35244
rect -258 35237 -254 35244
rect -259 35223 -254 35237
rect -258 35198 -254 35223
rect -234 35198 -230 35628
rect -210 35198 -206 35628
rect -186 35198 -182 35628
rect -162 35198 -158 35628
rect -138 35198 -134 35628
rect -114 35198 -110 35628
rect -90 35198 -86 35628
rect -66 35198 -62 35628
rect -42 35198 -38 35628
rect -18 35198 -14 35628
rect 6 35198 10 35628
rect 30 35198 34 35628
rect 54 35198 58 35628
rect 78 35198 82 35628
rect 102 35198 106 35628
rect 126 35198 130 35628
rect 150 35198 154 35628
rect 163 35501 168 35511
rect 174 35501 178 35628
rect 173 35487 178 35501
rect 163 35477 168 35487
rect 173 35463 178 35477
rect 174 35198 178 35463
rect 198 35435 202 35628
rect 198 35414 205 35435
rect 222 35414 226 35628
rect 246 35414 250 35628
rect 270 35414 274 35628
rect 294 35414 298 35628
rect 318 35414 322 35628
rect 342 35414 346 35628
rect 366 35414 370 35628
rect 390 35414 394 35628
rect 414 35414 418 35628
rect 438 35414 442 35628
rect 462 35414 466 35628
rect 486 35414 490 35628
rect 510 35414 514 35628
rect 534 35414 538 35628
rect 558 35414 562 35628
rect 582 35414 586 35628
rect 606 35414 610 35628
rect 630 35414 634 35628
rect 654 35414 658 35628
rect 678 35414 682 35628
rect 702 35414 706 35628
rect 726 35414 730 35628
rect 750 35414 754 35628
rect 774 35414 778 35628
rect 798 35414 802 35628
rect 822 35414 826 35628
rect 846 35414 850 35628
rect 870 35414 874 35628
rect 894 35414 898 35628
rect 918 35414 922 35628
rect 942 35414 946 35628
rect 966 35414 970 35628
rect 990 35414 994 35628
rect 1014 35414 1018 35628
rect 1038 35414 1042 35628
rect 1062 35414 1066 35628
rect 1086 35414 1090 35628
rect 1110 35414 1114 35628
rect 1134 35414 1138 35628
rect 1158 35414 1162 35628
rect 1182 35414 1186 35628
rect 1206 35414 1210 35628
rect 1230 35414 1234 35628
rect 1254 35414 1258 35628
rect 1278 35414 1282 35628
rect 1285 35627 1299 35628
rect 1291 35621 1296 35627
rect 1301 35607 1306 35621
rect 1302 35414 1306 35607
rect 1315 35501 1320 35511
rect 1325 35487 1330 35501
rect 1326 35414 1330 35487
rect 1339 35414 1347 35415
rect 181 35412 1347 35414
rect 181 35411 195 35412
rect 198 35387 205 35412
rect 198 35198 202 35387
rect 211 35213 216 35223
rect 222 35213 226 35412
rect 221 35199 226 35213
rect 211 35198 245 35199
rect -2393 35196 245 35198
rect -2371 35174 -2366 35196
rect -2348 35174 -2343 35196
rect -2325 35174 -2320 35196
rect -2072 35194 -2036 35195
rect -2072 35188 -2054 35194
rect -2309 35180 -2301 35188
rect -2317 35174 -2309 35180
rect -2092 35179 -2062 35184
rect -2000 35175 -1992 35196
rect -1938 35195 -1906 35196
rect -1920 35194 -1906 35195
rect -1806 35188 -1680 35194
rect -1854 35179 -1806 35184
rect -1655 35180 -1647 35188
rect -1982 35175 -1966 35176
rect -2000 35174 -1966 35175
rect -1846 35174 -1806 35177
rect -1663 35174 -1655 35180
rect -1642 35174 -1637 35196
rect -1619 35174 -1614 35196
rect -1530 35174 -1526 35196
rect -1506 35174 -1502 35196
rect -1482 35174 -1478 35196
rect -1458 35174 -1454 35196
rect -1434 35174 -1430 35196
rect -1410 35174 -1406 35196
rect -1386 35174 -1382 35196
rect -1362 35174 -1358 35196
rect -1338 35174 -1334 35196
rect -1314 35174 -1310 35196
rect -1290 35174 -1286 35196
rect -1266 35174 -1262 35196
rect -1242 35174 -1238 35196
rect -1218 35174 -1214 35196
rect -1194 35174 -1190 35196
rect -1170 35174 -1166 35196
rect -1146 35174 -1142 35196
rect -1122 35174 -1118 35196
rect -1098 35174 -1094 35196
rect -1074 35174 -1070 35196
rect -1050 35174 -1046 35196
rect -1026 35174 -1022 35196
rect -1002 35174 -998 35196
rect -978 35174 -974 35196
rect -954 35174 -950 35196
rect -930 35174 -926 35196
rect -906 35174 -902 35196
rect -882 35174 -878 35196
rect -858 35174 -854 35196
rect -834 35174 -830 35196
rect -810 35174 -806 35196
rect -786 35174 -782 35196
rect -762 35174 -758 35196
rect -738 35174 -734 35196
rect -714 35174 -710 35196
rect -690 35174 -686 35196
rect -666 35174 -662 35196
rect -642 35174 -638 35196
rect -618 35174 -614 35196
rect -594 35174 -590 35196
rect -570 35174 -566 35196
rect -546 35174 -542 35196
rect -522 35174 -518 35196
rect -498 35174 -494 35196
rect -474 35174 -470 35196
rect -450 35174 -446 35196
rect -426 35195 -422 35196
rect -2393 35172 -429 35174
rect -2371 35150 -2366 35172
rect -2348 35150 -2343 35172
rect -2325 35150 -2320 35172
rect -2000 35170 -1966 35172
rect -2309 35152 -2301 35160
rect -2062 35159 -2054 35166
rect -2092 35152 -2084 35159
rect -2062 35152 -2026 35154
rect -2317 35150 -2309 35152
rect -2062 35150 -2012 35152
rect -2000 35150 -1992 35170
rect -1982 35169 -1966 35170
rect -1846 35168 -1806 35172
rect -1846 35161 -1798 35166
rect -1806 35159 -1798 35161
rect -1854 35157 -1846 35159
rect -1854 35152 -1806 35157
rect -1655 35152 -1647 35160
rect -1864 35150 -1796 35151
rect -1663 35150 -1655 35152
rect -1642 35150 -1637 35172
rect -1619 35150 -1614 35172
rect -1530 35150 -1526 35172
rect -1506 35150 -1502 35172
rect -1482 35150 -1478 35172
rect -1458 35150 -1454 35172
rect -1434 35150 -1430 35172
rect -1410 35150 -1406 35172
rect -1386 35150 -1382 35172
rect -1362 35150 -1358 35172
rect -1338 35150 -1334 35172
rect -1314 35150 -1310 35172
rect -1290 35150 -1286 35172
rect -1266 35150 -1262 35172
rect -1242 35150 -1238 35172
rect -1218 35150 -1214 35172
rect -1194 35150 -1190 35172
rect -1170 35150 -1166 35172
rect -1146 35150 -1142 35172
rect -1122 35150 -1118 35172
rect -1098 35150 -1094 35172
rect -1074 35150 -1070 35172
rect -1050 35150 -1046 35172
rect -1026 35150 -1022 35172
rect -1002 35150 -998 35172
rect -978 35150 -974 35172
rect -954 35150 -950 35172
rect -930 35150 -926 35172
rect -906 35150 -902 35172
rect -882 35150 -878 35172
rect -858 35150 -854 35172
rect -834 35150 -830 35172
rect -810 35150 -806 35172
rect -786 35150 -782 35172
rect -762 35150 -758 35172
rect -738 35150 -734 35172
rect -714 35150 -710 35172
rect -690 35150 -686 35172
rect -666 35150 -662 35172
rect -642 35150 -638 35172
rect -618 35150 -614 35172
rect -594 35150 -590 35172
rect -570 35150 -566 35172
rect -546 35150 -542 35172
rect -522 35150 -518 35172
rect -498 35150 -494 35172
rect -474 35150 -470 35172
rect -450 35150 -446 35172
rect -443 35171 -429 35172
rect -426 35171 -419 35195
rect -426 35150 -422 35171
rect -402 35150 -398 35196
rect -378 35150 -374 35196
rect -354 35150 -350 35196
rect -330 35150 -326 35196
rect -306 35150 -302 35196
rect -282 35150 -278 35196
rect -258 35150 -254 35196
rect -234 35171 -230 35196
rect -2393 35148 -237 35150
rect -2371 35102 -2366 35148
rect -2348 35102 -2343 35148
rect -2325 35102 -2320 35148
rect -2317 35144 -2309 35148
rect -2062 35144 -2054 35148
rect -2154 35140 -2138 35142
rect -2057 35140 -2054 35144
rect -2292 35134 -2054 35140
rect -2052 35134 -2044 35144
rect -2092 35118 -2062 35120
rect -2094 35114 -2062 35118
rect -2000 35102 -1992 35148
rect -1846 35141 -1806 35148
rect -1663 35144 -1655 35148
rect -1846 35134 -1680 35140
rect -1854 35118 -1806 35120
rect -1854 35114 -1680 35118
rect -1642 35102 -1637 35148
rect -1619 35102 -1614 35148
rect -1530 35102 -1526 35148
rect -1506 35102 -1502 35148
rect -1482 35102 -1478 35148
rect -1458 35102 -1454 35148
rect -1434 35102 -1430 35148
rect -1410 35102 -1406 35148
rect -1386 35102 -1382 35148
rect -1362 35102 -1358 35148
rect -1338 35102 -1334 35148
rect -1314 35102 -1310 35148
rect -1290 35102 -1286 35148
rect -1266 35102 -1262 35148
rect -1242 35102 -1238 35148
rect -1218 35102 -1214 35148
rect -1194 35102 -1190 35148
rect -1170 35102 -1166 35148
rect -1157 35117 -1152 35127
rect -1146 35117 -1142 35148
rect -1147 35103 -1142 35117
rect -1157 35102 -1123 35103
rect -2393 35100 -1123 35102
rect -2371 35078 -2366 35100
rect -2348 35078 -2343 35100
rect -2325 35078 -2320 35100
rect -2072 35098 -2036 35099
rect -2072 35092 -2054 35098
rect -2309 35084 -2301 35092
rect -2317 35078 -2309 35084
rect -2092 35083 -2062 35088
rect -2000 35079 -1992 35100
rect -1938 35099 -1906 35100
rect -1920 35098 -1906 35099
rect -1806 35092 -1680 35098
rect -1854 35083 -1806 35088
rect -1655 35084 -1647 35092
rect -1982 35079 -1966 35080
rect -2000 35078 -1966 35079
rect -1846 35078 -1806 35081
rect -1663 35078 -1655 35084
rect -1642 35078 -1637 35100
rect -1619 35078 -1614 35100
rect -1530 35078 -1526 35100
rect -1506 35078 -1502 35100
rect -1482 35078 -1478 35100
rect -1458 35078 -1454 35100
rect -1434 35078 -1430 35100
rect -1410 35078 -1406 35100
rect -1386 35078 -1382 35100
rect -1362 35078 -1358 35100
rect -1338 35078 -1334 35100
rect -1314 35078 -1310 35100
rect -1290 35078 -1286 35100
rect -1266 35078 -1262 35100
rect -1242 35078 -1238 35100
rect -1218 35078 -1214 35100
rect -1194 35078 -1190 35100
rect -1170 35078 -1166 35100
rect -1157 35093 -1152 35100
rect -1147 35079 -1142 35093
rect -1146 35078 -1142 35079
rect -1122 35078 -1118 35148
rect -1098 35078 -1094 35148
rect -1074 35078 -1070 35148
rect -1050 35078 -1046 35148
rect -1026 35078 -1022 35148
rect -1002 35078 -998 35148
rect -978 35078 -974 35148
rect -954 35078 -950 35148
rect -930 35078 -926 35148
rect -906 35078 -902 35148
rect -882 35078 -878 35148
rect -858 35078 -854 35148
rect -834 35078 -830 35148
rect -810 35078 -806 35148
rect -786 35078 -782 35148
rect -762 35078 -758 35148
rect -738 35078 -734 35148
rect -714 35078 -710 35148
rect -690 35078 -686 35148
rect -666 35078 -662 35148
rect -642 35078 -638 35148
rect -618 35078 -614 35148
rect -594 35078 -590 35148
rect -570 35078 -566 35148
rect -546 35078 -542 35148
rect -522 35078 -518 35148
rect -498 35078 -494 35148
rect -474 35078 -470 35148
rect -450 35078 -446 35148
rect -426 35078 -422 35148
rect -402 35078 -398 35148
rect -378 35078 -374 35148
rect -354 35078 -350 35148
rect -330 35078 -326 35148
rect -306 35078 -302 35148
rect -282 35078 -278 35148
rect -258 35078 -254 35148
rect -251 35147 -237 35148
rect -234 35147 -227 35171
rect -234 35078 -230 35147
rect -210 35078 -206 35196
rect -186 35078 -182 35196
rect -173 35165 -168 35175
rect -162 35165 -158 35196
rect -163 35151 -158 35165
rect -162 35078 -158 35151
rect -138 35099 -134 35196
rect -2393 35076 -141 35078
rect -2371 35054 -2366 35076
rect -2348 35054 -2343 35076
rect -2325 35054 -2320 35076
rect -2000 35074 -1966 35076
rect -2309 35056 -2301 35064
rect -2062 35063 -2054 35070
rect -2092 35056 -2084 35063
rect -2062 35056 -2026 35058
rect -2317 35054 -2309 35056
rect -2062 35054 -2012 35056
rect -2000 35054 -1992 35074
rect -1982 35073 -1966 35074
rect -1846 35072 -1806 35076
rect -1846 35065 -1798 35070
rect -1806 35063 -1798 35065
rect -1854 35061 -1846 35063
rect -1854 35056 -1806 35061
rect -1655 35056 -1647 35064
rect -1864 35054 -1796 35055
rect -1663 35054 -1655 35056
rect -1642 35054 -1637 35076
rect -1619 35054 -1614 35076
rect -1530 35054 -1526 35076
rect -1506 35054 -1502 35076
rect -1482 35054 -1478 35076
rect -1458 35054 -1454 35076
rect -1434 35054 -1430 35076
rect -1410 35054 -1406 35076
rect -1386 35054 -1382 35076
rect -1362 35054 -1358 35076
rect -1338 35054 -1334 35076
rect -1314 35054 -1310 35076
rect -1290 35054 -1286 35076
rect -1266 35054 -1262 35076
rect -1242 35054 -1238 35076
rect -1218 35054 -1214 35076
rect -1194 35054 -1190 35076
rect -1170 35054 -1166 35076
rect -1146 35054 -1142 35076
rect -1122 35054 -1118 35076
rect -1098 35054 -1094 35076
rect -1074 35054 -1070 35076
rect -1050 35054 -1046 35076
rect -1026 35054 -1022 35076
rect -1002 35054 -998 35076
rect -978 35054 -974 35076
rect -954 35054 -950 35076
rect -930 35054 -926 35076
rect -906 35054 -902 35076
rect -882 35054 -878 35076
rect -858 35054 -854 35076
rect -834 35054 -830 35076
rect -810 35054 -806 35076
rect -786 35054 -782 35076
rect -762 35054 -758 35076
rect -738 35054 -734 35076
rect -714 35054 -710 35076
rect -690 35054 -686 35076
rect -666 35054 -662 35076
rect -642 35054 -638 35076
rect -618 35054 -614 35076
rect -594 35054 -590 35076
rect -570 35054 -566 35076
rect -546 35054 -542 35076
rect -522 35054 -518 35076
rect -498 35054 -494 35076
rect -474 35054 -470 35076
rect -450 35054 -446 35076
rect -426 35054 -422 35076
rect -402 35054 -398 35076
rect -378 35054 -374 35076
rect -354 35054 -350 35076
rect -330 35054 -326 35076
rect -306 35054 -302 35076
rect -282 35054 -278 35076
rect -258 35054 -254 35076
rect -234 35054 -230 35076
rect -210 35054 -206 35076
rect -186 35054 -182 35076
rect -162 35055 -158 35076
rect -155 35075 -141 35076
rect -138 35075 -131 35099
rect -173 35054 -139 35055
rect -2393 35052 -139 35054
rect -2371 35006 -2366 35052
rect -2348 35006 -2343 35052
rect -2325 35006 -2320 35052
rect -2317 35048 -2309 35052
rect -2062 35048 -2054 35052
rect -2154 35044 -2138 35046
rect -2057 35044 -2054 35048
rect -2292 35038 -2054 35044
rect -2052 35038 -2044 35048
rect -2092 35022 -2062 35024
rect -2094 35018 -2062 35022
rect -2000 35006 -1992 35052
rect -1846 35045 -1806 35052
rect -1663 35048 -1655 35052
rect -1846 35038 -1680 35044
rect -1854 35022 -1806 35024
rect -1854 35018 -1680 35022
rect -1642 35006 -1637 35052
rect -1619 35006 -1614 35052
rect -1530 35006 -1526 35052
rect -1506 35006 -1502 35052
rect -1482 35006 -1478 35052
rect -1458 35006 -1454 35052
rect -1434 35006 -1430 35052
rect -1410 35006 -1406 35052
rect -1386 35006 -1382 35052
rect -1362 35006 -1358 35052
rect -1338 35006 -1334 35052
rect -1314 35006 -1310 35052
rect -1290 35006 -1286 35052
rect -1266 35006 -1262 35052
rect -1242 35006 -1238 35052
rect -1218 35006 -1214 35052
rect -1194 35006 -1190 35052
rect -1170 35006 -1166 35052
rect -1146 35006 -1142 35052
rect -1122 35051 -1118 35052
rect -2393 35004 -1125 35006
rect -2371 34982 -2366 35004
rect -2348 34982 -2343 35004
rect -2325 34982 -2320 35004
rect -2072 35002 -2036 35003
rect -2072 34996 -2054 35002
rect -2309 34988 -2301 34996
rect -2317 34982 -2309 34988
rect -2092 34987 -2062 34992
rect -2000 34983 -1992 35004
rect -1938 35003 -1906 35004
rect -1920 35002 -1906 35003
rect -1806 34996 -1680 35002
rect -1854 34987 -1806 34992
rect -1655 34988 -1647 34996
rect -1982 34983 -1966 34984
rect -2000 34982 -1966 34983
rect -1846 34982 -1806 34985
rect -1663 34982 -1655 34988
rect -1642 34982 -1637 35004
rect -1619 34982 -1614 35004
rect -1530 34982 -1526 35004
rect -1506 34982 -1502 35004
rect -1482 34982 -1478 35004
rect -1458 34982 -1454 35004
rect -1434 34982 -1430 35004
rect -1410 34982 -1406 35004
rect -1386 34982 -1382 35004
rect -1362 34982 -1358 35004
rect -1338 34982 -1334 35004
rect -1314 34982 -1310 35004
rect -1290 34982 -1286 35004
rect -1266 34982 -1262 35004
rect -1242 34982 -1238 35004
rect -1218 34982 -1214 35004
rect -1194 34982 -1190 35004
rect -1170 34982 -1166 35004
rect -1146 34982 -1142 35004
rect -1139 35003 -1125 35004
rect -1122 35003 -1115 35051
rect -1122 34982 -1118 35003
rect -1098 34982 -1094 35052
rect -1074 34982 -1070 35052
rect -1050 34982 -1046 35052
rect -1026 34982 -1022 35052
rect -1002 34982 -998 35052
rect -978 34982 -974 35052
rect -954 34982 -950 35052
rect -930 34982 -926 35052
rect -906 34982 -902 35052
rect -882 34982 -878 35052
rect -858 34982 -854 35052
rect -834 34982 -830 35052
rect -810 34982 -806 35052
rect -786 34982 -782 35052
rect -762 34982 -758 35052
rect -738 34982 -734 35052
rect -714 34982 -710 35052
rect -690 34982 -686 35052
rect -666 34982 -662 35052
rect -642 34982 -638 35052
rect -618 34982 -614 35052
rect -594 34982 -590 35052
rect -570 34982 -566 35052
rect -546 34982 -542 35052
rect -522 34982 -518 35052
rect -498 34982 -494 35052
rect -474 34982 -470 35052
rect -450 34982 -446 35052
rect -426 34982 -422 35052
rect -402 34982 -398 35052
rect -378 34982 -374 35052
rect -354 34982 -350 35052
rect -330 34982 -326 35052
rect -306 34982 -302 35052
rect -282 34982 -278 35052
rect -258 34982 -254 35052
rect -234 34982 -230 35052
rect -210 34982 -206 35052
rect -186 34982 -182 35052
rect -173 35045 -168 35052
rect -162 35045 -158 35052
rect -163 35031 -158 35045
rect -162 34983 -158 35031
rect -173 34982 -139 34983
rect -2393 34980 -139 34982
rect -2371 34958 -2366 34980
rect -2348 34958 -2343 34980
rect -2325 34958 -2320 34980
rect -2000 34978 -1966 34980
rect -2309 34960 -2301 34968
rect -2062 34967 -2054 34974
rect -2092 34960 -2084 34967
rect -2062 34960 -2026 34962
rect -2317 34958 -2309 34960
rect -2062 34958 -2012 34960
rect -2000 34958 -1992 34978
rect -1982 34977 -1966 34978
rect -1846 34976 -1806 34980
rect -1846 34969 -1798 34974
rect -1806 34967 -1798 34969
rect -1854 34965 -1846 34967
rect -1854 34960 -1806 34965
rect -1655 34960 -1647 34968
rect -1864 34958 -1796 34959
rect -1663 34958 -1655 34960
rect -1642 34958 -1637 34980
rect -1619 34958 -1614 34980
rect -1530 34958 -1526 34980
rect -1506 34958 -1502 34980
rect -1482 34958 -1478 34980
rect -1458 34958 -1454 34980
rect -1434 34958 -1430 34980
rect -1410 34958 -1406 34980
rect -1386 34958 -1382 34980
rect -1362 34958 -1358 34980
rect -1338 34958 -1334 34980
rect -1314 34958 -1310 34980
rect -1290 34958 -1286 34980
rect -1266 34958 -1262 34980
rect -1242 34958 -1238 34980
rect -1218 34958 -1214 34980
rect -1194 34958 -1190 34980
rect -1170 34958 -1166 34980
rect -1146 34958 -1142 34980
rect -1122 34959 -1118 34980
rect -1133 34958 -1099 34959
rect -2393 34956 -1099 34958
rect -2371 34886 -2366 34956
rect -2348 34886 -2343 34956
rect -2325 34886 -2320 34956
rect -2317 34952 -2309 34956
rect -2062 34952 -2054 34956
rect -2154 34948 -2138 34950
rect -2057 34948 -2054 34952
rect -2292 34942 -2054 34948
rect -2052 34942 -2044 34952
rect -2092 34926 -2062 34928
rect -2094 34922 -2062 34926
rect -2309 34892 -2301 34898
rect -2317 34886 -2309 34892
rect -2000 34886 -1992 34956
rect -1846 34949 -1806 34956
rect -1663 34952 -1655 34956
rect -1846 34942 -1680 34948
rect -1854 34926 -1806 34928
rect -1854 34922 -1680 34926
rect -1655 34892 -1647 34898
rect -1663 34886 -1655 34892
rect -1642 34886 -1637 34956
rect -1619 34886 -1614 34956
rect -1530 34886 -1526 34956
rect -1506 34886 -1502 34956
rect -1482 34886 -1478 34956
rect -1458 34886 -1454 34956
rect -1434 34886 -1430 34956
rect -1410 34886 -1406 34956
rect -1386 34886 -1382 34956
rect -1362 34886 -1358 34956
rect -1338 34886 -1334 34956
rect -1314 34886 -1310 34956
rect -1290 34886 -1286 34956
rect -1266 34886 -1262 34956
rect -1242 34886 -1238 34956
rect -1218 34886 -1214 34956
rect -1194 34886 -1190 34956
rect -1170 34886 -1166 34956
rect -1146 34886 -1142 34956
rect -1133 34949 -1128 34956
rect -1122 34949 -1118 34956
rect -1123 34935 -1118 34949
rect -1122 34886 -1118 34935
rect -1098 34886 -1094 34980
rect -1074 34886 -1070 34980
rect -1050 34886 -1046 34980
rect -1026 34886 -1022 34980
rect -1002 34886 -998 34980
rect -978 34886 -974 34980
rect -954 34886 -950 34980
rect -930 34886 -926 34980
rect -906 34886 -902 34980
rect -882 34886 -878 34980
rect -858 34886 -854 34980
rect -834 34886 -830 34980
rect -810 34886 -806 34980
rect -786 34886 -782 34980
rect -762 34886 -758 34980
rect -738 34886 -734 34980
rect -714 34886 -710 34980
rect -690 34886 -686 34980
rect -666 34886 -662 34980
rect -642 34886 -638 34980
rect -618 34886 -614 34980
rect -594 34886 -590 34980
rect -570 34886 -566 34980
rect -546 34886 -542 34980
rect -522 34886 -518 34980
rect -498 34886 -494 34980
rect -474 34886 -470 34980
rect -450 34886 -446 34980
rect -426 34886 -422 34980
rect -402 34886 -398 34980
rect -378 34886 -374 34980
rect -354 34886 -350 34980
rect -330 34886 -326 34980
rect -306 34886 -302 34980
rect -282 34886 -278 34980
rect -258 34886 -254 34980
rect -234 34886 -230 34980
rect -210 34886 -206 34980
rect -186 34886 -182 34980
rect -173 34973 -168 34980
rect -162 34973 -158 34980
rect -138 34979 -134 35075
rect -163 34959 -158 34973
rect -149 34969 -141 34973
rect -155 34959 -149 34969
rect -162 34886 -158 34959
rect -138 34955 -131 34979
rect -138 34907 -134 34955
rect -2393 34884 -141 34886
rect -2371 34790 -2366 34884
rect -2348 34790 -2343 34884
rect -2325 34822 -2320 34884
rect -2317 34882 -2309 34884
rect -2000 34883 -1966 34884
rect -2000 34882 -1982 34883
rect -1663 34882 -1655 34884
rect -2028 34874 -2018 34876
rect -2309 34864 -2301 34870
rect -2091 34864 -2061 34871
rect -2317 34854 -2309 34864
rect -2044 34862 -2028 34864
rect -2026 34862 -2014 34874
rect -2084 34856 -2061 34862
rect -2044 34860 -2014 34862
rect -2292 34846 -2054 34855
rect -2325 34814 -2317 34822
rect -2325 34794 -2320 34814
rect -2317 34806 -2309 34814
rect -2325 34790 -2317 34794
rect -2000 34790 -1992 34882
rect -1982 34881 -1966 34882
rect -1980 34864 -1932 34871
rect -1655 34864 -1647 34870
rect -1846 34846 -1680 34855
rect -1663 34854 -1655 34864
rect -1671 34814 -1663 34822
rect -1663 34806 -1655 34814
rect -1671 34790 -1663 34794
rect -1642 34790 -1637 34884
rect -1619 34790 -1614 34884
rect -1530 34790 -1526 34884
rect -1506 34790 -1502 34884
rect -1482 34790 -1478 34884
rect -1458 34790 -1454 34884
rect -1434 34790 -1430 34884
rect -1410 34790 -1406 34884
rect -1386 34790 -1382 34884
rect -1362 34790 -1358 34884
rect -1338 34790 -1334 34884
rect -1314 34790 -1310 34884
rect -1290 34790 -1286 34884
rect -1266 34790 -1262 34884
rect -1242 34790 -1238 34884
rect -1218 34790 -1214 34884
rect -1194 34790 -1190 34884
rect -1170 34790 -1166 34884
rect -1146 34790 -1142 34884
rect -1122 34790 -1118 34884
rect -1098 34883 -1094 34884
rect -1098 34859 -1091 34883
rect -1098 34790 -1094 34859
rect -1074 34790 -1070 34884
rect -1050 34790 -1046 34884
rect -1026 34790 -1022 34884
rect -1002 34790 -998 34884
rect -989 34805 -984 34815
rect -978 34805 -974 34884
rect -979 34791 -974 34805
rect -989 34790 -955 34791
rect -2393 34788 -955 34790
rect -2371 34742 -2366 34788
rect -2348 34742 -2343 34788
rect -2325 34780 -2317 34788
rect -2018 34787 -2004 34788
rect -2000 34787 -1992 34788
rect -2072 34786 -1928 34787
rect -2072 34780 -2053 34786
rect -2325 34764 -2320 34780
rect -2317 34778 -2309 34780
rect -2309 34766 -2301 34778
rect -2092 34771 -2062 34776
rect -2317 34764 -2309 34766
rect -2325 34752 -2317 34764
rect -2098 34758 -2096 34769
rect -2092 34758 -2084 34771
rect -2000 34770 -1992 34786
rect -1972 34780 -1928 34786
rect -1924 34780 -1918 34788
rect -1671 34780 -1663 34788
rect -1663 34778 -1655 34780
rect -2083 34760 -2062 34769
rect -2027 34768 -1992 34770
rect -2018 34760 -2002 34768
rect -2000 34760 -1992 34768
rect -2100 34753 -2096 34758
rect -2083 34753 -2053 34758
rect -2003 34756 -1990 34760
rect -1972 34758 -1964 34767
rect -1928 34766 -1924 34769
rect -1655 34766 -1647 34778
rect -1663 34764 -1655 34766
rect -2325 34742 -2320 34752
rect -2317 34750 -2309 34752
rect -2309 34742 -2301 34750
rect -2004 34746 -2003 34756
rect -2062 34742 -2012 34744
rect -2000 34742 -1992 34756
rect -1972 34753 -1924 34758
rect -1864 34753 -1796 34759
rect -1671 34752 -1663 34764
rect -1663 34750 -1655 34752
rect -1864 34742 -1796 34743
rect -1655 34742 -1647 34750
rect -1642 34742 -1637 34788
rect -1619 34742 -1614 34788
rect -1530 34742 -1526 34788
rect -1506 34742 -1502 34788
rect -1482 34742 -1478 34788
rect -1458 34742 -1454 34788
rect -1434 34742 -1430 34788
rect -1410 34743 -1406 34788
rect -1421 34742 -1387 34743
rect -2393 34740 -1387 34742
rect -2371 34694 -2366 34740
rect -2348 34694 -2343 34740
rect -2325 34736 -2320 34740
rect -2309 34738 -2301 34740
rect -2317 34736 -2309 34738
rect -2325 34724 -2317 34736
rect -2325 34694 -2320 34724
rect -2317 34722 -2309 34724
rect -2092 34710 -2062 34712
rect -2094 34706 -2062 34710
rect -2000 34694 -1992 34740
rect -1655 34738 -1647 34740
rect -1663 34736 -1655 34738
rect -1671 34724 -1663 34736
rect -1663 34722 -1655 34724
rect -1854 34710 -1806 34712
rect -1854 34706 -1680 34710
rect -1642 34694 -1637 34740
rect -1619 34694 -1614 34740
rect -1530 34694 -1526 34740
rect -1506 34694 -1502 34740
rect -1482 34694 -1478 34740
rect -1458 34694 -1454 34740
rect -1434 34694 -1430 34740
rect -1421 34733 -1416 34740
rect -1410 34733 -1406 34740
rect -1411 34719 -1406 34733
rect -1410 34694 -1406 34719
rect -1386 34694 -1382 34788
rect -1362 34694 -1358 34788
rect -1338 34694 -1334 34788
rect -1314 34694 -1310 34788
rect -1290 34694 -1286 34788
rect -1266 34694 -1262 34788
rect -1242 34694 -1238 34788
rect -1218 34694 -1214 34788
rect -1194 34694 -1190 34788
rect -1170 34694 -1166 34788
rect -1157 34709 -1152 34719
rect -1146 34709 -1142 34788
rect -1147 34695 -1142 34709
rect -1157 34694 -1123 34695
rect -2393 34692 -1123 34694
rect -2371 34670 -2366 34692
rect -2348 34670 -2343 34692
rect -2325 34670 -2320 34692
rect -2072 34690 -2036 34691
rect -2072 34684 -2054 34690
rect -2309 34676 -2301 34684
rect -2317 34670 -2309 34676
rect -2092 34675 -2062 34680
rect -2000 34671 -1992 34692
rect -1938 34691 -1906 34692
rect -1920 34690 -1906 34691
rect -1806 34684 -1680 34690
rect -1854 34675 -1806 34680
rect -1655 34676 -1647 34684
rect -1982 34671 -1966 34672
rect -2000 34670 -1966 34671
rect -1846 34670 -1806 34673
rect -1663 34670 -1655 34676
rect -1642 34670 -1637 34692
rect -1619 34670 -1614 34692
rect -1530 34670 -1526 34692
rect -1506 34670 -1502 34692
rect -1482 34670 -1478 34692
rect -1458 34670 -1454 34692
rect -1434 34670 -1430 34692
rect -1410 34670 -1406 34692
rect -1386 34670 -1382 34692
rect -1362 34670 -1358 34692
rect -1338 34670 -1334 34692
rect -1314 34670 -1310 34692
rect -1290 34670 -1286 34692
rect -1266 34670 -1262 34692
rect -1242 34670 -1238 34692
rect -1218 34670 -1214 34692
rect -1194 34670 -1190 34692
rect -1170 34670 -1166 34692
rect -1157 34685 -1152 34692
rect -1147 34671 -1142 34685
rect -1146 34670 -1142 34671
rect -1122 34670 -1118 34788
rect -1098 34670 -1094 34788
rect -1074 34670 -1070 34788
rect -1050 34670 -1046 34788
rect -1026 34670 -1022 34788
rect -1002 34670 -998 34788
rect -989 34781 -984 34788
rect -979 34767 -974 34781
rect -978 34670 -974 34767
rect -954 34739 -950 34884
rect -941 34757 -936 34767
rect -930 34757 -926 34884
rect -931 34743 -926 34757
rect -954 34718 -947 34739
rect -930 34718 -926 34743
rect -906 34718 -902 34884
rect -882 34718 -878 34884
rect -858 34718 -854 34884
rect -834 34718 -830 34884
rect -821 34829 -816 34839
rect -810 34829 -806 34884
rect -811 34815 -806 34829
rect -810 34718 -806 34815
rect -786 34763 -782 34884
rect -786 34739 -779 34763
rect -786 34718 -782 34739
rect -762 34718 -758 34884
rect -738 34718 -734 34884
rect -714 34718 -710 34884
rect -690 34718 -686 34884
rect -666 34718 -662 34884
rect -642 34718 -638 34884
rect -618 34718 -614 34884
rect -594 34718 -590 34884
rect -570 34718 -566 34884
rect -546 34718 -542 34884
rect -522 34718 -518 34884
rect -498 34718 -494 34884
rect -474 34718 -470 34884
rect -450 34718 -446 34884
rect -426 34718 -422 34884
rect -402 34718 -398 34884
rect -378 34718 -374 34884
rect -354 34718 -350 34884
rect -330 34718 -326 34884
rect -306 34718 -302 34884
rect -282 34718 -278 34884
rect -258 34718 -254 34884
rect -234 34718 -230 34884
rect -210 34718 -206 34884
rect -186 34718 -182 34884
rect -162 34718 -158 34884
rect -155 34883 -141 34884
rect -138 34883 -131 34907
rect -138 34718 -134 34883
rect -114 34718 -110 35196
rect -90 34718 -86 35196
rect -66 34718 -62 35196
rect -42 34718 -38 35196
rect -18 34718 -14 35196
rect 6 34718 10 35196
rect 30 34718 34 35196
rect 54 34718 58 35196
rect 78 34718 82 35196
rect 102 35031 106 35196
rect 91 35030 125 35031
rect 126 35030 130 35196
rect 150 35030 154 35196
rect 174 35030 178 35196
rect 198 35030 202 35196
rect 211 35189 216 35196
rect 221 35175 226 35189
rect 222 35030 226 35175
rect 246 35147 250 35412
rect 246 35126 253 35147
rect 270 35126 274 35412
rect 294 35126 298 35412
rect 318 35126 322 35412
rect 342 35126 346 35412
rect 366 35126 370 35412
rect 390 35126 394 35412
rect 414 35126 418 35412
rect 438 35126 442 35412
rect 462 35126 466 35412
rect 486 35126 490 35412
rect 510 35126 514 35412
rect 534 35126 538 35412
rect 558 35126 562 35412
rect 582 35126 586 35412
rect 606 35126 610 35412
rect 630 35126 634 35412
rect 654 35126 658 35412
rect 678 35126 682 35412
rect 702 35126 706 35412
rect 726 35126 730 35412
rect 750 35126 754 35412
rect 774 35126 778 35412
rect 798 35126 802 35412
rect 822 35126 826 35412
rect 846 35126 850 35412
rect 870 35319 874 35412
rect 859 35318 893 35319
rect 894 35318 898 35412
rect 918 35318 922 35412
rect 942 35318 946 35412
rect 966 35318 970 35412
rect 990 35318 994 35412
rect 1014 35318 1018 35412
rect 1038 35318 1042 35412
rect 1062 35318 1066 35412
rect 1086 35318 1090 35412
rect 1110 35318 1114 35412
rect 1134 35318 1138 35412
rect 1158 35318 1162 35412
rect 1182 35318 1186 35412
rect 1206 35318 1210 35412
rect 1230 35318 1234 35412
rect 1254 35318 1258 35412
rect 1278 35318 1282 35412
rect 1302 35318 1306 35412
rect 1326 35318 1330 35412
rect 1333 35411 1347 35412
rect 1339 35405 1344 35411
rect 1349 35391 1354 35405
rect 1339 35333 1344 35343
rect 1350 35333 1354 35391
rect 1349 35319 1354 35333
rect 1363 35329 1371 35333
rect 1357 35319 1363 35329
rect 1339 35318 1371 35319
rect 859 35316 1371 35318
rect 859 35309 864 35316
rect 870 35309 874 35316
rect 869 35295 874 35309
rect 859 35285 864 35295
rect 869 35271 874 35285
rect 870 35126 874 35271
rect 894 35243 898 35316
rect 894 35222 901 35243
rect 918 35222 922 35316
rect 942 35222 946 35316
rect 966 35222 970 35316
rect 990 35222 994 35316
rect 1014 35222 1018 35316
rect 1038 35222 1042 35316
rect 1062 35222 1066 35316
rect 1086 35222 1090 35316
rect 1110 35222 1114 35316
rect 1134 35222 1138 35316
rect 1158 35222 1162 35316
rect 1182 35222 1186 35316
rect 1206 35222 1210 35316
rect 1230 35222 1234 35316
rect 1254 35222 1258 35316
rect 1278 35222 1282 35316
rect 1302 35222 1306 35316
rect 1326 35222 1330 35316
rect 1339 35309 1344 35316
rect 1357 35315 1371 35316
rect 1349 35295 1354 35309
rect 1350 35222 1354 35295
rect 1363 35222 1371 35223
rect 877 35220 1371 35222
rect 877 35219 891 35220
rect 894 35195 901 35220
rect 894 35126 898 35195
rect 918 35126 922 35220
rect 942 35126 946 35220
rect 966 35126 970 35220
rect 990 35126 994 35220
rect 1014 35126 1018 35220
rect 1038 35126 1042 35220
rect 1062 35126 1066 35220
rect 1086 35126 1090 35220
rect 1110 35126 1114 35220
rect 1134 35126 1138 35220
rect 1158 35126 1162 35220
rect 1182 35126 1186 35220
rect 1206 35126 1210 35220
rect 1230 35126 1234 35220
rect 1254 35126 1258 35220
rect 1278 35126 1282 35220
rect 1302 35126 1306 35220
rect 1326 35126 1330 35220
rect 1350 35126 1354 35220
rect 1357 35219 1371 35220
rect 1363 35213 1368 35219
rect 1373 35199 1378 35213
rect 1363 35141 1368 35151
rect 1374 35141 1378 35199
rect 1373 35127 1378 35141
rect 1387 35137 1395 35141
rect 1381 35127 1387 35137
rect 1363 35126 1395 35127
rect 229 35124 1395 35126
rect 229 35123 243 35124
rect 246 35099 253 35124
rect 246 35030 250 35099
rect 270 35030 274 35124
rect 294 35030 298 35124
rect 318 35030 322 35124
rect 342 35030 346 35124
rect 366 35030 370 35124
rect 390 35030 394 35124
rect 414 35030 418 35124
rect 438 35030 442 35124
rect 462 35030 466 35124
rect 486 35030 490 35124
rect 510 35030 514 35124
rect 534 35030 538 35124
rect 558 35030 562 35124
rect 582 35030 586 35124
rect 606 35030 610 35124
rect 630 35030 634 35124
rect 654 35030 658 35124
rect 678 35030 682 35124
rect 702 35030 706 35124
rect 726 35030 730 35124
rect 750 35030 754 35124
rect 774 35030 778 35124
rect 798 35030 802 35124
rect 822 35030 826 35124
rect 846 35030 850 35124
rect 870 35030 874 35124
rect 894 35030 898 35124
rect 918 35030 922 35124
rect 942 35030 946 35124
rect 966 35030 970 35124
rect 990 35030 994 35124
rect 1014 35030 1018 35124
rect 1038 35030 1042 35124
rect 1062 35030 1066 35124
rect 1086 35030 1090 35124
rect 1110 35030 1114 35124
rect 1134 35030 1138 35124
rect 1158 35030 1162 35124
rect 1182 35030 1186 35124
rect 1206 35030 1210 35124
rect 1230 35030 1234 35124
rect 1254 35030 1258 35124
rect 1278 35030 1282 35124
rect 1302 35030 1306 35124
rect 1326 35030 1330 35124
rect 1350 35030 1354 35124
rect 1363 35117 1368 35124
rect 1381 35123 1395 35124
rect 1373 35103 1378 35117
rect 1363 35069 1368 35079
rect 1374 35069 1378 35103
rect 1373 35055 1378 35069
rect 1387 35065 1395 35069
rect 1381 35055 1387 35065
rect 1363 35030 1395 35031
rect 91 35028 1395 35030
rect 91 35021 96 35028
rect 102 35021 106 35028
rect 101 35007 106 35021
rect 91 34997 96 35007
rect 101 34983 106 34997
rect 102 34718 106 34983
rect 126 34955 130 35028
rect 126 34907 133 34955
rect 126 34718 130 34907
rect 150 34718 154 35028
rect 174 34718 178 35028
rect 198 34718 202 35028
rect 222 34718 226 35028
rect 246 34718 250 35028
rect 270 34718 274 35028
rect 294 34718 298 35028
rect 318 34718 322 35028
rect 342 34718 346 35028
rect 366 34718 370 35028
rect 390 34718 394 35028
rect 414 34718 418 35028
rect 438 34718 442 35028
rect 462 34718 466 35028
rect 486 34718 490 35028
rect 510 34718 514 35028
rect 534 34718 538 35028
rect 558 34718 562 35028
rect 582 34718 586 35028
rect 606 34718 610 35028
rect 630 34718 634 35028
rect 654 34718 658 35028
rect 678 34718 682 35028
rect 702 34718 706 35028
rect 726 34718 730 35028
rect 750 34718 754 35028
rect 774 34718 778 35028
rect 798 34718 802 35028
rect 811 34901 816 34911
rect 822 34901 826 35028
rect 821 34887 826 34901
rect 811 34877 816 34887
rect 821 34863 826 34877
rect 822 34718 826 34863
rect 846 34835 850 35028
rect 846 34814 853 34835
rect 870 34814 874 35028
rect 894 34814 898 35028
rect 918 34814 922 35028
rect 942 34814 946 35028
rect 966 34814 970 35028
rect 990 34814 994 35028
rect 1014 34814 1018 35028
rect 1038 34814 1042 35028
rect 1062 34814 1066 35028
rect 1086 34814 1090 35028
rect 1110 34814 1114 35028
rect 1134 34814 1138 35028
rect 1158 34814 1162 35028
rect 1182 34814 1186 35028
rect 1206 34814 1210 35028
rect 1230 34814 1234 35028
rect 1254 34814 1258 35028
rect 1278 34814 1282 35028
rect 1302 34814 1306 35028
rect 1326 34814 1330 35028
rect 1350 34814 1354 35028
rect 1363 35021 1368 35028
rect 1381 35027 1395 35028
rect 1373 35007 1378 35021
rect 1374 34814 1378 35007
rect 1387 34901 1392 34911
rect 1397 34887 1402 34901
rect 1398 34814 1402 34887
rect 1411 34814 1419 34815
rect 829 34812 1419 34814
rect 829 34811 843 34812
rect 846 34787 853 34812
rect 846 34718 850 34787
rect 870 34718 874 34812
rect 894 34718 898 34812
rect 918 34718 922 34812
rect 942 34718 946 34812
rect 966 34718 970 34812
rect 990 34718 994 34812
rect 1014 34718 1018 34812
rect 1038 34718 1042 34812
rect 1062 34718 1066 34812
rect 1086 34718 1090 34812
rect 1110 34718 1114 34812
rect 1134 34718 1138 34812
rect 1158 34718 1162 34812
rect 1182 34718 1186 34812
rect 1206 34718 1210 34812
rect 1230 34718 1234 34812
rect 1254 34718 1258 34812
rect 1278 34718 1282 34812
rect 1302 34718 1306 34812
rect 1326 34718 1330 34812
rect 1350 34718 1354 34812
rect 1374 34718 1378 34812
rect 1398 34718 1402 34812
rect 1405 34811 1419 34812
rect 1411 34805 1416 34811
rect 1421 34791 1426 34805
rect 1422 34718 1426 34791
rect 1435 34718 1443 34719
rect -971 34716 1443 34718
rect -971 34715 -957 34716
rect -954 34691 -947 34716
rect -954 34670 -950 34691
rect -930 34670 -926 34716
rect -906 34691 -902 34716
rect -2393 34668 -909 34670
rect -2371 34646 -2366 34668
rect -2348 34646 -2343 34668
rect -2325 34646 -2320 34668
rect -2000 34666 -1966 34668
rect -2309 34648 -2301 34656
rect -2062 34655 -2054 34662
rect -2092 34648 -2084 34655
rect -2062 34648 -2026 34650
rect -2317 34646 -2309 34648
rect -2062 34646 -2012 34648
rect -2000 34646 -1992 34666
rect -1982 34665 -1966 34666
rect -1846 34664 -1806 34668
rect -1846 34657 -1798 34662
rect -1806 34655 -1798 34657
rect -1854 34653 -1846 34655
rect -1854 34648 -1806 34653
rect -1655 34648 -1647 34656
rect -1864 34646 -1796 34647
rect -1663 34646 -1655 34648
rect -1642 34646 -1637 34668
rect -1619 34646 -1614 34668
rect -1530 34646 -1526 34668
rect -1506 34646 -1502 34668
rect -1482 34646 -1478 34668
rect -1458 34646 -1454 34668
rect -1434 34646 -1430 34668
rect -1410 34646 -1406 34668
rect -1386 34667 -1382 34668
rect -2393 34644 -1389 34646
rect -2371 34574 -2366 34644
rect -2348 34574 -2343 34644
rect -2325 34574 -2320 34644
rect -2317 34640 -2309 34644
rect -2062 34640 -2054 34644
rect -2154 34636 -2138 34638
rect -2057 34636 -2054 34640
rect -2292 34630 -2054 34636
rect -2052 34630 -2044 34640
rect -2092 34614 -2062 34616
rect -2094 34610 -2062 34614
rect -2309 34580 -2301 34586
rect -2317 34574 -2309 34580
rect -2000 34574 -1992 34644
rect -1846 34637 -1806 34644
rect -1663 34640 -1655 34644
rect -1846 34630 -1680 34636
rect -1854 34614 -1806 34616
rect -1854 34610 -1680 34614
rect -1655 34580 -1647 34586
rect -1663 34574 -1655 34580
rect -1642 34574 -1637 34644
rect -1619 34574 -1614 34644
rect -1530 34574 -1526 34644
rect -1506 34574 -1502 34644
rect -1482 34574 -1478 34644
rect -1458 34574 -1454 34644
rect -1434 34574 -1430 34644
rect -1410 34574 -1406 34644
rect -1403 34643 -1389 34644
rect -1386 34643 -1379 34667
rect -1386 34574 -1382 34643
rect -1362 34574 -1358 34668
rect -1338 34574 -1334 34668
rect -1314 34574 -1310 34668
rect -1290 34574 -1286 34668
rect -1266 34574 -1262 34668
rect -1242 34574 -1238 34668
rect -1218 34574 -1214 34668
rect -1194 34574 -1190 34668
rect -1170 34574 -1166 34668
rect -1146 34574 -1142 34668
rect -1122 34643 -1118 34668
rect -1122 34595 -1115 34643
rect -1122 34574 -1118 34595
rect -1098 34574 -1094 34668
rect -1074 34574 -1070 34668
rect -1050 34574 -1046 34668
rect -1026 34574 -1022 34668
rect -1002 34574 -998 34668
rect -978 34574 -974 34668
rect -954 34574 -950 34668
rect -930 34574 -926 34668
rect -923 34667 -909 34668
rect -906 34667 -899 34691
rect -906 34574 -902 34667
rect -882 34574 -878 34716
rect -858 34574 -854 34716
rect -834 34574 -830 34716
rect -810 34574 -806 34716
rect -786 34574 -782 34716
rect -762 34574 -758 34716
rect -738 34574 -734 34716
rect -714 34574 -710 34716
rect -690 34574 -686 34716
rect -666 34574 -662 34716
rect -642 34574 -638 34716
rect -618 34574 -614 34716
rect -594 34574 -590 34716
rect -570 34574 -566 34716
rect -546 34574 -542 34716
rect -522 34574 -518 34716
rect -498 34574 -494 34716
rect -474 34574 -470 34716
rect -450 34574 -446 34716
rect -426 34574 -422 34716
rect -402 34574 -398 34716
rect -378 34574 -374 34716
rect -354 34574 -350 34716
rect -330 34574 -326 34716
rect -306 34574 -302 34716
rect -282 34574 -278 34716
rect -258 34574 -254 34716
rect -234 34574 -230 34716
rect -210 34574 -206 34716
rect -186 34574 -182 34716
rect -162 34574 -158 34716
rect -149 34637 -144 34647
rect -138 34637 -134 34716
rect -139 34623 -134 34637
rect -138 34574 -134 34623
rect -114 34574 -110 34716
rect -90 34574 -86 34716
rect -66 34574 -62 34716
rect -42 34574 -38 34716
rect -18 34574 -14 34716
rect 6 34574 10 34716
rect 30 34574 34 34716
rect 54 34574 58 34716
rect 78 34574 82 34716
rect 102 34574 106 34716
rect 126 34574 130 34716
rect 150 34574 154 34716
rect 174 34574 178 34716
rect 198 34574 202 34716
rect 222 34574 226 34716
rect 246 34574 250 34716
rect 270 34574 274 34716
rect 294 34574 298 34716
rect 318 34574 322 34716
rect 342 34574 346 34716
rect 366 34574 370 34716
rect 390 34574 394 34716
rect 414 34574 418 34716
rect 438 34574 442 34716
rect 462 34574 466 34716
rect 486 34574 490 34716
rect 510 34574 514 34716
rect 534 34574 538 34716
rect 547 34661 552 34671
rect 558 34661 562 34716
rect 557 34647 562 34661
rect 558 34574 562 34647
rect 582 34595 586 34716
rect -2393 34572 579 34574
rect -2371 34358 -2366 34572
rect -2348 34358 -2343 34572
rect -2325 34510 -2320 34572
rect -2317 34570 -2309 34572
rect -2000 34571 -1966 34572
rect -2000 34570 -1982 34571
rect -1663 34570 -1655 34572
rect -2028 34562 -2018 34564
rect -2309 34552 -2301 34558
rect -2091 34552 -2061 34559
rect -2317 34542 -2309 34552
rect -2044 34550 -2028 34552
rect -2026 34550 -2014 34562
rect -2084 34544 -2061 34550
rect -2044 34548 -2014 34550
rect -2292 34534 -2054 34543
rect -2325 34502 -2317 34510
rect -2325 34482 -2320 34502
rect -2317 34494 -2309 34502
rect -2325 34466 -2317 34482
rect -2325 34450 -2320 34466
rect -2309 34454 -2301 34466
rect -2317 34450 -2309 34454
rect -2103 34450 -2096 34452
rect -2083 34450 -2053 34452
rect -2325 34438 -2317 34450
rect -2103 34441 -2053 34450
rect -2018 34448 -2017 34454
rect -2003 34448 -2002 34450
rect -2026 34444 -2017 34448
rect -2325 34422 -2320 34438
rect -2309 34426 -2301 34438
rect -2017 34434 -2012 34444
rect -2317 34422 -2309 34426
rect -2325 34410 -2317 34422
rect -2325 34390 -2320 34410
rect -2325 34382 -2317 34390
rect -2325 34362 -2320 34382
rect -2317 34374 -2309 34382
rect -2325 34358 -2317 34362
rect -2000 34358 -1992 34570
rect -1982 34569 -1966 34570
rect -1980 34552 -1932 34559
rect -1655 34552 -1647 34558
rect -1846 34534 -1680 34543
rect -1663 34542 -1655 34552
rect -1671 34502 -1663 34510
rect -1663 34494 -1655 34502
rect -1671 34466 -1663 34482
rect -1655 34454 -1647 34466
rect -1972 34450 -1924 34452
rect -1663 34450 -1655 34454
rect -1972 34441 -1922 34450
rect -1671 34438 -1663 34450
rect -1655 34426 -1647 34438
rect -1663 34422 -1655 34426
rect -1671 34410 -1663 34422
rect -1671 34382 -1663 34390
rect -1663 34374 -1655 34382
rect -1671 34358 -1663 34362
rect -1642 34358 -1637 34572
rect -1619 34358 -1614 34572
rect -1530 34358 -1526 34572
rect -1506 34358 -1502 34572
rect -1482 34358 -1478 34572
rect -1458 34358 -1454 34572
rect -1434 34358 -1430 34572
rect -1410 34358 -1406 34572
rect -1386 34358 -1382 34572
rect -1362 34358 -1358 34572
rect -1338 34358 -1334 34572
rect -1314 34358 -1310 34572
rect -1290 34358 -1286 34572
rect -1266 34358 -1262 34572
rect -1242 34358 -1238 34572
rect -1218 34358 -1214 34572
rect -1194 34358 -1190 34572
rect -1170 34358 -1166 34572
rect -1146 34358 -1142 34572
rect -1122 34358 -1118 34572
rect -1098 34358 -1094 34572
rect -1074 34358 -1070 34572
rect -1050 34358 -1046 34572
rect -1026 34358 -1022 34572
rect -1002 34479 -998 34572
rect -1013 34478 -979 34479
rect -978 34478 -974 34572
rect -954 34478 -950 34572
rect -930 34478 -926 34572
rect -906 34478 -902 34572
rect -882 34478 -878 34572
rect -869 34517 -864 34527
rect -858 34517 -854 34572
rect -859 34503 -854 34517
rect -858 34478 -854 34503
rect -834 34478 -830 34572
rect -810 34478 -806 34572
rect -786 34478 -782 34572
rect -762 34478 -758 34572
rect -738 34478 -734 34572
rect -714 34478 -710 34572
rect -690 34478 -686 34572
rect -666 34478 -662 34572
rect -642 34478 -638 34572
rect -618 34478 -614 34572
rect -594 34478 -590 34572
rect -570 34478 -566 34572
rect -546 34478 -542 34572
rect -522 34478 -518 34572
rect -498 34478 -494 34572
rect -474 34478 -470 34572
rect -450 34478 -446 34572
rect -426 34478 -422 34572
rect -402 34478 -398 34572
rect -378 34478 -374 34572
rect -354 34478 -350 34572
rect -330 34478 -326 34572
rect -306 34478 -302 34572
rect -282 34478 -278 34572
rect -258 34478 -254 34572
rect -234 34478 -230 34572
rect -210 34478 -206 34572
rect -186 34478 -182 34572
rect -162 34478 -158 34572
rect -138 34478 -134 34572
rect -114 34571 -110 34572
rect -114 34547 -107 34571
rect -114 34478 -110 34547
rect -90 34478 -86 34572
rect -66 34478 -62 34572
rect -42 34478 -38 34572
rect -18 34478 -14 34572
rect 6 34478 10 34572
rect 30 34478 34 34572
rect 54 34478 58 34572
rect 78 34478 82 34572
rect 102 34478 106 34572
rect 126 34478 130 34572
rect 150 34478 154 34572
rect 174 34478 178 34572
rect 198 34478 202 34572
rect 222 34478 226 34572
rect 246 34478 250 34572
rect 270 34478 274 34572
rect 294 34478 298 34572
rect 318 34478 322 34572
rect 342 34478 346 34572
rect 366 34478 370 34572
rect 390 34478 394 34572
rect 414 34478 418 34572
rect 438 34478 442 34572
rect 462 34478 466 34572
rect 486 34478 490 34572
rect 510 34478 514 34572
rect 534 34478 538 34572
rect 558 34478 562 34572
rect 565 34571 579 34572
rect 582 34571 589 34595
rect 582 34478 586 34571
rect 606 34478 610 34716
rect 630 34478 634 34716
rect 654 34478 658 34716
rect 678 34478 682 34716
rect 702 34478 706 34716
rect 726 34478 730 34716
rect 750 34478 754 34716
rect 774 34478 778 34716
rect 798 34478 802 34716
rect 811 34589 816 34599
rect 822 34589 826 34716
rect 821 34575 826 34589
rect 811 34565 816 34575
rect 821 34551 826 34565
rect 822 34478 826 34551
rect 846 34523 850 34716
rect -1013 34476 843 34478
rect -1013 34469 -1008 34476
rect -1002 34469 -998 34476
rect -1003 34455 -998 34469
rect -1013 34445 -1008 34455
rect -1003 34431 -998 34445
rect -1002 34358 -998 34431
rect -978 34403 -974 34476
rect -2393 34356 -981 34358
rect -2371 34310 -2366 34356
rect -2348 34310 -2343 34356
rect -2325 34350 -2317 34356
rect -2018 34354 -2004 34356
rect -2325 34334 -2320 34350
rect -2317 34346 -2309 34350
rect -2069 34348 -2053 34350
rect -2309 34334 -2301 34346
rect -2096 34337 -2095 34343
rect -2000 34338 -1992 34356
rect -1671 34350 -1663 34356
rect -1663 34346 -1655 34350
rect -1977 34339 -1929 34345
rect -2112 34334 -2095 34337
rect -2325 34322 -2317 34334
rect -2325 34310 -2320 34322
rect -2317 34318 -2309 34322
rect -2112 34321 -2096 34334
rect -2059 34330 -2053 34337
rect -2027 34336 -1992 34338
rect -2059 34326 -2045 34330
rect -2018 34328 -2017 34330
rect -2083 34321 -2053 34322
rect -2019 34320 -2017 34324
rect -2309 34310 -2301 34318
rect -2017 34314 -2009 34320
rect -2000 34314 -1992 34336
rect -1972 34322 -1929 34337
rect -1655 34334 -1647 34346
rect -1671 34322 -1663 34334
rect -1972 34321 -1924 34322
rect -1663 34318 -1655 34322
rect -2033 34310 -1992 34314
rect -1655 34310 -1647 34318
rect -1642 34310 -1637 34356
rect -1619 34310 -1614 34356
rect -1530 34310 -1526 34356
rect -1506 34310 -1502 34356
rect -1482 34310 -1478 34356
rect -1458 34310 -1454 34356
rect -1434 34310 -1430 34356
rect -1410 34310 -1406 34356
rect -1386 34310 -1382 34356
rect -1362 34310 -1358 34356
rect -1338 34310 -1334 34356
rect -1314 34310 -1310 34356
rect -1290 34310 -1286 34356
rect -1266 34310 -1262 34356
rect -1242 34310 -1238 34356
rect -1218 34310 -1214 34356
rect -1194 34310 -1190 34356
rect -1170 34310 -1166 34356
rect -1146 34310 -1142 34356
rect -1122 34310 -1118 34356
rect -1098 34310 -1094 34356
rect -1074 34310 -1070 34356
rect -1050 34310 -1046 34356
rect -1026 34310 -1022 34356
rect -1002 34310 -998 34356
rect -995 34355 -981 34356
rect -978 34355 -971 34403
rect -978 34310 -974 34355
rect -954 34310 -950 34476
rect -930 34310 -926 34476
rect -906 34310 -902 34476
rect -882 34310 -878 34476
rect -858 34310 -854 34476
rect -834 34451 -830 34476
rect -834 34427 -827 34451
rect -834 34310 -830 34427
rect -810 34310 -806 34476
rect -786 34310 -782 34476
rect -762 34310 -758 34476
rect -738 34310 -734 34476
rect -714 34310 -710 34476
rect -690 34310 -686 34476
rect -666 34310 -662 34476
rect -642 34310 -638 34476
rect -618 34310 -614 34476
rect -594 34310 -590 34476
rect -570 34310 -566 34476
rect -546 34310 -542 34476
rect -522 34310 -518 34476
rect -498 34310 -494 34476
rect -474 34310 -470 34476
rect -450 34310 -446 34476
rect -426 34310 -422 34476
rect -402 34310 -398 34476
rect -378 34310 -374 34476
rect -354 34310 -350 34476
rect -330 34310 -326 34476
rect -306 34383 -302 34476
rect -293 34397 -288 34407
rect -282 34397 -278 34476
rect -283 34383 -278 34397
rect -317 34382 -283 34383
rect -282 34382 -278 34383
rect -258 34382 -254 34476
rect -234 34382 -230 34476
rect -210 34382 -206 34476
rect -186 34382 -182 34476
rect -162 34382 -158 34476
rect -138 34382 -134 34476
rect -114 34382 -110 34476
rect -90 34382 -86 34476
rect -66 34382 -62 34476
rect -42 34382 -38 34476
rect -18 34382 -14 34476
rect 6 34382 10 34476
rect 30 34382 34 34476
rect 54 34382 58 34476
rect 78 34382 82 34476
rect 102 34382 106 34476
rect 126 34382 130 34476
rect 150 34382 154 34476
rect 174 34382 178 34476
rect 198 34382 202 34476
rect 222 34382 226 34476
rect 246 34382 250 34476
rect 270 34382 274 34476
rect 294 34382 298 34476
rect 318 34382 322 34476
rect 342 34382 346 34476
rect 366 34382 370 34476
rect 390 34382 394 34476
rect 414 34382 418 34476
rect 438 34382 442 34476
rect 462 34382 466 34476
rect 486 34382 490 34476
rect 510 34382 514 34476
rect 534 34382 538 34476
rect 558 34382 562 34476
rect 582 34382 586 34476
rect 606 34382 610 34476
rect 630 34382 634 34476
rect 654 34382 658 34476
rect 678 34382 682 34476
rect 702 34382 706 34476
rect 726 34382 730 34476
rect 750 34382 754 34476
rect 774 34382 778 34476
rect 798 34382 802 34476
rect 822 34382 826 34476
rect 829 34475 843 34476
rect 846 34475 853 34523
rect 846 34382 850 34475
rect 870 34382 874 34716
rect 894 34382 898 34716
rect 918 34382 922 34716
rect 942 34382 946 34716
rect 966 34382 970 34716
rect 990 34382 994 34716
rect 1014 34382 1018 34716
rect 1038 34382 1042 34716
rect 1062 34382 1066 34716
rect 1086 34382 1090 34716
rect 1110 34382 1114 34716
rect 1134 34382 1138 34716
rect 1158 34382 1162 34716
rect 1182 34382 1186 34716
rect 1206 34382 1210 34716
rect 1230 34382 1234 34716
rect 1254 34382 1258 34716
rect 1278 34382 1282 34716
rect 1302 34382 1306 34716
rect 1326 34382 1330 34716
rect 1350 34382 1354 34716
rect 1374 34382 1378 34716
rect 1398 34382 1402 34716
rect 1422 34382 1426 34716
rect 1429 34715 1443 34716
rect 1435 34709 1440 34715
rect 1445 34695 1450 34709
rect 1446 34382 1450 34695
rect 1459 34589 1464 34599
rect 1469 34575 1474 34589
rect 1470 34382 1474 34575
rect 1483 34469 1488 34479
rect 1493 34455 1498 34469
rect 1494 34382 1498 34455
rect 1507 34382 1515 34383
rect -317 34380 1515 34382
rect -317 34373 -312 34380
rect -306 34373 -302 34380
rect -307 34359 -302 34373
rect -317 34349 -312 34359
rect -307 34335 -302 34349
rect -306 34310 -302 34335
rect -282 34310 -278 34380
rect -258 34331 -254 34380
rect -2393 34308 -261 34310
rect -2371 34214 -2366 34308
rect -2348 34214 -2343 34308
rect -2325 34306 -2320 34308
rect -2309 34306 -2301 34308
rect -2325 34294 -2317 34306
rect -2325 34274 -2320 34294
rect -2317 34290 -2309 34294
rect -2325 34266 -2317 34274
rect -2325 34214 -2320 34266
rect -2317 34258 -2309 34266
rect -2117 34257 -2095 34267
rect -2045 34264 -2037 34278
rect -2309 34218 -2301 34228
rect -2087 34224 -2076 34232
rect -2017 34228 -2015 34235
rect -2317 34214 -2309 34218
rect -2092 34216 -2087 34224
rect -2092 34214 -2077 34215
rect -2000 34214 -1992 34308
rect -1655 34306 -1647 34308
rect -1671 34294 -1663 34306
rect -1663 34290 -1655 34294
rect -1969 34257 -1929 34269
rect -1671 34266 -1663 34274
rect -1663 34258 -1655 34266
rect -1655 34218 -1647 34228
rect -1928 34214 -1924 34215
rect -1854 34214 -1680 34215
rect -1663 34214 -1655 34218
rect -1642 34214 -1637 34308
rect -1619 34214 -1614 34308
rect -1530 34214 -1526 34308
rect -1506 34214 -1502 34308
rect -1482 34214 -1478 34308
rect -1458 34214 -1454 34308
rect -1445 34277 -1440 34287
rect -1434 34277 -1430 34308
rect -1435 34263 -1430 34277
rect -1434 34214 -1430 34263
rect -1410 34214 -1406 34308
rect -1386 34214 -1382 34308
rect -1362 34214 -1358 34308
rect -1338 34214 -1334 34308
rect -1314 34214 -1310 34308
rect -1290 34214 -1286 34308
rect -1266 34214 -1262 34308
rect -1242 34214 -1238 34308
rect -1218 34214 -1214 34308
rect -1194 34214 -1190 34308
rect -1170 34214 -1166 34308
rect -1146 34214 -1142 34308
rect -1122 34214 -1118 34308
rect -1098 34214 -1094 34308
rect -1074 34214 -1070 34308
rect -1050 34214 -1046 34308
rect -1026 34214 -1022 34308
rect -1002 34214 -998 34308
rect -978 34214 -974 34308
rect -954 34214 -950 34308
rect -930 34214 -926 34308
rect -906 34214 -902 34308
rect -882 34214 -878 34308
rect -858 34214 -854 34308
rect -834 34214 -830 34308
rect -810 34214 -806 34308
rect -786 34214 -782 34308
rect -762 34214 -758 34308
rect -738 34214 -734 34308
rect -714 34214 -710 34308
rect -690 34214 -686 34308
rect -666 34214 -662 34308
rect -642 34214 -638 34308
rect -618 34214 -614 34308
rect -594 34214 -590 34308
rect -570 34214 -566 34308
rect -546 34214 -542 34308
rect -522 34214 -518 34308
rect -498 34214 -494 34308
rect -474 34214 -470 34308
rect -450 34214 -446 34308
rect -426 34214 -422 34308
rect -402 34214 -398 34308
rect -378 34214 -374 34308
rect -354 34214 -350 34308
rect -330 34214 -326 34308
rect -306 34214 -302 34308
rect -282 34307 -278 34308
rect -275 34307 -261 34308
rect -258 34307 -251 34331
rect -282 34259 -275 34307
rect -282 34214 -278 34259
rect -258 34214 -254 34307
rect -234 34214 -230 34380
rect -210 34214 -206 34380
rect -186 34214 -182 34380
rect -162 34214 -158 34380
rect -138 34214 -134 34380
rect -114 34214 -110 34380
rect -90 34214 -86 34380
rect -66 34214 -62 34380
rect -42 34214 -38 34380
rect -18 34214 -14 34380
rect 6 34214 10 34380
rect 30 34214 34 34380
rect 43 34253 48 34263
rect 54 34253 58 34380
rect 53 34239 58 34253
rect 43 34229 48 34239
rect 53 34215 58 34229
rect 54 34214 58 34215
rect 78 34214 82 34380
rect 102 34214 106 34380
rect 126 34214 130 34380
rect 150 34214 154 34380
rect 174 34214 178 34380
rect 198 34214 202 34380
rect 222 34214 226 34380
rect 246 34214 250 34380
rect 270 34214 274 34380
rect 294 34214 298 34380
rect 318 34214 322 34380
rect 342 34214 346 34380
rect 366 34214 370 34380
rect 390 34214 394 34380
rect 414 34214 418 34380
rect 438 34214 442 34380
rect 462 34214 466 34380
rect 486 34214 490 34380
rect 510 34214 514 34380
rect 534 34214 538 34380
rect 558 34214 562 34380
rect 582 34214 586 34380
rect 606 34214 610 34380
rect 630 34214 634 34380
rect 654 34214 658 34380
rect 678 34214 682 34380
rect 702 34214 706 34380
rect 726 34214 730 34380
rect 750 34214 754 34380
rect 774 34214 778 34380
rect 798 34214 802 34380
rect 822 34214 826 34380
rect 846 34214 850 34380
rect 870 34214 874 34380
rect 894 34214 898 34380
rect 918 34214 922 34380
rect 942 34214 946 34380
rect 966 34214 970 34380
rect 990 34214 994 34380
rect 1014 34214 1018 34380
rect 1038 34214 1042 34380
rect 1062 34214 1066 34380
rect 1086 34214 1090 34380
rect 1110 34214 1114 34380
rect 1134 34214 1138 34380
rect 1158 34214 1162 34380
rect 1182 34214 1186 34380
rect 1206 34214 1210 34380
rect 1219 34301 1224 34311
rect 1230 34301 1234 34380
rect 1229 34287 1234 34301
rect 1230 34215 1234 34287
rect 1254 34235 1258 34380
rect 1219 34214 1251 34215
rect -2393 34212 1251 34214
rect -2371 34190 -2366 34212
rect -2348 34190 -2343 34212
rect -2325 34190 -2320 34212
rect -2092 34207 -2037 34212
rect -2021 34207 -1969 34212
rect -1921 34207 -1913 34212
rect -1854 34208 -1680 34212
rect -2100 34205 -2092 34206
rect -2309 34190 -2301 34200
rect -2100 34199 -2087 34205
rect -2051 34192 -2026 34194
rect -2062 34190 -2012 34192
rect -2000 34190 -1992 34207
rect -1969 34199 -1921 34206
rect -1969 34190 -1964 34199
rect -1864 34190 -1796 34191
rect -1655 34190 -1647 34200
rect -1642 34190 -1637 34212
rect -1619 34190 -1614 34212
rect -1530 34190 -1526 34212
rect -1506 34190 -1502 34212
rect -1482 34190 -1478 34212
rect -1458 34190 -1454 34212
rect -1434 34190 -1430 34212
rect -1410 34211 -1406 34212
rect -2393 34188 -1413 34190
rect -2371 34142 -2366 34188
rect -2348 34142 -2343 34188
rect -2325 34142 -2320 34188
rect -2317 34184 -2309 34188
rect -2105 34181 -2092 34184
rect -2092 34158 -2062 34160
rect -2094 34154 -2062 34158
rect -2000 34142 -1992 34188
rect -1663 34184 -1655 34188
rect -1969 34181 -1921 34184
rect -1854 34158 -1806 34160
rect -1854 34154 -1680 34158
rect -1642 34142 -1637 34188
rect -1619 34142 -1614 34188
rect -1530 34142 -1526 34188
rect -1506 34142 -1502 34188
rect -1482 34142 -1478 34188
rect -1458 34142 -1454 34188
rect -1434 34142 -1430 34188
rect -1427 34187 -1413 34188
rect -1410 34187 -1403 34211
rect -1410 34142 -1406 34187
rect -1386 34142 -1382 34212
rect -1362 34142 -1358 34212
rect -1338 34142 -1334 34212
rect -1314 34142 -1310 34212
rect -1290 34142 -1286 34212
rect -1266 34142 -1262 34212
rect -1242 34142 -1238 34212
rect -1218 34142 -1214 34212
rect -1194 34142 -1190 34212
rect -1170 34142 -1166 34212
rect -1146 34142 -1142 34212
rect -1122 34142 -1118 34212
rect -1098 34142 -1094 34212
rect -1074 34142 -1070 34212
rect -1050 34142 -1046 34212
rect -1026 34142 -1022 34212
rect -1002 34142 -998 34212
rect -978 34142 -974 34212
rect -954 34142 -950 34212
rect -930 34142 -926 34212
rect -906 34142 -902 34212
rect -893 34157 -888 34167
rect -882 34157 -878 34212
rect -883 34143 -878 34157
rect -893 34142 -859 34143
rect -2393 34140 -859 34142
rect -2371 34118 -2366 34140
rect -2348 34118 -2343 34140
rect -2325 34118 -2320 34140
rect -2072 34138 -2036 34139
rect -2072 34132 -2054 34138
rect -2309 34124 -2301 34132
rect -2317 34118 -2309 34124
rect -2092 34123 -2062 34128
rect -2000 34119 -1992 34140
rect -1938 34139 -1906 34140
rect -1920 34138 -1906 34139
rect -1806 34132 -1680 34138
rect -1854 34123 -1806 34128
rect -1655 34124 -1647 34132
rect -1982 34119 -1966 34120
rect -2000 34118 -1966 34119
rect -1846 34118 -1806 34121
rect -1663 34118 -1655 34124
rect -1642 34118 -1637 34140
rect -1619 34118 -1614 34140
rect -1530 34118 -1526 34140
rect -1506 34118 -1502 34140
rect -1482 34118 -1478 34140
rect -1458 34118 -1454 34140
rect -1434 34118 -1430 34140
rect -1410 34118 -1406 34140
rect -1386 34118 -1382 34140
rect -1362 34118 -1358 34140
rect -1338 34118 -1334 34140
rect -1314 34118 -1310 34140
rect -1290 34118 -1286 34140
rect -1266 34118 -1262 34140
rect -1242 34118 -1238 34140
rect -1218 34118 -1214 34140
rect -1194 34118 -1190 34140
rect -1170 34118 -1166 34140
rect -1146 34118 -1142 34140
rect -1122 34118 -1118 34140
rect -1098 34118 -1094 34140
rect -1074 34118 -1070 34140
rect -1050 34118 -1046 34140
rect -1026 34118 -1022 34140
rect -1002 34118 -998 34140
rect -978 34118 -974 34140
rect -954 34118 -950 34140
rect -930 34118 -926 34140
rect -906 34118 -902 34140
rect -893 34133 -888 34140
rect -883 34119 -878 34133
rect -882 34118 -878 34119
rect -858 34118 -854 34212
rect -834 34118 -830 34212
rect -810 34118 -806 34212
rect -786 34118 -782 34212
rect -762 34118 -758 34212
rect -738 34118 -734 34212
rect -714 34118 -710 34212
rect -690 34118 -686 34212
rect -666 34118 -662 34212
rect -642 34118 -638 34212
rect -618 34118 -614 34212
rect -594 34118 -590 34212
rect -570 34119 -566 34212
rect -581 34118 -547 34119
rect -2393 34116 -547 34118
rect -2371 34094 -2366 34116
rect -2348 34094 -2343 34116
rect -2325 34094 -2320 34116
rect -2000 34114 -1966 34116
rect -2309 34096 -2301 34104
rect -2062 34103 -2054 34110
rect -2092 34096 -2084 34103
rect -2062 34096 -2026 34098
rect -2317 34094 -2309 34096
rect -2062 34094 -2012 34096
rect -2000 34094 -1992 34114
rect -1982 34113 -1966 34114
rect -1846 34112 -1806 34116
rect -1846 34105 -1798 34110
rect -1806 34103 -1798 34105
rect -1854 34101 -1846 34103
rect -1854 34096 -1806 34101
rect -1655 34096 -1647 34104
rect -1864 34094 -1796 34095
rect -1663 34094 -1655 34096
rect -1642 34094 -1637 34116
rect -1619 34094 -1614 34116
rect -1530 34094 -1526 34116
rect -1506 34094 -1502 34116
rect -1482 34094 -1478 34116
rect -1458 34094 -1454 34116
rect -1434 34094 -1430 34116
rect -1410 34094 -1406 34116
rect -1386 34094 -1382 34116
rect -1362 34094 -1358 34116
rect -1338 34094 -1334 34116
rect -1314 34094 -1310 34116
rect -1290 34094 -1286 34116
rect -1266 34094 -1262 34116
rect -1242 34094 -1238 34116
rect -1218 34094 -1214 34116
rect -1194 34094 -1190 34116
rect -1170 34094 -1166 34116
rect -1146 34094 -1142 34116
rect -1122 34094 -1118 34116
rect -1098 34094 -1094 34116
rect -1074 34094 -1070 34116
rect -1050 34094 -1046 34116
rect -1026 34094 -1022 34116
rect -1002 34094 -998 34116
rect -978 34094 -974 34116
rect -954 34094 -950 34116
rect -930 34094 -926 34116
rect -906 34094 -902 34116
rect -882 34094 -878 34116
rect -858 34094 -854 34116
rect -834 34094 -830 34116
rect -810 34094 -806 34116
rect -786 34094 -782 34116
rect -762 34094 -758 34116
rect -738 34094 -734 34116
rect -714 34094 -710 34116
rect -690 34094 -686 34116
rect -666 34094 -662 34116
rect -642 34094 -638 34116
rect -618 34094 -614 34116
rect -594 34094 -590 34116
rect -581 34109 -576 34116
rect -570 34109 -566 34116
rect -571 34095 -566 34109
rect -570 34094 -566 34095
rect -546 34094 -542 34212
rect -522 34094 -518 34212
rect -498 34094 -494 34212
rect -474 34094 -470 34212
rect -450 34094 -446 34212
rect -426 34094 -422 34212
rect -402 34094 -398 34212
rect -378 34094 -374 34212
rect -354 34094 -350 34212
rect -330 34094 -326 34212
rect -306 34094 -302 34212
rect -282 34094 -278 34212
rect -258 34094 -254 34212
rect -234 34094 -230 34212
rect -210 34094 -206 34212
rect -186 34094 -182 34212
rect -162 34094 -158 34212
rect -138 34095 -134 34212
rect -149 34094 -115 34095
rect -2393 34092 -115 34094
rect -2371 34046 -2366 34092
rect -2348 34046 -2343 34092
rect -2325 34046 -2320 34092
rect -2317 34088 -2309 34092
rect -2062 34088 -2054 34092
rect -2154 34084 -2138 34086
rect -2057 34084 -2054 34088
rect -2292 34078 -2054 34084
rect -2052 34078 -2044 34088
rect -2092 34062 -2062 34064
rect -2094 34058 -2062 34062
rect -2000 34046 -1992 34092
rect -1846 34085 -1806 34092
rect -1663 34088 -1655 34092
rect -1846 34078 -1680 34084
rect -1854 34062 -1806 34064
rect -1854 34058 -1680 34062
rect -1642 34046 -1637 34092
rect -1619 34046 -1614 34092
rect -1530 34046 -1526 34092
rect -1506 34046 -1502 34092
rect -1482 34046 -1478 34092
rect -1458 34046 -1454 34092
rect -1434 34046 -1430 34092
rect -1410 34046 -1406 34092
rect -1386 34046 -1382 34092
rect -1362 34046 -1358 34092
rect -1338 34046 -1334 34092
rect -1314 34046 -1310 34092
rect -1290 34046 -1286 34092
rect -1266 34046 -1262 34092
rect -1242 34046 -1238 34092
rect -1218 34046 -1214 34092
rect -1194 34046 -1190 34092
rect -1170 34046 -1166 34092
rect -1146 34046 -1142 34092
rect -1122 34046 -1118 34092
rect -1098 34046 -1094 34092
rect -1074 34046 -1070 34092
rect -1050 34046 -1046 34092
rect -1026 34046 -1022 34092
rect -1002 34046 -998 34092
rect -978 34046 -974 34092
rect -954 34046 -950 34092
rect -930 34046 -926 34092
rect -906 34046 -902 34092
rect -882 34046 -878 34092
rect -858 34091 -854 34092
rect -2393 34044 -861 34046
rect -2371 34022 -2366 34044
rect -2348 34022 -2343 34044
rect -2325 34022 -2320 34044
rect -2072 34042 -2036 34043
rect -2072 34036 -2054 34042
rect -2309 34028 -2301 34036
rect -2317 34022 -2309 34028
rect -2092 34027 -2062 34032
rect -2000 34023 -1992 34044
rect -1938 34043 -1906 34044
rect -1920 34042 -1906 34043
rect -1806 34036 -1680 34042
rect -1854 34027 -1806 34032
rect -1655 34028 -1647 34036
rect -1982 34023 -1966 34024
rect -2000 34022 -1966 34023
rect -1846 34022 -1806 34025
rect -1663 34022 -1655 34028
rect -1642 34022 -1637 34044
rect -1619 34022 -1614 34044
rect -1530 34022 -1526 34044
rect -1506 34022 -1502 34044
rect -1482 34022 -1478 34044
rect -1458 34022 -1454 34044
rect -1434 34023 -1430 34044
rect -1445 34022 -1411 34023
rect -2393 34020 -1411 34022
rect -2371 33998 -2366 34020
rect -2348 33998 -2343 34020
rect -2325 33998 -2320 34020
rect -2000 34018 -1966 34020
rect -2309 34000 -2301 34008
rect -2062 34007 -2054 34014
rect -2092 34000 -2084 34007
rect -2062 34000 -2026 34002
rect -2317 33998 -2309 34000
rect -2062 33998 -2012 34000
rect -2000 33998 -1992 34018
rect -1982 34017 -1966 34018
rect -1846 34016 -1806 34020
rect -1846 34009 -1798 34014
rect -1806 34007 -1798 34009
rect -1854 34005 -1846 34007
rect -1854 34000 -1806 34005
rect -1655 34000 -1647 34008
rect -1864 33998 -1796 33999
rect -1663 33998 -1655 34000
rect -1642 33998 -1637 34020
rect -1619 33998 -1614 34020
rect -1530 33998 -1526 34020
rect -1506 33998 -1502 34020
rect -1482 33998 -1478 34020
rect -1458 33998 -1454 34020
rect -1445 34013 -1440 34020
rect -1434 34013 -1430 34020
rect -1435 33999 -1430 34013
rect -1434 33998 -1430 33999
rect -1410 33998 -1406 34044
rect -1386 33998 -1382 34044
rect -1362 33998 -1358 34044
rect -1338 33998 -1334 34044
rect -1314 33998 -1310 34044
rect -1290 33998 -1286 34044
rect -1266 33998 -1262 34044
rect -1242 33998 -1238 34044
rect -1218 33998 -1214 34044
rect -1194 33998 -1190 34044
rect -1170 33998 -1166 34044
rect -1146 33998 -1142 34044
rect -1122 33998 -1118 34044
rect -1098 33998 -1094 34044
rect -1074 33998 -1070 34044
rect -1050 33998 -1046 34044
rect -1026 33998 -1022 34044
rect -1002 33998 -998 34044
rect -978 33998 -974 34044
rect -954 33998 -950 34044
rect -930 33998 -926 34044
rect -906 33998 -902 34044
rect -882 33998 -878 34044
rect -875 34043 -861 34044
rect -858 34043 -851 34091
rect -858 33998 -854 34043
rect -834 33998 -830 34092
rect -810 33998 -806 34092
rect -786 33998 -782 34092
rect -762 33998 -758 34092
rect -738 33998 -734 34092
rect -714 33998 -710 34092
rect -690 33998 -686 34092
rect -666 33998 -662 34092
rect -642 33998 -638 34092
rect -618 33998 -614 34092
rect -594 33998 -590 34092
rect -570 33998 -566 34092
rect -546 34043 -542 34092
rect -546 34019 -539 34043
rect -546 33998 -542 34019
rect -522 33998 -518 34092
rect -498 33998 -494 34092
rect -474 33998 -470 34092
rect -450 33998 -446 34092
rect -426 33998 -422 34092
rect -402 33998 -398 34092
rect -378 33998 -374 34092
rect -354 33998 -350 34092
rect -330 33998 -326 34092
rect -306 33998 -302 34092
rect -282 33998 -278 34092
rect -258 33998 -254 34092
rect -234 33998 -230 34092
rect -210 33998 -206 34092
rect -186 33998 -182 34092
rect -162 33999 -158 34092
rect -149 34085 -144 34092
rect -138 34085 -134 34092
rect -139 34071 -134 34085
rect -173 33998 -139 33999
rect -2393 33996 -139 33998
rect -2371 33950 -2366 33996
rect -2348 33950 -2343 33996
rect -2325 33950 -2320 33996
rect -2317 33992 -2309 33996
rect -2062 33992 -2054 33996
rect -2154 33988 -2138 33990
rect -2057 33988 -2054 33992
rect -2292 33982 -2054 33988
rect -2052 33982 -2044 33992
rect -2092 33966 -2062 33968
rect -2094 33962 -2062 33966
rect -2000 33950 -1992 33996
rect -1846 33989 -1806 33996
rect -1663 33992 -1655 33996
rect -1846 33982 -1680 33988
rect -1854 33966 -1806 33968
rect -1854 33962 -1680 33966
rect -1642 33950 -1637 33996
rect -1619 33950 -1614 33996
rect -1530 33950 -1526 33996
rect -1506 33950 -1502 33996
rect -1482 33950 -1478 33996
rect -1458 33950 -1454 33996
rect -1434 33950 -1430 33996
rect -1410 33950 -1406 33996
rect -1386 33950 -1382 33996
rect -1362 33950 -1358 33996
rect -1338 33950 -1334 33996
rect -1314 33950 -1310 33996
rect -1290 33950 -1286 33996
rect -1266 33950 -1262 33996
rect -1242 33950 -1238 33996
rect -1218 33950 -1214 33996
rect -1205 33965 -1200 33975
rect -1194 33965 -1190 33996
rect -1195 33951 -1190 33965
rect -1205 33950 -1171 33951
rect -2393 33948 -1171 33950
rect -2371 33902 -2366 33948
rect -2348 33902 -2343 33948
rect -2325 33902 -2320 33948
rect -2309 33932 -2301 33942
rect -2317 33926 -2309 33932
rect -2097 33926 -2095 33935
rect -2309 33904 -2301 33914
rect -2097 33912 -2095 33916
rect -2292 33911 -2095 33912
rect -2097 33909 -2095 33911
rect -2084 33904 -2083 33947
rect -2069 33940 -2054 33942
rect -2054 33924 -2018 33926
rect -2054 33922 -2004 33924
rect -2059 33918 -2045 33922
rect -2054 33916 -2049 33918
rect -2317 33902 -2309 33904
rect -2084 33902 -2054 33904
rect -2044 33902 -2039 33916
rect -2025 33906 -2014 33912
rect -2000 33906 -1992 33948
rect -1920 33946 -1906 33948
rect -1977 33931 -1929 33937
rect -1655 33932 -1647 33942
rect -1977 33921 -1966 33931
rect -1663 33926 -1655 33932
rect -1977 33909 -1929 33911
rect -2033 33902 -1992 33906
rect -1655 33904 -1647 33914
rect -1663 33902 -1655 33904
rect -1642 33902 -1637 33948
rect -1619 33902 -1614 33948
rect -1530 33902 -1526 33948
rect -1506 33902 -1502 33948
rect -1482 33902 -1478 33948
rect -1458 33902 -1454 33948
rect -1434 33902 -1430 33948
rect -1410 33947 -1406 33948
rect -1410 33923 -1403 33947
rect -1410 33902 -1406 33923
rect -1386 33902 -1382 33948
rect -1362 33902 -1358 33948
rect -1338 33902 -1334 33948
rect -1314 33902 -1310 33948
rect -1290 33902 -1286 33948
rect -1266 33902 -1262 33948
rect -1242 33902 -1238 33948
rect -1218 33902 -1214 33948
rect -1205 33941 -1200 33948
rect -1195 33927 -1190 33941
rect -1194 33902 -1190 33927
rect -1170 33902 -1166 33996
rect -1146 33902 -1142 33996
rect -1122 33902 -1118 33996
rect -1098 33902 -1094 33996
rect -1074 33902 -1070 33996
rect -1050 33902 -1046 33996
rect -1026 33902 -1022 33996
rect -1002 33902 -998 33996
rect -978 33902 -974 33996
rect -954 33902 -950 33996
rect -930 33902 -926 33996
rect -906 33902 -902 33996
rect -882 33902 -878 33996
rect -858 33902 -854 33996
rect -834 33902 -830 33996
rect -810 33902 -806 33996
rect -786 33902 -782 33996
rect -762 33902 -758 33996
rect -738 33902 -734 33996
rect -714 33902 -710 33996
rect -690 33902 -686 33996
rect -666 33902 -662 33996
rect -642 33902 -638 33996
rect -618 33902 -614 33996
rect -594 33902 -590 33996
rect -570 33902 -566 33996
rect -546 33902 -542 33996
rect -522 33902 -518 33996
rect -498 33902 -494 33996
rect -474 33902 -470 33996
rect -450 33902 -446 33996
rect -426 33902 -422 33996
rect -402 33902 -398 33996
rect -378 33902 -374 33996
rect -354 33902 -350 33996
rect -330 33902 -326 33996
rect -306 33902 -302 33996
rect -282 33902 -278 33996
rect -258 33902 -254 33996
rect -234 33902 -230 33996
rect -210 33902 -206 33996
rect -186 33902 -182 33996
rect -173 33989 -168 33996
rect -162 33989 -158 33996
rect -163 33975 -158 33989
rect -162 33902 -158 33975
rect -138 33923 -134 34071
rect -114 34019 -110 34212
rect -114 33995 -107 34019
rect -2393 33900 -141 33902
rect -2371 33806 -2366 33900
rect -2348 33806 -2343 33900
rect -2325 33866 -2320 33900
rect -2317 33898 -2309 33900
rect -2084 33887 -2083 33900
rect -2084 33886 -2054 33887
rect -2325 33858 -2317 33866
rect -2325 33806 -2320 33858
rect -2317 33850 -2309 33858
rect -2117 33849 -2095 33859
rect -2045 33856 -2037 33870
rect -2309 33810 -2301 33818
rect -2317 33806 -2309 33810
rect -2000 33806 -1992 33900
rect -1663 33898 -1655 33900
rect -1969 33849 -1929 33861
rect -1671 33858 -1663 33866
rect -1663 33850 -1655 33858
rect -1655 33810 -1647 33818
rect -1663 33806 -1655 33810
rect -1642 33806 -1637 33900
rect -1619 33806 -1614 33900
rect -1530 33806 -1526 33900
rect -1506 33806 -1502 33900
rect -1482 33806 -1478 33900
rect -1458 33806 -1454 33900
rect -1434 33806 -1430 33900
rect -1410 33806 -1406 33900
rect -1386 33806 -1382 33900
rect -1362 33806 -1358 33900
rect -1338 33806 -1334 33900
rect -1314 33806 -1310 33900
rect -1290 33806 -1286 33900
rect -1266 33806 -1262 33900
rect -1242 33806 -1238 33900
rect -1218 33806 -1214 33900
rect -1194 33806 -1190 33900
rect -1170 33899 -1166 33900
rect -1170 33878 -1163 33899
rect -1146 33878 -1142 33900
rect -1122 33878 -1118 33900
rect -1098 33878 -1094 33900
rect -1074 33878 -1070 33900
rect -1050 33878 -1046 33900
rect -1026 33878 -1022 33900
rect -1002 33878 -998 33900
rect -978 33878 -974 33900
rect -954 33878 -950 33900
rect -930 33878 -926 33900
rect -906 33878 -902 33900
rect -882 33878 -878 33900
rect -858 33878 -854 33900
rect -834 33878 -830 33900
rect -810 33878 -806 33900
rect -786 33878 -782 33900
rect -762 33878 -758 33900
rect -738 33878 -734 33900
rect -714 33878 -710 33900
rect -690 33878 -686 33900
rect -666 33878 -662 33900
rect -642 33878 -638 33900
rect -618 33878 -614 33900
rect -594 33878 -590 33900
rect -570 33878 -566 33900
rect -546 33878 -542 33900
rect -522 33878 -518 33900
rect -498 33878 -494 33900
rect -474 33878 -470 33900
rect -450 33878 -446 33900
rect -426 33878 -422 33900
rect -402 33878 -398 33900
rect -378 33878 -374 33900
rect -354 33878 -350 33900
rect -330 33878 -326 33900
rect -306 33878 -302 33900
rect -282 33878 -278 33900
rect -258 33878 -254 33900
rect -234 33878 -230 33900
rect -210 33878 -206 33900
rect -186 33878 -182 33900
rect -162 33878 -158 33900
rect -155 33899 -141 33900
rect -138 33899 -131 33923
rect -138 33878 -134 33899
rect -114 33878 -110 33995
rect -90 33878 -86 34212
rect -66 33878 -62 34212
rect -42 33878 -38 34212
rect -18 33878 -14 34212
rect 6 33878 10 34212
rect 30 33878 34 34212
rect 54 33878 58 34212
rect 78 34187 82 34212
rect 78 34166 85 34187
rect 102 34166 106 34212
rect 126 34166 130 34212
rect 150 34166 154 34212
rect 174 34166 178 34212
rect 198 34166 202 34212
rect 222 34166 226 34212
rect 246 34166 250 34212
rect 270 34166 274 34212
rect 283 34181 288 34191
rect 294 34181 298 34212
rect 293 34167 298 34181
rect 294 34166 298 34167
rect 318 34166 322 34212
rect 342 34166 346 34212
rect 366 34166 370 34212
rect 390 34166 394 34212
rect 414 34166 418 34212
rect 438 34166 442 34212
rect 462 34166 466 34212
rect 486 34166 490 34212
rect 510 34166 514 34212
rect 534 34166 538 34212
rect 558 34166 562 34212
rect 582 34166 586 34212
rect 606 34166 610 34212
rect 630 34166 634 34212
rect 654 34166 658 34212
rect 678 34166 682 34212
rect 702 34166 706 34212
rect 726 34166 730 34212
rect 750 34166 754 34212
rect 774 34166 778 34212
rect 798 34166 802 34212
rect 822 34166 826 34212
rect 846 34166 850 34212
rect 870 34166 874 34212
rect 894 34166 898 34212
rect 918 34166 922 34212
rect 942 34166 946 34212
rect 966 34166 970 34212
rect 990 34166 994 34212
rect 1014 34166 1018 34212
rect 1038 34166 1042 34212
rect 1062 34166 1066 34212
rect 1086 34166 1090 34212
rect 1110 34166 1114 34212
rect 1134 34166 1138 34212
rect 1158 34166 1162 34212
rect 1182 34166 1186 34212
rect 1206 34166 1210 34212
rect 1219 34205 1224 34212
rect 1230 34205 1234 34212
rect 1237 34211 1251 34212
rect 1254 34211 1261 34235
rect 1229 34191 1234 34205
rect 1230 34166 1234 34191
rect 1254 34166 1258 34211
rect 1278 34166 1282 34380
rect 1302 34166 1306 34380
rect 1326 34166 1330 34380
rect 1350 34166 1354 34380
rect 1374 34166 1378 34380
rect 1398 34166 1402 34380
rect 1422 34166 1426 34380
rect 1446 34166 1450 34380
rect 1470 34166 1474 34380
rect 1494 34166 1498 34380
rect 1501 34379 1515 34380
rect 1507 34373 1512 34379
rect 1517 34359 1522 34373
rect 1518 34166 1522 34359
rect 1531 34253 1536 34263
rect 1541 34239 1546 34253
rect 1542 34166 1546 34239
rect 1555 34166 1563 34167
rect 61 34164 1563 34166
rect 61 34163 75 34164
rect 78 34139 85 34164
rect 78 33878 82 34139
rect 102 33878 106 34164
rect 126 33878 130 34164
rect 150 33878 154 34164
rect 174 33878 178 34164
rect 198 33878 202 34164
rect 222 34071 226 34164
rect 211 34070 245 34071
rect 246 34070 250 34164
rect 270 34070 274 34164
rect 294 34070 298 34164
rect 318 34115 322 34164
rect 318 34091 325 34115
rect 318 34070 322 34091
rect 342 34070 346 34164
rect 366 34070 370 34164
rect 390 34070 394 34164
rect 414 34070 418 34164
rect 438 34070 442 34164
rect 462 34070 466 34164
rect 486 34070 490 34164
rect 510 34070 514 34164
rect 534 34070 538 34164
rect 558 34070 562 34164
rect 582 34070 586 34164
rect 606 34070 610 34164
rect 630 34070 634 34164
rect 654 34070 658 34164
rect 678 34070 682 34164
rect 702 34070 706 34164
rect 726 34070 730 34164
rect 750 34070 754 34164
rect 774 34070 778 34164
rect 798 34070 802 34164
rect 822 34070 826 34164
rect 846 34070 850 34164
rect 870 34070 874 34164
rect 894 34070 898 34164
rect 918 34070 922 34164
rect 942 34070 946 34164
rect 966 34070 970 34164
rect 990 34070 994 34164
rect 1014 34070 1018 34164
rect 1038 34070 1042 34164
rect 1062 34070 1066 34164
rect 1086 34070 1090 34164
rect 1110 34070 1114 34164
rect 1134 34070 1138 34164
rect 1158 34070 1162 34164
rect 1182 34070 1186 34164
rect 1206 34070 1210 34164
rect 1230 34070 1234 34164
rect 1254 34139 1258 34164
rect 1254 34115 1261 34139
rect 1254 34070 1258 34115
rect 1278 34070 1282 34164
rect 1302 34070 1306 34164
rect 1326 34070 1330 34164
rect 1350 34070 1354 34164
rect 1374 34070 1378 34164
rect 1398 34070 1402 34164
rect 1422 34070 1426 34164
rect 1446 34070 1450 34164
rect 1470 34070 1474 34164
rect 1494 34070 1498 34164
rect 1518 34070 1522 34164
rect 1542 34070 1546 34164
rect 1549 34163 1563 34164
rect 1555 34157 1560 34163
rect 1565 34143 1570 34157
rect 1566 34070 1570 34143
rect 1579 34070 1587 34071
rect 211 34068 1587 34070
rect 211 34061 216 34068
rect 222 34061 226 34068
rect 221 34047 226 34061
rect 211 34037 216 34047
rect 221 34023 226 34037
rect 222 33878 226 34023
rect 246 33995 250 34068
rect 246 33974 253 33995
rect 270 33974 274 34068
rect 294 33974 298 34068
rect 318 33974 322 34068
rect 342 33974 346 34068
rect 366 33974 370 34068
rect 390 33974 394 34068
rect 414 33974 418 34068
rect 438 33974 442 34068
rect 462 33974 466 34068
rect 486 33974 490 34068
rect 510 33974 514 34068
rect 534 33974 538 34068
rect 558 33974 562 34068
rect 582 33974 586 34068
rect 606 33974 610 34068
rect 630 33974 634 34068
rect 654 33974 658 34068
rect 678 33974 682 34068
rect 702 33974 706 34068
rect 726 33974 730 34068
rect 750 33974 754 34068
rect 774 33974 778 34068
rect 798 33974 802 34068
rect 822 33974 826 34068
rect 846 33974 850 34068
rect 870 33974 874 34068
rect 894 33974 898 34068
rect 918 33974 922 34068
rect 942 33974 946 34068
rect 966 33974 970 34068
rect 990 33974 994 34068
rect 1014 33974 1018 34068
rect 1038 33974 1042 34068
rect 1062 33974 1066 34068
rect 1086 33974 1090 34068
rect 1110 33974 1114 34068
rect 1134 33974 1138 34068
rect 1158 33974 1162 34068
rect 1182 33974 1186 34068
rect 1206 33974 1210 34068
rect 1230 33974 1234 34068
rect 1254 33974 1258 34068
rect 1278 33974 1282 34068
rect 1302 33974 1306 34068
rect 1326 33974 1330 34068
rect 1350 33974 1354 34068
rect 1374 33974 1378 34068
rect 1398 33974 1402 34068
rect 1422 33974 1426 34068
rect 1446 33974 1450 34068
rect 1470 33974 1474 34068
rect 1494 33974 1498 34068
rect 1518 33974 1522 34068
rect 1542 33974 1546 34068
rect 1566 33974 1570 34068
rect 1573 34067 1587 34068
rect 1579 34061 1584 34067
rect 1589 34047 1594 34061
rect 1590 33974 1594 34047
rect 1603 33974 1611 33975
rect 229 33972 1611 33974
rect 229 33971 243 33972
rect 246 33947 253 33972
rect 246 33878 250 33947
rect 270 33878 274 33972
rect 294 33878 298 33972
rect 318 33878 322 33972
rect 342 33878 346 33972
rect 366 33878 370 33972
rect 390 33878 394 33972
rect 414 33878 418 33972
rect 438 33878 442 33972
rect 462 33878 466 33972
rect 486 33878 490 33972
rect 510 33878 514 33972
rect 534 33878 538 33972
rect 558 33878 562 33972
rect 582 33878 586 33972
rect 606 33878 610 33972
rect 630 33878 634 33972
rect 654 33878 658 33972
rect 678 33878 682 33972
rect 702 33878 706 33972
rect 726 33878 730 33972
rect 750 33878 754 33972
rect 774 33878 778 33972
rect 798 33878 802 33972
rect 822 33878 826 33972
rect 846 33878 850 33972
rect 870 33878 874 33972
rect 894 33878 898 33972
rect 918 33878 922 33972
rect 942 33878 946 33972
rect 966 33878 970 33972
rect 990 33878 994 33972
rect 1014 33878 1018 33972
rect 1038 33878 1042 33972
rect 1062 33878 1066 33972
rect 1086 33878 1090 33972
rect 1110 33878 1114 33972
rect 1134 33878 1138 33972
rect 1158 33878 1162 33972
rect 1182 33878 1186 33972
rect 1206 33878 1210 33972
rect 1230 33879 1234 33972
rect 1219 33878 1253 33879
rect -1187 33876 1253 33878
rect -1187 33875 -1173 33876
rect -1170 33851 -1163 33876
rect -1170 33806 -1166 33851
rect -1146 33806 -1142 33876
rect -1122 33806 -1118 33876
rect -1098 33806 -1094 33876
rect -1074 33806 -1070 33876
rect -1050 33806 -1046 33876
rect -1026 33806 -1022 33876
rect -1002 33806 -998 33876
rect -978 33806 -974 33876
rect -954 33806 -950 33876
rect -930 33806 -926 33876
rect -906 33806 -902 33876
rect -882 33806 -878 33876
rect -858 33806 -854 33876
rect -834 33806 -830 33876
rect -810 33806 -806 33876
rect -786 33806 -782 33876
rect -762 33806 -758 33876
rect -738 33806 -734 33876
rect -714 33806 -710 33876
rect -690 33806 -686 33876
rect -666 33806 -662 33876
rect -642 33806 -638 33876
rect -618 33806 -614 33876
rect -594 33806 -590 33876
rect -570 33806 -566 33876
rect -546 33806 -542 33876
rect -522 33806 -518 33876
rect -498 33806 -494 33876
rect -474 33806 -470 33876
rect -450 33806 -446 33876
rect -426 33806 -422 33876
rect -402 33806 -398 33876
rect -378 33806 -374 33876
rect -354 33806 -350 33876
rect -330 33806 -326 33876
rect -306 33806 -302 33876
rect -282 33806 -278 33876
rect -258 33806 -254 33876
rect -234 33806 -230 33876
rect -210 33806 -206 33876
rect -186 33806 -182 33876
rect -162 33806 -158 33876
rect -138 33806 -134 33876
rect -114 33806 -110 33876
rect -90 33806 -86 33876
rect -66 33806 -62 33876
rect -42 33806 -38 33876
rect -18 33806 -14 33876
rect 6 33806 10 33876
rect 30 33806 34 33876
rect 54 33806 58 33876
rect 78 33806 82 33876
rect 102 33806 106 33876
rect 126 33806 130 33876
rect 150 33806 154 33876
rect 174 33806 178 33876
rect 198 33806 202 33876
rect 222 33806 226 33876
rect 246 33806 250 33876
rect 270 33806 274 33876
rect 294 33806 298 33876
rect 318 33806 322 33876
rect 342 33806 346 33876
rect 366 33806 370 33876
rect 390 33806 394 33876
rect 414 33806 418 33876
rect 438 33806 442 33876
rect 462 33806 466 33876
rect 486 33806 490 33876
rect 510 33806 514 33876
rect 534 33806 538 33876
rect 558 33806 562 33876
rect 582 33806 586 33876
rect 606 33806 610 33876
rect 630 33806 634 33876
rect 654 33806 658 33876
rect 678 33806 682 33876
rect 702 33806 706 33876
rect 726 33806 730 33876
rect 750 33806 754 33876
rect 763 33821 768 33831
rect 774 33821 778 33876
rect 773 33807 778 33821
rect 763 33806 797 33807
rect -2393 33804 -2026 33806
rect -2021 33804 797 33806
rect -2371 33710 -2366 33804
rect -2348 33710 -2343 33804
rect -2325 33742 -2320 33804
rect -2317 33802 -2309 33804
rect -2309 33782 -2301 33790
rect -2317 33774 -2309 33782
rect -2123 33777 -2116 33782
rect -2123 33775 -2092 33777
rect -2091 33776 -2087 33792
rect -2026 33784 -2021 33796
rect -2037 33780 -2021 33784
rect -2292 33773 -2087 33775
rect -2123 33771 -2116 33773
rect -2325 33734 -2317 33742
rect -2325 33714 -2320 33734
rect -2317 33726 -2309 33734
rect -2325 33710 -2317 33714
rect -2000 33710 -1992 33804
rect -1663 33802 -1655 33804
rect -1969 33776 -1932 33792
rect -1655 33782 -1647 33790
rect -1969 33773 -1680 33775
rect -1663 33774 -1655 33782
rect -1671 33734 -1663 33742
rect -1663 33726 -1655 33734
rect -1671 33710 -1663 33714
rect -1642 33710 -1637 33804
rect -1619 33710 -1614 33804
rect -1530 33710 -1526 33804
rect -1506 33710 -1502 33804
rect -1482 33710 -1478 33804
rect -1458 33710 -1454 33804
rect -1434 33710 -1430 33804
rect -1410 33710 -1406 33804
rect -1386 33710 -1382 33804
rect -1362 33710 -1358 33804
rect -1338 33710 -1334 33804
rect -1314 33710 -1310 33804
rect -1290 33710 -1286 33804
rect -1266 33710 -1262 33804
rect -1242 33710 -1238 33804
rect -1218 33710 -1214 33804
rect -1194 33710 -1190 33804
rect -1170 33710 -1166 33804
rect -1146 33710 -1142 33804
rect -1122 33710 -1118 33804
rect -1098 33710 -1094 33804
rect -1074 33710 -1070 33804
rect -1050 33710 -1046 33804
rect -1026 33710 -1022 33804
rect -1002 33710 -998 33804
rect -978 33710 -974 33804
rect -954 33710 -950 33804
rect -930 33710 -926 33804
rect -906 33710 -902 33804
rect -882 33710 -878 33804
rect -858 33710 -854 33804
rect -834 33710 -830 33804
rect -810 33710 -806 33804
rect -786 33710 -782 33804
rect -762 33710 -758 33804
rect -738 33710 -734 33804
rect -714 33710 -710 33804
rect -690 33710 -686 33804
rect -666 33710 -662 33804
rect -642 33710 -638 33804
rect -618 33710 -614 33804
rect -594 33710 -590 33804
rect -570 33710 -566 33804
rect -546 33710 -542 33804
rect -522 33710 -518 33804
rect -498 33710 -494 33804
rect -474 33710 -470 33804
rect -450 33710 -446 33804
rect -426 33710 -422 33804
rect -402 33710 -398 33804
rect -378 33710 -374 33804
rect -354 33710 -350 33804
rect -330 33710 -326 33804
rect -306 33710 -302 33804
rect -282 33710 -278 33804
rect -258 33710 -254 33804
rect -234 33710 -230 33804
rect -210 33710 -206 33804
rect -186 33710 -182 33804
rect -162 33710 -158 33804
rect -138 33710 -134 33804
rect -114 33710 -110 33804
rect -90 33710 -86 33804
rect -66 33710 -62 33804
rect -42 33710 -38 33804
rect -18 33710 -14 33804
rect 6 33710 10 33804
rect 30 33710 34 33804
rect 54 33710 58 33804
rect 78 33710 82 33804
rect 102 33710 106 33804
rect 126 33710 130 33804
rect 150 33710 154 33804
rect 174 33710 178 33804
rect 198 33710 202 33804
rect 222 33710 226 33804
rect 246 33710 250 33804
rect 270 33710 274 33804
rect 294 33710 298 33804
rect 318 33710 322 33804
rect 342 33710 346 33804
rect 366 33710 370 33804
rect 390 33710 394 33804
rect 414 33710 418 33804
rect 438 33710 442 33804
rect 462 33710 466 33804
rect 486 33710 490 33804
rect 510 33710 514 33804
rect 534 33710 538 33804
rect 558 33710 562 33804
rect 582 33710 586 33804
rect 606 33710 610 33804
rect 630 33710 634 33804
rect 654 33710 658 33804
rect 678 33710 682 33804
rect 702 33710 706 33804
rect 726 33710 730 33804
rect 750 33710 754 33804
rect 763 33797 768 33804
rect 773 33783 778 33797
rect 774 33710 778 33783
rect 798 33755 802 33876
rect -2393 33708 795 33710
rect -2371 33662 -2366 33708
rect -2348 33662 -2343 33708
rect -2325 33700 -2317 33708
rect -2018 33707 -2004 33708
rect -2000 33707 -1992 33708
rect -2072 33706 -1928 33707
rect -2072 33700 -2053 33706
rect -2325 33684 -2320 33700
rect -2317 33698 -2309 33700
rect -2309 33686 -2301 33698
rect -2092 33691 -2062 33696
rect -2317 33684 -2309 33686
rect -2325 33672 -2317 33684
rect -2098 33678 -2096 33689
rect -2092 33678 -2084 33691
rect -2000 33690 -1992 33706
rect -1972 33700 -1928 33706
rect -1924 33700 -1918 33708
rect -1671 33700 -1663 33708
rect -1663 33698 -1655 33700
rect -2083 33680 -2062 33689
rect -2027 33688 -1992 33690
rect -2018 33680 -2002 33688
rect -2000 33680 -1992 33688
rect -2100 33673 -2096 33678
rect -2083 33673 -2053 33678
rect -2003 33676 -1990 33680
rect -1972 33678 -1964 33687
rect -1928 33686 -1924 33689
rect -1655 33686 -1647 33698
rect -1663 33684 -1655 33686
rect -2325 33662 -2320 33672
rect -2317 33670 -2309 33672
rect -2309 33662 -2301 33670
rect -2004 33666 -2003 33676
rect -2062 33662 -2012 33664
rect -2000 33662 -1992 33676
rect -1972 33673 -1924 33678
rect -1864 33673 -1796 33679
rect -1671 33672 -1663 33684
rect -1663 33670 -1655 33672
rect -1864 33662 -1796 33663
rect -1655 33662 -1647 33670
rect -1642 33662 -1637 33708
rect -1619 33662 -1614 33708
rect -1530 33662 -1526 33708
rect -1506 33662 -1502 33708
rect -1482 33662 -1478 33708
rect -1458 33662 -1454 33708
rect -1434 33662 -1430 33708
rect -1410 33662 -1406 33708
rect -1386 33662 -1382 33708
rect -1362 33662 -1358 33708
rect -1338 33662 -1334 33708
rect -1314 33662 -1310 33708
rect -1290 33662 -1286 33708
rect -1266 33662 -1262 33708
rect -1242 33662 -1238 33708
rect -1218 33662 -1214 33708
rect -1194 33662 -1190 33708
rect -1170 33662 -1166 33708
rect -1146 33662 -1142 33708
rect -1122 33662 -1118 33708
rect -1098 33662 -1094 33708
rect -1074 33662 -1070 33708
rect -1050 33662 -1046 33708
rect -1026 33662 -1022 33708
rect -1002 33662 -998 33708
rect -978 33662 -974 33708
rect -954 33662 -950 33708
rect -930 33662 -926 33708
rect -906 33662 -902 33708
rect -882 33662 -878 33708
rect -858 33662 -854 33708
rect -834 33662 -830 33708
rect -810 33662 -806 33708
rect -786 33662 -782 33708
rect -762 33662 -758 33708
rect -738 33662 -734 33708
rect -714 33662 -710 33708
rect -690 33662 -686 33708
rect -666 33662 -662 33708
rect -642 33662 -638 33708
rect -618 33662 -614 33708
rect -594 33662 -590 33708
rect -570 33662 -566 33708
rect -546 33662 -542 33708
rect -522 33662 -518 33708
rect -498 33662 -494 33708
rect -474 33662 -470 33708
rect -450 33662 -446 33708
rect -426 33662 -422 33708
rect -402 33662 -398 33708
rect -378 33662 -374 33708
rect -354 33662 -350 33708
rect -330 33662 -326 33708
rect -306 33662 -302 33708
rect -282 33662 -278 33708
rect -258 33662 -254 33708
rect -234 33662 -230 33708
rect -210 33662 -206 33708
rect -186 33662 -182 33708
rect -162 33662 -158 33708
rect -138 33662 -134 33708
rect -114 33662 -110 33708
rect -90 33662 -86 33708
rect -66 33662 -62 33708
rect -42 33662 -38 33708
rect -18 33662 -14 33708
rect 6 33662 10 33708
rect 30 33662 34 33708
rect 54 33662 58 33708
rect 78 33662 82 33708
rect 102 33662 106 33708
rect 126 33662 130 33708
rect 150 33662 154 33708
rect 174 33662 178 33708
rect 198 33662 202 33708
rect 222 33662 226 33708
rect 246 33662 250 33708
rect 259 33677 264 33687
rect 270 33677 274 33708
rect 269 33663 274 33677
rect 270 33662 274 33663
rect 294 33662 298 33708
rect 318 33662 322 33708
rect 342 33662 346 33708
rect 366 33662 370 33708
rect 390 33662 394 33708
rect 414 33662 418 33708
rect 438 33662 442 33708
rect 462 33662 466 33708
rect 486 33662 490 33708
rect 510 33662 514 33708
rect 534 33662 538 33708
rect 558 33662 562 33708
rect 582 33662 586 33708
rect 606 33662 610 33708
rect 630 33662 634 33708
rect 654 33662 658 33708
rect 678 33662 682 33708
rect 702 33662 706 33708
rect 726 33662 730 33708
rect 750 33662 754 33708
rect 774 33662 778 33708
rect 781 33707 795 33708
rect 798 33707 805 33755
rect 798 33662 802 33707
rect 822 33662 826 33876
rect 846 33662 850 33876
rect 870 33662 874 33876
rect 894 33662 898 33876
rect 918 33662 922 33876
rect 942 33662 946 33876
rect 966 33662 970 33876
rect 990 33662 994 33876
rect 1014 33662 1018 33876
rect 1027 33749 1032 33759
rect 1038 33749 1042 33876
rect 1037 33735 1042 33749
rect 1038 33662 1042 33735
rect 1062 33683 1066 33876
rect -2393 33660 1059 33662
rect -2371 33590 -2366 33660
rect -2348 33590 -2343 33660
rect -2325 33656 -2320 33660
rect -2309 33658 -2301 33660
rect -2317 33656 -2309 33658
rect -2325 33644 -2317 33656
rect -2325 33596 -2320 33644
rect -2317 33642 -2309 33644
rect -2092 33630 -2062 33632
rect -2094 33626 -2062 33630
rect -2084 33604 -2054 33606
rect -2325 33590 -2317 33596
rect -2000 33590 -1992 33660
rect -1655 33658 -1647 33660
rect -1663 33656 -1655 33658
rect -1671 33644 -1663 33656
rect -1663 33642 -1655 33644
rect -1854 33630 -1806 33632
rect -1854 33626 -1680 33630
rect -1768 33606 -1700 33609
rect -1846 33604 -1700 33606
rect -1674 33590 -1663 33596
rect -1642 33590 -1637 33660
rect -1619 33590 -1614 33660
rect -1530 33590 -1526 33660
rect -1506 33590 -1502 33660
rect -1482 33590 -1478 33660
rect -1458 33590 -1454 33660
rect -1434 33590 -1430 33660
rect -1410 33590 -1406 33660
rect -1386 33590 -1382 33660
rect -1362 33590 -1358 33660
rect -1338 33590 -1334 33660
rect -1314 33590 -1310 33660
rect -1290 33590 -1286 33660
rect -1266 33590 -1262 33660
rect -1242 33590 -1238 33660
rect -1218 33590 -1214 33660
rect -1194 33590 -1190 33660
rect -1170 33590 -1166 33660
rect -1146 33590 -1142 33660
rect -1122 33590 -1118 33660
rect -1098 33590 -1094 33660
rect -1074 33590 -1070 33660
rect -1050 33590 -1046 33660
rect -1026 33590 -1022 33660
rect -1002 33590 -998 33660
rect -978 33590 -974 33660
rect -954 33590 -950 33660
rect -930 33590 -926 33660
rect -906 33590 -902 33660
rect -882 33590 -878 33660
rect -858 33590 -854 33660
rect -834 33590 -830 33660
rect -810 33590 -806 33660
rect -786 33590 -782 33660
rect -762 33590 -758 33660
rect -738 33590 -734 33660
rect -714 33590 -710 33660
rect -690 33590 -686 33660
rect -666 33590 -662 33660
rect -642 33590 -638 33660
rect -618 33590 -614 33660
rect -594 33590 -590 33660
rect -570 33590 -566 33660
rect -546 33590 -542 33660
rect -522 33590 -518 33660
rect -498 33590 -494 33660
rect -474 33590 -470 33660
rect -450 33590 -446 33660
rect -426 33590 -422 33660
rect -402 33590 -398 33660
rect -378 33590 -374 33660
rect -354 33590 -350 33660
rect -330 33590 -326 33660
rect -306 33590 -302 33660
rect -282 33590 -278 33660
rect -258 33590 -254 33660
rect -234 33590 -230 33660
rect -210 33590 -206 33660
rect -186 33590 -182 33660
rect -162 33590 -158 33660
rect -138 33590 -134 33660
rect -114 33590 -110 33660
rect -90 33590 -86 33660
rect -66 33590 -62 33660
rect -42 33590 -38 33660
rect -18 33590 -14 33660
rect 6 33590 10 33660
rect 30 33590 34 33660
rect 54 33590 58 33660
rect 78 33590 82 33660
rect 102 33590 106 33660
rect 126 33590 130 33660
rect 150 33590 154 33660
rect 174 33590 178 33660
rect 198 33590 202 33660
rect 222 33590 226 33660
rect 246 33590 250 33660
rect 270 33590 274 33660
rect 294 33611 298 33660
rect -2393 33588 -1946 33590
rect -1932 33588 291 33590
rect -2371 33566 -2366 33588
rect -2348 33566 -2343 33588
rect -2325 33586 -2317 33588
rect -2054 33586 -2004 33588
rect -2000 33586 -1966 33588
rect -2325 33568 -2320 33586
rect -2317 33580 -2306 33586
rect -2307 33570 -2306 33580
rect -2084 33575 -2054 33580
rect -2084 33568 -2054 33569
rect -2325 33566 -2317 33568
rect -2024 33566 -2014 33575
rect -2000 33566 -1992 33586
rect -1982 33585 -1966 33586
rect -1663 33580 -1658 33588
rect -1846 33575 -1798 33580
rect -1784 33568 -1780 33573
rect -1923 33566 -1889 33567
rect -1674 33566 -1663 33568
rect -1642 33566 -1637 33588
rect -1619 33566 -1614 33588
rect -1530 33566 -1526 33588
rect -1506 33566 -1502 33588
rect -1482 33566 -1478 33588
rect -1458 33566 -1454 33588
rect -1434 33566 -1430 33588
rect -1410 33566 -1406 33588
rect -1386 33566 -1382 33588
rect -1362 33566 -1358 33588
rect -1338 33566 -1334 33588
rect -1314 33566 -1310 33588
rect -1290 33566 -1286 33588
rect -1266 33566 -1262 33588
rect -1242 33566 -1238 33588
rect -1218 33566 -1214 33588
rect -1194 33566 -1190 33588
rect -1170 33566 -1166 33588
rect -1146 33566 -1142 33588
rect -1122 33566 -1118 33588
rect -1098 33566 -1094 33588
rect -1074 33566 -1070 33588
rect -1050 33566 -1046 33588
rect -1026 33566 -1022 33588
rect -1002 33566 -998 33588
rect -978 33566 -974 33588
rect -954 33566 -950 33588
rect -930 33566 -926 33588
rect -906 33566 -902 33588
rect -882 33566 -878 33588
rect -858 33566 -854 33588
rect -834 33566 -830 33588
rect -810 33566 -806 33588
rect -786 33566 -782 33588
rect -762 33566 -758 33588
rect -738 33566 -734 33588
rect -714 33566 -710 33588
rect -690 33566 -686 33588
rect -666 33566 -662 33588
rect -642 33566 -638 33588
rect -618 33566 -614 33588
rect -594 33566 -590 33588
rect -570 33566 -566 33588
rect -546 33566 -542 33588
rect -522 33566 -518 33588
rect -498 33566 -494 33588
rect -474 33566 -470 33588
rect -450 33566 -446 33588
rect -426 33566 -422 33588
rect -402 33566 -398 33588
rect -378 33566 -374 33588
rect -354 33566 -350 33588
rect -330 33566 -326 33588
rect -306 33566 -302 33588
rect -282 33566 -278 33588
rect -258 33566 -254 33588
rect -234 33566 -230 33588
rect -210 33566 -206 33588
rect -186 33566 -182 33588
rect -162 33566 -158 33588
rect -138 33566 -134 33588
rect -114 33566 -110 33588
rect -90 33566 -86 33588
rect -66 33566 -62 33588
rect -42 33567 -38 33588
rect -53 33566 -19 33567
rect -2393 33564 -19 33566
rect -2371 33494 -2366 33564
rect -2348 33494 -2343 33564
rect -2325 33558 -2317 33564
rect -2154 33562 -2138 33564
rect -2325 33510 -2320 33558
rect -2317 33552 -2306 33558
rect -2149 33555 -2138 33562
rect -2154 33550 -2138 33552
rect -2084 33550 -2054 33564
rect -2153 33532 -2147 33534
rect -2153 33530 -2101 33532
rect -2153 33524 -2054 33530
rect -2307 33514 -2306 33522
rect -2325 33502 -2314 33510
rect -2104 33506 -2101 33510
rect -2104 33504 -2101 33505
rect -2000 33504 -1992 33564
rect -1674 33561 -1663 33564
rect -1846 33550 -1798 33554
rect -1663 33552 -1658 33561
rect -1758 33527 -1692 33533
rect -1758 33524 -1710 33527
rect -1750 33515 -1702 33522
rect -1917 33508 -1901 33514
rect -1828 33510 -1792 33514
rect -1916 33504 -1914 33508
rect -1750 33507 -1710 33513
rect -1700 33507 -1692 33527
rect -1674 33516 -1665 33525
rect -1674 33504 -1666 33513
rect -2325 33494 -2320 33502
rect -2314 33494 -2306 33502
rect -2139 33495 -2123 33504
rect -2111 33497 -2016 33504
rect -2139 33494 -2111 33495
rect -2104 33494 -2101 33497
rect -2021 33494 -2016 33497
rect -2000 33497 -1818 33504
rect -1802 33497 -1776 33504
rect -1760 33497 -1710 33504
rect -1666 33497 -1658 33504
rect -2000 33494 -1992 33497
rect -1758 33495 -1755 33497
rect -1758 33494 -1757 33495
rect -1710 33494 -1702 33495
rect -1674 33494 -1665 33497
rect -1642 33494 -1637 33564
rect -1619 33494 -1614 33564
rect -1530 33494 -1526 33564
rect -1506 33494 -1502 33564
rect -1482 33494 -1478 33564
rect -1458 33494 -1454 33564
rect -1434 33494 -1430 33564
rect -1410 33494 -1406 33564
rect -1386 33494 -1382 33564
rect -1362 33494 -1358 33564
rect -1338 33494 -1334 33564
rect -1314 33494 -1310 33564
rect -1290 33494 -1286 33564
rect -1266 33494 -1262 33564
rect -1242 33494 -1238 33564
rect -1218 33494 -1214 33564
rect -1194 33494 -1190 33564
rect -1170 33494 -1166 33564
rect -1146 33494 -1142 33564
rect -1122 33494 -1118 33564
rect -1098 33494 -1094 33564
rect -1074 33494 -1070 33564
rect -1050 33494 -1046 33564
rect -1026 33494 -1022 33564
rect -1002 33494 -998 33564
rect -978 33494 -974 33564
rect -954 33494 -950 33564
rect -930 33494 -926 33564
rect -906 33494 -902 33564
rect -882 33494 -878 33564
rect -858 33494 -854 33564
rect -845 33509 -840 33519
rect -834 33509 -830 33564
rect -835 33495 -830 33509
rect -834 33494 -830 33495
rect -810 33494 -806 33564
rect -786 33494 -782 33564
rect -762 33494 -758 33564
rect -738 33494 -734 33564
rect -714 33494 -710 33564
rect -690 33494 -686 33564
rect -666 33494 -662 33564
rect -642 33494 -638 33564
rect -618 33494 -614 33564
rect -594 33494 -590 33564
rect -570 33494 -566 33564
rect -546 33494 -542 33564
rect -522 33494 -518 33564
rect -498 33494 -494 33564
rect -474 33494 -470 33564
rect -450 33494 -446 33564
rect -426 33494 -422 33564
rect -402 33494 -398 33564
rect -378 33494 -374 33564
rect -354 33494 -350 33564
rect -330 33494 -326 33564
rect -306 33494 -302 33564
rect -282 33494 -278 33564
rect -258 33494 -254 33564
rect -234 33494 -230 33564
rect -210 33494 -206 33564
rect -186 33494 -182 33564
rect -162 33494 -158 33564
rect -138 33494 -134 33564
rect -114 33494 -110 33564
rect -90 33494 -86 33564
rect -66 33494 -62 33564
rect -53 33557 -48 33564
rect -42 33557 -38 33564
rect -43 33543 -38 33557
rect -42 33494 -38 33543
rect -18 33494 -14 33588
rect 6 33494 10 33588
rect 30 33494 34 33588
rect 54 33494 58 33588
rect 78 33494 82 33588
rect 102 33494 106 33588
rect 126 33494 130 33588
rect 150 33494 154 33588
rect 174 33494 178 33588
rect 198 33494 202 33588
rect 222 33494 226 33588
rect 246 33494 250 33588
rect 270 33495 274 33588
rect 277 33587 291 33588
rect 294 33587 301 33611
rect 259 33494 293 33495
rect -2393 33492 293 33494
rect -2371 33422 -2366 33492
rect -2348 33422 -2343 33492
rect -2325 33482 -2320 33492
rect -2307 33486 -2306 33492
rect -2139 33488 -2111 33492
rect -2325 33474 -2314 33482
rect -2141 33479 -2119 33483
rect -2325 33454 -2320 33474
rect -2314 33466 -2306 33474
rect -2149 33467 -2141 33474
rect -2307 33458 -2306 33466
rect -2104 33464 -2101 33492
rect -2076 33488 -2046 33491
rect -2076 33475 -2054 33483
rect -2021 33480 -2016 33492
rect -2084 33473 -2036 33474
rect -2000 33473 -1992 33492
rect -1931 33488 -1895 33492
rect -1768 33484 -1760 33492
rect -1758 33488 -1757 33492
rect -1750 33488 -1702 33492
rect -1674 33488 -1665 33492
rect -1768 33483 -1764 33484
rect -1758 33483 -1755 33488
rect -1932 33473 -1917 33482
rect -2084 33470 -1917 33473
rect -1916 33473 -1905 33475
rect -1758 33474 -1754 33483
rect -1750 33476 -1710 33483
rect -1674 33476 -1666 33485
rect -1758 33473 -1692 33474
rect -1916 33471 -1692 33473
rect -1916 33470 -1690 33471
rect -2084 33466 -2054 33470
rect -2046 33466 -1932 33470
rect -1921 33466 -1710 33470
rect -1680 33468 -1672 33471
rect -1666 33469 -1658 33476
rect -2054 33464 -2046 33465
rect -2155 33458 -2139 33464
rect -2076 33458 -2046 33464
rect -2325 33446 -2314 33454
rect -2149 33448 -2139 33458
rect -2076 33448 -2054 33456
rect -2325 33426 -2320 33446
rect -2314 33438 -2306 33446
rect -2104 33443 -2054 33446
rect -2084 33440 -2054 33443
rect -2307 33430 -2306 33438
rect -2325 33422 -2314 33426
rect -2000 33422 -1992 33466
rect -1710 33464 -1702 33465
rect -1750 33458 -1702 33464
rect -1680 33460 -1665 33468
rect -1919 33456 -1916 33458
rect -1680 33456 -1672 33460
rect -1932 33454 -1916 33456
rect -1750 33448 -1710 33456
rect -1674 33448 -1666 33456
rect -1837 33440 -1789 33446
rect -1760 33444 -1692 33447
rect -1764 33440 -1692 33444
rect -1666 33440 -1658 33448
rect -1680 33432 -1665 33440
rect -1926 33422 -1892 33425
rect -1680 33422 -1672 33432
rect -1671 33422 -1666 33428
rect -1642 33422 -1637 33492
rect -1619 33422 -1614 33492
rect -1530 33422 -1526 33492
rect -1506 33422 -1502 33492
rect -1482 33422 -1478 33492
rect -1458 33422 -1454 33492
rect -1434 33422 -1430 33492
rect -1410 33422 -1406 33492
rect -1386 33422 -1382 33492
rect -1362 33422 -1358 33492
rect -1338 33422 -1334 33492
rect -1314 33422 -1310 33492
rect -1290 33422 -1286 33492
rect -1266 33422 -1262 33492
rect -1242 33422 -1238 33492
rect -1218 33422 -1214 33492
rect -1194 33422 -1190 33492
rect -1170 33422 -1166 33492
rect -1146 33422 -1142 33492
rect -1122 33422 -1118 33492
rect -1098 33422 -1094 33492
rect -1074 33422 -1070 33492
rect -1050 33422 -1046 33492
rect -1026 33422 -1022 33492
rect -1002 33422 -998 33492
rect -978 33422 -974 33492
rect -954 33422 -950 33492
rect -930 33422 -926 33492
rect -906 33422 -902 33492
rect -882 33422 -878 33492
rect -858 33422 -854 33492
rect -834 33422 -830 33492
rect -810 33443 -806 33492
rect -2393 33420 -813 33422
rect -2371 33398 -2366 33420
rect -2348 33398 -2343 33420
rect -2325 33414 -2314 33420
rect -2325 33398 -2320 33414
rect -2314 33410 -2309 33414
rect -2070 33412 -2046 33413
rect -2309 33398 -2298 33410
rect -2046 33407 -2038 33411
rect -2068 33398 -2046 33407
rect -2011 33400 -2003 33402
rect -2000 33400 -1992 33420
rect -1908 33418 -1894 33420
rect -1923 33408 -1916 33415
rect -1810 33412 -1801 33414
rect -1934 33402 -1923 33404
rect -1916 33401 -1909 33408
rect -1852 33407 -1804 33411
rect -2025 33399 -1991 33400
rect -2025 33398 -1975 33399
rect -1829 33398 -1804 33407
rect -1680 33398 -1672 33420
rect -1671 33414 -1666 33420
rect -1666 33412 -1655 33414
rect -1655 33400 -1650 33412
rect -1666 33398 -1655 33400
rect -1642 33398 -1637 33420
rect -1619 33398 -1614 33420
rect -1530 33398 -1526 33420
rect -1506 33398 -1502 33420
rect -1482 33398 -1478 33420
rect -1458 33398 -1454 33420
rect -1434 33398 -1430 33420
rect -1410 33398 -1406 33420
rect -1386 33398 -1382 33420
rect -1362 33398 -1358 33420
rect -1338 33398 -1334 33420
rect -1314 33398 -1310 33420
rect -1290 33398 -1286 33420
rect -1266 33398 -1262 33420
rect -1242 33398 -1238 33420
rect -1218 33398 -1214 33420
rect -1194 33398 -1190 33420
rect -1170 33398 -1166 33420
rect -1146 33398 -1142 33420
rect -1122 33398 -1118 33420
rect -1098 33398 -1094 33420
rect -1074 33398 -1070 33420
rect -1050 33398 -1046 33420
rect -1026 33398 -1022 33420
rect -1002 33398 -998 33420
rect -978 33398 -974 33420
rect -954 33398 -950 33420
rect -930 33398 -926 33420
rect -906 33398 -902 33420
rect -882 33398 -878 33420
rect -858 33398 -854 33420
rect -834 33398 -830 33420
rect -827 33419 -813 33420
rect -810 33419 -803 33443
rect -810 33398 -806 33419
rect -786 33398 -782 33492
rect -762 33398 -758 33492
rect -738 33398 -734 33492
rect -714 33398 -710 33492
rect -690 33398 -686 33492
rect -666 33398 -662 33492
rect -642 33398 -638 33492
rect -618 33398 -614 33492
rect -594 33398 -590 33492
rect -570 33398 -566 33492
rect -546 33398 -542 33492
rect -522 33398 -518 33492
rect -498 33398 -494 33492
rect -474 33398 -470 33492
rect -450 33398 -446 33492
rect -426 33398 -422 33492
rect -402 33398 -398 33492
rect -378 33398 -374 33492
rect -354 33398 -350 33492
rect -330 33398 -326 33492
rect -306 33398 -302 33492
rect -282 33398 -278 33492
rect -258 33398 -254 33492
rect -234 33398 -230 33492
rect -210 33398 -206 33492
rect -186 33398 -182 33492
rect -162 33398 -158 33492
rect -138 33398 -134 33492
rect -114 33398 -110 33492
rect -90 33398 -86 33492
rect -66 33398 -62 33492
rect -42 33398 -38 33492
rect -18 33491 -14 33492
rect -18 33467 -11 33491
rect -18 33398 -14 33467
rect 6 33398 10 33492
rect 30 33398 34 33492
rect 54 33398 58 33492
rect 78 33398 82 33492
rect 102 33398 106 33492
rect 126 33398 130 33492
rect 150 33398 154 33492
rect 174 33398 178 33492
rect 187 33437 192 33447
rect 198 33437 202 33492
rect 197 33423 202 33437
rect 187 33413 192 33423
rect 197 33399 202 33413
rect 198 33398 202 33399
rect 222 33398 226 33492
rect 246 33398 250 33492
rect 259 33485 264 33492
rect 270 33485 274 33492
rect 269 33471 274 33485
rect 270 33398 274 33471
rect 294 33419 298 33587
rect -2393 33396 291 33398
rect -2371 33302 -2366 33396
rect -2348 33302 -2343 33396
rect -2325 33386 -2314 33396
rect -2068 33395 -2046 33396
rect -2025 33394 -2003 33396
rect -2076 33391 -2046 33393
rect -2076 33389 -2068 33391
rect -2068 33386 -2046 33389
rect -2325 33370 -2320 33386
rect -2314 33382 -2309 33386
rect -2046 33382 -2038 33386
rect -2309 33370 -2298 33382
rect -2325 33358 -2314 33370
rect -2076 33364 -2046 33366
rect -2325 33338 -2320 33358
rect -2314 33354 -2309 33358
rect -2325 33330 -2317 33338
rect -2060 33332 -2030 33335
rect -2325 33302 -2320 33330
rect -2317 33322 -2309 33330
rect -2060 33319 -2038 33330
rect -2033 33323 -2030 33332
rect -2028 33328 -2027 33332
rect -2068 33314 -2038 33317
rect -2000 33302 -1992 33396
rect -1923 33394 -1909 33396
rect -1829 33395 -1804 33396
rect -1680 33394 -1672 33396
rect -1804 33393 -1781 33394
rect -1829 33391 -1781 33393
rect -1750 33391 -1702 33394
rect -1804 33389 -1796 33391
rect -1829 33386 -1804 33389
rect -1671 33386 -1666 33396
rect -1852 33384 -1829 33386
rect -1666 33384 -1655 33386
rect -1852 33382 -1804 33384
rect -1829 33368 -1804 33380
rect -1655 33372 -1650 33384
rect -1666 33370 -1655 33372
rect -1829 33364 -1794 33367
rect -1671 33358 -1666 33370
rect -1666 33356 -1655 33358
rect -1912 33347 -1884 33349
rect -1852 33341 -1804 33345
rect -1844 33332 -1796 33335
rect -1671 33330 -1663 33338
rect -1844 33319 -1804 33330
rect -1663 33322 -1655 33330
rect -1852 33314 -1680 33318
rect -1642 33302 -1637 33396
rect -1619 33302 -1614 33396
rect -1530 33302 -1526 33396
rect -1506 33302 -1502 33396
rect -1482 33302 -1478 33396
rect -1458 33302 -1454 33396
rect -1434 33302 -1430 33396
rect -1410 33302 -1406 33396
rect -1386 33302 -1382 33396
rect -1362 33302 -1358 33396
rect -1338 33302 -1334 33396
rect -1314 33302 -1310 33396
rect -1290 33302 -1286 33396
rect -1266 33302 -1262 33396
rect -1242 33302 -1238 33396
rect -1218 33302 -1214 33396
rect -1194 33302 -1190 33396
rect -1170 33302 -1166 33396
rect -1146 33302 -1142 33396
rect -1133 33365 -1128 33375
rect -1122 33365 -1118 33396
rect -1123 33351 -1118 33365
rect -1122 33302 -1118 33351
rect -1098 33302 -1094 33396
rect -1074 33302 -1070 33396
rect -1050 33302 -1046 33396
rect -1026 33302 -1022 33396
rect -1002 33302 -998 33396
rect -978 33302 -974 33396
rect -954 33302 -950 33396
rect -930 33302 -926 33396
rect -906 33302 -902 33396
rect -882 33302 -878 33396
rect -858 33302 -854 33396
rect -834 33302 -830 33396
rect -810 33302 -806 33396
rect -797 33341 -792 33351
rect -786 33341 -782 33396
rect -787 33327 -782 33341
rect -786 33302 -782 33327
rect -762 33302 -758 33396
rect -738 33302 -734 33396
rect -714 33302 -710 33396
rect -690 33302 -686 33396
rect -666 33302 -662 33396
rect -642 33302 -638 33396
rect -618 33302 -614 33396
rect -594 33302 -590 33396
rect -570 33302 -566 33396
rect -546 33302 -542 33396
rect -522 33302 -518 33396
rect -498 33302 -494 33396
rect -474 33302 -470 33396
rect -450 33302 -446 33396
rect -426 33302 -422 33396
rect -402 33302 -398 33396
rect -378 33302 -374 33396
rect -354 33302 -350 33396
rect -330 33302 -326 33396
rect -306 33302 -302 33396
rect -282 33302 -278 33396
rect -258 33302 -254 33396
rect -234 33302 -230 33396
rect -210 33302 -206 33396
rect -186 33302 -182 33396
rect -162 33302 -158 33396
rect -138 33302 -134 33396
rect -114 33302 -110 33396
rect -90 33302 -86 33396
rect -66 33302 -62 33396
rect -42 33302 -38 33396
rect -18 33302 -14 33396
rect 6 33302 10 33396
rect 30 33302 34 33396
rect 54 33302 58 33396
rect 78 33302 82 33396
rect 102 33302 106 33396
rect 126 33302 130 33396
rect 150 33302 154 33396
rect 174 33302 178 33396
rect 198 33302 202 33396
rect 222 33371 226 33396
rect 222 33323 229 33371
rect 222 33302 226 33323
rect 246 33302 250 33396
rect 270 33302 274 33396
rect 277 33395 291 33396
rect 294 33395 301 33419
rect 294 33302 298 33395
rect 318 33302 322 33660
rect 342 33302 346 33660
rect 366 33302 370 33660
rect 390 33302 394 33660
rect 414 33302 418 33660
rect 438 33302 442 33660
rect 462 33302 466 33660
rect 486 33302 490 33660
rect 499 33317 504 33327
rect 510 33317 514 33660
rect 509 33303 514 33317
rect 499 33302 533 33303
rect -2393 33300 533 33302
rect -2371 33278 -2366 33300
rect -2348 33278 -2343 33300
rect -2325 33278 -2320 33300
rect -2309 33282 -2301 33292
rect -2068 33283 -2062 33288
rect -2317 33278 -2309 33282
rect -2060 33278 -2050 33283
rect -2000 33278 -1992 33300
rect -1806 33292 -1680 33298
rect -1854 33283 -1806 33288
rect -1655 33282 -1647 33292
rect -1972 33278 -1964 33279
rect -1958 33278 -1942 33280
rect -1844 33278 -1806 33281
rect -1663 33278 -1655 33282
rect -1642 33278 -1637 33300
rect -1619 33278 -1614 33300
rect -1530 33278 -1526 33300
rect -1506 33278 -1502 33300
rect -1482 33278 -1478 33300
rect -1458 33278 -1454 33300
rect -1434 33278 -1430 33300
rect -1410 33278 -1406 33300
rect -1386 33278 -1382 33300
rect -1362 33278 -1358 33300
rect -1338 33278 -1334 33300
rect -1314 33278 -1310 33300
rect -1290 33278 -1286 33300
rect -1266 33278 -1262 33300
rect -1242 33278 -1238 33300
rect -1218 33278 -1214 33300
rect -1194 33278 -1190 33300
rect -1170 33278 -1166 33300
rect -1146 33278 -1142 33300
rect -1122 33278 -1118 33300
rect -1098 33299 -1094 33300
rect -2393 33276 -1101 33278
rect -2371 33254 -2366 33276
rect -2348 33254 -2343 33276
rect -2325 33254 -2320 33276
rect -2060 33270 -2050 33276
rect -2309 33254 -2301 33264
rect -2060 33263 -2030 33270
rect -2000 33266 -1992 33276
rect -1972 33274 -1942 33276
rect -1958 33273 -1942 33274
rect -1844 33272 -1806 33276
rect -2068 33256 -2062 33263
rect -2062 33254 -2036 33256
rect -2393 33252 -2036 33254
rect -2030 33254 -2012 33256
rect -2004 33254 -1990 33266
rect -1844 33265 -1798 33270
rect -1806 33263 -1798 33265
rect -1854 33261 -1844 33263
rect -1854 33256 -1806 33261
rect -1864 33254 -1796 33255
rect -1655 33254 -1647 33264
rect -1642 33254 -1637 33276
rect -1619 33254 -1614 33276
rect -1530 33254 -1526 33276
rect -1506 33254 -1502 33276
rect -1482 33254 -1478 33276
rect -1458 33254 -1454 33276
rect -1434 33254 -1430 33276
rect -1410 33254 -1406 33276
rect -1386 33254 -1382 33276
rect -1362 33254 -1358 33276
rect -1338 33254 -1334 33276
rect -1314 33254 -1310 33276
rect -1290 33254 -1286 33276
rect -1266 33254 -1262 33276
rect -1242 33254 -1238 33276
rect -1218 33254 -1214 33276
rect -1194 33254 -1190 33276
rect -1170 33254 -1166 33276
rect -1146 33254 -1142 33276
rect -1122 33254 -1118 33276
rect -1115 33275 -1101 33276
rect -1098 33275 -1091 33299
rect -1098 33254 -1094 33275
rect -1074 33254 -1070 33300
rect -1050 33254 -1046 33300
rect -1026 33254 -1022 33300
rect -1002 33254 -998 33300
rect -978 33254 -974 33300
rect -954 33254 -950 33300
rect -930 33254 -926 33300
rect -906 33254 -902 33300
rect -882 33254 -878 33300
rect -858 33254 -854 33300
rect -834 33254 -830 33300
rect -810 33254 -806 33300
rect -786 33254 -782 33300
rect -762 33275 -758 33300
rect -2030 33252 -765 33254
rect -2371 33206 -2366 33252
rect -2348 33206 -2343 33252
rect -2325 33206 -2320 33252
rect -2317 33248 -2309 33252
rect -2060 33248 -2050 33252
rect -2060 33246 -2036 33248
rect -2060 33244 -2030 33246
rect -2292 33238 -2030 33244
rect -2092 33222 -2062 33224
rect -2094 33218 -2062 33222
rect -2000 33206 -1992 33252
rect -1844 33245 -1806 33252
rect -1663 33248 -1655 33252
rect -1844 33238 -1680 33244
rect -1854 33222 -1806 33224
rect -1854 33218 -1680 33222
rect -1642 33206 -1637 33252
rect -1619 33206 -1614 33252
rect -1530 33206 -1526 33252
rect -1506 33206 -1502 33252
rect -1482 33206 -1478 33252
rect -1458 33206 -1454 33252
rect -1434 33206 -1430 33252
rect -1410 33206 -1406 33252
rect -1386 33206 -1382 33252
rect -1362 33206 -1358 33252
rect -1338 33206 -1334 33252
rect -1314 33206 -1310 33252
rect -1290 33206 -1286 33252
rect -1266 33206 -1262 33252
rect -1242 33206 -1238 33252
rect -1218 33206 -1214 33252
rect -1194 33206 -1190 33252
rect -1170 33206 -1166 33252
rect -1146 33206 -1142 33252
rect -1122 33206 -1118 33252
rect -1098 33206 -1094 33252
rect -1074 33206 -1070 33252
rect -1050 33206 -1046 33252
rect -1026 33206 -1022 33252
rect -1002 33206 -998 33252
rect -978 33206 -974 33252
rect -954 33206 -950 33252
rect -930 33206 -926 33252
rect -906 33206 -902 33252
rect -882 33206 -878 33252
rect -858 33206 -854 33252
rect -834 33206 -830 33252
rect -810 33206 -806 33252
rect -786 33206 -782 33252
rect -779 33251 -765 33252
rect -762 33251 -755 33275
rect -762 33206 -758 33251
rect -738 33206 -734 33300
rect -714 33206 -710 33300
rect -690 33206 -686 33300
rect -666 33206 -662 33300
rect -642 33206 -638 33300
rect -618 33206 -614 33300
rect -594 33206 -590 33300
rect -570 33206 -566 33300
rect -546 33206 -542 33300
rect -522 33206 -518 33300
rect -498 33206 -494 33300
rect -474 33206 -470 33300
rect -450 33206 -446 33300
rect -426 33206 -422 33300
rect -402 33206 -398 33300
rect -378 33206 -374 33300
rect -354 33206 -350 33300
rect -330 33206 -326 33300
rect -306 33206 -302 33300
rect -282 33206 -278 33300
rect -258 33206 -254 33300
rect -234 33206 -230 33300
rect -210 33206 -206 33300
rect -186 33206 -182 33300
rect -162 33206 -158 33300
rect -138 33206 -134 33300
rect -114 33206 -110 33300
rect -90 33206 -86 33300
rect -66 33206 -62 33300
rect -42 33206 -38 33300
rect -18 33206 -14 33300
rect 6 33206 10 33300
rect 30 33206 34 33300
rect 54 33206 58 33300
rect 78 33206 82 33300
rect 102 33206 106 33300
rect 126 33206 130 33300
rect 150 33206 154 33300
rect 174 33206 178 33300
rect 198 33206 202 33300
rect 222 33206 226 33300
rect 246 33206 250 33300
rect 270 33206 274 33300
rect 294 33206 298 33300
rect 318 33206 322 33300
rect 342 33206 346 33300
rect 366 33206 370 33300
rect 390 33206 394 33300
rect 414 33206 418 33300
rect 438 33206 442 33300
rect 462 33206 466 33300
rect 486 33206 490 33300
rect 499 33293 504 33300
rect 509 33279 514 33293
rect 510 33206 514 33279
rect 534 33251 538 33660
rect -2393 33204 531 33206
rect -2371 33182 -2366 33204
rect -2348 33182 -2343 33204
rect -2325 33182 -2320 33204
rect -2072 33202 -2036 33203
rect -2072 33196 -2054 33202
rect -2309 33188 -2301 33196
rect -2317 33182 -2309 33188
rect -2092 33187 -2062 33192
rect -2000 33183 -1992 33204
rect -1938 33203 -1906 33204
rect -1920 33202 -1906 33203
rect -1806 33196 -1680 33202
rect -1854 33187 -1806 33192
rect -1655 33188 -1647 33196
rect -1982 33183 -1966 33184
rect -2000 33182 -1966 33183
rect -1846 33182 -1806 33185
rect -1663 33182 -1655 33188
rect -1642 33182 -1637 33204
rect -1619 33182 -1614 33204
rect -1530 33182 -1526 33204
rect -1506 33182 -1502 33204
rect -1482 33182 -1478 33204
rect -1458 33182 -1454 33204
rect -1434 33182 -1430 33204
rect -1410 33182 -1406 33204
rect -1386 33182 -1382 33204
rect -1362 33182 -1358 33204
rect -1338 33182 -1334 33204
rect -1314 33182 -1310 33204
rect -1290 33182 -1286 33204
rect -1266 33182 -1262 33204
rect -1242 33182 -1238 33204
rect -1218 33182 -1214 33204
rect -1194 33182 -1190 33204
rect -1170 33182 -1166 33204
rect -1146 33182 -1142 33204
rect -1122 33182 -1118 33204
rect -1098 33183 -1094 33204
rect -1109 33182 -1075 33183
rect -2393 33180 -1075 33182
rect -2371 33158 -2366 33180
rect -2348 33158 -2343 33180
rect -2325 33158 -2320 33180
rect -2000 33178 -1966 33180
rect -2309 33160 -2301 33168
rect -2062 33167 -2054 33174
rect -2092 33160 -2084 33167
rect -2062 33160 -2026 33162
rect -2317 33158 -2309 33160
rect -2062 33158 -2012 33160
rect -2000 33158 -1992 33178
rect -1982 33177 -1966 33178
rect -1846 33176 -1806 33180
rect -1846 33169 -1798 33174
rect -1806 33167 -1798 33169
rect -1854 33165 -1846 33167
rect -1854 33160 -1806 33165
rect -1655 33160 -1647 33168
rect -1864 33158 -1796 33159
rect -1663 33158 -1655 33160
rect -1642 33158 -1637 33180
rect -1619 33158 -1614 33180
rect -1530 33158 -1526 33180
rect -1506 33158 -1502 33180
rect -1482 33158 -1478 33180
rect -1458 33158 -1454 33180
rect -1434 33158 -1430 33180
rect -1410 33158 -1406 33180
rect -1386 33158 -1382 33180
rect -1362 33158 -1358 33180
rect -1338 33158 -1334 33180
rect -1314 33158 -1310 33180
rect -1290 33158 -1286 33180
rect -1266 33158 -1262 33180
rect -1242 33158 -1238 33180
rect -1218 33158 -1214 33180
rect -1194 33158 -1190 33180
rect -1170 33158 -1166 33180
rect -1146 33158 -1142 33180
rect -1122 33158 -1118 33180
rect -1109 33173 -1104 33180
rect -1098 33173 -1094 33180
rect -1099 33159 -1094 33173
rect -1098 33158 -1094 33159
rect -1074 33158 -1070 33204
rect -1050 33158 -1046 33204
rect -1026 33158 -1022 33204
rect -1002 33158 -998 33204
rect -978 33158 -974 33204
rect -954 33158 -950 33204
rect -930 33158 -926 33204
rect -906 33158 -902 33204
rect -882 33158 -878 33204
rect -858 33158 -854 33204
rect -834 33158 -830 33204
rect -810 33158 -806 33204
rect -786 33158 -782 33204
rect -762 33158 -758 33204
rect -738 33158 -734 33204
rect -714 33158 -710 33204
rect -690 33158 -686 33204
rect -666 33158 -662 33204
rect -642 33158 -638 33204
rect -618 33158 -614 33204
rect -594 33158 -590 33204
rect -570 33158 -566 33204
rect -546 33158 -542 33204
rect -522 33158 -518 33204
rect -498 33158 -494 33204
rect -474 33158 -470 33204
rect -450 33158 -446 33204
rect -426 33158 -422 33204
rect -402 33158 -398 33204
rect -378 33158 -374 33204
rect -354 33158 -350 33204
rect -330 33158 -326 33204
rect -306 33158 -302 33204
rect -282 33158 -278 33204
rect -258 33158 -254 33204
rect -234 33158 -230 33204
rect -210 33158 -206 33204
rect -186 33158 -182 33204
rect -162 33158 -158 33204
rect -138 33158 -134 33204
rect -114 33158 -110 33204
rect -90 33158 -86 33204
rect -66 33158 -62 33204
rect -42 33158 -38 33204
rect -18 33158 -14 33204
rect 6 33158 10 33204
rect 30 33158 34 33204
rect 54 33158 58 33204
rect 78 33158 82 33204
rect 102 33158 106 33204
rect 126 33159 130 33204
rect 115 33158 149 33159
rect -2393 33156 149 33158
rect -2371 33110 -2366 33156
rect -2348 33110 -2343 33156
rect -2325 33110 -2320 33156
rect -2317 33152 -2309 33156
rect -2062 33152 -2054 33156
rect -2154 33148 -2138 33150
rect -2057 33148 -2054 33152
rect -2292 33142 -2054 33148
rect -2052 33142 -2044 33152
rect -2092 33126 -2062 33128
rect -2094 33122 -2062 33126
rect -2000 33110 -1992 33156
rect -1846 33149 -1806 33156
rect -1663 33152 -1655 33156
rect -1846 33142 -1680 33148
rect -1854 33126 -1806 33128
rect -1854 33122 -1680 33126
rect -1642 33110 -1637 33156
rect -1619 33110 -1614 33156
rect -1530 33110 -1526 33156
rect -1506 33110 -1502 33156
rect -1482 33110 -1478 33156
rect -1458 33110 -1454 33156
rect -1434 33110 -1430 33156
rect -1410 33110 -1406 33156
rect -1386 33110 -1382 33156
rect -1362 33110 -1358 33156
rect -1338 33110 -1334 33156
rect -1314 33110 -1310 33156
rect -1290 33110 -1286 33156
rect -1266 33110 -1262 33156
rect -1242 33110 -1238 33156
rect -1218 33110 -1214 33156
rect -1194 33110 -1190 33156
rect -1170 33110 -1166 33156
rect -1146 33110 -1142 33156
rect -1122 33110 -1118 33156
rect -1098 33110 -1094 33156
rect -1074 33110 -1070 33156
rect -1050 33110 -1046 33156
rect -1026 33110 -1022 33156
rect -1002 33110 -998 33156
rect -978 33110 -974 33156
rect -954 33110 -950 33156
rect -930 33110 -926 33156
rect -906 33110 -902 33156
rect -882 33110 -878 33156
rect -858 33110 -854 33156
rect -834 33110 -830 33156
rect -810 33110 -806 33156
rect -786 33110 -782 33156
rect -762 33110 -758 33156
rect -738 33110 -734 33156
rect -714 33110 -710 33156
rect -690 33110 -686 33156
rect -666 33110 -662 33156
rect -642 33110 -638 33156
rect -618 33110 -614 33156
rect -594 33110 -590 33156
rect -570 33110 -566 33156
rect -546 33110 -542 33156
rect -522 33110 -518 33156
rect -498 33110 -494 33156
rect -474 33110 -470 33156
rect -450 33110 -446 33156
rect -426 33110 -422 33156
rect -402 33110 -398 33156
rect -378 33110 -374 33156
rect -354 33110 -350 33156
rect -330 33110 -326 33156
rect -306 33110 -302 33156
rect -282 33110 -278 33156
rect -258 33110 -254 33156
rect -234 33110 -230 33156
rect -210 33110 -206 33156
rect -186 33110 -182 33156
rect -162 33110 -158 33156
rect -138 33110 -134 33156
rect -114 33110 -110 33156
rect -90 33110 -86 33156
rect -66 33110 -62 33156
rect -42 33110 -38 33156
rect -18 33110 -14 33156
rect 6 33110 10 33156
rect 30 33110 34 33156
rect 54 33110 58 33156
rect 78 33110 82 33156
rect 102 33110 106 33156
rect 115 33149 120 33156
rect 126 33149 130 33156
rect 125 33135 130 33149
rect 126 33110 130 33135
rect 150 33110 154 33204
rect 174 33110 178 33204
rect 198 33110 202 33204
rect 222 33110 226 33204
rect 246 33110 250 33204
rect 270 33110 274 33204
rect 294 33110 298 33204
rect 318 33110 322 33204
rect 342 33110 346 33204
rect 366 33110 370 33204
rect 390 33110 394 33204
rect 414 33110 418 33204
rect 438 33110 442 33204
rect 462 33110 466 33204
rect 486 33110 490 33204
rect 510 33110 514 33204
rect 517 33203 531 33204
rect 534 33203 541 33251
rect 534 33110 538 33203
rect 558 33110 562 33660
rect 582 33110 586 33660
rect 606 33110 610 33660
rect 630 33110 634 33660
rect 654 33231 658 33660
rect 643 33230 677 33231
rect 678 33230 682 33660
rect 702 33230 706 33660
rect 726 33230 730 33660
rect 750 33230 754 33660
rect 774 33230 778 33660
rect 798 33230 802 33660
rect 822 33230 826 33660
rect 846 33230 850 33660
rect 870 33230 874 33660
rect 894 33230 898 33660
rect 918 33230 922 33660
rect 942 33230 946 33660
rect 966 33230 970 33660
rect 990 33230 994 33660
rect 1014 33230 1018 33660
rect 1038 33230 1042 33660
rect 1045 33659 1059 33660
rect 1062 33659 1069 33683
rect 1062 33230 1066 33659
rect 1086 33230 1090 33876
rect 1099 33389 1104 33399
rect 1110 33389 1114 33876
rect 1109 33375 1114 33389
rect 1110 33230 1114 33375
rect 1134 33323 1138 33876
rect 1134 33299 1141 33323
rect 1134 33230 1138 33299
rect 1158 33230 1162 33876
rect 1182 33230 1186 33876
rect 1206 33230 1210 33876
rect 1219 33869 1224 33876
rect 1230 33869 1234 33876
rect 1229 33855 1234 33869
rect 1230 33615 1234 33855
rect 1254 33803 1258 33972
rect 1254 33779 1261 33803
rect 1219 33614 1253 33615
rect 1254 33614 1258 33779
rect 1278 33614 1282 33972
rect 1302 33614 1306 33972
rect 1326 33614 1330 33972
rect 1350 33614 1354 33972
rect 1374 33614 1378 33972
rect 1387 33893 1392 33903
rect 1398 33893 1402 33972
rect 1397 33879 1402 33893
rect 1398 33614 1402 33879
rect 1422 33827 1426 33972
rect 1422 33803 1429 33827
rect 1422 33614 1426 33803
rect 1446 33614 1450 33972
rect 1470 33614 1474 33972
rect 1494 33614 1498 33972
rect 1518 33614 1522 33972
rect 1542 33735 1546 33972
rect 1531 33734 1565 33735
rect 1566 33734 1570 33972
rect 1590 33734 1594 33972
rect 1597 33971 1611 33972
rect 1603 33965 1608 33971
rect 1613 33951 1618 33965
rect 1614 33734 1618 33951
rect 1627 33821 1632 33831
rect 1637 33807 1642 33821
rect 1638 33734 1642 33807
rect 1651 33734 1659 33735
rect 1531 33732 1659 33734
rect 1531 33725 1536 33732
rect 1542 33725 1546 33732
rect 1541 33711 1546 33725
rect 1531 33701 1536 33711
rect 1541 33687 1546 33701
rect 1542 33614 1546 33687
rect 1566 33659 1570 33732
rect 1219 33612 1563 33614
rect 1219 33605 1224 33612
rect 1230 33605 1234 33612
rect 1229 33591 1234 33605
rect 1219 33581 1224 33591
rect 1229 33567 1234 33581
rect 1230 33230 1234 33567
rect 1254 33539 1258 33612
rect 1254 33491 1261 33539
rect 1254 33230 1258 33491
rect 1278 33230 1282 33612
rect 1302 33230 1306 33612
rect 1326 33230 1330 33612
rect 1350 33230 1354 33612
rect 1374 33230 1378 33612
rect 1398 33230 1402 33612
rect 1422 33230 1426 33612
rect 1446 33230 1450 33612
rect 1470 33230 1474 33612
rect 1494 33230 1498 33612
rect 1518 33230 1522 33612
rect 1542 33230 1546 33612
rect 1549 33611 1563 33612
rect 1566 33611 1573 33659
rect 1566 33230 1570 33611
rect 1590 33230 1594 33732
rect 1614 33230 1618 33732
rect 1638 33230 1642 33732
rect 1645 33731 1659 33732
rect 1651 33725 1656 33731
rect 1661 33711 1666 33725
rect 1651 33653 1656 33663
rect 1662 33653 1666 33711
rect 1661 33639 1666 33653
rect 1675 33649 1683 33653
rect 1669 33639 1675 33649
rect 1651 33605 1656 33615
rect 1661 33591 1666 33605
rect 1662 33230 1666 33591
rect 1675 33437 1680 33447
rect 1685 33423 1690 33437
rect 1675 33245 1680 33255
rect 1686 33245 1690 33423
rect 1699 33317 1704 33327
rect 1709 33303 1714 33317
rect 1699 33269 1704 33279
rect 1710 33269 1714 33303
rect 1709 33255 1714 33269
rect 1685 33231 1690 33245
rect 1675 33230 1709 33231
rect 643 33228 1709 33230
rect 643 33221 648 33228
rect 654 33221 658 33228
rect 653 33207 658 33221
rect 643 33197 648 33207
rect 653 33183 658 33197
rect 654 33110 658 33183
rect 678 33155 682 33228
rect -2393 33108 675 33110
rect -2371 33086 -2366 33108
rect -2348 33086 -2343 33108
rect -2325 33086 -2320 33108
rect -2072 33106 -2036 33107
rect -2072 33100 -2054 33106
rect -2309 33092 -2301 33100
rect -2317 33086 -2309 33092
rect -2092 33091 -2062 33096
rect -2000 33087 -1992 33108
rect -1938 33107 -1906 33108
rect -1920 33106 -1906 33107
rect -1806 33100 -1680 33106
rect -1854 33091 -1806 33096
rect -1655 33092 -1647 33100
rect -1982 33087 -1966 33088
rect -2000 33086 -1966 33087
rect -1846 33086 -1806 33089
rect -1663 33086 -1655 33092
rect -1642 33086 -1637 33108
rect -1619 33086 -1614 33108
rect -1530 33086 -1526 33108
rect -1506 33086 -1502 33108
rect -1482 33086 -1478 33108
rect -1458 33086 -1454 33108
rect -1434 33086 -1430 33108
rect -1410 33086 -1406 33108
rect -1386 33086 -1382 33108
rect -1362 33086 -1358 33108
rect -1338 33086 -1334 33108
rect -1314 33086 -1310 33108
rect -1290 33086 -1286 33108
rect -1266 33086 -1262 33108
rect -1242 33086 -1238 33108
rect -1218 33086 -1214 33108
rect -1194 33086 -1190 33108
rect -1170 33086 -1166 33108
rect -1146 33086 -1142 33108
rect -1122 33086 -1118 33108
rect -1098 33086 -1094 33108
rect -1074 33107 -1070 33108
rect -2393 33084 -1077 33086
rect -2371 33062 -2366 33084
rect -2348 33062 -2343 33084
rect -2325 33062 -2320 33084
rect -2000 33082 -1966 33084
rect -2309 33064 -2301 33072
rect -2062 33071 -2054 33078
rect -2092 33064 -2084 33071
rect -2062 33064 -2026 33066
rect -2317 33062 -2309 33064
rect -2062 33062 -2012 33064
rect -2000 33062 -1992 33082
rect -1982 33081 -1966 33082
rect -1846 33080 -1806 33084
rect -1846 33073 -1798 33078
rect -1806 33071 -1798 33073
rect -1854 33069 -1846 33071
rect -1854 33064 -1806 33069
rect -1655 33064 -1647 33072
rect -1864 33062 -1796 33063
rect -1663 33062 -1655 33064
rect -1642 33062 -1637 33084
rect -1619 33062 -1614 33084
rect -1530 33062 -1526 33084
rect -1506 33062 -1502 33084
rect -1482 33062 -1478 33084
rect -1458 33062 -1454 33084
rect -1434 33062 -1430 33084
rect -1410 33062 -1406 33084
rect -1386 33062 -1382 33084
rect -1362 33062 -1358 33084
rect -1338 33062 -1334 33084
rect -1314 33062 -1310 33084
rect -1290 33062 -1286 33084
rect -1266 33062 -1262 33084
rect -1242 33062 -1238 33084
rect -1218 33062 -1214 33084
rect -1194 33062 -1190 33084
rect -1170 33062 -1166 33084
rect -1146 33062 -1142 33084
rect -1122 33062 -1118 33084
rect -1098 33062 -1094 33084
rect -1091 33083 -1077 33084
rect -1074 33083 -1067 33107
rect -1074 33062 -1070 33083
rect -1050 33062 -1046 33108
rect -1026 33062 -1022 33108
rect -1002 33062 -998 33108
rect -978 33062 -974 33108
rect -954 33062 -950 33108
rect -930 33062 -926 33108
rect -906 33062 -902 33108
rect -882 33062 -878 33108
rect -858 33062 -854 33108
rect -834 33062 -830 33108
rect -810 33062 -806 33108
rect -786 33062 -782 33108
rect -762 33062 -758 33108
rect -738 33062 -734 33108
rect -714 33062 -710 33108
rect -690 33062 -686 33108
rect -666 33062 -662 33108
rect -642 33062 -638 33108
rect -618 33062 -614 33108
rect -594 33062 -590 33108
rect -570 33062 -566 33108
rect -546 33062 -542 33108
rect -522 33062 -518 33108
rect -498 33062 -494 33108
rect -474 33062 -470 33108
rect -450 33062 -446 33108
rect -426 33062 -422 33108
rect -402 33062 -398 33108
rect -378 33062 -374 33108
rect -354 33062 -350 33108
rect -330 33062 -326 33108
rect -306 33062 -302 33108
rect -282 33062 -278 33108
rect -258 33062 -254 33108
rect -245 33077 -240 33087
rect -234 33077 -230 33108
rect -235 33063 -230 33077
rect -234 33062 -230 33063
rect -210 33062 -206 33108
rect -186 33062 -182 33108
rect -162 33062 -158 33108
rect -138 33062 -134 33108
rect -114 33062 -110 33108
rect -90 33062 -86 33108
rect -66 33062 -62 33108
rect -42 33062 -38 33108
rect -18 33062 -14 33108
rect 6 33062 10 33108
rect 30 33062 34 33108
rect 54 33062 58 33108
rect 78 33062 82 33108
rect 102 33062 106 33108
rect 126 33062 130 33108
rect 150 33083 154 33108
rect -2393 33060 147 33062
rect -2371 32990 -2366 33060
rect -2348 32990 -2343 33060
rect -2325 32990 -2320 33060
rect -2317 33056 -2309 33060
rect -2062 33056 -2054 33060
rect -2154 33052 -2138 33054
rect -2057 33052 -2054 33056
rect -2292 33046 -2054 33052
rect -2052 33046 -2044 33056
rect -2092 33030 -2062 33032
rect -2094 33026 -2062 33030
rect -2309 32996 -2301 33002
rect -2317 32990 -2309 32996
rect -2000 32990 -1992 33060
rect -1846 33053 -1806 33060
rect -1663 33056 -1655 33060
rect -1846 33046 -1680 33052
rect -1854 33030 -1806 33032
rect -1854 33026 -1680 33030
rect -1655 32996 -1647 33002
rect -1663 32990 -1655 32996
rect -1642 32990 -1637 33060
rect -1619 32990 -1614 33060
rect -1530 32990 -1526 33060
rect -1506 32990 -1502 33060
rect -1482 32990 -1478 33060
rect -1458 32990 -1454 33060
rect -1434 32990 -1430 33060
rect -1410 32990 -1406 33060
rect -1386 32990 -1382 33060
rect -1362 32990 -1358 33060
rect -1338 32990 -1334 33060
rect -1314 32990 -1310 33060
rect -1290 32990 -1286 33060
rect -1266 32990 -1262 33060
rect -1242 32990 -1238 33060
rect -1218 32990 -1214 33060
rect -1194 32990 -1190 33060
rect -1170 32990 -1166 33060
rect -1146 32990 -1142 33060
rect -1122 32990 -1118 33060
rect -1098 32990 -1094 33060
rect -1074 32990 -1070 33060
rect -1050 32990 -1046 33060
rect -1026 32990 -1022 33060
rect -1002 32990 -998 33060
rect -978 32990 -974 33060
rect -954 32990 -950 33060
rect -930 32990 -926 33060
rect -906 32990 -902 33060
rect -882 32990 -878 33060
rect -858 32990 -854 33060
rect -834 32990 -830 33060
rect -810 32990 -806 33060
rect -786 32990 -782 33060
rect -762 32990 -758 33060
rect -738 32990 -734 33060
rect -714 32990 -710 33060
rect -690 32990 -686 33060
rect -666 32990 -662 33060
rect -642 32990 -638 33060
rect -618 32990 -614 33060
rect -594 32990 -590 33060
rect -570 32990 -566 33060
rect -546 32990 -542 33060
rect -522 32990 -518 33060
rect -498 32990 -494 33060
rect -474 32990 -470 33060
rect -450 32990 -446 33060
rect -426 32990 -422 33060
rect -402 33015 -398 33060
rect -413 33014 -379 33015
rect -378 33014 -374 33060
rect -354 33014 -350 33060
rect -330 33014 -326 33060
rect -306 33014 -302 33060
rect -282 33014 -278 33060
rect -258 33014 -254 33060
rect -234 33014 -230 33060
rect -210 33014 -206 33060
rect -186 33014 -182 33060
rect -162 33014 -158 33060
rect -138 33014 -134 33060
rect -114 33014 -110 33060
rect -90 33014 -86 33060
rect -66 33014 -62 33060
rect -42 33014 -38 33060
rect -18 33014 -14 33060
rect 6 33014 10 33060
rect 30 33014 34 33060
rect 54 33014 58 33060
rect 78 33014 82 33060
rect 102 33014 106 33060
rect 126 33014 130 33060
rect 133 33059 147 33060
rect 150 33059 157 33083
rect 150 33014 154 33059
rect 174 33014 178 33108
rect 198 33014 202 33108
rect 222 33014 226 33108
rect 246 33014 250 33108
rect 270 33014 274 33108
rect 294 33014 298 33108
rect 318 33014 322 33108
rect 342 33014 346 33108
rect 366 33014 370 33108
rect 390 33014 394 33108
rect 414 33014 418 33108
rect 438 33014 442 33108
rect 462 33014 466 33108
rect 486 33014 490 33108
rect 510 33014 514 33108
rect 534 33014 538 33108
rect 558 33014 562 33108
rect 582 33014 586 33108
rect 606 33014 610 33108
rect 630 33014 634 33108
rect 654 33014 658 33108
rect 661 33107 675 33108
rect 678 33107 685 33155
rect 678 33014 682 33107
rect 702 33014 706 33228
rect 726 33014 730 33228
rect 750 33014 754 33228
rect 774 33014 778 33228
rect 798 33014 802 33228
rect 822 33014 826 33228
rect 846 33014 850 33228
rect 870 33014 874 33228
rect 894 33014 898 33228
rect 918 33014 922 33228
rect 942 33014 946 33228
rect 966 33014 970 33228
rect 979 33053 984 33063
rect 990 33053 994 33228
rect 989 33039 994 33053
rect 990 33014 994 33039
rect 1014 33014 1018 33228
rect 1038 33014 1042 33228
rect 1062 33014 1066 33228
rect 1086 33014 1090 33228
rect 1110 33014 1114 33228
rect 1134 33014 1138 33228
rect 1158 33135 1162 33228
rect 1147 33134 1181 33135
rect 1182 33134 1186 33228
rect 1206 33134 1210 33228
rect 1230 33134 1234 33228
rect 1254 33134 1258 33228
rect 1278 33134 1282 33228
rect 1302 33134 1306 33228
rect 1326 33134 1330 33228
rect 1350 33134 1354 33228
rect 1374 33134 1378 33228
rect 1398 33134 1402 33228
rect 1422 33134 1426 33228
rect 1446 33134 1450 33228
rect 1470 33134 1474 33228
rect 1494 33134 1498 33228
rect 1518 33134 1522 33228
rect 1542 33134 1546 33228
rect 1566 33134 1570 33228
rect 1590 33134 1594 33228
rect 1614 33134 1618 33228
rect 1638 33134 1642 33228
rect 1662 33134 1666 33228
rect 1675 33221 1680 33228
rect 1685 33207 1690 33221
rect 1686 33134 1690 33207
rect 1699 33134 1707 33135
rect 1147 33132 1707 33134
rect 1147 33125 1152 33132
rect 1158 33125 1162 33132
rect 1157 33111 1162 33125
rect 1147 33101 1152 33111
rect 1157 33087 1162 33101
rect 1158 33014 1162 33087
rect 1182 33059 1186 33132
rect -413 33012 1179 33014
rect -413 33005 -408 33012
rect -402 33005 -398 33012
rect -403 32991 -398 33005
rect -413 32990 -379 32991
rect -2393 32988 -379 32990
rect -2371 32894 -2366 32988
rect -2348 32894 -2343 32988
rect -2325 32926 -2320 32988
rect -2317 32986 -2309 32988
rect -2000 32987 -1966 32988
rect -2000 32986 -1982 32987
rect -1663 32986 -1655 32988
rect -2028 32978 -2018 32980
rect -2309 32968 -2301 32974
rect -2091 32968 -2061 32975
rect -2317 32958 -2309 32968
rect -2044 32966 -2028 32968
rect -2026 32966 -2014 32978
rect -2084 32960 -2061 32966
rect -2044 32964 -2014 32966
rect -2292 32950 -2054 32959
rect -2325 32918 -2317 32926
rect -2325 32898 -2320 32918
rect -2317 32910 -2309 32918
rect -2325 32894 -2317 32898
rect -2000 32894 -1992 32986
rect -1982 32985 -1966 32986
rect -1980 32968 -1932 32975
rect -1655 32968 -1647 32974
rect -1846 32950 -1680 32959
rect -1663 32958 -1655 32968
rect -1671 32918 -1663 32926
rect -1663 32910 -1655 32918
rect -1671 32894 -1663 32898
rect -1642 32894 -1637 32988
rect -1619 32894 -1614 32988
rect -1530 32894 -1526 32988
rect -1506 32894 -1502 32988
rect -1482 32894 -1478 32988
rect -1458 32894 -1454 32988
rect -1434 32894 -1430 32988
rect -1410 32894 -1406 32988
rect -1386 32894 -1382 32988
rect -1362 32894 -1358 32988
rect -1338 32894 -1334 32988
rect -1314 32894 -1310 32988
rect -1290 32894 -1286 32988
rect -1266 32894 -1262 32988
rect -1242 32894 -1238 32988
rect -1218 32894 -1214 32988
rect -1194 32894 -1190 32988
rect -1170 32894 -1166 32988
rect -1146 32894 -1142 32988
rect -1122 32894 -1118 32988
rect -1098 32894 -1094 32988
rect -1074 32894 -1070 32988
rect -1050 32894 -1046 32988
rect -1026 32894 -1022 32988
rect -1002 32894 -998 32988
rect -978 32894 -974 32988
rect -954 32894 -950 32988
rect -930 32894 -926 32988
rect -906 32894 -902 32988
rect -882 32894 -878 32988
rect -858 32894 -854 32988
rect -834 32894 -830 32988
rect -810 32894 -806 32988
rect -786 32894 -782 32988
rect -762 32894 -758 32988
rect -738 32894 -734 32988
rect -714 32894 -710 32988
rect -690 32894 -686 32988
rect -666 32894 -662 32988
rect -642 32894 -638 32988
rect -618 32894 -614 32988
rect -594 32894 -590 32988
rect -570 32894 -566 32988
rect -546 32894 -542 32988
rect -522 32894 -518 32988
rect -498 32894 -494 32988
rect -474 32894 -470 32988
rect -450 32894 -446 32988
rect -426 32894 -422 32988
rect -413 32981 -408 32988
rect -403 32967 -398 32981
rect -402 32894 -398 32967
rect -378 32939 -374 33012
rect -2393 32892 -381 32894
rect -2371 32846 -2366 32892
rect -2348 32846 -2343 32892
rect -2325 32884 -2317 32892
rect -2018 32891 -2004 32892
rect -2000 32891 -1992 32892
rect -2072 32890 -1928 32891
rect -2072 32884 -2053 32890
rect -2325 32868 -2320 32884
rect -2317 32882 -2309 32884
rect -2309 32870 -2301 32882
rect -2092 32875 -2062 32880
rect -2317 32868 -2309 32870
rect -2325 32856 -2317 32868
rect -2098 32862 -2096 32873
rect -2092 32862 -2084 32875
rect -2000 32874 -1992 32890
rect -1972 32884 -1928 32890
rect -1924 32884 -1918 32892
rect -1671 32884 -1663 32892
rect -1663 32882 -1655 32884
rect -2083 32864 -2062 32873
rect -2027 32872 -1992 32874
rect -2018 32864 -2002 32872
rect -2000 32864 -1992 32872
rect -2100 32857 -2096 32862
rect -2083 32857 -2053 32862
rect -2003 32860 -1990 32864
rect -1972 32862 -1964 32871
rect -1928 32870 -1924 32873
rect -1655 32870 -1647 32882
rect -1663 32868 -1655 32870
rect -2325 32846 -2320 32856
rect -2317 32854 -2309 32856
rect -2309 32846 -2301 32854
rect -2004 32850 -2003 32860
rect -2062 32846 -2012 32848
rect -2000 32846 -1992 32860
rect -1972 32857 -1924 32862
rect -1864 32857 -1796 32863
rect -1671 32856 -1663 32868
rect -1663 32854 -1655 32856
rect -1864 32846 -1796 32847
rect -1655 32846 -1647 32854
rect -1642 32846 -1637 32892
rect -1619 32846 -1614 32892
rect -1530 32846 -1526 32892
rect -1506 32846 -1502 32892
rect -1482 32846 -1478 32892
rect -1458 32846 -1454 32892
rect -1434 32846 -1430 32892
rect -1410 32846 -1406 32892
rect -1386 32846 -1382 32892
rect -1362 32846 -1358 32892
rect -1338 32846 -1334 32892
rect -1314 32846 -1310 32892
rect -1290 32846 -1286 32892
rect -1266 32846 -1262 32892
rect -1242 32846 -1238 32892
rect -1218 32846 -1214 32892
rect -1194 32846 -1190 32892
rect -1170 32846 -1166 32892
rect -1146 32846 -1142 32892
rect -1122 32846 -1118 32892
rect -1098 32846 -1094 32892
rect -1074 32846 -1070 32892
rect -1050 32846 -1046 32892
rect -1026 32846 -1022 32892
rect -1002 32846 -998 32892
rect -978 32846 -974 32892
rect -954 32846 -950 32892
rect -930 32846 -926 32892
rect -906 32846 -902 32892
rect -882 32846 -878 32892
rect -858 32846 -854 32892
rect -834 32846 -830 32892
rect -810 32846 -806 32892
rect -786 32846 -782 32892
rect -762 32846 -758 32892
rect -738 32846 -734 32892
rect -714 32846 -710 32892
rect -690 32846 -686 32892
rect -666 32846 -662 32892
rect -642 32846 -638 32892
rect -618 32846 -614 32892
rect -594 32846 -590 32892
rect -570 32846 -566 32892
rect -546 32846 -542 32892
rect -522 32846 -518 32892
rect -498 32846 -494 32892
rect -474 32846 -470 32892
rect -450 32846 -446 32892
rect -426 32846 -422 32892
rect -402 32846 -398 32892
rect -395 32891 -381 32892
rect -378 32891 -371 32939
rect -378 32846 -374 32891
rect -354 32846 -350 33012
rect -330 32846 -326 33012
rect -306 32846 -302 33012
rect -282 32846 -278 33012
rect -258 32846 -254 33012
rect -234 32846 -230 33012
rect -210 33011 -206 33012
rect -210 32987 -203 33011
rect -210 32846 -206 32987
rect -186 32846 -182 33012
rect -162 32846 -158 33012
rect -138 32846 -134 33012
rect -114 32919 -110 33012
rect -125 32918 -91 32919
rect -90 32918 -86 33012
rect -66 32918 -62 33012
rect -42 32918 -38 33012
rect -18 32918 -14 33012
rect 6 32918 10 33012
rect 30 32918 34 33012
rect 54 32918 58 33012
rect 78 32918 82 33012
rect 102 32918 106 33012
rect 126 32918 130 33012
rect 150 32918 154 33012
rect 174 32918 178 33012
rect 198 32918 202 33012
rect 222 32918 226 33012
rect 246 32918 250 33012
rect 270 32918 274 33012
rect 294 32918 298 33012
rect 318 32918 322 33012
rect 342 32918 346 33012
rect 366 32918 370 33012
rect 390 32918 394 33012
rect 414 32918 418 33012
rect 438 32918 442 33012
rect 462 32918 466 33012
rect 486 32918 490 33012
rect 510 32918 514 33012
rect 534 32918 538 33012
rect 558 32918 562 33012
rect 582 32918 586 33012
rect 606 32918 610 33012
rect 630 32918 634 33012
rect 654 32918 658 33012
rect 678 32918 682 33012
rect 702 32918 706 33012
rect 726 32918 730 33012
rect 750 32918 754 33012
rect 774 32918 778 33012
rect 798 32918 802 33012
rect 822 32918 826 33012
rect 846 32918 850 33012
rect 870 32918 874 33012
rect 894 32918 898 33012
rect 918 32918 922 33012
rect 942 32918 946 33012
rect 966 32918 970 33012
rect 990 32918 994 33012
rect 1014 32987 1018 33012
rect 1014 32963 1021 32987
rect 1014 32918 1018 32963
rect 1038 32918 1042 33012
rect 1062 32918 1066 33012
rect 1086 32918 1090 33012
rect 1110 32918 1114 33012
rect 1134 32918 1138 33012
rect 1147 32933 1152 32943
rect 1158 32933 1162 33012
rect 1165 33011 1179 33012
rect 1182 33011 1189 33059
rect 1157 32919 1162 32933
rect 1158 32918 1162 32919
rect 1182 32918 1186 33011
rect 1206 32918 1210 33132
rect 1230 32918 1234 33132
rect 1254 32918 1258 33132
rect 1278 32918 1282 33132
rect 1302 32918 1306 33132
rect 1326 32918 1330 33132
rect 1350 32918 1354 33132
rect 1374 32918 1378 33132
rect 1398 32918 1402 33132
rect 1422 32918 1426 33132
rect 1446 32918 1450 33132
rect 1470 32918 1474 33132
rect 1494 32918 1498 33132
rect 1518 32918 1522 33132
rect 1542 32918 1546 33132
rect 1566 32918 1570 33132
rect 1590 32918 1594 33132
rect 1614 32918 1618 33132
rect 1638 32918 1642 33132
rect 1662 32918 1666 33132
rect 1686 32918 1690 33132
rect 1693 33131 1707 33132
rect 1699 33125 1704 33131
rect 1709 33111 1714 33125
rect 1710 32918 1714 33111
rect 1723 33005 1728 33015
rect 1733 32991 1738 33005
rect 1734 32918 1738 32991
rect 1747 32918 1755 32919
rect -125 32916 1755 32918
rect -125 32909 -120 32916
rect -114 32909 -110 32916
rect -115 32895 -110 32909
rect -125 32885 -120 32895
rect -115 32871 -110 32885
rect -114 32846 -110 32871
rect -90 32847 -86 32916
rect -101 32846 -67 32847
rect -2393 32844 -67 32846
rect -2371 32798 -2366 32844
rect -2348 32798 -2343 32844
rect -2325 32840 -2320 32844
rect -2309 32842 -2301 32844
rect -2317 32840 -2309 32842
rect -2325 32828 -2317 32840
rect -2325 32798 -2320 32828
rect -2317 32826 -2309 32828
rect -2092 32814 -2062 32816
rect -2094 32810 -2062 32814
rect -2000 32798 -1992 32844
rect -1655 32842 -1647 32844
rect -1663 32840 -1655 32842
rect -1671 32828 -1663 32840
rect -1663 32826 -1655 32828
rect -1854 32814 -1806 32816
rect -1854 32810 -1680 32814
rect -1642 32798 -1637 32844
rect -1619 32798 -1614 32844
rect -1530 32798 -1526 32844
rect -1506 32798 -1502 32844
rect -1482 32798 -1478 32844
rect -1458 32798 -1454 32844
rect -1434 32798 -1430 32844
rect -1410 32798 -1406 32844
rect -1386 32798 -1382 32844
rect -1362 32798 -1358 32844
rect -1338 32798 -1334 32844
rect -1314 32798 -1310 32844
rect -1290 32798 -1286 32844
rect -1266 32798 -1262 32844
rect -1242 32798 -1238 32844
rect -1218 32798 -1214 32844
rect -1194 32798 -1190 32844
rect -1170 32798 -1166 32844
rect -1146 32798 -1142 32844
rect -1122 32798 -1118 32844
rect -1098 32798 -1094 32844
rect -1074 32798 -1070 32844
rect -1050 32798 -1046 32844
rect -1026 32798 -1022 32844
rect -1002 32798 -998 32844
rect -978 32798 -974 32844
rect -954 32798 -950 32844
rect -930 32798 -926 32844
rect -906 32798 -902 32844
rect -882 32798 -878 32844
rect -858 32798 -854 32844
rect -834 32798 -830 32844
rect -810 32798 -806 32844
rect -786 32798 -782 32844
rect -762 32798 -758 32844
rect -738 32798 -734 32844
rect -714 32798 -710 32844
rect -690 32798 -686 32844
rect -666 32798 -662 32844
rect -642 32798 -638 32844
rect -618 32798 -614 32844
rect -594 32798 -590 32844
rect -570 32798 -566 32844
rect -546 32798 -542 32844
rect -522 32798 -518 32844
rect -498 32798 -494 32844
rect -474 32798 -470 32844
rect -450 32798 -446 32844
rect -426 32798 -422 32844
rect -402 32798 -398 32844
rect -378 32798 -374 32844
rect -354 32798 -350 32844
rect -330 32798 -326 32844
rect -306 32798 -302 32844
rect -282 32798 -278 32844
rect -258 32798 -254 32844
rect -234 32798 -230 32844
rect -210 32798 -206 32844
rect -186 32798 -182 32844
rect -162 32798 -158 32844
rect -138 32798 -134 32844
rect -114 32798 -110 32844
rect -101 32837 -96 32844
rect -90 32843 -86 32844
rect -90 32837 -83 32843
rect -91 32823 -83 32837
rect -2393 32796 -93 32798
rect -2371 32774 -2366 32796
rect -2348 32774 -2343 32796
rect -2325 32774 -2320 32796
rect -2072 32794 -2036 32795
rect -2072 32788 -2054 32794
rect -2309 32780 -2301 32788
rect -2317 32774 -2309 32780
rect -2092 32779 -2062 32784
rect -2000 32775 -1992 32796
rect -1938 32795 -1906 32796
rect -1920 32794 -1906 32795
rect -1806 32788 -1680 32794
rect -1854 32779 -1806 32784
rect -1655 32780 -1647 32788
rect -1982 32775 -1966 32776
rect -2000 32774 -1966 32775
rect -1846 32774 -1806 32777
rect -1663 32774 -1655 32780
rect -1642 32774 -1637 32796
rect -1619 32774 -1614 32796
rect -1530 32774 -1526 32796
rect -1506 32774 -1502 32796
rect -1482 32774 -1478 32796
rect -1458 32774 -1454 32796
rect -1434 32774 -1430 32796
rect -1410 32774 -1406 32796
rect -1386 32774 -1382 32796
rect -1362 32774 -1358 32796
rect -1338 32774 -1334 32796
rect -1314 32774 -1310 32796
rect -1290 32774 -1286 32796
rect -1266 32774 -1262 32796
rect -1242 32774 -1238 32796
rect -1218 32774 -1214 32796
rect -1194 32774 -1190 32796
rect -1170 32774 -1166 32796
rect -1146 32774 -1142 32796
rect -1122 32774 -1118 32796
rect -1098 32774 -1094 32796
rect -1074 32774 -1070 32796
rect -1050 32774 -1046 32796
rect -1026 32774 -1022 32796
rect -1002 32774 -998 32796
rect -978 32774 -974 32796
rect -954 32774 -950 32796
rect -930 32774 -926 32796
rect -906 32774 -902 32796
rect -882 32774 -878 32796
rect -858 32774 -854 32796
rect -834 32774 -830 32796
rect -810 32774 -806 32796
rect -786 32774 -782 32796
rect -762 32774 -758 32796
rect -738 32774 -734 32796
rect -714 32774 -710 32796
rect -690 32774 -686 32796
rect -666 32774 -662 32796
rect -642 32774 -638 32796
rect -618 32774 -614 32796
rect -594 32774 -590 32796
rect -570 32774 -566 32796
rect -546 32774 -542 32796
rect -522 32774 -518 32796
rect -498 32774 -494 32796
rect -474 32774 -470 32796
rect -450 32774 -446 32796
rect -426 32774 -422 32796
rect -402 32774 -398 32796
rect -378 32774 -374 32796
rect -354 32774 -350 32796
rect -330 32774 -326 32796
rect -306 32774 -302 32796
rect -282 32774 -278 32796
rect -258 32774 -254 32796
rect -234 32774 -230 32796
rect -210 32774 -206 32796
rect -186 32774 -182 32796
rect -162 32774 -158 32796
rect -138 32774 -134 32796
rect -114 32774 -110 32796
rect -107 32795 -93 32796
rect -90 32795 -83 32823
rect -90 32774 -86 32795
rect -66 32774 -62 32916
rect -42 32774 -38 32916
rect -18 32774 -14 32916
rect 6 32774 10 32916
rect 30 32774 34 32916
rect 54 32774 58 32916
rect 78 32774 82 32916
rect 102 32774 106 32916
rect 126 32774 130 32916
rect 150 32774 154 32916
rect 174 32774 178 32916
rect 198 32774 202 32916
rect 222 32774 226 32916
rect 246 32774 250 32916
rect 270 32774 274 32916
rect 294 32774 298 32916
rect 318 32774 322 32916
rect 342 32774 346 32916
rect 366 32774 370 32916
rect 390 32774 394 32916
rect 414 32774 418 32916
rect 438 32774 442 32916
rect 462 32774 466 32916
rect 486 32774 490 32916
rect 510 32774 514 32916
rect 534 32774 538 32916
rect 558 32774 562 32916
rect 582 32774 586 32916
rect 606 32774 610 32916
rect 630 32774 634 32916
rect 654 32774 658 32916
rect 678 32774 682 32916
rect 702 32774 706 32916
rect 726 32774 730 32916
rect 750 32774 754 32916
rect 774 32774 778 32916
rect 798 32774 802 32916
rect 822 32774 826 32916
rect 846 32774 850 32916
rect 870 32774 874 32916
rect 894 32774 898 32916
rect 918 32774 922 32916
rect 942 32774 946 32916
rect 966 32774 970 32916
rect 990 32774 994 32916
rect 1014 32774 1018 32916
rect 1038 32774 1042 32916
rect 1062 32774 1066 32916
rect 1086 32774 1090 32916
rect 1110 32774 1114 32916
rect 1134 32774 1138 32916
rect 1158 32774 1162 32916
rect 1182 32867 1186 32916
rect 1182 32843 1189 32867
rect 1182 32774 1186 32843
rect 1206 32774 1210 32916
rect 1230 32774 1234 32916
rect 1254 32823 1258 32916
rect 1243 32822 1277 32823
rect 1278 32822 1282 32916
rect 1302 32822 1306 32916
rect 1326 32822 1330 32916
rect 1350 32822 1354 32916
rect 1374 32822 1378 32916
rect 1398 32822 1402 32916
rect 1422 32822 1426 32916
rect 1446 32822 1450 32916
rect 1470 32822 1474 32916
rect 1494 32822 1498 32916
rect 1518 32822 1522 32916
rect 1542 32822 1546 32916
rect 1566 32822 1570 32916
rect 1590 32822 1594 32916
rect 1614 32822 1618 32916
rect 1638 32822 1642 32916
rect 1662 32822 1666 32916
rect 1686 32822 1690 32916
rect 1710 32822 1714 32916
rect 1734 32822 1738 32916
rect 1741 32915 1755 32916
rect 1747 32909 1752 32915
rect 1757 32895 1762 32909
rect 1747 32861 1752 32871
rect 1758 32861 1762 32895
rect 1757 32847 1762 32861
rect 1747 32822 1779 32823
rect 1243 32820 1779 32822
rect 1243 32813 1248 32820
rect 1254 32813 1258 32820
rect 1253 32799 1258 32813
rect 1243 32789 1248 32799
rect 1253 32775 1258 32789
rect 1254 32774 1258 32775
rect 1278 32774 1282 32820
rect 1302 32774 1306 32820
rect 1326 32775 1330 32820
rect 1315 32774 1349 32775
rect -2393 32772 1349 32774
rect -2371 32750 -2366 32772
rect -2348 32750 -2343 32772
rect -2325 32750 -2320 32772
rect -2000 32770 -1966 32772
rect -2309 32752 -2301 32760
rect -2062 32759 -2054 32766
rect -2092 32752 -2084 32759
rect -2062 32752 -2026 32754
rect -2317 32750 -2309 32752
rect -2062 32750 -2012 32752
rect -2000 32750 -1992 32770
rect -1982 32769 -1966 32770
rect -1846 32768 -1806 32772
rect -1846 32761 -1798 32766
rect -1806 32759 -1798 32761
rect -1854 32757 -1846 32759
rect -1854 32752 -1806 32757
rect -1655 32752 -1647 32760
rect -1864 32750 -1796 32751
rect -1663 32750 -1655 32752
rect -1642 32750 -1637 32772
rect -1619 32750 -1614 32772
rect -1530 32750 -1526 32772
rect -1506 32750 -1502 32772
rect -1482 32750 -1478 32772
rect -1458 32750 -1454 32772
rect -1434 32750 -1430 32772
rect -1410 32750 -1406 32772
rect -1386 32750 -1382 32772
rect -1362 32750 -1358 32772
rect -1338 32750 -1334 32772
rect -1314 32750 -1310 32772
rect -1290 32750 -1286 32772
rect -1266 32750 -1262 32772
rect -1242 32750 -1238 32772
rect -1218 32750 -1214 32772
rect -1194 32750 -1190 32772
rect -1170 32750 -1166 32772
rect -1146 32750 -1142 32772
rect -1122 32750 -1118 32772
rect -1098 32750 -1094 32772
rect -1074 32750 -1070 32772
rect -1050 32750 -1046 32772
rect -1026 32750 -1022 32772
rect -1002 32750 -998 32772
rect -978 32750 -974 32772
rect -954 32750 -950 32772
rect -930 32750 -926 32772
rect -906 32750 -902 32772
rect -882 32750 -878 32772
rect -858 32750 -854 32772
rect -834 32750 -830 32772
rect -810 32750 -806 32772
rect -786 32750 -782 32772
rect -762 32750 -758 32772
rect -738 32750 -734 32772
rect -714 32750 -710 32772
rect -690 32750 -686 32772
rect -666 32750 -662 32772
rect -642 32750 -638 32772
rect -618 32750 -614 32772
rect -594 32750 -590 32772
rect -570 32750 -566 32772
rect -546 32750 -542 32772
rect -522 32750 -518 32772
rect -498 32750 -494 32772
rect -474 32750 -470 32772
rect -450 32750 -446 32772
rect -426 32750 -422 32772
rect -402 32750 -398 32772
rect -378 32750 -374 32772
rect -354 32750 -350 32772
rect -330 32750 -326 32772
rect -306 32750 -302 32772
rect -282 32750 -278 32772
rect -258 32750 -254 32772
rect -234 32750 -230 32772
rect -210 32750 -206 32772
rect -186 32750 -182 32772
rect -162 32750 -158 32772
rect -138 32750 -134 32772
rect -114 32750 -110 32772
rect -90 32750 -86 32772
rect -66 32771 -62 32772
rect -2393 32748 -69 32750
rect -2371 32702 -2366 32748
rect -2348 32702 -2343 32748
rect -2325 32702 -2320 32748
rect -2317 32744 -2309 32748
rect -2062 32744 -2054 32748
rect -2154 32740 -2138 32742
rect -2057 32740 -2054 32744
rect -2292 32734 -2054 32740
rect -2052 32734 -2044 32744
rect -2092 32718 -2062 32720
rect -2094 32714 -2062 32718
rect -2000 32702 -1992 32748
rect -1846 32741 -1806 32748
rect -1663 32744 -1655 32748
rect -1846 32734 -1680 32740
rect -1854 32718 -1806 32720
rect -1854 32714 -1680 32718
rect -1642 32702 -1637 32748
rect -1619 32702 -1614 32748
rect -1530 32702 -1526 32748
rect -1506 32702 -1502 32748
rect -1482 32702 -1478 32748
rect -1458 32702 -1454 32748
rect -1434 32702 -1430 32748
rect -1410 32702 -1406 32748
rect -1386 32702 -1382 32748
rect -1362 32702 -1358 32748
rect -1338 32702 -1334 32748
rect -1314 32702 -1310 32748
rect -1290 32702 -1286 32748
rect -1266 32702 -1262 32748
rect -1242 32702 -1238 32748
rect -1218 32702 -1214 32748
rect -1194 32702 -1190 32748
rect -1170 32702 -1166 32748
rect -1146 32702 -1142 32748
rect -1122 32702 -1118 32748
rect -1098 32702 -1094 32748
rect -1074 32702 -1070 32748
rect -1050 32702 -1046 32748
rect -1026 32702 -1022 32748
rect -1002 32702 -998 32748
rect -978 32702 -974 32748
rect -954 32702 -950 32748
rect -930 32702 -926 32748
rect -906 32702 -902 32748
rect -882 32702 -878 32748
rect -858 32702 -854 32748
rect -834 32702 -830 32748
rect -810 32702 -806 32748
rect -786 32702 -782 32748
rect -762 32702 -758 32748
rect -738 32702 -734 32748
rect -714 32702 -710 32748
rect -690 32702 -686 32748
rect -666 32702 -662 32748
rect -642 32702 -638 32748
rect -618 32702 -614 32748
rect -594 32702 -590 32748
rect -570 32702 -566 32748
rect -546 32702 -542 32748
rect -522 32702 -518 32748
rect -498 32702 -494 32748
rect -474 32702 -470 32748
rect -450 32702 -446 32748
rect -426 32702 -422 32748
rect -402 32702 -398 32748
rect -378 32702 -374 32748
rect -354 32702 -350 32748
rect -330 32702 -326 32748
rect -306 32702 -302 32748
rect -282 32702 -278 32748
rect -258 32702 -254 32748
rect -234 32702 -230 32748
rect -210 32702 -206 32748
rect -186 32702 -182 32748
rect -162 32702 -158 32748
rect -138 32702 -134 32748
rect -114 32702 -110 32748
rect -90 32702 -86 32748
rect -83 32747 -69 32748
rect -66 32747 -59 32771
rect -66 32702 -62 32747
rect -42 32702 -38 32772
rect -18 32702 -14 32772
rect 6 32702 10 32772
rect 30 32702 34 32772
rect 54 32702 58 32772
rect 78 32702 82 32772
rect 102 32702 106 32772
rect 126 32702 130 32772
rect 150 32702 154 32772
rect 174 32702 178 32772
rect 198 32702 202 32772
rect 222 32702 226 32772
rect 246 32702 250 32772
rect 270 32702 274 32772
rect 294 32702 298 32772
rect 318 32702 322 32772
rect 342 32702 346 32772
rect 366 32702 370 32772
rect 390 32702 394 32772
rect 414 32702 418 32772
rect 438 32702 442 32772
rect 462 32702 466 32772
rect 486 32702 490 32772
rect 510 32702 514 32772
rect 534 32702 538 32772
rect 558 32702 562 32772
rect 582 32702 586 32772
rect 606 32702 610 32772
rect 630 32702 634 32772
rect 654 32702 658 32772
rect 678 32702 682 32772
rect 702 32702 706 32772
rect 726 32702 730 32772
rect 750 32702 754 32772
rect 774 32702 778 32772
rect 798 32702 802 32772
rect 822 32702 826 32772
rect 846 32702 850 32772
rect 870 32702 874 32772
rect 894 32702 898 32772
rect 918 32702 922 32772
rect 942 32702 946 32772
rect 966 32702 970 32772
rect 990 32702 994 32772
rect 1014 32702 1018 32772
rect 1038 32702 1042 32772
rect 1062 32702 1066 32772
rect 1075 32717 1080 32727
rect 1086 32717 1090 32772
rect 1085 32703 1090 32717
rect 1075 32702 1109 32703
rect -2393 32700 1109 32702
rect -2371 32678 -2366 32700
rect -2348 32678 -2343 32700
rect -2325 32678 -2320 32700
rect -2072 32698 -2036 32699
rect -2072 32692 -2054 32698
rect -2309 32684 -2301 32692
rect -2317 32678 -2309 32684
rect -2092 32683 -2062 32688
rect -2000 32679 -1992 32700
rect -1938 32699 -1906 32700
rect -1920 32698 -1906 32699
rect -1806 32692 -1680 32698
rect -1854 32683 -1806 32688
rect -1655 32684 -1647 32692
rect -1982 32679 -1966 32680
rect -2000 32678 -1966 32679
rect -1846 32678 -1806 32681
rect -1663 32678 -1655 32684
rect -1642 32678 -1637 32700
rect -1619 32678 -1614 32700
rect -1530 32678 -1526 32700
rect -1506 32678 -1502 32700
rect -1482 32678 -1478 32700
rect -1458 32678 -1454 32700
rect -1434 32678 -1430 32700
rect -1410 32678 -1406 32700
rect -1386 32678 -1382 32700
rect -1362 32678 -1358 32700
rect -1338 32678 -1334 32700
rect -1314 32678 -1310 32700
rect -1290 32678 -1286 32700
rect -1266 32678 -1262 32700
rect -1242 32678 -1238 32700
rect -1218 32678 -1214 32700
rect -1194 32678 -1190 32700
rect -1170 32678 -1166 32700
rect -1146 32678 -1142 32700
rect -1122 32678 -1118 32700
rect -1098 32678 -1094 32700
rect -1074 32678 -1070 32700
rect -1050 32678 -1046 32700
rect -1026 32678 -1022 32700
rect -1002 32678 -998 32700
rect -978 32678 -974 32700
rect -954 32678 -950 32700
rect -930 32678 -926 32700
rect -906 32678 -902 32700
rect -882 32678 -878 32700
rect -858 32678 -854 32700
rect -834 32678 -830 32700
rect -810 32678 -806 32700
rect -786 32678 -782 32700
rect -762 32678 -758 32700
rect -738 32678 -734 32700
rect -714 32678 -710 32700
rect -690 32678 -686 32700
rect -666 32678 -662 32700
rect -642 32678 -638 32700
rect -618 32678 -614 32700
rect -594 32678 -590 32700
rect -570 32678 -566 32700
rect -546 32678 -542 32700
rect -522 32678 -518 32700
rect -498 32678 -494 32700
rect -474 32678 -470 32700
rect -450 32678 -446 32700
rect -426 32678 -422 32700
rect -402 32678 -398 32700
rect -378 32678 -374 32700
rect -354 32678 -350 32700
rect -330 32678 -326 32700
rect -306 32678 -302 32700
rect -282 32678 -278 32700
rect -258 32678 -254 32700
rect -234 32678 -230 32700
rect -210 32678 -206 32700
rect -186 32678 -182 32700
rect -162 32678 -158 32700
rect -138 32678 -134 32700
rect -114 32678 -110 32700
rect -90 32678 -86 32700
rect -66 32678 -62 32700
rect -42 32678 -38 32700
rect -18 32678 -14 32700
rect 6 32678 10 32700
rect 30 32678 34 32700
rect 54 32678 58 32700
rect 78 32678 82 32700
rect 102 32678 106 32700
rect 126 32678 130 32700
rect 150 32678 154 32700
rect 174 32678 178 32700
rect 198 32678 202 32700
rect 222 32678 226 32700
rect 246 32678 250 32700
rect 270 32678 274 32700
rect 294 32678 298 32700
rect 318 32678 322 32700
rect 342 32678 346 32700
rect 366 32678 370 32700
rect 390 32678 394 32700
rect 414 32678 418 32700
rect 438 32678 442 32700
rect 462 32678 466 32700
rect 486 32678 490 32700
rect 510 32678 514 32700
rect 534 32678 538 32700
rect 558 32678 562 32700
rect 582 32678 586 32700
rect 606 32678 610 32700
rect 630 32678 634 32700
rect 654 32678 658 32700
rect 678 32678 682 32700
rect 702 32678 706 32700
rect 726 32678 730 32700
rect 750 32678 754 32700
rect 774 32678 778 32700
rect 798 32678 802 32700
rect 822 32678 826 32700
rect 846 32678 850 32700
rect 870 32678 874 32700
rect 894 32678 898 32700
rect 918 32678 922 32700
rect 942 32678 946 32700
rect 966 32678 970 32700
rect 990 32678 994 32700
rect 1014 32678 1018 32700
rect 1038 32678 1042 32700
rect 1062 32678 1066 32700
rect 1075 32693 1080 32700
rect 1085 32679 1090 32693
rect 1086 32678 1090 32679
rect 1110 32678 1114 32772
rect 1134 32678 1138 32772
rect 1158 32678 1162 32772
rect 1182 32678 1186 32772
rect 1206 32678 1210 32772
rect 1230 32678 1234 32772
rect 1254 32678 1258 32772
rect 1278 32747 1282 32772
rect 1278 32726 1285 32747
rect 1302 32726 1306 32772
rect 1315 32765 1320 32772
rect 1326 32765 1330 32772
rect 1325 32751 1330 32765
rect 1315 32741 1320 32751
rect 1325 32727 1330 32741
rect 1326 32726 1330 32727
rect 1350 32726 1354 32820
rect 1374 32726 1378 32820
rect 1398 32726 1402 32820
rect 1422 32726 1426 32820
rect 1446 32726 1450 32820
rect 1470 32726 1474 32820
rect 1494 32726 1498 32820
rect 1518 32726 1522 32820
rect 1542 32726 1546 32820
rect 1566 32726 1570 32820
rect 1590 32726 1594 32820
rect 1614 32726 1618 32820
rect 1638 32726 1642 32820
rect 1662 32726 1666 32820
rect 1686 32726 1690 32820
rect 1710 32726 1714 32820
rect 1734 32726 1738 32820
rect 1747 32813 1752 32820
rect 1765 32819 1779 32820
rect 1757 32799 1762 32813
rect 1758 32726 1762 32799
rect 1771 32726 1779 32727
rect 1261 32724 1779 32726
rect 1261 32723 1275 32724
rect 1278 32699 1285 32724
rect 1278 32678 1282 32699
rect 1302 32678 1306 32724
rect 1326 32678 1330 32724
rect 1350 32699 1354 32724
rect -2393 32676 1347 32678
rect -2371 32654 -2366 32676
rect -2348 32654 -2343 32676
rect -2325 32654 -2320 32676
rect -2000 32674 -1966 32676
rect -2309 32656 -2301 32664
rect -2062 32663 -2054 32670
rect -2092 32656 -2084 32663
rect -2062 32656 -2026 32658
rect -2317 32654 -2309 32656
rect -2062 32654 -2012 32656
rect -2000 32654 -1992 32674
rect -1982 32673 -1966 32674
rect -1846 32672 -1806 32676
rect -1846 32665 -1798 32670
rect -1806 32663 -1798 32665
rect -1854 32661 -1846 32663
rect -1854 32656 -1806 32661
rect -1655 32656 -1647 32664
rect -1864 32654 -1796 32655
rect -1663 32654 -1655 32656
rect -1642 32654 -1637 32676
rect -1619 32654 -1614 32676
rect -1530 32654 -1526 32676
rect -1506 32654 -1502 32676
rect -1482 32654 -1478 32676
rect -1458 32654 -1454 32676
rect -1434 32654 -1430 32676
rect -1410 32654 -1406 32676
rect -1386 32654 -1382 32676
rect -1362 32654 -1358 32676
rect -1338 32654 -1334 32676
rect -1314 32654 -1310 32676
rect -1290 32654 -1286 32676
rect -1266 32654 -1262 32676
rect -1242 32654 -1238 32676
rect -1218 32654 -1214 32676
rect -1194 32654 -1190 32676
rect -1170 32654 -1166 32676
rect -1146 32654 -1142 32676
rect -1122 32654 -1118 32676
rect -1098 32654 -1094 32676
rect -1074 32654 -1070 32676
rect -1050 32654 -1046 32676
rect -1026 32654 -1022 32676
rect -1002 32654 -998 32676
rect -978 32654 -974 32676
rect -954 32654 -950 32676
rect -930 32654 -926 32676
rect -906 32654 -902 32676
rect -882 32654 -878 32676
rect -858 32654 -854 32676
rect -834 32654 -830 32676
rect -810 32654 -806 32676
rect -786 32654 -782 32676
rect -762 32654 -758 32676
rect -738 32654 -734 32676
rect -714 32654 -710 32676
rect -690 32654 -686 32676
rect -666 32654 -662 32676
rect -642 32654 -638 32676
rect -618 32654 -614 32676
rect -594 32654 -590 32676
rect -570 32654 -566 32676
rect -546 32654 -542 32676
rect -522 32654 -518 32676
rect -498 32654 -494 32676
rect -474 32654 -470 32676
rect -450 32654 -446 32676
rect -426 32654 -422 32676
rect -402 32654 -398 32676
rect -378 32654 -374 32676
rect -354 32654 -350 32676
rect -330 32654 -326 32676
rect -306 32654 -302 32676
rect -282 32654 -278 32676
rect -258 32654 -254 32676
rect -234 32654 -230 32676
rect -210 32654 -206 32676
rect -186 32654 -182 32676
rect -162 32654 -158 32676
rect -138 32654 -134 32676
rect -114 32654 -110 32676
rect -90 32654 -86 32676
rect -66 32654 -62 32676
rect -42 32654 -38 32676
rect -18 32654 -14 32676
rect 6 32654 10 32676
rect 30 32654 34 32676
rect 54 32654 58 32676
rect 78 32654 82 32676
rect 102 32654 106 32676
rect 126 32654 130 32676
rect 150 32654 154 32676
rect 174 32654 178 32676
rect 198 32654 202 32676
rect 222 32654 226 32676
rect 246 32654 250 32676
rect 270 32654 274 32676
rect 294 32654 298 32676
rect 318 32654 322 32676
rect 342 32654 346 32676
rect 366 32654 370 32676
rect 390 32654 394 32676
rect 414 32654 418 32676
rect 438 32654 442 32676
rect 462 32654 466 32676
rect 486 32654 490 32676
rect 510 32654 514 32676
rect 534 32654 538 32676
rect 558 32654 562 32676
rect 582 32654 586 32676
rect 606 32654 610 32676
rect 630 32654 634 32676
rect 654 32654 658 32676
rect 678 32654 682 32676
rect 702 32654 706 32676
rect 726 32654 730 32676
rect 750 32654 754 32676
rect 774 32654 778 32676
rect 798 32654 802 32676
rect 822 32654 826 32676
rect 846 32654 850 32676
rect 870 32654 874 32676
rect 894 32654 898 32676
rect 918 32654 922 32676
rect 942 32654 946 32676
rect 966 32654 970 32676
rect 990 32654 994 32676
rect 1014 32654 1018 32676
rect 1038 32654 1042 32676
rect 1062 32654 1066 32676
rect 1086 32654 1090 32676
rect 1110 32654 1114 32676
rect 1134 32654 1138 32676
rect 1158 32654 1162 32676
rect 1182 32654 1186 32676
rect 1206 32654 1210 32676
rect 1230 32654 1234 32676
rect 1254 32654 1258 32676
rect 1278 32654 1282 32676
rect 1302 32654 1306 32676
rect 1326 32654 1330 32676
rect 1333 32675 1347 32676
rect -2393 32652 1347 32654
rect -2371 32606 -2366 32652
rect -2348 32606 -2343 32652
rect -2325 32606 -2320 32652
rect -2317 32648 -2309 32652
rect -2062 32648 -2054 32652
rect -2154 32644 -2138 32646
rect -2057 32644 -2054 32648
rect -2292 32638 -2054 32644
rect -2052 32638 -2044 32648
rect -2092 32622 -2062 32624
rect -2094 32618 -2062 32622
rect -2000 32606 -1992 32652
rect -1846 32645 -1806 32652
rect -1663 32648 -1655 32652
rect -1846 32638 -1680 32644
rect -1854 32622 -1806 32624
rect -1854 32618 -1680 32622
rect -1642 32606 -1637 32652
rect -1619 32606 -1614 32652
rect -1530 32606 -1526 32652
rect -1506 32606 -1502 32652
rect -1482 32606 -1478 32652
rect -1458 32606 -1454 32652
rect -1434 32606 -1430 32652
rect -1410 32606 -1406 32652
rect -1386 32606 -1382 32652
rect -1362 32606 -1358 32652
rect -1338 32606 -1334 32652
rect -1314 32606 -1310 32652
rect -1290 32606 -1286 32652
rect -1266 32606 -1262 32652
rect -1242 32606 -1238 32652
rect -1218 32606 -1214 32652
rect -1194 32606 -1190 32652
rect -1170 32606 -1166 32652
rect -1146 32606 -1142 32652
rect -1122 32606 -1118 32652
rect -1098 32606 -1094 32652
rect -1074 32606 -1070 32652
rect -1050 32606 -1046 32652
rect -1026 32606 -1022 32652
rect -1002 32606 -998 32652
rect -978 32606 -974 32652
rect -954 32606 -950 32652
rect -930 32606 -926 32652
rect -906 32606 -902 32652
rect -882 32606 -878 32652
rect -858 32606 -854 32652
rect -834 32606 -830 32652
rect -810 32606 -806 32652
rect -786 32606 -782 32652
rect -762 32606 -758 32652
rect -738 32606 -734 32652
rect -714 32606 -710 32652
rect -690 32606 -686 32652
rect -666 32606 -662 32652
rect -642 32606 -638 32652
rect -618 32606 -614 32652
rect -594 32606 -590 32652
rect -570 32606 -566 32652
rect -546 32606 -542 32652
rect -522 32606 -518 32652
rect -498 32606 -494 32652
rect -474 32606 -470 32652
rect -450 32606 -446 32652
rect -426 32606 -422 32652
rect -402 32606 -398 32652
rect -378 32606 -374 32652
rect -354 32606 -350 32652
rect -330 32606 -326 32652
rect -306 32606 -302 32652
rect -282 32606 -278 32652
rect -258 32606 -254 32652
rect -234 32606 -230 32652
rect -210 32606 -206 32652
rect -186 32606 -182 32652
rect -162 32606 -158 32652
rect -138 32606 -134 32652
rect -114 32606 -110 32652
rect -90 32606 -86 32652
rect -66 32606 -62 32652
rect -42 32606 -38 32652
rect -18 32606 -14 32652
rect 6 32606 10 32652
rect 30 32606 34 32652
rect 54 32606 58 32652
rect 78 32606 82 32652
rect 102 32606 106 32652
rect 126 32606 130 32652
rect 150 32606 154 32652
rect 174 32606 178 32652
rect 198 32606 202 32652
rect 222 32606 226 32652
rect 246 32606 250 32652
rect 270 32606 274 32652
rect 294 32606 298 32652
rect 318 32606 322 32652
rect 342 32606 346 32652
rect 366 32606 370 32652
rect 390 32606 394 32652
rect 414 32606 418 32652
rect 438 32606 442 32652
rect 462 32606 466 32652
rect 486 32606 490 32652
rect 510 32606 514 32652
rect 534 32606 538 32652
rect 558 32606 562 32652
rect 582 32606 586 32652
rect 606 32606 610 32652
rect 630 32606 634 32652
rect 654 32606 658 32652
rect 678 32606 682 32652
rect 702 32606 706 32652
rect 726 32606 730 32652
rect 750 32606 754 32652
rect 774 32606 778 32652
rect 798 32606 802 32652
rect 822 32606 826 32652
rect 846 32606 850 32652
rect 870 32606 874 32652
rect 894 32606 898 32652
rect 918 32606 922 32652
rect 942 32606 946 32652
rect 966 32606 970 32652
rect 990 32606 994 32652
rect 1003 32621 1008 32631
rect 1014 32621 1018 32652
rect 1013 32607 1018 32621
rect 1003 32606 1037 32607
rect -2393 32604 1037 32606
rect -2371 32582 -2366 32604
rect -2348 32582 -2343 32604
rect -2325 32582 -2320 32604
rect -2072 32602 -2036 32603
rect -2072 32596 -2054 32602
rect -2309 32588 -2301 32596
rect -2317 32582 -2309 32588
rect -2092 32587 -2062 32592
rect -2000 32583 -1992 32604
rect -1938 32603 -1906 32604
rect -1920 32602 -1906 32603
rect -1806 32596 -1680 32602
rect -1854 32587 -1806 32592
rect -1655 32588 -1647 32596
rect -1982 32583 -1966 32584
rect -2000 32582 -1966 32583
rect -1846 32582 -1806 32585
rect -1663 32582 -1655 32588
rect -1642 32582 -1637 32604
rect -1619 32582 -1614 32604
rect -1530 32582 -1526 32604
rect -1506 32582 -1502 32604
rect -1482 32582 -1478 32604
rect -1458 32582 -1454 32604
rect -1434 32582 -1430 32604
rect -1410 32582 -1406 32604
rect -1386 32582 -1382 32604
rect -1362 32582 -1358 32604
rect -1338 32582 -1334 32604
rect -1314 32582 -1310 32604
rect -1290 32582 -1286 32604
rect -1266 32582 -1262 32604
rect -1242 32582 -1238 32604
rect -1218 32582 -1214 32604
rect -1194 32582 -1190 32604
rect -1170 32582 -1166 32604
rect -1146 32582 -1142 32604
rect -1122 32582 -1118 32604
rect -1098 32582 -1094 32604
rect -1074 32582 -1070 32604
rect -1050 32582 -1046 32604
rect -1026 32582 -1022 32604
rect -1002 32582 -998 32604
rect -978 32582 -974 32604
rect -954 32582 -950 32604
rect -930 32582 -926 32604
rect -906 32582 -902 32604
rect -882 32582 -878 32604
rect -858 32582 -854 32604
rect -834 32582 -830 32604
rect -810 32582 -806 32604
rect -786 32582 -782 32604
rect -762 32582 -758 32604
rect -738 32582 -734 32604
rect -714 32582 -710 32604
rect -690 32582 -686 32604
rect -666 32582 -662 32604
rect -642 32582 -638 32604
rect -618 32582 -614 32604
rect -594 32582 -590 32604
rect -570 32582 -566 32604
rect -546 32582 -542 32604
rect -522 32582 -518 32604
rect -498 32582 -494 32604
rect -474 32582 -470 32604
rect -450 32582 -446 32604
rect -426 32582 -422 32604
rect -402 32582 -398 32604
rect -378 32582 -374 32604
rect -354 32582 -350 32604
rect -330 32582 -326 32604
rect -306 32582 -302 32604
rect -282 32582 -278 32604
rect -258 32582 -254 32604
rect -234 32582 -230 32604
rect -210 32582 -206 32604
rect -186 32582 -182 32604
rect -162 32582 -158 32604
rect -138 32582 -134 32604
rect -114 32582 -110 32604
rect -90 32582 -86 32604
rect -66 32582 -62 32604
rect -42 32582 -38 32604
rect -18 32582 -14 32604
rect 6 32582 10 32604
rect 30 32582 34 32604
rect 54 32582 58 32604
rect 78 32582 82 32604
rect 102 32582 106 32604
rect 126 32582 130 32604
rect 150 32582 154 32604
rect 174 32582 178 32604
rect 198 32582 202 32604
rect 222 32582 226 32604
rect 246 32582 250 32604
rect 270 32582 274 32604
rect 294 32582 298 32604
rect 318 32582 322 32604
rect 342 32582 346 32604
rect 366 32582 370 32604
rect 390 32582 394 32604
rect 414 32582 418 32604
rect 438 32582 442 32604
rect 462 32582 466 32604
rect 486 32582 490 32604
rect 510 32582 514 32604
rect 534 32582 538 32604
rect 558 32582 562 32604
rect 582 32582 586 32604
rect 606 32582 610 32604
rect 630 32582 634 32604
rect 654 32582 658 32604
rect 678 32582 682 32604
rect 702 32582 706 32604
rect 726 32582 730 32604
rect 750 32582 754 32604
rect 774 32582 778 32604
rect 798 32582 802 32604
rect 822 32582 826 32604
rect 846 32582 850 32604
rect 870 32582 874 32604
rect 894 32582 898 32604
rect 918 32582 922 32604
rect 942 32582 946 32604
rect 966 32582 970 32604
rect 990 32582 994 32604
rect 1003 32597 1008 32604
rect 1013 32583 1018 32597
rect 1014 32582 1018 32583
rect 1038 32582 1042 32652
rect 1062 32582 1066 32652
rect 1086 32582 1090 32652
rect 1110 32651 1114 32652
rect 1110 32630 1117 32651
rect 1134 32630 1138 32652
rect 1158 32630 1162 32652
rect 1182 32630 1186 32652
rect 1206 32630 1210 32652
rect 1230 32630 1234 32652
rect 1254 32630 1258 32652
rect 1278 32630 1282 32652
rect 1302 32630 1306 32652
rect 1326 32630 1330 32652
rect 1333 32651 1347 32652
rect 1350 32651 1357 32699
rect 1350 32630 1354 32651
rect 1374 32630 1378 32724
rect 1398 32630 1402 32724
rect 1422 32630 1426 32724
rect 1446 32630 1450 32724
rect 1470 32630 1474 32724
rect 1494 32630 1498 32724
rect 1518 32630 1522 32724
rect 1542 32630 1546 32724
rect 1566 32630 1570 32724
rect 1590 32630 1594 32724
rect 1614 32630 1618 32724
rect 1638 32630 1642 32724
rect 1662 32630 1666 32724
rect 1686 32630 1690 32724
rect 1710 32630 1714 32724
rect 1734 32630 1738 32724
rect 1747 32645 1752 32655
rect 1758 32645 1762 32724
rect 1765 32723 1779 32724
rect 1771 32717 1776 32723
rect 1781 32703 1786 32717
rect 1771 32669 1776 32679
rect 1782 32669 1786 32703
rect 1781 32655 1786 32669
rect 1757 32631 1762 32645
rect 1747 32630 1781 32631
rect 1093 32628 1781 32630
rect 1093 32627 1107 32628
rect 1110 32603 1117 32628
rect 1110 32582 1114 32603
rect 1134 32582 1138 32628
rect 1158 32582 1162 32628
rect 1182 32582 1186 32628
rect 1206 32582 1210 32628
rect 1230 32582 1234 32628
rect 1254 32582 1258 32628
rect 1278 32582 1282 32628
rect 1302 32582 1306 32628
rect 1326 32582 1330 32628
rect 1350 32582 1354 32628
rect 1374 32582 1378 32628
rect 1398 32582 1402 32628
rect 1422 32582 1426 32628
rect 1446 32582 1450 32628
rect 1470 32582 1474 32628
rect 1494 32582 1498 32628
rect 1518 32582 1522 32628
rect 1542 32582 1546 32628
rect 1566 32582 1570 32628
rect 1590 32582 1594 32628
rect 1614 32582 1618 32628
rect 1638 32582 1642 32628
rect 1662 32582 1666 32628
rect 1686 32582 1690 32628
rect 1710 32582 1714 32628
rect 1734 32582 1738 32628
rect 1747 32621 1752 32628
rect 1757 32607 1762 32621
rect 1758 32583 1762 32607
rect 1747 32582 1781 32583
rect -2393 32580 1781 32582
rect -2371 32558 -2366 32580
rect -2348 32558 -2343 32580
rect -2325 32558 -2320 32580
rect -2000 32578 -1966 32580
rect -2309 32560 -2301 32568
rect -2062 32567 -2054 32574
rect -2092 32560 -2084 32567
rect -2062 32560 -2026 32562
rect -2317 32558 -2309 32560
rect -2062 32558 -2012 32560
rect -2000 32558 -1992 32578
rect -1982 32577 -1966 32578
rect -1846 32576 -1806 32580
rect -1846 32569 -1798 32574
rect -1806 32567 -1798 32569
rect -1854 32565 -1846 32567
rect -1854 32560 -1806 32565
rect -1655 32560 -1647 32568
rect -1864 32558 -1796 32559
rect -1663 32558 -1655 32560
rect -1642 32558 -1637 32580
rect -1619 32558 -1614 32580
rect -1530 32558 -1526 32580
rect -1506 32558 -1502 32580
rect -1482 32558 -1478 32580
rect -1458 32558 -1454 32580
rect -1434 32558 -1430 32580
rect -1410 32558 -1406 32580
rect -1386 32558 -1382 32580
rect -1362 32558 -1358 32580
rect -1338 32558 -1334 32580
rect -1314 32558 -1310 32580
rect -1290 32558 -1286 32580
rect -1266 32558 -1262 32580
rect -1242 32558 -1238 32580
rect -1218 32558 -1214 32580
rect -1194 32558 -1190 32580
rect -1170 32558 -1166 32580
rect -1146 32558 -1142 32580
rect -1122 32558 -1118 32580
rect -1098 32558 -1094 32580
rect -1074 32558 -1070 32580
rect -1050 32558 -1046 32580
rect -1026 32558 -1022 32580
rect -1002 32558 -998 32580
rect -978 32558 -974 32580
rect -954 32558 -950 32580
rect -930 32558 -926 32580
rect -906 32558 -902 32580
rect -882 32558 -878 32580
rect -858 32558 -854 32580
rect -834 32558 -830 32580
rect -810 32558 -806 32580
rect -786 32558 -782 32580
rect -762 32558 -758 32580
rect -738 32558 -734 32580
rect -714 32558 -710 32580
rect -690 32558 -686 32580
rect -666 32558 -662 32580
rect -642 32558 -638 32580
rect -618 32558 -614 32580
rect -594 32558 -590 32580
rect -570 32558 -566 32580
rect -546 32558 -542 32580
rect -522 32558 -518 32580
rect -498 32558 -494 32580
rect -474 32558 -470 32580
rect -450 32558 -446 32580
rect -426 32558 -422 32580
rect -402 32558 -398 32580
rect -378 32558 -374 32580
rect -354 32558 -350 32580
rect -330 32558 -326 32580
rect -306 32558 -302 32580
rect -282 32558 -278 32580
rect -258 32558 -254 32580
rect -234 32558 -230 32580
rect -210 32558 -206 32580
rect -186 32558 -182 32580
rect -162 32558 -158 32580
rect -138 32558 -134 32580
rect -114 32558 -110 32580
rect -90 32558 -86 32580
rect -66 32558 -62 32580
rect -42 32558 -38 32580
rect -18 32558 -14 32580
rect 6 32558 10 32580
rect 30 32558 34 32580
rect 54 32558 58 32580
rect 78 32558 82 32580
rect 102 32558 106 32580
rect 126 32558 130 32580
rect 150 32558 154 32580
rect 174 32558 178 32580
rect 198 32558 202 32580
rect 222 32558 226 32580
rect 246 32558 250 32580
rect 270 32558 274 32580
rect 294 32558 298 32580
rect 318 32558 322 32580
rect 342 32558 346 32580
rect 366 32558 370 32580
rect 390 32558 394 32580
rect 414 32558 418 32580
rect 438 32558 442 32580
rect 462 32558 466 32580
rect 486 32558 490 32580
rect 510 32558 514 32580
rect 534 32558 538 32580
rect 558 32558 562 32580
rect 582 32558 586 32580
rect 606 32558 610 32580
rect 630 32559 634 32580
rect 619 32558 653 32559
rect -2393 32556 653 32558
rect -2371 32510 -2366 32556
rect -2348 32510 -2343 32556
rect -2325 32510 -2320 32556
rect -2317 32552 -2309 32556
rect -2062 32552 -2054 32556
rect -2154 32548 -2138 32550
rect -2057 32548 -2054 32552
rect -2292 32542 -2054 32548
rect -2052 32542 -2044 32552
rect -2092 32526 -2062 32528
rect -2094 32522 -2062 32526
rect -2000 32510 -1992 32556
rect -1846 32549 -1806 32556
rect -1663 32552 -1655 32556
rect -1846 32542 -1680 32548
rect -1854 32526 -1806 32528
rect -1854 32522 -1680 32526
rect -1642 32510 -1637 32556
rect -1619 32510 -1614 32556
rect -1530 32510 -1526 32556
rect -1506 32510 -1502 32556
rect -1482 32510 -1478 32556
rect -1458 32510 -1454 32556
rect -1434 32510 -1430 32556
rect -1410 32510 -1406 32556
rect -1386 32510 -1382 32556
rect -1362 32510 -1358 32556
rect -1338 32510 -1334 32556
rect -1314 32510 -1310 32556
rect -1290 32510 -1286 32556
rect -1266 32510 -1262 32556
rect -1242 32510 -1238 32556
rect -1218 32510 -1214 32556
rect -1194 32510 -1190 32556
rect -1170 32510 -1166 32556
rect -1146 32510 -1142 32556
rect -1122 32510 -1118 32556
rect -1098 32510 -1094 32556
rect -1074 32510 -1070 32556
rect -1050 32510 -1046 32556
rect -1026 32510 -1022 32556
rect -1002 32510 -998 32556
rect -978 32510 -974 32556
rect -954 32510 -950 32556
rect -930 32510 -926 32556
rect -906 32510 -902 32556
rect -882 32510 -878 32556
rect -858 32510 -854 32556
rect -834 32510 -830 32556
rect -821 32525 -816 32535
rect -810 32525 -806 32556
rect -811 32511 -806 32525
rect -821 32510 -787 32511
rect -2393 32508 -787 32510
rect -2371 32486 -2366 32508
rect -2348 32486 -2343 32508
rect -2325 32486 -2320 32508
rect -2072 32506 -2036 32507
rect -2072 32500 -2054 32506
rect -2309 32492 -2301 32500
rect -2317 32486 -2309 32492
rect -2092 32491 -2062 32496
rect -2000 32487 -1992 32508
rect -1938 32507 -1906 32508
rect -1920 32506 -1906 32507
rect -1806 32500 -1680 32506
rect -1854 32491 -1806 32496
rect -1655 32492 -1647 32500
rect -1982 32487 -1966 32488
rect -2000 32486 -1966 32487
rect -1846 32486 -1806 32489
rect -1663 32486 -1655 32492
rect -1642 32486 -1637 32508
rect -1619 32486 -1614 32508
rect -1530 32486 -1526 32508
rect -1506 32486 -1502 32508
rect -1482 32486 -1478 32508
rect -1458 32486 -1454 32508
rect -1434 32486 -1430 32508
rect -1410 32486 -1406 32508
rect -1386 32486 -1382 32508
rect -1362 32487 -1358 32508
rect -1373 32486 -1339 32487
rect -2393 32484 -1339 32486
rect -2371 32462 -2366 32484
rect -2348 32462 -2343 32484
rect -2325 32462 -2320 32484
rect -2000 32482 -1966 32484
rect -2309 32464 -2301 32472
rect -2062 32471 -2054 32478
rect -2092 32464 -2084 32471
rect -2062 32464 -2026 32466
rect -2317 32462 -2309 32464
rect -2062 32462 -2012 32464
rect -2000 32462 -1992 32482
rect -1982 32481 -1966 32482
rect -1846 32480 -1806 32484
rect -1846 32473 -1798 32478
rect -1806 32471 -1798 32473
rect -1854 32469 -1846 32471
rect -1854 32464 -1806 32469
rect -1655 32464 -1647 32472
rect -1864 32462 -1796 32463
rect -1663 32462 -1655 32464
rect -1642 32462 -1637 32484
rect -1619 32462 -1614 32484
rect -1530 32462 -1526 32484
rect -1506 32462 -1502 32484
rect -1482 32462 -1478 32484
rect -1458 32462 -1454 32484
rect -1434 32462 -1430 32484
rect -1410 32462 -1406 32484
rect -1386 32462 -1382 32484
rect -1373 32477 -1368 32484
rect -1362 32477 -1358 32484
rect -1363 32463 -1358 32477
rect -1362 32462 -1358 32463
rect -1338 32462 -1334 32508
rect -1314 32462 -1310 32508
rect -1290 32462 -1286 32508
rect -1266 32462 -1262 32508
rect -1242 32462 -1238 32508
rect -1218 32462 -1214 32508
rect -1194 32462 -1190 32508
rect -1170 32462 -1166 32508
rect -1146 32462 -1142 32508
rect -1122 32462 -1118 32508
rect -1098 32462 -1094 32508
rect -1074 32462 -1070 32508
rect -1050 32462 -1046 32508
rect -1026 32462 -1022 32508
rect -1002 32462 -998 32508
rect -978 32462 -974 32508
rect -954 32462 -950 32508
rect -930 32462 -926 32508
rect -906 32462 -902 32508
rect -882 32462 -878 32508
rect -858 32462 -854 32508
rect -834 32462 -830 32508
rect -821 32501 -816 32508
rect -811 32487 -806 32501
rect -810 32462 -806 32487
rect -786 32462 -782 32556
rect -762 32462 -758 32556
rect -738 32462 -734 32556
rect -714 32462 -710 32556
rect -690 32462 -686 32556
rect -666 32462 -662 32556
rect -642 32462 -638 32556
rect -618 32462 -614 32556
rect -594 32462 -590 32556
rect -570 32462 -566 32556
rect -546 32462 -542 32556
rect -522 32462 -518 32556
rect -498 32462 -494 32556
rect -474 32462 -470 32556
rect -450 32462 -446 32556
rect -426 32462 -422 32556
rect -402 32462 -398 32556
rect -378 32462 -374 32556
rect -354 32462 -350 32556
rect -330 32462 -326 32556
rect -306 32462 -302 32556
rect -282 32462 -278 32556
rect -258 32462 -254 32556
rect -234 32462 -230 32556
rect -210 32462 -206 32556
rect -186 32462 -182 32556
rect -162 32462 -158 32556
rect -138 32462 -134 32556
rect -114 32462 -110 32556
rect -90 32462 -86 32556
rect -66 32462 -62 32556
rect -42 32462 -38 32556
rect -18 32462 -14 32556
rect 6 32462 10 32556
rect 30 32462 34 32556
rect 54 32462 58 32556
rect 78 32462 82 32556
rect 102 32462 106 32556
rect 126 32462 130 32556
rect 150 32462 154 32556
rect 174 32462 178 32556
rect 198 32462 202 32556
rect 222 32462 226 32556
rect 246 32462 250 32556
rect 270 32462 274 32556
rect 294 32462 298 32556
rect 318 32462 322 32556
rect 342 32462 346 32556
rect 366 32462 370 32556
rect 390 32462 394 32556
rect 414 32462 418 32556
rect 438 32462 442 32556
rect 462 32462 466 32556
rect 486 32462 490 32556
rect 510 32462 514 32556
rect 534 32462 538 32556
rect 558 32462 562 32556
rect 582 32462 586 32556
rect 606 32462 610 32556
rect 619 32549 624 32556
rect 630 32549 634 32556
rect 629 32535 634 32549
rect 630 32462 634 32535
rect 654 32483 658 32580
rect -2393 32460 651 32462
rect -2371 32390 -2366 32460
rect -2348 32390 -2343 32460
rect -2325 32390 -2320 32460
rect -2317 32456 -2309 32460
rect -2062 32456 -2054 32460
rect -2154 32452 -2138 32454
rect -2057 32452 -2054 32456
rect -2292 32446 -2054 32452
rect -2052 32446 -2044 32456
rect -2092 32430 -2062 32432
rect -2094 32426 -2062 32430
rect -2309 32396 -2301 32402
rect -2317 32390 -2309 32396
rect -2000 32390 -1992 32460
rect -1846 32453 -1806 32460
rect -1663 32456 -1655 32460
rect -1846 32446 -1680 32452
rect -1854 32430 -1806 32432
rect -1854 32426 -1680 32430
rect -1655 32396 -1647 32402
rect -1663 32390 -1655 32396
rect -1642 32390 -1637 32460
rect -1619 32390 -1614 32460
rect -1530 32390 -1526 32460
rect -1506 32390 -1502 32460
rect -1482 32390 -1478 32460
rect -1458 32390 -1454 32460
rect -1434 32390 -1430 32460
rect -1410 32390 -1406 32460
rect -1386 32390 -1382 32460
rect -1362 32390 -1358 32460
rect -1338 32411 -1334 32460
rect -2393 32388 -1341 32390
rect -2371 32294 -2366 32388
rect -2348 32294 -2343 32388
rect -2325 32326 -2320 32388
rect -2317 32386 -2309 32388
rect -2000 32387 -1966 32388
rect -2000 32386 -1982 32387
rect -1663 32386 -1655 32388
rect -2028 32378 -2018 32380
rect -2309 32368 -2301 32374
rect -2091 32368 -2061 32375
rect -2317 32358 -2309 32368
rect -2044 32366 -2028 32368
rect -2026 32366 -2014 32378
rect -2084 32360 -2061 32366
rect -2044 32364 -2014 32366
rect -2292 32350 -2054 32359
rect -2325 32318 -2317 32326
rect -2325 32298 -2320 32318
rect -2317 32310 -2309 32318
rect -2325 32294 -2317 32298
rect -2000 32294 -1992 32386
rect -1982 32385 -1966 32386
rect -1980 32368 -1932 32375
rect -1655 32368 -1647 32374
rect -1846 32350 -1680 32359
rect -1663 32358 -1655 32368
rect -1671 32318 -1663 32326
rect -1663 32310 -1655 32318
rect -1671 32294 -1663 32298
rect -1642 32294 -1637 32388
rect -1619 32294 -1614 32388
rect -1530 32294 -1526 32388
rect -1506 32294 -1502 32388
rect -1482 32294 -1478 32388
rect -1458 32294 -1454 32388
rect -1434 32294 -1430 32388
rect -1410 32294 -1406 32388
rect -1386 32294 -1382 32388
rect -1362 32294 -1358 32388
rect -1355 32387 -1341 32388
rect -1338 32387 -1331 32411
rect -1338 32294 -1334 32387
rect -1314 32294 -1310 32460
rect -1290 32294 -1286 32460
rect -1266 32294 -1262 32460
rect -1242 32294 -1238 32460
rect -1218 32294 -1214 32460
rect -1194 32294 -1190 32460
rect -1170 32294 -1166 32460
rect -1146 32294 -1142 32460
rect -1122 32294 -1118 32460
rect -1098 32294 -1094 32460
rect -1074 32294 -1070 32460
rect -1050 32294 -1046 32460
rect -1026 32294 -1022 32460
rect -1002 32294 -998 32460
rect -978 32294 -974 32460
rect -954 32294 -950 32460
rect -930 32294 -926 32460
rect -906 32294 -902 32460
rect -882 32294 -878 32460
rect -858 32294 -854 32460
rect -834 32294 -830 32460
rect -810 32294 -806 32460
rect -786 32459 -782 32460
rect -786 32411 -779 32459
rect -786 32294 -782 32411
rect -762 32294 -758 32460
rect -738 32294 -734 32460
rect -714 32294 -710 32460
rect -690 32294 -686 32460
rect -666 32294 -662 32460
rect -642 32294 -638 32460
rect -618 32294 -614 32460
rect -594 32294 -590 32460
rect -570 32294 -566 32460
rect -546 32294 -542 32460
rect -522 32294 -518 32460
rect -498 32294 -494 32460
rect -474 32294 -470 32460
rect -450 32294 -446 32460
rect -426 32294 -422 32460
rect -402 32294 -398 32460
rect -378 32294 -374 32460
rect -354 32294 -350 32460
rect -330 32294 -326 32460
rect -306 32294 -302 32460
rect -282 32294 -278 32460
rect -258 32294 -254 32460
rect -234 32294 -230 32460
rect -210 32294 -206 32460
rect -186 32294 -182 32460
rect -162 32294 -158 32460
rect -138 32294 -134 32460
rect -114 32294 -110 32460
rect -90 32294 -86 32460
rect -77 32333 -72 32343
rect -66 32333 -62 32460
rect -67 32319 -62 32333
rect -66 32294 -62 32319
rect -42 32294 -38 32460
rect -18 32294 -14 32460
rect 6 32294 10 32460
rect 30 32294 34 32460
rect 54 32294 58 32460
rect 78 32294 82 32460
rect 102 32294 106 32460
rect 126 32294 130 32460
rect 150 32294 154 32460
rect 174 32294 178 32460
rect 198 32294 202 32460
rect 222 32294 226 32460
rect 246 32294 250 32460
rect 259 32405 264 32415
rect 270 32405 274 32460
rect 269 32391 274 32405
rect 259 32381 264 32391
rect 269 32367 274 32381
rect 270 32294 274 32367
rect 294 32339 298 32460
rect -2393 32292 -1969 32294
rect -1955 32292 291 32294
rect -2371 32246 -2366 32292
rect -2348 32246 -2343 32292
rect -2325 32282 -2317 32292
rect -2080 32290 -1969 32292
rect -2080 32284 -2053 32290
rect -2325 32266 -2320 32282
rect -2309 32270 -2301 32282
rect -2070 32275 -2040 32282
rect -2000 32274 -1992 32290
rect -1972 32286 -1969 32290
rect -1972 32284 -1955 32286
rect -1955 32274 -1850 32283
rect -1671 32282 -1663 32292
rect -2317 32266 -2309 32270
rect -2070 32267 -2053 32273
rect -2027 32272 -1992 32274
rect -1969 32272 -1955 32273
rect -2325 32254 -2317 32266
rect -2292 32257 -2053 32266
rect -2325 32246 -2320 32254
rect -2309 32246 -2301 32254
rect -2000 32246 -1992 32272
rect -1655 32270 -1647 32282
rect -1663 32266 -1655 32270
rect -1972 32258 -1924 32265
rect -1945 32257 -1929 32258
rect -1860 32257 -1680 32266
rect -1671 32254 -1663 32266
rect -1978 32246 -1942 32247
rect -1655 32246 -1647 32254
rect -1642 32246 -1637 32292
rect -1619 32246 -1614 32292
rect -1530 32246 -1526 32292
rect -1506 32246 -1502 32292
rect -1482 32246 -1478 32292
rect -1458 32246 -1454 32292
rect -1434 32246 -1430 32292
rect -1410 32246 -1406 32292
rect -1386 32246 -1382 32292
rect -1362 32246 -1358 32292
rect -1338 32246 -1334 32292
rect -1314 32246 -1310 32292
rect -1290 32246 -1286 32292
rect -1266 32246 -1262 32292
rect -1242 32246 -1238 32292
rect -1218 32246 -1214 32292
rect -1194 32246 -1190 32292
rect -1170 32246 -1166 32292
rect -1146 32246 -1142 32292
rect -1122 32246 -1118 32292
rect -1098 32246 -1094 32292
rect -1074 32246 -1070 32292
rect -1050 32246 -1046 32292
rect -1026 32246 -1022 32292
rect -1002 32246 -998 32292
rect -978 32246 -974 32292
rect -954 32246 -950 32292
rect -930 32246 -926 32292
rect -906 32246 -902 32292
rect -882 32246 -878 32292
rect -858 32246 -854 32292
rect -834 32246 -830 32292
rect -810 32246 -806 32292
rect -786 32246 -782 32292
rect -762 32246 -758 32292
rect -738 32246 -734 32292
rect -714 32246 -710 32292
rect -690 32246 -686 32292
rect -666 32246 -662 32292
rect -642 32246 -638 32292
rect -618 32246 -614 32292
rect -594 32246 -590 32292
rect -570 32246 -566 32292
rect -546 32246 -542 32292
rect -522 32246 -518 32292
rect -498 32246 -494 32292
rect -474 32246 -470 32292
rect -450 32246 -446 32292
rect -426 32246 -422 32292
rect -402 32246 -398 32292
rect -378 32246 -374 32292
rect -354 32246 -350 32292
rect -330 32246 -326 32292
rect -306 32246 -302 32292
rect -282 32246 -278 32292
rect -258 32246 -254 32292
rect -234 32246 -230 32292
rect -210 32246 -206 32292
rect -186 32246 -182 32292
rect -162 32247 -158 32292
rect -173 32246 -139 32247
rect -2393 32244 -139 32246
rect -2371 32150 -2366 32244
rect -2348 32150 -2343 32244
rect -2325 32238 -2320 32244
rect -2309 32242 -2301 32244
rect -2317 32238 -2309 32242
rect -2325 32226 -2317 32238
rect -2325 32206 -2320 32226
rect -2062 32206 -2032 32207
rect -2000 32206 -1992 32244
rect -1655 32242 -1647 32244
rect -1663 32238 -1655 32242
rect -1671 32226 -1663 32238
rect -1942 32208 -1937 32220
rect -1850 32217 -1822 32218
rect -1850 32213 -1802 32217
rect -2325 32198 -2317 32206
rect -2062 32204 -1961 32206
rect -2325 32178 -2320 32198
rect -2317 32190 -2309 32198
rect -2062 32191 -2040 32202
rect -2032 32197 -1961 32204
rect -1947 32198 -1942 32206
rect -1842 32204 -1794 32207
rect -2070 32186 -2022 32190
rect -2325 32164 -2317 32178
rect -2072 32170 -2032 32171
rect -2102 32164 -2032 32170
rect -2325 32150 -2320 32164
rect -2317 32162 -2309 32164
rect -2309 32150 -2301 32162
rect -2070 32155 -2062 32160
rect -2000 32150 -1992 32197
rect -1942 32196 -1937 32198
rect -1932 32188 -1927 32196
rect -1912 32193 -1896 32199
rect -1842 32191 -1802 32202
rect -1671 32198 -1663 32206
rect -1663 32190 -1655 32198
rect -1850 32186 -1680 32190
rect -1924 32172 -1921 32174
rect -1806 32164 -1680 32170
rect -1671 32164 -1663 32178
rect -1663 32162 -1655 32164
rect -1854 32155 -1806 32160
rect -1974 32150 -1964 32151
rect -1960 32150 -1944 32152
rect -1842 32150 -1806 32153
rect -1655 32150 -1647 32162
rect -1642 32150 -1637 32244
rect -1619 32150 -1614 32244
rect -1530 32150 -1526 32244
rect -1506 32150 -1502 32244
rect -1482 32150 -1478 32244
rect -1458 32150 -1454 32244
rect -1434 32150 -1430 32244
rect -1410 32150 -1406 32244
rect -1386 32150 -1382 32244
rect -1362 32150 -1358 32244
rect -1338 32150 -1334 32244
rect -1314 32150 -1310 32244
rect -1290 32150 -1286 32244
rect -1266 32150 -1262 32244
rect -1242 32150 -1238 32244
rect -1218 32150 -1214 32244
rect -1194 32150 -1190 32244
rect -1170 32150 -1166 32244
rect -1146 32150 -1142 32244
rect -1122 32150 -1118 32244
rect -1098 32150 -1094 32244
rect -1074 32150 -1070 32244
rect -1050 32150 -1046 32244
rect -1026 32150 -1022 32244
rect -1002 32150 -998 32244
rect -978 32150 -974 32244
rect -954 32150 -950 32244
rect -930 32150 -926 32244
rect -906 32150 -902 32244
rect -882 32150 -878 32244
rect -858 32150 -854 32244
rect -834 32150 -830 32244
rect -810 32150 -806 32244
rect -786 32151 -782 32244
rect -797 32150 -763 32151
rect -2393 32148 -763 32150
rect -2371 32126 -2366 32148
rect -2348 32126 -2343 32148
rect -2325 32136 -2317 32148
rect -2325 32126 -2320 32136
rect -2317 32134 -2309 32136
rect -2062 32135 -2032 32142
rect -2309 32126 -2301 32134
rect -2070 32128 -2062 32135
rect -2000 32130 -1992 32148
rect -1974 32146 -1944 32148
rect -1960 32145 -1944 32146
rect -1842 32144 -1806 32148
rect -1842 32137 -1798 32142
rect -1806 32135 -1798 32137
rect -1671 32136 -1663 32148
rect -1854 32133 -1842 32135
rect -1663 32134 -1655 32136
rect -2062 32126 -2036 32128
rect -2393 32124 -2036 32126
rect -2032 32126 -2012 32128
rect -2004 32126 -1974 32130
rect -1854 32128 -1806 32133
rect -1864 32126 -1796 32127
rect -1655 32126 -1647 32134
rect -1642 32126 -1637 32148
rect -1619 32126 -1614 32148
rect -1530 32126 -1526 32148
rect -1506 32126 -1502 32148
rect -1482 32126 -1478 32148
rect -1458 32126 -1454 32148
rect -1434 32126 -1430 32148
rect -1410 32126 -1406 32148
rect -1386 32126 -1382 32148
rect -1362 32126 -1358 32148
rect -1338 32126 -1334 32148
rect -1314 32126 -1310 32148
rect -1290 32126 -1286 32148
rect -1266 32126 -1262 32148
rect -1242 32126 -1238 32148
rect -1218 32126 -1214 32148
rect -1194 32126 -1190 32148
rect -1170 32126 -1166 32148
rect -1146 32126 -1142 32148
rect -1122 32126 -1118 32148
rect -1098 32126 -1094 32148
rect -1074 32126 -1070 32148
rect -1050 32126 -1046 32148
rect -1026 32126 -1022 32148
rect -1002 32126 -998 32148
rect -978 32126 -974 32148
rect -954 32126 -950 32148
rect -930 32126 -926 32148
rect -906 32126 -902 32148
rect -882 32126 -878 32148
rect -858 32126 -854 32148
rect -834 32126 -830 32148
rect -810 32126 -806 32148
rect -797 32141 -792 32148
rect -786 32141 -782 32148
rect -787 32127 -782 32141
rect -786 32126 -782 32127
rect -762 32126 -758 32244
rect -738 32126 -734 32244
rect -714 32126 -710 32244
rect -690 32126 -686 32244
rect -666 32126 -662 32244
rect -642 32126 -638 32244
rect -618 32126 -614 32244
rect -594 32126 -590 32244
rect -570 32126 -566 32244
rect -546 32126 -542 32244
rect -522 32126 -518 32244
rect -498 32126 -494 32244
rect -474 32126 -470 32244
rect -450 32126 -446 32244
rect -426 32126 -422 32244
rect -402 32126 -398 32244
rect -378 32126 -374 32244
rect -354 32126 -350 32244
rect -330 32126 -326 32244
rect -306 32126 -302 32244
rect -282 32126 -278 32244
rect -258 32126 -254 32244
rect -234 32126 -230 32244
rect -210 32126 -206 32244
rect -186 32126 -182 32244
rect -173 32237 -168 32244
rect -162 32237 -158 32244
rect -163 32223 -158 32237
rect -162 32126 -158 32223
rect -138 32171 -134 32292
rect -138 32147 -131 32171
rect -138 32126 -134 32147
rect -114 32126 -110 32292
rect -90 32126 -86 32292
rect -66 32126 -62 32292
rect -42 32267 -38 32292
rect -42 32243 -35 32267
rect -42 32126 -38 32243
rect -18 32126 -14 32292
rect 6 32126 10 32292
rect 30 32126 34 32292
rect 54 32126 58 32292
rect 78 32126 82 32292
rect 102 32126 106 32292
rect 126 32126 130 32292
rect 150 32126 154 32292
rect 174 32126 178 32292
rect 198 32126 202 32292
rect 222 32126 226 32292
rect 246 32126 250 32292
rect 270 32126 274 32292
rect 277 32291 291 32292
rect 294 32291 301 32339
rect 294 32126 298 32291
rect 318 32126 322 32460
rect 342 32126 346 32460
rect 366 32126 370 32460
rect 390 32126 394 32460
rect 414 32319 418 32460
rect 403 32318 437 32319
rect 438 32318 442 32460
rect 462 32318 466 32460
rect 486 32318 490 32460
rect 510 32318 514 32460
rect 534 32318 538 32460
rect 558 32318 562 32460
rect 582 32318 586 32460
rect 606 32318 610 32460
rect 630 32318 634 32460
rect 637 32459 651 32460
rect 654 32459 661 32483
rect 654 32318 658 32459
rect 678 32318 682 32580
rect 702 32318 706 32580
rect 726 32318 730 32580
rect 750 32318 754 32580
rect 774 32318 778 32580
rect 798 32318 802 32580
rect 822 32318 826 32580
rect 846 32318 850 32580
rect 870 32318 874 32580
rect 894 32318 898 32580
rect 918 32318 922 32580
rect 942 32318 946 32580
rect 966 32318 970 32580
rect 990 32318 994 32580
rect 1014 32318 1018 32580
rect 1038 32555 1042 32580
rect 1038 32534 1045 32555
rect 1062 32534 1066 32580
rect 1086 32534 1090 32580
rect 1110 32534 1114 32580
rect 1134 32534 1138 32580
rect 1158 32534 1162 32580
rect 1182 32534 1186 32580
rect 1206 32534 1210 32580
rect 1230 32534 1234 32580
rect 1254 32534 1258 32580
rect 1278 32534 1282 32580
rect 1302 32534 1306 32580
rect 1326 32534 1330 32580
rect 1350 32534 1354 32580
rect 1374 32534 1378 32580
rect 1398 32534 1402 32580
rect 1422 32534 1426 32580
rect 1446 32534 1450 32580
rect 1470 32534 1474 32580
rect 1494 32534 1498 32580
rect 1518 32534 1522 32580
rect 1542 32534 1546 32580
rect 1566 32534 1570 32580
rect 1590 32534 1594 32580
rect 1614 32534 1618 32580
rect 1638 32534 1642 32580
rect 1662 32534 1666 32580
rect 1686 32534 1690 32580
rect 1710 32534 1714 32580
rect 1734 32534 1738 32580
rect 1747 32573 1752 32580
rect 1758 32573 1762 32580
rect 1757 32559 1762 32573
rect 1771 32569 1779 32573
rect 1765 32559 1771 32569
rect 1747 32534 1779 32535
rect 1021 32532 1779 32534
rect 1021 32531 1035 32532
rect 1038 32507 1045 32532
rect 1038 32318 1042 32507
rect 1062 32318 1066 32532
rect 1086 32318 1090 32532
rect 1110 32318 1114 32532
rect 1134 32318 1138 32532
rect 1158 32318 1162 32532
rect 1182 32318 1186 32532
rect 1206 32318 1210 32532
rect 1230 32318 1234 32532
rect 1254 32318 1258 32532
rect 1278 32318 1282 32532
rect 1302 32318 1306 32532
rect 1326 32318 1330 32532
rect 1350 32318 1354 32532
rect 1374 32318 1378 32532
rect 1398 32318 1402 32532
rect 1422 32318 1426 32532
rect 1446 32318 1450 32532
rect 1470 32318 1474 32532
rect 1494 32318 1498 32532
rect 1518 32318 1522 32532
rect 1542 32318 1546 32532
rect 1566 32318 1570 32532
rect 1590 32318 1594 32532
rect 1614 32318 1618 32532
rect 1638 32318 1642 32532
rect 1662 32318 1666 32532
rect 1686 32318 1690 32532
rect 1710 32318 1714 32532
rect 1734 32318 1738 32532
rect 1747 32525 1752 32532
rect 1765 32531 1779 32532
rect 1757 32511 1762 32525
rect 1747 32453 1752 32463
rect 1758 32453 1762 32511
rect 1757 32439 1762 32453
rect 1771 32449 1779 32453
rect 1765 32439 1771 32449
rect 1747 32405 1752 32415
rect 1757 32391 1762 32405
rect 1758 32318 1762 32391
rect 1771 32318 1779 32319
rect 403 32316 1779 32318
rect 403 32309 408 32316
rect 414 32309 418 32316
rect 413 32295 418 32309
rect 403 32285 408 32295
rect 413 32271 418 32285
rect 414 32126 418 32271
rect 438 32243 442 32316
rect 438 32222 445 32243
rect 462 32222 466 32316
rect 486 32222 490 32316
rect 510 32222 514 32316
rect 534 32222 538 32316
rect 558 32222 562 32316
rect 582 32222 586 32316
rect 606 32222 610 32316
rect 630 32222 634 32316
rect 654 32222 658 32316
rect 678 32222 682 32316
rect 702 32222 706 32316
rect 726 32222 730 32316
rect 750 32222 754 32316
rect 774 32222 778 32316
rect 798 32222 802 32316
rect 822 32222 826 32316
rect 846 32222 850 32316
rect 870 32222 874 32316
rect 894 32222 898 32316
rect 918 32222 922 32316
rect 942 32222 946 32316
rect 966 32222 970 32316
rect 990 32222 994 32316
rect 1014 32222 1018 32316
rect 1038 32223 1042 32316
rect 1027 32222 1061 32223
rect 421 32220 1061 32222
rect 421 32219 435 32220
rect 438 32195 445 32220
rect 438 32126 442 32195
rect 462 32126 466 32220
rect 486 32126 490 32220
rect 510 32126 514 32220
rect 534 32126 538 32220
rect 558 32126 562 32220
rect 582 32126 586 32220
rect 606 32126 610 32220
rect 630 32126 634 32220
rect 654 32126 658 32220
rect 678 32126 682 32220
rect 702 32126 706 32220
rect 726 32126 730 32220
rect 750 32126 754 32220
rect 774 32126 778 32220
rect 798 32126 802 32220
rect 822 32126 826 32220
rect 846 32126 850 32220
rect 870 32126 874 32220
rect 894 32126 898 32220
rect 918 32126 922 32220
rect 942 32126 946 32220
rect 966 32126 970 32220
rect 990 32126 994 32220
rect 1003 32189 1008 32199
rect 1014 32189 1018 32220
rect 1027 32213 1032 32220
rect 1038 32213 1042 32220
rect 1037 32199 1042 32213
rect 1013 32175 1018 32189
rect 1003 32165 1008 32175
rect 1013 32151 1018 32165
rect 1014 32126 1018 32151
rect 1038 32127 1042 32199
rect 1062 32147 1066 32316
rect 1027 32126 1059 32127
rect -2032 32124 1059 32126
rect -2371 32054 -2366 32124
rect -2348 32054 -2343 32124
rect -2325 32120 -2320 32124
rect -2309 32122 -2301 32124
rect -2317 32120 -2309 32122
rect -2325 32108 -2317 32120
rect -2052 32118 -2036 32120
rect -2052 32116 -2032 32118
rect -2062 32110 -2032 32116
rect -2325 32054 -2320 32108
rect -2317 32106 -2309 32108
rect -2092 32094 -2062 32096
rect -2094 32090 -2062 32094
rect -2309 32060 -2301 32066
rect -2317 32054 -2309 32060
rect -2000 32054 -1992 32124
rect -1904 32117 -1874 32124
rect -1842 32117 -1806 32124
rect -1655 32122 -1647 32124
rect -1663 32120 -1655 32122
rect -1842 32110 -1680 32116
rect -1671 32108 -1663 32120
rect -1663 32106 -1655 32108
rect -1854 32094 -1806 32096
rect -1854 32090 -1680 32094
rect -1655 32060 -1647 32066
rect -1663 32054 -1655 32060
rect -1642 32054 -1637 32124
rect -1619 32054 -1614 32124
rect -1530 32054 -1526 32124
rect -1506 32054 -1502 32124
rect -1482 32054 -1478 32124
rect -1458 32054 -1454 32124
rect -1434 32054 -1430 32124
rect -1410 32054 -1406 32124
rect -1386 32054 -1382 32124
rect -1362 32054 -1358 32124
rect -1338 32054 -1334 32124
rect -1314 32054 -1310 32124
rect -1290 32054 -1286 32124
rect -1266 32054 -1262 32124
rect -1242 32054 -1238 32124
rect -1218 32054 -1214 32124
rect -1194 32054 -1190 32124
rect -1170 32054 -1166 32124
rect -1146 32054 -1142 32124
rect -1122 32054 -1118 32124
rect -1098 32054 -1094 32124
rect -1074 32054 -1070 32124
rect -1050 32054 -1046 32124
rect -1026 32054 -1022 32124
rect -1002 32054 -998 32124
rect -978 32054 -974 32124
rect -954 32054 -950 32124
rect -930 32054 -926 32124
rect -906 32054 -902 32124
rect -882 32054 -878 32124
rect -858 32054 -854 32124
rect -834 32054 -830 32124
rect -810 32054 -806 32124
rect -786 32054 -782 32124
rect -762 32075 -758 32124
rect -2393 32052 -765 32054
rect -2371 31838 -2366 32052
rect -2348 31838 -2343 32052
rect -2325 31990 -2320 32052
rect -2317 32050 -2309 32052
rect -2000 32051 -1966 32052
rect -2000 32050 -1982 32051
rect -1663 32050 -1655 32052
rect -2028 32042 -2018 32044
rect -2309 32032 -2301 32038
rect -2091 32032 -2061 32039
rect -2317 32022 -2309 32032
rect -2044 32030 -2028 32032
rect -2026 32030 -2014 32042
rect -2084 32024 -2061 32030
rect -2044 32028 -2014 32030
rect -2292 32014 -2054 32023
rect -2325 31982 -2317 31990
rect -2325 31962 -2320 31982
rect -2317 31974 -2309 31982
rect -2325 31946 -2317 31962
rect -2325 31930 -2320 31946
rect -2309 31934 -2301 31946
rect -2317 31930 -2309 31934
rect -2103 31930 -2096 31932
rect -2083 31930 -2053 31932
rect -2325 31918 -2317 31930
rect -2103 31921 -2053 31930
rect -2018 31928 -2017 31934
rect -2003 31928 -2002 31930
rect -2026 31924 -2017 31928
rect -2325 31902 -2320 31918
rect -2309 31906 -2301 31918
rect -2017 31914 -2012 31924
rect -2317 31902 -2309 31906
rect -2325 31890 -2317 31902
rect -2325 31870 -2320 31890
rect -2325 31862 -2317 31870
rect -2325 31842 -2320 31862
rect -2317 31854 -2309 31862
rect -2325 31838 -2317 31842
rect -2000 31838 -1992 32050
rect -1982 32049 -1966 32050
rect -1980 32032 -1932 32039
rect -1655 32032 -1647 32038
rect -1846 32014 -1680 32023
rect -1663 32022 -1655 32032
rect -1671 31982 -1663 31990
rect -1663 31974 -1655 31982
rect -1671 31946 -1663 31962
rect -1655 31934 -1647 31946
rect -1972 31930 -1924 31932
rect -1663 31930 -1655 31934
rect -1972 31921 -1922 31930
rect -1671 31918 -1663 31930
rect -1655 31906 -1647 31918
rect -1663 31902 -1655 31906
rect -1671 31890 -1663 31902
rect -1671 31862 -1663 31870
rect -1663 31854 -1655 31862
rect -1926 31838 -1892 31841
rect -1671 31838 -1663 31842
rect -1642 31838 -1637 32052
rect -1619 31838 -1614 32052
rect -1530 31838 -1526 32052
rect -1506 31838 -1502 32052
rect -1482 31838 -1478 32052
rect -1458 31838 -1454 32052
rect -1434 31838 -1430 32052
rect -1410 31838 -1406 32052
rect -1386 31838 -1382 32052
rect -1362 31838 -1358 32052
rect -1338 31838 -1334 32052
rect -1314 31838 -1310 32052
rect -1290 31838 -1286 32052
rect -1266 31838 -1262 32052
rect -1242 31838 -1238 32052
rect -1218 31838 -1214 32052
rect -1194 31838 -1190 32052
rect -1170 31959 -1166 32052
rect -1181 31958 -1147 31959
rect -1146 31958 -1142 32052
rect -1122 31958 -1118 32052
rect -1098 31958 -1094 32052
rect -1074 31958 -1070 32052
rect -1050 31958 -1046 32052
rect -1026 31958 -1022 32052
rect -1002 31958 -998 32052
rect -978 31958 -974 32052
rect -954 31958 -950 32052
rect -930 31958 -926 32052
rect -906 31958 -902 32052
rect -882 31958 -878 32052
rect -858 31958 -854 32052
rect -834 31958 -830 32052
rect -810 31958 -806 32052
rect -786 31958 -782 32052
rect -779 32051 -765 32052
rect -762 32051 -755 32075
rect -762 31958 -758 32051
rect -738 31958 -734 32124
rect -714 31958 -710 32124
rect -690 31958 -686 32124
rect -666 31958 -662 32124
rect -642 31958 -638 32124
rect -618 31958 -614 32124
rect -594 31958 -590 32124
rect -570 31958 -566 32124
rect -546 31958 -542 32124
rect -522 31958 -518 32124
rect -509 31997 -504 32007
rect -498 31997 -494 32124
rect -499 31983 -494 31997
rect -498 31958 -494 31983
rect -474 31958 -470 32124
rect -450 31958 -446 32124
rect -426 31958 -422 32124
rect -402 31958 -398 32124
rect -378 31958 -374 32124
rect -354 31958 -350 32124
rect -330 31958 -326 32124
rect -306 31958 -302 32124
rect -282 31958 -278 32124
rect -258 31958 -254 32124
rect -234 31958 -230 32124
rect -210 31958 -206 32124
rect -186 31958 -182 32124
rect -162 31958 -158 32124
rect -138 31958 -134 32124
rect -114 31958 -110 32124
rect -90 31958 -86 32124
rect -66 31958 -62 32124
rect -42 31958 -38 32124
rect -18 31958 -14 32124
rect 6 31958 10 32124
rect 30 31958 34 32124
rect 54 31958 58 32124
rect 78 31958 82 32124
rect 102 31958 106 32124
rect 126 31958 130 32124
rect 150 31958 154 32124
rect 174 31958 178 32124
rect 198 31958 202 32124
rect 222 31958 226 32124
rect 246 31958 250 32124
rect 270 31958 274 32124
rect 294 31958 298 32124
rect 318 31958 322 32124
rect 342 31958 346 32124
rect 366 31958 370 32124
rect 390 31958 394 32124
rect 414 31958 418 32124
rect 438 31958 442 32124
rect 462 31958 466 32124
rect 486 31958 490 32124
rect 510 31958 514 32124
rect 534 31958 538 32124
rect 558 31958 562 32124
rect 582 31958 586 32124
rect 606 31958 610 32124
rect 630 31958 634 32124
rect 654 31958 658 32124
rect 678 31958 682 32124
rect 702 31958 706 32124
rect 726 31958 730 32124
rect 750 31958 754 32124
rect 774 31958 778 32124
rect 798 31958 802 32124
rect 822 31958 826 32124
rect 846 31958 850 32124
rect 870 31958 874 32124
rect 894 31958 898 32124
rect 918 31958 922 32124
rect 942 31958 946 32124
rect 966 31958 970 32124
rect 990 31958 994 32124
rect 1014 31958 1018 32124
rect 1027 32117 1032 32124
rect 1038 32123 1042 32124
rect 1045 32123 1059 32124
rect 1062 32123 1069 32147
rect 1038 32117 1045 32123
rect 1037 32103 1045 32117
rect 1038 32075 1045 32103
rect 1038 31958 1042 32075
rect 1062 32051 1066 32123
rect 1062 32027 1069 32051
rect 1062 31958 1066 32027
rect 1086 31958 1090 32316
rect 1110 31958 1114 32316
rect 1123 32069 1128 32079
rect 1134 32069 1138 32316
rect 1133 32055 1138 32069
rect 1123 32045 1128 32055
rect 1133 32031 1138 32045
rect 1134 31958 1138 32031
rect 1158 32003 1162 32316
rect -1181 31956 1155 31958
rect -1181 31949 -1176 31956
rect -1170 31949 -1166 31956
rect -1171 31935 -1166 31949
rect -1181 31925 -1176 31935
rect -1171 31911 -1166 31925
rect -1170 31838 -1166 31911
rect -1146 31883 -1142 31956
rect -2393 31836 -1149 31838
rect -2371 31790 -2366 31836
rect -2348 31790 -2343 31836
rect -2325 31830 -2317 31836
rect -2053 31834 -1972 31836
rect -2325 31814 -2320 31830
rect -2317 31826 -2309 31830
rect -2069 31826 -2068 31827
rect -2309 31814 -2301 31826
rect -2069 31819 -2038 31826
rect -2069 31817 -2068 31819
rect -2000 31818 -1992 31834
rect -1926 31831 -1924 31836
rect -1916 31828 -1914 31831
rect -1671 31830 -1663 31836
rect -1982 31818 -1916 31827
rect -1663 31826 -1655 31830
rect -2325 31802 -2317 31814
rect -2068 31811 -2053 31817
rect -2027 31816 -1992 31818
rect -2076 31802 -2053 31809
rect -2011 31808 -2002 31816
rect -2000 31808 -1992 31816
rect -1655 31814 -1647 31826
rect -2003 31806 -1992 31808
rect -2325 31790 -2320 31802
rect -2317 31798 -2309 31802
rect -2309 31790 -2301 31798
rect -2015 31794 -2003 31806
rect -2000 31790 -1992 31806
rect -1972 31802 -1924 31809
rect -1862 31801 -1680 31810
rect -1671 31802 -1663 31814
rect -1663 31798 -1655 31802
rect -1976 31790 -1940 31791
rect -1655 31790 -1647 31798
rect -1642 31790 -1637 31836
rect -1619 31790 -1614 31836
rect -1530 31790 -1526 31836
rect -1506 31790 -1502 31836
rect -1482 31790 -1478 31836
rect -1458 31790 -1454 31836
rect -1434 31790 -1430 31836
rect -1410 31791 -1406 31836
rect -1421 31790 -1387 31791
rect -2393 31788 -1387 31790
rect -2371 31694 -2366 31788
rect -2348 31694 -2343 31788
rect -2325 31786 -2320 31788
rect -2309 31786 -2301 31788
rect -2325 31774 -2317 31786
rect -2325 31754 -2320 31774
rect -2317 31770 -2309 31774
rect -2325 31746 -2317 31754
rect -2060 31748 -2030 31751
rect -2325 31694 -2320 31746
rect -2317 31738 -2309 31746
rect -2060 31735 -2038 31746
rect -2033 31739 -2030 31748
rect -2028 31744 -2027 31748
rect -2068 31730 -2038 31733
rect -2309 31698 -2301 31706
rect -2317 31694 -2309 31698
rect -2000 31694 -1992 31788
rect -1655 31786 -1647 31788
rect -1671 31774 -1663 31786
rect -1663 31770 -1655 31774
rect -1912 31763 -1884 31765
rect -1852 31757 -1804 31761
rect -1844 31748 -1796 31751
rect -1671 31746 -1663 31754
rect -1844 31735 -1804 31746
rect -1663 31738 -1655 31746
rect -1852 31730 -1680 31734
rect -1655 31698 -1647 31706
rect -1663 31694 -1655 31698
rect -1642 31694 -1637 31788
rect -1619 31694 -1614 31788
rect -1530 31694 -1526 31788
rect -1506 31694 -1502 31788
rect -1482 31694 -1478 31788
rect -1458 31694 -1454 31788
rect -1434 31694 -1430 31788
rect -1421 31781 -1416 31788
rect -1410 31781 -1406 31788
rect -1411 31767 -1406 31781
rect -1410 31694 -1406 31767
rect -1386 31715 -1382 31836
rect -2393 31692 -2020 31694
rect -2012 31692 -1389 31694
rect -2371 31358 -2366 31692
rect -2348 31358 -2343 31692
rect -2325 31630 -2320 31692
rect -2317 31690 -2309 31692
rect -2062 31679 -2061 31680
rect -2060 31679 -2049 31692
rect -2309 31670 -2301 31678
rect -2068 31672 -2061 31679
rect -2020 31672 -2012 31684
rect -2317 31662 -2309 31670
rect -2124 31663 -2108 31665
rect -2060 31663 -2049 31672
rect -2020 31670 -2004 31672
rect -2000 31670 -1992 31692
rect -1972 31690 -1958 31692
rect -1663 31690 -1655 31692
rect -1958 31689 -1942 31690
rect -1980 31672 -1932 31679
rect -1655 31670 -1647 31678
rect -2292 31662 -2049 31663
rect -2036 31662 -2030 31670
rect -2020 31668 -1992 31670
rect -2292 31655 -2030 31662
rect -2292 31654 -2049 31655
rect -2031 31654 -2030 31655
rect -2026 31654 -2020 31660
rect -2325 31622 -2317 31630
rect -2325 31602 -2320 31622
rect -2317 31614 -2309 31622
rect -2325 31586 -2317 31602
rect -2325 31570 -2320 31586
rect -2309 31574 -2301 31586
rect -2317 31570 -2309 31574
rect -2103 31570 -2096 31572
rect -2083 31570 -2053 31572
rect -2325 31558 -2317 31570
rect -2103 31561 -2053 31570
rect -2018 31568 -2017 31574
rect -2003 31568 -2002 31570
rect -2026 31564 -2017 31568
rect -2325 31542 -2320 31558
rect -2309 31546 -2301 31558
rect -2017 31554 -2012 31564
rect -2317 31542 -2309 31546
rect -2325 31530 -2317 31542
rect -2325 31510 -2320 31530
rect -2325 31502 -2317 31510
rect -2325 31482 -2320 31502
rect -2317 31494 -2309 31502
rect -2325 31466 -2317 31482
rect -2325 31450 -2320 31466
rect -2309 31454 -2301 31466
rect -2317 31450 -2309 31454
rect -2103 31450 -2096 31452
rect -2083 31450 -2053 31452
rect -2325 31438 -2317 31450
rect -2103 31441 -2053 31450
rect -2018 31448 -2017 31454
rect -2003 31448 -2002 31450
rect -2026 31444 -2017 31448
rect -2325 31422 -2320 31438
rect -2309 31426 -2301 31438
rect -2017 31434 -2012 31444
rect -2317 31422 -2309 31426
rect -2325 31410 -2317 31422
rect -2325 31390 -2320 31410
rect -2325 31382 -2317 31390
rect -2325 31362 -2320 31382
rect -2317 31374 -2309 31382
rect -2325 31358 -2317 31362
rect -2000 31358 -1992 31668
rect -1844 31654 -1680 31663
rect -1663 31662 -1655 31670
rect -1671 31622 -1663 31630
rect -1663 31614 -1655 31622
rect -1671 31586 -1663 31602
rect -1655 31574 -1647 31586
rect -1972 31570 -1924 31572
rect -1663 31570 -1655 31574
rect -1972 31561 -1922 31570
rect -1671 31558 -1663 31570
rect -1655 31546 -1647 31558
rect -1663 31542 -1655 31546
rect -1671 31530 -1663 31542
rect -1671 31502 -1663 31510
rect -1663 31494 -1655 31502
rect -1671 31466 -1663 31482
rect -1655 31454 -1647 31466
rect -1972 31450 -1924 31452
rect -1663 31450 -1655 31454
rect -1972 31441 -1922 31450
rect -1671 31438 -1663 31450
rect -1655 31426 -1647 31438
rect -1663 31422 -1655 31426
rect -1671 31410 -1663 31422
rect -1671 31382 -1663 31390
rect -1663 31374 -1655 31382
rect -1671 31358 -1663 31362
rect -1642 31358 -1637 31692
rect -1619 31358 -1614 31692
rect -1530 31358 -1526 31692
rect -1506 31358 -1502 31692
rect -1482 31358 -1478 31692
rect -1458 31358 -1454 31692
rect -1434 31358 -1430 31692
rect -1410 31358 -1406 31692
rect -1403 31691 -1389 31692
rect -1386 31691 -1379 31715
rect -1386 31358 -1382 31691
rect -1362 31358 -1358 31836
rect -1338 31358 -1334 31836
rect -1314 31358 -1310 31836
rect -1290 31358 -1286 31836
rect -1266 31358 -1262 31836
rect -1242 31358 -1238 31836
rect -1218 31358 -1214 31836
rect -1194 31358 -1190 31836
rect -1170 31358 -1166 31836
rect -1163 31835 -1149 31836
rect -1146 31835 -1139 31883
rect -1157 31637 -1152 31647
rect -1146 31637 -1142 31835
rect -1147 31623 -1142 31637
rect -1146 31358 -1142 31623
rect -1122 31571 -1118 31956
rect -1122 31547 -1115 31571
rect -1122 31358 -1118 31547
rect -1098 31358 -1094 31956
rect -1074 31358 -1070 31956
rect -1050 31479 -1046 31956
rect -1061 31478 -1027 31479
rect -1026 31478 -1022 31956
rect -1002 31478 -998 31956
rect -978 31478 -974 31956
rect -954 31478 -950 31956
rect -930 31478 -926 31956
rect -906 31478 -902 31956
rect -882 31478 -878 31956
rect -858 31478 -854 31956
rect -834 31478 -830 31956
rect -810 31478 -806 31956
rect -786 31478 -782 31956
rect -762 31478 -758 31956
rect -738 31478 -734 31956
rect -714 31478 -710 31956
rect -690 31478 -686 31956
rect -666 31478 -662 31956
rect -642 31478 -638 31956
rect -618 31478 -614 31956
rect -594 31478 -590 31956
rect -570 31478 -566 31956
rect -546 31478 -542 31956
rect -522 31478 -518 31956
rect -498 31478 -494 31956
rect -474 31931 -470 31956
rect -474 31907 -467 31931
rect -474 31478 -470 31907
rect -450 31478 -446 31956
rect -426 31478 -422 31956
rect -402 31478 -398 31956
rect -378 31478 -374 31956
rect -354 31719 -350 31956
rect -365 31718 -331 31719
rect -330 31718 -326 31956
rect -306 31718 -302 31956
rect -282 31718 -278 31956
rect -258 31718 -254 31956
rect -234 31718 -230 31956
rect -210 31718 -206 31956
rect -186 31718 -182 31956
rect -162 31718 -158 31956
rect -138 31718 -134 31956
rect -114 31718 -110 31956
rect -90 31718 -86 31956
rect -66 31718 -62 31956
rect -42 31718 -38 31956
rect -18 31718 -14 31956
rect 6 31718 10 31956
rect 30 31718 34 31956
rect 54 31863 58 31956
rect 43 31862 77 31863
rect 78 31862 82 31956
rect 102 31862 106 31956
rect 126 31862 130 31956
rect 150 31862 154 31956
rect 163 31877 168 31887
rect 174 31877 178 31956
rect 173 31863 178 31877
rect 174 31862 178 31863
rect 198 31862 202 31956
rect 222 31862 226 31956
rect 246 31862 250 31956
rect 270 31862 274 31956
rect 294 31862 298 31956
rect 318 31862 322 31956
rect 342 31862 346 31956
rect 366 31862 370 31956
rect 390 31862 394 31956
rect 414 31862 418 31956
rect 438 31862 442 31956
rect 462 31862 466 31956
rect 486 31862 490 31956
rect 510 31862 514 31956
rect 534 31862 538 31956
rect 558 31862 562 31956
rect 582 31862 586 31956
rect 606 31862 610 31956
rect 630 31862 634 31956
rect 654 31862 658 31956
rect 678 31862 682 31956
rect 702 31862 706 31956
rect 726 31862 730 31956
rect 750 31862 754 31956
rect 774 31862 778 31956
rect 798 31862 802 31956
rect 822 31862 826 31956
rect 846 31862 850 31956
rect 870 31862 874 31956
rect 894 31862 898 31956
rect 918 31862 922 31956
rect 942 31862 946 31956
rect 966 31862 970 31956
rect 990 31862 994 31956
rect 1014 31862 1018 31956
rect 1038 31862 1042 31956
rect 1062 31862 1066 31956
rect 1086 31862 1090 31956
rect 1110 31862 1114 31956
rect 1134 31862 1138 31956
rect 1141 31955 1155 31956
rect 1158 31955 1165 32003
rect 1158 31862 1162 31955
rect 1182 31862 1186 32316
rect 1206 31862 1210 32316
rect 1230 31862 1234 32316
rect 1254 31862 1258 32316
rect 1278 31862 1282 32316
rect 1302 31862 1306 32316
rect 1326 31862 1330 32316
rect 1350 31862 1354 32316
rect 1374 31862 1378 32316
rect 1398 31862 1402 32316
rect 1422 31862 1426 32316
rect 1446 31862 1450 32316
rect 1470 31862 1474 32316
rect 1494 31862 1498 32316
rect 1518 31862 1522 32316
rect 1542 31862 1546 32316
rect 1566 31862 1570 32316
rect 1590 31862 1594 32316
rect 1614 31862 1618 32316
rect 1638 31862 1642 32316
rect 1662 31862 1666 32316
rect 1686 31862 1690 32316
rect 1710 31862 1714 32316
rect 1734 31862 1738 32316
rect 1758 31862 1762 32316
rect 1765 32315 1779 32316
rect 1771 32309 1776 32315
rect 1781 32295 1786 32309
rect 1782 31862 1786 32295
rect 1795 32189 1800 32199
rect 1805 32175 1810 32189
rect 1806 31862 1810 32175
rect 1819 32069 1824 32079
rect 1829 32055 1834 32069
rect 1830 31862 1834 32055
rect 1843 31949 1848 31959
rect 1853 31935 1858 31949
rect 1854 31862 1858 31935
rect 1867 31862 1875 31863
rect 43 31860 1875 31862
rect 43 31853 48 31860
rect 54 31853 58 31860
rect 53 31839 58 31853
rect 43 31829 48 31839
rect 53 31815 58 31829
rect 54 31718 58 31815
rect 78 31787 82 31860
rect 78 31766 85 31787
rect 102 31766 106 31860
rect 126 31766 130 31860
rect 150 31766 154 31860
rect 174 31766 178 31860
rect 198 31811 202 31860
rect 198 31787 205 31811
rect 198 31766 202 31787
rect 222 31766 226 31860
rect 246 31766 250 31860
rect 270 31766 274 31860
rect 294 31766 298 31860
rect 318 31766 322 31860
rect 342 31766 346 31860
rect 366 31766 370 31860
rect 390 31766 394 31860
rect 414 31766 418 31860
rect 438 31766 442 31860
rect 462 31766 466 31860
rect 486 31766 490 31860
rect 510 31766 514 31860
rect 534 31766 538 31860
rect 558 31766 562 31860
rect 582 31766 586 31860
rect 606 31766 610 31860
rect 630 31766 634 31860
rect 654 31766 658 31860
rect 678 31766 682 31860
rect 702 31766 706 31860
rect 726 31766 730 31860
rect 750 31766 754 31860
rect 774 31766 778 31860
rect 798 31766 802 31860
rect 822 31766 826 31860
rect 846 31766 850 31860
rect 870 31766 874 31860
rect 894 31766 898 31860
rect 918 31766 922 31860
rect 942 31766 946 31860
rect 966 31767 970 31860
rect 955 31766 989 31767
rect 61 31764 989 31766
rect 61 31763 75 31764
rect 78 31739 85 31764
rect 78 31718 82 31739
rect 102 31718 106 31764
rect 126 31718 130 31764
rect 150 31718 154 31764
rect 174 31718 178 31764
rect 198 31718 202 31764
rect 222 31718 226 31764
rect 246 31718 250 31764
rect 270 31718 274 31764
rect 294 31718 298 31764
rect 318 31718 322 31764
rect 342 31718 346 31764
rect 366 31718 370 31764
rect 390 31718 394 31764
rect 414 31718 418 31764
rect 438 31718 442 31764
rect 462 31718 466 31764
rect 486 31718 490 31764
rect 510 31718 514 31764
rect 534 31718 538 31764
rect 558 31718 562 31764
rect 582 31718 586 31764
rect 606 31718 610 31764
rect 630 31718 634 31764
rect 654 31718 658 31764
rect 678 31718 682 31764
rect 702 31718 706 31764
rect 726 31718 730 31764
rect 750 31718 754 31764
rect 774 31718 778 31764
rect 798 31718 802 31764
rect 822 31718 826 31764
rect 846 31718 850 31764
rect 870 31718 874 31764
rect 894 31718 898 31764
rect 918 31718 922 31764
rect 942 31718 946 31764
rect 955 31757 960 31764
rect 966 31757 970 31764
rect 965 31743 970 31757
rect 966 31718 970 31743
rect 990 31718 994 31860
rect 1014 31718 1018 31860
rect 1038 31718 1042 31860
rect 1062 31718 1066 31860
rect 1086 31718 1090 31860
rect 1110 31718 1114 31860
rect 1134 31718 1138 31860
rect 1158 31718 1162 31860
rect 1182 31718 1186 31860
rect 1206 31718 1210 31860
rect 1230 31718 1234 31860
rect 1254 31718 1258 31860
rect 1278 31718 1282 31860
rect 1302 31718 1306 31860
rect 1326 31718 1330 31860
rect 1350 31718 1354 31860
rect 1374 31718 1378 31860
rect 1387 31805 1392 31815
rect 1398 31805 1402 31860
rect 1397 31791 1402 31805
rect 1398 31718 1402 31791
rect 1422 31739 1426 31860
rect -365 31716 1419 31718
rect -365 31709 -360 31716
rect -354 31709 -350 31716
rect -355 31695 -350 31709
rect -365 31685 -360 31695
rect -355 31671 -350 31685
rect -354 31478 -350 31671
rect -330 31643 -326 31716
rect -330 31595 -323 31643
rect -330 31478 -326 31595
rect -317 31517 -312 31527
rect -306 31517 -302 31716
rect -307 31503 -302 31517
rect -306 31478 -302 31503
rect -282 31478 -278 31716
rect -258 31478 -254 31716
rect -234 31478 -230 31716
rect -210 31478 -206 31716
rect -186 31478 -182 31716
rect -162 31478 -158 31716
rect -138 31478 -134 31716
rect -114 31478 -110 31716
rect -90 31478 -86 31716
rect -66 31478 -62 31716
rect -42 31478 -38 31716
rect -18 31478 -14 31716
rect 6 31478 10 31716
rect 30 31478 34 31716
rect 54 31478 58 31716
rect 78 31478 82 31716
rect 102 31478 106 31716
rect 126 31478 130 31716
rect 150 31478 154 31716
rect 174 31478 178 31716
rect 198 31478 202 31716
rect 222 31478 226 31716
rect 246 31478 250 31716
rect 270 31478 274 31716
rect 294 31478 298 31716
rect 318 31478 322 31716
rect 342 31478 346 31716
rect 366 31478 370 31716
rect 390 31478 394 31716
rect 414 31478 418 31716
rect 438 31478 442 31716
rect 462 31478 466 31716
rect 486 31478 490 31716
rect 510 31478 514 31716
rect 534 31478 538 31716
rect 558 31478 562 31716
rect 582 31478 586 31716
rect 606 31478 610 31716
rect 630 31478 634 31716
rect 654 31478 658 31716
rect 678 31478 682 31716
rect 702 31478 706 31716
rect 726 31478 730 31716
rect 750 31478 754 31716
rect 774 31478 778 31716
rect 798 31478 802 31716
rect 822 31478 826 31716
rect 835 31589 840 31599
rect 846 31589 850 31716
rect 845 31575 850 31589
rect 835 31565 840 31575
rect 845 31551 850 31565
rect 846 31478 850 31551
rect 870 31523 874 31716
rect -1061 31476 867 31478
rect -1061 31469 -1056 31476
rect -1050 31469 -1046 31476
rect -1051 31455 -1046 31469
rect -1061 31445 -1056 31455
rect -1051 31431 -1046 31445
rect -1050 31358 -1046 31431
rect -1026 31403 -1022 31476
rect -2393 31356 -1029 31358
rect -2371 31310 -2366 31356
rect -2348 31310 -2343 31356
rect -2325 31350 -2317 31356
rect -2018 31354 -2004 31356
rect -2325 31334 -2320 31350
rect -2317 31346 -2309 31350
rect -2069 31348 -2053 31350
rect -2309 31334 -2301 31346
rect -2096 31337 -2095 31343
rect -2000 31338 -1992 31356
rect -1671 31350 -1663 31356
rect -1663 31346 -1655 31350
rect -1977 31339 -1929 31345
rect -2112 31334 -2095 31337
rect -2325 31322 -2317 31334
rect -2325 31310 -2320 31322
rect -2317 31318 -2309 31322
rect -2112 31321 -2096 31334
rect -2059 31330 -2053 31337
rect -2027 31336 -1992 31338
rect -2059 31326 -2045 31330
rect -2018 31328 -2017 31330
rect -2083 31321 -2053 31322
rect -2019 31320 -2017 31324
rect -2309 31310 -2301 31318
rect -2017 31314 -2009 31320
rect -2000 31314 -1992 31336
rect -1972 31322 -1929 31337
rect -1655 31334 -1647 31346
rect -1671 31322 -1663 31334
rect -1972 31321 -1924 31322
rect -1663 31318 -1655 31322
rect -2033 31310 -1992 31314
rect -1655 31310 -1647 31318
rect -1642 31310 -1637 31356
rect -1619 31310 -1614 31356
rect -1530 31311 -1526 31356
rect -1541 31310 -1507 31311
rect -2393 31308 -1507 31310
rect -2371 31214 -2366 31308
rect -2348 31214 -2343 31308
rect -2325 31306 -2320 31308
rect -2309 31306 -2301 31308
rect -2325 31294 -2317 31306
rect -2325 31274 -2320 31294
rect -2317 31290 -2309 31294
rect -2325 31266 -2317 31274
rect -2325 31214 -2320 31266
rect -2317 31258 -2309 31266
rect -2117 31257 -2095 31267
rect -2045 31264 -2037 31278
rect -2309 31218 -2301 31228
rect -2087 31224 -2076 31232
rect -2017 31228 -2015 31235
rect -2317 31214 -2309 31218
rect -2092 31216 -2087 31224
rect -2092 31214 -2077 31215
rect -2000 31214 -1992 31308
rect -1655 31306 -1647 31308
rect -1671 31294 -1663 31306
rect -1663 31290 -1655 31294
rect -1969 31257 -1929 31269
rect -1671 31266 -1663 31274
rect -1663 31258 -1655 31266
rect -1655 31218 -1647 31228
rect -1928 31214 -1924 31215
rect -1854 31214 -1680 31215
rect -1663 31214 -1655 31218
rect -1642 31214 -1637 31308
rect -1619 31214 -1614 31308
rect -1541 31301 -1536 31308
rect -1530 31301 -1526 31308
rect -1531 31287 -1526 31301
rect -1530 31214 -1526 31287
rect -1506 31235 -1502 31356
rect -2393 31212 -1509 31214
rect -2371 31190 -2366 31212
rect -2348 31190 -2343 31212
rect -2325 31190 -2320 31212
rect -2092 31207 -2037 31212
rect -2021 31207 -1969 31212
rect -1921 31207 -1913 31212
rect -1854 31208 -1680 31212
rect -2100 31205 -2092 31206
rect -2309 31190 -2301 31200
rect -2100 31199 -2087 31205
rect -2051 31192 -2026 31194
rect -2062 31190 -2012 31192
rect -2000 31190 -1992 31207
rect -1969 31199 -1921 31206
rect -1969 31190 -1964 31199
rect -1864 31190 -1796 31191
rect -1655 31190 -1647 31200
rect -1642 31190 -1637 31212
rect -1619 31190 -1614 31212
rect -1530 31190 -1526 31212
rect -1523 31211 -1509 31212
rect -1506 31211 -1499 31235
rect -1506 31190 -1502 31211
rect -1482 31190 -1478 31356
rect -1458 31190 -1454 31356
rect -1434 31190 -1430 31356
rect -1410 31190 -1406 31356
rect -1386 31190 -1382 31356
rect -1362 31190 -1358 31356
rect -1338 31190 -1334 31356
rect -1314 31190 -1310 31356
rect -1290 31190 -1286 31356
rect -1266 31190 -1262 31356
rect -1242 31190 -1238 31356
rect -1218 31190 -1214 31356
rect -1194 31190 -1190 31356
rect -1170 31190 -1166 31356
rect -1146 31190 -1142 31356
rect -1122 31190 -1118 31356
rect -1098 31190 -1094 31356
rect -1074 31190 -1070 31356
rect -1050 31190 -1046 31356
rect -1043 31355 -1029 31356
rect -1026 31355 -1019 31403
rect -1026 31190 -1022 31355
rect -1002 31190 -998 31476
rect -978 31190 -974 31476
rect -954 31190 -950 31476
rect -930 31190 -926 31476
rect -906 31190 -902 31476
rect -893 31397 -888 31407
rect -882 31397 -878 31476
rect -883 31383 -878 31397
rect -882 31190 -878 31383
rect -858 31331 -854 31476
rect -858 31307 -851 31331
rect -858 31190 -854 31307
rect -834 31190 -830 31476
rect -810 31190 -806 31476
rect -786 31190 -782 31476
rect -762 31190 -758 31476
rect -738 31190 -734 31476
rect -714 31190 -710 31476
rect -690 31190 -686 31476
rect -666 31190 -662 31476
rect -642 31191 -638 31476
rect -653 31190 -619 31191
rect -2393 31188 -619 31190
rect -2371 31142 -2366 31188
rect -2348 31142 -2343 31188
rect -2325 31142 -2320 31188
rect -2317 31184 -2309 31188
rect -2105 31181 -2092 31184
rect -2092 31158 -2062 31160
rect -2094 31154 -2062 31158
rect -2000 31142 -1992 31188
rect -1663 31184 -1655 31188
rect -1969 31181 -1921 31184
rect -1854 31158 -1806 31160
rect -1854 31154 -1680 31158
rect -1642 31142 -1637 31188
rect -1619 31142 -1614 31188
rect -1530 31142 -1526 31188
rect -1506 31142 -1502 31188
rect -1482 31142 -1478 31188
rect -1458 31142 -1454 31188
rect -1434 31142 -1430 31188
rect -1410 31142 -1406 31188
rect -1386 31142 -1382 31188
rect -1362 31142 -1358 31188
rect -1338 31142 -1334 31188
rect -1314 31142 -1310 31188
rect -1290 31142 -1286 31188
rect -1266 31142 -1262 31188
rect -1242 31142 -1238 31188
rect -1218 31142 -1214 31188
rect -1194 31142 -1190 31188
rect -1170 31142 -1166 31188
rect -1146 31142 -1142 31188
rect -1122 31142 -1118 31188
rect -1098 31142 -1094 31188
rect -1074 31142 -1070 31188
rect -1050 31142 -1046 31188
rect -1026 31142 -1022 31188
rect -1002 31142 -998 31188
rect -978 31142 -974 31188
rect -954 31142 -950 31188
rect -930 31142 -926 31188
rect -906 31142 -902 31188
rect -882 31142 -878 31188
rect -858 31142 -854 31188
rect -834 31142 -830 31188
rect -810 31142 -806 31188
rect -786 31142 -782 31188
rect -762 31142 -758 31188
rect -738 31142 -734 31188
rect -714 31142 -710 31188
rect -690 31142 -686 31188
rect -666 31142 -662 31188
rect -653 31181 -648 31188
rect -642 31181 -638 31188
rect -643 31167 -638 31181
rect -642 31142 -638 31167
rect -618 31142 -614 31476
rect -594 31142 -590 31476
rect -581 31205 -576 31215
rect -570 31205 -566 31476
rect -571 31191 -566 31205
rect -570 31142 -566 31191
rect -546 31142 -542 31476
rect -522 31142 -518 31476
rect -498 31142 -494 31476
rect -474 31142 -470 31476
rect -450 31142 -446 31476
rect -426 31142 -422 31476
rect -402 31142 -398 31476
rect -378 31383 -374 31476
rect -389 31382 -355 31383
rect -354 31382 -350 31476
rect -330 31382 -326 31476
rect -306 31382 -302 31476
rect -282 31451 -278 31476
rect -282 31427 -275 31451
rect -282 31382 -278 31427
rect -258 31382 -254 31476
rect -234 31382 -230 31476
rect -210 31382 -206 31476
rect -186 31382 -182 31476
rect -162 31382 -158 31476
rect -138 31382 -134 31476
rect -114 31382 -110 31476
rect -90 31382 -86 31476
rect -66 31382 -62 31476
rect -42 31382 -38 31476
rect -18 31382 -14 31476
rect 6 31382 10 31476
rect 30 31382 34 31476
rect 54 31382 58 31476
rect 78 31382 82 31476
rect 102 31382 106 31476
rect 126 31382 130 31476
rect 150 31382 154 31476
rect 174 31382 178 31476
rect 198 31382 202 31476
rect 222 31382 226 31476
rect 246 31382 250 31476
rect 270 31382 274 31476
rect 294 31382 298 31476
rect 318 31382 322 31476
rect 342 31382 346 31476
rect 366 31382 370 31476
rect 390 31382 394 31476
rect 414 31382 418 31476
rect 438 31382 442 31476
rect 462 31382 466 31476
rect 486 31382 490 31476
rect 510 31382 514 31476
rect 534 31382 538 31476
rect 558 31382 562 31476
rect 582 31382 586 31476
rect 606 31382 610 31476
rect 630 31382 634 31476
rect 654 31382 658 31476
rect 678 31382 682 31476
rect 702 31382 706 31476
rect 726 31382 730 31476
rect 750 31382 754 31476
rect 774 31382 778 31476
rect 798 31382 802 31476
rect 822 31382 826 31476
rect 846 31382 850 31476
rect 853 31475 867 31476
rect 870 31475 877 31523
rect 870 31382 874 31475
rect 894 31382 898 31716
rect 918 31382 922 31716
rect 942 31382 946 31716
rect 966 31382 970 31716
rect 990 31691 994 31716
rect 990 31667 997 31691
rect 990 31382 994 31667
rect 1014 31382 1018 31716
rect 1038 31382 1042 31716
rect 1062 31382 1066 31716
rect 1086 31382 1090 31716
rect 1110 31382 1114 31716
rect 1134 31382 1138 31716
rect 1158 31382 1162 31716
rect 1182 31382 1186 31716
rect 1206 31382 1210 31716
rect 1230 31382 1234 31716
rect 1254 31382 1258 31716
rect 1278 31382 1282 31716
rect 1302 31382 1306 31716
rect 1326 31382 1330 31716
rect 1350 31382 1354 31716
rect 1374 31382 1378 31716
rect 1398 31382 1402 31716
rect 1405 31715 1419 31716
rect 1422 31715 1429 31739
rect 1422 31382 1426 31715
rect 1446 31382 1450 31860
rect 1470 31382 1474 31860
rect 1494 31382 1498 31860
rect 1518 31382 1522 31860
rect 1542 31382 1546 31860
rect 1566 31382 1570 31860
rect 1590 31382 1594 31860
rect 1614 31382 1618 31860
rect 1638 31382 1642 31860
rect 1662 31382 1666 31860
rect 1686 31382 1690 31860
rect 1710 31382 1714 31860
rect 1734 31382 1738 31860
rect 1758 31382 1762 31860
rect 1782 31382 1786 31860
rect 1806 31382 1810 31860
rect 1830 31382 1834 31860
rect 1854 31382 1858 31860
rect 1861 31859 1875 31860
rect 1867 31853 1872 31859
rect 1877 31839 1882 31853
rect 1878 31382 1882 31839
rect 1891 31709 1896 31719
rect 1901 31695 1906 31709
rect 1902 31382 1906 31695
rect 1915 31589 1920 31599
rect 1925 31575 1930 31589
rect 1926 31382 1930 31575
rect 1939 31469 1944 31479
rect 1949 31455 1954 31469
rect 1950 31382 1954 31455
rect 1963 31382 1971 31383
rect -389 31380 1971 31382
rect -389 31373 -384 31380
rect -378 31373 -374 31380
rect -379 31359 -374 31373
rect -389 31349 -384 31359
rect -379 31335 -374 31349
rect -378 31142 -374 31335
rect -354 31307 -350 31380
rect -354 31286 -347 31307
rect -330 31286 -326 31380
rect -306 31286 -302 31380
rect -282 31286 -278 31380
rect -258 31286 -254 31380
rect -234 31286 -230 31380
rect -210 31286 -206 31380
rect -186 31286 -182 31380
rect -162 31286 -158 31380
rect -138 31286 -134 31380
rect -114 31286 -110 31380
rect -90 31286 -86 31380
rect -66 31286 -62 31380
rect -42 31286 -38 31380
rect -18 31286 -14 31380
rect 6 31286 10 31380
rect 30 31286 34 31380
rect 54 31286 58 31380
rect 78 31286 82 31380
rect 102 31286 106 31380
rect 126 31286 130 31380
rect 150 31286 154 31380
rect 174 31286 178 31380
rect 198 31286 202 31380
rect 222 31286 226 31380
rect 246 31286 250 31380
rect 270 31286 274 31380
rect 294 31286 298 31380
rect 318 31286 322 31380
rect 342 31286 346 31380
rect 366 31286 370 31380
rect 390 31286 394 31380
rect 414 31286 418 31380
rect 438 31286 442 31380
rect 462 31286 466 31380
rect 486 31286 490 31380
rect 510 31286 514 31380
rect 534 31286 538 31380
rect 558 31286 562 31380
rect 582 31286 586 31380
rect 606 31286 610 31380
rect 630 31286 634 31380
rect 654 31286 658 31380
rect 678 31286 682 31380
rect 702 31286 706 31380
rect 726 31286 730 31380
rect 750 31286 754 31380
rect 774 31286 778 31380
rect 798 31286 802 31380
rect 822 31286 826 31380
rect 846 31286 850 31380
rect 870 31286 874 31380
rect 894 31286 898 31380
rect 918 31286 922 31380
rect 942 31286 946 31380
rect 966 31286 970 31380
rect 990 31286 994 31380
rect 1014 31286 1018 31380
rect 1038 31286 1042 31380
rect 1062 31286 1066 31380
rect 1086 31286 1090 31380
rect 1110 31286 1114 31380
rect 1134 31286 1138 31380
rect 1158 31286 1162 31380
rect 1182 31286 1186 31380
rect 1206 31286 1210 31380
rect 1230 31286 1234 31380
rect 1254 31286 1258 31380
rect 1278 31286 1282 31380
rect 1302 31286 1306 31380
rect 1326 31286 1330 31380
rect 1350 31286 1354 31380
rect 1374 31286 1378 31380
rect 1398 31286 1402 31380
rect 1422 31286 1426 31380
rect 1446 31286 1450 31380
rect 1470 31286 1474 31380
rect 1494 31286 1498 31380
rect 1518 31286 1522 31380
rect 1542 31286 1546 31380
rect 1566 31286 1570 31380
rect 1590 31286 1594 31380
rect 1614 31286 1618 31380
rect 1638 31286 1642 31380
rect 1662 31286 1666 31380
rect 1686 31286 1690 31380
rect 1710 31286 1714 31380
rect 1734 31286 1738 31380
rect 1758 31286 1762 31380
rect 1782 31286 1786 31380
rect 1806 31286 1810 31380
rect 1830 31286 1834 31380
rect 1854 31286 1858 31380
rect 1878 31286 1882 31380
rect 1902 31286 1906 31380
rect 1926 31286 1930 31380
rect 1950 31286 1954 31380
rect 1957 31379 1971 31380
rect 1963 31373 1968 31379
rect 1973 31359 1978 31373
rect 1974 31287 1978 31359
rect 1963 31286 1995 31287
rect -371 31284 1995 31286
rect -371 31283 -357 31284
rect -354 31259 -347 31284
rect -354 31142 -350 31259
rect -330 31142 -326 31284
rect -306 31142 -302 31284
rect -282 31142 -278 31284
rect -258 31142 -254 31284
rect -234 31142 -230 31284
rect -221 31253 -216 31263
rect -210 31253 -206 31284
rect -211 31239 -206 31253
rect -221 31229 -216 31239
rect -211 31215 -206 31229
rect -210 31142 -206 31215
rect -186 31187 -182 31284
rect -2393 31140 -189 31142
rect -2371 31118 -2366 31140
rect -2348 31118 -2343 31140
rect -2325 31118 -2320 31140
rect -2072 31138 -2036 31139
rect -2072 31132 -2054 31138
rect -2309 31124 -2301 31132
rect -2317 31118 -2309 31124
rect -2092 31123 -2062 31128
rect -2000 31119 -1992 31140
rect -1938 31139 -1906 31140
rect -1920 31138 -1906 31139
rect -1806 31132 -1680 31138
rect -1854 31123 -1806 31128
rect -1655 31124 -1647 31132
rect -1982 31119 -1966 31120
rect -2000 31118 -1966 31119
rect -1846 31118 -1806 31121
rect -1663 31118 -1655 31124
rect -1642 31118 -1637 31140
rect -1619 31118 -1614 31140
rect -1530 31118 -1526 31140
rect -1506 31118 -1502 31140
rect -1482 31118 -1478 31140
rect -1458 31118 -1454 31140
rect -1434 31118 -1430 31140
rect -1410 31118 -1406 31140
rect -1386 31118 -1382 31140
rect -1362 31118 -1358 31140
rect -1338 31118 -1334 31140
rect -1314 31118 -1310 31140
rect -1290 31118 -1286 31140
rect -1266 31118 -1262 31140
rect -1242 31118 -1238 31140
rect -1218 31118 -1214 31140
rect -1194 31118 -1190 31140
rect -1170 31118 -1166 31140
rect -1146 31118 -1142 31140
rect -1122 31118 -1118 31140
rect -1098 31118 -1094 31140
rect -1074 31118 -1070 31140
rect -1050 31118 -1046 31140
rect -1026 31118 -1022 31140
rect -1002 31118 -998 31140
rect -978 31118 -974 31140
rect -954 31118 -950 31140
rect -930 31118 -926 31140
rect -906 31118 -902 31140
rect -882 31118 -878 31140
rect -858 31118 -854 31140
rect -834 31118 -830 31140
rect -810 31118 -806 31140
rect -786 31118 -782 31140
rect -762 31118 -758 31140
rect -738 31118 -734 31140
rect -714 31118 -710 31140
rect -690 31118 -686 31140
rect -666 31118 -662 31140
rect -642 31118 -638 31140
rect -618 31118 -614 31140
rect -594 31118 -590 31140
rect -570 31118 -566 31140
rect -546 31139 -542 31140
rect -2393 31116 -549 31118
rect -2371 31094 -2366 31116
rect -2348 31094 -2343 31116
rect -2325 31094 -2320 31116
rect -2000 31114 -1966 31116
rect -2309 31096 -2301 31104
rect -2062 31103 -2054 31110
rect -2092 31096 -2084 31103
rect -2062 31096 -2026 31098
rect -2317 31094 -2309 31096
rect -2062 31094 -2012 31096
rect -2000 31094 -1992 31114
rect -1982 31113 -1966 31114
rect -1846 31112 -1806 31116
rect -1846 31105 -1798 31110
rect -1806 31103 -1798 31105
rect -1854 31101 -1846 31103
rect -1854 31096 -1806 31101
rect -1655 31096 -1647 31104
rect -1864 31094 -1796 31095
rect -1663 31094 -1655 31096
rect -1642 31094 -1637 31116
rect -1619 31094 -1614 31116
rect -1530 31094 -1526 31116
rect -1506 31094 -1502 31116
rect -1482 31094 -1478 31116
rect -1458 31094 -1454 31116
rect -1434 31094 -1430 31116
rect -1410 31094 -1406 31116
rect -1386 31094 -1382 31116
rect -1362 31094 -1358 31116
rect -1338 31094 -1334 31116
rect -1314 31094 -1310 31116
rect -1290 31094 -1286 31116
rect -1266 31094 -1262 31116
rect -1242 31094 -1238 31116
rect -1218 31094 -1214 31116
rect -1194 31094 -1190 31116
rect -1170 31094 -1166 31116
rect -1146 31094 -1142 31116
rect -1122 31094 -1118 31116
rect -1098 31094 -1094 31116
rect -1074 31094 -1070 31116
rect -1050 31094 -1046 31116
rect -1026 31094 -1022 31116
rect -1002 31094 -998 31116
rect -978 31094 -974 31116
rect -954 31094 -950 31116
rect -930 31094 -926 31116
rect -906 31094 -902 31116
rect -882 31094 -878 31116
rect -858 31094 -854 31116
rect -834 31094 -830 31116
rect -810 31094 -806 31116
rect -786 31094 -782 31116
rect -762 31094 -758 31116
rect -738 31094 -734 31116
rect -714 31094 -710 31116
rect -690 31094 -686 31116
rect -666 31094 -662 31116
rect -642 31094 -638 31116
rect -618 31115 -614 31116
rect -2393 31092 -621 31094
rect -2371 31046 -2366 31092
rect -2348 31046 -2343 31092
rect -2325 31046 -2320 31092
rect -2317 31088 -2309 31092
rect -2062 31088 -2054 31092
rect -2154 31084 -2138 31086
rect -2057 31084 -2054 31088
rect -2292 31078 -2054 31084
rect -2052 31078 -2044 31088
rect -2092 31062 -2062 31064
rect -2094 31058 -2062 31062
rect -2000 31046 -1992 31092
rect -1846 31085 -1806 31092
rect -1663 31088 -1655 31092
rect -1846 31078 -1680 31084
rect -1854 31062 -1806 31064
rect -1854 31058 -1680 31062
rect -1642 31046 -1637 31092
rect -1619 31046 -1614 31092
rect -1530 31046 -1526 31092
rect -1506 31046 -1502 31092
rect -1482 31046 -1478 31092
rect -1458 31046 -1454 31092
rect -1434 31046 -1430 31092
rect -1410 31046 -1406 31092
rect -1386 31046 -1382 31092
rect -1362 31046 -1358 31092
rect -1338 31046 -1334 31092
rect -1314 31046 -1310 31092
rect -1290 31046 -1286 31092
rect -1266 31046 -1262 31092
rect -1242 31046 -1238 31092
rect -1218 31046 -1214 31092
rect -1194 31046 -1190 31092
rect -1170 31046 -1166 31092
rect -1146 31046 -1142 31092
rect -1122 31046 -1118 31092
rect -1098 31046 -1094 31092
rect -1074 31046 -1070 31092
rect -1050 31046 -1046 31092
rect -1026 31046 -1022 31092
rect -1002 31046 -998 31092
rect -978 31046 -974 31092
rect -954 31046 -950 31092
rect -930 31046 -926 31092
rect -906 31046 -902 31092
rect -882 31046 -878 31092
rect -858 31046 -854 31092
rect -834 31046 -830 31092
rect -810 31046 -806 31092
rect -786 31046 -782 31092
rect -762 31046 -758 31092
rect -738 31046 -734 31092
rect -714 31046 -710 31092
rect -690 31046 -686 31092
rect -666 31046 -662 31092
rect -642 31046 -638 31092
rect -635 31091 -621 31092
rect -618 31091 -611 31115
rect -618 31046 -614 31091
rect -594 31046 -590 31116
rect -570 31046 -566 31116
rect -563 31115 -549 31116
rect -546 31115 -539 31139
rect -546 31046 -542 31115
rect -522 31046 -518 31140
rect -498 31046 -494 31140
rect -474 31046 -470 31140
rect -450 31046 -446 31140
rect -426 31046 -422 31140
rect -402 31046 -398 31140
rect -378 31046 -374 31140
rect -354 31046 -350 31140
rect -330 31046 -326 31140
rect -306 31046 -302 31140
rect -282 31046 -278 31140
rect -258 31046 -254 31140
rect -234 31046 -230 31140
rect -210 31046 -206 31140
rect -203 31139 -189 31140
rect -186 31139 -179 31187
rect -186 31046 -182 31139
rect -162 31046 -158 31284
rect -138 31046 -134 31284
rect -114 31046 -110 31284
rect -90 31046 -86 31284
rect -66 31046 -62 31284
rect -42 31046 -38 31284
rect -18 31046 -14 31284
rect 6 31046 10 31284
rect 30 31046 34 31284
rect 54 31046 58 31284
rect 78 31046 82 31284
rect 102 31046 106 31284
rect 126 31046 130 31284
rect 150 31046 154 31284
rect 174 31046 178 31284
rect 198 31046 202 31284
rect 222 31046 226 31284
rect 246 31046 250 31284
rect 270 31046 274 31284
rect 294 31046 298 31284
rect 318 31046 322 31284
rect 342 31046 346 31284
rect 366 31046 370 31284
rect 390 31046 394 31284
rect 414 31046 418 31284
rect 438 31046 442 31284
rect 462 31046 466 31284
rect 486 31046 490 31284
rect 510 31046 514 31284
rect 534 31046 538 31284
rect 558 31046 562 31284
rect 582 31046 586 31284
rect 606 31046 610 31284
rect 630 31046 634 31284
rect 654 31046 658 31284
rect 678 31046 682 31284
rect 702 31046 706 31284
rect 726 31046 730 31284
rect 750 31046 754 31284
rect 774 31046 778 31284
rect 798 31046 802 31284
rect 822 31046 826 31284
rect 846 31046 850 31284
rect 870 31046 874 31284
rect 894 31167 898 31284
rect 883 31166 917 31167
rect 918 31166 922 31284
rect 942 31166 946 31284
rect 966 31166 970 31284
rect 990 31166 994 31284
rect 1014 31166 1018 31284
rect 1038 31166 1042 31284
rect 1062 31166 1066 31284
rect 1086 31166 1090 31284
rect 1110 31166 1114 31284
rect 1134 31166 1138 31284
rect 1158 31166 1162 31284
rect 1182 31166 1186 31284
rect 1206 31166 1210 31284
rect 1230 31166 1234 31284
rect 1254 31166 1258 31284
rect 1278 31166 1282 31284
rect 1302 31166 1306 31284
rect 1326 31166 1330 31284
rect 1350 31166 1354 31284
rect 1374 31166 1378 31284
rect 1398 31166 1402 31284
rect 1422 31166 1426 31284
rect 1446 31166 1450 31284
rect 1470 31166 1474 31284
rect 1494 31166 1498 31284
rect 1518 31166 1522 31284
rect 1542 31166 1546 31284
rect 1566 31166 1570 31284
rect 1590 31166 1594 31284
rect 1614 31166 1618 31284
rect 1638 31166 1642 31284
rect 1662 31166 1666 31284
rect 1686 31166 1690 31284
rect 1710 31166 1714 31284
rect 1734 31166 1738 31284
rect 1758 31166 1762 31284
rect 1782 31166 1786 31284
rect 1806 31166 1810 31284
rect 1830 31166 1834 31284
rect 1854 31166 1858 31284
rect 1878 31166 1882 31284
rect 1902 31166 1906 31284
rect 1926 31166 1930 31284
rect 1950 31166 1954 31284
rect 1963 31277 1968 31284
rect 1974 31277 1978 31284
rect 1981 31283 1995 31284
rect 1973 31263 1978 31277
rect 1963 31253 1968 31263
rect 1973 31239 1978 31253
rect 1974 31166 1978 31239
rect 1987 31166 1995 31167
rect 883 31164 1995 31166
rect 883 31157 888 31164
rect 894 31157 898 31164
rect 893 31143 898 31157
rect 883 31133 888 31143
rect 893 31119 898 31133
rect 894 31046 898 31119
rect 918 31091 922 31164
rect -2393 31044 915 31046
rect -2371 31022 -2366 31044
rect -2348 31022 -2343 31044
rect -2325 31022 -2320 31044
rect -2072 31042 -2036 31043
rect -2072 31036 -2054 31042
rect -2309 31028 -2301 31036
rect -2317 31022 -2309 31028
rect -2092 31027 -2062 31032
rect -2000 31023 -1992 31044
rect -1938 31043 -1906 31044
rect -1920 31042 -1906 31043
rect -1806 31036 -1680 31042
rect -1854 31027 -1806 31032
rect -1655 31028 -1647 31036
rect -1982 31023 -1966 31024
rect -2000 31022 -1966 31023
rect -1846 31022 -1806 31025
rect -1663 31022 -1655 31028
rect -1642 31022 -1637 31044
rect -1619 31022 -1614 31044
rect -1530 31022 -1526 31044
rect -1506 31022 -1502 31044
rect -1482 31022 -1478 31044
rect -1458 31022 -1454 31044
rect -1434 31022 -1430 31044
rect -1410 31022 -1406 31044
rect -1386 31022 -1382 31044
rect -1362 31022 -1358 31044
rect -1338 31022 -1334 31044
rect -1314 31022 -1310 31044
rect -1290 31022 -1286 31044
rect -1266 31022 -1262 31044
rect -1242 31022 -1238 31044
rect -1218 31022 -1214 31044
rect -1194 31022 -1190 31044
rect -1170 31022 -1166 31044
rect -1146 31022 -1142 31044
rect -1122 31022 -1118 31044
rect -1098 31022 -1094 31044
rect -1074 31022 -1070 31044
rect -1050 31022 -1046 31044
rect -1026 31022 -1022 31044
rect -1002 31022 -998 31044
rect -978 31022 -974 31044
rect -954 31022 -950 31044
rect -930 31022 -926 31044
rect -906 31022 -902 31044
rect -882 31022 -878 31044
rect -858 31022 -854 31044
rect -834 31022 -830 31044
rect -810 31022 -806 31044
rect -786 31022 -782 31044
rect -762 31022 -758 31044
rect -738 31022 -734 31044
rect -714 31022 -710 31044
rect -690 31022 -686 31044
rect -666 31022 -662 31044
rect -642 31022 -638 31044
rect -618 31022 -614 31044
rect -594 31022 -590 31044
rect -570 31022 -566 31044
rect -546 31022 -542 31044
rect -522 31022 -518 31044
rect -498 31022 -494 31044
rect -474 31022 -470 31044
rect -450 31022 -446 31044
rect -426 31022 -422 31044
rect -402 31022 -398 31044
rect -378 31022 -374 31044
rect -354 31022 -350 31044
rect -330 31022 -326 31044
rect -306 31022 -302 31044
rect -282 31022 -278 31044
rect -258 31022 -254 31044
rect -234 31022 -230 31044
rect -210 31022 -206 31044
rect -186 31022 -182 31044
rect -162 31022 -158 31044
rect -138 31022 -134 31044
rect -114 31022 -110 31044
rect -90 31022 -86 31044
rect -66 31022 -62 31044
rect -42 31022 -38 31044
rect -18 31022 -14 31044
rect 6 31022 10 31044
rect 30 31022 34 31044
rect 54 31022 58 31044
rect 78 31022 82 31044
rect 102 31022 106 31044
rect 126 31022 130 31044
rect 150 31022 154 31044
rect 174 31022 178 31044
rect 198 31022 202 31044
rect 222 31022 226 31044
rect 246 31022 250 31044
rect 270 31022 274 31044
rect 294 31022 298 31044
rect 318 31022 322 31044
rect 342 31022 346 31044
rect 366 31022 370 31044
rect 390 31022 394 31044
rect 414 31022 418 31044
rect 438 31022 442 31044
rect 462 31022 466 31044
rect 486 31023 490 31044
rect 475 31022 509 31023
rect -2393 31020 509 31022
rect -2371 30998 -2366 31020
rect -2348 30998 -2343 31020
rect -2325 30998 -2320 31020
rect -2000 31018 -1966 31020
rect -2309 31000 -2301 31008
rect -2062 31007 -2054 31014
rect -2092 31000 -2084 31007
rect -2062 31000 -2026 31002
rect -2317 30998 -2309 31000
rect -2062 30998 -2012 31000
rect -2000 30998 -1992 31018
rect -1982 31017 -1966 31018
rect -1846 31016 -1806 31020
rect -1846 31009 -1798 31014
rect -1806 31007 -1798 31009
rect -1854 31005 -1846 31007
rect -1854 31000 -1806 31005
rect -1655 31000 -1647 31008
rect -1864 30998 -1796 30999
rect -1663 30998 -1655 31000
rect -1642 30998 -1637 31020
rect -1619 30998 -1614 31020
rect -1530 30998 -1526 31020
rect -1506 30998 -1502 31020
rect -1482 30998 -1478 31020
rect -1458 30998 -1454 31020
rect -1434 30998 -1430 31020
rect -1410 30998 -1406 31020
rect -1386 30998 -1382 31020
rect -1362 30998 -1358 31020
rect -1338 30998 -1334 31020
rect -1314 30998 -1310 31020
rect -1290 30998 -1286 31020
rect -1266 30998 -1262 31020
rect -1242 30998 -1238 31020
rect -1218 30998 -1214 31020
rect -1194 30998 -1190 31020
rect -1170 30998 -1166 31020
rect -1146 30998 -1142 31020
rect -1122 30998 -1118 31020
rect -1098 30998 -1094 31020
rect -1074 30998 -1070 31020
rect -1050 30998 -1046 31020
rect -1026 30998 -1022 31020
rect -1002 30998 -998 31020
rect -978 30998 -974 31020
rect -954 30998 -950 31020
rect -930 30998 -926 31020
rect -906 30998 -902 31020
rect -882 30998 -878 31020
rect -858 30998 -854 31020
rect -834 30998 -830 31020
rect -810 30998 -806 31020
rect -786 30998 -782 31020
rect -762 30998 -758 31020
rect -738 30998 -734 31020
rect -714 30998 -710 31020
rect -690 30998 -686 31020
rect -666 30998 -662 31020
rect -642 30998 -638 31020
rect -618 30998 -614 31020
rect -594 30998 -590 31020
rect -570 30998 -566 31020
rect -546 30998 -542 31020
rect -522 30998 -518 31020
rect -498 30998 -494 31020
rect -474 30998 -470 31020
rect -450 30998 -446 31020
rect -426 30998 -422 31020
rect -402 30998 -398 31020
rect -378 30998 -374 31020
rect -354 30998 -350 31020
rect -330 30998 -326 31020
rect -306 30998 -302 31020
rect -282 30998 -278 31020
rect -258 30998 -254 31020
rect -234 30998 -230 31020
rect -210 30998 -206 31020
rect -186 30998 -182 31020
rect -162 30998 -158 31020
rect -138 30998 -134 31020
rect -114 30998 -110 31020
rect -90 30998 -86 31020
rect -66 30998 -62 31020
rect -42 30998 -38 31020
rect -18 30998 -14 31020
rect 6 30998 10 31020
rect 30 30998 34 31020
rect 54 30998 58 31020
rect 78 30998 82 31020
rect 102 30998 106 31020
rect 126 30998 130 31020
rect 150 30998 154 31020
rect 174 30998 178 31020
rect 198 30998 202 31020
rect 222 30998 226 31020
rect 246 30998 250 31020
rect 270 30998 274 31020
rect 294 30998 298 31020
rect 318 30998 322 31020
rect 342 30998 346 31020
rect 366 30998 370 31020
rect 390 30998 394 31020
rect 414 30998 418 31020
rect 438 30998 442 31020
rect 462 30998 466 31020
rect 475 31013 480 31020
rect 486 31013 490 31020
rect 485 30999 490 31013
rect 486 30998 490 30999
rect 510 30998 514 31044
rect 534 30998 538 31044
rect 558 30998 562 31044
rect 582 30998 586 31044
rect 606 30998 610 31044
rect 630 30998 634 31044
rect 654 30998 658 31044
rect 678 30998 682 31044
rect 702 30998 706 31044
rect 726 30998 730 31044
rect 750 30998 754 31044
rect 774 30998 778 31044
rect 798 30998 802 31044
rect 822 30998 826 31044
rect 846 30998 850 31044
rect 870 30998 874 31044
rect 894 30998 898 31044
rect 901 31043 915 31044
rect 918 31043 925 31091
rect 918 30998 922 31043
rect 942 30998 946 31164
rect 966 30998 970 31164
rect 990 30998 994 31164
rect 1014 30998 1018 31164
rect 1038 30998 1042 31164
rect 1062 30998 1066 31164
rect 1086 30998 1090 31164
rect 1110 30998 1114 31164
rect 1134 30998 1138 31164
rect 1158 30998 1162 31164
rect 1182 31071 1186 31164
rect 1171 31070 1205 31071
rect 1206 31070 1210 31164
rect 1230 31070 1234 31164
rect 1254 31070 1258 31164
rect 1278 31070 1282 31164
rect 1302 31070 1306 31164
rect 1326 31070 1330 31164
rect 1350 31070 1354 31164
rect 1374 31070 1378 31164
rect 1398 31070 1402 31164
rect 1422 31070 1426 31164
rect 1446 31070 1450 31164
rect 1470 31070 1474 31164
rect 1494 31070 1498 31164
rect 1518 31070 1522 31164
rect 1542 31070 1546 31164
rect 1566 31070 1570 31164
rect 1590 31070 1594 31164
rect 1614 31070 1618 31164
rect 1638 31070 1642 31164
rect 1662 31070 1666 31164
rect 1686 31070 1690 31164
rect 1710 31070 1714 31164
rect 1734 31070 1738 31164
rect 1758 31070 1762 31164
rect 1782 31070 1786 31164
rect 1806 31070 1810 31164
rect 1830 31070 1834 31164
rect 1854 31070 1858 31164
rect 1878 31070 1882 31164
rect 1902 31070 1906 31164
rect 1926 31070 1930 31164
rect 1950 31070 1954 31164
rect 1963 31085 1968 31095
rect 1974 31085 1978 31164
rect 1981 31163 1995 31164
rect 1987 31157 1992 31163
rect 1997 31143 2002 31157
rect 1987 31109 1992 31119
rect 1998 31109 2002 31143
rect 1997 31095 2002 31109
rect 1973 31071 1978 31085
rect 1963 31070 1997 31071
rect 1171 31068 1997 31070
rect 1171 31061 1176 31068
rect 1182 31061 1186 31068
rect 1181 31047 1186 31061
rect 1171 31037 1176 31047
rect 1181 31023 1186 31037
rect 1182 30998 1186 31023
rect 1206 30998 1210 31068
rect 1230 30998 1234 31068
rect 1254 30998 1258 31068
rect 1278 30998 1282 31068
rect 1302 30998 1306 31068
rect 1326 30998 1330 31068
rect 1350 30998 1354 31068
rect 1374 30998 1378 31068
rect 1398 30998 1402 31068
rect 1422 30998 1426 31068
rect 1446 30998 1450 31068
rect 1470 30998 1474 31068
rect 1494 30998 1498 31068
rect 1518 30998 1522 31068
rect 1542 30998 1546 31068
rect 1566 30998 1570 31068
rect 1590 30998 1594 31068
rect 1614 30998 1618 31068
rect 1638 30998 1642 31068
rect 1662 30998 1666 31068
rect 1686 30998 1690 31068
rect 1710 30998 1714 31068
rect 1734 30998 1738 31068
rect 1758 30998 1762 31068
rect 1782 30998 1786 31068
rect 1806 30998 1810 31068
rect 1830 30998 1834 31068
rect 1854 30998 1858 31068
rect 1878 30998 1882 31068
rect 1902 30998 1906 31068
rect 1926 30998 1930 31068
rect 1950 30998 1954 31068
rect 1963 31061 1968 31068
rect 1973 31047 1978 31061
rect 1974 30999 1978 31047
rect 1963 30998 1995 30999
rect -2393 30996 1995 30998
rect -2371 30950 -2366 30996
rect -2348 30950 -2343 30996
rect -2325 30950 -2320 30996
rect -2317 30992 -2309 30996
rect -2062 30992 -2054 30996
rect -2154 30988 -2138 30990
rect -2057 30988 -2054 30992
rect -2292 30982 -2054 30988
rect -2052 30982 -2044 30992
rect -2092 30966 -2062 30968
rect -2094 30962 -2062 30966
rect -2000 30950 -1992 30996
rect -1846 30989 -1806 30996
rect -1663 30992 -1655 30996
rect -1846 30982 -1680 30988
rect -1854 30966 -1806 30968
rect -1854 30962 -1680 30966
rect -1642 30950 -1637 30996
rect -1619 30950 -1614 30996
rect -1530 30950 -1526 30996
rect -1506 30950 -1502 30996
rect -1482 30950 -1478 30996
rect -1458 30950 -1454 30996
rect -1434 30950 -1430 30996
rect -1410 30950 -1406 30996
rect -1386 30950 -1382 30996
rect -1362 30950 -1358 30996
rect -1338 30950 -1334 30996
rect -1314 30950 -1310 30996
rect -1290 30950 -1286 30996
rect -1266 30950 -1262 30996
rect -1242 30950 -1238 30996
rect -1218 30950 -1214 30996
rect -1194 30950 -1190 30996
rect -1170 30950 -1166 30996
rect -1146 30950 -1142 30996
rect -1122 30950 -1118 30996
rect -1098 30950 -1094 30996
rect -1074 30950 -1070 30996
rect -1050 30950 -1046 30996
rect -1026 30950 -1022 30996
rect -1002 30950 -998 30996
rect -978 30950 -974 30996
rect -954 30950 -950 30996
rect -930 30950 -926 30996
rect -906 30950 -902 30996
rect -882 30950 -878 30996
rect -858 30950 -854 30996
rect -834 30950 -830 30996
rect -810 30950 -806 30996
rect -786 30950 -782 30996
rect -762 30950 -758 30996
rect -738 30950 -734 30996
rect -714 30950 -710 30996
rect -690 30950 -686 30996
rect -666 30950 -662 30996
rect -642 30950 -638 30996
rect -618 30950 -614 30996
rect -594 30950 -590 30996
rect -570 30950 -566 30996
rect -546 30950 -542 30996
rect -522 30950 -518 30996
rect -498 30950 -494 30996
rect -474 30950 -470 30996
rect -450 30950 -446 30996
rect -426 30950 -422 30996
rect -402 30950 -398 30996
rect -378 30950 -374 30996
rect -354 30950 -350 30996
rect -330 30950 -326 30996
rect -306 30950 -302 30996
rect -282 30950 -278 30996
rect -258 30950 -254 30996
rect -234 30950 -230 30996
rect -210 30950 -206 30996
rect -186 30950 -182 30996
rect -162 30950 -158 30996
rect -138 30950 -134 30996
rect -114 30950 -110 30996
rect -90 30950 -86 30996
rect -66 30950 -62 30996
rect -42 30950 -38 30996
rect -18 30950 -14 30996
rect 6 30950 10 30996
rect 30 30950 34 30996
rect 54 30950 58 30996
rect 78 30950 82 30996
rect 102 30950 106 30996
rect 126 30950 130 30996
rect 150 30950 154 30996
rect 174 30950 178 30996
rect 198 30950 202 30996
rect 222 30950 226 30996
rect 246 30950 250 30996
rect 270 30950 274 30996
rect 294 30950 298 30996
rect 318 30950 322 30996
rect 342 30950 346 30996
rect 366 30950 370 30996
rect 390 30950 394 30996
rect 414 30950 418 30996
rect 438 30950 442 30996
rect 462 30950 466 30996
rect 486 30950 490 30996
rect 510 30950 514 30996
rect 534 30950 538 30996
rect 558 30950 562 30996
rect 571 30965 576 30975
rect 582 30965 586 30996
rect 581 30951 586 30965
rect 571 30950 605 30951
rect -2393 30948 605 30950
rect -2371 30926 -2366 30948
rect -2348 30926 -2343 30948
rect -2325 30926 -2320 30948
rect -2072 30946 -2036 30947
rect -2072 30940 -2054 30946
rect -2309 30932 -2301 30940
rect -2317 30926 -2309 30932
rect -2092 30931 -2062 30936
rect -2000 30927 -1992 30948
rect -1938 30947 -1906 30948
rect -1920 30946 -1906 30947
rect -1806 30940 -1680 30946
rect -1854 30931 -1806 30936
rect -1655 30932 -1647 30940
rect -1982 30927 -1966 30928
rect -2000 30926 -1966 30927
rect -1846 30926 -1806 30929
rect -1663 30926 -1655 30932
rect -1642 30926 -1637 30948
rect -1619 30926 -1614 30948
rect -1530 30926 -1526 30948
rect -1506 30926 -1502 30948
rect -1482 30926 -1478 30948
rect -1458 30926 -1454 30948
rect -1434 30926 -1430 30948
rect -1410 30926 -1406 30948
rect -1386 30926 -1382 30948
rect -1362 30926 -1358 30948
rect -1338 30926 -1334 30948
rect -1314 30926 -1310 30948
rect -1290 30926 -1286 30948
rect -1266 30926 -1262 30948
rect -1242 30926 -1238 30948
rect -1218 30926 -1214 30948
rect -1194 30926 -1190 30948
rect -1170 30926 -1166 30948
rect -1146 30926 -1142 30948
rect -1122 30926 -1118 30948
rect -1098 30926 -1094 30948
rect -1074 30926 -1070 30948
rect -1050 30926 -1046 30948
rect -1026 30926 -1022 30948
rect -1002 30926 -998 30948
rect -978 30926 -974 30948
rect -954 30926 -950 30948
rect -930 30926 -926 30948
rect -906 30926 -902 30948
rect -882 30926 -878 30948
rect -858 30926 -854 30948
rect -834 30926 -830 30948
rect -810 30926 -806 30948
rect -786 30926 -782 30948
rect -762 30926 -758 30948
rect -738 30926 -734 30948
rect -714 30926 -710 30948
rect -690 30926 -686 30948
rect -666 30926 -662 30948
rect -642 30926 -638 30948
rect -618 30926 -614 30948
rect -594 30926 -590 30948
rect -570 30926 -566 30948
rect -546 30926 -542 30948
rect -522 30926 -518 30948
rect -498 30926 -494 30948
rect -474 30926 -470 30948
rect -450 30926 -446 30948
rect -426 30926 -422 30948
rect -402 30926 -398 30948
rect -378 30926 -374 30948
rect -354 30926 -350 30948
rect -330 30926 -326 30948
rect -306 30926 -302 30948
rect -282 30926 -278 30948
rect -258 30926 -254 30948
rect -234 30926 -230 30948
rect -210 30926 -206 30948
rect -186 30926 -182 30948
rect -162 30926 -158 30948
rect -138 30926 -134 30948
rect -114 30926 -110 30948
rect -90 30926 -86 30948
rect -66 30926 -62 30948
rect -42 30926 -38 30948
rect -18 30926 -14 30948
rect 6 30926 10 30948
rect 30 30926 34 30948
rect 54 30926 58 30948
rect 78 30926 82 30948
rect 102 30926 106 30948
rect 126 30926 130 30948
rect 150 30926 154 30948
rect 174 30926 178 30948
rect 198 30926 202 30948
rect 222 30926 226 30948
rect 246 30926 250 30948
rect 270 30926 274 30948
rect 294 30926 298 30948
rect 318 30926 322 30948
rect 342 30926 346 30948
rect 366 30926 370 30948
rect 390 30926 394 30948
rect 414 30926 418 30948
rect 438 30926 442 30948
rect 462 30926 466 30948
rect 486 30926 490 30948
rect 510 30947 514 30948
rect -2393 30924 507 30926
rect -2371 30902 -2366 30924
rect -2348 30902 -2343 30924
rect -2325 30902 -2320 30924
rect -2000 30922 -1966 30924
rect -2309 30904 -2301 30912
rect -2062 30911 -2054 30918
rect -2092 30904 -2084 30911
rect -2062 30904 -2026 30906
rect -2317 30902 -2309 30904
rect -2062 30902 -2012 30904
rect -2000 30902 -1992 30922
rect -1982 30921 -1966 30922
rect -1846 30920 -1806 30924
rect -1846 30913 -1798 30918
rect -1806 30911 -1798 30913
rect -1854 30909 -1846 30911
rect -1854 30904 -1806 30909
rect -1655 30904 -1647 30912
rect -1864 30902 -1796 30903
rect -1663 30902 -1655 30904
rect -1642 30902 -1637 30924
rect -1619 30902 -1614 30924
rect -1530 30902 -1526 30924
rect -1506 30902 -1502 30924
rect -1482 30902 -1478 30924
rect -1458 30902 -1454 30924
rect -1434 30902 -1430 30924
rect -1410 30902 -1406 30924
rect -1386 30902 -1382 30924
rect -1362 30902 -1358 30924
rect -1338 30902 -1334 30924
rect -1314 30902 -1310 30924
rect -1290 30902 -1286 30924
rect -1266 30902 -1262 30924
rect -1242 30902 -1238 30924
rect -1218 30902 -1214 30924
rect -1194 30902 -1190 30924
rect -1170 30902 -1166 30924
rect -1146 30902 -1142 30924
rect -1122 30902 -1118 30924
rect -1098 30902 -1094 30924
rect -1074 30902 -1070 30924
rect -1050 30902 -1046 30924
rect -1026 30902 -1022 30924
rect -1002 30902 -998 30924
rect -978 30902 -974 30924
rect -954 30902 -950 30924
rect -930 30902 -926 30924
rect -906 30902 -902 30924
rect -882 30902 -878 30924
rect -858 30902 -854 30924
rect -834 30902 -830 30924
rect -810 30902 -806 30924
rect -786 30902 -782 30924
rect -762 30902 -758 30924
rect -738 30902 -734 30924
rect -714 30902 -710 30924
rect -690 30902 -686 30924
rect -666 30902 -662 30924
rect -642 30902 -638 30924
rect -618 30902 -614 30924
rect -594 30902 -590 30924
rect -570 30902 -566 30924
rect -546 30902 -542 30924
rect -522 30902 -518 30924
rect -498 30902 -494 30924
rect -474 30902 -470 30924
rect -450 30902 -446 30924
rect -426 30902 -422 30924
rect -402 30902 -398 30924
rect -378 30902 -374 30924
rect -354 30902 -350 30924
rect -330 30902 -326 30924
rect -306 30902 -302 30924
rect -282 30902 -278 30924
rect -258 30902 -254 30924
rect -234 30902 -230 30924
rect -210 30902 -206 30924
rect -186 30902 -182 30924
rect -162 30902 -158 30924
rect -138 30902 -134 30924
rect -114 30902 -110 30924
rect -90 30902 -86 30924
rect -66 30902 -62 30924
rect -42 30902 -38 30924
rect -18 30902 -14 30924
rect 6 30902 10 30924
rect 30 30902 34 30924
rect 54 30902 58 30924
rect 78 30902 82 30924
rect 102 30902 106 30924
rect 126 30902 130 30924
rect 150 30902 154 30924
rect 174 30902 178 30924
rect 198 30902 202 30924
rect 222 30902 226 30924
rect 246 30902 250 30924
rect 270 30902 274 30924
rect 294 30902 298 30924
rect 318 30902 322 30924
rect 342 30902 346 30924
rect 366 30902 370 30924
rect 390 30902 394 30924
rect 414 30902 418 30924
rect 438 30902 442 30924
rect 462 30902 466 30924
rect 486 30902 490 30924
rect 493 30923 507 30924
rect 510 30923 517 30947
rect 510 30902 514 30923
rect 534 30902 538 30948
rect 558 30902 562 30948
rect 571 30941 576 30948
rect 581 30927 586 30941
rect 582 30902 586 30927
rect 606 30902 610 30996
rect 630 30903 634 30996
rect 619 30902 653 30903
rect -2393 30900 653 30902
rect -2371 30854 -2366 30900
rect -2348 30854 -2343 30900
rect -2325 30854 -2320 30900
rect -2317 30896 -2309 30900
rect -2062 30896 -2054 30900
rect -2154 30892 -2138 30894
rect -2057 30892 -2054 30896
rect -2292 30886 -2054 30892
rect -2052 30886 -2044 30896
rect -2092 30870 -2062 30872
rect -2094 30866 -2062 30870
rect -2000 30854 -1992 30900
rect -1846 30893 -1806 30900
rect -1663 30896 -1655 30900
rect -1846 30886 -1680 30892
rect -1854 30870 -1806 30872
rect -1854 30866 -1680 30870
rect -1642 30854 -1637 30900
rect -1619 30854 -1614 30900
rect -1530 30854 -1526 30900
rect -1506 30854 -1502 30900
rect -1482 30854 -1478 30900
rect -1458 30854 -1454 30900
rect -1434 30854 -1430 30900
rect -1410 30854 -1406 30900
rect -1386 30854 -1382 30900
rect -1362 30854 -1358 30900
rect -1338 30854 -1334 30900
rect -1314 30854 -1310 30900
rect -1290 30854 -1286 30900
rect -1266 30854 -1262 30900
rect -1242 30854 -1238 30900
rect -1218 30854 -1214 30900
rect -1194 30854 -1190 30900
rect -1170 30854 -1166 30900
rect -1146 30854 -1142 30900
rect -1122 30854 -1118 30900
rect -1098 30854 -1094 30900
rect -1074 30854 -1070 30900
rect -1050 30854 -1046 30900
rect -1026 30854 -1022 30900
rect -1002 30854 -998 30900
rect -978 30854 -974 30900
rect -954 30854 -950 30900
rect -930 30854 -926 30900
rect -906 30854 -902 30900
rect -882 30854 -878 30900
rect -858 30854 -854 30900
rect -834 30854 -830 30900
rect -810 30854 -806 30900
rect -786 30854 -782 30900
rect -762 30854 -758 30900
rect -738 30854 -734 30900
rect -714 30854 -710 30900
rect -690 30854 -686 30900
rect -666 30854 -662 30900
rect -642 30854 -638 30900
rect -618 30854 -614 30900
rect -594 30854 -590 30900
rect -570 30854 -566 30900
rect -546 30854 -542 30900
rect -522 30854 -518 30900
rect -498 30854 -494 30900
rect -474 30854 -470 30900
rect -450 30854 -446 30900
rect -426 30854 -422 30900
rect -402 30854 -398 30900
rect -378 30854 -374 30900
rect -354 30854 -350 30900
rect -330 30854 -326 30900
rect -306 30854 -302 30900
rect -282 30854 -278 30900
rect -258 30854 -254 30900
rect -234 30854 -230 30900
rect -210 30854 -206 30900
rect -186 30854 -182 30900
rect -162 30854 -158 30900
rect -138 30854 -134 30900
rect -114 30854 -110 30900
rect -90 30854 -86 30900
rect -66 30854 -62 30900
rect -42 30854 -38 30900
rect -18 30854 -14 30900
rect 6 30854 10 30900
rect 30 30854 34 30900
rect 54 30854 58 30900
rect 78 30854 82 30900
rect 102 30854 106 30900
rect 126 30854 130 30900
rect 150 30854 154 30900
rect 174 30854 178 30900
rect 198 30854 202 30900
rect 222 30854 226 30900
rect 246 30854 250 30900
rect 270 30854 274 30900
rect 294 30854 298 30900
rect 318 30854 322 30900
rect 342 30854 346 30900
rect 366 30854 370 30900
rect 390 30854 394 30900
rect 414 30854 418 30900
rect 438 30854 442 30900
rect 462 30854 466 30900
rect 486 30854 490 30900
rect 510 30854 514 30900
rect 534 30854 538 30900
rect 558 30854 562 30900
rect 582 30854 586 30900
rect 606 30899 610 30900
rect -2393 30852 603 30854
rect -2371 30830 -2366 30852
rect -2348 30830 -2343 30852
rect -2325 30830 -2320 30852
rect -2072 30850 -2036 30851
rect -2072 30844 -2054 30850
rect -2309 30836 -2301 30844
rect -2317 30830 -2309 30836
rect -2092 30835 -2062 30840
rect -2000 30831 -1992 30852
rect -1938 30851 -1906 30852
rect -1920 30850 -1906 30851
rect -1806 30844 -1680 30850
rect -1854 30835 -1806 30840
rect -1655 30836 -1647 30844
rect -1982 30831 -1966 30832
rect -2000 30830 -1966 30831
rect -1846 30830 -1806 30833
rect -1663 30830 -1655 30836
rect -1642 30830 -1637 30852
rect -1619 30830 -1614 30852
rect -1530 30830 -1526 30852
rect -1506 30830 -1502 30852
rect -1482 30830 -1478 30852
rect -1458 30830 -1454 30852
rect -1434 30830 -1430 30852
rect -1410 30830 -1406 30852
rect -1386 30830 -1382 30852
rect -1362 30830 -1358 30852
rect -1338 30830 -1334 30852
rect -1314 30830 -1310 30852
rect -1290 30830 -1286 30852
rect -1266 30830 -1262 30852
rect -1242 30830 -1238 30852
rect -1218 30830 -1214 30852
rect -1194 30830 -1190 30852
rect -1170 30830 -1166 30852
rect -1146 30830 -1142 30852
rect -1122 30830 -1118 30852
rect -1098 30830 -1094 30852
rect -1074 30830 -1070 30852
rect -1050 30830 -1046 30852
rect -1026 30830 -1022 30852
rect -1002 30830 -998 30852
rect -978 30830 -974 30852
rect -954 30830 -950 30852
rect -930 30830 -926 30852
rect -906 30830 -902 30852
rect -882 30830 -878 30852
rect -858 30830 -854 30852
rect -834 30830 -830 30852
rect -810 30830 -806 30852
rect -786 30830 -782 30852
rect -762 30830 -758 30852
rect -738 30830 -734 30852
rect -714 30830 -710 30852
rect -690 30830 -686 30852
rect -666 30830 -662 30852
rect -642 30830 -638 30852
rect -618 30830 -614 30852
rect -594 30830 -590 30852
rect -570 30830 -566 30852
rect -546 30830 -542 30852
rect -522 30830 -518 30852
rect -498 30830 -494 30852
rect -474 30830 -470 30852
rect -450 30831 -446 30852
rect -461 30830 -427 30831
rect -2393 30828 -427 30830
rect -2371 30806 -2366 30828
rect -2348 30806 -2343 30828
rect -2325 30806 -2320 30828
rect -2000 30826 -1966 30828
rect -2309 30808 -2301 30816
rect -2062 30815 -2054 30822
rect -2092 30808 -2084 30815
rect -2062 30808 -2026 30810
rect -2317 30806 -2309 30808
rect -2062 30806 -2012 30808
rect -2000 30806 -1992 30826
rect -1982 30825 -1966 30826
rect -1846 30824 -1806 30828
rect -1846 30817 -1798 30822
rect -1806 30815 -1798 30817
rect -1854 30813 -1846 30815
rect -1854 30808 -1806 30813
rect -1655 30808 -1647 30816
rect -1864 30806 -1796 30807
rect -1663 30806 -1655 30808
rect -1642 30806 -1637 30828
rect -1619 30806 -1614 30828
rect -1530 30806 -1526 30828
rect -1506 30806 -1502 30828
rect -1482 30806 -1478 30828
rect -1458 30806 -1454 30828
rect -1434 30806 -1430 30828
rect -1410 30806 -1406 30828
rect -1386 30806 -1382 30828
rect -1362 30806 -1358 30828
rect -1338 30806 -1334 30828
rect -1314 30806 -1310 30828
rect -1290 30806 -1286 30828
rect -1266 30806 -1262 30828
rect -1242 30806 -1238 30828
rect -1218 30806 -1214 30828
rect -1194 30806 -1190 30828
rect -1170 30806 -1166 30828
rect -1146 30806 -1142 30828
rect -1122 30806 -1118 30828
rect -1098 30806 -1094 30828
rect -1074 30806 -1070 30828
rect -1050 30806 -1046 30828
rect -1026 30806 -1022 30828
rect -1002 30806 -998 30828
rect -978 30806 -974 30828
rect -954 30806 -950 30828
rect -930 30806 -926 30828
rect -906 30806 -902 30828
rect -882 30806 -878 30828
rect -858 30806 -854 30828
rect -834 30806 -830 30828
rect -810 30806 -806 30828
rect -786 30806 -782 30828
rect -762 30806 -758 30828
rect -738 30806 -734 30828
rect -714 30806 -710 30828
rect -690 30806 -686 30828
rect -666 30806 -662 30828
rect -642 30806 -638 30828
rect -618 30806 -614 30828
rect -594 30806 -590 30828
rect -570 30806 -566 30828
rect -546 30806 -542 30828
rect -522 30806 -518 30828
rect -498 30806 -494 30828
rect -474 30806 -470 30828
rect -461 30821 -456 30828
rect -450 30821 -446 30828
rect -451 30807 -446 30821
rect -450 30806 -446 30807
rect -426 30806 -422 30852
rect -402 30806 -398 30852
rect -378 30806 -374 30852
rect -354 30806 -350 30852
rect -330 30806 -326 30852
rect -306 30806 -302 30852
rect -282 30806 -278 30852
rect -258 30806 -254 30852
rect -234 30806 -230 30852
rect -210 30806 -206 30852
rect -186 30806 -182 30852
rect -162 30806 -158 30852
rect -138 30806 -134 30852
rect -114 30806 -110 30852
rect -90 30806 -86 30852
rect -66 30806 -62 30852
rect -42 30806 -38 30852
rect -18 30806 -14 30852
rect 6 30806 10 30852
rect 30 30806 34 30852
rect 54 30806 58 30852
rect 78 30806 82 30852
rect 102 30806 106 30852
rect 126 30806 130 30852
rect 150 30806 154 30852
rect 174 30806 178 30852
rect 198 30806 202 30852
rect 222 30806 226 30852
rect 246 30806 250 30852
rect 270 30806 274 30852
rect 294 30806 298 30852
rect 318 30806 322 30852
rect 342 30806 346 30852
rect 366 30806 370 30852
rect 390 30806 394 30852
rect 414 30806 418 30852
rect 438 30806 442 30852
rect 462 30806 466 30852
rect 486 30806 490 30852
rect 510 30806 514 30852
rect 534 30806 538 30852
rect 558 30806 562 30852
rect 582 30806 586 30852
rect 589 30851 603 30852
rect 606 30851 613 30899
rect 619 30893 624 30900
rect 630 30893 634 30900
rect 629 30879 634 30893
rect 606 30806 610 30851
rect 630 30806 634 30879
rect 654 30827 658 30996
rect -2393 30804 651 30806
rect -2371 30734 -2366 30804
rect -2348 30734 -2343 30804
rect -2325 30734 -2320 30804
rect -2317 30800 -2309 30804
rect -2062 30800 -2054 30804
rect -2154 30796 -2138 30798
rect -2057 30796 -2054 30800
rect -2292 30790 -2054 30796
rect -2052 30790 -2044 30800
rect -2092 30774 -2062 30776
rect -2094 30770 -2062 30774
rect -2309 30740 -2301 30746
rect -2317 30734 -2309 30740
rect -2000 30734 -1992 30804
rect -1846 30797 -1806 30804
rect -1663 30800 -1655 30804
rect -1846 30790 -1680 30796
rect -1854 30774 -1806 30776
rect -1854 30770 -1680 30774
rect -1655 30740 -1647 30746
rect -1663 30734 -1655 30740
rect -1642 30734 -1637 30804
rect -1619 30734 -1614 30804
rect -1530 30734 -1526 30804
rect -1506 30734 -1502 30804
rect -1482 30734 -1478 30804
rect -1458 30734 -1454 30804
rect -1434 30734 -1430 30804
rect -1410 30734 -1406 30804
rect -1386 30734 -1382 30804
rect -1362 30734 -1358 30804
rect -1338 30734 -1334 30804
rect -1314 30734 -1310 30804
rect -1290 30734 -1286 30804
rect -1266 30734 -1262 30804
rect -1242 30734 -1238 30804
rect -1218 30734 -1214 30804
rect -1194 30734 -1190 30804
rect -1170 30734 -1166 30804
rect -1146 30734 -1142 30804
rect -1122 30734 -1118 30804
rect -1098 30734 -1094 30804
rect -1074 30734 -1070 30804
rect -1050 30734 -1046 30804
rect -1026 30734 -1022 30804
rect -1002 30734 -998 30804
rect -978 30734 -974 30804
rect -954 30734 -950 30804
rect -930 30734 -926 30804
rect -906 30734 -902 30804
rect -882 30734 -878 30804
rect -858 30759 -854 30804
rect -869 30758 -835 30759
rect -834 30758 -830 30804
rect -810 30758 -806 30804
rect -786 30758 -782 30804
rect -762 30758 -758 30804
rect -738 30758 -734 30804
rect -714 30758 -710 30804
rect -690 30758 -686 30804
rect -666 30758 -662 30804
rect -642 30758 -638 30804
rect -618 30758 -614 30804
rect -594 30758 -590 30804
rect -570 30758 -566 30804
rect -546 30758 -542 30804
rect -522 30758 -518 30804
rect -498 30758 -494 30804
rect -474 30758 -470 30804
rect -450 30758 -446 30804
rect -426 30758 -422 30804
rect -402 30758 -398 30804
rect -378 30758 -374 30804
rect -354 30758 -350 30804
rect -330 30758 -326 30804
rect -306 30758 -302 30804
rect -282 30758 -278 30804
rect -258 30758 -254 30804
rect -234 30758 -230 30804
rect -210 30758 -206 30804
rect -186 30758 -182 30804
rect -162 30758 -158 30804
rect -138 30758 -134 30804
rect -114 30758 -110 30804
rect -90 30758 -86 30804
rect -66 30758 -62 30804
rect -42 30758 -38 30804
rect -18 30758 -14 30804
rect 6 30758 10 30804
rect 30 30758 34 30804
rect 54 30758 58 30804
rect 78 30758 82 30804
rect 102 30758 106 30804
rect 126 30758 130 30804
rect 150 30758 154 30804
rect 174 30758 178 30804
rect 198 30758 202 30804
rect 222 30758 226 30804
rect 246 30758 250 30804
rect 270 30758 274 30804
rect 294 30758 298 30804
rect 318 30758 322 30804
rect 342 30758 346 30804
rect 366 30758 370 30804
rect 390 30758 394 30804
rect 414 30758 418 30804
rect 438 30758 442 30804
rect 462 30758 466 30804
rect 486 30758 490 30804
rect 510 30758 514 30804
rect 534 30758 538 30804
rect 558 30758 562 30804
rect 582 30758 586 30804
rect 606 30758 610 30804
rect 630 30758 634 30804
rect 637 30803 651 30804
rect 654 30803 661 30827
rect 654 30758 658 30803
rect 678 30758 682 30996
rect 702 30758 706 30996
rect 726 30758 730 30996
rect 750 30758 754 30996
rect 774 30758 778 30996
rect 798 30758 802 30996
rect 822 30758 826 30996
rect 846 30758 850 30996
rect 870 30758 874 30996
rect 894 30758 898 30996
rect 918 30758 922 30996
rect 942 30758 946 30996
rect 966 30758 970 30996
rect 990 30758 994 30996
rect 1014 30879 1018 30996
rect 1003 30878 1037 30879
rect 1038 30878 1042 30996
rect 1062 30878 1066 30996
rect 1086 30878 1090 30996
rect 1110 30878 1114 30996
rect 1134 30878 1138 30996
rect 1158 30878 1162 30996
rect 1182 30878 1186 30996
rect 1206 30995 1210 30996
rect 1206 30974 1213 30995
rect 1230 30974 1234 30996
rect 1254 30974 1258 30996
rect 1278 30974 1282 30996
rect 1302 30974 1306 30996
rect 1326 30974 1330 30996
rect 1350 30974 1354 30996
rect 1374 30974 1378 30996
rect 1398 30974 1402 30996
rect 1422 30974 1426 30996
rect 1446 30974 1450 30996
rect 1470 30974 1474 30996
rect 1494 30974 1498 30996
rect 1518 30974 1522 30996
rect 1542 30974 1546 30996
rect 1566 30974 1570 30996
rect 1590 30974 1594 30996
rect 1614 30974 1618 30996
rect 1638 30974 1642 30996
rect 1662 30974 1666 30996
rect 1686 30974 1690 30996
rect 1710 30974 1714 30996
rect 1734 30974 1738 30996
rect 1758 30974 1762 30996
rect 1782 30974 1786 30996
rect 1806 30974 1810 30996
rect 1830 30974 1834 30996
rect 1854 30974 1858 30996
rect 1878 30974 1882 30996
rect 1902 30974 1906 30996
rect 1926 30974 1930 30996
rect 1950 30974 1954 30996
rect 1963 30989 1968 30996
rect 1974 30989 1978 30996
rect 1981 30995 1995 30996
rect 1973 30975 1978 30989
rect 1987 30985 1995 30989
rect 1981 30975 1987 30985
rect 1963 30974 1995 30975
rect 1189 30972 1995 30974
rect 1189 30971 1203 30972
rect 1206 30947 1213 30972
rect 1206 30878 1210 30947
rect 1230 30878 1234 30972
rect 1254 30878 1258 30972
rect 1278 30878 1282 30972
rect 1302 30878 1306 30972
rect 1326 30878 1330 30972
rect 1350 30878 1354 30972
rect 1374 30878 1378 30972
rect 1398 30878 1402 30972
rect 1422 30878 1426 30972
rect 1446 30878 1450 30972
rect 1470 30878 1474 30972
rect 1494 30878 1498 30972
rect 1518 30878 1522 30972
rect 1542 30878 1546 30972
rect 1566 30878 1570 30972
rect 1590 30878 1594 30972
rect 1614 30878 1618 30972
rect 1638 30878 1642 30972
rect 1662 30878 1666 30972
rect 1686 30878 1690 30972
rect 1710 30878 1714 30972
rect 1734 30878 1738 30972
rect 1758 30878 1762 30972
rect 1782 30878 1786 30972
rect 1806 30878 1810 30972
rect 1830 30878 1834 30972
rect 1854 30878 1858 30972
rect 1878 30878 1882 30972
rect 1902 30878 1906 30972
rect 1926 30878 1930 30972
rect 1950 30878 1954 30972
rect 1963 30965 1968 30972
rect 1981 30971 1995 30972
rect 1973 30951 1978 30965
rect 1963 30917 1968 30927
rect 1974 30917 1978 30951
rect 1973 30903 1978 30917
rect 1987 30913 1995 30917
rect 1981 30903 1987 30913
rect 1963 30878 1995 30879
rect 1003 30876 1995 30878
rect 1003 30869 1008 30876
rect 1014 30869 1018 30876
rect 1013 30855 1018 30869
rect 1003 30845 1008 30855
rect 1013 30831 1018 30845
rect 1014 30758 1018 30831
rect 1027 30797 1032 30807
rect 1038 30803 1042 30876
rect 1038 30797 1045 30803
rect 1037 30783 1045 30797
rect -869 30756 1035 30758
rect -869 30749 -864 30756
rect -858 30749 -854 30756
rect -859 30735 -854 30749
rect -869 30734 -835 30735
rect -2393 30732 -835 30734
rect -2371 30638 -2366 30732
rect -2348 30638 -2343 30732
rect -2325 30670 -2320 30732
rect -2317 30730 -2309 30732
rect -2000 30731 -1966 30732
rect -2000 30730 -1982 30731
rect -1663 30730 -1655 30732
rect -2028 30722 -2018 30724
rect -2309 30712 -2301 30718
rect -2091 30712 -2061 30719
rect -2317 30702 -2309 30712
rect -2044 30710 -2028 30712
rect -2026 30710 -2014 30722
rect -2084 30704 -2061 30710
rect -2044 30708 -2014 30710
rect -2292 30694 -2054 30703
rect -2325 30662 -2317 30670
rect -2325 30642 -2320 30662
rect -2317 30654 -2309 30662
rect -2325 30638 -2317 30642
rect -2000 30638 -1992 30730
rect -1982 30729 -1966 30730
rect -1980 30712 -1932 30719
rect -1655 30712 -1647 30718
rect -1846 30694 -1680 30703
rect -1663 30702 -1655 30712
rect -1671 30662 -1663 30670
rect -1663 30654 -1655 30662
rect -1671 30638 -1663 30642
rect -1642 30638 -1637 30732
rect -1619 30638 -1614 30732
rect -1530 30638 -1526 30732
rect -1506 30638 -1502 30732
rect -1482 30638 -1478 30732
rect -1458 30638 -1454 30732
rect -1434 30638 -1430 30732
rect -1410 30638 -1406 30732
rect -1386 30638 -1382 30732
rect -1362 30638 -1358 30732
rect -1338 30638 -1334 30732
rect -1314 30638 -1310 30732
rect -1290 30638 -1286 30732
rect -1266 30638 -1262 30732
rect -1242 30638 -1238 30732
rect -1218 30638 -1214 30732
rect -1194 30638 -1190 30732
rect -1170 30638 -1166 30732
rect -1146 30638 -1142 30732
rect -1122 30638 -1118 30732
rect -1098 30638 -1094 30732
rect -1074 30638 -1070 30732
rect -1050 30638 -1046 30732
rect -1026 30638 -1022 30732
rect -1002 30638 -998 30732
rect -978 30638 -974 30732
rect -954 30638 -950 30732
rect -930 30638 -926 30732
rect -906 30638 -902 30732
rect -882 30638 -878 30732
rect -869 30725 -864 30732
rect -859 30711 -854 30725
rect -858 30638 -854 30711
rect -834 30683 -830 30756
rect -2393 30636 -837 30638
rect -2371 30590 -2366 30636
rect -2348 30590 -2343 30636
rect -2325 30628 -2317 30636
rect -2018 30635 -2004 30636
rect -2000 30635 -1992 30636
rect -2072 30634 -1928 30635
rect -2072 30628 -2053 30634
rect -2325 30612 -2320 30628
rect -2317 30626 -2309 30628
rect -2309 30614 -2301 30626
rect -2092 30619 -2062 30624
rect -2317 30612 -2309 30614
rect -2325 30600 -2317 30612
rect -2098 30606 -2096 30617
rect -2092 30606 -2084 30619
rect -2000 30618 -1992 30634
rect -1972 30628 -1928 30634
rect -1924 30628 -1918 30636
rect -1671 30628 -1663 30636
rect -1663 30626 -1655 30628
rect -2083 30608 -2062 30617
rect -2027 30616 -1992 30618
rect -2018 30608 -2002 30616
rect -2000 30608 -1992 30616
rect -2100 30601 -2096 30606
rect -2083 30601 -2053 30606
rect -2003 30604 -1990 30608
rect -1972 30606 -1964 30615
rect -1928 30614 -1924 30617
rect -1655 30614 -1647 30626
rect -1663 30612 -1655 30614
rect -2325 30590 -2320 30600
rect -2317 30598 -2309 30600
rect -2309 30590 -2301 30598
rect -2004 30594 -2003 30604
rect -2062 30590 -2012 30592
rect -2000 30590 -1992 30604
rect -1972 30601 -1924 30606
rect -1864 30601 -1796 30607
rect -1671 30600 -1663 30612
rect -1663 30598 -1655 30600
rect -1864 30590 -1796 30591
rect -1655 30590 -1647 30598
rect -1642 30590 -1637 30636
rect -1619 30590 -1614 30636
rect -1530 30590 -1526 30636
rect -1506 30590 -1502 30636
rect -1482 30590 -1478 30636
rect -1458 30590 -1454 30636
rect -1434 30590 -1430 30636
rect -1410 30590 -1406 30636
rect -1386 30590 -1382 30636
rect -1362 30590 -1358 30636
rect -1338 30590 -1334 30636
rect -1325 30605 -1320 30615
rect -1314 30605 -1310 30636
rect -1315 30591 -1310 30605
rect -1314 30590 -1310 30591
rect -1290 30590 -1286 30636
rect -1266 30590 -1262 30636
rect -1242 30590 -1238 30636
rect -1218 30590 -1214 30636
rect -1194 30590 -1190 30636
rect -1170 30590 -1166 30636
rect -1146 30590 -1142 30636
rect -1122 30590 -1118 30636
rect -1098 30590 -1094 30636
rect -1074 30590 -1070 30636
rect -1050 30590 -1046 30636
rect -1026 30590 -1022 30636
rect -1002 30590 -998 30636
rect -978 30590 -974 30636
rect -954 30590 -950 30636
rect -930 30590 -926 30636
rect -906 30590 -902 30636
rect -882 30590 -878 30636
rect -858 30590 -854 30636
rect -851 30635 -837 30636
rect -834 30635 -827 30683
rect -834 30590 -830 30635
rect -810 30590 -806 30756
rect -786 30590 -782 30756
rect -762 30590 -758 30756
rect -738 30590 -734 30756
rect -714 30590 -710 30756
rect -690 30590 -686 30756
rect -666 30590 -662 30756
rect -642 30590 -638 30756
rect -618 30590 -614 30756
rect -594 30590 -590 30756
rect -570 30590 -566 30756
rect -546 30590 -542 30756
rect -522 30590 -518 30756
rect -498 30590 -494 30756
rect -474 30590 -470 30756
rect -450 30590 -446 30756
rect -426 30755 -422 30756
rect -426 30731 -419 30755
rect -426 30590 -422 30731
rect -402 30590 -398 30756
rect -378 30590 -374 30756
rect -354 30590 -350 30756
rect -330 30590 -326 30756
rect -306 30590 -302 30756
rect -282 30590 -278 30756
rect -258 30590 -254 30756
rect -234 30590 -230 30756
rect -210 30590 -206 30756
rect -186 30590 -182 30756
rect -162 30590 -158 30756
rect -138 30590 -134 30756
rect -114 30590 -110 30756
rect -90 30590 -86 30756
rect -66 30590 -62 30756
rect -42 30590 -38 30756
rect -18 30590 -14 30756
rect 6 30590 10 30756
rect 30 30590 34 30756
rect 54 30590 58 30756
rect 78 30590 82 30756
rect 102 30590 106 30756
rect 126 30590 130 30756
rect 150 30590 154 30756
rect 174 30590 178 30756
rect 198 30590 202 30756
rect 222 30590 226 30756
rect 246 30590 250 30756
rect 270 30590 274 30756
rect 294 30590 298 30756
rect 318 30590 322 30756
rect 342 30590 346 30756
rect 366 30590 370 30756
rect 390 30590 394 30756
rect 414 30590 418 30756
rect 438 30590 442 30756
rect 462 30590 466 30756
rect 486 30590 490 30756
rect 510 30590 514 30756
rect 534 30590 538 30756
rect 558 30590 562 30756
rect 582 30590 586 30756
rect 606 30590 610 30756
rect 630 30590 634 30756
rect 654 30590 658 30756
rect 678 30590 682 30756
rect 702 30590 706 30756
rect 726 30590 730 30756
rect 750 30590 754 30756
rect 774 30590 778 30756
rect 798 30590 802 30756
rect 822 30590 826 30756
rect 846 30590 850 30756
rect 859 30677 864 30687
rect 870 30677 874 30756
rect 869 30663 874 30677
rect 870 30590 874 30663
rect 894 30611 898 30756
rect -2393 30588 891 30590
rect -2371 30542 -2366 30588
rect -2348 30542 -2343 30588
rect -2325 30584 -2320 30588
rect -2309 30586 -2301 30588
rect -2317 30584 -2309 30586
rect -2325 30572 -2317 30584
rect -2325 30542 -2320 30572
rect -2317 30570 -2309 30572
rect -2092 30558 -2062 30560
rect -2094 30554 -2062 30558
rect -2000 30542 -1992 30588
rect -1655 30586 -1647 30588
rect -1663 30584 -1655 30586
rect -1671 30572 -1663 30584
rect -1663 30570 -1655 30572
rect -1854 30558 -1806 30560
rect -1854 30554 -1680 30558
rect -1642 30542 -1637 30588
rect -1619 30542 -1614 30588
rect -1530 30542 -1526 30588
rect -1506 30542 -1502 30588
rect -1482 30542 -1478 30588
rect -1458 30542 -1454 30588
rect -1434 30542 -1430 30588
rect -1410 30542 -1406 30588
rect -1386 30542 -1382 30588
rect -1362 30542 -1358 30588
rect -1338 30542 -1334 30588
rect -1314 30542 -1310 30588
rect -1290 30542 -1286 30588
rect -1266 30542 -1262 30588
rect -1242 30542 -1238 30588
rect -1218 30542 -1214 30588
rect -1194 30542 -1190 30588
rect -1170 30542 -1166 30588
rect -1146 30542 -1142 30588
rect -1122 30542 -1118 30588
rect -1098 30542 -1094 30588
rect -1074 30542 -1070 30588
rect -1050 30542 -1046 30588
rect -1026 30542 -1022 30588
rect -1002 30542 -998 30588
rect -978 30542 -974 30588
rect -954 30542 -950 30588
rect -930 30542 -926 30588
rect -906 30542 -902 30588
rect -882 30542 -878 30588
rect -858 30542 -854 30588
rect -834 30542 -830 30588
rect -810 30542 -806 30588
rect -786 30542 -782 30588
rect -762 30542 -758 30588
rect -738 30542 -734 30588
rect -714 30542 -710 30588
rect -690 30542 -686 30588
rect -666 30542 -662 30588
rect -642 30542 -638 30588
rect -618 30542 -614 30588
rect -594 30542 -590 30588
rect -570 30542 -566 30588
rect -546 30542 -542 30588
rect -522 30542 -518 30588
rect -498 30542 -494 30588
rect -474 30542 -470 30588
rect -450 30542 -446 30588
rect -426 30542 -422 30588
rect -402 30542 -398 30588
rect -378 30542 -374 30588
rect -354 30542 -350 30588
rect -330 30542 -326 30588
rect -317 30557 -312 30567
rect -306 30557 -302 30588
rect -307 30543 -302 30557
rect -317 30542 -283 30543
rect -2393 30540 -283 30542
rect -2371 30518 -2366 30540
rect -2348 30518 -2343 30540
rect -2325 30518 -2320 30540
rect -2072 30538 -2036 30539
rect -2072 30532 -2054 30538
rect -2309 30524 -2301 30532
rect -2317 30518 -2309 30524
rect -2092 30523 -2062 30528
rect -2000 30519 -1992 30540
rect -1938 30539 -1906 30540
rect -1920 30538 -1906 30539
rect -1806 30532 -1680 30538
rect -1854 30523 -1806 30528
rect -1655 30524 -1647 30532
rect -1982 30519 -1966 30520
rect -2000 30518 -1966 30519
rect -1846 30518 -1806 30521
rect -1663 30518 -1655 30524
rect -1642 30518 -1637 30540
rect -1619 30518 -1614 30540
rect -1530 30518 -1526 30540
rect -1506 30518 -1502 30540
rect -1482 30518 -1478 30540
rect -1458 30518 -1454 30540
rect -1434 30518 -1430 30540
rect -1410 30518 -1406 30540
rect -1386 30518 -1382 30540
rect -1362 30518 -1358 30540
rect -1338 30518 -1334 30540
rect -1314 30518 -1310 30540
rect -1290 30539 -1286 30540
rect -2393 30516 -1293 30518
rect -2371 30494 -2366 30516
rect -2348 30494 -2343 30516
rect -2325 30494 -2320 30516
rect -2000 30514 -1966 30516
rect -2309 30496 -2301 30504
rect -2062 30503 -2054 30510
rect -2092 30496 -2084 30503
rect -2062 30496 -2026 30498
rect -2317 30494 -2309 30496
rect -2062 30494 -2012 30496
rect -2000 30494 -1992 30514
rect -1982 30513 -1966 30514
rect -1846 30512 -1806 30516
rect -1846 30505 -1798 30510
rect -1806 30503 -1798 30505
rect -1854 30501 -1846 30503
rect -1854 30496 -1806 30501
rect -1655 30496 -1647 30504
rect -1864 30494 -1796 30495
rect -1663 30494 -1655 30496
rect -1642 30494 -1637 30516
rect -1619 30494 -1614 30516
rect -1530 30494 -1526 30516
rect -1506 30494 -1502 30516
rect -1482 30494 -1478 30516
rect -1458 30494 -1454 30516
rect -1434 30494 -1430 30516
rect -1410 30494 -1406 30516
rect -1386 30494 -1382 30516
rect -1362 30494 -1358 30516
rect -1338 30494 -1334 30516
rect -1314 30494 -1310 30516
rect -1307 30515 -1293 30516
rect -1290 30515 -1283 30539
rect -1290 30494 -1286 30515
rect -1266 30494 -1262 30540
rect -1242 30494 -1238 30540
rect -1218 30494 -1214 30540
rect -1194 30494 -1190 30540
rect -1170 30494 -1166 30540
rect -1146 30494 -1142 30540
rect -1122 30494 -1118 30540
rect -1098 30494 -1094 30540
rect -1074 30494 -1070 30540
rect -1050 30494 -1046 30540
rect -1026 30494 -1022 30540
rect -1002 30494 -998 30540
rect -978 30494 -974 30540
rect -954 30494 -950 30540
rect -930 30494 -926 30540
rect -906 30494 -902 30540
rect -882 30494 -878 30540
rect -858 30494 -854 30540
rect -834 30494 -830 30540
rect -810 30494 -806 30540
rect -786 30494 -782 30540
rect -762 30494 -758 30540
rect -738 30494 -734 30540
rect -714 30494 -710 30540
rect -690 30494 -686 30540
rect -666 30494 -662 30540
rect -642 30494 -638 30540
rect -618 30494 -614 30540
rect -594 30494 -590 30540
rect -570 30494 -566 30540
rect -546 30494 -542 30540
rect -533 30509 -528 30519
rect -522 30509 -518 30540
rect -523 30495 -518 30509
rect -522 30494 -518 30495
rect -498 30494 -494 30540
rect -474 30494 -470 30540
rect -450 30494 -446 30540
rect -426 30494 -422 30540
rect -402 30494 -398 30540
rect -378 30494 -374 30540
rect -354 30494 -350 30540
rect -330 30494 -326 30540
rect -317 30533 -312 30540
rect -307 30519 -302 30533
rect -306 30494 -302 30519
rect -282 30494 -278 30588
rect -258 30494 -254 30588
rect -234 30494 -230 30588
rect -210 30494 -206 30588
rect -186 30494 -182 30588
rect -162 30494 -158 30588
rect -138 30494 -134 30588
rect -114 30494 -110 30588
rect -90 30494 -86 30588
rect -66 30494 -62 30588
rect -42 30494 -38 30588
rect -18 30494 -14 30588
rect 6 30494 10 30588
rect 30 30494 34 30588
rect 54 30494 58 30588
rect 78 30494 82 30588
rect 102 30494 106 30588
rect 126 30494 130 30588
rect 150 30494 154 30588
rect 174 30494 178 30588
rect 198 30494 202 30588
rect 222 30494 226 30588
rect 246 30494 250 30588
rect 270 30494 274 30588
rect 294 30494 298 30588
rect 318 30494 322 30588
rect 342 30494 346 30588
rect 366 30494 370 30588
rect 390 30494 394 30588
rect 414 30494 418 30588
rect 438 30494 442 30588
rect 462 30494 466 30588
rect 486 30494 490 30588
rect 510 30494 514 30588
rect 534 30494 538 30588
rect 558 30494 562 30588
rect 582 30494 586 30588
rect 606 30494 610 30588
rect 630 30494 634 30588
rect 654 30494 658 30588
rect 678 30494 682 30588
rect 702 30494 706 30588
rect 726 30494 730 30588
rect 750 30494 754 30588
rect 774 30494 778 30588
rect 798 30494 802 30588
rect 822 30494 826 30588
rect 846 30494 850 30588
rect 870 30494 874 30588
rect 877 30587 891 30588
rect 894 30587 901 30611
rect 894 30494 898 30587
rect 918 30494 922 30756
rect 942 30494 946 30756
rect 966 30494 970 30756
rect 990 30494 994 30756
rect 1014 30494 1018 30756
rect 1021 30755 1035 30756
rect 1038 30755 1045 30783
rect 1038 30663 1042 30755
rect 1062 30731 1066 30876
rect 1062 30707 1069 30731
rect 1027 30662 1061 30663
rect 1062 30662 1066 30707
rect 1086 30662 1090 30876
rect 1110 30662 1114 30876
rect 1134 30662 1138 30876
rect 1158 30662 1162 30876
rect 1182 30662 1186 30876
rect 1206 30662 1210 30876
rect 1230 30662 1234 30876
rect 1254 30662 1258 30876
rect 1278 30662 1282 30876
rect 1302 30662 1306 30876
rect 1326 30662 1330 30876
rect 1350 30662 1354 30876
rect 1374 30662 1378 30876
rect 1398 30662 1402 30876
rect 1422 30662 1426 30876
rect 1446 30662 1450 30876
rect 1470 30662 1474 30876
rect 1494 30662 1498 30876
rect 1518 30662 1522 30876
rect 1542 30662 1546 30876
rect 1566 30662 1570 30876
rect 1590 30662 1594 30876
rect 1614 30662 1618 30876
rect 1638 30662 1642 30876
rect 1662 30662 1666 30876
rect 1686 30662 1690 30876
rect 1710 30662 1714 30876
rect 1734 30662 1738 30876
rect 1758 30662 1762 30876
rect 1782 30662 1786 30876
rect 1806 30662 1810 30876
rect 1830 30662 1834 30876
rect 1854 30662 1858 30876
rect 1878 30662 1882 30876
rect 1902 30662 1906 30876
rect 1926 30662 1930 30876
rect 1950 30662 1954 30876
rect 1963 30869 1968 30876
rect 1981 30875 1995 30876
rect 1973 30855 1978 30869
rect 1974 30662 1978 30855
rect 1987 30749 1992 30759
rect 1997 30735 2002 30749
rect 1998 30662 2002 30735
rect 2011 30662 2019 30663
rect 1027 30660 2019 30662
rect 1027 30653 1032 30660
rect 1038 30653 1042 30660
rect 1037 30639 1042 30653
rect 1027 30629 1032 30639
rect 1037 30615 1042 30629
rect 1038 30494 1042 30615
rect 1062 30587 1066 30660
rect 1062 30566 1069 30587
rect 1086 30566 1090 30660
rect 1110 30566 1114 30660
rect 1134 30566 1138 30660
rect 1158 30566 1162 30660
rect 1182 30566 1186 30660
rect 1206 30566 1210 30660
rect 1230 30566 1234 30660
rect 1254 30566 1258 30660
rect 1278 30566 1282 30660
rect 1302 30566 1306 30660
rect 1326 30566 1330 30660
rect 1350 30566 1354 30660
rect 1374 30566 1378 30660
rect 1398 30566 1402 30660
rect 1422 30566 1426 30660
rect 1446 30566 1450 30660
rect 1470 30566 1474 30660
rect 1494 30566 1498 30660
rect 1518 30566 1522 30660
rect 1542 30566 1546 30660
rect 1566 30566 1570 30660
rect 1590 30566 1594 30660
rect 1614 30566 1618 30660
rect 1638 30566 1642 30660
rect 1662 30566 1666 30660
rect 1686 30566 1690 30660
rect 1710 30566 1714 30660
rect 1734 30566 1738 30660
rect 1758 30566 1762 30660
rect 1782 30566 1786 30660
rect 1806 30566 1810 30660
rect 1830 30566 1834 30660
rect 1854 30566 1858 30660
rect 1878 30566 1882 30660
rect 1902 30566 1906 30660
rect 1926 30566 1930 30660
rect 1950 30566 1954 30660
rect 1974 30566 1978 30660
rect 1998 30566 2002 30660
rect 2005 30659 2019 30660
rect 2011 30653 2016 30659
rect 2021 30639 2026 30653
rect 2011 30581 2016 30591
rect 2022 30581 2026 30639
rect 2021 30567 2026 30581
rect 2035 30577 2043 30581
rect 2029 30567 2035 30577
rect 2011 30566 2043 30567
rect 1045 30564 2043 30566
rect 1045 30563 1059 30564
rect 1062 30539 1069 30564
rect 1062 30494 1066 30539
rect 1086 30494 1090 30564
rect 1110 30494 1114 30564
rect 1134 30494 1138 30564
rect 1158 30494 1162 30564
rect 1182 30494 1186 30564
rect 1206 30494 1210 30564
rect 1230 30494 1234 30564
rect 1254 30494 1258 30564
rect 1278 30494 1282 30564
rect 1302 30494 1306 30564
rect 1326 30494 1330 30564
rect 1350 30494 1354 30564
rect 1374 30494 1378 30564
rect 1398 30494 1402 30564
rect 1422 30494 1426 30564
rect 1446 30494 1450 30564
rect 1470 30494 1474 30564
rect 1494 30494 1498 30564
rect 1518 30494 1522 30564
rect 1542 30494 1546 30564
rect 1566 30494 1570 30564
rect 1590 30494 1594 30564
rect 1614 30494 1618 30564
rect 1638 30494 1642 30564
rect 1662 30494 1666 30564
rect 1686 30494 1690 30564
rect 1710 30494 1714 30564
rect 1734 30494 1738 30564
rect 1758 30494 1762 30564
rect 1782 30494 1786 30564
rect 1806 30494 1810 30564
rect 1830 30494 1834 30564
rect 1854 30494 1858 30564
rect 1878 30494 1882 30564
rect 1902 30494 1906 30564
rect 1926 30494 1930 30564
rect 1950 30494 1954 30564
rect 1974 30494 1978 30564
rect 1998 30494 2002 30564
rect 2011 30557 2016 30564
rect 2029 30563 2043 30564
rect 2021 30543 2026 30557
rect 2022 30495 2026 30543
rect 2011 30494 2043 30495
rect -2393 30492 2043 30494
rect -2371 30422 -2366 30492
rect -2348 30422 -2343 30492
rect -2325 30422 -2320 30492
rect -2317 30488 -2309 30492
rect -2062 30488 -2054 30492
rect -2154 30484 -2138 30486
rect -2057 30484 -2054 30488
rect -2292 30478 -2054 30484
rect -2052 30478 -2044 30488
rect -2092 30462 -2062 30464
rect -2094 30458 -2062 30462
rect -2309 30428 -2301 30434
rect -2317 30422 -2309 30428
rect -2000 30422 -1992 30492
rect -1846 30485 -1806 30492
rect -1663 30488 -1655 30492
rect -1846 30478 -1680 30484
rect -1854 30462 -1806 30464
rect -1854 30458 -1680 30462
rect -1655 30428 -1647 30434
rect -1663 30422 -1655 30428
rect -1642 30422 -1637 30492
rect -1619 30422 -1614 30492
rect -1530 30422 -1526 30492
rect -1506 30422 -1502 30492
rect -1482 30422 -1478 30492
rect -1458 30422 -1454 30492
rect -1434 30422 -1430 30492
rect -1410 30422 -1406 30492
rect -1386 30422 -1382 30492
rect -1362 30422 -1358 30492
rect -1338 30422 -1334 30492
rect -1314 30422 -1310 30492
rect -1290 30422 -1286 30492
rect -1266 30422 -1262 30492
rect -1242 30422 -1238 30492
rect -1218 30422 -1214 30492
rect -1194 30422 -1190 30492
rect -1170 30422 -1166 30492
rect -1146 30422 -1142 30492
rect -1122 30422 -1118 30492
rect -1098 30422 -1094 30492
rect -1074 30422 -1070 30492
rect -1050 30422 -1046 30492
rect -1026 30422 -1022 30492
rect -1002 30422 -998 30492
rect -978 30422 -974 30492
rect -954 30422 -950 30492
rect -930 30422 -926 30492
rect -906 30422 -902 30492
rect -882 30422 -878 30492
rect -858 30422 -854 30492
rect -834 30422 -830 30492
rect -810 30422 -806 30492
rect -786 30422 -782 30492
rect -762 30422 -758 30492
rect -738 30422 -734 30492
rect -714 30422 -710 30492
rect -690 30422 -686 30492
rect -666 30422 -662 30492
rect -642 30422 -638 30492
rect -618 30422 -614 30492
rect -594 30422 -590 30492
rect -570 30422 -566 30492
rect -546 30422 -542 30492
rect -522 30422 -518 30492
rect -498 30443 -494 30492
rect -2393 30420 -501 30422
rect -2371 30326 -2366 30420
rect -2348 30326 -2343 30420
rect -2325 30358 -2320 30420
rect -2317 30418 -2309 30420
rect -2000 30419 -1966 30420
rect -2000 30418 -1982 30419
rect -1663 30418 -1655 30420
rect -2028 30410 -2018 30412
rect -2309 30400 -2301 30406
rect -2091 30400 -2061 30407
rect -2317 30390 -2309 30400
rect -2044 30398 -2028 30400
rect -2026 30398 -2014 30410
rect -2084 30392 -2061 30398
rect -2044 30396 -2014 30398
rect -2292 30382 -2054 30391
rect -2325 30350 -2317 30358
rect -2325 30330 -2320 30350
rect -2317 30342 -2309 30350
rect -2325 30326 -2317 30330
rect -2000 30326 -1992 30418
rect -1982 30417 -1966 30418
rect -1980 30400 -1932 30407
rect -1655 30400 -1647 30406
rect -1846 30382 -1680 30391
rect -1663 30390 -1655 30400
rect -1671 30350 -1663 30358
rect -1663 30342 -1655 30350
rect -1671 30326 -1663 30330
rect -1642 30326 -1637 30420
rect -1619 30326 -1614 30420
rect -1530 30326 -1526 30420
rect -1506 30326 -1502 30420
rect -1482 30326 -1478 30420
rect -1458 30326 -1454 30420
rect -1434 30326 -1430 30420
rect -1410 30326 -1406 30420
rect -1386 30326 -1382 30420
rect -1362 30326 -1358 30420
rect -1338 30326 -1334 30420
rect -1314 30326 -1310 30420
rect -1290 30326 -1286 30420
rect -1266 30326 -1262 30420
rect -1242 30326 -1238 30420
rect -1218 30326 -1214 30420
rect -1194 30326 -1190 30420
rect -1170 30326 -1166 30420
rect -1146 30326 -1142 30420
rect -1122 30326 -1118 30420
rect -1098 30326 -1094 30420
rect -1074 30326 -1070 30420
rect -1050 30326 -1046 30420
rect -1026 30326 -1022 30420
rect -1002 30326 -998 30420
rect -978 30326 -974 30420
rect -954 30326 -950 30420
rect -930 30326 -926 30420
rect -906 30326 -902 30420
rect -882 30326 -878 30420
rect -858 30326 -854 30420
rect -834 30326 -830 30420
rect -821 30365 -816 30375
rect -810 30365 -806 30420
rect -811 30351 -806 30365
rect -810 30326 -806 30351
rect -786 30326 -782 30420
rect -762 30326 -758 30420
rect -738 30326 -734 30420
rect -714 30326 -710 30420
rect -690 30326 -686 30420
rect -666 30326 -662 30420
rect -642 30326 -638 30420
rect -618 30326 -614 30420
rect -594 30326 -590 30420
rect -570 30326 -566 30420
rect -546 30326 -542 30420
rect -522 30326 -518 30420
rect -515 30419 -501 30420
rect -498 30419 -491 30443
rect -498 30326 -494 30419
rect -474 30326 -470 30492
rect -450 30326 -446 30492
rect -426 30326 -422 30492
rect -402 30326 -398 30492
rect -378 30326 -374 30492
rect -354 30326 -350 30492
rect -330 30326 -326 30492
rect -306 30326 -302 30492
rect -282 30491 -278 30492
rect -282 30443 -275 30491
rect -282 30326 -278 30443
rect -258 30326 -254 30492
rect -234 30326 -230 30492
rect -210 30326 -206 30492
rect -186 30326 -182 30492
rect -162 30326 -158 30492
rect -138 30326 -134 30492
rect -114 30326 -110 30492
rect -90 30326 -86 30492
rect -66 30326 -62 30492
rect -42 30326 -38 30492
rect -18 30326 -14 30492
rect 6 30326 10 30492
rect 30 30326 34 30492
rect 54 30326 58 30492
rect 78 30326 82 30492
rect 102 30326 106 30492
rect 126 30326 130 30492
rect 150 30326 154 30492
rect 174 30326 178 30492
rect 198 30326 202 30492
rect 211 30341 216 30351
rect 222 30341 226 30492
rect 221 30327 226 30341
rect 211 30326 245 30327
rect -2393 30324 245 30326
rect -2371 30278 -2366 30324
rect -2348 30278 -2343 30324
rect -2325 30316 -2317 30324
rect -2018 30323 -2004 30324
rect -2000 30323 -1992 30324
rect -2072 30322 -1928 30323
rect -2072 30316 -2053 30322
rect -2325 30300 -2320 30316
rect -2317 30314 -2309 30316
rect -2309 30302 -2301 30314
rect -2092 30307 -2062 30312
rect -2317 30300 -2309 30302
rect -2325 30288 -2317 30300
rect -2098 30294 -2096 30305
rect -2092 30294 -2084 30307
rect -2000 30306 -1992 30322
rect -1972 30316 -1928 30322
rect -1924 30316 -1918 30324
rect -1671 30316 -1663 30324
rect -1663 30314 -1655 30316
rect -2083 30296 -2062 30305
rect -2027 30304 -1992 30306
rect -2018 30296 -2002 30304
rect -2000 30296 -1992 30304
rect -2100 30289 -2096 30294
rect -2083 30289 -2053 30294
rect -2003 30292 -1990 30296
rect -1972 30294 -1964 30303
rect -1928 30302 -1924 30305
rect -1655 30302 -1647 30314
rect -1663 30300 -1655 30302
rect -2325 30278 -2320 30288
rect -2317 30286 -2309 30288
rect -2309 30278 -2301 30286
rect -2004 30282 -2003 30292
rect -2062 30278 -2012 30280
rect -2000 30278 -1992 30292
rect -1972 30289 -1924 30294
rect -1864 30289 -1796 30295
rect -1671 30288 -1663 30300
rect -1663 30286 -1655 30288
rect -1864 30278 -1796 30279
rect -1655 30278 -1647 30286
rect -1642 30278 -1637 30324
rect -1619 30278 -1614 30324
rect -1530 30278 -1526 30324
rect -1506 30278 -1502 30324
rect -1482 30278 -1478 30324
rect -1458 30278 -1454 30324
rect -1434 30278 -1430 30324
rect -1410 30278 -1406 30324
rect -1386 30278 -1382 30324
rect -1362 30278 -1358 30324
rect -1338 30278 -1334 30324
rect -1314 30278 -1310 30324
rect -1290 30278 -1286 30324
rect -1266 30278 -1262 30324
rect -1242 30278 -1238 30324
rect -1218 30278 -1214 30324
rect -1194 30278 -1190 30324
rect -1170 30278 -1166 30324
rect -1146 30278 -1142 30324
rect -1122 30278 -1118 30324
rect -1098 30278 -1094 30324
rect -1074 30278 -1070 30324
rect -1050 30278 -1046 30324
rect -1026 30278 -1022 30324
rect -1002 30278 -998 30324
rect -978 30278 -974 30324
rect -954 30278 -950 30324
rect -930 30278 -926 30324
rect -906 30278 -902 30324
rect -882 30278 -878 30324
rect -858 30278 -854 30324
rect -834 30278 -830 30324
rect -810 30278 -806 30324
rect -786 30299 -782 30324
rect -2393 30276 -789 30278
rect -2371 30230 -2366 30276
rect -2348 30230 -2343 30276
rect -2325 30272 -2320 30276
rect -2309 30274 -2301 30276
rect -2317 30272 -2309 30274
rect -2325 30260 -2317 30272
rect -2325 30230 -2320 30260
rect -2317 30258 -2309 30260
rect -2092 30246 -2062 30248
rect -2094 30242 -2062 30246
rect -2000 30230 -1992 30276
rect -1655 30274 -1647 30276
rect -1663 30272 -1655 30274
rect -1671 30260 -1663 30272
rect -1663 30258 -1655 30260
rect -1854 30246 -1806 30248
rect -1854 30242 -1680 30246
rect -1642 30230 -1637 30276
rect -1619 30230 -1614 30276
rect -1530 30230 -1526 30276
rect -1506 30230 -1502 30276
rect -1482 30230 -1478 30276
rect -1458 30230 -1454 30276
rect -1434 30230 -1430 30276
rect -1410 30230 -1406 30276
rect -1386 30230 -1382 30276
rect -1362 30230 -1358 30276
rect -1338 30230 -1334 30276
rect -1314 30230 -1310 30276
rect -1290 30230 -1286 30276
rect -1266 30230 -1262 30276
rect -1242 30230 -1238 30276
rect -1218 30230 -1214 30276
rect -1194 30230 -1190 30276
rect -1170 30230 -1166 30276
rect -1146 30230 -1142 30276
rect -1122 30230 -1118 30276
rect -1098 30230 -1094 30276
rect -1074 30230 -1070 30276
rect -1050 30230 -1046 30276
rect -1026 30230 -1022 30276
rect -1002 30230 -998 30276
rect -978 30230 -974 30276
rect -954 30230 -950 30276
rect -930 30230 -926 30276
rect -906 30230 -902 30276
rect -882 30230 -878 30276
rect -858 30230 -854 30276
rect -834 30230 -830 30276
rect -810 30230 -806 30276
rect -803 30275 -789 30276
rect -786 30275 -779 30299
rect -786 30230 -782 30275
rect -773 30245 -768 30255
rect -762 30245 -758 30324
rect -763 30231 -758 30245
rect -773 30230 -739 30231
rect -2393 30228 -739 30230
rect -2371 30182 -2366 30228
rect -2348 30182 -2343 30228
rect -2325 30182 -2320 30228
rect -2309 30212 -2301 30222
rect -2317 30206 -2309 30212
rect -2097 30206 -2095 30215
rect -2309 30184 -2301 30194
rect -2097 30192 -2095 30196
rect -2292 30191 -2095 30192
rect -2097 30189 -2095 30191
rect -2084 30184 -2083 30227
rect -2069 30220 -2054 30222
rect -2054 30204 -2018 30206
rect -2054 30202 -2004 30204
rect -2059 30198 -2045 30202
rect -2054 30196 -2049 30198
rect -2317 30182 -2309 30184
rect -2084 30182 -2054 30184
rect -2044 30182 -2039 30196
rect -2025 30186 -2014 30192
rect -2000 30186 -1992 30228
rect -1920 30226 -1906 30228
rect -1977 30211 -1929 30217
rect -1655 30212 -1647 30222
rect -1977 30201 -1966 30211
rect -1663 30206 -1655 30212
rect -1977 30189 -1929 30191
rect -2033 30182 -1992 30186
rect -1655 30184 -1647 30194
rect -1663 30182 -1655 30184
rect -1642 30182 -1637 30228
rect -1619 30182 -1614 30228
rect -1530 30182 -1526 30228
rect -1506 30182 -1502 30228
rect -1482 30182 -1478 30228
rect -1458 30182 -1454 30228
rect -1434 30182 -1430 30228
rect -1410 30182 -1406 30228
rect -1386 30182 -1382 30228
rect -1362 30182 -1358 30228
rect -1338 30182 -1334 30228
rect -1314 30182 -1310 30228
rect -1290 30182 -1286 30228
rect -1266 30182 -1262 30228
rect -1242 30182 -1238 30228
rect -1218 30182 -1214 30228
rect -1194 30182 -1190 30228
rect -1170 30182 -1166 30228
rect -1146 30182 -1142 30228
rect -1122 30182 -1118 30228
rect -1098 30182 -1094 30228
rect -1074 30182 -1070 30228
rect -1050 30182 -1046 30228
rect -1026 30182 -1022 30228
rect -1002 30182 -998 30228
rect -978 30182 -974 30228
rect -954 30182 -950 30228
rect -930 30182 -926 30228
rect -906 30182 -902 30228
rect -882 30182 -878 30228
rect -858 30182 -854 30228
rect -834 30182 -830 30228
rect -810 30182 -806 30228
rect -786 30182 -782 30228
rect -773 30221 -768 30228
rect -763 30207 -758 30221
rect -762 30182 -758 30207
rect -738 30182 -734 30324
rect -714 30182 -710 30324
rect -690 30182 -686 30324
rect -666 30182 -662 30324
rect -642 30182 -638 30324
rect -618 30182 -614 30324
rect -594 30182 -590 30324
rect -570 30182 -566 30324
rect -546 30183 -542 30324
rect -557 30182 -523 30183
rect -2393 30180 -523 30182
rect -2371 30086 -2366 30180
rect -2348 30086 -2343 30180
rect -2325 30146 -2320 30180
rect -2317 30178 -2309 30180
rect -2084 30167 -2083 30180
rect -2084 30166 -2054 30167
rect -2325 30138 -2317 30146
rect -2325 30086 -2320 30138
rect -2317 30130 -2309 30138
rect -2117 30129 -2095 30139
rect -2045 30136 -2037 30150
rect -2309 30090 -2301 30100
rect -2087 30096 -2076 30104
rect -2017 30100 -2015 30107
rect -2317 30086 -2309 30090
rect -2092 30088 -2087 30096
rect -2092 30086 -2077 30087
rect -2000 30086 -1992 30180
rect -1663 30178 -1655 30180
rect -1969 30129 -1929 30141
rect -1671 30138 -1663 30146
rect -1663 30130 -1655 30138
rect -1655 30090 -1647 30100
rect -1928 30086 -1924 30087
rect -1854 30086 -1680 30087
rect -1663 30086 -1655 30090
rect -1642 30086 -1637 30180
rect -1619 30086 -1614 30180
rect -1530 30086 -1526 30180
rect -1506 30086 -1502 30180
rect -1482 30086 -1478 30180
rect -1458 30086 -1454 30180
rect -1434 30086 -1430 30180
rect -1410 30086 -1406 30180
rect -1386 30086 -1382 30180
rect -1362 30086 -1358 30180
rect -1338 30086 -1334 30180
rect -1314 30086 -1310 30180
rect -1290 30086 -1286 30180
rect -1266 30086 -1262 30180
rect -1242 30086 -1238 30180
rect -1218 30086 -1214 30180
rect -1194 30086 -1190 30180
rect -1170 30086 -1166 30180
rect -1146 30086 -1142 30180
rect -1122 30086 -1118 30180
rect -1098 30086 -1094 30180
rect -1074 30086 -1070 30180
rect -1050 30086 -1046 30180
rect -1026 30086 -1022 30180
rect -1002 30086 -998 30180
rect -978 30086 -974 30180
rect -954 30087 -950 30180
rect -965 30086 -931 30087
rect -2393 30084 -931 30086
rect -2371 30062 -2366 30084
rect -2348 30062 -2343 30084
rect -2325 30062 -2320 30084
rect -2092 30079 -2037 30084
rect -2021 30079 -1969 30084
rect -1921 30079 -1913 30084
rect -1854 30080 -1680 30084
rect -2100 30077 -2092 30078
rect -2309 30062 -2301 30072
rect -2100 30071 -2087 30077
rect -2051 30064 -2026 30066
rect -2062 30062 -2012 30064
rect -2000 30062 -1992 30079
rect -1969 30071 -1921 30078
rect -1969 30062 -1964 30071
rect -1864 30062 -1796 30063
rect -1655 30062 -1647 30072
rect -1642 30062 -1637 30084
rect -1619 30062 -1614 30084
rect -1530 30062 -1526 30084
rect -1506 30062 -1502 30084
rect -1482 30062 -1478 30084
rect -1458 30062 -1454 30084
rect -1434 30062 -1430 30084
rect -1410 30062 -1406 30084
rect -1386 30062 -1382 30084
rect -1362 30062 -1358 30084
rect -1338 30062 -1334 30084
rect -1314 30062 -1310 30084
rect -1290 30062 -1286 30084
rect -1266 30062 -1262 30084
rect -1242 30062 -1238 30084
rect -1218 30062 -1214 30084
rect -1194 30062 -1190 30084
rect -1170 30062 -1166 30084
rect -1146 30062 -1142 30084
rect -1122 30062 -1118 30084
rect -1098 30062 -1094 30084
rect -1074 30062 -1070 30084
rect -1050 30062 -1046 30084
rect -1026 30062 -1022 30084
rect -1002 30062 -998 30084
rect -978 30062 -974 30084
rect -965 30077 -960 30084
rect -954 30077 -950 30084
rect -955 30063 -950 30077
rect -954 30062 -950 30063
rect -930 30062 -926 30180
rect -906 30062 -902 30180
rect -882 30062 -878 30180
rect -858 30062 -854 30180
rect -834 30062 -830 30180
rect -810 30062 -806 30180
rect -786 30062 -782 30180
rect -762 30062 -758 30180
rect -738 30179 -734 30180
rect -738 30158 -731 30179
rect -714 30158 -710 30180
rect -690 30158 -686 30180
rect -666 30158 -662 30180
rect -642 30158 -638 30180
rect -618 30158 -614 30180
rect -594 30158 -590 30180
rect -570 30158 -566 30180
rect -557 30173 -552 30180
rect -546 30173 -542 30180
rect -547 30159 -542 30173
rect -546 30158 -542 30159
rect -522 30158 -518 30324
rect -498 30158 -494 30324
rect -474 30158 -470 30324
rect -450 30158 -446 30324
rect -426 30158 -422 30324
rect -402 30158 -398 30324
rect -378 30158 -374 30324
rect -354 30158 -350 30324
rect -330 30158 -326 30324
rect -306 30158 -302 30324
rect -282 30158 -278 30324
rect -258 30158 -254 30324
rect -234 30158 -230 30324
rect -210 30158 -206 30324
rect -186 30158 -182 30324
rect -162 30158 -158 30324
rect -138 30158 -134 30324
rect -114 30158 -110 30324
rect -90 30158 -86 30324
rect -66 30158 -62 30324
rect -42 30158 -38 30324
rect -18 30158 -14 30324
rect 6 30158 10 30324
rect 30 30158 34 30324
rect 54 30158 58 30324
rect 78 30158 82 30324
rect 102 30158 106 30324
rect 126 30158 130 30324
rect 150 30158 154 30324
rect 174 30158 178 30324
rect 198 30158 202 30324
rect 211 30317 216 30324
rect 221 30303 226 30317
rect 222 30158 226 30303
rect 246 30275 250 30492
rect 246 30254 253 30275
rect 270 30254 274 30492
rect 294 30254 298 30492
rect 318 30254 322 30492
rect 342 30254 346 30492
rect 366 30254 370 30492
rect 390 30254 394 30492
rect 414 30254 418 30492
rect 438 30254 442 30492
rect 462 30254 466 30492
rect 486 30254 490 30492
rect 510 30254 514 30492
rect 534 30254 538 30492
rect 558 30254 562 30492
rect 582 30254 586 30492
rect 606 30254 610 30492
rect 630 30254 634 30492
rect 654 30254 658 30492
rect 678 30254 682 30492
rect 702 30254 706 30492
rect 726 30254 730 30492
rect 750 30254 754 30492
rect 774 30254 778 30492
rect 798 30254 802 30492
rect 822 30254 826 30492
rect 846 30254 850 30492
rect 870 30254 874 30492
rect 894 30254 898 30492
rect 918 30254 922 30492
rect 942 30254 946 30492
rect 966 30254 970 30492
rect 990 30254 994 30492
rect 1014 30254 1018 30492
rect 1038 30254 1042 30492
rect 1062 30254 1066 30492
rect 1086 30254 1090 30492
rect 1110 30254 1114 30492
rect 1134 30254 1138 30492
rect 1158 30254 1162 30492
rect 1182 30254 1186 30492
rect 1206 30254 1210 30492
rect 1230 30254 1234 30492
rect 1254 30254 1258 30492
rect 1278 30254 1282 30492
rect 1302 30254 1306 30492
rect 1326 30254 1330 30492
rect 1350 30254 1354 30492
rect 1374 30254 1378 30492
rect 1398 30254 1402 30492
rect 1422 30254 1426 30492
rect 1446 30254 1450 30492
rect 1470 30254 1474 30492
rect 1494 30254 1498 30492
rect 1518 30254 1522 30492
rect 1542 30254 1546 30492
rect 1566 30254 1570 30492
rect 1590 30254 1594 30492
rect 1614 30254 1618 30492
rect 1638 30254 1642 30492
rect 1662 30254 1666 30492
rect 1686 30254 1690 30492
rect 1710 30254 1714 30492
rect 1734 30254 1738 30492
rect 1758 30254 1762 30492
rect 1782 30254 1786 30492
rect 1806 30254 1810 30492
rect 1830 30254 1834 30492
rect 1854 30254 1858 30492
rect 1878 30254 1882 30492
rect 1902 30254 1906 30492
rect 1926 30254 1930 30492
rect 1950 30254 1954 30492
rect 1974 30254 1978 30492
rect 1987 30269 1992 30279
rect 1998 30269 2002 30492
rect 2011 30485 2016 30492
rect 2022 30485 2026 30492
rect 2029 30491 2043 30492
rect 2021 30471 2026 30485
rect 2035 30481 2043 30485
rect 2029 30471 2035 30481
rect 2011 30413 2016 30423
rect 2419 30413 2424 30423
rect 2659 30413 2664 30423
rect 2899 30413 2904 30423
rect 3139 30413 3144 30423
rect 3859 30413 3864 30423
rect 4099 30413 4104 30423
rect 4339 30413 4344 30423
rect 4579 30413 4584 30423
rect 4819 30413 4824 30423
rect 7219 30413 7224 30423
rect 10099 30413 10104 30423
rect 10339 30413 10344 30423
rect 10579 30413 10584 30423
rect 10819 30413 10824 30423
rect 11059 30413 11064 30423
rect 11299 30413 11304 30423
rect 2021 30399 2026 30413
rect 2035 30409 2043 30413
rect 2029 30399 2035 30409
rect 2429 30399 2434 30413
rect 2669 30399 2674 30413
rect 2909 30399 2914 30413
rect 3149 30399 3154 30413
rect 3869 30399 3874 30413
rect 4109 30399 4114 30413
rect 4349 30399 4354 30413
rect 4589 30399 4594 30413
rect 4829 30399 4834 30413
rect 7229 30399 7234 30413
rect 10109 30399 10114 30413
rect 10349 30399 10354 30413
rect 10589 30399 10594 30413
rect 10829 30399 10834 30413
rect 11069 30399 11074 30413
rect 11309 30399 11314 30413
rect 2011 30341 2016 30351
rect 2021 30327 2026 30341
rect 2035 30337 2043 30341
rect 2029 30327 2035 30337
rect 2011 30293 2016 30303
rect 2022 30293 2026 30327
rect 2406 30323 2413 30347
rect 2646 30323 2653 30347
rect 2886 30323 2893 30347
rect 3126 30323 3133 30347
rect 3846 30323 3853 30347
rect 4086 30323 4093 30347
rect 4326 30323 4333 30347
rect 4566 30323 4573 30347
rect 4806 30323 4813 30347
rect 7206 30323 7213 30347
rect 10086 30323 10093 30347
rect 10326 30323 10333 30347
rect 10566 30323 10573 30347
rect 10806 30323 10813 30347
rect 11046 30323 11053 30347
rect 11286 30323 11293 30347
rect 2021 30279 2026 30293
rect 1997 30255 2002 30269
rect 1987 30254 2021 30255
rect 229 30252 2021 30254
rect 229 30251 243 30252
rect 246 30227 253 30252
rect 246 30158 250 30227
rect 270 30158 274 30252
rect 294 30158 298 30252
rect 318 30158 322 30252
rect 342 30158 346 30252
rect 366 30158 370 30252
rect 390 30158 394 30252
rect 414 30158 418 30252
rect 438 30158 442 30252
rect 462 30158 466 30252
rect 486 30158 490 30252
rect 510 30158 514 30252
rect 534 30158 538 30252
rect 558 30158 562 30252
rect 582 30158 586 30252
rect 606 30158 610 30252
rect 630 30158 634 30252
rect 654 30158 658 30252
rect 678 30158 682 30252
rect 702 30158 706 30252
rect 726 30158 730 30252
rect 750 30158 754 30252
rect 774 30158 778 30252
rect 798 30158 802 30252
rect 822 30158 826 30252
rect 846 30158 850 30252
rect 870 30158 874 30252
rect 894 30158 898 30252
rect 918 30158 922 30252
rect 942 30158 946 30252
rect 966 30158 970 30252
rect 990 30158 994 30252
rect 1014 30158 1018 30252
rect 1038 30158 1042 30252
rect 1062 30158 1066 30252
rect 1086 30158 1090 30252
rect 1110 30158 1114 30252
rect 1134 30158 1138 30252
rect 1158 30158 1162 30252
rect 1182 30158 1186 30252
rect 1206 30158 1210 30252
rect 1230 30158 1234 30252
rect 1254 30158 1258 30252
rect 1278 30158 1282 30252
rect 1302 30158 1306 30252
rect 1326 30158 1330 30252
rect 1350 30158 1354 30252
rect 1374 30158 1378 30252
rect 1398 30158 1402 30252
rect 1422 30158 1426 30252
rect 1446 30158 1450 30252
rect 1470 30158 1474 30252
rect 1494 30158 1498 30252
rect 1518 30158 1522 30252
rect 1542 30158 1546 30252
rect 1566 30158 1570 30252
rect 1590 30158 1594 30252
rect 1614 30158 1618 30252
rect 1638 30158 1642 30252
rect 1662 30158 1666 30252
rect 1686 30158 1690 30252
rect 1710 30158 1714 30252
rect 1734 30158 1738 30252
rect 1758 30158 1762 30252
rect 1782 30158 1786 30252
rect 1806 30158 1810 30252
rect 1830 30158 1834 30252
rect 1854 30158 1858 30252
rect 1878 30159 1882 30252
rect 1867 30158 1901 30159
rect -755 30156 1901 30158
rect -755 30155 -741 30156
rect -738 30131 -731 30156
rect -738 30062 -734 30131
rect -714 30062 -710 30156
rect -690 30062 -686 30156
rect -666 30062 -662 30156
rect -642 30062 -638 30156
rect -618 30062 -614 30156
rect -594 30062 -590 30156
rect -570 30062 -566 30156
rect -546 30062 -542 30156
rect -522 30107 -518 30156
rect -522 30083 -515 30107
rect -522 30062 -518 30083
rect -498 30062 -494 30156
rect -474 30062 -470 30156
rect -450 30062 -446 30156
rect -426 30062 -422 30156
rect -402 30062 -398 30156
rect -378 30062 -374 30156
rect -354 30062 -350 30156
rect -330 30062 -326 30156
rect -306 30062 -302 30156
rect -282 30062 -278 30156
rect -258 30062 -254 30156
rect -234 30062 -230 30156
rect -210 30062 -206 30156
rect -186 30062 -182 30156
rect -162 30062 -158 30156
rect -138 30062 -134 30156
rect -114 30062 -110 30156
rect -90 30062 -86 30156
rect -66 30062 -62 30156
rect -42 30062 -38 30156
rect -18 30062 -14 30156
rect 6 30062 10 30156
rect 30 30062 34 30156
rect 54 30062 58 30156
rect 78 30062 82 30156
rect 102 30062 106 30156
rect 126 30062 130 30156
rect 150 30062 154 30156
rect 174 30062 178 30156
rect 198 30062 202 30156
rect 222 30062 226 30156
rect 246 30062 250 30156
rect 270 30062 274 30156
rect 294 30062 298 30156
rect 318 30062 322 30156
rect 342 30062 346 30156
rect 366 30062 370 30156
rect 390 30062 394 30156
rect 414 30062 418 30156
rect 438 30062 442 30156
rect 462 30062 466 30156
rect 486 30062 490 30156
rect 510 30062 514 30156
rect 534 30062 538 30156
rect 558 30062 562 30156
rect 582 30062 586 30156
rect 606 30062 610 30156
rect 630 30062 634 30156
rect 654 30062 658 30156
rect 678 30062 682 30156
rect 702 30062 706 30156
rect 726 30062 730 30156
rect 750 30062 754 30156
rect 774 30062 778 30156
rect 798 30062 802 30156
rect 822 30062 826 30156
rect 846 30062 850 30156
rect 870 30062 874 30156
rect 894 30062 898 30156
rect 907 30125 912 30135
rect 918 30125 922 30156
rect 917 30111 922 30125
rect 907 30101 912 30111
rect 917 30087 922 30101
rect 918 30062 922 30087
rect 942 30062 946 30156
rect 966 30062 970 30156
rect 990 30062 994 30156
rect 1014 30062 1018 30156
rect 1038 30062 1042 30156
rect 1062 30062 1066 30156
rect 1086 30062 1090 30156
rect 1110 30062 1114 30156
rect 1134 30062 1138 30156
rect 1158 30062 1162 30156
rect 1182 30062 1186 30156
rect 1206 30062 1210 30156
rect 1230 30062 1234 30156
rect 1254 30062 1258 30156
rect 1278 30062 1282 30156
rect 1302 30062 1306 30156
rect 1326 30062 1330 30156
rect 1350 30062 1354 30156
rect 1374 30062 1378 30156
rect 1398 30062 1402 30156
rect 1422 30062 1426 30156
rect 1446 30062 1450 30156
rect 1470 30062 1474 30156
rect 1494 30062 1498 30156
rect 1518 30062 1522 30156
rect 1542 30062 1546 30156
rect 1566 30062 1570 30156
rect 1590 30062 1594 30156
rect 1614 30062 1618 30156
rect 1638 30062 1642 30156
rect 1662 30062 1666 30156
rect 1686 30062 1690 30156
rect 1710 30062 1714 30156
rect 1734 30062 1738 30156
rect 1758 30062 1762 30156
rect 1782 30062 1786 30156
rect 1806 30062 1810 30156
rect 1830 30062 1834 30156
rect 1854 30062 1858 30156
rect 1867 30149 1872 30156
rect 1878 30149 1882 30156
rect 1877 30135 1882 30149
rect 1878 30062 1882 30135
rect 1902 30083 1906 30252
rect -2393 30060 1899 30062
rect -2371 30014 -2366 30060
rect -2348 30014 -2343 30060
rect -2325 30014 -2320 30060
rect -2317 30056 -2309 30060
rect -2105 30053 -2092 30056
rect -2092 30030 -2062 30032
rect -2094 30026 -2062 30030
rect -2000 30014 -1992 30060
rect -1663 30056 -1655 30060
rect -1969 30053 -1921 30056
rect -1854 30030 -1806 30032
rect -1854 30026 -1680 30030
rect -1642 30014 -1637 30060
rect -1619 30014 -1614 30060
rect -1530 30014 -1526 30060
rect -1517 30029 -1512 30039
rect -1506 30029 -1502 30060
rect -1507 30015 -1502 30029
rect -1517 30014 -1483 30015
rect -2393 30012 -1483 30014
rect -2371 29966 -2366 30012
rect -2348 29966 -2343 30012
rect -2325 29966 -2320 30012
rect -2309 29996 -2301 30006
rect -2317 29990 -2309 29996
rect -2097 29990 -2095 29999
rect -2309 29968 -2301 29978
rect -2097 29976 -2095 29980
rect -2292 29975 -2095 29976
rect -2097 29973 -2095 29975
rect -2084 29968 -2083 30011
rect -2069 30004 -2054 30006
rect -2054 29988 -2018 29990
rect -2054 29986 -2004 29988
rect -2059 29982 -2045 29986
rect -2054 29980 -2049 29982
rect -2317 29966 -2309 29968
rect -2084 29966 -2054 29968
rect -2044 29966 -2039 29980
rect -2025 29970 -2014 29976
rect -2000 29970 -1992 30012
rect -1920 30010 -1906 30012
rect -1977 29995 -1929 30001
rect -1655 29996 -1647 30006
rect -1977 29985 -1966 29995
rect -1663 29990 -1655 29996
rect -1977 29973 -1929 29975
rect -2033 29966 -1992 29970
rect -1655 29968 -1647 29978
rect -1663 29966 -1655 29968
rect -1642 29966 -1637 30012
rect -1619 29966 -1614 30012
rect -1530 29966 -1526 30012
rect -1517 30005 -1512 30012
rect -1507 29991 -1502 30005
rect -1506 29966 -1502 29991
rect -1482 29966 -1478 30060
rect -1458 29966 -1454 30060
rect -1434 29966 -1430 30060
rect -1410 29966 -1406 30060
rect -1386 29966 -1382 30060
rect -1362 29966 -1358 30060
rect -1338 29966 -1334 30060
rect -1314 29966 -1310 30060
rect -1290 29966 -1286 30060
rect -1266 29966 -1262 30060
rect -1242 29966 -1238 30060
rect -1218 29966 -1214 30060
rect -1194 29966 -1190 30060
rect -1170 29966 -1166 30060
rect -1146 29966 -1142 30060
rect -1122 29966 -1118 30060
rect -1098 29966 -1094 30060
rect -1074 29966 -1070 30060
rect -1050 29966 -1046 30060
rect -1026 29966 -1022 30060
rect -1002 29966 -998 30060
rect -978 29966 -974 30060
rect -954 29966 -950 30060
rect -930 30011 -926 30060
rect -930 29987 -923 30011
rect -930 29966 -926 29987
rect -906 29966 -902 30060
rect -882 29966 -878 30060
rect -858 29966 -854 30060
rect -834 29966 -830 30060
rect -810 29966 -806 30060
rect -786 29966 -782 30060
rect -762 29966 -758 30060
rect -738 29966 -734 30060
rect -714 29966 -710 30060
rect -690 29966 -686 30060
rect -666 29966 -662 30060
rect -642 29966 -638 30060
rect -618 29966 -614 30060
rect -594 29966 -590 30060
rect -570 29966 -566 30060
rect -546 29966 -542 30060
rect -522 29967 -518 30060
rect -533 29966 -499 29967
rect -2393 29964 -499 29966
rect -2371 29870 -2366 29964
rect -2348 29870 -2343 29964
rect -2325 29930 -2320 29964
rect -2317 29962 -2309 29964
rect -2084 29951 -2083 29964
rect -2084 29950 -2054 29951
rect -2325 29922 -2317 29930
rect -2325 29870 -2320 29922
rect -2317 29914 -2309 29922
rect -2117 29913 -2095 29923
rect -2045 29920 -2037 29934
rect -2309 29874 -2301 29884
rect -2087 29880 -2076 29888
rect -2017 29884 -2015 29891
rect -2317 29870 -2309 29874
rect -2092 29872 -2087 29880
rect -2092 29870 -2077 29871
rect -2000 29870 -1992 29964
rect -1663 29962 -1655 29964
rect -1969 29913 -1929 29925
rect -1671 29922 -1663 29930
rect -1663 29914 -1655 29922
rect -1655 29874 -1647 29884
rect -1928 29870 -1924 29871
rect -1854 29870 -1680 29871
rect -1663 29870 -1655 29874
rect -1642 29870 -1637 29964
rect -1619 29870 -1614 29964
rect -1530 29870 -1526 29964
rect -1506 29870 -1502 29964
rect -1482 29963 -1478 29964
rect -1482 29942 -1475 29963
rect -1458 29942 -1454 29964
rect -1434 29942 -1430 29964
rect -1410 29942 -1406 29964
rect -1386 29942 -1382 29964
rect -1362 29942 -1358 29964
rect -1338 29942 -1334 29964
rect -1314 29942 -1310 29964
rect -1290 29942 -1286 29964
rect -1266 29942 -1262 29964
rect -1242 29942 -1238 29964
rect -1218 29942 -1214 29964
rect -1194 29942 -1190 29964
rect -1170 29942 -1166 29964
rect -1146 29942 -1142 29964
rect -1122 29942 -1118 29964
rect -1098 29942 -1094 29964
rect -1074 29942 -1070 29964
rect -1050 29942 -1046 29964
rect -1026 29942 -1022 29964
rect -1002 29942 -998 29964
rect -978 29942 -974 29964
rect -954 29942 -950 29964
rect -930 29942 -926 29964
rect -906 29942 -902 29964
rect -882 29942 -878 29964
rect -858 29942 -854 29964
rect -834 29942 -830 29964
rect -810 29942 -806 29964
rect -786 29942 -782 29964
rect -762 29942 -758 29964
rect -738 29942 -734 29964
rect -714 29942 -710 29964
rect -690 29942 -686 29964
rect -666 29942 -662 29964
rect -642 29942 -638 29964
rect -618 29942 -614 29964
rect -594 29942 -590 29964
rect -570 29942 -566 29964
rect -546 29942 -542 29964
rect -533 29957 -528 29964
rect -522 29957 -518 29964
rect -523 29943 -518 29957
rect -522 29942 -518 29943
rect -498 29942 -494 30060
rect -474 29942 -470 30060
rect -450 29942 -446 30060
rect -426 29942 -422 30060
rect -402 29942 -398 30060
rect -378 29942 -374 30060
rect -354 29942 -350 30060
rect -330 29942 -326 30060
rect -306 29942 -302 30060
rect -282 29942 -278 30060
rect -258 29942 -254 30060
rect -234 29942 -230 30060
rect -210 29942 -206 30060
rect -186 29942 -182 30060
rect -162 29942 -158 30060
rect -138 29942 -134 30060
rect -114 29942 -110 30060
rect -90 29942 -86 30060
rect -66 29942 -62 30060
rect -42 29942 -38 30060
rect -18 29942 -14 30060
rect 6 29942 10 30060
rect 30 29942 34 30060
rect 54 29942 58 30060
rect 78 29942 82 30060
rect 102 29942 106 30060
rect 126 29942 130 30060
rect 150 29942 154 30060
rect 174 29943 178 30060
rect 163 29942 197 29943
rect -1499 29940 197 29942
rect -1499 29939 -1485 29940
rect -1482 29915 -1475 29940
rect -1482 29870 -1478 29915
rect -1458 29870 -1454 29940
rect -1434 29870 -1430 29940
rect -1410 29870 -1406 29940
rect -1386 29870 -1382 29940
rect -1362 29870 -1358 29940
rect -1338 29870 -1334 29940
rect -1314 29870 -1310 29940
rect -1290 29870 -1286 29940
rect -1266 29870 -1262 29940
rect -1242 29870 -1238 29940
rect -1218 29870 -1214 29940
rect -1194 29870 -1190 29940
rect -1170 29870 -1166 29940
rect -1146 29870 -1142 29940
rect -1122 29870 -1118 29940
rect -1098 29870 -1094 29940
rect -1074 29870 -1070 29940
rect -1050 29870 -1046 29940
rect -1026 29870 -1022 29940
rect -1002 29870 -998 29940
rect -978 29870 -974 29940
rect -954 29870 -950 29940
rect -930 29870 -926 29940
rect -906 29870 -902 29940
rect -882 29870 -878 29940
rect -858 29870 -854 29940
rect -834 29870 -830 29940
rect -810 29870 -806 29940
rect -786 29870 -782 29940
rect -762 29870 -758 29940
rect -738 29870 -734 29940
rect -714 29870 -710 29940
rect -690 29870 -686 29940
rect -666 29870 -662 29940
rect -642 29870 -638 29940
rect -618 29870 -614 29940
rect -594 29870 -590 29940
rect -570 29870 -566 29940
rect -546 29870 -542 29940
rect -522 29870 -518 29940
rect -498 29891 -494 29940
rect -2393 29868 -501 29870
rect -2371 29846 -2366 29868
rect -2348 29846 -2343 29868
rect -2325 29846 -2320 29868
rect -2092 29863 -2037 29868
rect -2021 29863 -1969 29868
rect -1921 29863 -1913 29868
rect -1854 29864 -1680 29868
rect -2100 29861 -2092 29862
rect -2309 29846 -2301 29856
rect -2100 29855 -2087 29861
rect -2051 29848 -2026 29850
rect -2062 29846 -2012 29848
rect -2000 29846 -1992 29863
rect -1969 29855 -1921 29862
rect -1969 29846 -1964 29855
rect -1864 29846 -1796 29847
rect -1655 29846 -1647 29856
rect -1642 29846 -1637 29868
rect -1619 29846 -1614 29868
rect -1530 29846 -1526 29868
rect -1506 29846 -1502 29868
rect -1482 29846 -1478 29868
rect -1458 29846 -1454 29868
rect -1434 29846 -1430 29868
rect -1410 29846 -1406 29868
rect -1386 29846 -1382 29868
rect -1362 29846 -1358 29868
rect -1338 29846 -1334 29868
rect -1314 29846 -1310 29868
rect -1290 29846 -1286 29868
rect -1266 29846 -1262 29868
rect -1242 29846 -1238 29868
rect -1218 29846 -1214 29868
rect -1194 29846 -1190 29868
rect -1170 29846 -1166 29868
rect -1146 29846 -1142 29868
rect -1122 29846 -1118 29868
rect -1098 29846 -1094 29868
rect -1074 29846 -1070 29868
rect -1050 29846 -1046 29868
rect -1026 29846 -1022 29868
rect -1002 29846 -998 29868
rect -978 29846 -974 29868
rect -954 29846 -950 29868
rect -930 29846 -926 29868
rect -906 29846 -902 29868
rect -882 29846 -878 29868
rect -858 29846 -854 29868
rect -834 29846 -830 29868
rect -810 29846 -806 29868
rect -786 29846 -782 29868
rect -762 29846 -758 29868
rect -738 29846 -734 29868
rect -714 29846 -710 29868
rect -690 29846 -686 29868
rect -666 29846 -662 29868
rect -642 29846 -638 29868
rect -618 29846 -614 29868
rect -594 29846 -590 29868
rect -570 29846 -566 29868
rect -546 29846 -542 29868
rect -522 29846 -518 29868
rect -515 29867 -501 29868
rect -498 29867 -491 29891
rect -498 29846 -494 29867
rect -474 29846 -470 29940
rect -450 29846 -446 29940
rect -426 29846 -422 29940
rect -402 29846 -398 29940
rect -378 29846 -374 29940
rect -354 29846 -350 29940
rect -330 29846 -326 29940
rect -306 29846 -302 29940
rect -282 29846 -278 29940
rect -258 29846 -254 29940
rect -234 29846 -230 29940
rect -210 29846 -206 29940
rect -186 29846 -182 29940
rect -162 29846 -158 29940
rect -138 29846 -134 29940
rect -114 29846 -110 29940
rect -90 29846 -86 29940
rect -66 29846 -62 29940
rect -42 29846 -38 29940
rect -18 29846 -14 29940
rect 6 29846 10 29940
rect 30 29846 34 29940
rect 54 29846 58 29940
rect 78 29846 82 29940
rect 102 29846 106 29940
rect 126 29846 130 29940
rect 150 29846 154 29940
rect 163 29933 168 29940
rect 174 29933 178 29940
rect 173 29919 178 29933
rect 174 29846 178 29919
rect 198 29867 202 30060
rect -2393 29844 195 29846
rect -2371 29798 -2366 29844
rect -2348 29798 -2343 29844
rect -2325 29798 -2320 29844
rect -2317 29840 -2309 29844
rect -2105 29837 -2092 29840
rect -2092 29814 -2062 29816
rect -2094 29810 -2062 29814
rect -2000 29798 -1992 29844
rect -1663 29840 -1655 29844
rect -1969 29837 -1921 29840
rect -1854 29814 -1806 29816
rect -1854 29810 -1680 29814
rect -1926 29798 -1892 29801
rect -1642 29798 -1637 29844
rect -1619 29798 -1614 29844
rect -1530 29798 -1526 29844
rect -1506 29798 -1502 29844
rect -1482 29798 -1478 29844
rect -1458 29798 -1454 29844
rect -1434 29798 -1430 29844
rect -1410 29798 -1406 29844
rect -1386 29798 -1382 29844
rect -1362 29798 -1358 29844
rect -1338 29798 -1334 29844
rect -1314 29798 -1310 29844
rect -1290 29798 -1286 29844
rect -1266 29798 -1262 29844
rect -1242 29798 -1238 29844
rect -1218 29798 -1214 29844
rect -1194 29798 -1190 29844
rect -1170 29798 -1166 29844
rect -1146 29798 -1142 29844
rect -1122 29798 -1118 29844
rect -1098 29798 -1094 29844
rect -1074 29798 -1070 29844
rect -1050 29798 -1046 29844
rect -1026 29798 -1022 29844
rect -1002 29798 -998 29844
rect -978 29798 -974 29844
rect -954 29798 -950 29844
rect -930 29798 -926 29844
rect -906 29798 -902 29844
rect -882 29798 -878 29844
rect -858 29798 -854 29844
rect -834 29798 -830 29844
rect -810 29798 -806 29844
rect -786 29798 -782 29844
rect -762 29798 -758 29844
rect -738 29798 -734 29844
rect -714 29798 -710 29844
rect -690 29798 -686 29844
rect -666 29798 -662 29844
rect -642 29798 -638 29844
rect -618 29798 -614 29844
rect -594 29798 -590 29844
rect -570 29798 -566 29844
rect -546 29798 -542 29844
rect -522 29798 -518 29844
rect -498 29798 -494 29844
rect -474 29798 -470 29844
rect -450 29798 -446 29844
rect -426 29798 -422 29844
rect -402 29798 -398 29844
rect -378 29798 -374 29844
rect -354 29798 -350 29844
rect -330 29798 -326 29844
rect -306 29798 -302 29844
rect -282 29798 -278 29844
rect -258 29798 -254 29844
rect -234 29798 -230 29844
rect -210 29798 -206 29844
rect -186 29798 -182 29844
rect -162 29798 -158 29844
rect -138 29798 -134 29844
rect -114 29798 -110 29844
rect -90 29798 -86 29844
rect -66 29798 -62 29844
rect -42 29798 -38 29844
rect -18 29798 -14 29844
rect 6 29798 10 29844
rect 30 29798 34 29844
rect 54 29798 58 29844
rect 78 29798 82 29844
rect 102 29798 106 29844
rect 126 29798 130 29844
rect 139 29813 144 29823
rect 150 29813 154 29844
rect 149 29799 154 29813
rect 139 29798 173 29799
rect -2393 29796 173 29798
rect -2371 29774 -2366 29796
rect -2348 29774 -2343 29796
rect -2325 29774 -2320 29796
rect -2054 29795 -1906 29796
rect -2054 29794 -2036 29795
rect -2309 29780 -2301 29790
rect -2317 29774 -2309 29780
rect -2068 29779 -2038 29786
rect -2000 29778 -1992 29795
rect -1920 29794 -1906 29795
rect -1846 29788 -1794 29796
rect -1852 29781 -1804 29786
rect -1902 29779 -1804 29781
rect -1655 29780 -1647 29790
rect -2000 29776 -1975 29778
rect -1902 29777 -1852 29779
rect -2025 29774 -1975 29776
rect -1846 29774 -1804 29777
rect -1663 29774 -1655 29780
rect -1642 29774 -1637 29796
rect -1619 29774 -1614 29796
rect -1530 29774 -1526 29796
rect -1506 29774 -1502 29796
rect -1482 29774 -1478 29796
rect -1458 29774 -1454 29796
rect -1434 29774 -1430 29796
rect -1410 29774 -1406 29796
rect -1386 29774 -1382 29796
rect -1362 29774 -1358 29796
rect -1338 29774 -1334 29796
rect -1314 29774 -1310 29796
rect -1290 29774 -1286 29796
rect -1266 29774 -1262 29796
rect -1242 29774 -1238 29796
rect -1218 29775 -1214 29796
rect -1229 29774 -1195 29775
rect -2393 29772 -1195 29774
rect -2371 29750 -2366 29772
rect -2348 29750 -2343 29772
rect -2325 29750 -2320 29772
rect -2054 29771 -2038 29772
rect -2000 29771 -1966 29772
rect -1846 29771 -1804 29772
rect -2000 29770 -1975 29771
rect -2076 29762 -2054 29769
rect -2309 29752 -2301 29762
rect -2044 29759 -2038 29764
rect -2028 29762 -2001 29769
rect -2054 29752 -2038 29759
rect -2015 29761 -2001 29762
rect -2015 29752 -2014 29761
rect -2317 29750 -2309 29752
rect -2044 29750 -2028 29752
rect -2000 29750 -1992 29770
rect -1982 29769 -1975 29770
rect -1862 29769 -1798 29770
rect -1985 29762 -1796 29769
rect -1862 29761 -1798 29762
rect -1852 29752 -1804 29759
rect -1655 29752 -1647 29762
rect -1976 29750 -1940 29751
rect -1663 29750 -1655 29752
rect -1642 29750 -1637 29772
rect -1619 29750 -1614 29772
rect -1530 29750 -1526 29772
rect -1506 29750 -1502 29772
rect -1482 29750 -1478 29772
rect -1458 29750 -1454 29772
rect -1434 29750 -1430 29772
rect -1410 29750 -1406 29772
rect -1386 29750 -1382 29772
rect -1362 29750 -1358 29772
rect -1338 29750 -1334 29772
rect -1314 29750 -1310 29772
rect -1290 29750 -1286 29772
rect -1266 29750 -1262 29772
rect -1242 29750 -1238 29772
rect -1229 29765 -1224 29772
rect -1218 29765 -1214 29772
rect -1219 29751 -1214 29765
rect -1218 29750 -1214 29751
rect -1194 29750 -1190 29796
rect -1170 29750 -1166 29796
rect -1146 29750 -1142 29796
rect -1122 29750 -1118 29796
rect -1098 29750 -1094 29796
rect -1074 29750 -1070 29796
rect -1050 29750 -1046 29796
rect -1026 29750 -1022 29796
rect -1002 29750 -998 29796
rect -978 29750 -974 29796
rect -954 29750 -950 29796
rect -930 29750 -926 29796
rect -906 29750 -902 29796
rect -882 29750 -878 29796
rect -858 29750 -854 29796
rect -834 29750 -830 29796
rect -810 29750 -806 29796
rect -786 29750 -782 29796
rect -762 29750 -758 29796
rect -738 29750 -734 29796
rect -714 29750 -710 29796
rect -690 29750 -686 29796
rect -666 29750 -662 29796
rect -642 29750 -638 29796
rect -618 29750 -614 29796
rect -594 29750 -590 29796
rect -570 29750 -566 29796
rect -546 29750 -542 29796
rect -522 29750 -518 29796
rect -498 29750 -494 29796
rect -474 29750 -470 29796
rect -450 29750 -446 29796
rect -426 29750 -422 29796
rect -402 29750 -398 29796
rect -378 29750 -374 29796
rect -354 29750 -350 29796
rect -330 29750 -326 29796
rect -306 29750 -302 29796
rect -282 29750 -278 29796
rect -258 29750 -254 29796
rect -234 29750 -230 29796
rect -210 29750 -206 29796
rect -186 29750 -182 29796
rect -162 29750 -158 29796
rect -138 29750 -134 29796
rect -114 29750 -110 29796
rect -90 29750 -86 29796
rect -66 29750 -62 29796
rect -42 29750 -38 29796
rect -18 29750 -14 29796
rect 6 29750 10 29796
rect 30 29750 34 29796
rect 54 29750 58 29796
rect 78 29750 82 29796
rect 102 29750 106 29796
rect 126 29750 130 29796
rect 139 29789 144 29796
rect 149 29775 154 29789
rect 150 29750 154 29775
rect 174 29750 178 29844
rect 181 29843 195 29844
rect 198 29843 205 29867
rect 198 29750 202 29843
rect 222 29750 226 30060
rect 246 29750 250 30060
rect 270 29750 274 30060
rect 294 29750 298 30060
rect 318 29750 322 30060
rect 342 29750 346 30060
rect 366 29750 370 30060
rect 379 29861 384 29871
rect 390 29861 394 30060
rect 389 29847 394 29861
rect 390 29750 394 29847
rect 414 29795 418 30060
rect 414 29771 421 29795
rect 414 29750 418 29771
rect 438 29750 442 30060
rect 462 29750 466 30060
rect 486 29750 490 30060
rect 510 29750 514 30060
rect 534 29750 538 30060
rect 558 29750 562 30060
rect 582 29750 586 30060
rect 606 29750 610 30060
rect 630 29750 634 30060
rect 654 29750 658 30060
rect 678 29750 682 30060
rect 702 29750 706 30060
rect 726 29750 730 30060
rect 750 29750 754 30060
rect 774 29750 778 30060
rect 798 29750 802 30060
rect 822 29750 826 30060
rect 846 29750 850 30060
rect 870 29750 874 30060
rect 894 29750 898 30060
rect 918 29750 922 30060
rect 942 30059 946 30060
rect 942 30038 949 30059
rect 966 30038 970 30060
rect 990 30038 994 30060
rect 1014 30038 1018 30060
rect 1038 30038 1042 30060
rect 1062 30038 1066 30060
rect 1086 30038 1090 30060
rect 1110 30038 1114 30060
rect 1134 30038 1138 30060
rect 1158 30038 1162 30060
rect 1182 30038 1186 30060
rect 1206 30038 1210 30060
rect 1230 30038 1234 30060
rect 1254 30038 1258 30060
rect 1278 30038 1282 30060
rect 1302 30038 1306 30060
rect 1326 30038 1330 30060
rect 1350 30038 1354 30060
rect 1374 30038 1378 30060
rect 1398 30038 1402 30060
rect 1422 30038 1426 30060
rect 1446 30038 1450 30060
rect 1470 30038 1474 30060
rect 1494 30038 1498 30060
rect 1518 30038 1522 30060
rect 1542 30038 1546 30060
rect 1566 30038 1570 30060
rect 1590 30038 1594 30060
rect 1614 30038 1618 30060
rect 1638 30038 1642 30060
rect 1662 30038 1666 30060
rect 1686 30038 1690 30060
rect 1710 30038 1714 30060
rect 1734 30038 1738 30060
rect 1758 30038 1762 30060
rect 1782 30038 1786 30060
rect 1806 30038 1810 30060
rect 1830 30038 1834 30060
rect 1854 30038 1858 30060
rect 1878 30038 1882 30060
rect 1885 30059 1899 30060
rect 1902 30059 1909 30083
rect 1902 30038 1906 30059
rect 1926 30038 1930 30252
rect 1950 30038 1954 30252
rect 1974 30038 1978 30252
rect 1987 30245 1992 30252
rect 1997 30231 2002 30245
rect 1998 30038 2002 30231
rect 2011 30125 2016 30135
rect 2021 30111 2026 30125
rect 2011 30053 2016 30063
rect 2022 30053 2026 30111
rect 2021 30039 2026 30053
rect 2035 30049 2043 30053
rect 2029 30039 2035 30049
rect 2011 30038 2043 30039
rect 925 30036 2043 30038
rect 925 30035 939 30036
rect 942 30011 949 30036
rect 942 29750 946 30011
rect 966 29750 970 30036
rect 990 29750 994 30036
rect 1014 29750 1018 30036
rect 1038 29750 1042 30036
rect 1062 29750 1066 30036
rect 1086 29750 1090 30036
rect 1110 29750 1114 30036
rect 1134 29750 1138 30036
rect 1158 29750 1162 30036
rect 1182 29750 1186 30036
rect 1206 29750 1210 30036
rect 1230 29750 1234 30036
rect 1254 29750 1258 30036
rect 1278 29750 1282 30036
rect 1302 29750 1306 30036
rect 1326 29750 1330 30036
rect 1350 29750 1354 30036
rect 1374 29750 1378 30036
rect 1398 29750 1402 30036
rect 1422 29750 1426 30036
rect 1446 29750 1450 30036
rect 1470 29750 1474 30036
rect 1494 29750 1498 30036
rect 1518 29750 1522 30036
rect 1531 29909 1536 29919
rect 1542 29909 1546 30036
rect 1541 29895 1546 29909
rect 1531 29885 1536 29895
rect 1541 29871 1546 29885
rect 1542 29750 1546 29871
rect 1566 29843 1570 30036
rect 1566 29822 1573 29843
rect 1590 29822 1594 30036
rect 1614 29822 1618 30036
rect 1638 29822 1642 30036
rect 1662 29822 1666 30036
rect 1686 29822 1690 30036
rect 1710 29822 1714 30036
rect 1734 29822 1738 30036
rect 1758 29822 1762 30036
rect 1782 29822 1786 30036
rect 1806 29822 1810 30036
rect 1830 29822 1834 30036
rect 1854 29822 1858 30036
rect 1878 29822 1882 30036
rect 1902 29822 1906 30036
rect 1926 29822 1930 30036
rect 1950 29822 1954 30036
rect 1974 29822 1978 30036
rect 1998 29822 2002 30036
rect 2011 30029 2016 30036
rect 2029 30035 2043 30036
rect 2021 30015 2026 30029
rect 2022 29822 2026 30015
rect 2035 29909 2040 29919
rect 2045 29895 2050 29909
rect 2035 29837 2040 29847
rect 2046 29837 2050 29895
rect 2045 29823 2050 29837
rect 2059 29833 2067 29837
rect 2053 29823 2059 29833
rect 2035 29822 2067 29823
rect 1549 29820 2067 29822
rect 1549 29819 1563 29820
rect 1566 29795 1573 29820
rect 1566 29750 1570 29795
rect 1590 29750 1594 29820
rect 1614 29750 1618 29820
rect 1638 29750 1642 29820
rect 1662 29750 1666 29820
rect 1686 29750 1690 29820
rect 1710 29750 1714 29820
rect 1734 29750 1738 29820
rect 1758 29750 1762 29820
rect 1782 29750 1786 29820
rect 1806 29750 1810 29820
rect 1830 29750 1834 29820
rect 1854 29750 1858 29820
rect 1878 29750 1882 29820
rect 1902 29750 1906 29820
rect 1926 29750 1930 29820
rect 1950 29750 1954 29820
rect 1974 29750 1978 29820
rect 1998 29750 2002 29820
rect 2022 29750 2026 29820
rect 2035 29813 2040 29820
rect 2053 29819 2067 29820
rect 2045 29799 2050 29813
rect 2046 29751 2050 29799
rect 2035 29750 2067 29751
rect -2393 29748 2067 29750
rect -2371 29678 -2366 29748
rect -2348 29678 -2343 29748
rect -2325 29714 -2320 29748
rect -2317 29746 -2309 29748
rect -2076 29735 -2054 29742
rect -2325 29706 -2317 29714
rect -2060 29708 -2030 29711
rect -2325 29678 -2320 29706
rect -2317 29698 -2309 29706
rect -2060 29695 -2038 29706
rect -2033 29699 -2030 29708
rect -2028 29704 -2027 29708
rect -2068 29690 -2038 29693
rect -2000 29678 -1992 29748
rect -1846 29744 -1804 29748
rect -1663 29746 -1655 29748
rect -1846 29734 -1794 29743
rect -1912 29723 -1884 29725
rect -1852 29717 -1804 29721
rect -1844 29708 -1796 29711
rect -1671 29706 -1663 29714
rect -1844 29695 -1804 29706
rect -1663 29698 -1655 29706
rect -1852 29690 -1680 29694
rect -1642 29678 -1637 29748
rect -1619 29678 -1614 29748
rect -1530 29678 -1526 29748
rect -1506 29678 -1502 29748
rect -1482 29678 -1478 29748
rect -1458 29678 -1454 29748
rect -1434 29678 -1430 29748
rect -1410 29678 -1406 29748
rect -1386 29678 -1382 29748
rect -1362 29678 -1358 29748
rect -1338 29678 -1334 29748
rect -1314 29678 -1310 29748
rect -1290 29678 -1286 29748
rect -1266 29678 -1262 29748
rect -1242 29678 -1238 29748
rect -1218 29678 -1214 29748
rect -1194 29699 -1190 29748
rect -2393 29676 -1197 29678
rect -2371 29654 -2366 29676
rect -2348 29654 -2343 29676
rect -2325 29654 -2320 29676
rect -2309 29658 -2301 29668
rect -2068 29659 -2062 29664
rect -2317 29654 -2309 29658
rect -2060 29654 -2050 29659
rect -2000 29654 -1992 29676
rect -1806 29668 -1680 29674
rect -1854 29659 -1806 29664
rect -1655 29658 -1647 29668
rect -1972 29654 -1964 29655
rect -1958 29654 -1942 29656
rect -1844 29654 -1806 29657
rect -1663 29654 -1655 29658
rect -1642 29654 -1637 29676
rect -1619 29654 -1614 29676
rect -1530 29654 -1526 29676
rect -1506 29654 -1502 29676
rect -1482 29654 -1478 29676
rect -1458 29654 -1454 29676
rect -1434 29654 -1430 29676
rect -1410 29654 -1406 29676
rect -1386 29654 -1382 29676
rect -1362 29654 -1358 29676
rect -1338 29654 -1334 29676
rect -1314 29654 -1310 29676
rect -1290 29654 -1286 29676
rect -1266 29654 -1262 29676
rect -1242 29654 -1238 29676
rect -1218 29654 -1214 29676
rect -1211 29675 -1197 29676
rect -1194 29675 -1187 29699
rect -1194 29654 -1190 29675
rect -1170 29654 -1166 29748
rect -1146 29654 -1142 29748
rect -1122 29654 -1118 29748
rect -1098 29654 -1094 29748
rect -1074 29654 -1070 29748
rect -1050 29654 -1046 29748
rect -1026 29654 -1022 29748
rect -1002 29654 -998 29748
rect -978 29654 -974 29748
rect -954 29654 -950 29748
rect -930 29654 -926 29748
rect -906 29654 -902 29748
rect -882 29654 -878 29748
rect -858 29654 -854 29748
rect -834 29654 -830 29748
rect -810 29654 -806 29748
rect -786 29654 -782 29748
rect -762 29654 -758 29748
rect -738 29654 -734 29748
rect -714 29654 -710 29748
rect -690 29654 -686 29748
rect -666 29654 -662 29748
rect -642 29654 -638 29748
rect -618 29654 -614 29748
rect -594 29654 -590 29748
rect -570 29654 -566 29748
rect -546 29654 -542 29748
rect -522 29654 -518 29748
rect -498 29654 -494 29748
rect -474 29654 -470 29748
rect -450 29654 -446 29748
rect -426 29654 -422 29748
rect -402 29654 -398 29748
rect -378 29654 -374 29748
rect -354 29654 -350 29748
rect -330 29654 -326 29748
rect -306 29654 -302 29748
rect -282 29654 -278 29748
rect -258 29654 -254 29748
rect -234 29654 -230 29748
rect -210 29654 -206 29748
rect -186 29654 -182 29748
rect -162 29654 -158 29748
rect -138 29654 -134 29748
rect -114 29654 -110 29748
rect -90 29654 -86 29748
rect -66 29654 -62 29748
rect -42 29654 -38 29748
rect -18 29654 -14 29748
rect 6 29654 10 29748
rect 30 29654 34 29748
rect 54 29654 58 29748
rect 78 29654 82 29748
rect 102 29654 106 29748
rect 126 29654 130 29748
rect 150 29654 154 29748
rect 174 29747 178 29748
rect 174 29726 181 29747
rect 198 29726 202 29748
rect 222 29726 226 29748
rect 246 29726 250 29748
rect 270 29726 274 29748
rect 294 29726 298 29748
rect 318 29726 322 29748
rect 342 29726 346 29748
rect 366 29726 370 29748
rect 390 29726 394 29748
rect 414 29726 418 29748
rect 438 29726 442 29748
rect 462 29726 466 29748
rect 486 29726 490 29748
rect 510 29726 514 29748
rect 534 29726 538 29748
rect 558 29726 562 29748
rect 582 29726 586 29748
rect 606 29726 610 29748
rect 630 29726 634 29748
rect 654 29726 658 29748
rect 678 29726 682 29748
rect 702 29726 706 29748
rect 726 29726 730 29748
rect 750 29726 754 29748
rect 774 29726 778 29748
rect 798 29726 802 29748
rect 822 29726 826 29748
rect 846 29726 850 29748
rect 870 29726 874 29748
rect 894 29726 898 29748
rect 918 29726 922 29748
rect 942 29726 946 29748
rect 966 29726 970 29748
rect 990 29726 994 29748
rect 1014 29726 1018 29748
rect 1038 29726 1042 29748
rect 1062 29726 1066 29748
rect 1086 29726 1090 29748
rect 1110 29726 1114 29748
rect 1134 29726 1138 29748
rect 1158 29726 1162 29748
rect 1182 29726 1186 29748
rect 1206 29726 1210 29748
rect 1230 29726 1234 29748
rect 1254 29726 1258 29748
rect 1278 29726 1282 29748
rect 1302 29726 1306 29748
rect 1326 29726 1330 29748
rect 1350 29726 1354 29748
rect 1374 29726 1378 29748
rect 1398 29726 1402 29748
rect 1422 29726 1426 29748
rect 1446 29726 1450 29748
rect 1470 29726 1474 29748
rect 1494 29726 1498 29748
rect 1518 29726 1522 29748
rect 1542 29726 1546 29748
rect 1566 29726 1570 29748
rect 1590 29726 1594 29748
rect 1614 29726 1618 29748
rect 1638 29726 1642 29748
rect 1662 29726 1666 29748
rect 1686 29726 1690 29748
rect 1710 29726 1714 29748
rect 1734 29726 1738 29748
rect 1758 29726 1762 29748
rect 1782 29726 1786 29748
rect 1806 29726 1810 29748
rect 1830 29726 1834 29748
rect 1854 29726 1858 29748
rect 1878 29726 1882 29748
rect 1902 29726 1906 29748
rect 1926 29726 1930 29748
rect 1950 29726 1954 29748
rect 1974 29726 1978 29748
rect 1998 29726 2002 29748
rect 2022 29727 2026 29748
rect 2035 29741 2040 29748
rect 2046 29741 2050 29748
rect 2053 29747 2067 29748
rect 2045 29727 2050 29741
rect 2059 29737 2067 29741
rect 2053 29727 2059 29737
rect 2011 29726 2045 29727
rect 157 29724 2045 29726
rect 157 29723 171 29724
rect 174 29699 181 29724
rect 174 29654 178 29699
rect 198 29654 202 29724
rect 222 29654 226 29724
rect 246 29654 250 29724
rect 270 29654 274 29724
rect 294 29654 298 29724
rect 318 29654 322 29724
rect 342 29654 346 29724
rect 366 29654 370 29724
rect 390 29654 394 29724
rect 414 29654 418 29724
rect 438 29654 442 29724
rect 462 29654 466 29724
rect 486 29654 490 29724
rect 510 29654 514 29724
rect 534 29654 538 29724
rect 558 29654 562 29724
rect 582 29654 586 29724
rect 606 29654 610 29724
rect 630 29654 634 29724
rect 654 29654 658 29724
rect 678 29654 682 29724
rect 702 29654 706 29724
rect 726 29654 730 29724
rect 750 29654 754 29724
rect 774 29654 778 29724
rect 798 29654 802 29724
rect 822 29654 826 29724
rect 846 29654 850 29724
rect 870 29654 874 29724
rect 894 29654 898 29724
rect 918 29654 922 29724
rect 942 29654 946 29724
rect 966 29654 970 29724
rect 990 29654 994 29724
rect 1014 29654 1018 29724
rect 1038 29654 1042 29724
rect 1062 29654 1066 29724
rect 1086 29654 1090 29724
rect 1110 29654 1114 29724
rect 1134 29654 1138 29724
rect 1158 29654 1162 29724
rect 1182 29654 1186 29724
rect 1206 29654 1210 29724
rect 1230 29654 1234 29724
rect 1254 29654 1258 29724
rect 1278 29654 1282 29724
rect 1302 29654 1306 29724
rect 1326 29654 1330 29724
rect 1350 29654 1354 29724
rect 1374 29654 1378 29724
rect 1398 29654 1402 29724
rect 1422 29654 1426 29724
rect 1446 29654 1450 29724
rect 1470 29654 1474 29724
rect 1494 29654 1498 29724
rect 1518 29654 1522 29724
rect 1542 29654 1546 29724
rect 1566 29654 1570 29724
rect 1590 29654 1594 29724
rect 1614 29654 1618 29724
rect 1638 29654 1642 29724
rect 1662 29654 1666 29724
rect 1686 29654 1690 29724
rect 1710 29654 1714 29724
rect 1734 29654 1738 29724
rect 1758 29654 1762 29724
rect 1782 29654 1786 29724
rect 1806 29654 1810 29724
rect 1830 29654 1834 29724
rect 1854 29654 1858 29724
rect 1878 29654 1882 29724
rect 1902 29654 1906 29724
rect 1926 29654 1930 29724
rect 1939 29693 1944 29703
rect 1950 29693 1954 29724
rect 1949 29679 1954 29693
rect 1939 29669 1944 29679
rect 1949 29655 1954 29669
rect 1950 29654 1954 29655
rect 1974 29654 1978 29724
rect 1998 29654 2002 29724
rect 2011 29717 2016 29724
rect 2022 29717 2026 29724
rect 2021 29703 2026 29717
rect 2011 29693 2016 29703
rect 2021 29679 2026 29693
rect 2022 29655 2026 29679
rect 2011 29654 2045 29655
rect -2393 29652 2045 29654
rect -2371 29630 -2366 29652
rect -2348 29630 -2343 29652
rect -2325 29630 -2320 29652
rect -2060 29646 -2050 29652
rect -2309 29630 -2301 29640
rect -2060 29639 -2030 29646
rect -2000 29642 -1992 29652
rect -1972 29650 -1942 29652
rect -1958 29649 -1942 29650
rect -1844 29648 -1806 29652
rect -2068 29632 -2062 29639
rect -2062 29630 -2036 29632
rect -2393 29628 -2036 29630
rect -2030 29630 -2012 29632
rect -2004 29630 -1990 29642
rect -1844 29641 -1798 29646
rect -1806 29639 -1798 29641
rect -1854 29637 -1844 29639
rect -1854 29632 -1806 29637
rect -1864 29630 -1796 29631
rect -1655 29630 -1647 29640
rect -1642 29630 -1637 29652
rect -1619 29630 -1614 29652
rect -1530 29630 -1526 29652
rect -1506 29630 -1502 29652
rect -1482 29630 -1478 29652
rect -1458 29630 -1454 29652
rect -1434 29630 -1430 29652
rect -1410 29630 -1406 29652
rect -1386 29630 -1382 29652
rect -1362 29630 -1358 29652
rect -1338 29630 -1334 29652
rect -1314 29630 -1310 29652
rect -1290 29630 -1286 29652
rect -1266 29630 -1262 29652
rect -1242 29630 -1238 29652
rect -1218 29630 -1214 29652
rect -1194 29630 -1190 29652
rect -1170 29630 -1166 29652
rect -1146 29630 -1142 29652
rect -1122 29630 -1118 29652
rect -1098 29630 -1094 29652
rect -1074 29630 -1070 29652
rect -1050 29630 -1046 29652
rect -1026 29630 -1022 29652
rect -1002 29630 -998 29652
rect -978 29630 -974 29652
rect -954 29630 -950 29652
rect -930 29630 -926 29652
rect -906 29630 -902 29652
rect -882 29630 -878 29652
rect -858 29630 -854 29652
rect -834 29630 -830 29652
rect -810 29630 -806 29652
rect -786 29630 -782 29652
rect -762 29630 -758 29652
rect -738 29630 -734 29652
rect -714 29630 -710 29652
rect -690 29630 -686 29652
rect -666 29630 -662 29652
rect -642 29630 -638 29652
rect -618 29630 -614 29652
rect -594 29630 -590 29652
rect -570 29630 -566 29652
rect -546 29630 -542 29652
rect -522 29630 -518 29652
rect -498 29630 -494 29652
rect -474 29630 -470 29652
rect -450 29630 -446 29652
rect -426 29630 -422 29652
rect -402 29630 -398 29652
rect -378 29630 -374 29652
rect -354 29630 -350 29652
rect -330 29630 -326 29652
rect -306 29630 -302 29652
rect -282 29630 -278 29652
rect -258 29630 -254 29652
rect -234 29630 -230 29652
rect -210 29630 -206 29652
rect -186 29630 -182 29652
rect -162 29630 -158 29652
rect -138 29630 -134 29652
rect -114 29630 -110 29652
rect -90 29630 -86 29652
rect -66 29630 -62 29652
rect -42 29630 -38 29652
rect -18 29630 -14 29652
rect 6 29630 10 29652
rect 30 29630 34 29652
rect 54 29630 58 29652
rect 78 29630 82 29652
rect 102 29630 106 29652
rect 126 29630 130 29652
rect 150 29630 154 29652
rect 174 29630 178 29652
rect 198 29630 202 29652
rect 222 29630 226 29652
rect 246 29630 250 29652
rect 270 29630 274 29652
rect 294 29630 298 29652
rect 318 29630 322 29652
rect 342 29630 346 29652
rect 366 29630 370 29652
rect 390 29630 394 29652
rect 414 29630 418 29652
rect 438 29630 442 29652
rect 462 29630 466 29652
rect 486 29630 490 29652
rect 510 29630 514 29652
rect 534 29630 538 29652
rect 558 29630 562 29652
rect 582 29630 586 29652
rect 606 29630 610 29652
rect 630 29630 634 29652
rect 654 29630 658 29652
rect 678 29630 682 29652
rect 702 29630 706 29652
rect 726 29630 730 29652
rect 750 29630 754 29652
rect 774 29630 778 29652
rect 798 29630 802 29652
rect 822 29630 826 29652
rect 846 29630 850 29652
rect 870 29630 874 29652
rect 894 29630 898 29652
rect 918 29630 922 29652
rect 942 29630 946 29652
rect 966 29630 970 29652
rect 990 29630 994 29652
rect 1014 29630 1018 29652
rect 1038 29630 1042 29652
rect 1062 29630 1066 29652
rect 1086 29630 1090 29652
rect 1110 29630 1114 29652
rect 1134 29630 1138 29652
rect 1158 29630 1162 29652
rect 1182 29630 1186 29652
rect 1206 29630 1210 29652
rect 1230 29630 1234 29652
rect 1254 29630 1258 29652
rect 1278 29630 1282 29652
rect 1302 29630 1306 29652
rect 1326 29630 1330 29652
rect 1350 29630 1354 29652
rect 1374 29630 1378 29652
rect 1398 29630 1402 29652
rect 1422 29630 1426 29652
rect 1446 29630 1450 29652
rect 1470 29630 1474 29652
rect 1494 29630 1498 29652
rect 1518 29630 1522 29652
rect 1542 29630 1546 29652
rect 1566 29630 1570 29652
rect 1590 29630 1594 29652
rect 1614 29630 1618 29652
rect 1638 29630 1642 29652
rect 1662 29630 1666 29652
rect 1686 29630 1690 29652
rect 1710 29630 1714 29652
rect 1734 29630 1738 29652
rect 1758 29630 1762 29652
rect 1782 29630 1786 29652
rect 1806 29630 1810 29652
rect 1830 29630 1834 29652
rect 1854 29630 1858 29652
rect 1878 29630 1882 29652
rect 1902 29630 1906 29652
rect 1926 29630 1930 29652
rect 1950 29630 1954 29652
rect 1974 29630 1978 29652
rect 1998 29631 2002 29652
rect 2011 29645 2016 29652
rect 2022 29645 2026 29652
rect 2021 29631 2026 29645
rect 2035 29641 2043 29645
rect 2029 29631 2035 29641
rect 1987 29630 2021 29631
rect -2030 29628 2021 29630
rect -2371 29582 -2366 29628
rect -2348 29582 -2343 29628
rect -2325 29582 -2320 29628
rect -2317 29624 -2309 29628
rect -2060 29624 -2050 29628
rect -2060 29622 -2036 29624
rect -2060 29620 -2030 29622
rect -2292 29614 -2030 29620
rect -2092 29598 -2062 29600
rect -2094 29594 -2062 29598
rect -2000 29582 -1992 29628
rect -1844 29621 -1806 29628
rect -1663 29624 -1655 29628
rect -1844 29614 -1680 29620
rect -1854 29598 -1806 29600
rect -1854 29594 -1680 29598
rect -1642 29582 -1637 29628
rect -1619 29582 -1614 29628
rect -1530 29582 -1526 29628
rect -1506 29582 -1502 29628
rect -1482 29582 -1478 29628
rect -1458 29582 -1454 29628
rect -1434 29582 -1430 29628
rect -1410 29582 -1406 29628
rect -1386 29582 -1382 29628
rect -1362 29582 -1358 29628
rect -1338 29582 -1334 29628
rect -1314 29582 -1310 29628
rect -1290 29582 -1286 29628
rect -1266 29582 -1262 29628
rect -1242 29582 -1238 29628
rect -1218 29582 -1214 29628
rect -1194 29582 -1190 29628
rect -1170 29582 -1166 29628
rect -1146 29582 -1142 29628
rect -1122 29582 -1118 29628
rect -1098 29582 -1094 29628
rect -1074 29582 -1070 29628
rect -1050 29582 -1046 29628
rect -1026 29582 -1022 29628
rect -1002 29582 -998 29628
rect -978 29582 -974 29628
rect -954 29582 -950 29628
rect -930 29582 -926 29628
rect -906 29582 -902 29628
rect -882 29582 -878 29628
rect -858 29582 -854 29628
rect -834 29582 -830 29628
rect -810 29582 -806 29628
rect -786 29582 -782 29628
rect -762 29582 -758 29628
rect -738 29582 -734 29628
rect -714 29582 -710 29628
rect -690 29582 -686 29628
rect -666 29582 -662 29628
rect -642 29582 -638 29628
rect -618 29582 -614 29628
rect -594 29582 -590 29628
rect -570 29582 -566 29628
rect -546 29582 -542 29628
rect -522 29582 -518 29628
rect -498 29582 -494 29628
rect -474 29582 -470 29628
rect -450 29582 -446 29628
rect -426 29582 -422 29628
rect -402 29582 -398 29628
rect -378 29582 -374 29628
rect -354 29582 -350 29628
rect -330 29582 -326 29628
rect -306 29582 -302 29628
rect -282 29582 -278 29628
rect -258 29582 -254 29628
rect -234 29582 -230 29628
rect -210 29582 -206 29628
rect -186 29582 -182 29628
rect -162 29582 -158 29628
rect -138 29582 -134 29628
rect -114 29582 -110 29628
rect -90 29582 -86 29628
rect -66 29582 -62 29628
rect -42 29582 -38 29628
rect -18 29582 -14 29628
rect 6 29582 10 29628
rect 30 29582 34 29628
rect 54 29582 58 29628
rect 78 29582 82 29628
rect 102 29582 106 29628
rect 126 29582 130 29628
rect 150 29582 154 29628
rect 174 29582 178 29628
rect 198 29582 202 29628
rect 222 29582 226 29628
rect 246 29582 250 29628
rect 270 29582 274 29628
rect 294 29582 298 29628
rect 318 29582 322 29628
rect 342 29582 346 29628
rect 366 29582 370 29628
rect 390 29582 394 29628
rect 414 29582 418 29628
rect 438 29582 442 29628
rect 462 29582 466 29628
rect 486 29582 490 29628
rect 510 29582 514 29628
rect 534 29582 538 29628
rect 558 29582 562 29628
rect 582 29582 586 29628
rect 606 29582 610 29628
rect 630 29582 634 29628
rect 654 29582 658 29628
rect 678 29582 682 29628
rect 702 29582 706 29628
rect 726 29582 730 29628
rect 750 29582 754 29628
rect 774 29582 778 29628
rect 798 29582 802 29628
rect 822 29582 826 29628
rect 846 29582 850 29628
rect 870 29582 874 29628
rect 894 29582 898 29628
rect 918 29582 922 29628
rect 942 29582 946 29628
rect 966 29582 970 29628
rect 990 29582 994 29628
rect 1014 29582 1018 29628
rect 1038 29582 1042 29628
rect 1062 29582 1066 29628
rect 1086 29582 1090 29628
rect 1110 29582 1114 29628
rect 1134 29582 1138 29628
rect 1158 29582 1162 29628
rect 1182 29582 1186 29628
rect 1206 29582 1210 29628
rect 1230 29582 1234 29628
rect 1254 29582 1258 29628
rect 1267 29597 1272 29607
rect 1278 29597 1282 29628
rect 1277 29583 1282 29597
rect 1267 29582 1301 29583
rect -2393 29580 1301 29582
rect -2371 29558 -2366 29580
rect -2348 29558 -2343 29580
rect -2325 29558 -2320 29580
rect -2072 29578 -2036 29579
rect -2072 29572 -2054 29578
rect -2309 29564 -2301 29572
rect -2317 29558 -2309 29564
rect -2092 29563 -2062 29568
rect -2000 29559 -1992 29580
rect -1938 29579 -1906 29580
rect -1920 29578 -1906 29579
rect -1806 29572 -1680 29578
rect -1854 29563 -1806 29568
rect -1655 29564 -1647 29572
rect -1982 29559 -1966 29560
rect -2000 29558 -1966 29559
rect -1846 29558 -1806 29561
rect -1663 29558 -1655 29564
rect -1642 29558 -1637 29580
rect -1619 29558 -1614 29580
rect -1530 29558 -1526 29580
rect -1506 29558 -1502 29580
rect -1482 29558 -1478 29580
rect -1458 29558 -1454 29580
rect -1434 29558 -1430 29580
rect -1410 29558 -1406 29580
rect -1386 29558 -1382 29580
rect -1362 29558 -1358 29580
rect -1338 29558 -1334 29580
rect -1314 29558 -1310 29580
rect -1290 29558 -1286 29580
rect -1266 29558 -1262 29580
rect -1242 29558 -1238 29580
rect -1218 29558 -1214 29580
rect -1194 29558 -1190 29580
rect -1170 29558 -1166 29580
rect -1146 29558 -1142 29580
rect -1122 29558 -1118 29580
rect -1098 29558 -1094 29580
rect -1074 29558 -1070 29580
rect -1050 29558 -1046 29580
rect -1026 29558 -1022 29580
rect -1002 29558 -998 29580
rect -978 29558 -974 29580
rect -954 29558 -950 29580
rect -930 29558 -926 29580
rect -906 29558 -902 29580
rect -882 29558 -878 29580
rect -858 29558 -854 29580
rect -834 29558 -830 29580
rect -810 29558 -806 29580
rect -786 29558 -782 29580
rect -762 29558 -758 29580
rect -738 29558 -734 29580
rect -714 29558 -710 29580
rect -690 29558 -686 29580
rect -666 29558 -662 29580
rect -642 29558 -638 29580
rect -618 29558 -614 29580
rect -594 29558 -590 29580
rect -570 29558 -566 29580
rect -546 29558 -542 29580
rect -522 29558 -518 29580
rect -498 29558 -494 29580
rect -474 29558 -470 29580
rect -450 29558 -446 29580
rect -426 29558 -422 29580
rect -402 29558 -398 29580
rect -378 29558 -374 29580
rect -354 29558 -350 29580
rect -330 29559 -326 29580
rect -341 29558 -307 29559
rect -2393 29556 -307 29558
rect -2371 29534 -2366 29556
rect -2348 29534 -2343 29556
rect -2325 29534 -2320 29556
rect -2000 29554 -1966 29556
rect -2309 29536 -2301 29544
rect -2062 29543 -2054 29550
rect -2092 29536 -2084 29543
rect -2062 29536 -2026 29538
rect -2317 29534 -2309 29536
rect -2062 29534 -2012 29536
rect -2000 29534 -1992 29554
rect -1982 29553 -1966 29554
rect -1846 29552 -1806 29556
rect -1846 29545 -1798 29550
rect -1806 29543 -1798 29545
rect -1854 29541 -1846 29543
rect -1854 29536 -1806 29541
rect -1655 29536 -1647 29544
rect -1864 29534 -1796 29535
rect -1663 29534 -1655 29536
rect -1642 29534 -1637 29556
rect -1619 29534 -1614 29556
rect -1530 29534 -1526 29556
rect -1506 29534 -1502 29556
rect -1482 29534 -1478 29556
rect -1458 29534 -1454 29556
rect -1434 29534 -1430 29556
rect -1410 29534 -1406 29556
rect -1386 29534 -1382 29556
rect -1362 29534 -1358 29556
rect -1338 29534 -1334 29556
rect -1314 29534 -1310 29556
rect -1290 29534 -1286 29556
rect -1266 29534 -1262 29556
rect -1242 29534 -1238 29556
rect -1218 29534 -1214 29556
rect -1194 29534 -1190 29556
rect -1170 29534 -1166 29556
rect -1146 29534 -1142 29556
rect -1122 29534 -1118 29556
rect -1098 29534 -1094 29556
rect -1074 29534 -1070 29556
rect -1050 29534 -1046 29556
rect -1026 29534 -1022 29556
rect -1002 29534 -998 29556
rect -978 29534 -974 29556
rect -954 29534 -950 29556
rect -930 29534 -926 29556
rect -906 29534 -902 29556
rect -882 29534 -878 29556
rect -858 29534 -854 29556
rect -834 29534 -830 29556
rect -810 29534 -806 29556
rect -786 29534 -782 29556
rect -762 29534 -758 29556
rect -738 29534 -734 29556
rect -714 29534 -710 29556
rect -690 29534 -686 29556
rect -666 29534 -662 29556
rect -642 29534 -638 29556
rect -618 29534 -614 29556
rect -594 29534 -590 29556
rect -570 29534 -566 29556
rect -546 29534 -542 29556
rect -522 29534 -518 29556
rect -498 29534 -494 29556
rect -474 29534 -470 29556
rect -450 29534 -446 29556
rect -426 29534 -422 29556
rect -402 29534 -398 29556
rect -378 29534 -374 29556
rect -354 29534 -350 29556
rect -341 29549 -336 29556
rect -330 29549 -326 29556
rect -331 29535 -326 29549
rect -330 29534 -326 29535
rect -306 29534 -302 29580
rect -282 29534 -278 29580
rect -258 29534 -254 29580
rect -234 29534 -230 29580
rect -210 29534 -206 29580
rect -186 29534 -182 29580
rect -162 29534 -158 29580
rect -138 29534 -134 29580
rect -114 29534 -110 29580
rect -90 29534 -86 29580
rect -66 29534 -62 29580
rect -42 29534 -38 29580
rect -18 29534 -14 29580
rect 6 29534 10 29580
rect 30 29534 34 29580
rect 54 29534 58 29580
rect 78 29534 82 29580
rect 102 29534 106 29580
rect 126 29534 130 29580
rect 150 29534 154 29580
rect 174 29534 178 29580
rect 198 29534 202 29580
rect 222 29534 226 29580
rect 246 29534 250 29580
rect 270 29534 274 29580
rect 294 29534 298 29580
rect 318 29534 322 29580
rect 342 29534 346 29580
rect 366 29534 370 29580
rect 390 29534 394 29580
rect 414 29534 418 29580
rect 438 29534 442 29580
rect 462 29534 466 29580
rect 486 29534 490 29580
rect 510 29534 514 29580
rect 534 29534 538 29580
rect 558 29534 562 29580
rect 582 29534 586 29580
rect 606 29534 610 29580
rect 630 29534 634 29580
rect 654 29534 658 29580
rect 678 29534 682 29580
rect 702 29534 706 29580
rect 726 29534 730 29580
rect 750 29534 754 29580
rect 774 29534 778 29580
rect 798 29534 802 29580
rect 822 29534 826 29580
rect 846 29534 850 29580
rect 870 29534 874 29580
rect 894 29534 898 29580
rect 918 29534 922 29580
rect 942 29534 946 29580
rect 966 29534 970 29580
rect 990 29534 994 29580
rect 1014 29534 1018 29580
rect 1038 29534 1042 29580
rect 1062 29534 1066 29580
rect 1086 29534 1090 29580
rect 1110 29534 1114 29580
rect 1134 29534 1138 29580
rect 1158 29534 1162 29580
rect 1182 29534 1186 29580
rect 1206 29534 1210 29580
rect 1230 29534 1234 29580
rect 1254 29534 1258 29580
rect 1267 29573 1272 29580
rect 1277 29559 1282 29573
rect 1278 29534 1282 29559
rect 1302 29534 1306 29628
rect 1326 29534 1330 29628
rect 1350 29534 1354 29628
rect 1374 29534 1378 29628
rect 1398 29534 1402 29628
rect 1422 29534 1426 29628
rect 1446 29534 1450 29628
rect 1470 29534 1474 29628
rect 1494 29534 1498 29628
rect 1518 29534 1522 29628
rect 1542 29534 1546 29628
rect 1566 29534 1570 29628
rect 1590 29534 1594 29628
rect 1614 29534 1618 29628
rect 1638 29534 1642 29628
rect 1662 29534 1666 29628
rect 1686 29534 1690 29628
rect 1710 29534 1714 29628
rect 1734 29534 1738 29628
rect 1758 29534 1762 29628
rect 1782 29534 1786 29628
rect 1806 29534 1810 29628
rect 1830 29534 1834 29628
rect 1854 29534 1858 29628
rect 1878 29534 1882 29628
rect 1902 29534 1906 29628
rect 1926 29534 1930 29628
rect 1950 29534 1954 29628
rect 1974 29627 1978 29628
rect 1974 29606 1981 29627
rect 1987 29621 1992 29628
rect 1998 29621 2002 29628
rect 1997 29607 2002 29621
rect 1987 29606 2021 29607
rect 1957 29604 2021 29606
rect 1957 29603 1971 29604
rect 1974 29579 1981 29604
rect 1987 29597 1992 29604
rect 1997 29583 2002 29597
rect 1974 29534 1978 29579
rect 1998 29535 2002 29583
rect 1987 29534 2019 29535
rect -2393 29532 2019 29534
rect -2371 29486 -2366 29532
rect -2348 29486 -2343 29532
rect -2325 29486 -2320 29532
rect -2317 29528 -2309 29532
rect -2062 29528 -2054 29532
rect -2154 29524 -2138 29526
rect -2057 29524 -2054 29528
rect -2292 29518 -2054 29524
rect -2052 29518 -2044 29528
rect -2092 29502 -2062 29504
rect -2094 29498 -2062 29502
rect -2000 29486 -1992 29532
rect -1846 29525 -1806 29532
rect -1663 29528 -1655 29532
rect -1846 29518 -1680 29524
rect -1854 29502 -1806 29504
rect -1854 29498 -1680 29502
rect -1642 29486 -1637 29532
rect -1619 29486 -1614 29532
rect -1530 29486 -1526 29532
rect -1506 29486 -1502 29532
rect -1482 29486 -1478 29532
rect -1458 29486 -1454 29532
rect -1434 29486 -1430 29532
rect -1410 29486 -1406 29532
rect -1386 29486 -1382 29532
rect -1362 29486 -1358 29532
rect -1338 29486 -1334 29532
rect -1314 29486 -1310 29532
rect -1290 29486 -1286 29532
rect -1266 29486 -1262 29532
rect -1242 29486 -1238 29532
rect -1218 29486 -1214 29532
rect -1194 29486 -1190 29532
rect -1170 29486 -1166 29532
rect -1146 29486 -1142 29532
rect -1122 29486 -1118 29532
rect -1098 29486 -1094 29532
rect -1074 29486 -1070 29532
rect -1050 29486 -1046 29532
rect -1026 29486 -1022 29532
rect -1002 29486 -998 29532
rect -978 29486 -974 29532
rect -954 29486 -950 29532
rect -930 29486 -926 29532
rect -906 29486 -902 29532
rect -882 29486 -878 29532
rect -858 29486 -854 29532
rect -834 29486 -830 29532
rect -810 29486 -806 29532
rect -786 29486 -782 29532
rect -762 29486 -758 29532
rect -738 29486 -734 29532
rect -714 29486 -710 29532
rect -690 29486 -686 29532
rect -666 29486 -662 29532
rect -642 29486 -638 29532
rect -618 29486 -614 29532
rect -594 29486 -590 29532
rect -570 29486 -566 29532
rect -546 29486 -542 29532
rect -522 29486 -518 29532
rect -498 29486 -494 29532
rect -474 29486 -470 29532
rect -450 29486 -446 29532
rect -426 29486 -422 29532
rect -402 29486 -398 29532
rect -378 29486 -374 29532
rect -354 29486 -350 29532
rect -330 29486 -326 29532
rect -306 29486 -302 29532
rect -282 29486 -278 29532
rect -258 29486 -254 29532
rect -234 29486 -230 29532
rect -210 29486 -206 29532
rect -186 29486 -182 29532
rect -162 29486 -158 29532
rect -138 29486 -134 29532
rect -114 29486 -110 29532
rect -90 29486 -86 29532
rect -66 29486 -62 29532
rect -42 29486 -38 29532
rect -18 29486 -14 29532
rect 6 29486 10 29532
rect 30 29486 34 29532
rect 54 29486 58 29532
rect 78 29486 82 29532
rect 102 29486 106 29532
rect 126 29486 130 29532
rect 150 29486 154 29532
rect 174 29486 178 29532
rect 198 29486 202 29532
rect 222 29486 226 29532
rect 246 29486 250 29532
rect 270 29486 274 29532
rect 294 29486 298 29532
rect 318 29486 322 29532
rect 342 29486 346 29532
rect 366 29486 370 29532
rect 390 29486 394 29532
rect 414 29486 418 29532
rect 438 29486 442 29532
rect 462 29486 466 29532
rect 486 29486 490 29532
rect 510 29486 514 29532
rect 534 29486 538 29532
rect 558 29486 562 29532
rect 582 29486 586 29532
rect 606 29486 610 29532
rect 630 29486 634 29532
rect 654 29486 658 29532
rect 678 29486 682 29532
rect 702 29486 706 29532
rect 726 29486 730 29532
rect 750 29486 754 29532
rect 774 29486 778 29532
rect 798 29486 802 29532
rect 822 29486 826 29532
rect 846 29486 850 29532
rect 870 29486 874 29532
rect 894 29486 898 29532
rect 918 29486 922 29532
rect 942 29486 946 29532
rect 966 29486 970 29532
rect 990 29486 994 29532
rect 1014 29486 1018 29532
rect 1038 29486 1042 29532
rect 1062 29486 1066 29532
rect 1086 29486 1090 29532
rect 1110 29486 1114 29532
rect 1134 29486 1138 29532
rect 1158 29486 1162 29532
rect 1182 29486 1186 29532
rect 1206 29486 1210 29532
rect 1230 29486 1234 29532
rect 1254 29486 1258 29532
rect 1278 29486 1282 29532
rect 1302 29531 1306 29532
rect -2393 29484 1299 29486
rect -2371 29462 -2366 29484
rect -2348 29462 -2343 29484
rect -2325 29462 -2320 29484
rect -2072 29482 -2036 29483
rect -2072 29476 -2054 29482
rect -2309 29468 -2301 29476
rect -2317 29462 -2309 29468
rect -2092 29467 -2062 29472
rect -2000 29463 -1992 29484
rect -1938 29483 -1906 29484
rect -1920 29482 -1906 29483
rect -1806 29476 -1680 29482
rect -1854 29467 -1806 29472
rect -1655 29468 -1647 29476
rect -1982 29463 -1966 29464
rect -2000 29462 -1966 29463
rect -1846 29462 -1806 29465
rect -1663 29462 -1655 29468
rect -1642 29462 -1637 29484
rect -1619 29462 -1614 29484
rect -1530 29462 -1526 29484
rect -1506 29462 -1502 29484
rect -1482 29462 -1478 29484
rect -1458 29462 -1454 29484
rect -1434 29462 -1430 29484
rect -1410 29462 -1406 29484
rect -1386 29462 -1382 29484
rect -1362 29462 -1358 29484
rect -1338 29462 -1334 29484
rect -1314 29462 -1310 29484
rect -1290 29462 -1286 29484
rect -1266 29462 -1262 29484
rect -1242 29462 -1238 29484
rect -1218 29462 -1214 29484
rect -1194 29462 -1190 29484
rect -1170 29462 -1166 29484
rect -1146 29462 -1142 29484
rect -1122 29462 -1118 29484
rect -1098 29462 -1094 29484
rect -1074 29462 -1070 29484
rect -1050 29462 -1046 29484
rect -1026 29462 -1022 29484
rect -1002 29462 -998 29484
rect -978 29462 -974 29484
rect -954 29462 -950 29484
rect -930 29462 -926 29484
rect -906 29462 -902 29484
rect -882 29462 -878 29484
rect -858 29462 -854 29484
rect -834 29462 -830 29484
rect -810 29462 -806 29484
rect -786 29462 -782 29484
rect -762 29462 -758 29484
rect -738 29463 -734 29484
rect -749 29462 -715 29463
rect -2393 29460 -715 29462
rect -2371 29438 -2366 29460
rect -2348 29438 -2343 29460
rect -2325 29438 -2320 29460
rect -2000 29458 -1966 29460
rect -2309 29440 -2301 29448
rect -2062 29447 -2054 29454
rect -2092 29440 -2084 29447
rect -2062 29440 -2026 29442
rect -2317 29438 -2309 29440
rect -2062 29438 -2012 29440
rect -2000 29438 -1992 29458
rect -1982 29457 -1966 29458
rect -1846 29456 -1806 29460
rect -1846 29449 -1798 29454
rect -1806 29447 -1798 29449
rect -1854 29445 -1846 29447
rect -1854 29440 -1806 29445
rect -1655 29440 -1647 29448
rect -1864 29438 -1796 29439
rect -1663 29438 -1655 29440
rect -1642 29438 -1637 29460
rect -1619 29438 -1614 29460
rect -1530 29438 -1526 29460
rect -1506 29438 -1502 29460
rect -1482 29438 -1478 29460
rect -1458 29438 -1454 29460
rect -1434 29438 -1430 29460
rect -1410 29438 -1406 29460
rect -1386 29438 -1382 29460
rect -1362 29438 -1358 29460
rect -1338 29438 -1334 29460
rect -1314 29438 -1310 29460
rect -1290 29438 -1286 29460
rect -1266 29438 -1262 29460
rect -1242 29438 -1238 29460
rect -1218 29438 -1214 29460
rect -1194 29438 -1190 29460
rect -1170 29438 -1166 29460
rect -1146 29438 -1142 29460
rect -1122 29438 -1118 29460
rect -1098 29438 -1094 29460
rect -1074 29438 -1070 29460
rect -1050 29438 -1046 29460
rect -1026 29438 -1022 29460
rect -1002 29438 -998 29460
rect -978 29438 -974 29460
rect -954 29438 -950 29460
rect -930 29438 -926 29460
rect -906 29438 -902 29460
rect -882 29438 -878 29460
rect -858 29438 -854 29460
rect -834 29438 -830 29460
rect -810 29438 -806 29460
rect -786 29438 -782 29460
rect -762 29438 -758 29460
rect -749 29453 -744 29460
rect -738 29453 -734 29460
rect -739 29439 -734 29453
rect -738 29438 -734 29439
rect -714 29438 -710 29484
rect -690 29438 -686 29484
rect -666 29438 -662 29484
rect -642 29438 -638 29484
rect -618 29438 -614 29484
rect -594 29438 -590 29484
rect -570 29438 -566 29484
rect -546 29438 -542 29484
rect -522 29438 -518 29484
rect -498 29438 -494 29484
rect -474 29438 -470 29484
rect -450 29438 -446 29484
rect -426 29438 -422 29484
rect -402 29438 -398 29484
rect -378 29438 -374 29484
rect -354 29438 -350 29484
rect -330 29438 -326 29484
rect -306 29483 -302 29484
rect -306 29459 -299 29483
rect -306 29438 -302 29459
rect -282 29438 -278 29484
rect -258 29438 -254 29484
rect -234 29438 -230 29484
rect -210 29438 -206 29484
rect -186 29438 -182 29484
rect -162 29438 -158 29484
rect -138 29438 -134 29484
rect -114 29438 -110 29484
rect -90 29438 -86 29484
rect -66 29438 -62 29484
rect -42 29438 -38 29484
rect -18 29438 -14 29484
rect 6 29438 10 29484
rect 30 29438 34 29484
rect 54 29438 58 29484
rect 78 29438 82 29484
rect 102 29438 106 29484
rect 126 29438 130 29484
rect 150 29438 154 29484
rect 174 29438 178 29484
rect 198 29438 202 29484
rect 222 29438 226 29484
rect 246 29438 250 29484
rect 270 29438 274 29484
rect 294 29438 298 29484
rect 318 29438 322 29484
rect 342 29438 346 29484
rect 366 29438 370 29484
rect 390 29438 394 29484
rect 414 29438 418 29484
rect 438 29438 442 29484
rect 462 29438 466 29484
rect 486 29438 490 29484
rect 510 29438 514 29484
rect 534 29438 538 29484
rect 558 29438 562 29484
rect 582 29438 586 29484
rect 606 29438 610 29484
rect 630 29438 634 29484
rect 654 29438 658 29484
rect 678 29438 682 29484
rect 702 29438 706 29484
rect 726 29438 730 29484
rect 750 29438 754 29484
rect 774 29438 778 29484
rect 798 29438 802 29484
rect 822 29438 826 29484
rect 846 29438 850 29484
rect 870 29438 874 29484
rect 894 29438 898 29484
rect 918 29438 922 29484
rect 942 29438 946 29484
rect 966 29438 970 29484
rect 990 29438 994 29484
rect 1014 29438 1018 29484
rect 1038 29438 1042 29484
rect 1062 29438 1066 29484
rect 1086 29438 1090 29484
rect 1110 29438 1114 29484
rect 1134 29438 1138 29484
rect 1158 29438 1162 29484
rect 1182 29438 1186 29484
rect 1206 29438 1210 29484
rect 1230 29438 1234 29484
rect 1254 29438 1258 29484
rect 1278 29438 1282 29484
rect 1285 29483 1299 29484
rect 1302 29483 1309 29531
rect 1302 29438 1306 29483
rect 1326 29438 1330 29532
rect 1350 29438 1354 29532
rect 1374 29438 1378 29532
rect 1398 29438 1402 29532
rect 1422 29438 1426 29532
rect 1446 29438 1450 29532
rect 1470 29438 1474 29532
rect 1494 29438 1498 29532
rect 1518 29438 1522 29532
rect 1542 29438 1546 29532
rect 1566 29438 1570 29532
rect 1590 29438 1594 29532
rect 1614 29438 1618 29532
rect 1638 29438 1642 29532
rect 1662 29438 1666 29532
rect 1686 29438 1690 29532
rect 1710 29438 1714 29532
rect 1734 29511 1738 29532
rect 1723 29510 1757 29511
rect 1758 29510 1762 29532
rect 1782 29510 1786 29532
rect 1806 29510 1810 29532
rect 1830 29510 1834 29532
rect 1854 29510 1858 29532
rect 1878 29510 1882 29532
rect 1902 29510 1906 29532
rect 1926 29510 1930 29532
rect 1950 29510 1954 29532
rect 1974 29510 1978 29532
rect 1987 29525 1992 29532
rect 1998 29525 2002 29532
rect 2005 29531 2019 29532
rect 1997 29511 2002 29525
rect 2011 29521 2019 29525
rect 2005 29511 2011 29521
rect 1987 29510 2019 29511
rect 1723 29508 2019 29510
rect 1723 29501 1728 29508
rect 1734 29501 1738 29508
rect 1733 29487 1738 29501
rect 1723 29477 1728 29487
rect 1733 29463 1738 29477
rect 1734 29438 1738 29463
rect 1758 29438 1762 29508
rect 1782 29438 1786 29508
rect 1806 29438 1810 29508
rect 1830 29438 1834 29508
rect 1854 29438 1858 29508
rect 1878 29438 1882 29508
rect 1902 29438 1906 29508
rect 1926 29438 1930 29508
rect 1950 29438 1954 29508
rect 1974 29438 1978 29508
rect 1987 29501 1992 29508
rect 2005 29507 2019 29508
rect 1997 29487 2002 29501
rect 1998 29439 2002 29487
rect 1987 29438 2019 29439
rect -2393 29436 2019 29438
rect -2371 29390 -2366 29436
rect -2348 29390 -2343 29436
rect -2325 29390 -2320 29436
rect -2317 29432 -2309 29436
rect -2062 29432 -2054 29436
rect -2154 29428 -2138 29430
rect -2057 29428 -2054 29432
rect -2292 29422 -2054 29428
rect -2052 29422 -2044 29432
rect -2092 29406 -2062 29408
rect -2094 29402 -2062 29406
rect -2000 29390 -1992 29436
rect -1846 29429 -1806 29436
rect -1663 29432 -1655 29436
rect -1846 29422 -1680 29428
rect -1854 29406 -1806 29408
rect -1854 29402 -1680 29406
rect -1642 29390 -1637 29436
rect -1619 29390 -1614 29436
rect -1530 29390 -1526 29436
rect -1506 29390 -1502 29436
rect -1482 29390 -1478 29436
rect -1458 29390 -1454 29436
rect -1434 29390 -1430 29436
rect -1410 29390 -1406 29436
rect -1386 29390 -1382 29436
rect -1362 29390 -1358 29436
rect -1338 29390 -1334 29436
rect -1314 29390 -1310 29436
rect -1290 29390 -1286 29436
rect -1266 29390 -1262 29436
rect -1242 29390 -1238 29436
rect -1218 29390 -1214 29436
rect -1194 29390 -1190 29436
rect -1170 29390 -1166 29436
rect -1146 29390 -1142 29436
rect -1122 29390 -1118 29436
rect -1098 29390 -1094 29436
rect -1074 29390 -1070 29436
rect -1050 29390 -1046 29436
rect -1026 29390 -1022 29436
rect -1002 29390 -998 29436
rect -978 29390 -974 29436
rect -954 29390 -950 29436
rect -930 29390 -926 29436
rect -906 29390 -902 29436
rect -882 29390 -878 29436
rect -858 29390 -854 29436
rect -834 29390 -830 29436
rect -810 29390 -806 29436
rect -786 29390 -782 29436
rect -762 29390 -758 29436
rect -738 29390 -734 29436
rect -725 29405 -720 29415
rect -714 29405 -710 29436
rect -715 29391 -710 29405
rect -725 29390 -691 29391
rect -2393 29388 -691 29390
rect -2371 29366 -2366 29388
rect -2348 29366 -2343 29388
rect -2325 29366 -2320 29388
rect -2072 29386 -2036 29387
rect -2072 29380 -2054 29386
rect -2309 29372 -2301 29380
rect -2317 29366 -2309 29372
rect -2092 29371 -2062 29376
rect -2000 29367 -1992 29388
rect -1938 29387 -1906 29388
rect -1920 29386 -1906 29387
rect -1806 29380 -1680 29386
rect -1854 29371 -1806 29376
rect -1655 29372 -1647 29380
rect -1982 29367 -1966 29368
rect -2000 29366 -1966 29367
rect -1846 29366 -1806 29369
rect -1663 29366 -1655 29372
rect -1642 29366 -1637 29388
rect -1619 29366 -1614 29388
rect -1530 29366 -1526 29388
rect -1506 29366 -1502 29388
rect -1482 29366 -1478 29388
rect -1458 29366 -1454 29388
rect -1434 29366 -1430 29388
rect -1410 29366 -1406 29388
rect -1386 29366 -1382 29388
rect -1362 29366 -1358 29388
rect -1338 29366 -1334 29388
rect -1314 29366 -1310 29388
rect -1290 29366 -1286 29388
rect -1266 29366 -1262 29388
rect -1242 29366 -1238 29388
rect -1218 29366 -1214 29388
rect -1194 29366 -1190 29388
rect -1170 29366 -1166 29388
rect -1146 29366 -1142 29388
rect -1122 29366 -1118 29388
rect -1098 29366 -1094 29388
rect -1074 29366 -1070 29388
rect -1050 29366 -1046 29388
rect -1026 29366 -1022 29388
rect -1002 29366 -998 29388
rect -978 29366 -974 29388
rect -954 29366 -950 29388
rect -930 29367 -926 29388
rect -941 29366 -907 29367
rect -2393 29364 -907 29366
rect -2371 29342 -2366 29364
rect -2348 29342 -2343 29364
rect -2325 29342 -2320 29364
rect -2000 29362 -1966 29364
rect -2309 29344 -2301 29352
rect -2062 29351 -2054 29358
rect -2092 29344 -2084 29351
rect -2062 29344 -2026 29346
rect -2317 29342 -2309 29344
rect -2062 29342 -2012 29344
rect -2000 29342 -1992 29362
rect -1982 29361 -1966 29362
rect -1846 29360 -1806 29364
rect -1846 29353 -1798 29358
rect -1806 29351 -1798 29353
rect -1854 29349 -1846 29351
rect -1854 29344 -1806 29349
rect -1655 29344 -1647 29352
rect -1864 29342 -1796 29343
rect -1663 29342 -1655 29344
rect -1642 29342 -1637 29364
rect -1619 29342 -1614 29364
rect -1530 29342 -1526 29364
rect -1506 29342 -1502 29364
rect -1482 29342 -1478 29364
rect -1458 29342 -1454 29364
rect -1434 29342 -1430 29364
rect -1410 29342 -1406 29364
rect -1386 29342 -1382 29364
rect -1362 29342 -1358 29364
rect -1338 29342 -1334 29364
rect -1314 29342 -1310 29364
rect -1290 29342 -1286 29364
rect -1266 29342 -1262 29364
rect -1242 29342 -1238 29364
rect -1218 29342 -1214 29364
rect -1194 29342 -1190 29364
rect -1170 29342 -1166 29364
rect -1146 29342 -1142 29364
rect -1122 29342 -1118 29364
rect -1098 29342 -1094 29364
rect -1074 29342 -1070 29364
rect -1050 29342 -1046 29364
rect -1026 29342 -1022 29364
rect -1002 29342 -998 29364
rect -978 29342 -974 29364
rect -954 29342 -950 29364
rect -941 29357 -936 29364
rect -930 29357 -926 29364
rect -931 29343 -926 29357
rect -930 29342 -926 29343
rect -906 29342 -902 29388
rect -882 29342 -878 29388
rect -858 29342 -854 29388
rect -834 29342 -830 29388
rect -810 29342 -806 29388
rect -786 29342 -782 29388
rect -762 29342 -758 29388
rect -738 29342 -734 29388
rect -725 29381 -720 29388
rect -715 29367 -707 29381
rect -714 29363 -707 29367
rect -714 29342 -710 29363
rect -690 29342 -686 29436
rect -666 29342 -662 29436
rect -642 29342 -638 29436
rect -618 29342 -614 29436
rect -594 29342 -590 29436
rect -570 29342 -566 29436
rect -546 29342 -542 29436
rect -522 29342 -518 29436
rect -498 29342 -494 29436
rect -474 29342 -470 29436
rect -450 29342 -446 29436
rect -426 29342 -422 29436
rect -402 29342 -398 29436
rect -378 29342 -374 29436
rect -354 29342 -350 29436
rect -330 29342 -326 29436
rect -306 29342 -302 29436
rect -282 29342 -278 29436
rect -258 29342 -254 29436
rect -234 29342 -230 29436
rect -210 29342 -206 29436
rect -186 29342 -182 29436
rect -162 29342 -158 29436
rect -138 29342 -134 29436
rect -114 29342 -110 29436
rect -90 29342 -86 29436
rect -66 29343 -62 29436
rect -77 29342 -43 29343
rect -2393 29340 -43 29342
rect -2371 29294 -2366 29340
rect -2348 29294 -2343 29340
rect -2325 29294 -2320 29340
rect -2317 29336 -2309 29340
rect -2062 29336 -2054 29340
rect -2154 29332 -2138 29334
rect -2057 29332 -2054 29336
rect -2292 29326 -2054 29332
rect -2052 29326 -2044 29336
rect -2092 29310 -2062 29312
rect -2094 29306 -2062 29310
rect -2000 29294 -1992 29340
rect -1846 29333 -1806 29340
rect -1663 29336 -1655 29340
rect -1846 29326 -1680 29332
rect -1854 29310 -1806 29312
rect -1854 29306 -1680 29310
rect -1642 29294 -1637 29340
rect -1619 29294 -1614 29340
rect -1530 29294 -1526 29340
rect -1506 29294 -1502 29340
rect -1482 29294 -1478 29340
rect -1458 29294 -1454 29340
rect -1434 29294 -1430 29340
rect -1410 29294 -1406 29340
rect -1386 29294 -1382 29340
rect -1362 29294 -1358 29340
rect -1338 29294 -1334 29340
rect -1314 29294 -1310 29340
rect -1290 29294 -1286 29340
rect -1266 29294 -1262 29340
rect -1242 29294 -1238 29340
rect -1218 29294 -1214 29340
rect -1194 29294 -1190 29340
rect -1170 29294 -1166 29340
rect -1146 29294 -1142 29340
rect -1122 29294 -1118 29340
rect -1098 29294 -1094 29340
rect -1074 29294 -1070 29340
rect -1050 29294 -1046 29340
rect -1026 29294 -1022 29340
rect -1002 29294 -998 29340
rect -978 29294 -974 29340
rect -954 29294 -950 29340
rect -930 29294 -926 29340
rect -906 29294 -902 29340
rect -882 29294 -878 29340
rect -858 29294 -854 29340
rect -834 29294 -830 29340
rect -810 29294 -806 29340
rect -786 29294 -782 29340
rect -762 29294 -758 29340
rect -738 29294 -734 29340
rect -714 29294 -710 29340
rect -690 29339 -686 29340
rect -2393 29292 -693 29294
rect -2371 29270 -2366 29292
rect -2348 29270 -2343 29292
rect -2325 29270 -2320 29292
rect -2072 29290 -2036 29291
rect -2072 29284 -2054 29290
rect -2309 29276 -2301 29284
rect -2317 29270 -2309 29276
rect -2092 29275 -2062 29280
rect -2000 29271 -1992 29292
rect -1938 29291 -1906 29292
rect -1920 29290 -1906 29291
rect -1806 29284 -1680 29290
rect -1854 29275 -1806 29280
rect -1655 29276 -1647 29284
rect -1982 29271 -1966 29272
rect -2000 29270 -1966 29271
rect -1846 29270 -1806 29273
rect -1663 29270 -1655 29276
rect -1642 29270 -1637 29292
rect -1619 29270 -1614 29292
rect -1530 29270 -1526 29292
rect -1506 29270 -1502 29292
rect -1482 29270 -1478 29292
rect -1458 29270 -1454 29292
rect -1434 29270 -1430 29292
rect -1410 29270 -1406 29292
rect -1386 29270 -1382 29292
rect -1362 29270 -1358 29292
rect -1338 29270 -1334 29292
rect -1314 29270 -1310 29292
rect -1290 29270 -1286 29292
rect -1266 29270 -1262 29292
rect -1242 29270 -1238 29292
rect -1218 29270 -1214 29292
rect -1194 29270 -1190 29292
rect -1170 29270 -1166 29292
rect -1146 29270 -1142 29292
rect -1122 29270 -1118 29292
rect -1098 29270 -1094 29292
rect -1074 29270 -1070 29292
rect -1050 29270 -1046 29292
rect -1026 29270 -1022 29292
rect -1002 29270 -998 29292
rect -978 29270 -974 29292
rect -954 29270 -950 29292
rect -930 29270 -926 29292
rect -906 29291 -902 29292
rect -2393 29268 -909 29270
rect -2371 29246 -2366 29268
rect -2348 29246 -2343 29268
rect -2325 29246 -2320 29268
rect -2000 29266 -1966 29268
rect -2309 29248 -2301 29256
rect -2062 29255 -2054 29262
rect -2092 29248 -2084 29255
rect -2062 29248 -2026 29250
rect -2317 29246 -2309 29248
rect -2062 29246 -2012 29248
rect -2000 29246 -1992 29266
rect -1982 29265 -1966 29266
rect -1846 29264 -1806 29268
rect -1846 29257 -1798 29262
rect -1806 29255 -1798 29257
rect -1854 29253 -1846 29255
rect -1854 29248 -1806 29253
rect -1655 29248 -1647 29256
rect -1864 29246 -1796 29247
rect -1663 29246 -1655 29248
rect -1642 29246 -1637 29268
rect -1619 29246 -1614 29268
rect -1530 29246 -1526 29268
rect -1506 29246 -1502 29268
rect -1482 29246 -1478 29268
rect -1458 29246 -1454 29268
rect -1434 29246 -1430 29268
rect -1410 29246 -1406 29268
rect -1386 29246 -1382 29268
rect -1362 29246 -1358 29268
rect -1338 29246 -1334 29268
rect -1314 29246 -1310 29268
rect -1290 29246 -1286 29268
rect -1266 29246 -1262 29268
rect -1242 29246 -1238 29268
rect -1218 29246 -1214 29268
rect -1194 29246 -1190 29268
rect -1170 29246 -1166 29268
rect -1146 29246 -1142 29268
rect -1122 29246 -1118 29268
rect -1098 29246 -1094 29268
rect -1074 29246 -1070 29268
rect -1050 29246 -1046 29268
rect -1026 29246 -1022 29268
rect -1002 29246 -998 29268
rect -978 29246 -974 29268
rect -954 29246 -950 29268
rect -930 29246 -926 29268
rect -923 29267 -909 29268
rect -906 29267 -899 29291
rect -906 29246 -902 29267
rect -882 29246 -878 29292
rect -858 29246 -854 29292
rect -834 29246 -830 29292
rect -810 29246 -806 29292
rect -786 29246 -782 29292
rect -762 29246 -758 29292
rect -738 29246 -734 29292
rect -714 29246 -710 29292
rect -707 29291 -693 29292
rect -690 29291 -683 29339
rect -690 29246 -686 29291
rect -666 29246 -662 29340
rect -642 29246 -638 29340
rect -618 29246 -614 29340
rect -594 29246 -590 29340
rect -570 29246 -566 29340
rect -546 29246 -542 29340
rect -522 29247 -518 29340
rect -533 29246 -499 29247
rect -2393 29244 -499 29246
rect -2371 29198 -2366 29244
rect -2348 29198 -2343 29244
rect -2325 29198 -2320 29244
rect -2317 29240 -2309 29244
rect -2062 29240 -2054 29244
rect -2154 29236 -2138 29238
rect -2057 29236 -2054 29240
rect -2292 29230 -2054 29236
rect -2052 29230 -2044 29240
rect -2092 29214 -2062 29216
rect -2094 29210 -2062 29214
rect -2000 29198 -1992 29244
rect -1846 29237 -1806 29244
rect -1663 29240 -1655 29244
rect -1846 29230 -1680 29236
rect -1854 29214 -1806 29216
rect -1854 29210 -1680 29214
rect -1642 29198 -1637 29244
rect -1619 29198 -1614 29244
rect -1530 29198 -1526 29244
rect -1506 29198 -1502 29244
rect -1482 29198 -1478 29244
rect -1458 29198 -1454 29244
rect -1434 29198 -1430 29244
rect -1410 29198 -1406 29244
rect -1386 29198 -1382 29244
rect -1362 29198 -1358 29244
rect -1338 29198 -1334 29244
rect -1314 29198 -1310 29244
rect -1290 29198 -1286 29244
rect -1266 29198 -1262 29244
rect -1242 29198 -1238 29244
rect -1218 29198 -1214 29244
rect -1194 29198 -1190 29244
rect -1170 29198 -1166 29244
rect -1146 29198 -1142 29244
rect -1122 29198 -1118 29244
rect -1098 29198 -1094 29244
rect -1074 29198 -1070 29244
rect -1050 29198 -1046 29244
rect -1026 29198 -1022 29244
rect -1002 29198 -998 29244
rect -978 29198 -974 29244
rect -954 29198 -950 29244
rect -930 29198 -926 29244
rect -906 29198 -902 29244
rect -882 29198 -878 29244
rect -858 29198 -854 29244
rect -834 29198 -830 29244
rect -810 29198 -806 29244
rect -786 29198 -782 29244
rect -762 29198 -758 29244
rect -738 29198 -734 29244
rect -714 29198 -710 29244
rect -690 29198 -686 29244
rect -666 29198 -662 29244
rect -642 29198 -638 29244
rect -618 29198 -614 29244
rect -594 29198 -590 29244
rect -570 29198 -566 29244
rect -546 29198 -542 29244
rect -533 29237 -528 29244
rect -522 29237 -518 29244
rect -523 29223 -518 29237
rect -522 29198 -518 29223
rect -498 29198 -494 29340
rect -474 29198 -470 29340
rect -450 29198 -446 29340
rect -426 29198 -422 29340
rect -402 29198 -398 29340
rect -378 29198 -374 29340
rect -354 29198 -350 29340
rect -330 29198 -326 29340
rect -306 29198 -302 29340
rect -282 29198 -278 29340
rect -258 29198 -254 29340
rect -234 29198 -230 29340
rect -210 29198 -206 29340
rect -186 29198 -182 29340
rect -162 29198 -158 29340
rect -138 29198 -134 29340
rect -114 29198 -110 29340
rect -90 29198 -86 29340
rect -77 29333 -72 29340
rect -66 29333 -62 29340
rect -67 29319 -62 29333
rect -77 29261 -72 29271
rect -66 29261 -62 29319
rect -42 29267 -38 29436
rect -67 29247 -62 29261
rect -53 29257 -45 29261
rect -59 29247 -53 29257
rect -66 29198 -62 29247
rect -42 29243 -35 29267
rect -42 29198 -38 29243
rect -18 29198 -14 29436
rect 6 29198 10 29436
rect 30 29198 34 29436
rect 54 29198 58 29436
rect 78 29198 82 29436
rect 102 29198 106 29436
rect 126 29198 130 29436
rect 150 29198 154 29436
rect 174 29198 178 29436
rect 198 29198 202 29436
rect 222 29198 226 29436
rect 246 29198 250 29436
rect 270 29198 274 29436
rect 294 29198 298 29436
rect 318 29198 322 29436
rect 342 29198 346 29436
rect 366 29198 370 29436
rect 390 29198 394 29436
rect 414 29198 418 29436
rect 438 29198 442 29436
rect 462 29198 466 29436
rect 486 29198 490 29436
rect 510 29198 514 29436
rect 534 29198 538 29436
rect 558 29198 562 29436
rect 582 29198 586 29436
rect 606 29198 610 29436
rect 630 29198 634 29436
rect 654 29198 658 29436
rect 678 29198 682 29436
rect 702 29319 706 29436
rect 691 29318 725 29319
rect 726 29318 730 29436
rect 750 29318 754 29436
rect 774 29318 778 29436
rect 798 29318 802 29436
rect 822 29318 826 29436
rect 846 29318 850 29436
rect 870 29318 874 29436
rect 894 29318 898 29436
rect 918 29318 922 29436
rect 942 29318 946 29436
rect 966 29318 970 29436
rect 990 29318 994 29436
rect 1014 29318 1018 29436
rect 1038 29318 1042 29436
rect 1062 29318 1066 29436
rect 1086 29318 1090 29436
rect 1110 29318 1114 29436
rect 1134 29318 1138 29436
rect 1158 29318 1162 29436
rect 1182 29318 1186 29436
rect 1206 29318 1210 29436
rect 1230 29318 1234 29436
rect 1254 29318 1258 29436
rect 1278 29318 1282 29436
rect 1302 29318 1306 29436
rect 1326 29318 1330 29436
rect 1350 29318 1354 29436
rect 1374 29318 1378 29436
rect 1398 29318 1402 29436
rect 1422 29318 1426 29436
rect 1446 29318 1450 29436
rect 1470 29318 1474 29436
rect 1494 29318 1498 29436
rect 1518 29318 1522 29436
rect 1542 29318 1546 29436
rect 1566 29318 1570 29436
rect 1590 29318 1594 29436
rect 1614 29318 1618 29436
rect 1638 29318 1642 29436
rect 1662 29318 1666 29436
rect 1686 29318 1690 29436
rect 1710 29318 1714 29436
rect 1734 29318 1738 29436
rect 1758 29435 1762 29436
rect 1758 29414 1765 29435
rect 1782 29414 1786 29436
rect 1806 29414 1810 29436
rect 1830 29414 1834 29436
rect 1854 29414 1858 29436
rect 1878 29414 1882 29436
rect 1902 29414 1906 29436
rect 1926 29414 1930 29436
rect 1950 29414 1954 29436
rect 1974 29414 1978 29436
rect 1987 29429 1992 29436
rect 1998 29429 2002 29436
rect 2005 29435 2019 29436
rect 1997 29415 2002 29429
rect 2011 29425 2019 29429
rect 2005 29415 2011 29425
rect 1987 29414 2019 29415
rect 1741 29412 2019 29414
rect 1741 29411 1755 29412
rect 1758 29387 1765 29412
rect 1758 29318 1762 29387
rect 1782 29318 1786 29412
rect 1806 29318 1810 29412
rect 1830 29318 1834 29412
rect 1854 29318 1858 29412
rect 1878 29318 1882 29412
rect 1902 29318 1906 29412
rect 1926 29318 1930 29412
rect 1950 29318 1954 29412
rect 1974 29318 1978 29412
rect 1987 29405 1992 29412
rect 2005 29411 2019 29412
rect 1997 29391 2002 29405
rect 1998 29318 2002 29391
rect 2011 29318 2019 29319
rect 691 29316 2019 29318
rect 691 29309 696 29316
rect 702 29309 706 29316
rect 701 29295 706 29309
rect 691 29285 696 29295
rect 701 29271 706 29285
rect 702 29198 706 29271
rect 726 29243 730 29316
rect -2393 29196 723 29198
rect -2371 29174 -2366 29196
rect -2348 29174 -2343 29196
rect -2325 29174 -2320 29196
rect -2072 29194 -2036 29195
rect -2072 29188 -2054 29194
rect -2309 29180 -2301 29188
rect -2317 29174 -2309 29180
rect -2092 29179 -2062 29184
rect -2000 29175 -1992 29196
rect -1938 29195 -1906 29196
rect -1920 29194 -1906 29195
rect -1806 29188 -1680 29194
rect -1854 29179 -1806 29184
rect -1655 29180 -1647 29188
rect -1982 29175 -1966 29176
rect -2000 29174 -1966 29175
rect -1846 29174 -1806 29177
rect -1663 29174 -1655 29180
rect -1642 29174 -1637 29196
rect -1619 29174 -1614 29196
rect -1530 29174 -1526 29196
rect -1506 29174 -1502 29196
rect -1482 29174 -1478 29196
rect -1458 29174 -1454 29196
rect -1434 29174 -1430 29196
rect -1410 29174 -1406 29196
rect -1386 29174 -1382 29196
rect -1362 29174 -1358 29196
rect -1338 29174 -1334 29196
rect -1314 29174 -1310 29196
rect -1290 29174 -1286 29196
rect -1266 29174 -1262 29196
rect -1242 29174 -1238 29196
rect -1218 29174 -1214 29196
rect -1194 29174 -1190 29196
rect -1170 29174 -1166 29196
rect -1146 29174 -1142 29196
rect -1122 29174 -1118 29196
rect -1098 29174 -1094 29196
rect -1074 29174 -1070 29196
rect -1050 29174 -1046 29196
rect -1026 29174 -1022 29196
rect -1002 29174 -998 29196
rect -978 29174 -974 29196
rect -954 29174 -950 29196
rect -930 29174 -926 29196
rect -906 29174 -902 29196
rect -882 29174 -878 29196
rect -858 29174 -854 29196
rect -834 29174 -830 29196
rect -810 29174 -806 29196
rect -786 29174 -782 29196
rect -762 29174 -758 29196
rect -738 29174 -734 29196
rect -714 29174 -710 29196
rect -690 29174 -686 29196
rect -666 29174 -662 29196
rect -642 29174 -638 29196
rect -618 29174 -614 29196
rect -594 29174 -590 29196
rect -570 29174 -566 29196
rect -546 29174 -542 29196
rect -522 29174 -518 29196
rect -498 29174 -494 29196
rect -474 29174 -470 29196
rect -450 29174 -446 29196
rect -426 29174 -422 29196
rect -402 29174 -398 29196
rect -378 29174 -374 29196
rect -354 29174 -350 29196
rect -330 29174 -326 29196
rect -306 29174 -302 29196
rect -282 29174 -278 29196
rect -258 29174 -254 29196
rect -234 29174 -230 29196
rect -210 29174 -206 29196
rect -186 29174 -182 29196
rect -162 29174 -158 29196
rect -138 29174 -134 29196
rect -114 29174 -110 29196
rect -90 29174 -86 29196
rect -66 29174 -62 29196
rect -42 29195 -38 29196
rect -2393 29172 -45 29174
rect -2371 29150 -2366 29172
rect -2348 29150 -2343 29172
rect -2325 29150 -2320 29172
rect -2000 29170 -1966 29172
rect -2309 29152 -2301 29160
rect -2062 29159 -2054 29166
rect -2092 29152 -2084 29159
rect -2062 29152 -2026 29154
rect -2317 29150 -2309 29152
rect -2062 29150 -2012 29152
rect -2000 29150 -1992 29170
rect -1982 29169 -1966 29170
rect -1846 29168 -1806 29172
rect -1846 29161 -1798 29166
rect -1806 29159 -1798 29161
rect -1854 29157 -1846 29159
rect -1854 29152 -1806 29157
rect -1655 29152 -1647 29160
rect -1864 29150 -1796 29151
rect -1663 29150 -1655 29152
rect -1642 29150 -1637 29172
rect -1619 29150 -1614 29172
rect -1530 29150 -1526 29172
rect -1506 29150 -1502 29172
rect -1482 29150 -1478 29172
rect -1458 29150 -1454 29172
rect -1434 29150 -1430 29172
rect -1410 29150 -1406 29172
rect -1386 29150 -1382 29172
rect -1362 29150 -1358 29172
rect -1338 29150 -1334 29172
rect -1314 29150 -1310 29172
rect -1290 29150 -1286 29172
rect -1266 29150 -1262 29172
rect -1242 29150 -1238 29172
rect -1218 29150 -1214 29172
rect -1194 29150 -1190 29172
rect -1170 29150 -1166 29172
rect -1146 29150 -1142 29172
rect -1122 29150 -1118 29172
rect -1098 29150 -1094 29172
rect -1074 29150 -1070 29172
rect -1050 29150 -1046 29172
rect -1026 29150 -1022 29172
rect -1002 29150 -998 29172
rect -978 29150 -974 29172
rect -954 29150 -950 29172
rect -930 29150 -926 29172
rect -906 29150 -902 29172
rect -882 29150 -878 29172
rect -858 29150 -854 29172
rect -834 29150 -830 29172
rect -810 29150 -806 29172
rect -786 29150 -782 29172
rect -762 29150 -758 29172
rect -738 29150 -734 29172
rect -714 29150 -710 29172
rect -690 29150 -686 29172
rect -666 29150 -662 29172
rect -642 29150 -638 29172
rect -618 29150 -614 29172
rect -594 29150 -590 29172
rect -570 29150 -566 29172
rect -546 29150 -542 29172
rect -522 29150 -518 29172
rect -498 29171 -494 29172
rect -2393 29148 -501 29150
rect -2371 29102 -2366 29148
rect -2348 29102 -2343 29148
rect -2325 29102 -2320 29148
rect -2317 29144 -2309 29148
rect -2062 29144 -2054 29148
rect -2154 29140 -2138 29142
rect -2057 29140 -2054 29144
rect -2292 29134 -2054 29140
rect -2052 29134 -2044 29144
rect -2092 29118 -2062 29120
rect -2094 29114 -2062 29118
rect -2000 29102 -1992 29148
rect -1846 29141 -1806 29148
rect -1663 29144 -1655 29148
rect -1846 29134 -1680 29140
rect -1854 29118 -1806 29120
rect -1854 29114 -1680 29118
rect -1642 29102 -1637 29148
rect -1619 29102 -1614 29148
rect -1530 29102 -1526 29148
rect -1506 29102 -1502 29148
rect -1482 29102 -1478 29148
rect -1458 29102 -1454 29148
rect -1434 29102 -1430 29148
rect -1410 29102 -1406 29148
rect -1386 29102 -1382 29148
rect -1362 29102 -1358 29148
rect -1338 29102 -1334 29148
rect -1314 29102 -1310 29148
rect -1290 29102 -1286 29148
rect -1266 29102 -1262 29148
rect -1242 29102 -1238 29148
rect -1218 29102 -1214 29148
rect -1194 29102 -1190 29148
rect -1170 29102 -1166 29148
rect -1146 29102 -1142 29148
rect -1122 29102 -1118 29148
rect -1098 29102 -1094 29148
rect -1074 29102 -1070 29148
rect -1050 29102 -1046 29148
rect -1026 29102 -1022 29148
rect -1002 29102 -998 29148
rect -978 29102 -974 29148
rect -954 29102 -950 29148
rect -930 29102 -926 29148
rect -906 29102 -902 29148
rect -882 29102 -878 29148
rect -858 29102 -854 29148
rect -834 29102 -830 29148
rect -810 29102 -806 29148
rect -786 29102 -782 29148
rect -762 29102 -758 29148
rect -738 29102 -734 29148
rect -714 29102 -710 29148
rect -690 29102 -686 29148
rect -666 29102 -662 29148
rect -642 29102 -638 29148
rect -618 29102 -614 29148
rect -594 29102 -590 29148
rect -570 29102 -566 29148
rect -546 29102 -542 29148
rect -522 29102 -518 29148
rect -515 29147 -501 29148
rect -498 29147 -491 29171
rect -498 29102 -494 29147
rect -474 29102 -470 29172
rect -450 29102 -446 29172
rect -426 29102 -422 29172
rect -402 29102 -398 29172
rect -378 29102 -374 29172
rect -354 29102 -350 29172
rect -330 29102 -326 29172
rect -306 29102 -302 29172
rect -282 29102 -278 29172
rect -258 29102 -254 29172
rect -234 29102 -230 29172
rect -210 29102 -206 29172
rect -186 29102 -182 29172
rect -162 29102 -158 29172
rect -138 29102 -134 29172
rect -114 29102 -110 29172
rect -90 29102 -86 29172
rect -66 29102 -62 29172
rect -59 29171 -45 29172
rect -42 29171 -35 29195
rect -42 29102 -38 29171
rect -18 29102 -14 29196
rect 6 29102 10 29196
rect 30 29102 34 29196
rect 54 29102 58 29196
rect 78 29102 82 29196
rect 102 29102 106 29196
rect 126 29102 130 29196
rect 150 29102 154 29196
rect 174 29102 178 29196
rect 198 29102 202 29196
rect 222 29102 226 29196
rect 246 29102 250 29196
rect 270 29102 274 29196
rect 294 29102 298 29196
rect 318 29102 322 29196
rect 342 29102 346 29196
rect 366 29102 370 29196
rect 390 29102 394 29196
rect 414 29102 418 29196
rect 438 29102 442 29196
rect 462 29102 466 29196
rect 486 29102 490 29196
rect 499 29117 504 29127
rect 510 29117 514 29196
rect 509 29103 514 29117
rect 499 29102 533 29103
rect -2393 29100 533 29102
rect -2371 29078 -2366 29100
rect -2348 29078 -2343 29100
rect -2325 29078 -2320 29100
rect -2072 29098 -2036 29099
rect -2072 29092 -2054 29098
rect -2309 29084 -2301 29092
rect -2317 29078 -2309 29084
rect -2092 29083 -2062 29088
rect -2000 29079 -1992 29100
rect -1938 29099 -1906 29100
rect -1920 29098 -1906 29099
rect -1806 29092 -1680 29098
rect -1854 29083 -1806 29088
rect -1655 29084 -1647 29092
rect -1982 29079 -1966 29080
rect -2000 29078 -1966 29079
rect -1846 29078 -1806 29081
rect -1663 29078 -1655 29084
rect -1642 29078 -1637 29100
rect -1619 29078 -1614 29100
rect -1530 29078 -1526 29100
rect -1506 29078 -1502 29100
rect -1482 29078 -1478 29100
rect -1458 29078 -1454 29100
rect -1434 29078 -1430 29100
rect -1410 29078 -1406 29100
rect -1386 29078 -1382 29100
rect -1362 29078 -1358 29100
rect -1338 29078 -1334 29100
rect -1314 29078 -1310 29100
rect -1290 29078 -1286 29100
rect -1266 29078 -1262 29100
rect -1242 29078 -1238 29100
rect -1218 29078 -1214 29100
rect -1194 29078 -1190 29100
rect -1170 29078 -1166 29100
rect -1146 29078 -1142 29100
rect -1122 29078 -1118 29100
rect -1098 29078 -1094 29100
rect -1074 29078 -1070 29100
rect -1050 29078 -1046 29100
rect -1026 29078 -1022 29100
rect -1002 29078 -998 29100
rect -978 29078 -974 29100
rect -954 29078 -950 29100
rect -930 29078 -926 29100
rect -906 29078 -902 29100
rect -882 29078 -878 29100
rect -858 29078 -854 29100
rect -834 29078 -830 29100
rect -810 29078 -806 29100
rect -786 29078 -782 29100
rect -762 29078 -758 29100
rect -738 29078 -734 29100
rect -714 29078 -710 29100
rect -690 29078 -686 29100
rect -666 29078 -662 29100
rect -642 29078 -638 29100
rect -618 29078 -614 29100
rect -594 29078 -590 29100
rect -570 29078 -566 29100
rect -546 29078 -542 29100
rect -522 29078 -518 29100
rect -498 29078 -494 29100
rect -474 29078 -470 29100
rect -450 29078 -446 29100
rect -426 29078 -422 29100
rect -402 29078 -398 29100
rect -378 29078 -374 29100
rect -354 29078 -350 29100
rect -330 29078 -326 29100
rect -306 29078 -302 29100
rect -282 29078 -278 29100
rect -258 29078 -254 29100
rect -234 29078 -230 29100
rect -210 29078 -206 29100
rect -186 29078 -182 29100
rect -162 29078 -158 29100
rect -138 29078 -134 29100
rect -114 29078 -110 29100
rect -90 29078 -86 29100
rect -66 29078 -62 29100
rect -42 29078 -38 29100
rect -18 29078 -14 29100
rect 6 29078 10 29100
rect 30 29078 34 29100
rect 54 29078 58 29100
rect 78 29078 82 29100
rect 102 29078 106 29100
rect 126 29078 130 29100
rect 150 29078 154 29100
rect 174 29078 178 29100
rect 198 29078 202 29100
rect 222 29078 226 29100
rect 246 29078 250 29100
rect 270 29078 274 29100
rect 294 29078 298 29100
rect 318 29078 322 29100
rect 342 29078 346 29100
rect 366 29078 370 29100
rect 390 29078 394 29100
rect 414 29078 418 29100
rect 438 29078 442 29100
rect 462 29078 466 29100
rect 486 29078 490 29100
rect 499 29093 504 29100
rect 509 29079 514 29093
rect 510 29078 514 29079
rect 534 29078 538 29196
rect 558 29078 562 29196
rect 582 29078 586 29196
rect 606 29078 610 29196
rect 630 29078 634 29196
rect 654 29078 658 29196
rect 678 29078 682 29196
rect 702 29078 706 29196
rect 709 29195 723 29196
rect 726 29195 733 29243
rect 726 29078 730 29195
rect 750 29078 754 29316
rect 774 29078 778 29316
rect 798 29078 802 29316
rect 822 29078 826 29316
rect 846 29078 850 29316
rect 870 29078 874 29316
rect 894 29078 898 29316
rect 918 29078 922 29316
rect 942 29078 946 29316
rect 966 29079 970 29316
rect 955 29078 989 29079
rect -2393 29076 989 29078
rect -2371 29054 -2366 29076
rect -2348 29054 -2343 29076
rect -2325 29054 -2320 29076
rect -2000 29074 -1966 29076
rect -2309 29056 -2301 29064
rect -2062 29063 -2054 29070
rect -2092 29056 -2084 29063
rect -2062 29056 -2026 29058
rect -2317 29054 -2309 29056
rect -2062 29054 -2012 29056
rect -2000 29054 -1992 29074
rect -1982 29073 -1966 29074
rect -1846 29072 -1806 29076
rect -1846 29065 -1798 29070
rect -1806 29063 -1798 29065
rect -1854 29061 -1846 29063
rect -1854 29056 -1806 29061
rect -1655 29056 -1647 29064
rect -1864 29054 -1796 29055
rect -1663 29054 -1655 29056
rect -1642 29054 -1637 29076
rect -1619 29054 -1614 29076
rect -1530 29054 -1526 29076
rect -1506 29054 -1502 29076
rect -1482 29054 -1478 29076
rect -1458 29054 -1454 29076
rect -1434 29054 -1430 29076
rect -1410 29054 -1406 29076
rect -1386 29054 -1382 29076
rect -1362 29054 -1358 29076
rect -1338 29054 -1334 29076
rect -1314 29054 -1310 29076
rect -1290 29054 -1286 29076
rect -1266 29054 -1262 29076
rect -1242 29054 -1238 29076
rect -1218 29054 -1214 29076
rect -1194 29054 -1190 29076
rect -1170 29054 -1166 29076
rect -1146 29054 -1142 29076
rect -1122 29054 -1118 29076
rect -1098 29054 -1094 29076
rect -1074 29054 -1070 29076
rect -1050 29054 -1046 29076
rect -1026 29054 -1022 29076
rect -1002 29054 -998 29076
rect -978 29054 -974 29076
rect -954 29054 -950 29076
rect -930 29054 -926 29076
rect -906 29054 -902 29076
rect -882 29054 -878 29076
rect -858 29054 -854 29076
rect -834 29054 -830 29076
rect -810 29054 -806 29076
rect -786 29054 -782 29076
rect -762 29054 -758 29076
rect -738 29054 -734 29076
rect -714 29054 -710 29076
rect -690 29054 -686 29076
rect -666 29054 -662 29076
rect -642 29054 -638 29076
rect -618 29054 -614 29076
rect -594 29054 -590 29076
rect -570 29054 -566 29076
rect -546 29054 -542 29076
rect -522 29054 -518 29076
rect -498 29054 -494 29076
rect -474 29054 -470 29076
rect -450 29054 -446 29076
rect -426 29054 -422 29076
rect -402 29054 -398 29076
rect -378 29054 -374 29076
rect -354 29054 -350 29076
rect -330 29054 -326 29076
rect -306 29054 -302 29076
rect -282 29054 -278 29076
rect -258 29054 -254 29076
rect -234 29054 -230 29076
rect -210 29054 -206 29076
rect -186 29054 -182 29076
rect -162 29054 -158 29076
rect -138 29054 -134 29076
rect -114 29054 -110 29076
rect -90 29054 -86 29076
rect -66 29054 -62 29076
rect -42 29054 -38 29076
rect -18 29054 -14 29076
rect 6 29054 10 29076
rect 30 29054 34 29076
rect 54 29054 58 29076
rect 78 29054 82 29076
rect 102 29054 106 29076
rect 126 29054 130 29076
rect 150 29054 154 29076
rect 174 29054 178 29076
rect 198 29054 202 29076
rect 222 29054 226 29076
rect 246 29054 250 29076
rect 270 29054 274 29076
rect 294 29054 298 29076
rect 318 29054 322 29076
rect 342 29054 346 29076
rect 366 29054 370 29076
rect 390 29054 394 29076
rect 414 29054 418 29076
rect 438 29054 442 29076
rect 462 29054 466 29076
rect 486 29054 490 29076
rect 510 29054 514 29076
rect 534 29054 538 29076
rect 558 29054 562 29076
rect 582 29054 586 29076
rect 606 29054 610 29076
rect 630 29054 634 29076
rect 654 29054 658 29076
rect 678 29054 682 29076
rect 702 29054 706 29076
rect 726 29054 730 29076
rect 750 29054 754 29076
rect 774 29054 778 29076
rect 798 29054 802 29076
rect 822 29054 826 29076
rect 846 29054 850 29076
rect 870 29054 874 29076
rect 894 29054 898 29076
rect 918 29054 922 29076
rect 942 29054 946 29076
rect 955 29069 960 29076
rect 966 29069 970 29076
rect 965 29055 970 29069
rect 966 29054 970 29055
rect 990 29054 994 29316
rect 1014 29054 1018 29316
rect 1038 29054 1042 29316
rect 1051 29165 1056 29175
rect 1062 29165 1066 29316
rect 1061 29151 1066 29165
rect 1062 29054 1066 29151
rect 1086 29099 1090 29316
rect 1086 29075 1093 29099
rect 1086 29054 1090 29075
rect 1110 29054 1114 29316
rect 1134 29054 1138 29316
rect 1158 29054 1162 29316
rect 1182 29054 1186 29316
rect 1206 29054 1210 29316
rect 1230 29223 1234 29316
rect 1219 29222 1253 29223
rect 1254 29222 1258 29316
rect 1278 29222 1282 29316
rect 1302 29222 1306 29316
rect 1326 29222 1330 29316
rect 1350 29222 1354 29316
rect 1374 29222 1378 29316
rect 1398 29222 1402 29316
rect 1422 29222 1426 29316
rect 1446 29222 1450 29316
rect 1470 29222 1474 29316
rect 1494 29222 1498 29316
rect 1518 29222 1522 29316
rect 1542 29222 1546 29316
rect 1566 29222 1570 29316
rect 1590 29222 1594 29316
rect 1614 29222 1618 29316
rect 1638 29222 1642 29316
rect 1662 29222 1666 29316
rect 1686 29222 1690 29316
rect 1710 29222 1714 29316
rect 1734 29222 1738 29316
rect 1758 29222 1762 29316
rect 1782 29222 1786 29316
rect 1806 29222 1810 29316
rect 1830 29222 1834 29316
rect 1854 29222 1858 29316
rect 1878 29222 1882 29316
rect 1902 29222 1906 29316
rect 1926 29222 1930 29316
rect 1950 29222 1954 29316
rect 1974 29222 1978 29316
rect 1998 29222 2002 29316
rect 2005 29315 2019 29316
rect 2011 29309 2016 29315
rect 2021 29295 2026 29309
rect 2022 29222 2026 29295
rect 2035 29222 2043 29223
rect 1219 29220 2043 29222
rect 1219 29213 1224 29220
rect 1230 29213 1234 29220
rect 1229 29199 1234 29213
rect 1219 29189 1224 29199
rect 1229 29175 1234 29189
rect 1230 29054 1234 29175
rect 1254 29147 1258 29220
rect 1254 29126 1261 29147
rect 1278 29126 1282 29220
rect 1302 29126 1306 29220
rect 1326 29126 1330 29220
rect 1350 29126 1354 29220
rect 1374 29126 1378 29220
rect 1398 29126 1402 29220
rect 1422 29126 1426 29220
rect 1446 29126 1450 29220
rect 1470 29126 1474 29220
rect 1494 29126 1498 29220
rect 1518 29126 1522 29220
rect 1542 29126 1546 29220
rect 1566 29126 1570 29220
rect 1590 29126 1594 29220
rect 1614 29126 1618 29220
rect 1638 29126 1642 29220
rect 1662 29126 1666 29220
rect 1686 29126 1690 29220
rect 1710 29126 1714 29220
rect 1734 29126 1738 29220
rect 1758 29126 1762 29220
rect 1782 29126 1786 29220
rect 1806 29126 1810 29220
rect 1830 29126 1834 29220
rect 1854 29126 1858 29220
rect 1878 29126 1882 29220
rect 1902 29126 1906 29220
rect 1926 29126 1930 29220
rect 1950 29126 1954 29220
rect 1974 29126 1978 29220
rect 1998 29126 2002 29220
rect 2022 29126 2026 29220
rect 2029 29219 2043 29220
rect 2035 29213 2040 29219
rect 2045 29199 2050 29213
rect 2035 29141 2040 29151
rect 2046 29141 2050 29199
rect 2045 29127 2050 29141
rect 2059 29137 2067 29141
rect 2053 29127 2059 29137
rect 2035 29126 2067 29127
rect 1237 29124 2067 29126
rect 1237 29123 1251 29124
rect 1254 29099 1261 29124
rect 1254 29054 1258 29099
rect 1278 29054 1282 29124
rect 1302 29054 1306 29124
rect 1326 29054 1330 29124
rect 1350 29054 1354 29124
rect 1374 29054 1378 29124
rect 1398 29054 1402 29124
rect 1422 29054 1426 29124
rect 1446 29054 1450 29124
rect 1470 29054 1474 29124
rect 1494 29054 1498 29124
rect 1518 29054 1522 29124
rect 1542 29054 1546 29124
rect 1566 29054 1570 29124
rect 1590 29054 1594 29124
rect 1614 29054 1618 29124
rect 1638 29054 1642 29124
rect 1662 29054 1666 29124
rect 1686 29054 1690 29124
rect 1710 29054 1714 29124
rect 1734 29054 1738 29124
rect 1758 29054 1762 29124
rect 1782 29054 1786 29124
rect 1806 29054 1810 29124
rect 1830 29054 1834 29124
rect 1854 29054 1858 29124
rect 1878 29054 1882 29124
rect 1902 29054 1906 29124
rect 1926 29054 1930 29124
rect 1950 29054 1954 29124
rect 1974 29054 1978 29124
rect 1998 29054 2002 29124
rect 2022 29054 2026 29124
rect 2035 29117 2040 29124
rect 2053 29123 2067 29124
rect 2045 29103 2050 29117
rect 2046 29055 2050 29103
rect 2035 29054 2067 29055
rect -2393 29052 2067 29054
rect -2371 29006 -2366 29052
rect -2348 29006 -2343 29052
rect -2325 29006 -2320 29052
rect -2317 29048 -2309 29052
rect -2062 29048 -2054 29052
rect -2154 29044 -2138 29046
rect -2057 29044 -2054 29048
rect -2292 29038 -2054 29044
rect -2052 29038 -2044 29048
rect -2092 29022 -2062 29024
rect -2094 29018 -2062 29022
rect -2000 29006 -1992 29052
rect -1846 29045 -1806 29052
rect -1663 29048 -1655 29052
rect -1846 29038 -1680 29044
rect -1854 29022 -1806 29024
rect -1854 29018 -1680 29022
rect -1642 29006 -1637 29052
rect -1619 29006 -1614 29052
rect -1530 29006 -1526 29052
rect -1506 29006 -1502 29052
rect -1482 29006 -1478 29052
rect -1458 29006 -1454 29052
rect -1434 29006 -1430 29052
rect -1410 29006 -1406 29052
rect -1386 29006 -1382 29052
rect -1362 29006 -1358 29052
rect -1338 29006 -1334 29052
rect -1314 29006 -1310 29052
rect -1290 29006 -1286 29052
rect -1266 29006 -1262 29052
rect -1242 29006 -1238 29052
rect -1218 29006 -1214 29052
rect -1194 29006 -1190 29052
rect -1170 29006 -1166 29052
rect -1146 29006 -1142 29052
rect -1122 29006 -1118 29052
rect -1109 29021 -1104 29031
rect -1098 29021 -1094 29052
rect -1099 29007 -1094 29021
rect -1109 29006 -1075 29007
rect -2393 29004 -1075 29006
rect -2371 28958 -2366 29004
rect -2348 28958 -2343 29004
rect -2325 28958 -2320 29004
rect -2309 28988 -2301 28998
rect -2317 28982 -2309 28988
rect -2097 28982 -2095 28991
rect -2309 28960 -2301 28970
rect -2097 28968 -2095 28972
rect -2292 28967 -2095 28968
rect -2097 28965 -2095 28967
rect -2084 28960 -2083 29003
rect -2069 28996 -2054 28998
rect -2054 28980 -2018 28982
rect -2054 28978 -2004 28980
rect -2059 28974 -2045 28978
rect -2054 28972 -2049 28974
rect -2317 28958 -2309 28960
rect -2084 28958 -2054 28960
rect -2044 28958 -2039 28972
rect -2025 28962 -2014 28968
rect -2000 28962 -1992 29004
rect -1920 29002 -1906 29004
rect -1977 28987 -1929 28993
rect -1655 28988 -1647 28998
rect -1977 28977 -1966 28987
rect -1663 28982 -1655 28988
rect -1977 28965 -1929 28967
rect -2033 28958 -1992 28962
rect -1655 28960 -1647 28970
rect -1663 28958 -1655 28960
rect -1642 28958 -1637 29004
rect -1619 28958 -1614 29004
rect -1530 28958 -1526 29004
rect -1506 28958 -1502 29004
rect -1482 28958 -1478 29004
rect -1458 28958 -1454 29004
rect -1434 28958 -1430 29004
rect -1410 28958 -1406 29004
rect -1386 28958 -1382 29004
rect -1362 28958 -1358 29004
rect -1338 28958 -1334 29004
rect -1314 28958 -1310 29004
rect -1290 28958 -1286 29004
rect -1266 28958 -1262 29004
rect -1242 28958 -1238 29004
rect -1218 28958 -1214 29004
rect -1194 28958 -1190 29004
rect -1170 28958 -1166 29004
rect -1146 28958 -1142 29004
rect -1122 28958 -1118 29004
rect -1109 28997 -1104 29004
rect -1099 28983 -1094 28997
rect -1098 28958 -1094 28983
rect -1074 28958 -1070 29052
rect -1050 28958 -1046 29052
rect -1026 28958 -1022 29052
rect -1002 28958 -998 29052
rect -978 28958 -974 29052
rect -954 28958 -950 29052
rect -930 28958 -926 29052
rect -906 28958 -902 29052
rect -882 28958 -878 29052
rect -858 28958 -854 29052
rect -834 28958 -830 29052
rect -810 28958 -806 29052
rect -786 28958 -782 29052
rect -762 28958 -758 29052
rect -738 28958 -734 29052
rect -714 28958 -710 29052
rect -690 28958 -686 29052
rect -666 28958 -662 29052
rect -642 28958 -638 29052
rect -618 28958 -614 29052
rect -594 28958 -590 29052
rect -570 28958 -566 29052
rect -546 28958 -542 29052
rect -522 28958 -518 29052
rect -498 28958 -494 29052
rect -474 28958 -470 29052
rect -450 28958 -446 29052
rect -426 28958 -422 29052
rect -402 28958 -398 29052
rect -378 28958 -374 29052
rect -354 28958 -350 29052
rect -330 28958 -326 29052
rect -306 28958 -302 29052
rect -282 28958 -278 29052
rect -258 28958 -254 29052
rect -234 28958 -230 29052
rect -210 28958 -206 29052
rect -186 28958 -182 29052
rect -162 28958 -158 29052
rect -138 28958 -134 29052
rect -114 28958 -110 29052
rect -90 28958 -86 29052
rect -66 28958 -62 29052
rect -42 28958 -38 29052
rect -18 28958 -14 29052
rect 6 28958 10 29052
rect 30 28958 34 29052
rect 54 28958 58 29052
rect 78 28958 82 29052
rect 102 28958 106 29052
rect 126 28958 130 29052
rect 150 28958 154 29052
rect 174 28958 178 29052
rect 198 28958 202 29052
rect 222 28958 226 29052
rect 246 28958 250 29052
rect 270 28958 274 29052
rect 294 28958 298 29052
rect 318 28958 322 29052
rect 342 28958 346 29052
rect 366 28958 370 29052
rect 390 28958 394 29052
rect 414 28958 418 29052
rect 438 28958 442 29052
rect 462 28958 466 29052
rect 486 28958 490 29052
rect 510 28958 514 29052
rect 534 29051 538 29052
rect 534 29030 541 29051
rect 558 29030 562 29052
rect 582 29030 586 29052
rect 606 29030 610 29052
rect 630 29030 634 29052
rect 654 29030 658 29052
rect 678 29030 682 29052
rect 702 29030 706 29052
rect 726 29030 730 29052
rect 750 29030 754 29052
rect 774 29030 778 29052
rect 798 29030 802 29052
rect 822 29030 826 29052
rect 846 29030 850 29052
rect 870 29030 874 29052
rect 894 29030 898 29052
rect 918 29030 922 29052
rect 942 29030 946 29052
rect 966 29030 970 29052
rect 990 29030 994 29052
rect 1014 29030 1018 29052
rect 1038 29030 1042 29052
rect 1062 29030 1066 29052
rect 1086 29030 1090 29052
rect 1110 29030 1114 29052
rect 1134 29030 1138 29052
rect 1158 29030 1162 29052
rect 1182 29030 1186 29052
rect 1206 29030 1210 29052
rect 1230 29030 1234 29052
rect 1254 29030 1258 29052
rect 1278 29030 1282 29052
rect 1302 29030 1306 29052
rect 1326 29030 1330 29052
rect 1350 29030 1354 29052
rect 1374 29030 1378 29052
rect 1398 29030 1402 29052
rect 1422 29030 1426 29052
rect 1446 29030 1450 29052
rect 1470 29030 1474 29052
rect 1494 29030 1498 29052
rect 1518 29030 1522 29052
rect 1542 29030 1546 29052
rect 1566 29030 1570 29052
rect 1590 29030 1594 29052
rect 1614 29030 1618 29052
rect 1638 29030 1642 29052
rect 1662 29030 1666 29052
rect 1686 29030 1690 29052
rect 1710 29030 1714 29052
rect 1734 29030 1738 29052
rect 1758 29030 1762 29052
rect 1782 29030 1786 29052
rect 1806 29030 1810 29052
rect 1830 29030 1834 29052
rect 1854 29030 1858 29052
rect 1878 29030 1882 29052
rect 1902 29030 1906 29052
rect 1926 29030 1930 29052
rect 1950 29030 1954 29052
rect 1974 29030 1978 29052
rect 1998 29030 2002 29052
rect 2022 29030 2026 29052
rect 2035 29045 2040 29052
rect 2046 29045 2050 29052
rect 2053 29051 2067 29052
rect 2045 29031 2050 29045
rect 2059 29041 2067 29045
rect 2053 29031 2059 29041
rect 2035 29030 2067 29031
rect 517 29028 2067 29030
rect 517 29027 531 29028
rect 534 29003 541 29028
rect 534 28958 538 29003
rect 558 28958 562 29028
rect 582 28958 586 29028
rect 606 28958 610 29028
rect 630 28958 634 29028
rect 654 28958 658 29028
rect 678 28958 682 29028
rect 702 28958 706 29028
rect 726 28958 730 29028
rect 750 28958 754 29028
rect 774 28958 778 29028
rect 798 28958 802 29028
rect 822 28958 826 29028
rect 846 28958 850 29028
rect 870 28958 874 29028
rect 894 28958 898 29028
rect 918 28958 922 29028
rect 942 28958 946 29028
rect 966 28958 970 29028
rect 990 29003 994 29028
rect 990 28979 997 29003
rect 990 28958 994 28979
rect 1014 28958 1018 29028
rect 1038 28958 1042 29028
rect 1062 28958 1066 29028
rect 1086 28958 1090 29028
rect 1110 28958 1114 29028
rect 1134 28958 1138 29028
rect 1158 28958 1162 29028
rect 1182 28958 1186 29028
rect 1206 28958 1210 29028
rect 1230 28958 1234 29028
rect 1254 28958 1258 29028
rect 1278 28958 1282 29028
rect 1302 28958 1306 29028
rect 1326 28958 1330 29028
rect 1350 28958 1354 29028
rect 1374 28958 1378 29028
rect 1398 28958 1402 29028
rect 1422 28958 1426 29028
rect 1446 28958 1450 29028
rect 1470 28958 1474 29028
rect 1494 28958 1498 29028
rect 1518 28958 1522 29028
rect 1542 28958 1546 29028
rect 1566 28958 1570 29028
rect 1590 28958 1594 29028
rect 1614 28958 1618 29028
rect 1638 28958 1642 29028
rect 1662 28958 1666 29028
rect 1686 28958 1690 29028
rect 1710 28958 1714 29028
rect 1734 28958 1738 29028
rect 1758 28958 1762 29028
rect 1782 28958 1786 29028
rect 1806 28958 1810 29028
rect 1830 28958 1834 29028
rect 1854 28958 1858 29028
rect 1878 28958 1882 29028
rect 1902 28958 1906 29028
rect 1926 28958 1930 29028
rect 1950 28958 1954 29028
rect 1974 28958 1978 29028
rect 1998 28958 2002 29028
rect 2022 28958 2026 29028
rect 2035 29021 2040 29028
rect 2053 29027 2067 29028
rect 2045 29007 2050 29021
rect 2046 28959 2050 29007
rect 2035 28958 2067 28959
rect -2393 28956 2067 28958
rect -2371 28862 -2366 28956
rect -2348 28862 -2343 28956
rect -2325 28922 -2320 28956
rect -2317 28954 -2309 28956
rect -2084 28943 -2083 28956
rect -2084 28942 -2054 28943
rect -2325 28914 -2317 28922
rect -2325 28862 -2320 28914
rect -2317 28906 -2309 28914
rect -2117 28905 -2095 28915
rect -2045 28912 -2037 28926
rect -2309 28866 -2301 28876
rect -2087 28872 -2076 28880
rect -2017 28876 -2015 28883
rect -2317 28862 -2309 28866
rect -2092 28864 -2087 28872
rect -2092 28862 -2077 28863
rect -2000 28862 -1992 28956
rect -1663 28954 -1655 28956
rect -1969 28905 -1929 28917
rect -1671 28914 -1663 28922
rect -1663 28906 -1655 28914
rect -1655 28866 -1647 28876
rect -1928 28862 -1924 28863
rect -1854 28862 -1680 28863
rect -1663 28862 -1655 28866
rect -1642 28862 -1637 28956
rect -1619 28862 -1614 28956
rect -1530 28862 -1526 28956
rect -1506 28862 -1502 28956
rect -1482 28862 -1478 28956
rect -1458 28862 -1454 28956
rect -1434 28862 -1430 28956
rect -1410 28862 -1406 28956
rect -1386 28862 -1382 28956
rect -1362 28862 -1358 28956
rect -1338 28862 -1334 28956
rect -1314 28862 -1310 28956
rect -1290 28862 -1286 28956
rect -1266 28862 -1262 28956
rect -1242 28862 -1238 28956
rect -1218 28862 -1214 28956
rect -1194 28862 -1190 28956
rect -1170 28862 -1166 28956
rect -1146 28862 -1142 28956
rect -1122 28862 -1118 28956
rect -1098 28862 -1094 28956
rect -1074 28955 -1070 28956
rect -1074 28934 -1067 28955
rect -1050 28934 -1046 28956
rect -1026 28934 -1022 28956
rect -1002 28934 -998 28956
rect -978 28934 -974 28956
rect -954 28934 -950 28956
rect -930 28934 -926 28956
rect -906 28934 -902 28956
rect -882 28934 -878 28956
rect -858 28934 -854 28956
rect -834 28934 -830 28956
rect -810 28934 -806 28956
rect -786 28934 -782 28956
rect -762 28934 -758 28956
rect -738 28934 -734 28956
rect -714 28934 -710 28956
rect -690 28934 -686 28956
rect -666 28934 -662 28956
rect -642 28934 -638 28956
rect -618 28934 -614 28956
rect -594 28934 -590 28956
rect -570 28934 -566 28956
rect -546 28934 -542 28956
rect -522 28934 -518 28956
rect -498 28934 -494 28956
rect -474 28934 -470 28956
rect -450 28934 -446 28956
rect -426 28934 -422 28956
rect -402 28934 -398 28956
rect -378 28934 -374 28956
rect -354 28934 -350 28956
rect -330 28934 -326 28956
rect -306 28934 -302 28956
rect -282 28934 -278 28956
rect -258 28934 -254 28956
rect -234 28934 -230 28956
rect -210 28934 -206 28956
rect -186 28934 -182 28956
rect -162 28934 -158 28956
rect -138 28934 -134 28956
rect -114 28934 -110 28956
rect -90 28934 -86 28956
rect -66 28934 -62 28956
rect -42 28934 -38 28956
rect -18 28934 -14 28956
rect 6 28934 10 28956
rect 30 28934 34 28956
rect 54 28934 58 28956
rect 78 28934 82 28956
rect 102 28934 106 28956
rect 126 28934 130 28956
rect 150 28934 154 28956
rect 174 28934 178 28956
rect 198 28934 202 28956
rect 222 28934 226 28956
rect 246 28934 250 28956
rect 270 28934 274 28956
rect 294 28934 298 28956
rect 318 28934 322 28956
rect 342 28934 346 28956
rect 366 28934 370 28956
rect 390 28934 394 28956
rect 414 28934 418 28956
rect 438 28934 442 28956
rect 462 28934 466 28956
rect 486 28934 490 28956
rect 510 28934 514 28956
rect 534 28934 538 28956
rect 558 28934 562 28956
rect 582 28934 586 28956
rect 606 28934 610 28956
rect 630 28934 634 28956
rect 654 28934 658 28956
rect 678 28934 682 28956
rect 702 28934 706 28956
rect 726 28934 730 28956
rect 750 28934 754 28956
rect 774 28934 778 28956
rect 798 28934 802 28956
rect 822 28934 826 28956
rect 846 28934 850 28956
rect 870 28934 874 28956
rect 894 28934 898 28956
rect 918 28934 922 28956
rect 942 28934 946 28956
rect 966 28934 970 28956
rect 990 28934 994 28956
rect 1014 28934 1018 28956
rect 1038 28934 1042 28956
rect 1062 28934 1066 28956
rect 1086 28934 1090 28956
rect 1110 28934 1114 28956
rect 1134 28934 1138 28956
rect 1158 28934 1162 28956
rect 1182 28934 1186 28956
rect 1206 28934 1210 28956
rect 1230 28934 1234 28956
rect 1254 28934 1258 28956
rect 1278 28934 1282 28956
rect 1302 28934 1306 28956
rect 1326 28934 1330 28956
rect 1350 28934 1354 28956
rect 1374 28934 1378 28956
rect 1398 28934 1402 28956
rect 1422 28934 1426 28956
rect 1446 28934 1450 28956
rect 1470 28934 1474 28956
rect 1494 28934 1498 28956
rect 1518 28934 1522 28956
rect 1542 28934 1546 28956
rect 1566 28934 1570 28956
rect 1590 28934 1594 28956
rect 1614 28934 1618 28956
rect 1638 28934 1642 28956
rect 1662 28934 1666 28956
rect 1686 28934 1690 28956
rect 1710 28934 1714 28956
rect 1734 28934 1738 28956
rect 1758 28934 1762 28956
rect 1782 28934 1786 28956
rect 1806 28934 1810 28956
rect 1830 28934 1834 28956
rect 1854 28934 1858 28956
rect 1878 28934 1882 28956
rect 1902 28934 1906 28956
rect 1926 28934 1930 28956
rect 1950 28934 1954 28956
rect 1974 28934 1978 28956
rect 1998 28934 2002 28956
rect 2022 28935 2026 28956
rect 2035 28949 2040 28956
rect 2046 28949 2050 28956
rect 2053 28955 2067 28956
rect 2045 28935 2050 28949
rect 2059 28945 2067 28949
rect 2053 28935 2059 28945
rect 2011 28934 2045 28935
rect -1091 28932 2045 28934
rect -1091 28931 -1077 28932
rect -1074 28907 -1067 28932
rect -1074 28862 -1070 28907
rect -1050 28862 -1046 28932
rect -1026 28862 -1022 28932
rect -1002 28862 -998 28932
rect -978 28862 -974 28932
rect -954 28862 -950 28932
rect -930 28862 -926 28932
rect -906 28862 -902 28932
rect -882 28862 -878 28932
rect -858 28862 -854 28932
rect -834 28862 -830 28932
rect -810 28862 -806 28932
rect -786 28862 -782 28932
rect -762 28862 -758 28932
rect -738 28862 -734 28932
rect -714 28862 -710 28932
rect -690 28862 -686 28932
rect -666 28862 -662 28932
rect -642 28862 -638 28932
rect -618 28862 -614 28932
rect -594 28862 -590 28932
rect -570 28862 -566 28932
rect -546 28862 -542 28932
rect -522 28862 -518 28932
rect -509 28901 -504 28911
rect -498 28901 -494 28932
rect -499 28887 -494 28901
rect -509 28877 -504 28887
rect -499 28863 -494 28877
rect -498 28862 -494 28863
rect -474 28862 -470 28932
rect -450 28862 -446 28932
rect -426 28862 -422 28932
rect -402 28862 -398 28932
rect -378 28862 -374 28932
rect -354 28862 -350 28932
rect -330 28862 -326 28932
rect -306 28862 -302 28932
rect -282 28862 -278 28932
rect -258 28862 -254 28932
rect -234 28862 -230 28932
rect -210 28862 -206 28932
rect -186 28862 -182 28932
rect -162 28862 -158 28932
rect -138 28862 -134 28932
rect -114 28862 -110 28932
rect -90 28862 -86 28932
rect -66 28862 -62 28932
rect -42 28862 -38 28932
rect -18 28862 -14 28932
rect 6 28862 10 28932
rect 30 28862 34 28932
rect 54 28862 58 28932
rect 78 28862 82 28932
rect 102 28862 106 28932
rect 126 28862 130 28932
rect 150 28862 154 28932
rect 174 28862 178 28932
rect 198 28862 202 28932
rect 222 28862 226 28932
rect 246 28862 250 28932
rect 270 28862 274 28932
rect 294 28862 298 28932
rect 318 28862 322 28932
rect 342 28862 346 28932
rect 366 28862 370 28932
rect 390 28862 394 28932
rect 414 28862 418 28932
rect 438 28862 442 28932
rect 462 28862 466 28932
rect 486 28862 490 28932
rect 510 28862 514 28932
rect 534 28862 538 28932
rect 558 28862 562 28932
rect 582 28862 586 28932
rect 606 28862 610 28932
rect 630 28862 634 28932
rect 654 28862 658 28932
rect 678 28862 682 28932
rect 702 28862 706 28932
rect 726 28862 730 28932
rect 750 28862 754 28932
rect 774 28862 778 28932
rect 798 28862 802 28932
rect 822 28862 826 28932
rect 846 28862 850 28932
rect 870 28862 874 28932
rect 894 28862 898 28932
rect 918 28862 922 28932
rect 942 28862 946 28932
rect 966 28862 970 28932
rect 990 28862 994 28932
rect 1014 28862 1018 28932
rect 1038 28862 1042 28932
rect 1062 28862 1066 28932
rect 1086 28862 1090 28932
rect 1110 28862 1114 28932
rect 1134 28862 1138 28932
rect 1158 28862 1162 28932
rect 1182 28862 1186 28932
rect 1206 28862 1210 28932
rect 1230 28862 1234 28932
rect 1254 28862 1258 28932
rect 1278 28862 1282 28932
rect 1302 28862 1306 28932
rect 1326 28862 1330 28932
rect 1350 28862 1354 28932
rect 1374 28862 1378 28932
rect 1398 28862 1402 28932
rect 1422 28862 1426 28932
rect 1446 28862 1450 28932
rect 1470 28862 1474 28932
rect 1494 28862 1498 28932
rect 1518 28862 1522 28932
rect 1542 28862 1546 28932
rect 1566 28862 1570 28932
rect 1590 28862 1594 28932
rect 1614 28862 1618 28932
rect 1638 28862 1642 28932
rect 1662 28862 1666 28932
rect 1686 28862 1690 28932
rect 1710 28862 1714 28932
rect 1734 28862 1738 28932
rect 1758 28862 1762 28932
rect 1782 28862 1786 28932
rect 1806 28862 1810 28932
rect 1830 28862 1834 28932
rect 1854 28862 1858 28932
rect 1878 28862 1882 28932
rect 1902 28862 1906 28932
rect 1926 28862 1930 28932
rect 1950 28862 1954 28932
rect 1974 28862 1978 28932
rect 1998 28862 2002 28932
rect 2011 28925 2016 28932
rect 2022 28925 2026 28932
rect 2021 28911 2026 28925
rect 2011 28901 2016 28911
rect 2021 28887 2026 28901
rect 2022 28863 2026 28887
rect 2011 28862 2045 28863
rect -2393 28860 2045 28862
rect -2371 28838 -2366 28860
rect -2348 28838 -2343 28860
rect -2325 28838 -2320 28860
rect -2092 28855 -2037 28860
rect -2021 28855 -1969 28860
rect -1921 28855 -1913 28860
rect -1854 28856 -1680 28860
rect -2100 28853 -2092 28854
rect -2309 28838 -2301 28848
rect -2100 28847 -2087 28853
rect -2051 28840 -2026 28842
rect -2062 28838 -2012 28840
rect -2000 28838 -1992 28855
rect -1969 28847 -1921 28854
rect -1969 28838 -1964 28847
rect -1864 28838 -1796 28839
rect -1655 28838 -1647 28848
rect -1642 28838 -1637 28860
rect -1619 28838 -1614 28860
rect -1530 28838 -1526 28860
rect -1506 28838 -1502 28860
rect -1482 28838 -1478 28860
rect -1458 28838 -1454 28860
rect -1434 28838 -1430 28860
rect -1410 28838 -1406 28860
rect -1386 28838 -1382 28860
rect -1362 28838 -1358 28860
rect -1338 28838 -1334 28860
rect -1314 28838 -1310 28860
rect -1290 28838 -1286 28860
rect -1266 28838 -1262 28860
rect -1242 28838 -1238 28860
rect -1218 28838 -1214 28860
rect -1194 28838 -1190 28860
rect -1170 28838 -1166 28860
rect -1146 28838 -1142 28860
rect -1122 28838 -1118 28860
rect -1098 28838 -1094 28860
rect -1074 28838 -1070 28860
rect -1050 28838 -1046 28860
rect -1026 28838 -1022 28860
rect -1002 28838 -998 28860
rect -978 28838 -974 28860
rect -954 28838 -950 28860
rect -930 28838 -926 28860
rect -906 28838 -902 28860
rect -882 28838 -878 28860
rect -858 28838 -854 28860
rect -834 28838 -830 28860
rect -810 28838 -806 28860
rect -786 28838 -782 28860
rect -762 28838 -758 28860
rect -738 28838 -734 28860
rect -714 28838 -710 28860
rect -690 28838 -686 28860
rect -666 28838 -662 28860
rect -642 28838 -638 28860
rect -618 28838 -614 28860
rect -594 28838 -590 28860
rect -570 28838 -566 28860
rect -546 28838 -542 28860
rect -522 28838 -518 28860
rect -498 28838 -494 28860
rect -474 28838 -470 28860
rect -450 28838 -446 28860
rect -426 28838 -422 28860
rect -402 28838 -398 28860
rect -378 28838 -374 28860
rect -354 28838 -350 28860
rect -330 28838 -326 28860
rect -306 28838 -302 28860
rect -282 28838 -278 28860
rect -258 28838 -254 28860
rect -234 28838 -230 28860
rect -210 28838 -206 28860
rect -186 28838 -182 28860
rect -162 28838 -158 28860
rect -138 28838 -134 28860
rect -114 28838 -110 28860
rect -90 28838 -86 28860
rect -66 28838 -62 28860
rect -42 28838 -38 28860
rect -18 28838 -14 28860
rect 6 28838 10 28860
rect 30 28838 34 28860
rect 54 28838 58 28860
rect 78 28838 82 28860
rect 102 28838 106 28860
rect 126 28839 130 28860
rect 115 28838 149 28839
rect -2393 28836 149 28838
rect -2371 28790 -2366 28836
rect -2348 28790 -2343 28836
rect -2325 28790 -2320 28836
rect -2317 28832 -2309 28836
rect -2105 28829 -2092 28832
rect -2092 28806 -2062 28808
rect -2094 28802 -2062 28806
rect -2000 28790 -1992 28836
rect -1663 28832 -1655 28836
rect -1969 28829 -1921 28832
rect -1854 28806 -1806 28808
rect -1854 28802 -1680 28806
rect -1642 28790 -1637 28836
rect -1619 28790 -1614 28836
rect -1530 28790 -1526 28836
rect -1506 28790 -1502 28836
rect -1482 28790 -1478 28836
rect -1458 28790 -1454 28836
rect -1434 28790 -1430 28836
rect -1410 28790 -1406 28836
rect -1386 28790 -1382 28836
rect -1362 28790 -1358 28836
rect -1338 28790 -1334 28836
rect -1314 28790 -1310 28836
rect -1290 28790 -1286 28836
rect -1266 28790 -1262 28836
rect -1242 28790 -1238 28836
rect -1218 28790 -1214 28836
rect -1194 28790 -1190 28836
rect -1170 28790 -1166 28836
rect -1157 28805 -1152 28815
rect -1146 28805 -1142 28836
rect -1147 28791 -1142 28805
rect -1157 28790 -1123 28791
rect -2393 28788 -1123 28790
rect -2371 28766 -2366 28788
rect -2348 28766 -2343 28788
rect -2325 28766 -2320 28788
rect -2072 28786 -2036 28787
rect -2072 28780 -2054 28786
rect -2309 28772 -2301 28780
rect -2317 28766 -2309 28772
rect -2092 28771 -2062 28776
rect -2000 28767 -1992 28788
rect -1938 28787 -1906 28788
rect -1920 28786 -1906 28787
rect -1806 28780 -1680 28786
rect -1854 28771 -1806 28776
rect -1655 28772 -1647 28780
rect -1982 28767 -1966 28768
rect -2000 28766 -1966 28767
rect -1846 28766 -1806 28769
rect -1663 28766 -1655 28772
rect -1642 28766 -1637 28788
rect -1619 28766 -1614 28788
rect -1530 28766 -1526 28788
rect -1506 28766 -1502 28788
rect -1482 28766 -1478 28788
rect -1458 28766 -1454 28788
rect -1434 28766 -1430 28788
rect -1410 28766 -1406 28788
rect -1386 28766 -1382 28788
rect -1362 28766 -1358 28788
rect -1338 28766 -1334 28788
rect -1314 28766 -1310 28788
rect -1290 28766 -1286 28788
rect -1266 28766 -1262 28788
rect -1242 28766 -1238 28788
rect -1218 28766 -1214 28788
rect -1194 28766 -1190 28788
rect -1170 28766 -1166 28788
rect -1157 28781 -1152 28788
rect -1147 28767 -1142 28781
rect -1146 28766 -1142 28767
rect -1122 28766 -1118 28836
rect -1098 28766 -1094 28836
rect -1074 28766 -1070 28836
rect -1050 28766 -1046 28836
rect -1026 28766 -1022 28836
rect -1002 28766 -998 28836
rect -978 28766 -974 28836
rect -954 28766 -950 28836
rect -930 28766 -926 28836
rect -906 28766 -902 28836
rect -882 28766 -878 28836
rect -858 28766 -854 28836
rect -834 28766 -830 28836
rect -810 28766 -806 28836
rect -786 28766 -782 28836
rect -762 28766 -758 28836
rect -738 28766 -734 28836
rect -714 28766 -710 28836
rect -690 28766 -686 28836
rect -666 28766 -662 28836
rect -642 28766 -638 28836
rect -618 28766 -614 28836
rect -594 28766 -590 28836
rect -570 28766 -566 28836
rect -546 28766 -542 28836
rect -522 28766 -518 28836
rect -498 28766 -494 28836
rect -474 28835 -470 28836
rect -474 28814 -467 28835
rect -450 28814 -446 28836
rect -426 28814 -422 28836
rect -402 28814 -398 28836
rect -378 28814 -374 28836
rect -354 28814 -350 28836
rect -330 28814 -326 28836
rect -306 28814 -302 28836
rect -282 28814 -278 28836
rect -258 28814 -254 28836
rect -234 28814 -230 28836
rect -210 28814 -206 28836
rect -186 28814 -182 28836
rect -162 28814 -158 28836
rect -138 28814 -134 28836
rect -114 28814 -110 28836
rect -90 28814 -86 28836
rect -66 28814 -62 28836
rect -42 28814 -38 28836
rect -18 28814 -14 28836
rect 6 28814 10 28836
rect 30 28814 34 28836
rect 54 28814 58 28836
rect 78 28814 82 28836
rect 102 28814 106 28836
rect 115 28829 120 28836
rect 126 28829 130 28836
rect 125 28815 130 28829
rect 126 28814 130 28815
rect 150 28814 154 28860
rect 174 28814 178 28860
rect 198 28814 202 28860
rect 222 28814 226 28860
rect 246 28814 250 28860
rect 270 28814 274 28860
rect 294 28814 298 28860
rect 318 28814 322 28860
rect 342 28814 346 28860
rect 366 28814 370 28860
rect 390 28814 394 28860
rect 414 28814 418 28860
rect 438 28814 442 28860
rect 462 28814 466 28860
rect 486 28814 490 28860
rect 510 28814 514 28860
rect 534 28814 538 28860
rect 558 28814 562 28860
rect 582 28814 586 28860
rect 606 28814 610 28860
rect 630 28814 634 28860
rect 654 28814 658 28860
rect 678 28814 682 28860
rect 702 28814 706 28860
rect 726 28814 730 28860
rect 750 28814 754 28860
rect 774 28814 778 28860
rect 798 28814 802 28860
rect 822 28814 826 28860
rect 846 28814 850 28860
rect 870 28814 874 28860
rect 894 28814 898 28860
rect 918 28814 922 28860
rect 942 28814 946 28860
rect 966 28814 970 28860
rect 990 28814 994 28860
rect 1014 28814 1018 28860
rect 1038 28814 1042 28860
rect 1062 28814 1066 28860
rect 1086 28814 1090 28860
rect 1110 28814 1114 28860
rect 1134 28814 1138 28860
rect 1158 28814 1162 28860
rect 1182 28814 1186 28860
rect 1206 28814 1210 28860
rect 1230 28814 1234 28860
rect 1254 28814 1258 28860
rect 1278 28814 1282 28860
rect 1302 28814 1306 28860
rect 1326 28814 1330 28860
rect 1350 28814 1354 28860
rect 1374 28814 1378 28860
rect 1398 28814 1402 28860
rect 1422 28814 1426 28860
rect 1446 28814 1450 28860
rect 1470 28814 1474 28860
rect 1494 28814 1498 28860
rect 1518 28814 1522 28860
rect 1542 28814 1546 28860
rect 1566 28814 1570 28860
rect 1590 28814 1594 28860
rect 1614 28814 1618 28860
rect 1638 28814 1642 28860
rect 1662 28814 1666 28860
rect 1686 28814 1690 28860
rect 1710 28814 1714 28860
rect 1734 28814 1738 28860
rect 1758 28814 1762 28860
rect 1782 28814 1786 28860
rect 1806 28814 1810 28860
rect 1830 28814 1834 28860
rect 1854 28814 1858 28860
rect 1878 28814 1882 28860
rect 1902 28814 1906 28860
rect 1926 28814 1930 28860
rect 1950 28814 1954 28860
rect 1974 28814 1978 28860
rect 1998 28814 2002 28860
rect 2011 28853 2016 28860
rect 2022 28853 2026 28860
rect 2021 28839 2026 28853
rect 2035 28849 2043 28853
rect 2029 28839 2035 28849
rect 2011 28814 2043 28815
rect -491 28812 2043 28814
rect -491 28811 -477 28812
rect -474 28787 -467 28812
rect -474 28766 -470 28787
rect -450 28766 -446 28812
rect -426 28766 -422 28812
rect -402 28766 -398 28812
rect -378 28766 -374 28812
rect -354 28766 -350 28812
rect -330 28766 -326 28812
rect -306 28766 -302 28812
rect -282 28766 -278 28812
rect -258 28766 -254 28812
rect -234 28766 -230 28812
rect -210 28766 -206 28812
rect -186 28766 -182 28812
rect -162 28766 -158 28812
rect -138 28766 -134 28812
rect -114 28766 -110 28812
rect -90 28766 -86 28812
rect -66 28766 -62 28812
rect -42 28766 -38 28812
rect -18 28766 -14 28812
rect 6 28766 10 28812
rect 30 28766 34 28812
rect 54 28766 58 28812
rect 78 28766 82 28812
rect 102 28766 106 28812
rect 126 28766 130 28812
rect 150 28766 154 28812
rect 174 28766 178 28812
rect 198 28766 202 28812
rect 222 28766 226 28812
rect 246 28766 250 28812
rect 270 28766 274 28812
rect 294 28766 298 28812
rect 318 28766 322 28812
rect 342 28766 346 28812
rect 366 28766 370 28812
rect 390 28766 394 28812
rect 414 28766 418 28812
rect 438 28766 442 28812
rect 462 28766 466 28812
rect 486 28766 490 28812
rect 510 28766 514 28812
rect 534 28766 538 28812
rect 558 28766 562 28812
rect 582 28766 586 28812
rect 606 28766 610 28812
rect 630 28766 634 28812
rect 654 28766 658 28812
rect 678 28766 682 28812
rect 702 28766 706 28812
rect 726 28766 730 28812
rect 750 28766 754 28812
rect 774 28766 778 28812
rect 798 28766 802 28812
rect 822 28766 826 28812
rect 846 28766 850 28812
rect 870 28766 874 28812
rect 894 28766 898 28812
rect 918 28766 922 28812
rect 942 28766 946 28812
rect 966 28766 970 28812
rect 990 28766 994 28812
rect 1014 28766 1018 28812
rect 1038 28766 1042 28812
rect 1062 28766 1066 28812
rect 1086 28766 1090 28812
rect 1110 28766 1114 28812
rect 1134 28766 1138 28812
rect 1158 28766 1162 28812
rect 1182 28766 1186 28812
rect 1206 28766 1210 28812
rect 1230 28766 1234 28812
rect 1254 28766 1258 28812
rect 1278 28766 1282 28812
rect 1302 28766 1306 28812
rect 1326 28766 1330 28812
rect 1350 28766 1354 28812
rect 1374 28766 1378 28812
rect 1398 28766 1402 28812
rect 1422 28766 1426 28812
rect 1446 28766 1450 28812
rect 1470 28766 1474 28812
rect 1494 28766 1498 28812
rect 1518 28766 1522 28812
rect 1542 28766 1546 28812
rect 1566 28766 1570 28812
rect 1590 28766 1594 28812
rect 1614 28766 1618 28812
rect 1638 28766 1642 28812
rect 1662 28766 1666 28812
rect 1686 28766 1690 28812
rect 1710 28766 1714 28812
rect 1734 28766 1738 28812
rect 1758 28766 1762 28812
rect 1782 28766 1786 28812
rect 1806 28766 1810 28812
rect 1830 28766 1834 28812
rect 1854 28766 1858 28812
rect 1878 28766 1882 28812
rect 1902 28766 1906 28812
rect 1926 28766 1930 28812
rect 1950 28766 1954 28812
rect 1974 28766 1978 28812
rect 1998 28766 2002 28812
rect 2011 28805 2016 28812
rect 2029 28811 2043 28812
rect 2021 28791 2026 28805
rect 2022 28767 2026 28791
rect 2011 28766 2043 28767
rect -2393 28764 2043 28766
rect -2371 28742 -2366 28764
rect -2348 28742 -2343 28764
rect -2325 28742 -2320 28764
rect -2000 28762 -1966 28764
rect -2309 28744 -2301 28752
rect -2062 28751 -2054 28758
rect -2092 28744 -2084 28751
rect -2062 28744 -2026 28746
rect -2317 28742 -2309 28744
rect -2062 28742 -2012 28744
rect -2000 28742 -1992 28762
rect -1982 28761 -1966 28762
rect -1846 28760 -1806 28764
rect -1846 28753 -1798 28758
rect -1806 28751 -1798 28753
rect -1854 28749 -1846 28751
rect -1854 28744 -1806 28749
rect -1655 28744 -1647 28752
rect -1864 28742 -1796 28743
rect -1663 28742 -1655 28744
rect -1642 28742 -1637 28764
rect -1619 28742 -1614 28764
rect -1530 28742 -1526 28764
rect -1506 28742 -1502 28764
rect -1482 28742 -1478 28764
rect -1458 28742 -1454 28764
rect -1434 28742 -1430 28764
rect -1410 28742 -1406 28764
rect -1386 28742 -1382 28764
rect -1362 28742 -1358 28764
rect -1338 28742 -1334 28764
rect -1314 28742 -1310 28764
rect -1290 28742 -1286 28764
rect -1266 28742 -1262 28764
rect -1242 28742 -1238 28764
rect -1218 28742 -1214 28764
rect -1194 28742 -1190 28764
rect -1170 28742 -1166 28764
rect -1146 28742 -1142 28764
rect -1122 28742 -1118 28764
rect -1098 28742 -1094 28764
rect -1074 28742 -1070 28764
rect -1050 28742 -1046 28764
rect -1026 28742 -1022 28764
rect -1002 28742 -998 28764
rect -978 28742 -974 28764
rect -954 28742 -950 28764
rect -930 28742 -926 28764
rect -906 28742 -902 28764
rect -882 28742 -878 28764
rect -858 28742 -854 28764
rect -834 28742 -830 28764
rect -810 28742 -806 28764
rect -786 28742 -782 28764
rect -762 28742 -758 28764
rect -738 28742 -734 28764
rect -714 28742 -710 28764
rect -690 28742 -686 28764
rect -666 28742 -662 28764
rect -642 28742 -638 28764
rect -618 28742 -614 28764
rect -594 28742 -590 28764
rect -570 28742 -566 28764
rect -546 28742 -542 28764
rect -522 28742 -518 28764
rect -498 28742 -494 28764
rect -474 28742 -470 28764
rect -450 28742 -446 28764
rect -426 28742 -422 28764
rect -402 28742 -398 28764
rect -378 28742 -374 28764
rect -354 28742 -350 28764
rect -330 28742 -326 28764
rect -306 28742 -302 28764
rect -282 28742 -278 28764
rect -258 28742 -254 28764
rect -234 28742 -230 28764
rect -210 28742 -206 28764
rect -186 28742 -182 28764
rect -162 28742 -158 28764
rect -138 28742 -134 28764
rect -114 28742 -110 28764
rect -90 28742 -86 28764
rect -66 28742 -62 28764
rect -42 28742 -38 28764
rect -18 28742 -14 28764
rect 6 28742 10 28764
rect 30 28742 34 28764
rect 54 28742 58 28764
rect 78 28742 82 28764
rect 102 28742 106 28764
rect 126 28742 130 28764
rect 150 28763 154 28764
rect -2393 28740 147 28742
rect -2371 28694 -2366 28740
rect -2348 28694 -2343 28740
rect -2325 28694 -2320 28740
rect -2317 28736 -2309 28740
rect -2062 28736 -2054 28740
rect -2154 28732 -2138 28734
rect -2057 28732 -2054 28736
rect -2292 28726 -2054 28732
rect -2052 28726 -2044 28736
rect -2092 28710 -2062 28712
rect -2094 28706 -2062 28710
rect -2000 28694 -1992 28740
rect -1846 28733 -1806 28740
rect -1663 28736 -1655 28740
rect -1846 28726 -1680 28732
rect -1854 28710 -1806 28712
rect -1854 28706 -1680 28710
rect -1642 28694 -1637 28740
rect -1619 28694 -1614 28740
rect -1530 28694 -1526 28740
rect -1506 28694 -1502 28740
rect -1482 28694 -1478 28740
rect -1458 28694 -1454 28740
rect -1434 28694 -1430 28740
rect -1410 28694 -1406 28740
rect -1386 28694 -1382 28740
rect -1362 28694 -1358 28740
rect -1338 28694 -1334 28740
rect -1314 28694 -1310 28740
rect -1290 28694 -1286 28740
rect -1266 28694 -1262 28740
rect -1242 28694 -1238 28740
rect -1218 28694 -1214 28740
rect -1194 28694 -1190 28740
rect -1170 28694 -1166 28740
rect -1146 28694 -1142 28740
rect -1122 28739 -1118 28740
rect -2393 28692 -1125 28694
rect -2371 28670 -2366 28692
rect -2348 28670 -2343 28692
rect -2325 28670 -2320 28692
rect -2072 28690 -2036 28691
rect -2072 28684 -2054 28690
rect -2309 28676 -2301 28684
rect -2317 28670 -2309 28676
rect -2092 28675 -2062 28680
rect -2000 28671 -1992 28692
rect -1938 28691 -1906 28692
rect -1920 28690 -1906 28691
rect -1806 28684 -1680 28690
rect -1854 28675 -1806 28680
rect -1655 28676 -1647 28684
rect -1982 28671 -1966 28672
rect -2000 28670 -1966 28671
rect -1846 28670 -1806 28673
rect -1663 28670 -1655 28676
rect -1642 28670 -1637 28692
rect -1619 28670 -1614 28692
rect -1530 28670 -1526 28692
rect -1506 28670 -1502 28692
rect -1482 28670 -1478 28692
rect -1458 28670 -1454 28692
rect -1434 28670 -1430 28692
rect -1410 28670 -1406 28692
rect -1386 28670 -1382 28692
rect -1362 28670 -1358 28692
rect -1338 28670 -1334 28692
rect -1314 28670 -1310 28692
rect -1290 28670 -1286 28692
rect -1266 28670 -1262 28692
rect -1242 28670 -1238 28692
rect -1218 28670 -1214 28692
rect -1194 28670 -1190 28692
rect -1170 28670 -1166 28692
rect -1146 28670 -1142 28692
rect -1139 28691 -1125 28692
rect -1122 28691 -1115 28739
rect -1122 28670 -1118 28691
rect -1098 28670 -1094 28740
rect -1074 28670 -1070 28740
rect -1050 28670 -1046 28740
rect -1026 28670 -1022 28740
rect -1002 28670 -998 28740
rect -978 28670 -974 28740
rect -954 28670 -950 28740
rect -930 28670 -926 28740
rect -906 28670 -902 28740
rect -882 28670 -878 28740
rect -858 28670 -854 28740
rect -834 28670 -830 28740
rect -810 28670 -806 28740
rect -786 28670 -782 28740
rect -762 28670 -758 28740
rect -738 28671 -734 28740
rect -749 28670 -715 28671
rect -2393 28668 -715 28670
rect -2371 28646 -2366 28668
rect -2348 28646 -2343 28668
rect -2325 28646 -2320 28668
rect -2000 28666 -1966 28668
rect -2309 28648 -2301 28656
rect -2062 28655 -2054 28662
rect -2092 28648 -2084 28655
rect -2062 28648 -2026 28650
rect -2317 28646 -2309 28648
rect -2062 28646 -2012 28648
rect -2000 28646 -1992 28666
rect -1982 28665 -1966 28666
rect -1846 28664 -1806 28668
rect -1846 28657 -1798 28662
rect -1806 28655 -1798 28657
rect -1854 28653 -1846 28655
rect -1854 28648 -1806 28653
rect -1655 28648 -1647 28656
rect -1864 28646 -1796 28647
rect -1663 28646 -1655 28648
rect -1642 28646 -1637 28668
rect -1619 28646 -1614 28668
rect -1530 28646 -1526 28668
rect -1506 28646 -1502 28668
rect -1482 28646 -1478 28668
rect -1458 28646 -1454 28668
rect -1434 28646 -1430 28668
rect -1410 28646 -1406 28668
rect -1386 28646 -1382 28668
rect -1362 28646 -1358 28668
rect -1338 28646 -1334 28668
rect -1314 28646 -1310 28668
rect -1290 28646 -1286 28668
rect -1266 28646 -1262 28668
rect -1242 28646 -1238 28668
rect -1218 28646 -1214 28668
rect -1194 28646 -1190 28668
rect -1170 28646 -1166 28668
rect -1146 28646 -1142 28668
rect -1122 28646 -1118 28668
rect -1098 28646 -1094 28668
rect -1074 28646 -1070 28668
rect -1050 28646 -1046 28668
rect -1026 28646 -1022 28668
rect -1002 28647 -998 28668
rect -1013 28646 -979 28647
rect -2393 28644 -979 28646
rect -2371 28598 -2366 28644
rect -2348 28598 -2343 28644
rect -2325 28598 -2320 28644
rect -2317 28640 -2309 28644
rect -2062 28640 -2054 28644
rect -2154 28636 -2138 28638
rect -2057 28636 -2054 28640
rect -2292 28630 -2054 28636
rect -2052 28630 -2044 28640
rect -2092 28614 -2062 28616
rect -2094 28610 -2062 28614
rect -2000 28598 -1992 28644
rect -1846 28637 -1806 28644
rect -1663 28640 -1655 28644
rect -1846 28630 -1680 28636
rect -1854 28614 -1806 28616
rect -1854 28610 -1680 28614
rect -1642 28598 -1637 28644
rect -1619 28598 -1614 28644
rect -1530 28598 -1526 28644
rect -1506 28598 -1502 28644
rect -1482 28598 -1478 28644
rect -1458 28598 -1454 28644
rect -1434 28598 -1430 28644
rect -1410 28598 -1406 28644
rect -1386 28598 -1382 28644
rect -1362 28598 -1358 28644
rect -1338 28598 -1334 28644
rect -1314 28598 -1310 28644
rect -1290 28598 -1286 28644
rect -1266 28598 -1262 28644
rect -1242 28598 -1238 28644
rect -1218 28598 -1214 28644
rect -1194 28598 -1190 28644
rect -1170 28598 -1166 28644
rect -1146 28598 -1142 28644
rect -1122 28598 -1118 28644
rect -1098 28598 -1094 28644
rect -1074 28598 -1070 28644
rect -1050 28598 -1046 28644
rect -1026 28598 -1022 28644
rect -1013 28637 -1008 28644
rect -1002 28637 -998 28644
rect -1003 28623 -998 28637
rect -1002 28598 -998 28623
rect -978 28598 -974 28668
rect -954 28598 -950 28668
rect -930 28598 -926 28668
rect -906 28598 -902 28668
rect -882 28598 -878 28668
rect -858 28598 -854 28668
rect -834 28598 -830 28668
rect -810 28598 -806 28668
rect -786 28598 -782 28668
rect -762 28598 -758 28668
rect -749 28661 -744 28668
rect -738 28661 -734 28668
rect -739 28647 -734 28661
rect -738 28598 -734 28647
rect -714 28598 -710 28740
rect -690 28598 -686 28740
rect -666 28598 -662 28740
rect -642 28598 -638 28740
rect -618 28598 -614 28740
rect -594 28598 -590 28740
rect -570 28598 -566 28740
rect -546 28598 -542 28740
rect -522 28598 -518 28740
rect -498 28598 -494 28740
rect -474 28598 -470 28740
rect -450 28598 -446 28740
rect -426 28598 -422 28740
rect -402 28598 -398 28740
rect -378 28598 -374 28740
rect -354 28598 -350 28740
rect -330 28598 -326 28740
rect -306 28598 -302 28740
rect -282 28598 -278 28740
rect -258 28598 -254 28740
rect -234 28598 -230 28740
rect -210 28598 -206 28740
rect -186 28598 -182 28740
rect -162 28598 -158 28740
rect -138 28598 -134 28740
rect -114 28598 -110 28740
rect -90 28598 -86 28740
rect -66 28598 -62 28740
rect -42 28598 -38 28740
rect -18 28598 -14 28740
rect 6 28598 10 28740
rect 30 28598 34 28740
rect 54 28598 58 28740
rect 78 28598 82 28740
rect 102 28598 106 28740
rect 126 28598 130 28740
rect 133 28739 147 28740
rect 150 28739 157 28763
rect 150 28598 154 28739
rect 174 28598 178 28764
rect 198 28598 202 28764
rect 222 28598 226 28764
rect 246 28598 250 28764
rect 270 28598 274 28764
rect 294 28598 298 28764
rect 318 28598 322 28764
rect 342 28598 346 28764
rect 366 28598 370 28764
rect 390 28598 394 28764
rect 414 28598 418 28764
rect 438 28598 442 28764
rect 462 28598 466 28764
rect 486 28598 490 28764
rect 510 28598 514 28764
rect 534 28598 538 28764
rect 558 28598 562 28764
rect 582 28598 586 28764
rect 606 28598 610 28764
rect 630 28598 634 28764
rect 654 28598 658 28764
rect 678 28598 682 28764
rect 702 28598 706 28764
rect 726 28598 730 28764
rect 750 28598 754 28764
rect 774 28598 778 28764
rect 798 28598 802 28764
rect 822 28598 826 28764
rect 846 28598 850 28764
rect 870 28598 874 28764
rect 894 28598 898 28764
rect 918 28598 922 28764
rect 942 28598 946 28764
rect 966 28598 970 28764
rect 990 28598 994 28764
rect 1014 28598 1018 28764
rect 1038 28598 1042 28764
rect 1062 28598 1066 28764
rect 1086 28598 1090 28764
rect 1110 28598 1114 28764
rect 1134 28598 1138 28764
rect 1158 28598 1162 28764
rect 1182 28598 1186 28764
rect 1206 28598 1210 28764
rect 1230 28598 1234 28764
rect 1254 28598 1258 28764
rect 1278 28598 1282 28764
rect 1302 28598 1306 28764
rect 1326 28598 1330 28764
rect 1350 28598 1354 28764
rect 1374 28598 1378 28764
rect 1398 28598 1402 28764
rect 1422 28598 1426 28764
rect 1446 28598 1450 28764
rect 1459 28613 1464 28623
rect 1470 28613 1474 28764
rect 1469 28599 1474 28613
rect 1459 28598 1493 28599
rect -2393 28596 1493 28598
rect -2371 28574 -2366 28596
rect -2348 28574 -2343 28596
rect -2325 28574 -2320 28596
rect -2072 28594 -2036 28595
rect -2072 28588 -2054 28594
rect -2309 28580 -2301 28588
rect -2317 28574 -2309 28580
rect -2092 28579 -2062 28584
rect -2000 28575 -1992 28596
rect -1938 28595 -1906 28596
rect -1920 28594 -1906 28595
rect -1806 28588 -1680 28594
rect -1854 28579 -1806 28584
rect -1655 28580 -1647 28588
rect -1982 28575 -1966 28576
rect -2000 28574 -1966 28575
rect -1846 28574 -1806 28577
rect -1663 28574 -1655 28580
rect -1642 28574 -1637 28596
rect -1619 28574 -1614 28596
rect -1530 28574 -1526 28596
rect -1506 28574 -1502 28596
rect -1482 28574 -1478 28596
rect -1458 28574 -1454 28596
rect -1434 28574 -1430 28596
rect -1410 28574 -1406 28596
rect -1386 28574 -1382 28596
rect -1362 28575 -1358 28596
rect -1373 28574 -1339 28575
rect -2393 28572 -1339 28574
rect -2371 28550 -2366 28572
rect -2348 28550 -2343 28572
rect -2325 28550 -2320 28572
rect -2000 28570 -1966 28572
rect -2309 28552 -2301 28560
rect -2062 28559 -2054 28566
rect -2092 28552 -2084 28559
rect -2062 28552 -2026 28554
rect -2317 28550 -2309 28552
rect -2062 28550 -2012 28552
rect -2000 28550 -1992 28570
rect -1982 28569 -1966 28570
rect -1846 28568 -1806 28572
rect -1846 28561 -1798 28566
rect -1806 28559 -1798 28561
rect -1854 28557 -1846 28559
rect -1854 28552 -1806 28557
rect -1655 28552 -1647 28560
rect -1864 28550 -1796 28551
rect -1663 28550 -1655 28552
rect -1642 28550 -1637 28572
rect -1619 28550 -1614 28572
rect -1530 28550 -1526 28572
rect -1506 28550 -1502 28572
rect -1482 28550 -1478 28572
rect -1458 28550 -1454 28572
rect -1434 28550 -1430 28572
rect -1410 28550 -1406 28572
rect -1386 28550 -1382 28572
rect -1373 28565 -1368 28572
rect -1362 28565 -1358 28572
rect -1363 28551 -1358 28565
rect -1362 28550 -1358 28551
rect -1338 28550 -1334 28596
rect -1314 28550 -1310 28596
rect -1290 28550 -1286 28596
rect -1266 28550 -1262 28596
rect -1242 28550 -1238 28596
rect -1218 28550 -1214 28596
rect -1194 28550 -1190 28596
rect -1170 28550 -1166 28596
rect -1146 28550 -1142 28596
rect -1122 28550 -1118 28596
rect -1098 28550 -1094 28596
rect -1074 28550 -1070 28596
rect -1050 28550 -1046 28596
rect -1026 28550 -1022 28596
rect -1002 28550 -998 28596
rect -978 28571 -974 28596
rect -2393 28548 -981 28550
rect -2371 28502 -2366 28548
rect -2348 28502 -2343 28548
rect -2325 28502 -2320 28548
rect -2317 28544 -2309 28548
rect -2062 28544 -2054 28548
rect -2154 28540 -2138 28542
rect -2057 28540 -2054 28544
rect -2292 28534 -2054 28540
rect -2052 28534 -2044 28544
rect -2092 28518 -2062 28520
rect -2094 28514 -2062 28518
rect -2000 28502 -1992 28548
rect -1846 28541 -1806 28548
rect -1663 28544 -1655 28548
rect -1846 28534 -1680 28540
rect -1854 28518 -1806 28520
rect -1854 28514 -1680 28518
rect -1642 28502 -1637 28548
rect -1619 28502 -1614 28548
rect -1530 28502 -1526 28548
rect -1506 28502 -1502 28548
rect -1482 28502 -1478 28548
rect -1458 28502 -1454 28548
rect -1434 28502 -1430 28548
rect -1410 28502 -1406 28548
rect -1386 28502 -1382 28548
rect -1362 28502 -1358 28548
rect -1338 28502 -1334 28548
rect -1314 28502 -1310 28548
rect -1290 28502 -1286 28548
rect -1266 28502 -1262 28548
rect -1242 28502 -1238 28548
rect -1218 28502 -1214 28548
rect -1194 28502 -1190 28548
rect -1170 28502 -1166 28548
rect -1146 28502 -1142 28548
rect -1122 28502 -1118 28548
rect -1098 28502 -1094 28548
rect -1074 28502 -1070 28548
rect -1050 28502 -1046 28548
rect -1026 28502 -1022 28548
rect -1002 28502 -998 28548
rect -995 28547 -981 28548
rect -978 28547 -971 28571
rect -978 28502 -974 28547
rect -954 28502 -950 28596
rect -930 28502 -926 28596
rect -906 28502 -902 28596
rect -882 28502 -878 28596
rect -858 28502 -854 28596
rect -834 28502 -830 28596
rect -810 28502 -806 28596
rect -786 28502 -782 28596
rect -762 28502 -758 28596
rect -738 28502 -734 28596
rect -714 28595 -710 28596
rect -714 28571 -707 28595
rect -714 28502 -710 28571
rect -690 28502 -686 28596
rect -666 28502 -662 28596
rect -642 28502 -638 28596
rect -618 28502 -614 28596
rect -594 28502 -590 28596
rect -570 28502 -566 28596
rect -546 28502 -542 28596
rect -522 28502 -518 28596
rect -498 28502 -494 28596
rect -474 28502 -470 28596
rect -450 28502 -446 28596
rect -426 28502 -422 28596
rect -402 28502 -398 28596
rect -378 28502 -374 28596
rect -354 28502 -350 28596
rect -330 28502 -326 28596
rect -306 28502 -302 28596
rect -282 28502 -278 28596
rect -258 28502 -254 28596
rect -234 28502 -230 28596
rect -210 28502 -206 28596
rect -186 28502 -182 28596
rect -162 28502 -158 28596
rect -138 28502 -134 28596
rect -114 28502 -110 28596
rect -90 28502 -86 28596
rect -66 28502 -62 28596
rect -42 28502 -38 28596
rect -18 28502 -14 28596
rect 6 28502 10 28596
rect 30 28502 34 28596
rect 54 28502 58 28596
rect 78 28502 82 28596
rect 102 28502 106 28596
rect 126 28502 130 28596
rect 150 28502 154 28596
rect 174 28502 178 28596
rect 198 28502 202 28596
rect 222 28502 226 28596
rect 246 28502 250 28596
rect 270 28502 274 28596
rect 294 28502 298 28596
rect 318 28502 322 28596
rect 342 28502 346 28596
rect 366 28502 370 28596
rect 390 28502 394 28596
rect 414 28502 418 28596
rect 438 28502 442 28596
rect 462 28502 466 28596
rect 486 28502 490 28596
rect 510 28502 514 28596
rect 534 28502 538 28596
rect 558 28502 562 28596
rect 582 28502 586 28596
rect 606 28502 610 28596
rect 630 28502 634 28596
rect 654 28502 658 28596
rect 678 28502 682 28596
rect 702 28502 706 28596
rect 726 28502 730 28596
rect 750 28502 754 28596
rect 774 28502 778 28596
rect 798 28502 802 28596
rect 822 28502 826 28596
rect 846 28502 850 28596
rect 870 28502 874 28596
rect 894 28502 898 28596
rect 918 28502 922 28596
rect 942 28502 946 28596
rect 966 28502 970 28596
rect 990 28502 994 28596
rect 1014 28502 1018 28596
rect 1038 28502 1042 28596
rect 1062 28502 1066 28596
rect 1086 28502 1090 28596
rect 1110 28502 1114 28596
rect 1134 28502 1138 28596
rect 1158 28502 1162 28596
rect 1182 28502 1186 28596
rect 1206 28502 1210 28596
rect 1230 28502 1234 28596
rect 1254 28502 1258 28596
rect 1278 28502 1282 28596
rect 1302 28502 1306 28596
rect 1326 28502 1330 28596
rect 1350 28502 1354 28596
rect 1374 28502 1378 28596
rect 1398 28502 1402 28596
rect 1411 28517 1416 28527
rect 1422 28517 1426 28596
rect 1421 28503 1426 28517
rect 1411 28502 1445 28503
rect -2393 28500 1445 28502
rect -2371 28478 -2366 28500
rect -2348 28478 -2343 28500
rect -2325 28478 -2320 28500
rect -2072 28498 -2036 28499
rect -2072 28492 -2054 28498
rect -2309 28484 -2301 28492
rect -2317 28478 -2309 28484
rect -2092 28483 -2062 28488
rect -2000 28479 -1992 28500
rect -1938 28499 -1906 28500
rect -1920 28498 -1906 28499
rect -1806 28492 -1680 28498
rect -1854 28483 -1806 28488
rect -1655 28484 -1647 28492
rect -1982 28479 -1966 28480
rect -2000 28478 -1966 28479
rect -1846 28478 -1806 28481
rect -1663 28478 -1655 28484
rect -1642 28478 -1637 28500
rect -1619 28478 -1614 28500
rect -1530 28478 -1526 28500
rect -1506 28478 -1502 28500
rect -1482 28478 -1478 28500
rect -1458 28478 -1454 28500
rect -1434 28478 -1430 28500
rect -1410 28478 -1406 28500
rect -1386 28478 -1382 28500
rect -1362 28478 -1358 28500
rect -1338 28499 -1334 28500
rect -2393 28476 -1341 28478
rect -2371 28454 -2366 28476
rect -2348 28454 -2343 28476
rect -2325 28454 -2320 28476
rect -2000 28474 -1966 28476
rect -2309 28456 -2301 28464
rect -2062 28463 -2054 28470
rect -2092 28456 -2084 28463
rect -2062 28456 -2026 28458
rect -2317 28454 -2309 28456
rect -2062 28454 -2012 28456
rect -2000 28454 -1992 28474
rect -1982 28473 -1966 28474
rect -1846 28472 -1806 28476
rect -1846 28465 -1798 28470
rect -1806 28463 -1798 28465
rect -1854 28461 -1846 28463
rect -1854 28456 -1806 28461
rect -1655 28456 -1647 28464
rect -1864 28454 -1796 28455
rect -1663 28454 -1655 28456
rect -1642 28454 -1637 28476
rect -1619 28454 -1614 28476
rect -1530 28454 -1526 28476
rect -1506 28454 -1502 28476
rect -1482 28454 -1478 28476
rect -1458 28454 -1454 28476
rect -1434 28454 -1430 28476
rect -1410 28454 -1406 28476
rect -1386 28454 -1382 28476
rect -1362 28454 -1358 28476
rect -1355 28475 -1341 28476
rect -1338 28475 -1331 28499
rect -1338 28454 -1334 28475
rect -1314 28454 -1310 28500
rect -1290 28454 -1286 28500
rect -1266 28454 -1262 28500
rect -1242 28454 -1238 28500
rect -1218 28454 -1214 28500
rect -1194 28454 -1190 28500
rect -1170 28454 -1166 28500
rect -1146 28454 -1142 28500
rect -1122 28454 -1118 28500
rect -1098 28454 -1094 28500
rect -1074 28454 -1070 28500
rect -1050 28454 -1046 28500
rect -1026 28454 -1022 28500
rect -1002 28454 -998 28500
rect -978 28454 -974 28500
rect -954 28454 -950 28500
rect -930 28454 -926 28500
rect -906 28454 -902 28500
rect -882 28454 -878 28500
rect -858 28454 -854 28500
rect -834 28454 -830 28500
rect -810 28454 -806 28500
rect -786 28454 -782 28500
rect -762 28454 -758 28500
rect -738 28454 -734 28500
rect -714 28454 -710 28500
rect -690 28454 -686 28500
rect -666 28454 -662 28500
rect -642 28454 -638 28500
rect -618 28454 -614 28500
rect -594 28454 -590 28500
rect -570 28454 -566 28500
rect -546 28454 -542 28500
rect -522 28454 -518 28500
rect -498 28454 -494 28500
rect -474 28454 -470 28500
rect -450 28454 -446 28500
rect -426 28454 -422 28500
rect -402 28454 -398 28500
rect -378 28454 -374 28500
rect -354 28454 -350 28500
rect -330 28454 -326 28500
rect -306 28454 -302 28500
rect -282 28454 -278 28500
rect -258 28454 -254 28500
rect -234 28454 -230 28500
rect -210 28454 -206 28500
rect -186 28454 -182 28500
rect -162 28454 -158 28500
rect -138 28454 -134 28500
rect -114 28454 -110 28500
rect -90 28454 -86 28500
rect -66 28454 -62 28500
rect -42 28454 -38 28500
rect -18 28454 -14 28500
rect 6 28454 10 28500
rect 30 28454 34 28500
rect 54 28454 58 28500
rect 78 28454 82 28500
rect 102 28454 106 28500
rect 126 28454 130 28500
rect 150 28454 154 28500
rect 174 28454 178 28500
rect 198 28454 202 28500
rect 222 28454 226 28500
rect 246 28454 250 28500
rect 270 28454 274 28500
rect 294 28454 298 28500
rect 318 28454 322 28500
rect 342 28454 346 28500
rect 366 28454 370 28500
rect 390 28454 394 28500
rect 414 28454 418 28500
rect 438 28454 442 28500
rect 462 28454 466 28500
rect 486 28454 490 28500
rect 510 28454 514 28500
rect 534 28454 538 28500
rect 558 28454 562 28500
rect 582 28454 586 28500
rect 606 28454 610 28500
rect 630 28454 634 28500
rect 654 28454 658 28500
rect 678 28454 682 28500
rect 702 28454 706 28500
rect 726 28454 730 28500
rect 750 28454 754 28500
rect 774 28454 778 28500
rect 798 28454 802 28500
rect 822 28454 826 28500
rect 846 28454 850 28500
rect 870 28454 874 28500
rect 894 28454 898 28500
rect 918 28454 922 28500
rect 942 28454 946 28500
rect 966 28454 970 28500
rect 990 28454 994 28500
rect 1014 28454 1018 28500
rect 1038 28454 1042 28500
rect 1062 28454 1066 28500
rect 1086 28454 1090 28500
rect 1110 28454 1114 28500
rect 1134 28454 1138 28500
rect 1158 28454 1162 28500
rect 1182 28454 1186 28500
rect 1206 28454 1210 28500
rect 1230 28454 1234 28500
rect 1254 28454 1258 28500
rect 1278 28454 1282 28500
rect 1302 28454 1306 28500
rect 1326 28454 1330 28500
rect 1350 28454 1354 28500
rect 1374 28454 1378 28500
rect 1398 28454 1402 28500
rect 1411 28493 1416 28500
rect 1421 28479 1426 28493
rect 1422 28454 1426 28479
rect 1446 28454 1450 28596
rect 1459 28589 1464 28596
rect 1469 28575 1474 28589
rect 1470 28454 1474 28575
rect 1494 28547 1498 28764
rect 1494 28526 1501 28547
rect 1518 28526 1522 28764
rect 1542 28526 1546 28764
rect 1566 28526 1570 28764
rect 1590 28526 1594 28764
rect 1614 28526 1618 28764
rect 1638 28526 1642 28764
rect 1662 28526 1666 28764
rect 1686 28526 1690 28764
rect 1710 28526 1714 28764
rect 1734 28526 1738 28764
rect 1758 28526 1762 28764
rect 1782 28526 1786 28764
rect 1806 28526 1810 28764
rect 1830 28526 1834 28764
rect 1854 28526 1858 28764
rect 1878 28526 1882 28764
rect 1902 28526 1906 28764
rect 1926 28719 1930 28764
rect 1915 28718 1949 28719
rect 1950 28718 1954 28764
rect 1974 28718 1978 28764
rect 1987 28733 1992 28743
rect 1998 28733 2002 28764
rect 2011 28757 2016 28764
rect 2022 28757 2026 28764
rect 2029 28763 2043 28764
rect 2021 28743 2026 28757
rect 1997 28719 2002 28733
rect 1987 28718 2021 28719
rect 1915 28716 2021 28718
rect 1915 28709 1920 28716
rect 1926 28709 1930 28716
rect 1925 28695 1930 28709
rect 1915 28685 1920 28695
rect 1925 28671 1930 28685
rect 1926 28526 1930 28671
rect 1950 28643 1954 28716
rect 1950 28622 1957 28643
rect 1974 28622 1978 28716
rect 1987 28709 1992 28716
rect 1997 28695 2002 28709
rect 1998 28622 2002 28695
rect 2011 28622 2019 28623
rect 1933 28620 2019 28622
rect 1933 28619 1947 28620
rect 1950 28595 1957 28620
rect 1950 28526 1954 28595
rect 1974 28526 1978 28620
rect 1998 28526 2002 28620
rect 2005 28619 2019 28620
rect 2011 28613 2016 28619
rect 2021 28599 2026 28613
rect 2011 28541 2016 28551
rect 2022 28541 2026 28599
rect 2021 28527 2026 28541
rect 2035 28537 2043 28541
rect 2029 28527 2035 28537
rect 2011 28526 2043 28527
rect 1477 28524 2043 28526
rect 1477 28523 1491 28524
rect 1494 28499 1501 28524
rect 1494 28454 1498 28499
rect 1518 28454 1522 28524
rect 1542 28454 1546 28524
rect 1566 28454 1570 28524
rect 1590 28454 1594 28524
rect 1614 28454 1618 28524
rect 1638 28454 1642 28524
rect 1662 28454 1666 28524
rect 1686 28454 1690 28524
rect 1710 28454 1714 28524
rect 1734 28454 1738 28524
rect 1758 28454 1762 28524
rect 1782 28454 1786 28524
rect 1806 28454 1810 28524
rect 1830 28454 1834 28524
rect 1854 28454 1858 28524
rect 1878 28454 1882 28524
rect 1902 28454 1906 28524
rect 1926 28454 1930 28524
rect 1950 28454 1954 28524
rect 1974 28454 1978 28524
rect 1998 28455 2002 28524
rect 2011 28517 2016 28524
rect 2029 28523 2043 28524
rect 2021 28503 2026 28517
rect 2011 28469 2016 28479
rect 2022 28469 2026 28503
rect 2021 28455 2026 28469
rect 2035 28465 2043 28469
rect 2029 28455 2035 28465
rect 1987 28454 2021 28455
rect -2393 28452 2021 28454
rect -2371 28406 -2366 28452
rect -2348 28406 -2343 28452
rect -2325 28406 -2320 28452
rect -2317 28448 -2309 28452
rect -2062 28448 -2054 28452
rect -2154 28444 -2138 28446
rect -2057 28444 -2054 28448
rect -2292 28438 -2054 28444
rect -2052 28438 -2044 28448
rect -2092 28422 -2062 28424
rect -2094 28418 -2062 28422
rect -2000 28406 -1992 28452
rect -1846 28445 -1806 28452
rect -1663 28448 -1655 28452
rect -1846 28438 -1680 28444
rect -1854 28422 -1806 28424
rect -1854 28418 -1680 28422
rect -1642 28406 -1637 28452
rect -1619 28406 -1614 28452
rect -1530 28406 -1526 28452
rect -1506 28406 -1502 28452
rect -1482 28406 -1478 28452
rect -1458 28406 -1454 28452
rect -1434 28406 -1430 28452
rect -1410 28406 -1406 28452
rect -1386 28406 -1382 28452
rect -1362 28406 -1358 28452
rect -1338 28406 -1334 28452
rect -1314 28406 -1310 28452
rect -1290 28406 -1286 28452
rect -1266 28406 -1262 28452
rect -1242 28406 -1238 28452
rect -1218 28406 -1214 28452
rect -1194 28406 -1190 28452
rect -1170 28406 -1166 28452
rect -1146 28406 -1142 28452
rect -1122 28406 -1118 28452
rect -1098 28406 -1094 28452
rect -1074 28406 -1070 28452
rect -1050 28406 -1046 28452
rect -1026 28406 -1022 28452
rect -1002 28406 -998 28452
rect -978 28406 -974 28452
rect -954 28406 -950 28452
rect -930 28406 -926 28452
rect -906 28406 -902 28452
rect -882 28406 -878 28452
rect -858 28406 -854 28452
rect -834 28406 -830 28452
rect -810 28406 -806 28452
rect -786 28406 -782 28452
rect -762 28406 -758 28452
rect -738 28406 -734 28452
rect -725 28421 -720 28431
rect -714 28421 -710 28452
rect -715 28407 -710 28421
rect -725 28406 -691 28407
rect -2393 28404 -691 28406
rect -2371 28358 -2366 28404
rect -2348 28358 -2343 28404
rect -2325 28358 -2320 28404
rect -2309 28388 -2301 28398
rect -2317 28382 -2309 28388
rect -2097 28382 -2095 28391
rect -2309 28360 -2301 28370
rect -2097 28368 -2095 28372
rect -2292 28367 -2095 28368
rect -2097 28365 -2095 28367
rect -2084 28360 -2083 28403
rect -2069 28396 -2054 28398
rect -2054 28380 -2018 28382
rect -2054 28378 -2004 28380
rect -2059 28374 -2045 28378
rect -2054 28372 -2049 28374
rect -2317 28358 -2309 28360
rect -2084 28358 -2054 28360
rect -2044 28358 -2039 28372
rect -2025 28362 -2014 28368
rect -2000 28362 -1992 28404
rect -1920 28402 -1906 28404
rect -1977 28387 -1929 28393
rect -1655 28388 -1647 28398
rect -1977 28377 -1966 28387
rect -1663 28382 -1655 28388
rect -1977 28365 -1929 28367
rect -2033 28358 -1992 28362
rect -1655 28360 -1647 28370
rect -1663 28358 -1655 28360
rect -1642 28358 -1637 28404
rect -1619 28358 -1614 28404
rect -1530 28358 -1526 28404
rect -1506 28358 -1502 28404
rect -1482 28358 -1478 28404
rect -1458 28358 -1454 28404
rect -1434 28358 -1430 28404
rect -1410 28358 -1406 28404
rect -1386 28358 -1382 28404
rect -1362 28358 -1358 28404
rect -1338 28358 -1334 28404
rect -1314 28358 -1310 28404
rect -1290 28358 -1286 28404
rect -1266 28358 -1262 28404
rect -1242 28358 -1238 28404
rect -1218 28358 -1214 28404
rect -1194 28358 -1190 28404
rect -1170 28358 -1166 28404
rect -1146 28358 -1142 28404
rect -1122 28358 -1118 28404
rect -1098 28358 -1094 28404
rect -1074 28358 -1070 28404
rect -1050 28358 -1046 28404
rect -1026 28358 -1022 28404
rect -1002 28358 -998 28404
rect -978 28358 -974 28404
rect -954 28358 -950 28404
rect -930 28358 -926 28404
rect -906 28358 -902 28404
rect -882 28358 -878 28404
rect -858 28358 -854 28404
rect -834 28358 -830 28404
rect -810 28358 -806 28404
rect -786 28358 -782 28404
rect -762 28358 -758 28404
rect -738 28358 -734 28404
rect -725 28397 -720 28404
rect -715 28383 -710 28397
rect -714 28358 -710 28383
rect -690 28358 -686 28452
rect -666 28358 -662 28452
rect -642 28358 -638 28452
rect -618 28358 -614 28452
rect -594 28358 -590 28452
rect -570 28358 -566 28452
rect -546 28358 -542 28452
rect -522 28358 -518 28452
rect -498 28358 -494 28452
rect -474 28358 -470 28452
rect -450 28358 -446 28452
rect -426 28358 -422 28452
rect -402 28358 -398 28452
rect -378 28358 -374 28452
rect -354 28358 -350 28452
rect -330 28358 -326 28452
rect -306 28358 -302 28452
rect -282 28358 -278 28452
rect -258 28358 -254 28452
rect -234 28358 -230 28452
rect -210 28358 -206 28452
rect -186 28358 -182 28452
rect -162 28358 -158 28452
rect -138 28358 -134 28452
rect -114 28358 -110 28452
rect -90 28358 -86 28452
rect -66 28358 -62 28452
rect -42 28358 -38 28452
rect -18 28358 -14 28452
rect 6 28358 10 28452
rect 30 28358 34 28452
rect 54 28358 58 28452
rect 78 28358 82 28452
rect 102 28358 106 28452
rect 126 28358 130 28452
rect 150 28358 154 28452
rect 174 28358 178 28452
rect 198 28358 202 28452
rect 222 28358 226 28452
rect 246 28358 250 28452
rect 270 28358 274 28452
rect 294 28358 298 28452
rect 318 28358 322 28452
rect 342 28358 346 28452
rect 366 28358 370 28452
rect 390 28358 394 28452
rect 414 28358 418 28452
rect 438 28358 442 28452
rect 462 28358 466 28452
rect 486 28358 490 28452
rect 510 28358 514 28452
rect 534 28358 538 28452
rect 558 28358 562 28452
rect 582 28358 586 28452
rect 606 28358 610 28452
rect 630 28358 634 28452
rect 654 28358 658 28452
rect 678 28358 682 28452
rect 702 28358 706 28452
rect 726 28358 730 28452
rect 750 28358 754 28452
rect 774 28358 778 28452
rect 798 28358 802 28452
rect 822 28358 826 28452
rect 846 28358 850 28452
rect 870 28358 874 28452
rect 894 28358 898 28452
rect 918 28358 922 28452
rect 942 28358 946 28452
rect 966 28358 970 28452
rect 990 28358 994 28452
rect 1014 28358 1018 28452
rect 1038 28358 1042 28452
rect 1062 28358 1066 28452
rect 1086 28358 1090 28452
rect 1110 28358 1114 28452
rect 1134 28358 1138 28452
rect 1158 28358 1162 28452
rect 1182 28358 1186 28452
rect 1206 28358 1210 28452
rect 1230 28358 1234 28452
rect 1254 28358 1258 28452
rect 1278 28358 1282 28452
rect 1302 28358 1306 28452
rect 1326 28358 1330 28452
rect 1350 28358 1354 28452
rect 1374 28358 1378 28452
rect 1398 28358 1402 28452
rect 1422 28358 1426 28452
rect 1446 28451 1450 28452
rect 1446 28430 1453 28451
rect 1470 28430 1474 28452
rect 1494 28430 1498 28452
rect 1518 28430 1522 28452
rect 1542 28430 1546 28452
rect 1566 28430 1570 28452
rect 1590 28430 1594 28452
rect 1614 28430 1618 28452
rect 1638 28430 1642 28452
rect 1662 28430 1666 28452
rect 1686 28430 1690 28452
rect 1710 28430 1714 28452
rect 1734 28430 1738 28452
rect 1758 28430 1762 28452
rect 1782 28430 1786 28452
rect 1806 28430 1810 28452
rect 1830 28430 1834 28452
rect 1854 28430 1858 28452
rect 1878 28430 1882 28452
rect 1902 28430 1906 28452
rect 1926 28430 1930 28452
rect 1950 28430 1954 28452
rect 1974 28430 1978 28452
rect 1987 28445 1992 28452
rect 1998 28445 2002 28452
rect 1997 28431 2002 28445
rect 1987 28430 2021 28431
rect 1429 28428 2021 28430
rect 1429 28427 1443 28428
rect 1446 28403 1453 28428
rect 1446 28358 1450 28403
rect 1470 28358 1474 28428
rect 1494 28358 1498 28428
rect 1518 28358 1522 28428
rect 1542 28358 1546 28428
rect 1566 28358 1570 28428
rect 1590 28358 1594 28428
rect 1614 28358 1618 28428
rect 1638 28358 1642 28428
rect 1662 28358 1666 28428
rect 1686 28358 1690 28428
rect 1710 28358 1714 28428
rect 1734 28358 1738 28428
rect 1758 28358 1762 28428
rect 1782 28358 1786 28428
rect 1806 28358 1810 28428
rect 1830 28358 1834 28428
rect 1854 28358 1858 28428
rect 1878 28359 1882 28428
rect 1867 28358 1901 28359
rect -2393 28356 1901 28358
rect -2371 28262 -2366 28356
rect -2348 28262 -2343 28356
rect -2325 28322 -2320 28356
rect -2317 28354 -2309 28356
rect -2084 28343 -2083 28356
rect -2084 28342 -2054 28343
rect -2325 28314 -2317 28322
rect -2325 28262 -2320 28314
rect -2317 28306 -2309 28314
rect -2117 28305 -2095 28315
rect -2045 28312 -2037 28326
rect -2309 28266 -2301 28276
rect -2087 28272 -2076 28280
rect -2017 28276 -2015 28283
rect -2317 28262 -2309 28266
rect -2092 28264 -2087 28272
rect -2092 28262 -2077 28263
rect -2000 28262 -1992 28356
rect -1663 28354 -1655 28356
rect -1969 28305 -1929 28317
rect -1671 28314 -1663 28322
rect -1663 28306 -1655 28314
rect -1655 28266 -1647 28276
rect -1928 28262 -1924 28263
rect -1854 28262 -1680 28263
rect -1663 28262 -1655 28266
rect -1642 28262 -1637 28356
rect -1619 28262 -1614 28356
rect -1530 28262 -1526 28356
rect -1506 28262 -1502 28356
rect -1482 28262 -1478 28356
rect -1458 28262 -1454 28356
rect -1434 28262 -1430 28356
rect -1410 28262 -1406 28356
rect -1386 28262 -1382 28356
rect -1362 28262 -1358 28356
rect -1338 28262 -1334 28356
rect -1314 28262 -1310 28356
rect -1290 28262 -1286 28356
rect -1266 28262 -1262 28356
rect -1242 28262 -1238 28356
rect -1218 28262 -1214 28356
rect -1194 28262 -1190 28356
rect -1170 28262 -1166 28356
rect -1146 28262 -1142 28356
rect -1122 28262 -1118 28356
rect -1098 28262 -1094 28356
rect -1074 28262 -1070 28356
rect -1050 28262 -1046 28356
rect -1026 28262 -1022 28356
rect -1002 28262 -998 28356
rect -978 28262 -974 28356
rect -954 28262 -950 28356
rect -930 28262 -926 28356
rect -906 28262 -902 28356
rect -882 28262 -878 28356
rect -858 28262 -854 28356
rect -834 28262 -830 28356
rect -810 28262 -806 28356
rect -786 28262 -782 28356
rect -762 28262 -758 28356
rect -738 28262 -734 28356
rect -714 28262 -710 28356
rect -690 28355 -686 28356
rect -690 28334 -683 28355
rect -666 28334 -662 28356
rect -642 28334 -638 28356
rect -618 28334 -614 28356
rect -594 28334 -590 28356
rect -570 28334 -566 28356
rect -546 28334 -542 28356
rect -522 28334 -518 28356
rect -498 28334 -494 28356
rect -474 28334 -470 28356
rect -450 28334 -446 28356
rect -426 28334 -422 28356
rect -402 28334 -398 28356
rect -378 28334 -374 28356
rect -354 28334 -350 28356
rect -330 28334 -326 28356
rect -306 28334 -302 28356
rect -282 28335 -278 28356
rect -293 28334 -259 28335
rect -707 28332 -259 28334
rect -707 28331 -693 28332
rect -690 28307 -683 28332
rect -690 28262 -686 28307
rect -666 28262 -662 28332
rect -642 28262 -638 28332
rect -618 28262 -614 28332
rect -594 28262 -590 28332
rect -570 28262 -566 28332
rect -546 28262 -542 28332
rect -522 28262 -518 28332
rect -498 28262 -494 28332
rect -474 28262 -470 28332
rect -450 28262 -446 28332
rect -426 28262 -422 28332
rect -402 28262 -398 28332
rect -378 28262 -374 28332
rect -354 28262 -350 28332
rect -330 28262 -326 28332
rect -306 28262 -302 28332
rect -293 28325 -288 28332
rect -282 28325 -278 28332
rect -283 28311 -278 28325
rect -293 28301 -288 28311
rect -282 28301 -278 28311
rect -283 28287 -278 28301
rect -293 28277 -288 28287
rect -283 28263 -278 28277
rect -282 28262 -278 28263
rect -258 28262 -254 28356
rect -234 28262 -230 28356
rect -210 28262 -206 28356
rect -186 28262 -182 28356
rect -162 28263 -158 28356
rect -173 28262 -139 28263
rect -2393 28260 -139 28262
rect -2371 28238 -2366 28260
rect -2348 28238 -2343 28260
rect -2325 28238 -2320 28260
rect -2092 28255 -2037 28260
rect -2021 28255 -1969 28260
rect -1921 28255 -1913 28260
rect -1854 28256 -1680 28260
rect -2100 28253 -2092 28254
rect -2309 28238 -2301 28248
rect -2100 28247 -2087 28253
rect -2051 28240 -2026 28242
rect -2062 28238 -2012 28240
rect -2000 28238 -1992 28255
rect -1969 28247 -1921 28254
rect -1969 28238 -1964 28247
rect -1864 28238 -1796 28239
rect -1655 28238 -1647 28248
rect -1642 28238 -1637 28260
rect -1619 28238 -1614 28260
rect -1530 28238 -1526 28260
rect -1506 28238 -1502 28260
rect -1482 28238 -1478 28260
rect -1458 28238 -1454 28260
rect -1434 28238 -1430 28260
rect -1410 28238 -1406 28260
rect -1386 28238 -1382 28260
rect -1362 28238 -1358 28260
rect -1338 28238 -1334 28260
rect -1314 28238 -1310 28260
rect -1290 28238 -1286 28260
rect -1266 28238 -1262 28260
rect -1242 28238 -1238 28260
rect -1218 28238 -1214 28260
rect -1194 28238 -1190 28260
rect -1170 28238 -1166 28260
rect -1146 28238 -1142 28260
rect -1122 28238 -1118 28260
rect -1098 28238 -1094 28260
rect -1074 28238 -1070 28260
rect -1050 28238 -1046 28260
rect -1026 28238 -1022 28260
rect -1002 28239 -998 28260
rect -1013 28238 -979 28239
rect -2393 28236 -979 28238
rect -2371 28190 -2366 28236
rect -2348 28190 -2343 28236
rect -2325 28190 -2320 28236
rect -2317 28232 -2309 28236
rect -2105 28229 -2092 28232
rect -2092 28206 -2062 28208
rect -2094 28202 -2062 28206
rect -2000 28190 -1992 28236
rect -1663 28232 -1655 28236
rect -1969 28229 -1921 28232
rect -1854 28206 -1806 28208
rect -1854 28202 -1680 28206
rect -1642 28190 -1637 28236
rect -1619 28190 -1614 28236
rect -1530 28190 -1526 28236
rect -1506 28190 -1502 28236
rect -1482 28190 -1478 28236
rect -1458 28190 -1454 28236
rect -1434 28190 -1430 28236
rect -1410 28190 -1406 28236
rect -1386 28190 -1382 28236
rect -1362 28190 -1358 28236
rect -1338 28190 -1334 28236
rect -1314 28190 -1310 28236
rect -1290 28190 -1286 28236
rect -1266 28190 -1262 28236
rect -1242 28190 -1238 28236
rect -1218 28190 -1214 28236
rect -1194 28190 -1190 28236
rect -1170 28190 -1166 28236
rect -1146 28190 -1142 28236
rect -1122 28190 -1118 28236
rect -1098 28190 -1094 28236
rect -1074 28190 -1070 28236
rect -1050 28190 -1046 28236
rect -1026 28190 -1022 28236
rect -1013 28229 -1008 28236
rect -1002 28229 -998 28236
rect -1003 28215 -998 28229
rect -1002 28190 -998 28215
rect -978 28190 -974 28260
rect -954 28190 -950 28260
rect -930 28190 -926 28260
rect -906 28190 -902 28260
rect -882 28190 -878 28260
rect -858 28190 -854 28260
rect -834 28190 -830 28260
rect -810 28190 -806 28260
rect -786 28190 -782 28260
rect -762 28190 -758 28260
rect -738 28190 -734 28260
rect -714 28190 -710 28260
rect -690 28190 -686 28260
rect -666 28190 -662 28260
rect -642 28190 -638 28260
rect -618 28190 -614 28260
rect -594 28190 -590 28260
rect -570 28190 -566 28260
rect -546 28190 -542 28260
rect -522 28190 -518 28260
rect -498 28190 -494 28260
rect -474 28190 -470 28260
rect -450 28190 -446 28260
rect -426 28190 -422 28260
rect -402 28190 -398 28260
rect -378 28190 -374 28260
rect -354 28190 -350 28260
rect -330 28190 -326 28260
rect -306 28190 -302 28260
rect -282 28190 -278 28260
rect -258 28259 -254 28260
rect -2393 28188 -261 28190
rect -2371 28166 -2366 28188
rect -2348 28166 -2343 28188
rect -2325 28166 -2320 28188
rect -2072 28186 -2036 28187
rect -2072 28180 -2054 28186
rect -2309 28172 -2301 28180
rect -2317 28166 -2309 28172
rect -2092 28171 -2062 28176
rect -2000 28167 -1992 28188
rect -1938 28187 -1906 28188
rect -1920 28186 -1906 28187
rect -1806 28180 -1680 28186
rect -1854 28171 -1806 28176
rect -1655 28172 -1647 28180
rect -1982 28167 -1966 28168
rect -2000 28166 -1966 28167
rect -1846 28166 -1806 28169
rect -1663 28166 -1655 28172
rect -1642 28166 -1637 28188
rect -1619 28166 -1614 28188
rect -1530 28166 -1526 28188
rect -1506 28166 -1502 28188
rect -1482 28166 -1478 28188
rect -1458 28166 -1454 28188
rect -1434 28166 -1430 28188
rect -1410 28166 -1406 28188
rect -1386 28166 -1382 28188
rect -1362 28166 -1358 28188
rect -1338 28166 -1334 28188
rect -1314 28166 -1310 28188
rect -1290 28166 -1286 28188
rect -1266 28166 -1262 28188
rect -1242 28166 -1238 28188
rect -1218 28166 -1214 28188
rect -1194 28166 -1190 28188
rect -1170 28166 -1166 28188
rect -1146 28166 -1142 28188
rect -1122 28166 -1118 28188
rect -1098 28166 -1094 28188
rect -1074 28166 -1070 28188
rect -1050 28166 -1046 28188
rect -1026 28166 -1022 28188
rect -1002 28166 -998 28188
rect -978 28166 -974 28188
rect -954 28166 -950 28188
rect -930 28166 -926 28188
rect -906 28166 -902 28188
rect -882 28166 -878 28188
rect -858 28166 -854 28188
rect -834 28166 -830 28188
rect -810 28166 -806 28188
rect -786 28166 -782 28188
rect -762 28166 -758 28188
rect -738 28166 -734 28188
rect -714 28166 -710 28188
rect -690 28166 -686 28188
rect -666 28166 -662 28188
rect -642 28166 -638 28188
rect -618 28166 -614 28188
rect -594 28166 -590 28188
rect -570 28166 -566 28188
rect -546 28166 -542 28188
rect -522 28166 -518 28188
rect -498 28166 -494 28188
rect -474 28166 -470 28188
rect -450 28166 -446 28188
rect -426 28166 -422 28188
rect -402 28166 -398 28188
rect -378 28166 -374 28188
rect -354 28166 -350 28188
rect -330 28166 -326 28188
rect -306 28166 -302 28188
rect -282 28166 -278 28188
rect -275 28187 -261 28188
rect -258 28187 -251 28259
rect -258 28166 -254 28187
rect -234 28166 -230 28260
rect -210 28166 -206 28260
rect -186 28166 -182 28260
rect -173 28253 -168 28260
rect -162 28253 -158 28260
rect -163 28239 -158 28253
rect -162 28166 -158 28239
rect -138 28187 -134 28356
rect -2393 28164 -141 28166
rect -2371 28142 -2366 28164
rect -2348 28142 -2343 28164
rect -2325 28142 -2320 28164
rect -2000 28162 -1966 28164
rect -2309 28144 -2301 28152
rect -2062 28151 -2054 28158
rect -2092 28144 -2084 28151
rect -2062 28144 -2026 28146
rect -2317 28142 -2309 28144
rect -2062 28142 -2012 28144
rect -2000 28142 -1992 28162
rect -1982 28161 -1966 28162
rect -1846 28160 -1806 28164
rect -1846 28153 -1798 28158
rect -1806 28151 -1798 28153
rect -1854 28149 -1846 28151
rect -1854 28144 -1806 28149
rect -1655 28144 -1647 28152
rect -1864 28142 -1796 28143
rect -1663 28142 -1655 28144
rect -1642 28142 -1637 28164
rect -1619 28142 -1614 28164
rect -1530 28142 -1526 28164
rect -1506 28142 -1502 28164
rect -1482 28142 -1478 28164
rect -1458 28142 -1454 28164
rect -1434 28142 -1430 28164
rect -1410 28142 -1406 28164
rect -1386 28142 -1382 28164
rect -1362 28142 -1358 28164
rect -1338 28142 -1334 28164
rect -1314 28142 -1310 28164
rect -1290 28142 -1286 28164
rect -1266 28142 -1262 28164
rect -1242 28142 -1238 28164
rect -1218 28142 -1214 28164
rect -1194 28142 -1190 28164
rect -1170 28142 -1166 28164
rect -1146 28142 -1142 28164
rect -1122 28142 -1118 28164
rect -1098 28142 -1094 28164
rect -1074 28142 -1070 28164
rect -1050 28142 -1046 28164
rect -1026 28142 -1022 28164
rect -1002 28142 -998 28164
rect -978 28163 -974 28164
rect -2393 28140 -981 28142
rect -2371 28094 -2366 28140
rect -2348 28094 -2343 28140
rect -2325 28094 -2320 28140
rect -2317 28136 -2309 28140
rect -2062 28136 -2054 28140
rect -2154 28132 -2138 28134
rect -2057 28132 -2054 28136
rect -2292 28126 -2054 28132
rect -2052 28126 -2044 28136
rect -2092 28110 -2062 28112
rect -2094 28106 -2062 28110
rect -2000 28094 -1992 28140
rect -1846 28133 -1806 28140
rect -1663 28136 -1655 28140
rect -1846 28126 -1680 28132
rect -1854 28110 -1806 28112
rect -1854 28106 -1680 28110
rect -1642 28094 -1637 28140
rect -1619 28094 -1614 28140
rect -1530 28094 -1526 28140
rect -1506 28094 -1502 28140
rect -1482 28094 -1478 28140
rect -1469 28109 -1464 28119
rect -1458 28109 -1454 28140
rect -1459 28095 -1454 28109
rect -1469 28094 -1435 28095
rect -2393 28092 -1435 28094
rect -2371 28070 -2366 28092
rect -2348 28070 -2343 28092
rect -2325 28070 -2320 28092
rect -2072 28090 -2036 28091
rect -2072 28084 -2054 28090
rect -2309 28076 -2301 28084
rect -2317 28070 -2309 28076
rect -2092 28075 -2062 28080
rect -2000 28071 -1992 28092
rect -1938 28091 -1906 28092
rect -1920 28090 -1906 28091
rect -1806 28084 -1680 28090
rect -1854 28075 -1806 28080
rect -1655 28076 -1647 28084
rect -1982 28071 -1966 28072
rect -2000 28070 -1966 28071
rect -1846 28070 -1806 28073
rect -1663 28070 -1655 28076
rect -1642 28070 -1637 28092
rect -1619 28070 -1614 28092
rect -1530 28070 -1526 28092
rect -1506 28070 -1502 28092
rect -1482 28070 -1478 28092
rect -1469 28085 -1464 28092
rect -1459 28071 -1454 28085
rect -1458 28070 -1454 28071
rect -1434 28070 -1430 28140
rect -1410 28070 -1406 28140
rect -1386 28070 -1382 28140
rect -1362 28070 -1358 28140
rect -1338 28070 -1334 28140
rect -1314 28070 -1310 28140
rect -1290 28070 -1286 28140
rect -1266 28070 -1262 28140
rect -1242 28070 -1238 28140
rect -1218 28070 -1214 28140
rect -1194 28070 -1190 28140
rect -1170 28070 -1166 28140
rect -1146 28070 -1142 28140
rect -1122 28070 -1118 28140
rect -1098 28070 -1094 28140
rect -1074 28070 -1070 28140
rect -1050 28070 -1046 28140
rect -1026 28070 -1022 28140
rect -1002 28070 -998 28140
rect -995 28139 -981 28140
rect -978 28139 -971 28163
rect -978 28070 -974 28139
rect -954 28070 -950 28164
rect -930 28071 -926 28164
rect -941 28070 -907 28071
rect -2393 28068 -907 28070
rect -2371 28046 -2366 28068
rect -2348 28046 -2343 28068
rect -2325 28046 -2320 28068
rect -2000 28066 -1966 28068
rect -2309 28048 -2301 28056
rect -2062 28055 -2054 28062
rect -2092 28048 -2084 28055
rect -2062 28048 -2026 28050
rect -2317 28046 -2309 28048
rect -2062 28046 -2012 28048
rect -2000 28046 -1992 28066
rect -1982 28065 -1966 28066
rect -1846 28064 -1806 28068
rect -1846 28057 -1798 28062
rect -1806 28055 -1798 28057
rect -1854 28053 -1846 28055
rect -1854 28048 -1806 28053
rect -1655 28048 -1647 28056
rect -1864 28046 -1796 28047
rect -1663 28046 -1655 28048
rect -1642 28046 -1637 28068
rect -1619 28046 -1614 28068
rect -1530 28046 -1526 28068
rect -1506 28046 -1502 28068
rect -1482 28046 -1478 28068
rect -1458 28046 -1454 28068
rect -1434 28046 -1430 28068
rect -1410 28046 -1406 28068
rect -1386 28046 -1382 28068
rect -1362 28046 -1358 28068
rect -1338 28046 -1334 28068
rect -1314 28046 -1310 28068
rect -1290 28046 -1286 28068
rect -1266 28046 -1262 28068
rect -1242 28046 -1238 28068
rect -1218 28046 -1214 28068
rect -1194 28046 -1190 28068
rect -1170 28046 -1166 28068
rect -1146 28046 -1142 28068
rect -1122 28046 -1118 28068
rect -1098 28046 -1094 28068
rect -1074 28046 -1070 28068
rect -1050 28046 -1046 28068
rect -1026 28046 -1022 28068
rect -1002 28046 -998 28068
rect -978 28046 -974 28068
rect -954 28046 -950 28068
rect -941 28061 -936 28068
rect -930 28061 -926 28068
rect -931 28047 -926 28061
rect -930 28046 -926 28047
rect -906 28046 -902 28164
rect -882 28046 -878 28164
rect -858 28046 -854 28164
rect -834 28046 -830 28164
rect -810 28046 -806 28164
rect -786 28046 -782 28164
rect -762 28046 -758 28164
rect -738 28046 -734 28164
rect -714 28046 -710 28164
rect -690 28046 -686 28164
rect -666 28046 -662 28164
rect -642 28046 -638 28164
rect -618 28046 -614 28164
rect -594 28046 -590 28164
rect -570 28046 -566 28164
rect -546 28046 -542 28164
rect -522 28046 -518 28164
rect -498 28046 -494 28164
rect -474 28046 -470 28164
rect -450 28046 -446 28164
rect -426 28046 -422 28164
rect -402 28046 -398 28164
rect -378 28046 -374 28164
rect -354 28046 -350 28164
rect -330 28046 -326 28164
rect -306 28046 -302 28164
rect -282 28046 -278 28164
rect -258 28046 -254 28164
rect -234 28046 -230 28164
rect -210 28046 -206 28164
rect -186 28046 -182 28164
rect -162 28046 -158 28164
rect -155 28163 -141 28164
rect -138 28163 -131 28187
rect -138 28046 -134 28163
rect -114 28046 -110 28356
rect -90 28046 -86 28356
rect -66 28046 -62 28356
rect -42 28046 -38 28356
rect -18 28046 -14 28356
rect 6 28046 10 28356
rect 30 28046 34 28356
rect 54 28046 58 28356
rect 78 28046 82 28356
rect 102 28046 106 28356
rect 126 28046 130 28356
rect 150 28046 154 28356
rect 174 28046 178 28356
rect 198 28046 202 28356
rect 222 28046 226 28356
rect 246 28046 250 28356
rect 270 28046 274 28356
rect 294 28046 298 28356
rect 318 28046 322 28356
rect 342 28046 346 28356
rect 366 28046 370 28356
rect 390 28046 394 28356
rect 414 28046 418 28356
rect 438 28046 442 28356
rect 462 28046 466 28356
rect 486 28046 490 28356
rect 510 28046 514 28356
rect 534 28046 538 28356
rect 558 28046 562 28356
rect 582 28046 586 28356
rect 606 28046 610 28356
rect 630 28046 634 28356
rect 654 28046 658 28356
rect 678 28046 682 28356
rect 702 28046 706 28356
rect 726 28046 730 28356
rect 750 28046 754 28356
rect 774 28046 778 28356
rect 798 28046 802 28356
rect 822 28046 826 28356
rect 846 28046 850 28356
rect 870 28215 874 28356
rect 859 28214 893 28215
rect 894 28214 898 28356
rect 918 28214 922 28356
rect 942 28214 946 28356
rect 966 28214 970 28356
rect 990 28214 994 28356
rect 1014 28214 1018 28356
rect 1038 28214 1042 28356
rect 1062 28214 1066 28356
rect 1086 28214 1090 28356
rect 1110 28214 1114 28356
rect 1134 28214 1138 28356
rect 1158 28214 1162 28356
rect 1182 28214 1186 28356
rect 1206 28214 1210 28356
rect 1230 28214 1234 28356
rect 1254 28214 1258 28356
rect 1278 28214 1282 28356
rect 1302 28214 1306 28356
rect 1326 28214 1330 28356
rect 1350 28214 1354 28356
rect 1374 28214 1378 28356
rect 1398 28214 1402 28356
rect 1422 28214 1426 28356
rect 1446 28214 1450 28356
rect 1470 28214 1474 28356
rect 1494 28214 1498 28356
rect 1518 28214 1522 28356
rect 1542 28214 1546 28356
rect 1566 28214 1570 28356
rect 1590 28214 1594 28356
rect 1614 28214 1618 28356
rect 1638 28214 1642 28356
rect 1662 28214 1666 28356
rect 1686 28214 1690 28356
rect 1710 28214 1714 28356
rect 1734 28214 1738 28356
rect 1758 28214 1762 28356
rect 1782 28214 1786 28356
rect 1806 28214 1810 28356
rect 1830 28214 1834 28356
rect 1854 28214 1858 28356
rect 1867 28349 1872 28356
rect 1878 28349 1882 28356
rect 1877 28335 1882 28349
rect 1878 28214 1882 28335
rect 1902 28283 1906 28428
rect 1902 28259 1909 28283
rect 1902 28214 1906 28259
rect 1926 28214 1930 28428
rect 1950 28214 1954 28428
rect 1974 28214 1978 28428
rect 1987 28421 1992 28428
rect 1997 28407 2002 28421
rect 1998 28214 2002 28407
rect 2011 28301 2016 28311
rect 2021 28287 2026 28301
rect 2022 28214 2026 28287
rect 2035 28214 2043 28215
rect 859 28212 2043 28214
rect 859 28205 864 28212
rect 870 28205 874 28212
rect 869 28191 874 28205
rect 859 28181 864 28191
rect 869 28167 874 28181
rect 870 28046 874 28167
rect 894 28139 898 28212
rect 894 28118 901 28139
rect 918 28118 922 28212
rect 942 28118 946 28212
rect 966 28118 970 28212
rect 990 28118 994 28212
rect 1014 28118 1018 28212
rect 1038 28118 1042 28212
rect 1062 28118 1066 28212
rect 1086 28118 1090 28212
rect 1110 28118 1114 28212
rect 1134 28118 1138 28212
rect 1158 28118 1162 28212
rect 1182 28118 1186 28212
rect 1206 28118 1210 28212
rect 1230 28118 1234 28212
rect 1254 28118 1258 28212
rect 1278 28118 1282 28212
rect 1302 28118 1306 28212
rect 1326 28118 1330 28212
rect 1350 28118 1354 28212
rect 1374 28118 1378 28212
rect 1398 28118 1402 28212
rect 1422 28118 1426 28212
rect 1446 28118 1450 28212
rect 1470 28118 1474 28212
rect 1494 28118 1498 28212
rect 1518 28118 1522 28212
rect 1542 28118 1546 28212
rect 1566 28118 1570 28212
rect 1590 28118 1594 28212
rect 1614 28118 1618 28212
rect 1638 28118 1642 28212
rect 1662 28118 1666 28212
rect 1686 28118 1690 28212
rect 1710 28118 1714 28212
rect 1734 28118 1738 28212
rect 1758 28118 1762 28212
rect 1782 28118 1786 28212
rect 1806 28118 1810 28212
rect 1830 28118 1834 28212
rect 1854 28118 1858 28212
rect 1878 28118 1882 28212
rect 1902 28118 1906 28212
rect 1926 28118 1930 28212
rect 1950 28118 1954 28212
rect 1974 28118 1978 28212
rect 1998 28118 2002 28212
rect 2011 28133 2016 28143
rect 2022 28133 2026 28212
rect 2029 28211 2043 28212
rect 2035 28205 2040 28211
rect 2045 28191 2050 28205
rect 2035 28157 2040 28167
rect 2046 28157 2050 28191
rect 2045 28143 2050 28157
rect 2021 28119 2026 28133
rect 2011 28118 2045 28119
rect 877 28116 2045 28118
rect 877 28115 891 28116
rect 894 28091 901 28116
rect 894 28046 898 28091
rect 918 28046 922 28116
rect 942 28046 946 28116
rect 966 28046 970 28116
rect 990 28046 994 28116
rect 1014 28046 1018 28116
rect 1038 28046 1042 28116
rect 1062 28046 1066 28116
rect 1086 28046 1090 28116
rect 1110 28046 1114 28116
rect 1134 28047 1138 28116
rect 1123 28046 1157 28047
rect -2393 28044 1157 28046
rect -2371 27998 -2366 28044
rect -2348 27998 -2343 28044
rect -2325 27998 -2320 28044
rect -2317 28040 -2309 28044
rect -2062 28040 -2054 28044
rect -2154 28036 -2138 28038
rect -2057 28036 -2054 28040
rect -2292 28030 -2054 28036
rect -2052 28030 -2044 28040
rect -2092 28014 -2062 28016
rect -2094 28010 -2062 28014
rect -2000 27998 -1992 28044
rect -1846 28037 -1806 28044
rect -1663 28040 -1655 28044
rect -1846 28030 -1680 28036
rect -1854 28014 -1806 28016
rect -1854 28010 -1680 28014
rect -1642 27998 -1637 28044
rect -1619 27998 -1614 28044
rect -1530 27998 -1526 28044
rect -1506 27998 -1502 28044
rect -1482 27998 -1478 28044
rect -1458 27998 -1454 28044
rect -1434 28043 -1430 28044
rect -2393 27996 -1437 27998
rect -2371 27974 -2366 27996
rect -2348 27974 -2343 27996
rect -2325 27974 -2320 27996
rect -2072 27994 -2036 27995
rect -2072 27988 -2054 27994
rect -2309 27980 -2301 27988
rect -2317 27974 -2309 27980
rect -2092 27979 -2062 27984
rect -2000 27975 -1992 27996
rect -1938 27995 -1906 27996
rect -1920 27994 -1906 27995
rect -1806 27988 -1680 27994
rect -1854 27979 -1806 27984
rect -1655 27980 -1647 27988
rect -1982 27975 -1966 27976
rect -2000 27974 -1966 27975
rect -1846 27974 -1806 27977
rect -1663 27974 -1655 27980
rect -1642 27974 -1637 27996
rect -1619 27974 -1614 27996
rect -1530 27974 -1526 27996
rect -1506 27974 -1502 27996
rect -1482 27974 -1478 27996
rect -1458 27974 -1454 27996
rect -1451 27995 -1437 27996
rect -1434 27995 -1427 28043
rect -1434 27974 -1430 27995
rect -1410 27974 -1406 28044
rect -1386 27974 -1382 28044
rect -1362 27974 -1358 28044
rect -1338 27974 -1334 28044
rect -1314 27975 -1310 28044
rect -1325 27974 -1291 27975
rect -2393 27972 -1291 27974
rect -2371 27950 -2366 27972
rect -2348 27950 -2343 27972
rect -2325 27950 -2320 27972
rect -2000 27970 -1966 27972
rect -2309 27952 -2301 27960
rect -2062 27959 -2054 27966
rect -2092 27952 -2084 27959
rect -2062 27952 -2026 27954
rect -2317 27950 -2309 27952
rect -2062 27950 -2012 27952
rect -2000 27950 -1992 27970
rect -1982 27969 -1966 27970
rect -1846 27968 -1806 27972
rect -1846 27961 -1798 27966
rect -1806 27959 -1798 27961
rect -1854 27957 -1846 27959
rect -1854 27952 -1806 27957
rect -1655 27952 -1647 27960
rect -1864 27950 -1796 27951
rect -1663 27950 -1655 27952
rect -1642 27950 -1637 27972
rect -1619 27950 -1614 27972
rect -1530 27950 -1526 27972
rect -1506 27950 -1502 27972
rect -1482 27950 -1478 27972
rect -1458 27950 -1454 27972
rect -1434 27950 -1430 27972
rect -1410 27950 -1406 27972
rect -1386 27950 -1382 27972
rect -1362 27950 -1358 27972
rect -1338 27950 -1334 27972
rect -1325 27965 -1320 27972
rect -1314 27965 -1310 27972
rect -1315 27951 -1310 27965
rect -1314 27950 -1310 27951
rect -1290 27950 -1286 28044
rect -1266 27950 -1262 28044
rect -1242 27950 -1238 28044
rect -1218 27950 -1214 28044
rect -1194 27950 -1190 28044
rect -1170 27951 -1166 28044
rect -1181 27950 -1147 27951
rect -2393 27948 -1147 27950
rect -2371 27902 -2366 27948
rect -2348 27902 -2343 27948
rect -2325 27902 -2320 27948
rect -2317 27944 -2309 27948
rect -2062 27944 -2054 27948
rect -2154 27940 -2138 27942
rect -2057 27940 -2054 27944
rect -2292 27934 -2054 27940
rect -2052 27934 -2044 27944
rect -2092 27918 -2062 27920
rect -2094 27914 -2062 27918
rect -2000 27902 -1992 27948
rect -1846 27941 -1806 27948
rect -1663 27944 -1655 27948
rect -1846 27934 -1680 27940
rect -1854 27918 -1806 27920
rect -1854 27914 -1680 27918
rect -1979 27902 -1945 27904
rect -1642 27902 -1637 27948
rect -1619 27902 -1614 27948
rect -1530 27902 -1526 27948
rect -1517 27917 -1512 27927
rect -1506 27917 -1502 27948
rect -1507 27903 -1502 27917
rect -1517 27902 -1483 27903
rect -2393 27900 -1483 27902
rect -2371 27854 -2366 27900
rect -2348 27854 -2343 27900
rect -2325 27854 -2320 27900
rect -2080 27899 -1906 27900
rect -2080 27898 -2036 27899
rect -2080 27892 -2054 27898
rect -2309 27884 -2301 27890
rect -2317 27874 -2309 27884
rect -2070 27883 -2040 27890
rect -2054 27875 -2040 27878
rect -2000 27873 -1992 27899
rect -1920 27898 -1906 27899
rect -1850 27892 -1846 27900
rect -1840 27892 -1792 27900
rect -1969 27880 -1966 27889
rect -1850 27885 -1802 27890
rect -1906 27883 -1802 27885
rect -1655 27884 -1647 27890
rect -1906 27882 -1850 27883
rect -1846 27875 -1802 27881
rect -1663 27874 -1655 27884
rect -1860 27873 -1798 27874
rect -2078 27866 -2070 27873
rect -2309 27856 -2301 27862
rect -2317 27854 -2309 27856
rect -2154 27854 -2145 27864
rect -2044 27863 -2040 27868
rect -2028 27866 -1945 27873
rect -1929 27866 -1794 27873
rect -2070 27856 -2040 27863
rect -2044 27854 -2028 27856
rect -2000 27854 -1992 27866
rect -1860 27865 -1798 27866
rect -1850 27856 -1802 27863
rect -1655 27856 -1647 27862
rect -1978 27854 -1942 27855
rect -1663 27854 -1655 27856
rect -1642 27854 -1637 27900
rect -1619 27854 -1614 27900
rect -1530 27854 -1526 27900
rect -1517 27893 -1512 27900
rect -1507 27879 -1502 27893
rect -1506 27854 -1502 27879
rect -1482 27854 -1478 27948
rect -1458 27854 -1454 27948
rect -1434 27854 -1430 27948
rect -1410 27854 -1406 27948
rect -1386 27854 -1382 27948
rect -1362 27854 -1358 27948
rect -1338 27854 -1334 27948
rect -1314 27854 -1310 27948
rect -1290 27899 -1286 27948
rect -1290 27875 -1283 27899
rect -1290 27854 -1286 27875
rect -1266 27854 -1262 27948
rect -1242 27854 -1238 27948
rect -1218 27854 -1214 27948
rect -1194 27854 -1190 27948
rect -1181 27941 -1176 27948
rect -1170 27941 -1166 27948
rect -1171 27927 -1166 27941
rect -1170 27854 -1166 27927
rect -1146 27875 -1142 28044
rect -2393 27852 -1149 27854
rect -2371 27758 -2366 27852
rect -2348 27758 -2343 27852
rect -2325 27814 -2320 27852
rect -2317 27846 -2309 27852
rect -2145 27848 -2138 27852
rect -2070 27848 -2054 27852
rect -2078 27839 -2054 27846
rect -2062 27814 -2032 27815
rect -2000 27814 -1992 27852
rect -1846 27848 -1802 27852
rect -1846 27838 -1792 27847
rect -1663 27846 -1655 27852
rect -1942 27816 -1937 27828
rect -1850 27825 -1822 27826
rect -1850 27821 -1802 27825
rect -2325 27806 -2317 27814
rect -2062 27812 -1961 27814
rect -2325 27786 -2320 27806
rect -2317 27798 -2309 27806
rect -2062 27799 -2040 27810
rect -2032 27805 -1961 27812
rect -1947 27806 -1942 27814
rect -1842 27812 -1794 27815
rect -2070 27794 -2022 27798
rect -2325 27770 -2317 27786
rect -2325 27758 -2320 27770
rect -2309 27758 -2301 27770
rect -2000 27758 -1992 27805
rect -1942 27804 -1937 27806
rect -1932 27796 -1927 27804
rect -1912 27801 -1896 27807
rect -1842 27799 -1802 27810
rect -1671 27806 -1663 27814
rect -1663 27798 -1655 27806
rect -1850 27794 -1680 27798
rect -1671 27770 -1663 27786
rect -1655 27758 -1647 27770
rect -1642 27758 -1637 27852
rect -1619 27758 -1614 27852
rect -1530 27758 -1526 27852
rect -1506 27758 -1502 27852
rect -1482 27851 -1478 27852
rect -1482 27830 -1475 27851
rect -1458 27830 -1454 27852
rect -1434 27830 -1430 27852
rect -1410 27830 -1406 27852
rect -1386 27830 -1382 27852
rect -1362 27830 -1358 27852
rect -1338 27830 -1334 27852
rect -1314 27830 -1310 27852
rect -1290 27830 -1286 27852
rect -1266 27830 -1262 27852
rect -1242 27830 -1238 27852
rect -1218 27830 -1214 27852
rect -1194 27830 -1190 27852
rect -1170 27830 -1166 27852
rect -1163 27851 -1149 27852
rect -1146 27851 -1139 27875
rect -1146 27830 -1142 27851
rect -1122 27830 -1118 28044
rect -1098 27830 -1094 28044
rect -1074 27830 -1070 28044
rect -1050 27830 -1046 28044
rect -1026 27830 -1022 28044
rect -1002 27830 -998 28044
rect -978 27830 -974 28044
rect -954 27830 -950 28044
rect -930 27830 -926 28044
rect -906 27995 -902 28044
rect -906 27971 -899 27995
rect -906 27830 -902 27971
rect -882 27830 -878 28044
rect -858 27831 -854 28044
rect -869 27830 -835 27831
rect -1499 27828 -835 27830
rect -1499 27827 -1485 27828
rect -1482 27803 -1475 27828
rect -1482 27758 -1478 27803
rect -1458 27758 -1454 27828
rect -1434 27758 -1430 27828
rect -1410 27758 -1406 27828
rect -1386 27758 -1382 27828
rect -1362 27758 -1358 27828
rect -1338 27758 -1334 27828
rect -1314 27758 -1310 27828
rect -1301 27773 -1296 27783
rect -1290 27773 -1286 27828
rect -1291 27759 -1286 27773
rect -1301 27758 -1267 27759
rect -2393 27756 -1267 27758
rect -2371 27662 -2366 27756
rect -2348 27662 -2343 27756
rect -2325 27754 -2320 27756
rect -2317 27754 -2309 27756
rect -2325 27742 -2317 27754
rect -2061 27743 -2046 27744
rect -2325 27726 -2320 27742
rect -2309 27730 -2301 27742
rect -2070 27736 -2046 27743
rect -2000 27738 -1992 27756
rect -1974 27754 -1960 27756
rect -1663 27754 -1655 27756
rect -1960 27753 -1944 27754
rect -1980 27738 -1932 27743
rect -1671 27742 -1663 27754
rect -2061 27734 -2046 27736
rect -2032 27736 -1932 27738
rect -2032 27734 -1980 27736
rect -2317 27726 -2309 27730
rect -2062 27728 -2061 27734
rect -2062 27726 -2051 27727
rect -2325 27714 -2317 27726
rect -2062 27719 -2032 27726
rect -2062 27718 -2051 27719
rect -2325 27694 -2320 27714
rect -2325 27686 -2317 27694
rect -2325 27666 -2320 27686
rect -2317 27678 -2309 27686
rect -2325 27662 -2317 27666
rect -2000 27662 -1992 27734
rect -1655 27730 -1647 27742
rect -1990 27718 -1924 27727
rect -1904 27725 -1874 27727
rect -1842 27718 -1680 27727
rect -1663 27726 -1655 27730
rect -1671 27714 -1663 27726
rect -1671 27686 -1663 27694
rect -1663 27678 -1655 27686
rect -1671 27662 -1663 27666
rect -1642 27662 -1637 27756
rect -1619 27662 -1614 27756
rect -1530 27662 -1526 27756
rect -1506 27662 -1502 27756
rect -1482 27662 -1478 27756
rect -1458 27662 -1454 27756
rect -1434 27662 -1430 27756
rect -1410 27662 -1406 27756
rect -1386 27662 -1382 27756
rect -1362 27662 -1358 27756
rect -1338 27662 -1334 27756
rect -1314 27662 -1310 27756
rect -1301 27749 -1296 27756
rect -1291 27735 -1286 27749
rect -1290 27662 -1286 27735
rect -1266 27707 -1262 27828
rect -2393 27660 -1969 27662
rect -1955 27660 -1269 27662
rect -2371 27614 -2366 27660
rect -2348 27614 -2343 27660
rect -2325 27650 -2317 27660
rect -2080 27658 -1969 27660
rect -2080 27652 -2053 27658
rect -2325 27634 -2320 27650
rect -2309 27638 -2301 27650
rect -2070 27643 -2040 27650
rect -2000 27642 -1992 27658
rect -1972 27654 -1969 27658
rect -1972 27652 -1955 27654
rect -1955 27642 -1850 27651
rect -1671 27650 -1663 27660
rect -2317 27634 -2309 27638
rect -2070 27635 -2053 27641
rect -2027 27640 -1992 27642
rect -1969 27640 -1955 27641
rect -2325 27622 -2317 27634
rect -2292 27625 -2053 27634
rect -2325 27614 -2320 27622
rect -2309 27614 -2301 27622
rect -2000 27614 -1992 27640
rect -1655 27638 -1647 27650
rect -1663 27634 -1655 27638
rect -1972 27626 -1924 27633
rect -1945 27625 -1929 27626
rect -1860 27625 -1680 27634
rect -1671 27622 -1663 27634
rect -1978 27614 -1942 27615
rect -1655 27614 -1647 27622
rect -1642 27614 -1637 27660
rect -1619 27614 -1614 27660
rect -1530 27614 -1526 27660
rect -1506 27614 -1502 27660
rect -1482 27614 -1478 27660
rect -1458 27614 -1454 27660
rect -1434 27614 -1430 27660
rect -1410 27614 -1406 27660
rect -1386 27614 -1382 27660
rect -1362 27614 -1358 27660
rect -1338 27614 -1334 27660
rect -1314 27614 -1310 27660
rect -1290 27614 -1286 27660
rect -1283 27659 -1269 27660
rect -1266 27659 -1259 27707
rect -1266 27614 -1262 27659
rect -1242 27614 -1238 27828
rect -1218 27614 -1214 27828
rect -1194 27614 -1190 27828
rect -1170 27614 -1166 27828
rect -1146 27614 -1142 27828
rect -1122 27614 -1118 27828
rect -1098 27614 -1094 27828
rect -1074 27614 -1070 27828
rect -1050 27614 -1046 27828
rect -1026 27614 -1022 27828
rect -1002 27614 -998 27828
rect -978 27614 -974 27828
rect -954 27614 -950 27828
rect -930 27614 -926 27828
rect -906 27614 -902 27828
rect -882 27614 -878 27828
rect -869 27821 -864 27828
rect -858 27821 -854 27828
rect -859 27807 -854 27821
rect -858 27614 -854 27807
rect -834 27755 -830 28044
rect -834 27731 -827 27755
rect -834 27614 -830 27731
rect -810 27614 -806 28044
rect -786 27614 -782 28044
rect -773 27701 -768 27711
rect -762 27701 -758 28044
rect -763 27687 -758 27701
rect -762 27614 -758 27687
rect -738 27635 -734 28044
rect -2393 27612 -741 27614
rect -2371 27518 -2366 27612
rect -2348 27518 -2343 27612
rect -2325 27606 -2320 27612
rect -2309 27610 -2301 27612
rect -2317 27606 -2309 27610
rect -2325 27594 -2317 27606
rect -2325 27574 -2320 27594
rect -2062 27574 -2032 27575
rect -2000 27574 -1992 27612
rect -1655 27610 -1647 27612
rect -1663 27606 -1655 27610
rect -1671 27594 -1663 27606
rect -1942 27576 -1937 27588
rect -1850 27585 -1822 27586
rect -1850 27581 -1802 27585
rect -2325 27566 -2317 27574
rect -2062 27572 -1961 27574
rect -2325 27546 -2320 27566
rect -2317 27558 -2309 27566
rect -2062 27559 -2040 27570
rect -2032 27565 -1961 27572
rect -1947 27566 -1942 27574
rect -1842 27572 -1794 27575
rect -2070 27554 -2022 27558
rect -2325 27532 -2317 27546
rect -2072 27538 -2032 27539
rect -2102 27532 -2032 27538
rect -2325 27518 -2320 27532
rect -2317 27530 -2309 27532
rect -2309 27518 -2301 27530
rect -2070 27523 -2062 27528
rect -2000 27518 -1992 27565
rect -1942 27564 -1937 27566
rect -1932 27556 -1927 27564
rect -1912 27561 -1896 27567
rect -1842 27559 -1802 27570
rect -1671 27566 -1663 27574
rect -1663 27558 -1655 27566
rect -1850 27554 -1680 27558
rect -1924 27540 -1921 27542
rect -1806 27532 -1680 27538
rect -1671 27532 -1663 27546
rect -1663 27530 -1655 27532
rect -1854 27523 -1806 27528
rect -1974 27518 -1964 27519
rect -1960 27518 -1944 27520
rect -1842 27518 -1806 27521
rect -1655 27518 -1647 27530
rect -1642 27518 -1637 27612
rect -1619 27518 -1614 27612
rect -1530 27518 -1526 27612
rect -1506 27518 -1502 27612
rect -1482 27518 -1478 27612
rect -1458 27518 -1454 27612
rect -1434 27518 -1430 27612
rect -1410 27518 -1406 27612
rect -1386 27518 -1382 27612
rect -1362 27518 -1358 27612
rect -1338 27518 -1334 27612
rect -1314 27518 -1310 27612
rect -1290 27518 -1286 27612
rect -1266 27518 -1262 27612
rect -1242 27518 -1238 27612
rect -1218 27518 -1214 27612
rect -1194 27518 -1190 27612
rect -1170 27518 -1166 27612
rect -1146 27518 -1142 27612
rect -1122 27518 -1118 27612
rect -1098 27518 -1094 27612
rect -1074 27518 -1070 27612
rect -1050 27518 -1046 27612
rect -1026 27518 -1022 27612
rect -1002 27518 -998 27612
rect -978 27518 -974 27612
rect -954 27518 -950 27612
rect -930 27518 -926 27612
rect -906 27518 -902 27612
rect -882 27518 -878 27612
rect -858 27518 -854 27612
rect -834 27518 -830 27612
rect -810 27518 -806 27612
rect -786 27518 -782 27612
rect -762 27518 -758 27612
rect -755 27611 -741 27612
rect -738 27611 -731 27635
rect -738 27518 -734 27611
rect -714 27518 -710 28044
rect -690 27518 -686 28044
rect -666 27518 -662 28044
rect -642 27518 -638 28044
rect -618 27518 -614 28044
rect -594 27518 -590 28044
rect -570 27518 -566 28044
rect -546 27518 -542 28044
rect -522 27518 -518 28044
rect -498 27518 -494 28044
rect -474 27518 -470 28044
rect -450 27518 -446 28044
rect -426 27518 -422 28044
rect -402 27518 -398 28044
rect -378 27518 -374 28044
rect -354 27518 -350 28044
rect -330 27518 -326 28044
rect -306 27518 -302 28044
rect -282 27518 -278 28044
rect -258 27518 -254 28044
rect -234 27518 -230 28044
rect -210 27518 -206 28044
rect -186 27518 -182 28044
rect -162 27518 -158 28044
rect -138 27518 -134 28044
rect -114 27518 -110 28044
rect -90 27518 -86 28044
rect -66 27518 -62 28044
rect -53 27845 -48 27855
rect -42 27845 -38 28044
rect -43 27831 -38 27845
rect -42 27518 -38 27831
rect -18 27779 -14 28044
rect -18 27755 -11 27779
rect -18 27518 -14 27755
rect 6 27518 10 28044
rect 30 27518 34 28044
rect 54 27518 58 28044
rect 78 27518 82 28044
rect 102 27518 106 28044
rect 126 27518 130 28044
rect 150 27518 154 28044
rect 174 27518 178 28044
rect 198 27518 202 28044
rect 222 27518 226 28044
rect 246 27518 250 28044
rect 270 27518 274 28044
rect 283 27605 288 27615
rect 294 27605 298 28044
rect 293 27591 298 27605
rect 294 27518 298 27591
rect 318 27539 322 28044
rect 307 27518 315 27519
rect -2393 27516 315 27518
rect -2371 27494 -2366 27516
rect -2348 27494 -2343 27516
rect -2325 27504 -2317 27516
rect -2325 27494 -2320 27504
rect -2317 27502 -2309 27504
rect -2062 27503 -2032 27510
rect -2309 27494 -2301 27502
rect -2070 27496 -2062 27503
rect -2000 27498 -1992 27516
rect -1974 27514 -1944 27516
rect -1960 27513 -1944 27514
rect -1842 27512 -1806 27516
rect -1842 27505 -1798 27510
rect -1806 27503 -1798 27505
rect -1671 27504 -1663 27516
rect -1854 27501 -1842 27503
rect -1663 27502 -1655 27504
rect -2062 27494 -2036 27496
rect -2393 27492 -2036 27494
rect -2032 27494 -2012 27496
rect -2004 27494 -1974 27498
rect -1854 27496 -1806 27501
rect -1864 27494 -1796 27495
rect -1655 27494 -1647 27502
rect -1642 27494 -1637 27516
rect -1619 27494 -1614 27516
rect -1530 27494 -1526 27516
rect -1506 27494 -1502 27516
rect -1482 27494 -1478 27516
rect -1458 27494 -1454 27516
rect -1434 27494 -1430 27516
rect -1410 27494 -1406 27516
rect -1386 27494 -1382 27516
rect -1362 27494 -1358 27516
rect -1338 27494 -1334 27516
rect -1314 27494 -1310 27516
rect -1290 27494 -1286 27516
rect -1266 27494 -1262 27516
rect -1242 27494 -1238 27516
rect -1218 27494 -1214 27516
rect -1194 27494 -1190 27516
rect -1170 27495 -1166 27516
rect -1181 27494 -1147 27495
rect -2032 27492 -1147 27494
rect -2371 27422 -2366 27492
rect -2348 27422 -2343 27492
rect -2325 27488 -2320 27492
rect -2309 27490 -2301 27492
rect -2317 27488 -2309 27490
rect -2325 27476 -2317 27488
rect -2052 27486 -2036 27488
rect -2052 27484 -2032 27486
rect -2062 27478 -2032 27484
rect -2325 27422 -2320 27476
rect -2317 27474 -2309 27476
rect -2092 27462 -2062 27464
rect -2094 27458 -2062 27462
rect -2309 27428 -2301 27434
rect -2317 27422 -2309 27428
rect -2000 27422 -1992 27492
rect -1904 27485 -1874 27492
rect -1842 27485 -1806 27492
rect -1655 27490 -1647 27492
rect -1663 27488 -1655 27490
rect -1842 27478 -1680 27484
rect -1671 27476 -1663 27488
rect -1663 27474 -1655 27476
rect -1854 27462 -1806 27464
rect -1854 27458 -1680 27462
rect -1655 27428 -1647 27434
rect -1663 27422 -1655 27428
rect -1642 27422 -1637 27492
rect -1619 27422 -1614 27492
rect -1530 27422 -1526 27492
rect -1506 27422 -1502 27492
rect -1482 27422 -1478 27492
rect -1458 27422 -1454 27492
rect -1434 27422 -1430 27492
rect -1410 27422 -1406 27492
rect -1386 27422 -1382 27492
rect -1362 27422 -1358 27492
rect -1338 27422 -1334 27492
rect -1314 27422 -1310 27492
rect -1290 27422 -1286 27492
rect -1266 27422 -1262 27492
rect -1242 27422 -1238 27492
rect -1218 27422 -1214 27492
rect -1194 27422 -1190 27492
rect -1181 27485 -1176 27492
rect -1170 27485 -1166 27492
rect -1171 27471 -1166 27485
rect -1170 27422 -1166 27471
rect -1146 27422 -1142 27516
rect -1122 27422 -1118 27516
rect -1098 27422 -1094 27516
rect -1074 27422 -1070 27516
rect -1050 27422 -1046 27516
rect -1026 27422 -1022 27516
rect -1002 27422 -998 27516
rect -978 27422 -974 27516
rect -954 27422 -950 27516
rect -930 27422 -926 27516
rect -906 27422 -902 27516
rect -882 27422 -878 27516
rect -858 27422 -854 27516
rect -834 27422 -830 27516
rect -810 27422 -806 27516
rect -786 27422 -782 27516
rect -762 27422 -758 27516
rect -738 27422 -734 27516
rect -714 27422 -710 27516
rect -690 27422 -686 27516
rect -666 27422 -662 27516
rect -642 27422 -638 27516
rect -618 27422 -614 27516
rect -594 27422 -590 27516
rect -570 27422 -566 27516
rect -546 27422 -542 27516
rect -522 27422 -518 27516
rect -498 27422 -494 27516
rect -474 27422 -470 27516
rect -450 27422 -446 27516
rect -426 27422 -422 27516
rect -402 27422 -398 27516
rect -378 27422 -374 27516
rect -354 27422 -350 27516
rect -330 27422 -326 27516
rect -306 27422 -302 27516
rect -282 27422 -278 27516
rect -258 27422 -254 27516
rect -234 27422 -230 27516
rect -210 27422 -206 27516
rect -186 27422 -182 27516
rect -162 27422 -158 27516
rect -138 27422 -134 27516
rect -114 27422 -110 27516
rect -90 27422 -86 27516
rect -66 27422 -62 27516
rect -42 27422 -38 27516
rect -18 27422 -14 27516
rect 6 27422 10 27516
rect 30 27422 34 27516
rect 54 27422 58 27516
rect 78 27422 82 27516
rect 102 27422 106 27516
rect 126 27422 130 27516
rect 150 27447 154 27516
rect 139 27446 173 27447
rect 174 27446 178 27516
rect 198 27446 202 27516
rect 222 27446 226 27516
rect 246 27446 250 27516
rect 270 27446 274 27516
rect 294 27446 298 27516
rect 301 27515 315 27516
rect 318 27515 325 27539
rect 307 27509 312 27515
rect 318 27509 322 27515
rect 317 27495 322 27509
rect 318 27446 322 27495
rect 342 27446 346 28044
rect 366 27446 370 28044
rect 390 27446 394 28044
rect 414 27446 418 28044
rect 438 27446 442 28044
rect 462 27446 466 28044
rect 486 27446 490 28044
rect 510 27687 514 28044
rect 499 27686 533 27687
rect 534 27686 538 28044
rect 558 27686 562 28044
rect 582 27686 586 28044
rect 606 27686 610 28044
rect 630 27686 634 28044
rect 654 27686 658 28044
rect 678 27686 682 28044
rect 702 27686 706 28044
rect 726 27686 730 28044
rect 750 27686 754 28044
rect 774 27686 778 28044
rect 798 27686 802 28044
rect 822 27686 826 28044
rect 846 27686 850 28044
rect 870 27686 874 28044
rect 894 27686 898 28044
rect 918 28023 922 28044
rect 907 28022 941 28023
rect 942 28022 946 28044
rect 966 28022 970 28044
rect 990 28022 994 28044
rect 1014 28022 1018 28044
rect 1038 28022 1042 28044
rect 1062 28022 1066 28044
rect 1086 28022 1090 28044
rect 1110 28022 1114 28044
rect 1123 28037 1128 28044
rect 1134 28037 1138 28044
rect 1133 28023 1138 28037
rect 1134 28022 1138 28023
rect 1158 28022 1162 28116
rect 1182 28022 1186 28116
rect 1206 28022 1210 28116
rect 1230 28022 1234 28116
rect 1254 28022 1258 28116
rect 1278 28022 1282 28116
rect 1302 28022 1306 28116
rect 1326 28022 1330 28116
rect 1350 28022 1354 28116
rect 1374 28022 1378 28116
rect 1398 28022 1402 28116
rect 1422 28022 1426 28116
rect 1446 28022 1450 28116
rect 1470 28022 1474 28116
rect 1494 28022 1498 28116
rect 1518 28022 1522 28116
rect 1542 28022 1546 28116
rect 1566 28022 1570 28116
rect 1590 28022 1594 28116
rect 1614 28022 1618 28116
rect 1638 28022 1642 28116
rect 1662 28022 1666 28116
rect 1686 28022 1690 28116
rect 1710 28022 1714 28116
rect 1734 28022 1738 28116
rect 1758 28022 1762 28116
rect 1782 28022 1786 28116
rect 1806 28022 1810 28116
rect 1830 28022 1834 28116
rect 1854 28022 1858 28116
rect 1878 28022 1882 28116
rect 1902 28022 1906 28116
rect 1926 28022 1930 28116
rect 1950 28022 1954 28116
rect 1974 28022 1978 28116
rect 1998 28022 2002 28116
rect 2011 28109 2016 28116
rect 2021 28095 2026 28109
rect 2022 28022 2026 28095
rect 2035 28022 2043 28023
rect 907 28020 2043 28022
rect 907 28013 912 28020
rect 918 28013 922 28020
rect 917 27999 922 28013
rect 907 27989 912 27999
rect 917 27975 922 27989
rect 918 27686 922 27975
rect 942 27947 946 28020
rect 942 27926 949 27947
rect 966 27926 970 28020
rect 990 27926 994 28020
rect 1014 27926 1018 28020
rect 1038 27926 1042 28020
rect 1062 27926 1066 28020
rect 1086 27926 1090 28020
rect 1110 27926 1114 28020
rect 1134 27926 1138 28020
rect 1158 27971 1162 28020
rect 1158 27947 1165 27971
rect 1158 27926 1162 27947
rect 1182 27926 1186 28020
rect 1206 27926 1210 28020
rect 1230 27926 1234 28020
rect 1254 27926 1258 28020
rect 1278 27926 1282 28020
rect 1302 27926 1306 28020
rect 1326 27926 1330 28020
rect 1350 27926 1354 28020
rect 1374 27926 1378 28020
rect 1398 27926 1402 28020
rect 1422 27926 1426 28020
rect 1446 27926 1450 28020
rect 1470 27926 1474 28020
rect 1494 27926 1498 28020
rect 1518 27926 1522 28020
rect 1542 27926 1546 28020
rect 1566 27926 1570 28020
rect 1590 27926 1594 28020
rect 1614 27926 1618 28020
rect 1638 27926 1642 28020
rect 1662 27926 1666 28020
rect 1686 27926 1690 28020
rect 1710 27926 1714 28020
rect 1734 27926 1738 28020
rect 1758 27926 1762 28020
rect 1782 27926 1786 28020
rect 1806 27926 1810 28020
rect 1830 27926 1834 28020
rect 1854 27926 1858 28020
rect 1878 27926 1882 28020
rect 1902 27926 1906 28020
rect 1926 27926 1930 28020
rect 1950 27926 1954 28020
rect 1974 27926 1978 28020
rect 1998 27926 2002 28020
rect 2022 27926 2026 28020
rect 2029 28019 2043 28020
rect 2035 28013 2040 28019
rect 2045 27999 2050 28013
rect 2046 27926 2050 27999
rect 2059 27926 2067 27927
rect 925 27924 2067 27926
rect 925 27923 939 27924
rect 942 27899 949 27924
rect 942 27686 946 27899
rect 966 27686 970 27924
rect 990 27686 994 27924
rect 1014 27686 1018 27924
rect 1038 27686 1042 27924
rect 1062 27686 1066 27924
rect 1086 27686 1090 27924
rect 1110 27686 1114 27924
rect 1134 27686 1138 27924
rect 1158 27686 1162 27924
rect 1182 27686 1186 27924
rect 1206 27686 1210 27924
rect 1230 27686 1234 27924
rect 1254 27686 1258 27924
rect 1278 27686 1282 27924
rect 1302 27686 1306 27924
rect 1326 27686 1330 27924
rect 1350 27686 1354 27924
rect 1374 27686 1378 27924
rect 1398 27686 1402 27924
rect 1422 27686 1426 27924
rect 1446 27686 1450 27924
rect 1470 27686 1474 27924
rect 1494 27686 1498 27924
rect 1518 27686 1522 27924
rect 1542 27686 1546 27924
rect 1566 27686 1570 27924
rect 1590 27686 1594 27924
rect 1614 27686 1618 27924
rect 1638 27686 1642 27924
rect 1662 27686 1666 27924
rect 1686 27686 1690 27924
rect 1710 27686 1714 27924
rect 1734 27686 1738 27924
rect 1758 27686 1762 27924
rect 1782 27686 1786 27924
rect 1806 27686 1810 27924
rect 1830 27686 1834 27924
rect 1854 27686 1858 27924
rect 1878 27686 1882 27924
rect 1902 27686 1906 27924
rect 1926 27686 1930 27924
rect 1950 27686 1954 27924
rect 1974 27686 1978 27924
rect 1998 27686 2002 27924
rect 2022 27686 2026 27924
rect 2046 27686 2050 27924
rect 2053 27923 2067 27924
rect 2059 27917 2064 27923
rect 2069 27903 2074 27917
rect 2070 27686 2074 27903
rect 2083 27773 2088 27783
rect 2093 27759 2098 27773
rect 2094 27686 2098 27759
rect 2107 27686 2115 27687
rect 499 27684 2115 27686
rect 499 27677 504 27684
rect 510 27677 514 27684
rect 509 27663 514 27677
rect 499 27653 504 27663
rect 509 27639 514 27653
rect 510 27446 514 27639
rect 534 27611 538 27684
rect 534 27590 541 27611
rect 558 27590 562 27684
rect 582 27590 586 27684
rect 606 27590 610 27684
rect 630 27590 634 27684
rect 654 27590 658 27684
rect 678 27590 682 27684
rect 702 27590 706 27684
rect 726 27590 730 27684
rect 750 27590 754 27684
rect 774 27590 778 27684
rect 798 27590 802 27684
rect 822 27590 826 27684
rect 846 27590 850 27684
rect 870 27590 874 27684
rect 894 27590 898 27684
rect 918 27590 922 27684
rect 942 27590 946 27684
rect 966 27590 970 27684
rect 990 27590 994 27684
rect 1014 27590 1018 27684
rect 1038 27590 1042 27684
rect 1062 27590 1066 27684
rect 1086 27590 1090 27684
rect 1110 27590 1114 27684
rect 1134 27591 1138 27684
rect 1123 27590 1157 27591
rect 517 27588 1157 27590
rect 517 27587 531 27588
rect 534 27563 541 27588
rect 534 27446 538 27563
rect 558 27446 562 27588
rect 582 27446 586 27588
rect 606 27446 610 27588
rect 630 27446 634 27588
rect 654 27446 658 27588
rect 678 27446 682 27588
rect 702 27446 706 27588
rect 726 27446 730 27588
rect 739 27557 744 27567
rect 750 27557 754 27588
rect 749 27543 754 27557
rect 739 27533 744 27543
rect 749 27519 754 27533
rect 750 27446 754 27519
rect 774 27491 778 27588
rect 139 27444 771 27446
rect 139 27437 144 27444
rect 150 27437 154 27444
rect 149 27423 154 27437
rect 139 27422 173 27423
rect -2393 27420 173 27422
rect -2371 27326 -2366 27420
rect -2348 27326 -2343 27420
rect -2325 27358 -2320 27420
rect -2317 27418 -2309 27420
rect -2000 27419 -1966 27420
rect -2000 27418 -1982 27419
rect -1663 27418 -1655 27420
rect -2028 27410 -2018 27412
rect -2309 27400 -2301 27406
rect -2091 27400 -2061 27407
rect -2317 27390 -2309 27400
rect -2044 27398 -2028 27400
rect -2026 27398 -2014 27410
rect -2084 27392 -2061 27398
rect -2044 27396 -2014 27398
rect -2292 27382 -2054 27391
rect -2325 27350 -2317 27358
rect -2325 27330 -2320 27350
rect -2317 27342 -2309 27350
rect -2325 27326 -2317 27330
rect -2000 27326 -1992 27418
rect -1982 27417 -1966 27418
rect -1980 27400 -1932 27407
rect -1655 27400 -1647 27406
rect -1846 27382 -1680 27391
rect -1663 27390 -1655 27400
rect -1671 27350 -1663 27358
rect -1663 27342 -1655 27350
rect -1926 27326 -1892 27329
rect -1671 27326 -1663 27330
rect -1642 27326 -1637 27420
rect -1619 27326 -1614 27420
rect -1530 27326 -1526 27420
rect -1506 27326 -1502 27420
rect -1482 27326 -1478 27420
rect -1458 27326 -1454 27420
rect -1434 27326 -1430 27420
rect -1410 27326 -1406 27420
rect -1386 27326 -1382 27420
rect -1362 27326 -1358 27420
rect -1338 27326 -1334 27420
rect -1314 27326 -1310 27420
rect -1290 27326 -1286 27420
rect -1266 27326 -1262 27420
rect -1242 27326 -1238 27420
rect -1218 27326 -1214 27420
rect -1194 27326 -1190 27420
rect -1170 27326 -1166 27420
rect -1146 27419 -1142 27420
rect -1146 27395 -1139 27419
rect -1146 27326 -1142 27395
rect -1122 27326 -1118 27420
rect -1098 27326 -1094 27420
rect -1074 27326 -1070 27420
rect -1050 27326 -1046 27420
rect -1026 27326 -1022 27420
rect -1002 27326 -998 27420
rect -978 27326 -974 27420
rect -954 27326 -950 27420
rect -930 27326 -926 27420
rect -906 27326 -902 27420
rect -882 27326 -878 27420
rect -858 27326 -854 27420
rect -834 27326 -830 27420
rect -810 27326 -806 27420
rect -786 27326 -782 27420
rect -762 27326 -758 27420
rect -738 27326 -734 27420
rect -714 27326 -710 27420
rect -690 27326 -686 27420
rect -666 27326 -662 27420
rect -642 27326 -638 27420
rect -618 27326 -614 27420
rect -594 27326 -590 27420
rect -570 27326 -566 27420
rect -546 27326 -542 27420
rect -522 27326 -518 27420
rect -498 27326 -494 27420
rect -474 27326 -470 27420
rect -450 27326 -446 27420
rect -426 27326 -422 27420
rect -402 27326 -398 27420
rect -378 27326 -374 27420
rect -365 27341 -360 27351
rect -354 27341 -350 27420
rect -355 27327 -350 27341
rect -365 27326 -331 27327
rect -2393 27324 -331 27326
rect -2371 27278 -2366 27324
rect -2348 27278 -2343 27324
rect -2325 27318 -2317 27324
rect -2053 27322 -1972 27324
rect -2325 27302 -2320 27318
rect -2317 27314 -2309 27318
rect -2069 27314 -2068 27315
rect -2309 27302 -2301 27314
rect -2069 27307 -2038 27314
rect -2069 27305 -2068 27307
rect -2000 27306 -1992 27322
rect -1926 27319 -1924 27324
rect -1916 27316 -1914 27319
rect -1671 27318 -1663 27324
rect -1982 27306 -1916 27315
rect -1663 27314 -1655 27318
rect -2325 27290 -2317 27302
rect -2068 27299 -2053 27305
rect -2027 27304 -1992 27306
rect -2076 27290 -2053 27297
rect -2011 27296 -2002 27304
rect -2000 27296 -1992 27304
rect -1655 27302 -1647 27314
rect -2003 27294 -1992 27296
rect -2325 27278 -2320 27290
rect -2317 27286 -2309 27290
rect -2309 27278 -2301 27286
rect -2015 27282 -2003 27294
rect -2000 27278 -1992 27294
rect -1972 27290 -1924 27297
rect -1862 27289 -1680 27298
rect -1671 27290 -1663 27302
rect -1663 27286 -1655 27290
rect -1976 27278 -1940 27279
rect -1655 27278 -1647 27286
rect -1642 27278 -1637 27324
rect -1619 27278 -1614 27324
rect -1530 27278 -1526 27324
rect -1506 27278 -1502 27324
rect -1482 27278 -1478 27324
rect -1458 27278 -1454 27324
rect -1434 27278 -1430 27324
rect -1410 27278 -1406 27324
rect -1386 27279 -1382 27324
rect -1397 27278 -1363 27279
rect -2393 27276 -1363 27278
rect -2371 27206 -2366 27276
rect -2348 27206 -2343 27276
rect -2325 27274 -2320 27276
rect -2309 27274 -2301 27276
rect -2325 27262 -2317 27274
rect -2325 27242 -2320 27262
rect -2317 27258 -2309 27262
rect -2325 27234 -2317 27242
rect -2060 27236 -2030 27239
rect -2325 27206 -2320 27234
rect -2317 27226 -2309 27234
rect -2060 27223 -2038 27234
rect -2033 27227 -2030 27236
rect -2028 27232 -2027 27236
rect -2068 27218 -2038 27221
rect -2000 27206 -1992 27276
rect -1655 27274 -1647 27276
rect -1671 27262 -1663 27274
rect -1663 27258 -1655 27262
rect -1912 27251 -1884 27253
rect -1852 27245 -1804 27249
rect -1844 27236 -1796 27239
rect -1671 27234 -1663 27242
rect -1844 27223 -1804 27234
rect -1663 27226 -1655 27234
rect -1852 27218 -1680 27222
rect -1642 27206 -1637 27276
rect -1619 27206 -1614 27276
rect -1530 27206 -1526 27276
rect -1506 27206 -1502 27276
rect -1482 27206 -1478 27276
rect -1458 27206 -1454 27276
rect -1434 27206 -1430 27276
rect -1410 27206 -1406 27276
rect -1397 27269 -1392 27276
rect -1386 27269 -1382 27276
rect -1387 27255 -1382 27269
rect -1386 27206 -1382 27255
rect -1362 27206 -1358 27324
rect -1338 27206 -1334 27324
rect -1314 27206 -1310 27324
rect -1290 27206 -1286 27324
rect -1266 27206 -1262 27324
rect -1242 27206 -1238 27324
rect -1218 27206 -1214 27324
rect -1194 27206 -1190 27324
rect -1170 27206 -1166 27324
rect -1146 27206 -1142 27324
rect -1122 27206 -1118 27324
rect -1098 27206 -1094 27324
rect -1074 27206 -1070 27324
rect -1050 27206 -1046 27324
rect -1026 27206 -1022 27324
rect -1002 27206 -998 27324
rect -978 27206 -974 27324
rect -954 27206 -950 27324
rect -930 27231 -926 27324
rect -941 27230 -907 27231
rect -906 27230 -902 27324
rect -882 27230 -878 27324
rect -858 27230 -854 27324
rect -834 27230 -830 27324
rect -810 27230 -806 27324
rect -786 27230 -782 27324
rect -762 27230 -758 27324
rect -738 27230 -734 27324
rect -714 27230 -710 27324
rect -690 27230 -686 27324
rect -666 27230 -662 27324
rect -642 27230 -638 27324
rect -618 27230 -614 27324
rect -594 27230 -590 27324
rect -570 27230 -566 27324
rect -546 27230 -542 27324
rect -522 27230 -518 27324
rect -498 27230 -494 27324
rect -474 27230 -470 27324
rect -450 27230 -446 27324
rect -426 27230 -422 27324
rect -402 27230 -398 27324
rect -378 27230 -374 27324
rect -365 27317 -360 27324
rect -355 27303 -350 27317
rect -354 27230 -350 27303
rect -330 27275 -326 27420
rect -330 27254 -323 27275
rect -306 27254 -302 27420
rect -282 27254 -278 27420
rect -258 27254 -254 27420
rect -234 27254 -230 27420
rect -210 27254 -206 27420
rect -186 27254 -182 27420
rect -162 27254 -158 27420
rect -138 27254 -134 27420
rect -114 27254 -110 27420
rect -90 27254 -86 27420
rect -66 27254 -62 27420
rect -42 27254 -38 27420
rect -18 27254 -14 27420
rect 6 27254 10 27420
rect 30 27254 34 27420
rect 54 27254 58 27420
rect 78 27254 82 27420
rect 102 27254 106 27420
rect 126 27254 130 27420
rect 139 27413 144 27420
rect 149 27399 154 27413
rect 150 27254 154 27399
rect 174 27371 178 27444
rect 174 27350 181 27371
rect 198 27350 202 27444
rect 222 27350 226 27444
rect 246 27350 250 27444
rect 270 27350 274 27444
rect 294 27350 298 27444
rect 318 27350 322 27444
rect 342 27443 346 27444
rect 342 27419 349 27443
rect 342 27350 346 27419
rect 366 27350 370 27444
rect 390 27350 394 27444
rect 414 27350 418 27444
rect 438 27350 442 27444
rect 462 27350 466 27444
rect 486 27350 490 27444
rect 510 27350 514 27444
rect 534 27350 538 27444
rect 558 27350 562 27444
rect 582 27350 586 27444
rect 606 27350 610 27444
rect 630 27350 634 27444
rect 654 27350 658 27444
rect 678 27350 682 27444
rect 702 27350 706 27444
rect 726 27350 730 27444
rect 750 27350 754 27444
rect 757 27443 771 27444
rect 774 27443 781 27491
rect 774 27350 778 27443
rect 798 27350 802 27588
rect 822 27350 826 27588
rect 846 27350 850 27588
rect 870 27350 874 27588
rect 894 27350 898 27588
rect 918 27350 922 27588
rect 942 27350 946 27588
rect 966 27350 970 27588
rect 990 27350 994 27588
rect 1014 27350 1018 27588
rect 1038 27350 1042 27588
rect 1062 27350 1066 27588
rect 1086 27350 1090 27588
rect 1110 27350 1114 27588
rect 1123 27581 1128 27588
rect 1134 27581 1138 27588
rect 1133 27567 1138 27581
rect 1134 27350 1138 27567
rect 1158 27515 1162 27684
rect 1158 27491 1165 27515
rect 1158 27350 1162 27491
rect 1182 27350 1186 27684
rect 1206 27350 1210 27684
rect 1230 27350 1234 27684
rect 1254 27350 1258 27684
rect 1278 27350 1282 27684
rect 1302 27350 1306 27684
rect 1326 27350 1330 27684
rect 1350 27350 1354 27684
rect 1374 27350 1378 27684
rect 1398 27350 1402 27684
rect 1422 27350 1426 27684
rect 1446 27350 1450 27684
rect 1470 27350 1474 27684
rect 1494 27350 1498 27684
rect 1518 27350 1522 27684
rect 1542 27350 1546 27684
rect 1566 27350 1570 27684
rect 1590 27350 1594 27684
rect 1614 27350 1618 27684
rect 1638 27350 1642 27684
rect 1662 27350 1666 27684
rect 1686 27350 1690 27684
rect 1710 27350 1714 27684
rect 1734 27350 1738 27684
rect 1758 27350 1762 27684
rect 1782 27350 1786 27684
rect 1806 27350 1810 27684
rect 1830 27350 1834 27684
rect 1854 27350 1858 27684
rect 1878 27350 1882 27684
rect 1902 27350 1906 27684
rect 1926 27350 1930 27684
rect 1950 27350 1954 27684
rect 1974 27350 1978 27684
rect 1998 27350 2002 27684
rect 2022 27350 2026 27684
rect 2046 27350 2050 27684
rect 2070 27350 2074 27684
rect 2094 27350 2098 27684
rect 2101 27683 2115 27684
rect 2107 27677 2112 27683
rect 2117 27663 2122 27677
rect 2118 27350 2122 27663
rect 2131 27557 2136 27567
rect 2141 27543 2146 27557
rect 2142 27350 2146 27543
rect 2155 27437 2160 27447
rect 2165 27423 2170 27437
rect 2155 27365 2160 27375
rect 2166 27365 2170 27423
rect 2165 27351 2170 27365
rect 2179 27361 2187 27365
rect 2173 27351 2179 27361
rect 2155 27350 2187 27351
rect 157 27348 2187 27350
rect 157 27347 171 27348
rect 174 27323 181 27348
rect 174 27254 178 27323
rect 198 27254 202 27348
rect 222 27254 226 27348
rect 246 27254 250 27348
rect 270 27254 274 27348
rect 294 27254 298 27348
rect 318 27254 322 27348
rect 342 27254 346 27348
rect 366 27254 370 27348
rect 390 27254 394 27348
rect 414 27254 418 27348
rect 438 27255 442 27348
rect 427 27254 461 27255
rect -347 27252 461 27254
rect -347 27251 -333 27252
rect -941 27228 -333 27230
rect -941 27221 -936 27228
rect -930 27221 -926 27228
rect -931 27207 -926 27221
rect -941 27206 -907 27207
rect -2393 27204 -907 27206
rect -2371 27182 -2366 27204
rect -2348 27182 -2343 27204
rect -2325 27182 -2320 27204
rect -2309 27186 -2301 27196
rect -2068 27187 -2062 27192
rect -2317 27182 -2309 27186
rect -2060 27182 -2050 27187
rect -2000 27182 -1992 27204
rect -1806 27196 -1680 27202
rect -1854 27187 -1806 27192
rect -1655 27186 -1647 27196
rect -1972 27182 -1964 27183
rect -1958 27182 -1942 27184
rect -1844 27182 -1806 27185
rect -1663 27182 -1655 27186
rect -1642 27182 -1637 27204
rect -1619 27182 -1614 27204
rect -1530 27182 -1526 27204
rect -1506 27182 -1502 27204
rect -1482 27182 -1478 27204
rect -1458 27182 -1454 27204
rect -1434 27182 -1430 27204
rect -1410 27182 -1406 27204
rect -1386 27182 -1382 27204
rect -1362 27203 -1358 27204
rect -2393 27180 -1365 27182
rect -2371 27158 -2366 27180
rect -2348 27158 -2343 27180
rect -2325 27158 -2320 27180
rect -2060 27174 -2050 27180
rect -2309 27158 -2301 27168
rect -2060 27167 -2030 27174
rect -2000 27170 -1992 27180
rect -1972 27178 -1942 27180
rect -1958 27177 -1942 27178
rect -1844 27176 -1806 27180
rect -2068 27160 -2062 27167
rect -2062 27158 -2036 27160
rect -2393 27156 -2036 27158
rect -2030 27158 -2012 27160
rect -2004 27158 -1990 27170
rect -1844 27169 -1798 27174
rect -1806 27167 -1798 27169
rect -1854 27165 -1844 27167
rect -1854 27160 -1806 27165
rect -1864 27158 -1796 27159
rect -1655 27158 -1647 27168
rect -1642 27158 -1637 27180
rect -1619 27158 -1614 27180
rect -1530 27158 -1526 27180
rect -1506 27158 -1502 27180
rect -1482 27158 -1478 27180
rect -1458 27158 -1454 27180
rect -1434 27158 -1430 27180
rect -1410 27158 -1406 27180
rect -1386 27158 -1382 27180
rect -1379 27179 -1365 27180
rect -1362 27179 -1355 27203
rect -1362 27158 -1358 27179
rect -1338 27158 -1334 27204
rect -1314 27158 -1310 27204
rect -1290 27158 -1286 27204
rect -1266 27158 -1262 27204
rect -1242 27158 -1238 27204
rect -1218 27158 -1214 27204
rect -1194 27158 -1190 27204
rect -1170 27158 -1166 27204
rect -1146 27158 -1142 27204
rect -1122 27158 -1118 27204
rect -1098 27158 -1094 27204
rect -1074 27158 -1070 27204
rect -1050 27158 -1046 27204
rect -1026 27158 -1022 27204
rect -1002 27158 -998 27204
rect -978 27158 -974 27204
rect -954 27158 -950 27204
rect -941 27197 -936 27204
rect -931 27183 -926 27197
rect -930 27158 -926 27183
rect -906 27158 -902 27228
rect -882 27158 -878 27228
rect -858 27158 -854 27228
rect -834 27158 -830 27228
rect -810 27158 -806 27228
rect -786 27158 -782 27228
rect -762 27158 -758 27228
rect -738 27158 -734 27228
rect -714 27158 -710 27228
rect -690 27158 -686 27228
rect -666 27158 -662 27228
rect -642 27158 -638 27228
rect -618 27158 -614 27228
rect -594 27158 -590 27228
rect -570 27158 -566 27228
rect -546 27158 -542 27228
rect -522 27158 -518 27228
rect -498 27158 -494 27228
rect -474 27158 -470 27228
rect -450 27158 -446 27228
rect -426 27158 -422 27228
rect -402 27158 -398 27228
rect -378 27158 -374 27228
rect -354 27158 -350 27228
rect -347 27227 -333 27228
rect -330 27227 -323 27252
rect -330 27158 -326 27227
rect -306 27158 -302 27252
rect -282 27158 -278 27252
rect -258 27158 -254 27252
rect -234 27158 -230 27252
rect -210 27158 -206 27252
rect -186 27158 -182 27252
rect -162 27158 -158 27252
rect -138 27158 -134 27252
rect -114 27158 -110 27252
rect -90 27158 -86 27252
rect -66 27158 -62 27252
rect -42 27158 -38 27252
rect -18 27158 -14 27252
rect 6 27158 10 27252
rect 30 27158 34 27252
rect 54 27158 58 27252
rect 78 27158 82 27252
rect 102 27158 106 27252
rect 126 27158 130 27252
rect 150 27158 154 27252
rect 174 27158 178 27252
rect 198 27158 202 27252
rect 222 27158 226 27252
rect 246 27158 250 27252
rect 270 27158 274 27252
rect 294 27158 298 27252
rect 318 27158 322 27252
rect 342 27158 346 27252
rect 366 27158 370 27252
rect 390 27158 394 27252
rect 414 27158 418 27252
rect 427 27245 432 27252
rect 438 27245 442 27252
rect 437 27231 442 27245
rect 438 27158 442 27231
rect 462 27179 466 27348
rect -2030 27156 459 27158
rect -2371 27110 -2366 27156
rect -2348 27110 -2343 27156
rect -2325 27110 -2320 27156
rect -2317 27152 -2309 27156
rect -2060 27152 -2050 27156
rect -2060 27150 -2036 27152
rect -2060 27148 -2030 27150
rect -2292 27142 -2030 27148
rect -2092 27126 -2062 27128
rect -2094 27122 -2062 27126
rect -2000 27110 -1992 27156
rect -1844 27149 -1806 27156
rect -1663 27152 -1655 27156
rect -1844 27142 -1680 27148
rect -1854 27126 -1806 27128
rect -1854 27122 -1680 27126
rect -1642 27110 -1637 27156
rect -1619 27110 -1614 27156
rect -1530 27110 -1526 27156
rect -1506 27110 -1502 27156
rect -1482 27110 -1478 27156
rect -1458 27110 -1454 27156
rect -1434 27110 -1430 27156
rect -1410 27110 -1406 27156
rect -1386 27110 -1382 27156
rect -1362 27110 -1358 27156
rect -1338 27110 -1334 27156
rect -1314 27110 -1310 27156
rect -1290 27110 -1286 27156
rect -1266 27110 -1262 27156
rect -1242 27110 -1238 27156
rect -1218 27110 -1214 27156
rect -1194 27110 -1190 27156
rect -1170 27110 -1166 27156
rect -1146 27110 -1142 27156
rect -1122 27110 -1118 27156
rect -1098 27110 -1094 27156
rect -1074 27110 -1070 27156
rect -1050 27110 -1046 27156
rect -1026 27110 -1022 27156
rect -1002 27110 -998 27156
rect -978 27110 -974 27156
rect -954 27110 -950 27156
rect -930 27110 -926 27156
rect -906 27155 -902 27156
rect -2393 27108 -909 27110
rect -2371 27086 -2366 27108
rect -2348 27086 -2343 27108
rect -2325 27086 -2320 27108
rect -2072 27106 -2036 27107
rect -2072 27100 -2054 27106
rect -2309 27092 -2301 27100
rect -2317 27086 -2309 27092
rect -2092 27091 -2062 27096
rect -2000 27087 -1992 27108
rect -1938 27107 -1906 27108
rect -1920 27106 -1906 27107
rect -1806 27100 -1680 27106
rect -1854 27091 -1806 27096
rect -1655 27092 -1647 27100
rect -1982 27087 -1966 27088
rect -2000 27086 -1966 27087
rect -1846 27086 -1806 27089
rect -1663 27086 -1655 27092
rect -1642 27086 -1637 27108
rect -1619 27086 -1614 27108
rect -1530 27086 -1526 27108
rect -1506 27086 -1502 27108
rect -1482 27086 -1478 27108
rect -1458 27086 -1454 27108
rect -1434 27086 -1430 27108
rect -1410 27086 -1406 27108
rect -1386 27086 -1382 27108
rect -1362 27086 -1358 27108
rect -1338 27086 -1334 27108
rect -1314 27086 -1310 27108
rect -1290 27086 -1286 27108
rect -1266 27086 -1262 27108
rect -1242 27086 -1238 27108
rect -1218 27086 -1214 27108
rect -1194 27086 -1190 27108
rect -1170 27086 -1166 27108
rect -1146 27086 -1142 27108
rect -1122 27086 -1118 27108
rect -1098 27086 -1094 27108
rect -1074 27086 -1070 27108
rect -1050 27086 -1046 27108
rect -1026 27086 -1022 27108
rect -1002 27086 -998 27108
rect -978 27086 -974 27108
rect -954 27086 -950 27108
rect -930 27086 -926 27108
rect -923 27107 -909 27108
rect -906 27107 -899 27155
rect -906 27086 -902 27107
rect -882 27086 -878 27156
rect -858 27086 -854 27156
rect -834 27086 -830 27156
rect -810 27087 -806 27156
rect -821 27086 -787 27087
rect -786 27086 -782 27156
rect -762 27086 -758 27156
rect -738 27086 -734 27156
rect -714 27086 -710 27156
rect -690 27086 -686 27156
rect -666 27086 -662 27156
rect -642 27086 -638 27156
rect -618 27086 -614 27156
rect -594 27086 -590 27156
rect -570 27086 -566 27156
rect -546 27086 -542 27156
rect -522 27086 -518 27156
rect -498 27086 -494 27156
rect -474 27086 -470 27156
rect -450 27086 -446 27156
rect -426 27086 -422 27156
rect -402 27086 -398 27156
rect -378 27086 -374 27156
rect -354 27086 -350 27156
rect -330 27135 -326 27156
rect -341 27134 -307 27135
rect -306 27134 -302 27156
rect -282 27134 -278 27156
rect -258 27134 -254 27156
rect -234 27134 -230 27156
rect -210 27134 -206 27156
rect -186 27134 -182 27156
rect -162 27134 -158 27156
rect -138 27134 -134 27156
rect -114 27134 -110 27156
rect -90 27134 -86 27156
rect -66 27134 -62 27156
rect -42 27134 -38 27156
rect -18 27134 -14 27156
rect 6 27134 10 27156
rect 30 27134 34 27156
rect 54 27134 58 27156
rect 78 27134 82 27156
rect 102 27134 106 27156
rect 126 27134 130 27156
rect 150 27134 154 27156
rect 174 27134 178 27156
rect 198 27134 202 27156
rect 222 27134 226 27156
rect 246 27134 250 27156
rect 270 27134 274 27156
rect 294 27134 298 27156
rect 318 27134 322 27156
rect 342 27134 346 27156
rect 366 27134 370 27156
rect 390 27134 394 27156
rect 414 27134 418 27156
rect 438 27134 442 27156
rect 445 27155 459 27156
rect 462 27155 469 27179
rect 462 27134 466 27155
rect 486 27134 490 27348
rect 510 27134 514 27348
rect 534 27134 538 27348
rect 558 27134 562 27348
rect 582 27134 586 27348
rect 606 27134 610 27348
rect 630 27134 634 27348
rect 654 27134 658 27348
rect 678 27134 682 27348
rect 702 27134 706 27348
rect 726 27134 730 27348
rect 750 27134 754 27348
rect 774 27134 778 27348
rect 798 27134 802 27348
rect 822 27134 826 27348
rect 846 27134 850 27348
rect 870 27134 874 27348
rect 894 27134 898 27348
rect 918 27134 922 27348
rect 942 27134 946 27348
rect 966 27134 970 27348
rect 990 27134 994 27348
rect 1014 27134 1018 27348
rect 1038 27134 1042 27348
rect 1062 27134 1066 27348
rect 1086 27134 1090 27348
rect 1110 27134 1114 27348
rect 1123 27173 1128 27183
rect 1134 27173 1138 27348
rect 1133 27159 1138 27173
rect 1134 27134 1138 27159
rect 1147 27149 1152 27159
rect 1158 27149 1162 27348
rect 1157 27135 1162 27149
rect 1182 27134 1186 27348
rect 1206 27134 1210 27348
rect 1230 27134 1234 27348
rect 1254 27134 1258 27348
rect 1278 27134 1282 27348
rect 1302 27134 1306 27348
rect 1326 27134 1330 27348
rect 1350 27134 1354 27348
rect 1374 27134 1378 27348
rect 1398 27134 1402 27348
rect 1422 27134 1426 27348
rect 1446 27134 1450 27348
rect 1470 27134 1474 27348
rect 1494 27134 1498 27348
rect 1518 27134 1522 27348
rect 1542 27134 1546 27348
rect 1555 27293 1560 27303
rect 1566 27293 1570 27348
rect 1565 27279 1570 27293
rect 1566 27134 1570 27279
rect 1590 27227 1594 27348
rect 1590 27203 1597 27227
rect 1590 27134 1594 27203
rect 1614 27134 1618 27348
rect 1638 27134 1642 27348
rect 1662 27134 1666 27348
rect 1686 27134 1690 27348
rect 1710 27134 1714 27348
rect 1734 27134 1738 27348
rect 1758 27134 1762 27348
rect 1782 27134 1786 27348
rect 1806 27134 1810 27348
rect 1830 27134 1834 27348
rect 1854 27134 1858 27348
rect 1878 27134 1882 27348
rect 1902 27134 1906 27348
rect 1926 27134 1930 27348
rect 1950 27134 1954 27348
rect 1974 27134 1978 27348
rect 1998 27134 2002 27348
rect 2022 27134 2026 27348
rect 2046 27134 2050 27348
rect 2070 27134 2074 27348
rect 2094 27134 2098 27348
rect 2118 27134 2122 27348
rect 2142 27134 2146 27348
rect 2155 27341 2160 27348
rect 2173 27347 2187 27348
rect 2165 27327 2170 27341
rect 2166 27134 2170 27327
rect 2179 27221 2184 27231
rect 2189 27207 2194 27221
rect 2190 27134 2194 27207
rect 2203 27134 2211 27135
rect -341 27132 2211 27134
rect -341 27125 -336 27132
rect -330 27125 -326 27132
rect -331 27111 -326 27125
rect -341 27086 -307 27087
rect -2393 27084 -307 27086
rect -2371 27062 -2366 27084
rect -2348 27062 -2343 27084
rect -2325 27062 -2320 27084
rect -2000 27082 -1966 27084
rect -2309 27064 -2301 27072
rect -2062 27071 -2054 27078
rect -2092 27064 -2084 27071
rect -2062 27064 -2026 27066
rect -2317 27062 -2309 27064
rect -2062 27062 -2012 27064
rect -2000 27062 -1992 27082
rect -1982 27081 -1966 27082
rect -1846 27080 -1806 27084
rect -1846 27073 -1798 27078
rect -1806 27071 -1798 27073
rect -1854 27069 -1846 27071
rect -1854 27064 -1806 27069
rect -1655 27064 -1647 27072
rect -1864 27062 -1796 27063
rect -1663 27062 -1655 27064
rect -1642 27062 -1637 27084
rect -1619 27062 -1614 27084
rect -1530 27062 -1526 27084
rect -1506 27062 -1502 27084
rect -1482 27062 -1478 27084
rect -1458 27062 -1454 27084
rect -1434 27062 -1430 27084
rect -1410 27062 -1406 27084
rect -1386 27062 -1382 27084
rect -1362 27062 -1358 27084
rect -1338 27062 -1334 27084
rect -1314 27062 -1310 27084
rect -1290 27062 -1286 27084
rect -1266 27062 -1262 27084
rect -1242 27062 -1238 27084
rect -1218 27062 -1214 27084
rect -1194 27062 -1190 27084
rect -1170 27062 -1166 27084
rect -1146 27062 -1142 27084
rect -1122 27062 -1118 27084
rect -1098 27062 -1094 27084
rect -1074 27062 -1070 27084
rect -1050 27062 -1046 27084
rect -1026 27062 -1022 27084
rect -1002 27062 -998 27084
rect -978 27062 -974 27084
rect -954 27062 -950 27084
rect -930 27062 -926 27084
rect -906 27062 -902 27084
rect -882 27062 -878 27084
rect -858 27062 -854 27084
rect -834 27062 -830 27084
rect -821 27077 -816 27084
rect -810 27077 -806 27084
rect -811 27063 -806 27077
rect -821 27062 -787 27063
rect -2393 27060 -787 27062
rect -2371 27014 -2366 27060
rect -2348 27014 -2343 27060
rect -2325 27014 -2320 27060
rect -2317 27056 -2309 27060
rect -2062 27056 -2054 27060
rect -2154 27052 -2138 27054
rect -2057 27052 -2054 27056
rect -2292 27046 -2054 27052
rect -2052 27046 -2044 27056
rect -2092 27030 -2062 27032
rect -2094 27026 -2062 27030
rect -2000 27014 -1992 27060
rect -1846 27053 -1806 27060
rect -1663 27056 -1655 27060
rect -1846 27046 -1680 27052
rect -1854 27030 -1806 27032
rect -1854 27026 -1680 27030
rect -1642 27014 -1637 27060
rect -1619 27014 -1614 27060
rect -1530 27014 -1526 27060
rect -1506 27014 -1502 27060
rect -1482 27014 -1478 27060
rect -1458 27014 -1454 27060
rect -1434 27014 -1430 27060
rect -1410 27014 -1406 27060
rect -1386 27014 -1382 27060
rect -1362 27014 -1358 27060
rect -1338 27014 -1334 27060
rect -1314 27014 -1310 27060
rect -1290 27014 -1286 27060
rect -1266 27014 -1262 27060
rect -1242 27014 -1238 27060
rect -1218 27014 -1214 27060
rect -1194 27014 -1190 27060
rect -1170 27014 -1166 27060
rect -1146 27014 -1142 27060
rect -1122 27014 -1118 27060
rect -1098 27014 -1094 27060
rect -1074 27014 -1070 27060
rect -1050 27014 -1046 27060
rect -1026 27014 -1022 27060
rect -1002 27014 -998 27060
rect -978 27014 -974 27060
rect -954 27014 -950 27060
rect -930 27014 -926 27060
rect -906 27014 -902 27060
rect -882 27014 -878 27060
rect -858 27014 -854 27060
rect -834 27014 -830 27060
rect -821 27053 -816 27060
rect -811 27039 -806 27053
rect -810 27014 -806 27039
rect -786 27014 -782 27084
rect -762 27014 -758 27084
rect -738 27014 -734 27084
rect -714 27014 -710 27084
rect -690 27014 -686 27084
rect -666 27014 -662 27084
rect -642 27014 -638 27084
rect -618 27014 -614 27084
rect -594 27014 -590 27084
rect -570 27014 -566 27084
rect -546 27014 -542 27084
rect -522 27014 -518 27084
rect -498 27014 -494 27084
rect -474 27014 -470 27084
rect -450 27014 -446 27084
rect -426 27014 -422 27084
rect -402 27014 -398 27084
rect -378 27014 -374 27084
rect -354 27014 -350 27084
rect -341 27077 -336 27084
rect -331 27063 -326 27077
rect -330 27014 -326 27063
rect -306 27059 -302 27132
rect -306 27035 -299 27059
rect -282 27014 -278 27132
rect -258 27014 -254 27132
rect -234 27014 -230 27132
rect -210 27039 -206 27132
rect -221 27038 -187 27039
rect -186 27038 -182 27132
rect -162 27038 -158 27132
rect -138 27038 -134 27132
rect -114 27038 -110 27132
rect -90 27038 -86 27132
rect -66 27038 -62 27132
rect -42 27038 -38 27132
rect -18 27038 -14 27132
rect 6 27038 10 27132
rect 30 27038 34 27132
rect 54 27038 58 27132
rect 78 27038 82 27132
rect 102 27038 106 27132
rect 126 27038 130 27132
rect 150 27038 154 27132
rect 174 27038 178 27132
rect 198 27038 202 27132
rect 222 27038 226 27132
rect 246 27038 250 27132
rect 270 27038 274 27132
rect 294 27038 298 27132
rect 318 27038 322 27132
rect 342 27038 346 27132
rect 366 27038 370 27132
rect 390 27038 394 27132
rect 414 27038 418 27132
rect 438 27038 442 27132
rect 462 27038 466 27132
rect 486 27038 490 27132
rect 510 27038 514 27132
rect 534 27038 538 27132
rect 558 27038 562 27132
rect 582 27038 586 27132
rect 606 27038 610 27132
rect 630 27038 634 27132
rect 654 27038 658 27132
rect 678 27038 682 27132
rect 702 27038 706 27132
rect 726 27038 730 27132
rect 750 27038 754 27132
rect 774 27038 778 27132
rect 798 27038 802 27132
rect 822 27038 826 27132
rect 846 27038 850 27132
rect 870 27038 874 27132
rect 894 27038 898 27132
rect 918 27038 922 27132
rect 942 27038 946 27132
rect 966 27038 970 27132
rect 990 27038 994 27132
rect 1014 27038 1018 27132
rect 1038 27038 1042 27132
rect 1062 27038 1066 27132
rect 1086 27038 1090 27132
rect 1110 27038 1114 27132
rect 1134 27038 1138 27132
rect 1147 27101 1152 27111
rect 1157 27087 1165 27101
rect 1158 27083 1165 27087
rect 1182 27083 1186 27132
rect 1158 27038 1162 27083
rect 1182 27059 1189 27083
rect 1206 27038 1210 27132
rect 1230 27038 1234 27132
rect 1254 27038 1258 27132
rect 1278 27038 1282 27132
rect 1302 27038 1306 27132
rect 1326 27038 1330 27132
rect 1350 27038 1354 27132
rect 1374 27038 1378 27132
rect 1398 27038 1402 27132
rect 1422 27038 1426 27132
rect 1446 27038 1450 27132
rect 1470 27038 1474 27132
rect 1494 27038 1498 27132
rect 1518 27038 1522 27132
rect 1542 27038 1546 27132
rect 1566 27038 1570 27132
rect 1590 27038 1594 27132
rect 1614 27038 1618 27132
rect 1638 27038 1642 27132
rect 1662 27038 1666 27132
rect 1686 27038 1690 27132
rect 1710 27038 1714 27132
rect 1734 27038 1738 27132
rect 1758 27038 1762 27132
rect 1782 27038 1786 27132
rect 1806 27038 1810 27132
rect 1830 27038 1834 27132
rect 1854 27038 1858 27132
rect 1878 27038 1882 27132
rect 1902 27038 1906 27132
rect 1926 27038 1930 27132
rect 1950 27038 1954 27132
rect 1974 27038 1978 27132
rect 1998 27038 2002 27132
rect 2022 27038 2026 27132
rect 2046 27038 2050 27132
rect 2070 27038 2074 27132
rect 2094 27038 2098 27132
rect 2118 27038 2122 27132
rect 2142 27038 2146 27132
rect 2166 27038 2170 27132
rect 2190 27038 2194 27132
rect 2197 27131 2211 27132
rect 2203 27125 2208 27131
rect 2213 27111 2218 27125
rect 2214 27038 2218 27111
rect 2227 27038 2235 27039
rect -221 27036 2235 27038
rect -221 27029 -216 27036
rect -210 27029 -206 27036
rect -211 27015 -206 27029
rect -221 27014 -187 27015
rect -2393 27012 -187 27014
rect -2371 26990 -2366 27012
rect -2348 26990 -2343 27012
rect -2325 26990 -2320 27012
rect -2072 27010 -2036 27011
rect -2072 27004 -2054 27010
rect -2309 26996 -2301 27004
rect -2317 26990 -2309 26996
rect -2092 26995 -2062 27000
rect -2000 26991 -1992 27012
rect -1938 27011 -1906 27012
rect -1920 27010 -1906 27011
rect -1806 27004 -1680 27010
rect -1854 26995 -1806 27000
rect -1655 26996 -1647 27004
rect -1982 26991 -1966 26992
rect -2000 26990 -1966 26991
rect -1846 26990 -1806 26993
rect -1663 26990 -1655 26996
rect -1642 26990 -1637 27012
rect -1619 26990 -1614 27012
rect -1530 26990 -1526 27012
rect -1506 26990 -1502 27012
rect -1482 26990 -1478 27012
rect -1458 26990 -1454 27012
rect -1434 26990 -1430 27012
rect -1410 26990 -1406 27012
rect -1386 26990 -1382 27012
rect -1362 26990 -1358 27012
rect -1338 26990 -1334 27012
rect -1314 26990 -1310 27012
rect -1290 26990 -1286 27012
rect -1266 26990 -1262 27012
rect -1242 26990 -1238 27012
rect -1218 26990 -1214 27012
rect -1194 26990 -1190 27012
rect -1170 26990 -1166 27012
rect -1146 26990 -1142 27012
rect -1122 26990 -1118 27012
rect -1098 26990 -1094 27012
rect -1074 26990 -1070 27012
rect -1050 26990 -1046 27012
rect -1026 26990 -1022 27012
rect -1002 26990 -998 27012
rect -978 26990 -974 27012
rect -954 26990 -950 27012
rect -930 26990 -926 27012
rect -906 26990 -902 27012
rect -882 26990 -878 27012
rect -858 26990 -854 27012
rect -834 26990 -830 27012
rect -810 26990 -806 27012
rect -786 27011 -782 27012
rect -786 26990 -779 27011
rect -762 26990 -758 27012
rect -738 26990 -734 27012
rect -714 26990 -710 27012
rect -690 26990 -686 27012
rect -666 26990 -662 27012
rect -642 26990 -638 27012
rect -618 26990 -614 27012
rect -594 26990 -590 27012
rect -570 26990 -566 27012
rect -546 26990 -542 27012
rect -522 26990 -518 27012
rect -498 26990 -494 27012
rect -474 26990 -470 27012
rect -450 26990 -446 27012
rect -426 26990 -422 27012
rect -402 26990 -398 27012
rect -378 26990 -374 27012
rect -354 26990 -350 27012
rect -330 26990 -326 27012
rect -2393 26988 -309 26990
rect -2371 26966 -2366 26988
rect -2348 26966 -2343 26988
rect -2325 26966 -2320 26988
rect -2000 26986 -1966 26988
rect -2309 26968 -2301 26976
rect -2062 26975 -2054 26982
rect -2092 26968 -2084 26975
rect -2062 26968 -2026 26970
rect -2317 26966 -2309 26968
rect -2062 26966 -2012 26968
rect -2000 26966 -1992 26986
rect -1982 26985 -1966 26986
rect -1846 26984 -1806 26988
rect -1846 26977 -1798 26982
rect -1806 26975 -1798 26977
rect -1854 26973 -1846 26975
rect -1854 26968 -1806 26973
rect -1655 26968 -1647 26976
rect -1864 26966 -1796 26967
rect -1663 26966 -1655 26968
rect -1642 26966 -1637 26988
rect -1619 26966 -1614 26988
rect -1530 26966 -1526 26988
rect -1506 26966 -1502 26988
rect -1482 26966 -1478 26988
rect -1458 26966 -1454 26988
rect -1434 26966 -1430 26988
rect -1410 26966 -1406 26988
rect -1386 26966 -1382 26988
rect -1362 26966 -1358 26988
rect -1338 26966 -1334 26988
rect -1314 26966 -1310 26988
rect -1290 26966 -1286 26988
rect -1266 26966 -1262 26988
rect -1242 26966 -1238 26988
rect -1218 26966 -1214 26988
rect -1194 26966 -1190 26988
rect -1170 26966 -1166 26988
rect -1146 26966 -1142 26988
rect -1122 26966 -1118 26988
rect -1098 26966 -1094 26988
rect -1074 26966 -1070 26988
rect -1050 26966 -1046 26988
rect -1026 26966 -1022 26988
rect -1002 26966 -998 26988
rect -978 26966 -974 26988
rect -954 26966 -950 26988
rect -930 26966 -926 26988
rect -906 26966 -902 26988
rect -882 26966 -878 26988
rect -858 26966 -854 26988
rect -834 26966 -830 26988
rect -810 26966 -806 26988
rect -803 26987 -789 26988
rect -2393 26964 -789 26966
rect -2371 26918 -2366 26964
rect -2348 26918 -2343 26964
rect -2325 26918 -2320 26964
rect -2317 26960 -2309 26964
rect -2062 26960 -2054 26964
rect -2154 26956 -2138 26958
rect -2057 26956 -2054 26960
rect -2292 26950 -2054 26956
rect -2052 26950 -2044 26960
rect -2092 26934 -2062 26936
rect -2094 26930 -2062 26934
rect -2000 26918 -1992 26964
rect -1846 26957 -1806 26964
rect -1663 26960 -1655 26964
rect -1846 26950 -1680 26956
rect -1854 26934 -1806 26936
rect -1854 26930 -1680 26934
rect -1642 26918 -1637 26964
rect -1619 26918 -1614 26964
rect -1530 26918 -1526 26964
rect -1506 26918 -1502 26964
rect -1482 26918 -1478 26964
rect -1458 26918 -1454 26964
rect -1434 26918 -1430 26964
rect -1410 26918 -1406 26964
rect -1386 26918 -1382 26964
rect -1362 26918 -1358 26964
rect -1338 26918 -1334 26964
rect -1314 26918 -1310 26964
rect -1290 26918 -1286 26964
rect -1266 26918 -1262 26964
rect -1242 26918 -1238 26964
rect -1218 26918 -1214 26964
rect -1194 26918 -1190 26964
rect -1170 26918 -1166 26964
rect -1146 26918 -1142 26964
rect -1122 26918 -1118 26964
rect -1098 26918 -1094 26964
rect -1074 26918 -1070 26964
rect -1050 26918 -1046 26964
rect -1026 26918 -1022 26964
rect -1002 26918 -998 26964
rect -978 26918 -974 26964
rect -954 26918 -950 26964
rect -930 26918 -926 26964
rect -906 26918 -902 26964
rect -882 26918 -878 26964
rect -858 26918 -854 26964
rect -834 26918 -830 26964
rect -810 26918 -806 26964
rect -803 26963 -789 26964
rect -786 26963 -779 26988
rect -786 26918 -782 26963
rect -762 26918 -758 26988
rect -738 26918 -734 26988
rect -714 26918 -710 26988
rect -690 26918 -686 26988
rect -666 26918 -662 26988
rect -642 26918 -638 26988
rect -618 26918 -614 26988
rect -594 26918 -590 26988
rect -570 26918 -566 26988
rect -546 26918 -542 26988
rect -522 26918 -518 26988
rect -498 26918 -494 26988
rect -474 26918 -470 26988
rect -450 26918 -446 26988
rect -426 26918 -422 26988
rect -402 26918 -398 26988
rect -378 26918 -374 26988
rect -354 26918 -350 26988
rect -330 26918 -326 26988
rect -323 26987 -309 26988
rect -306 26987 -299 27011
rect -306 26918 -302 26987
rect -282 26918 -278 27012
rect -258 26918 -254 27012
rect -234 26918 -230 27012
rect -221 27005 -216 27012
rect -211 26991 -206 27005
rect -210 26918 -206 26991
rect -186 26963 -182 27036
rect -2393 26916 -189 26918
rect -2371 26894 -2366 26916
rect -2348 26894 -2343 26916
rect -2325 26894 -2320 26916
rect -2072 26914 -2036 26915
rect -2072 26908 -2054 26914
rect -2309 26900 -2301 26908
rect -2317 26894 -2309 26900
rect -2092 26899 -2062 26904
rect -2000 26895 -1992 26916
rect -1938 26915 -1906 26916
rect -1920 26914 -1906 26915
rect -1806 26908 -1680 26914
rect -1854 26899 -1806 26904
rect -1655 26900 -1647 26908
rect -1982 26895 -1966 26896
rect -2000 26894 -1966 26895
rect -1846 26894 -1806 26897
rect -1663 26894 -1655 26900
rect -1642 26894 -1637 26916
rect -1619 26894 -1614 26916
rect -1530 26894 -1526 26916
rect -1506 26894 -1502 26916
rect -1482 26894 -1478 26916
rect -1458 26894 -1454 26916
rect -1434 26894 -1430 26916
rect -1410 26894 -1406 26916
rect -1386 26894 -1382 26916
rect -1362 26894 -1358 26916
rect -1338 26894 -1334 26916
rect -1314 26894 -1310 26916
rect -1290 26894 -1286 26916
rect -1266 26894 -1262 26916
rect -1242 26894 -1238 26916
rect -1218 26894 -1214 26916
rect -1194 26894 -1190 26916
rect -1170 26894 -1166 26916
rect -1146 26894 -1142 26916
rect -1122 26894 -1118 26916
rect -1098 26894 -1094 26916
rect -1074 26894 -1070 26916
rect -1050 26894 -1046 26916
rect -1026 26894 -1022 26916
rect -1002 26894 -998 26916
rect -978 26894 -974 26916
rect -954 26894 -950 26916
rect -930 26894 -926 26916
rect -906 26894 -902 26916
rect -882 26894 -878 26916
rect -858 26894 -854 26916
rect -834 26894 -830 26916
rect -810 26894 -806 26916
rect -786 26894 -782 26916
rect -762 26894 -758 26916
rect -738 26894 -734 26916
rect -714 26894 -710 26916
rect -690 26894 -686 26916
rect -666 26894 -662 26916
rect -642 26894 -638 26916
rect -618 26894 -614 26916
rect -594 26894 -590 26916
rect -570 26894 -566 26916
rect -546 26894 -542 26916
rect -522 26894 -518 26916
rect -498 26894 -494 26916
rect -474 26894 -470 26916
rect -450 26894 -446 26916
rect -426 26894 -422 26916
rect -402 26894 -398 26916
rect -378 26894 -374 26916
rect -354 26894 -350 26916
rect -330 26894 -326 26916
rect -306 26894 -302 26916
rect -282 26894 -278 26916
rect -258 26894 -254 26916
rect -234 26894 -230 26916
rect -210 26894 -206 26916
rect -203 26915 -189 26916
rect -186 26915 -179 26963
rect -186 26894 -182 26915
rect -162 26894 -158 27036
rect -138 26943 -134 27036
rect -149 26942 -115 26943
rect -114 26942 -110 27036
rect -90 26942 -86 27036
rect -66 26942 -62 27036
rect -42 26942 -38 27036
rect -18 26942 -14 27036
rect 6 26942 10 27036
rect 30 26942 34 27036
rect 54 26942 58 27036
rect 78 26942 82 27036
rect 102 26942 106 27036
rect 126 26942 130 27036
rect 150 26942 154 27036
rect 174 26942 178 27036
rect 198 26942 202 27036
rect 222 26942 226 27036
rect 246 26942 250 27036
rect 270 26942 274 27036
rect 294 26942 298 27036
rect 318 26942 322 27036
rect 342 26942 346 27036
rect 366 26942 370 27036
rect 390 26942 394 27036
rect 414 26942 418 27036
rect 438 26942 442 27036
rect 462 26942 466 27036
rect 486 26942 490 27036
rect 510 26942 514 27036
rect 534 26942 538 27036
rect 558 26942 562 27036
rect 582 26942 586 27036
rect 606 26942 610 27036
rect 619 26957 624 26967
rect 630 26957 634 27036
rect 629 26943 634 26957
rect 630 26942 634 26943
rect 654 26942 658 27036
rect 678 26942 682 27036
rect 702 26942 706 27036
rect 726 26942 730 27036
rect 750 26942 754 27036
rect 774 26942 778 27036
rect 798 26942 802 27036
rect 822 26942 826 27036
rect 846 26942 850 27036
rect 870 26942 874 27036
rect 894 26942 898 27036
rect 918 26942 922 27036
rect 942 26942 946 27036
rect 966 26942 970 27036
rect 990 26942 994 27036
rect 1014 26942 1018 27036
rect 1038 26942 1042 27036
rect 1062 26942 1066 27036
rect 1086 26942 1090 27036
rect 1110 26942 1114 27036
rect 1134 26942 1138 27036
rect 1158 26942 1162 27036
rect 1182 27011 1189 27035
rect 1182 26942 1186 27011
rect 1206 26942 1210 27036
rect 1230 26942 1234 27036
rect 1254 26942 1258 27036
rect 1278 26942 1282 27036
rect 1302 26942 1306 27036
rect 1326 26942 1330 27036
rect 1350 26942 1354 27036
rect 1374 26942 1378 27036
rect 1398 26942 1402 27036
rect 1422 26942 1426 27036
rect 1446 26942 1450 27036
rect 1470 26942 1474 27036
rect 1494 26942 1498 27036
rect 1518 26942 1522 27036
rect 1542 26942 1546 27036
rect 1566 26942 1570 27036
rect 1590 26942 1594 27036
rect 1614 26942 1618 27036
rect 1638 26942 1642 27036
rect 1662 26942 1666 27036
rect 1686 26942 1690 27036
rect 1710 26942 1714 27036
rect 1734 26942 1738 27036
rect 1758 26942 1762 27036
rect 1782 26942 1786 27036
rect 1806 26942 1810 27036
rect 1830 26942 1834 27036
rect 1854 26942 1858 27036
rect 1878 26942 1882 27036
rect 1902 26942 1906 27036
rect 1926 26942 1930 27036
rect 1950 26942 1954 27036
rect 1974 26942 1978 27036
rect 1998 26942 2002 27036
rect 2022 26942 2026 27036
rect 2046 26942 2050 27036
rect 2070 26942 2074 27036
rect 2094 26942 2098 27036
rect 2118 26942 2122 27036
rect 2142 26942 2146 27036
rect 2166 26942 2170 27036
rect 2190 26942 2194 27036
rect 2214 26942 2218 27036
rect 2221 27035 2235 27036
rect 2227 27029 2232 27035
rect 2237 27015 2242 27029
rect 2227 26981 2232 26991
rect 2238 26981 2242 27015
rect 2237 26967 2242 26981
rect 2227 26942 2259 26943
rect -149 26940 2259 26942
rect -149 26933 -144 26940
rect -138 26933 -134 26940
rect -139 26919 -134 26933
rect -149 26909 -144 26919
rect -139 26895 -134 26909
rect -138 26894 -134 26895
rect -114 26894 -110 26940
rect -90 26894 -86 26940
rect -66 26894 -62 26940
rect -42 26894 -38 26940
rect -18 26894 -14 26940
rect 6 26894 10 26940
rect 30 26894 34 26940
rect 54 26894 58 26940
rect 78 26894 82 26940
rect 102 26894 106 26940
rect 126 26894 130 26940
rect 150 26894 154 26940
rect 174 26894 178 26940
rect 198 26894 202 26940
rect 222 26894 226 26940
rect 246 26894 250 26940
rect 270 26895 274 26940
rect 259 26894 293 26895
rect -2393 26892 293 26894
rect -2371 26870 -2366 26892
rect -2348 26870 -2343 26892
rect -2325 26870 -2320 26892
rect -2000 26890 -1966 26892
rect -2309 26872 -2301 26880
rect -2062 26879 -2054 26886
rect -2092 26872 -2084 26879
rect -2062 26872 -2026 26874
rect -2317 26870 -2309 26872
rect -2062 26870 -2012 26872
rect -2000 26870 -1992 26890
rect -1982 26889 -1966 26890
rect -1846 26888 -1806 26892
rect -1846 26881 -1798 26886
rect -1806 26879 -1798 26881
rect -1854 26877 -1846 26879
rect -1854 26872 -1806 26877
rect -1655 26872 -1647 26880
rect -1864 26870 -1796 26871
rect -1663 26870 -1655 26872
rect -1642 26870 -1637 26892
rect -1619 26870 -1614 26892
rect -1530 26870 -1526 26892
rect -1506 26870 -1502 26892
rect -1482 26870 -1478 26892
rect -1458 26870 -1454 26892
rect -1434 26870 -1430 26892
rect -1410 26870 -1406 26892
rect -1386 26870 -1382 26892
rect -1362 26870 -1358 26892
rect -1338 26870 -1334 26892
rect -1314 26870 -1310 26892
rect -1290 26870 -1286 26892
rect -1266 26870 -1262 26892
rect -1242 26870 -1238 26892
rect -1218 26870 -1214 26892
rect -1194 26870 -1190 26892
rect -1170 26870 -1166 26892
rect -1146 26870 -1142 26892
rect -1122 26870 -1118 26892
rect -1098 26870 -1094 26892
rect -1074 26870 -1070 26892
rect -1050 26870 -1046 26892
rect -1026 26870 -1022 26892
rect -1002 26870 -998 26892
rect -978 26870 -974 26892
rect -954 26870 -950 26892
rect -930 26870 -926 26892
rect -906 26870 -902 26892
rect -882 26870 -878 26892
rect -858 26870 -854 26892
rect -834 26870 -830 26892
rect -810 26870 -806 26892
rect -786 26870 -782 26892
rect -762 26870 -758 26892
rect -738 26870 -734 26892
rect -714 26870 -710 26892
rect -690 26870 -686 26892
rect -666 26870 -662 26892
rect -642 26870 -638 26892
rect -618 26870 -614 26892
rect -594 26870 -590 26892
rect -570 26870 -566 26892
rect -546 26870 -542 26892
rect -522 26870 -518 26892
rect -498 26870 -494 26892
rect -474 26870 -470 26892
rect -450 26870 -446 26892
rect -426 26870 -422 26892
rect -402 26870 -398 26892
rect -378 26870 -374 26892
rect -354 26870 -350 26892
rect -330 26870 -326 26892
rect -306 26870 -302 26892
rect -282 26870 -278 26892
rect -258 26870 -254 26892
rect -234 26870 -230 26892
rect -210 26870 -206 26892
rect -186 26870 -182 26892
rect -162 26870 -158 26892
rect -138 26870 -134 26892
rect -114 26870 -110 26892
rect -90 26870 -86 26892
rect -66 26870 -62 26892
rect -42 26870 -38 26892
rect -18 26870 -14 26892
rect 6 26870 10 26892
rect 30 26870 34 26892
rect 54 26870 58 26892
rect 78 26870 82 26892
rect 102 26870 106 26892
rect 126 26870 130 26892
rect 150 26870 154 26892
rect 174 26870 178 26892
rect 198 26870 202 26892
rect 222 26870 226 26892
rect 246 26870 250 26892
rect 259 26885 264 26892
rect 270 26885 274 26892
rect 269 26871 274 26885
rect 270 26870 274 26871
rect 294 26870 298 26940
rect 318 26871 322 26940
rect 307 26870 341 26871
rect -2393 26868 341 26870
rect -2371 26822 -2366 26868
rect -2348 26822 -2343 26868
rect -2325 26822 -2320 26868
rect -2317 26864 -2309 26868
rect -2062 26864 -2054 26868
rect -2154 26860 -2138 26862
rect -2057 26860 -2054 26864
rect -2292 26854 -2054 26860
rect -2052 26854 -2044 26864
rect -2092 26838 -2062 26840
rect -2094 26834 -2062 26838
rect -2000 26822 -1992 26868
rect -1846 26861 -1806 26868
rect -1663 26864 -1655 26868
rect -1846 26854 -1680 26860
rect -1854 26838 -1806 26840
rect -1854 26834 -1680 26838
rect -1642 26822 -1637 26868
rect -1619 26822 -1614 26868
rect -1530 26822 -1526 26868
rect -1506 26822 -1502 26868
rect -1482 26822 -1478 26868
rect -1458 26822 -1454 26868
rect -1434 26822 -1430 26868
rect -1410 26822 -1406 26868
rect -1386 26822 -1382 26868
rect -1362 26822 -1358 26868
rect -1338 26822 -1334 26868
rect -1314 26822 -1310 26868
rect -1290 26822 -1286 26868
rect -1266 26822 -1262 26868
rect -1242 26822 -1238 26868
rect -1218 26822 -1214 26868
rect -1194 26822 -1190 26868
rect -1170 26822 -1166 26868
rect -1146 26822 -1142 26868
rect -1122 26822 -1118 26868
rect -1098 26822 -1094 26868
rect -1074 26822 -1070 26868
rect -1050 26822 -1046 26868
rect -1026 26822 -1022 26868
rect -1002 26822 -998 26868
rect -978 26822 -974 26868
rect -954 26822 -950 26868
rect -930 26822 -926 26868
rect -906 26822 -902 26868
rect -882 26822 -878 26868
rect -858 26822 -854 26868
rect -834 26822 -830 26868
rect -810 26822 -806 26868
rect -786 26822 -782 26868
rect -762 26822 -758 26868
rect -738 26822 -734 26868
rect -714 26822 -710 26868
rect -690 26822 -686 26868
rect -666 26822 -662 26868
rect -642 26822 -638 26868
rect -618 26822 -614 26868
rect -594 26822 -590 26868
rect -570 26822 -566 26868
rect -546 26822 -542 26868
rect -522 26822 -518 26868
rect -498 26822 -494 26868
rect -474 26822 -470 26868
rect -450 26822 -446 26868
rect -426 26822 -422 26868
rect -402 26822 -398 26868
rect -389 26837 -384 26847
rect -378 26837 -374 26868
rect -379 26823 -374 26837
rect -389 26822 -355 26823
rect -2393 26820 -355 26822
rect -2371 26774 -2366 26820
rect -2348 26774 -2343 26820
rect -2325 26774 -2320 26820
rect -2309 26804 -2301 26814
rect -2317 26798 -2309 26804
rect -2097 26798 -2095 26807
rect -2309 26776 -2301 26786
rect -2097 26784 -2095 26788
rect -2292 26783 -2095 26784
rect -2097 26781 -2095 26783
rect -2084 26776 -2083 26819
rect -2069 26812 -2054 26814
rect -2054 26796 -2018 26798
rect -2054 26794 -2004 26796
rect -2059 26790 -2045 26794
rect -2054 26788 -2049 26790
rect -2317 26774 -2309 26776
rect -2084 26774 -2054 26776
rect -2044 26774 -2039 26788
rect -2025 26778 -2014 26784
rect -2000 26778 -1992 26820
rect -1920 26818 -1906 26820
rect -1977 26803 -1929 26809
rect -1655 26804 -1647 26814
rect -1977 26793 -1966 26803
rect -1663 26798 -1655 26804
rect -1977 26781 -1929 26783
rect -2033 26774 -1992 26778
rect -1655 26776 -1647 26786
rect -1663 26774 -1655 26776
rect -1642 26774 -1637 26820
rect -1619 26774 -1614 26820
rect -1530 26774 -1526 26820
rect -1506 26774 -1502 26820
rect -1482 26774 -1478 26820
rect -1458 26774 -1454 26820
rect -1434 26774 -1430 26820
rect -1410 26774 -1406 26820
rect -1386 26774 -1382 26820
rect -1362 26774 -1358 26820
rect -1338 26774 -1334 26820
rect -1314 26774 -1310 26820
rect -1290 26774 -1286 26820
rect -1266 26774 -1262 26820
rect -1242 26774 -1238 26820
rect -1218 26774 -1214 26820
rect -1194 26774 -1190 26820
rect -1170 26774 -1166 26820
rect -1146 26774 -1142 26820
rect -1122 26774 -1118 26820
rect -1098 26774 -1094 26820
rect -1074 26774 -1070 26820
rect -1050 26774 -1046 26820
rect -1026 26774 -1022 26820
rect -1002 26774 -998 26820
rect -978 26774 -974 26820
rect -954 26774 -950 26820
rect -930 26774 -926 26820
rect -906 26774 -902 26820
rect -882 26774 -878 26820
rect -858 26774 -854 26820
rect -834 26774 -830 26820
rect -810 26774 -806 26820
rect -786 26774 -782 26820
rect -762 26774 -758 26820
rect -738 26774 -734 26820
rect -714 26774 -710 26820
rect -690 26774 -686 26820
rect -666 26774 -662 26820
rect -642 26774 -638 26820
rect -618 26774 -614 26820
rect -594 26774 -590 26820
rect -570 26774 -566 26820
rect -546 26774 -542 26820
rect -522 26774 -518 26820
rect -498 26774 -494 26820
rect -474 26774 -470 26820
rect -450 26774 -446 26820
rect -426 26774 -422 26820
rect -402 26774 -398 26820
rect -389 26813 -384 26820
rect -379 26799 -374 26813
rect -378 26774 -374 26799
rect -354 26774 -350 26868
rect -330 26774 -326 26868
rect -306 26774 -302 26868
rect -282 26774 -278 26868
rect -258 26774 -254 26868
rect -234 26774 -230 26868
rect -210 26774 -206 26868
rect -186 26774 -182 26868
rect -162 26774 -158 26868
rect -138 26774 -134 26868
rect -114 26867 -110 26868
rect -114 26846 -107 26867
rect -90 26846 -86 26868
rect -66 26846 -62 26868
rect -42 26846 -38 26868
rect -18 26846 -14 26868
rect 6 26846 10 26868
rect 30 26846 34 26868
rect 54 26846 58 26868
rect 78 26846 82 26868
rect 102 26846 106 26868
rect 126 26846 130 26868
rect 150 26846 154 26868
rect 174 26846 178 26868
rect 198 26846 202 26868
rect 222 26846 226 26868
rect 246 26846 250 26868
rect 270 26846 274 26868
rect 294 26846 298 26868
rect 307 26861 312 26868
rect 318 26861 322 26868
rect 317 26847 322 26861
rect 318 26846 322 26847
rect 342 26846 346 26940
rect 366 26846 370 26940
rect 390 26846 394 26940
rect 414 26846 418 26940
rect 438 26846 442 26940
rect 462 26846 466 26940
rect 486 26846 490 26940
rect 510 26846 514 26940
rect 534 26846 538 26940
rect 558 26846 562 26940
rect 582 26846 586 26940
rect 606 26846 610 26940
rect 630 26846 634 26940
rect 654 26891 658 26940
rect 654 26867 661 26891
rect 654 26846 658 26867
rect 678 26846 682 26940
rect 702 26846 706 26940
rect 726 26846 730 26940
rect 750 26846 754 26940
rect 774 26846 778 26940
rect 798 26846 802 26940
rect 822 26846 826 26940
rect 846 26846 850 26940
rect 870 26846 874 26940
rect 894 26846 898 26940
rect 918 26846 922 26940
rect 942 26846 946 26940
rect 966 26846 970 26940
rect 990 26846 994 26940
rect 1014 26846 1018 26940
rect 1038 26846 1042 26940
rect 1062 26846 1066 26940
rect 1086 26846 1090 26940
rect 1110 26846 1114 26940
rect 1134 26846 1138 26940
rect 1158 26846 1162 26940
rect 1182 26846 1186 26940
rect 1206 26846 1210 26940
rect 1230 26846 1234 26940
rect 1254 26846 1258 26940
rect 1278 26846 1282 26940
rect 1302 26846 1306 26940
rect 1326 26846 1330 26940
rect 1350 26846 1354 26940
rect 1374 26846 1378 26940
rect 1398 26846 1402 26940
rect 1422 26846 1426 26940
rect 1446 26846 1450 26940
rect 1470 26846 1474 26940
rect 1494 26846 1498 26940
rect 1518 26846 1522 26940
rect 1542 26846 1546 26940
rect 1566 26846 1570 26940
rect 1590 26846 1594 26940
rect 1614 26846 1618 26940
rect 1638 26846 1642 26940
rect 1662 26846 1666 26940
rect 1686 26846 1690 26940
rect 1710 26846 1714 26940
rect 1734 26846 1738 26940
rect 1758 26846 1762 26940
rect 1782 26846 1786 26940
rect 1806 26846 1810 26940
rect 1830 26846 1834 26940
rect 1854 26846 1858 26940
rect 1878 26846 1882 26940
rect 1902 26846 1906 26940
rect 1926 26846 1930 26940
rect 1950 26846 1954 26940
rect 1974 26846 1978 26940
rect 1998 26846 2002 26940
rect 2022 26846 2026 26940
rect 2046 26846 2050 26940
rect 2070 26846 2074 26940
rect 2094 26846 2098 26940
rect 2118 26846 2122 26940
rect 2142 26846 2146 26940
rect 2166 26846 2170 26940
rect 2190 26846 2194 26940
rect 2214 26846 2218 26940
rect 2227 26933 2232 26940
rect 2245 26939 2259 26940
rect 2237 26919 2242 26933
rect 2238 26846 2242 26919
rect 2251 26846 2259 26847
rect -131 26844 2259 26846
rect -131 26843 -117 26844
rect -114 26819 -107 26844
rect -114 26774 -110 26819
rect -90 26774 -86 26844
rect -66 26774 -62 26844
rect -42 26774 -38 26844
rect -18 26774 -14 26844
rect 6 26774 10 26844
rect 30 26774 34 26844
rect 54 26774 58 26844
rect 78 26774 82 26844
rect 102 26774 106 26844
rect 126 26774 130 26844
rect 150 26774 154 26844
rect 174 26774 178 26844
rect 198 26774 202 26844
rect 222 26774 226 26844
rect 246 26774 250 26844
rect 270 26774 274 26844
rect 294 26819 298 26844
rect 294 26795 301 26819
rect 294 26774 298 26795
rect 318 26774 322 26844
rect 342 26795 346 26844
rect -2393 26772 339 26774
rect -2371 26654 -2366 26772
rect -2348 26654 -2343 26772
rect -2325 26738 -2320 26772
rect -2317 26770 -2309 26772
rect -2084 26759 -2083 26772
rect -2084 26758 -2054 26759
rect -2325 26730 -2317 26738
rect -2325 26710 -2320 26730
rect -2317 26722 -2309 26730
rect -2117 26721 -2095 26731
rect -2045 26728 -2037 26742
rect -2325 26694 -2317 26710
rect -2325 26678 -2320 26694
rect -2309 26682 -2301 26694
rect -2317 26678 -2309 26682
rect -2117 26680 -2095 26687
rect -2069 26686 -2041 26694
rect -2017 26692 -2015 26694
rect -2325 26666 -2317 26678
rect -2125 26671 -2095 26678
rect -2047 26676 -2011 26678
rect -2059 26674 -2011 26676
rect -2000 26674 -1992 26772
rect -1663 26770 -1655 26772
rect -1969 26721 -1929 26733
rect -1671 26730 -1663 26738
rect -1663 26722 -1655 26730
rect -1671 26694 -1663 26710
rect -1655 26682 -1647 26694
rect -1663 26678 -1655 26682
rect -2125 26669 -2117 26671
rect -2059 26670 -2045 26674
rect -2021 26671 -1992 26674
rect -1977 26671 -1929 26678
rect -2325 26654 -2320 26666
rect -2309 26654 -2301 26666
rect -2131 26661 -2129 26666
rect -2125 26663 -2095 26669
rect -2021 26664 -2009 26668
rect -2125 26661 -2117 26663
rect -2133 26654 -2129 26661
rect -2117 26654 -2087 26661
rect -2025 26658 -2021 26664
rect -2000 26658 -1992 26671
rect -1969 26663 -1929 26669
rect -1671 26666 -1663 26678
rect -2033 26654 -1992 26658
rect -1969 26654 -1921 26661
rect -1655 26654 -1647 26666
rect -1642 26654 -1637 26772
rect -1619 26654 -1614 26772
rect -1530 26654 -1526 26772
rect -1506 26654 -1502 26772
rect -1482 26654 -1478 26772
rect -1458 26654 -1454 26772
rect -1434 26654 -1430 26772
rect -1410 26654 -1406 26772
rect -1386 26654 -1382 26772
rect -1362 26654 -1358 26772
rect -1338 26654 -1334 26772
rect -1314 26654 -1310 26772
rect -1290 26654 -1286 26772
rect -1266 26654 -1262 26772
rect -1242 26654 -1238 26772
rect -1218 26654 -1214 26772
rect -1194 26727 -1190 26772
rect -1205 26726 -1171 26727
rect -1170 26726 -1166 26772
rect -1146 26726 -1142 26772
rect -1122 26726 -1118 26772
rect -1098 26726 -1094 26772
rect -1074 26726 -1070 26772
rect -1050 26726 -1046 26772
rect -1026 26726 -1022 26772
rect -1002 26726 -998 26772
rect -978 26726 -974 26772
rect -954 26726 -950 26772
rect -930 26726 -926 26772
rect -906 26726 -902 26772
rect -882 26726 -878 26772
rect -858 26726 -854 26772
rect -834 26726 -830 26772
rect -810 26726 -806 26772
rect -786 26726 -782 26772
rect -762 26726 -758 26772
rect -738 26726 -734 26772
rect -714 26726 -710 26772
rect -690 26726 -686 26772
rect -666 26726 -662 26772
rect -642 26726 -638 26772
rect -618 26726 -614 26772
rect -594 26726 -590 26772
rect -570 26726 -566 26772
rect -546 26726 -542 26772
rect -522 26726 -518 26772
rect -498 26726 -494 26772
rect -474 26726 -470 26772
rect -450 26726 -446 26772
rect -426 26726 -422 26772
rect -402 26726 -398 26772
rect -378 26726 -374 26772
rect -354 26771 -350 26772
rect -354 26750 -347 26771
rect -330 26750 -326 26772
rect -306 26750 -302 26772
rect -282 26750 -278 26772
rect -258 26750 -254 26772
rect -234 26750 -230 26772
rect -210 26750 -206 26772
rect -186 26750 -182 26772
rect -162 26750 -158 26772
rect -138 26750 -134 26772
rect -114 26750 -110 26772
rect -90 26750 -86 26772
rect -66 26750 -62 26772
rect -42 26750 -38 26772
rect -18 26750 -14 26772
rect 6 26750 10 26772
rect 30 26750 34 26772
rect 54 26750 58 26772
rect 78 26750 82 26772
rect 102 26750 106 26772
rect 126 26750 130 26772
rect 150 26750 154 26772
rect 174 26750 178 26772
rect 198 26750 202 26772
rect 222 26750 226 26772
rect 246 26750 250 26772
rect 270 26750 274 26772
rect 294 26750 298 26772
rect 318 26750 322 26772
rect 325 26771 339 26772
rect 342 26771 349 26795
rect 342 26750 346 26771
rect 366 26750 370 26844
rect 390 26750 394 26844
rect 414 26750 418 26844
rect 438 26750 442 26844
rect 462 26750 466 26844
rect 486 26750 490 26844
rect 510 26750 514 26844
rect 534 26750 538 26844
rect 558 26750 562 26844
rect 582 26750 586 26844
rect 606 26750 610 26844
rect 630 26750 634 26844
rect 654 26750 658 26844
rect 678 26750 682 26844
rect 702 26750 706 26844
rect 726 26750 730 26844
rect 750 26750 754 26844
rect 774 26750 778 26844
rect 798 26750 802 26844
rect 822 26750 826 26844
rect 846 26750 850 26844
rect 870 26750 874 26844
rect 894 26750 898 26844
rect 918 26750 922 26844
rect 942 26750 946 26844
rect 966 26750 970 26844
rect 990 26750 994 26844
rect 1014 26750 1018 26844
rect 1038 26750 1042 26844
rect 1062 26750 1066 26844
rect 1086 26750 1090 26844
rect 1110 26750 1114 26844
rect 1134 26750 1138 26844
rect 1158 26750 1162 26844
rect 1182 26750 1186 26844
rect 1206 26750 1210 26844
rect 1230 26750 1234 26844
rect 1254 26750 1258 26844
rect 1278 26750 1282 26844
rect 1302 26750 1306 26844
rect 1326 26750 1330 26844
rect 1350 26750 1354 26844
rect 1374 26750 1378 26844
rect 1398 26750 1402 26844
rect 1422 26750 1426 26844
rect 1446 26750 1450 26844
rect 1470 26750 1474 26844
rect 1494 26750 1498 26844
rect 1518 26750 1522 26844
rect 1542 26750 1546 26844
rect 1566 26750 1570 26844
rect 1590 26750 1594 26844
rect 1614 26750 1618 26844
rect 1638 26750 1642 26844
rect 1662 26750 1666 26844
rect 1686 26750 1690 26844
rect 1710 26750 1714 26844
rect 1734 26750 1738 26844
rect 1758 26750 1762 26844
rect 1782 26750 1786 26844
rect 1806 26750 1810 26844
rect 1830 26750 1834 26844
rect 1854 26750 1858 26844
rect 1878 26750 1882 26844
rect 1902 26750 1906 26844
rect 1926 26750 1930 26844
rect 1950 26750 1954 26844
rect 1974 26750 1978 26844
rect 1998 26750 2002 26844
rect 2022 26750 2026 26844
rect 2046 26750 2050 26844
rect 2070 26750 2074 26844
rect 2094 26750 2098 26844
rect 2118 26750 2122 26844
rect 2142 26750 2146 26844
rect 2166 26750 2170 26844
rect 2179 26765 2184 26775
rect 2190 26765 2194 26844
rect 2189 26751 2194 26765
rect 2190 26750 2194 26751
rect 2214 26750 2218 26844
rect 2238 26750 2242 26844
rect 2245 26843 2259 26844
rect 2251 26837 2256 26843
rect 2261 26823 2266 26837
rect 2262 26751 2266 26823
rect 2251 26750 2283 26751
rect -371 26748 2283 26750
rect -371 26747 -357 26748
rect -1205 26724 -357 26726
rect -1205 26717 -1200 26724
rect -1194 26717 -1190 26724
rect -1195 26703 -1190 26717
rect -1205 26693 -1200 26703
rect -1195 26679 -1190 26693
rect -1194 26654 -1190 26679
rect -1170 26654 -1166 26724
rect -1146 26654 -1142 26724
rect -1122 26654 -1118 26724
rect -1098 26654 -1094 26724
rect -1074 26654 -1070 26724
rect -1050 26654 -1046 26724
rect -1026 26654 -1022 26724
rect -1002 26654 -998 26724
rect -978 26654 -974 26724
rect -954 26654 -950 26724
rect -930 26654 -926 26724
rect -906 26654 -902 26724
rect -882 26654 -878 26724
rect -858 26654 -854 26724
rect -834 26654 -830 26724
rect -810 26654 -806 26724
rect -786 26654 -782 26724
rect -762 26654 -758 26724
rect -738 26654 -734 26724
rect -714 26654 -710 26724
rect -690 26654 -686 26724
rect -666 26654 -662 26724
rect -642 26654 -638 26724
rect -618 26654 -614 26724
rect -594 26654 -590 26724
rect -570 26654 -566 26724
rect -546 26654 -542 26724
rect -522 26654 -518 26724
rect -498 26654 -494 26724
rect -474 26654 -470 26724
rect -450 26654 -446 26724
rect -426 26654 -422 26724
rect -402 26654 -398 26724
rect -378 26654 -374 26724
rect -371 26723 -357 26724
rect -354 26723 -347 26748
rect -354 26654 -350 26723
rect -330 26654 -326 26748
rect -306 26654 -302 26748
rect -282 26654 -278 26748
rect -258 26654 -254 26748
rect -234 26654 -230 26748
rect -210 26654 -206 26748
rect -186 26654 -182 26748
rect -162 26654 -158 26748
rect -138 26654 -134 26748
rect -114 26654 -110 26748
rect -90 26654 -86 26748
rect -66 26654 -62 26748
rect -42 26654 -38 26748
rect -18 26654 -14 26748
rect 6 26654 10 26748
rect 30 26654 34 26748
rect 54 26654 58 26748
rect 78 26654 82 26748
rect 102 26654 106 26748
rect 126 26654 130 26748
rect 150 26654 154 26748
rect 174 26654 178 26748
rect 198 26654 202 26748
rect 222 26654 226 26748
rect 246 26654 250 26748
rect 270 26654 274 26748
rect 294 26654 298 26748
rect 318 26654 322 26748
rect 342 26654 346 26748
rect 366 26654 370 26748
rect 390 26654 394 26748
rect 414 26654 418 26748
rect 438 26654 442 26748
rect 462 26654 466 26748
rect 486 26654 490 26748
rect 510 26654 514 26748
rect 534 26654 538 26748
rect 558 26654 562 26748
rect 582 26654 586 26748
rect 606 26654 610 26748
rect 630 26654 634 26748
rect 654 26654 658 26748
rect 678 26654 682 26748
rect 702 26654 706 26748
rect 726 26654 730 26748
rect 750 26654 754 26748
rect 774 26654 778 26748
rect 798 26654 802 26748
rect 822 26654 826 26748
rect 846 26654 850 26748
rect 870 26654 874 26748
rect 894 26654 898 26748
rect 918 26654 922 26748
rect 942 26654 946 26748
rect 966 26654 970 26748
rect 990 26654 994 26748
rect 1014 26654 1018 26748
rect 1038 26654 1042 26748
rect 1062 26654 1066 26748
rect 1086 26654 1090 26748
rect 1110 26654 1114 26748
rect 1134 26654 1138 26748
rect 1158 26654 1162 26748
rect 1182 26654 1186 26748
rect 1206 26654 1210 26748
rect 1230 26654 1234 26748
rect 1254 26654 1258 26748
rect 1278 26654 1282 26748
rect 1302 26654 1306 26748
rect 1326 26654 1330 26748
rect 1350 26654 1354 26748
rect 1374 26654 1378 26748
rect 1398 26654 1402 26748
rect 1422 26654 1426 26748
rect 1446 26654 1450 26748
rect 1470 26654 1474 26748
rect 1494 26654 1498 26748
rect 1518 26654 1522 26748
rect 1542 26654 1546 26748
rect 1566 26654 1570 26748
rect 1590 26654 1594 26748
rect 1614 26654 1618 26748
rect 1638 26654 1642 26748
rect 1662 26654 1666 26748
rect 1686 26654 1690 26748
rect 1710 26654 1714 26748
rect 1734 26654 1738 26748
rect 1758 26654 1762 26748
rect 1782 26654 1786 26748
rect 1806 26654 1810 26748
rect 1830 26654 1834 26748
rect 1854 26654 1858 26748
rect 1878 26654 1882 26748
rect 1902 26654 1906 26748
rect 1926 26654 1930 26748
rect 1950 26654 1954 26748
rect 1974 26654 1978 26748
rect 1998 26654 2002 26748
rect 2022 26654 2026 26748
rect 2046 26654 2050 26748
rect 2070 26654 2074 26748
rect 2094 26654 2098 26748
rect 2118 26654 2122 26748
rect 2142 26654 2146 26748
rect 2166 26654 2170 26748
rect 2190 26654 2194 26748
rect 2214 26699 2218 26748
rect 2214 26675 2221 26699
rect 2214 26654 2218 26675
rect 2238 26654 2242 26748
rect 2251 26741 2256 26748
rect 2262 26741 2266 26748
rect 2269 26747 2283 26748
rect 2261 26727 2266 26741
rect 2251 26717 2256 26727
rect 2261 26703 2266 26717
rect 2262 26655 2266 26703
rect 2251 26654 2283 26655
rect -2393 26652 2283 26654
rect -2371 26534 -2366 26652
rect -2348 26534 -2343 26652
rect -2325 26650 -2320 26652
rect -2317 26650 -2309 26652
rect -2131 26650 -2129 26652
rect -2125 26650 -2095 26652
rect -2325 26638 -2317 26650
rect -2117 26645 -2095 26650
rect -2325 26618 -2320 26638
rect -2325 26610 -2317 26618
rect -2325 26590 -2320 26610
rect -2317 26602 -2309 26610
rect -2117 26601 -2095 26611
rect -2045 26608 -2037 26622
rect -2325 26574 -2317 26590
rect -2325 26558 -2320 26574
rect -2309 26562 -2301 26574
rect -2317 26558 -2309 26562
rect -2117 26560 -2095 26567
rect -2069 26566 -2041 26574
rect -2017 26572 -2015 26574
rect -2325 26546 -2317 26558
rect -2125 26551 -2095 26558
rect -2047 26556 -2011 26558
rect -2059 26554 -2011 26556
rect -2000 26554 -1992 26652
rect -1663 26650 -1655 26652
rect -1671 26638 -1663 26650
rect -1969 26601 -1929 26613
rect -1671 26610 -1663 26618
rect -1663 26602 -1655 26610
rect -1671 26574 -1663 26590
rect -1655 26562 -1647 26574
rect -1663 26558 -1655 26562
rect -2125 26549 -2117 26551
rect -2059 26550 -2045 26554
rect -2021 26551 -1992 26554
rect -1977 26551 -1929 26558
rect -2325 26534 -2320 26546
rect -2309 26534 -2301 26546
rect -2131 26541 -2129 26546
rect -2125 26543 -2095 26549
rect -2021 26544 -2009 26548
rect -2125 26541 -2117 26543
rect -2133 26534 -2129 26541
rect -2117 26534 -2087 26541
rect -2025 26538 -2021 26544
rect -2000 26538 -1992 26551
rect -1969 26543 -1929 26549
rect -1671 26546 -1663 26558
rect -2033 26534 -1992 26538
rect -1969 26534 -1921 26541
rect -1655 26534 -1647 26546
rect -1642 26534 -1637 26652
rect -1619 26534 -1614 26652
rect -1589 26534 -1555 26535
rect -2393 26532 -1555 26534
rect -2371 26438 -2366 26532
rect -2348 26438 -2343 26532
rect -2325 26530 -2320 26532
rect -2317 26530 -2309 26532
rect -2131 26530 -2129 26532
rect -2125 26530 -2095 26532
rect -2325 26518 -2317 26530
rect -2117 26525 -2095 26530
rect -2325 26498 -2320 26518
rect -2325 26490 -2317 26498
rect -2325 26438 -2320 26490
rect -2317 26482 -2309 26490
rect -2117 26481 -2095 26491
rect -2045 26488 -2037 26502
rect -2309 26442 -2301 26452
rect -2087 26448 -2076 26456
rect -2017 26452 -2015 26459
rect -2317 26438 -2309 26442
rect -2092 26440 -2087 26448
rect -2092 26438 -2077 26439
rect -2000 26438 -1992 26532
rect -1663 26530 -1655 26532
rect -1671 26518 -1663 26530
rect -1969 26481 -1929 26493
rect -1671 26490 -1663 26498
rect -1663 26482 -1655 26490
rect -1655 26442 -1647 26452
rect -1928 26438 -1924 26439
rect -1854 26438 -1680 26439
rect -1663 26438 -1655 26442
rect -1642 26438 -1637 26532
rect -1619 26438 -1614 26532
rect -1554 26446 -1547 26459
rect -2393 26436 -1557 26438
rect -2371 26414 -2366 26436
rect -2348 26414 -2343 26436
rect -2325 26414 -2320 26436
rect -2092 26431 -2037 26436
rect -2021 26431 -1969 26436
rect -1921 26431 -1913 26436
rect -1854 26432 -1680 26436
rect -2100 26429 -2092 26430
rect -2309 26414 -2301 26424
rect -2100 26423 -2087 26429
rect -2051 26416 -2026 26418
rect -2062 26414 -2012 26416
rect -2000 26414 -1992 26431
rect -1969 26423 -1921 26430
rect -1969 26414 -1964 26423
rect -1864 26414 -1796 26415
rect -1655 26414 -1647 26424
rect -1642 26414 -1637 26436
rect -1619 26414 -1614 26436
rect -1571 26435 -1557 26436
rect -1554 26435 -1547 26436
rect -1530 26414 -1526 26652
rect -1506 26414 -1502 26652
rect -1482 26414 -1478 26652
rect -1458 26414 -1454 26652
rect -1434 26414 -1430 26652
rect -1410 26414 -1406 26652
rect -1386 26414 -1382 26652
rect -1362 26414 -1358 26652
rect -1338 26414 -1334 26652
rect -1314 26414 -1310 26652
rect -1290 26414 -1286 26652
rect -1266 26414 -1262 26652
rect -1242 26414 -1238 26652
rect -1218 26414 -1214 26652
rect -1194 26414 -1190 26652
rect -1170 26651 -1166 26652
rect -1170 26630 -1163 26651
rect -1146 26630 -1142 26652
rect -1122 26630 -1118 26652
rect -1098 26630 -1094 26652
rect -1074 26630 -1070 26652
rect -1050 26630 -1046 26652
rect -1026 26630 -1022 26652
rect -1002 26630 -998 26652
rect -978 26630 -974 26652
rect -954 26630 -950 26652
rect -930 26630 -926 26652
rect -906 26630 -902 26652
rect -882 26630 -878 26652
rect -858 26630 -854 26652
rect -834 26630 -830 26652
rect -810 26630 -806 26652
rect -786 26630 -782 26652
rect -762 26630 -758 26652
rect -738 26630 -734 26652
rect -714 26630 -710 26652
rect -690 26630 -686 26652
rect -666 26630 -662 26652
rect -642 26630 -638 26652
rect -618 26630 -614 26652
rect -594 26630 -590 26652
rect -570 26630 -566 26652
rect -546 26630 -542 26652
rect -522 26630 -518 26652
rect -498 26630 -494 26652
rect -474 26630 -470 26652
rect -450 26630 -446 26652
rect -426 26630 -422 26652
rect -402 26630 -398 26652
rect -378 26630 -374 26652
rect -354 26630 -350 26652
rect -330 26630 -326 26652
rect -306 26630 -302 26652
rect -282 26630 -278 26652
rect -258 26630 -254 26652
rect -234 26630 -230 26652
rect -210 26630 -206 26652
rect -186 26630 -182 26652
rect -162 26630 -158 26652
rect -138 26630 -134 26652
rect -114 26630 -110 26652
rect -90 26630 -86 26652
rect -66 26630 -62 26652
rect -42 26630 -38 26652
rect -18 26630 -14 26652
rect 6 26630 10 26652
rect 30 26630 34 26652
rect 54 26630 58 26652
rect 78 26630 82 26652
rect 102 26630 106 26652
rect 126 26630 130 26652
rect 150 26630 154 26652
rect 174 26630 178 26652
rect 198 26630 202 26652
rect 222 26630 226 26652
rect 246 26630 250 26652
rect 270 26630 274 26652
rect 294 26630 298 26652
rect 318 26630 322 26652
rect 342 26630 346 26652
rect 366 26630 370 26652
rect 390 26630 394 26652
rect 414 26630 418 26652
rect 438 26630 442 26652
rect 462 26630 466 26652
rect 486 26630 490 26652
rect 510 26630 514 26652
rect 534 26630 538 26652
rect 558 26630 562 26652
rect 582 26630 586 26652
rect 606 26630 610 26652
rect 630 26630 634 26652
rect 654 26630 658 26652
rect 678 26630 682 26652
rect 702 26630 706 26652
rect 726 26630 730 26652
rect 750 26630 754 26652
rect 774 26630 778 26652
rect 798 26630 802 26652
rect 822 26630 826 26652
rect 846 26630 850 26652
rect 870 26630 874 26652
rect 894 26631 898 26652
rect 883 26630 917 26631
rect -1187 26628 917 26630
rect -1187 26627 -1173 26628
rect -1170 26603 -1163 26628
rect -1170 26414 -1166 26603
rect -1146 26414 -1142 26628
rect -1122 26414 -1118 26628
rect -1098 26414 -1094 26628
rect -1074 26414 -1070 26628
rect -1050 26414 -1046 26628
rect -1026 26414 -1022 26628
rect -1002 26414 -998 26628
rect -989 26597 -984 26607
rect -978 26597 -974 26628
rect -979 26583 -974 26597
rect -989 26573 -984 26583
rect -979 26559 -974 26573
rect -978 26414 -974 26559
rect -954 26531 -950 26628
rect -954 26510 -947 26531
rect -930 26510 -926 26628
rect -906 26510 -902 26628
rect -882 26510 -878 26628
rect -858 26510 -854 26628
rect -834 26510 -830 26628
rect -810 26510 -806 26628
rect -786 26510 -782 26628
rect -762 26510 -758 26628
rect -738 26510 -734 26628
rect -714 26510 -710 26628
rect -690 26510 -686 26628
rect -666 26510 -662 26628
rect -642 26510 -638 26628
rect -618 26510 -614 26628
rect -594 26510 -590 26628
rect -570 26510 -566 26628
rect -546 26510 -542 26628
rect -522 26510 -518 26628
rect -498 26510 -494 26628
rect -474 26510 -470 26628
rect -450 26510 -446 26628
rect -426 26510 -422 26628
rect -402 26510 -398 26628
rect -378 26510 -374 26628
rect -354 26510 -350 26628
rect -330 26510 -326 26628
rect -306 26510 -302 26628
rect -282 26510 -278 26628
rect -258 26510 -254 26628
rect -234 26510 -230 26628
rect -210 26510 -206 26628
rect -186 26510 -182 26628
rect -162 26510 -158 26628
rect -138 26510 -134 26628
rect -114 26511 -110 26628
rect -125 26510 -91 26511
rect -971 26508 -91 26510
rect -971 26507 -957 26508
rect -954 26483 -947 26508
rect -954 26414 -950 26483
rect -930 26414 -926 26508
rect -906 26414 -902 26508
rect -882 26414 -878 26508
rect -858 26414 -854 26508
rect -834 26414 -830 26508
rect -810 26414 -806 26508
rect -786 26414 -782 26508
rect -762 26414 -758 26508
rect -749 26429 -744 26439
rect -738 26429 -734 26508
rect -739 26415 -734 26429
rect -738 26414 -734 26415
rect -714 26414 -710 26508
rect -690 26414 -686 26508
rect -666 26414 -662 26508
rect -642 26414 -638 26508
rect -618 26414 -614 26508
rect -594 26414 -590 26508
rect -570 26414 -566 26508
rect -546 26414 -542 26508
rect -522 26414 -518 26508
rect -498 26414 -494 26508
rect -474 26414 -470 26508
rect -450 26414 -446 26508
rect -426 26414 -422 26508
rect -402 26414 -398 26508
rect -378 26414 -374 26508
rect -354 26414 -350 26508
rect -330 26414 -326 26508
rect -306 26414 -302 26508
rect -282 26414 -278 26508
rect -258 26414 -254 26508
rect -234 26414 -230 26508
rect -210 26414 -206 26508
rect -186 26414 -182 26508
rect -162 26414 -158 26508
rect -138 26414 -134 26508
rect -125 26501 -120 26508
rect -114 26501 -110 26508
rect -115 26487 -110 26501
rect -114 26414 -110 26487
rect -90 26435 -86 26628
rect -2393 26412 -93 26414
rect -2371 26366 -2366 26412
rect -2348 26366 -2343 26412
rect -2325 26366 -2320 26412
rect -2317 26408 -2309 26412
rect -2105 26405 -2092 26408
rect -2092 26382 -2062 26384
rect -2094 26378 -2062 26382
rect -2000 26366 -1992 26412
rect -1663 26408 -1655 26412
rect -1969 26405 -1921 26408
rect -1854 26382 -1806 26384
rect -1854 26378 -1680 26382
rect -1642 26366 -1637 26412
rect -1619 26366 -1614 26412
rect -1530 26366 -1526 26412
rect -1506 26366 -1502 26412
rect -1482 26366 -1478 26412
rect -1458 26366 -1454 26412
rect -1434 26366 -1430 26412
rect -1410 26366 -1406 26412
rect -1386 26366 -1382 26412
rect -1362 26366 -1358 26412
rect -1338 26366 -1334 26412
rect -1314 26366 -1310 26412
rect -1290 26366 -1286 26412
rect -1266 26366 -1262 26412
rect -1242 26366 -1238 26412
rect -1218 26366 -1214 26412
rect -1194 26366 -1190 26412
rect -1170 26366 -1166 26412
rect -1146 26366 -1142 26412
rect -1122 26366 -1118 26412
rect -1098 26366 -1094 26412
rect -1074 26366 -1070 26412
rect -1050 26366 -1046 26412
rect -1026 26366 -1022 26412
rect -1002 26366 -998 26412
rect -978 26366 -974 26412
rect -954 26366 -950 26412
rect -930 26366 -926 26412
rect -906 26366 -902 26412
rect -882 26366 -878 26412
rect -858 26366 -854 26412
rect -834 26366 -830 26412
rect -810 26366 -806 26412
rect -786 26366 -782 26412
rect -762 26366 -758 26412
rect -738 26366 -734 26412
rect -714 26366 -710 26412
rect -690 26366 -686 26412
rect -666 26366 -662 26412
rect -642 26366 -638 26412
rect -618 26366 -614 26412
rect -594 26366 -590 26412
rect -570 26366 -566 26412
rect -546 26366 -542 26412
rect -522 26366 -518 26412
rect -498 26366 -494 26412
rect -474 26366 -470 26412
rect -450 26366 -446 26412
rect -426 26366 -422 26412
rect -402 26366 -398 26412
rect -378 26366 -374 26412
rect -354 26366 -350 26412
rect -330 26366 -326 26412
rect -306 26366 -302 26412
rect -282 26366 -278 26412
rect -258 26366 -254 26412
rect -234 26366 -230 26412
rect -210 26366 -206 26412
rect -186 26366 -182 26412
rect -162 26366 -158 26412
rect -138 26366 -134 26412
rect -114 26366 -110 26412
rect -107 26411 -93 26412
rect -90 26411 -83 26435
rect -90 26366 -86 26411
rect -66 26366 -62 26628
rect -42 26366 -38 26628
rect -18 26366 -14 26628
rect 6 26366 10 26628
rect 30 26366 34 26628
rect 54 26366 58 26628
rect 78 26366 82 26628
rect 102 26366 106 26628
rect 126 26366 130 26628
rect 150 26366 154 26628
rect 174 26366 178 26628
rect 198 26366 202 26628
rect 222 26366 226 26628
rect 246 26366 250 26628
rect 270 26366 274 26628
rect 294 26366 298 26628
rect 318 26366 322 26628
rect 342 26366 346 26628
rect 366 26366 370 26628
rect 390 26366 394 26628
rect 414 26366 418 26628
rect 438 26366 442 26628
rect 462 26366 466 26628
rect 486 26366 490 26628
rect 510 26366 514 26628
rect 534 26366 538 26628
rect 558 26366 562 26628
rect 582 26366 586 26628
rect 606 26366 610 26628
rect 630 26366 634 26628
rect 654 26366 658 26628
rect 678 26366 682 26628
rect 702 26366 706 26628
rect 726 26366 730 26628
rect 750 26366 754 26628
rect 774 26366 778 26628
rect 798 26366 802 26628
rect 822 26366 826 26628
rect 846 26366 850 26628
rect 870 26366 874 26628
rect 883 26621 888 26628
rect 894 26621 898 26628
rect 893 26607 898 26621
rect 894 26366 898 26607
rect 918 26555 922 26652
rect 918 26531 925 26555
rect 918 26366 922 26531
rect 942 26366 946 26652
rect 966 26366 970 26652
rect 990 26366 994 26652
rect 1014 26366 1018 26652
rect 1038 26366 1042 26652
rect 1062 26366 1066 26652
rect 1075 26477 1080 26487
rect 1086 26477 1090 26652
rect 1085 26463 1090 26477
rect 1075 26453 1080 26463
rect 1085 26439 1090 26453
rect 1086 26366 1090 26439
rect 1110 26411 1114 26652
rect -2393 26364 1107 26366
rect -2371 26342 -2366 26364
rect -2348 26342 -2343 26364
rect -2325 26342 -2320 26364
rect -2072 26362 -2036 26363
rect -2072 26356 -2054 26362
rect -2309 26348 -2301 26356
rect -2317 26342 -2309 26348
rect -2092 26347 -2062 26352
rect -2000 26343 -1992 26364
rect -1938 26363 -1906 26364
rect -1920 26362 -1906 26363
rect -1806 26356 -1680 26362
rect -1854 26347 -1806 26352
rect -1655 26348 -1647 26356
rect -1982 26343 -1966 26344
rect -2000 26342 -1966 26343
rect -1846 26342 -1806 26345
rect -1663 26342 -1655 26348
rect -1642 26342 -1637 26364
rect -1619 26342 -1614 26364
rect -1530 26342 -1526 26364
rect -1506 26342 -1502 26364
rect -1482 26342 -1478 26364
rect -1458 26342 -1454 26364
rect -1434 26342 -1430 26364
rect -1410 26342 -1406 26364
rect -1386 26342 -1382 26364
rect -1362 26342 -1358 26364
rect -1338 26342 -1334 26364
rect -1314 26342 -1310 26364
rect -1290 26342 -1286 26364
rect -1266 26342 -1262 26364
rect -1242 26342 -1238 26364
rect -1218 26342 -1214 26364
rect -1194 26342 -1190 26364
rect -1170 26342 -1166 26364
rect -1146 26342 -1142 26364
rect -1122 26342 -1118 26364
rect -1098 26342 -1094 26364
rect -1074 26342 -1070 26364
rect -1050 26342 -1046 26364
rect -1026 26342 -1022 26364
rect -1002 26342 -998 26364
rect -978 26342 -974 26364
rect -954 26342 -950 26364
rect -930 26342 -926 26364
rect -906 26342 -902 26364
rect -882 26342 -878 26364
rect -858 26342 -854 26364
rect -834 26342 -830 26364
rect -810 26342 -806 26364
rect -786 26342 -782 26364
rect -762 26342 -758 26364
rect -738 26343 -734 26364
rect -714 26363 -710 26364
rect -749 26342 -717 26343
rect -2393 26340 -717 26342
rect -2371 26318 -2366 26340
rect -2348 26318 -2343 26340
rect -2325 26318 -2320 26340
rect -2000 26338 -1966 26340
rect -2309 26320 -2301 26328
rect -2062 26327 -2054 26334
rect -2092 26320 -2084 26327
rect -2062 26320 -2026 26322
rect -2317 26318 -2309 26320
rect -2062 26318 -2012 26320
rect -2000 26318 -1992 26338
rect -1982 26337 -1966 26338
rect -1846 26336 -1806 26340
rect -1846 26329 -1798 26334
rect -1806 26327 -1798 26329
rect -1854 26325 -1846 26327
rect -1854 26320 -1806 26325
rect -1655 26320 -1647 26328
rect -1864 26318 -1796 26319
rect -1663 26318 -1655 26320
rect -1642 26318 -1637 26340
rect -1619 26318 -1614 26340
rect -1530 26318 -1526 26340
rect -1506 26318 -1502 26340
rect -1482 26318 -1478 26340
rect -1458 26318 -1454 26340
rect -1434 26318 -1430 26340
rect -1410 26318 -1406 26340
rect -1386 26318 -1382 26340
rect -1362 26318 -1358 26340
rect -1338 26318 -1334 26340
rect -1314 26318 -1310 26340
rect -1290 26318 -1286 26340
rect -1266 26318 -1262 26340
rect -1242 26318 -1238 26340
rect -1218 26318 -1214 26340
rect -1194 26318 -1190 26340
rect -1170 26318 -1166 26340
rect -1146 26318 -1142 26340
rect -1122 26318 -1118 26340
rect -1098 26318 -1094 26340
rect -1074 26318 -1070 26340
rect -1050 26318 -1046 26340
rect -1026 26318 -1022 26340
rect -1002 26318 -998 26340
rect -978 26318 -974 26340
rect -954 26318 -950 26340
rect -930 26318 -926 26340
rect -906 26318 -902 26340
rect -882 26318 -878 26340
rect -858 26318 -854 26340
rect -834 26318 -830 26340
rect -810 26318 -806 26340
rect -786 26318 -782 26340
rect -762 26318 -758 26340
rect -749 26333 -744 26340
rect -738 26333 -734 26340
rect -731 26339 -717 26340
rect -714 26339 -707 26363
rect -739 26319 -734 26333
rect -738 26318 -734 26319
rect -714 26318 -710 26339
rect -690 26318 -686 26364
rect -666 26318 -662 26364
rect -642 26318 -638 26364
rect -618 26318 -614 26364
rect -594 26318 -590 26364
rect -570 26318 -566 26364
rect -546 26318 -542 26364
rect -522 26318 -518 26364
rect -498 26318 -494 26364
rect -474 26318 -470 26364
rect -450 26318 -446 26364
rect -426 26318 -422 26364
rect -402 26318 -398 26364
rect -378 26318 -374 26364
rect -354 26318 -350 26364
rect -330 26318 -326 26364
rect -306 26318 -302 26364
rect -282 26318 -278 26364
rect -258 26318 -254 26364
rect -234 26318 -230 26364
rect -210 26318 -206 26364
rect -186 26318 -182 26364
rect -162 26318 -158 26364
rect -138 26318 -134 26364
rect -114 26318 -110 26364
rect -90 26318 -86 26364
rect -66 26318 -62 26364
rect -42 26318 -38 26364
rect -18 26318 -14 26364
rect 6 26318 10 26364
rect 30 26318 34 26364
rect 54 26318 58 26364
rect 78 26318 82 26364
rect 102 26318 106 26364
rect 126 26318 130 26364
rect 150 26318 154 26364
rect 174 26318 178 26364
rect 198 26318 202 26364
rect 222 26318 226 26364
rect 246 26318 250 26364
rect 270 26318 274 26364
rect 294 26318 298 26364
rect 318 26318 322 26364
rect 342 26318 346 26364
rect 366 26318 370 26364
rect 390 26318 394 26364
rect 414 26318 418 26364
rect 438 26318 442 26364
rect 462 26318 466 26364
rect 486 26318 490 26364
rect 510 26318 514 26364
rect 534 26318 538 26364
rect 558 26318 562 26364
rect 582 26318 586 26364
rect 606 26318 610 26364
rect 630 26318 634 26364
rect 654 26318 658 26364
rect 678 26318 682 26364
rect 702 26318 706 26364
rect 726 26318 730 26364
rect 750 26318 754 26364
rect 774 26318 778 26364
rect 798 26318 802 26364
rect 822 26318 826 26364
rect 846 26318 850 26364
rect 870 26318 874 26364
rect 894 26318 898 26364
rect 918 26318 922 26364
rect 942 26318 946 26364
rect 966 26318 970 26364
rect 990 26318 994 26364
rect 1014 26318 1018 26364
rect 1038 26318 1042 26364
rect 1062 26318 1066 26364
rect 1086 26318 1090 26364
rect 1093 26363 1107 26364
rect 1110 26363 1117 26411
rect 1110 26318 1114 26363
rect 1134 26318 1138 26652
rect 1158 26318 1162 26652
rect 1182 26318 1186 26652
rect 1206 26318 1210 26652
rect 1230 26318 1234 26652
rect 1254 26318 1258 26652
rect 1278 26318 1282 26652
rect 1302 26318 1306 26652
rect 1326 26318 1330 26652
rect 1350 26318 1354 26652
rect 1374 26318 1378 26652
rect 1398 26318 1402 26652
rect 1422 26318 1426 26652
rect 1446 26318 1450 26652
rect 1470 26318 1474 26652
rect 1494 26318 1498 26652
rect 1518 26318 1522 26652
rect 1542 26318 1546 26652
rect 1566 26318 1570 26652
rect 1590 26318 1594 26652
rect 1614 26318 1618 26652
rect 1638 26318 1642 26652
rect 1662 26318 1666 26652
rect 1686 26318 1690 26652
rect 1710 26318 1714 26652
rect 1734 26318 1738 26652
rect 1758 26318 1762 26652
rect 1782 26318 1786 26652
rect 1806 26391 1810 26652
rect 1795 26390 1829 26391
rect 1830 26390 1834 26652
rect 1854 26390 1858 26652
rect 1878 26390 1882 26652
rect 1902 26390 1906 26652
rect 1926 26390 1930 26652
rect 1950 26390 1954 26652
rect 1974 26390 1978 26652
rect 1998 26390 2002 26652
rect 2022 26390 2026 26652
rect 2046 26390 2050 26652
rect 2070 26390 2074 26652
rect 2094 26390 2098 26652
rect 2118 26390 2122 26652
rect 2142 26390 2146 26652
rect 2166 26390 2170 26652
rect 2190 26390 2194 26652
rect 2214 26390 2218 26652
rect 2238 26390 2242 26652
rect 2251 26645 2256 26652
rect 2262 26645 2266 26652
rect 2269 26651 2283 26652
rect 2261 26631 2266 26645
rect 2275 26641 2283 26645
rect 2269 26631 2275 26641
rect 2251 26597 2256 26607
rect 2261 26583 2266 26597
rect 2262 26390 2266 26583
rect 2275 26477 2280 26487
rect 2285 26463 2290 26477
rect 2275 26405 2280 26415
rect 2286 26405 2290 26463
rect 2285 26391 2290 26405
rect 2299 26401 2307 26405
rect 2293 26391 2299 26401
rect 2275 26390 2307 26391
rect 1795 26388 2307 26390
rect 1795 26381 1800 26388
rect 1806 26381 1810 26388
rect 1805 26367 1810 26381
rect 1795 26357 1800 26367
rect 1805 26343 1810 26357
rect 1806 26318 1810 26343
rect 1830 26318 1834 26388
rect 1854 26318 1858 26388
rect 1878 26318 1882 26388
rect 1902 26318 1906 26388
rect 1926 26318 1930 26388
rect 1950 26318 1954 26388
rect 1974 26318 1978 26388
rect 1998 26318 2002 26388
rect 2022 26318 2026 26388
rect 2046 26318 2050 26388
rect 2070 26318 2074 26388
rect 2094 26318 2098 26388
rect 2118 26318 2122 26388
rect 2142 26318 2146 26388
rect 2166 26318 2170 26388
rect 2190 26318 2194 26388
rect 2214 26318 2218 26388
rect 2238 26318 2242 26388
rect 2262 26318 2266 26388
rect 2275 26381 2280 26388
rect 2293 26387 2307 26388
rect 2285 26367 2290 26381
rect 2286 26319 2290 26367
rect 2275 26318 2307 26319
rect -2393 26316 2307 26318
rect -2371 26270 -2366 26316
rect -2348 26270 -2343 26316
rect -2325 26280 -2320 26316
rect -2317 26312 -2309 26316
rect -2062 26312 -2054 26316
rect -2154 26308 -2138 26310
rect -2057 26308 -2054 26312
rect -2292 26302 -2054 26308
rect -2052 26302 -2044 26312
rect -2092 26286 -2062 26288
rect -2094 26282 -2062 26286
rect -2325 26270 -2317 26280
rect -2095 26272 -2084 26276
rect -2000 26273 -1992 26316
rect -1846 26309 -1806 26316
rect -1663 26312 -1655 26316
rect -1846 26302 -1680 26308
rect -1854 26286 -1806 26288
rect -1854 26282 -1680 26286
rect -2119 26270 -2069 26272
rect -2054 26270 -1892 26273
rect -1671 26270 -1663 26280
rect -1642 26270 -1637 26316
rect -1619 26270 -1614 26316
rect -1530 26270 -1526 26316
rect -1506 26270 -1502 26316
rect -1482 26270 -1478 26316
rect -1458 26270 -1454 26316
rect -1434 26270 -1430 26316
rect -1410 26270 -1406 26316
rect -1386 26270 -1382 26316
rect -1362 26270 -1358 26316
rect -1338 26270 -1334 26316
rect -1314 26270 -1310 26316
rect -1290 26270 -1286 26316
rect -1266 26270 -1262 26316
rect -1242 26270 -1238 26316
rect -1218 26270 -1214 26316
rect -1194 26270 -1190 26316
rect -1170 26270 -1166 26316
rect -1146 26270 -1142 26316
rect -1122 26270 -1118 26316
rect -1098 26270 -1094 26316
rect -1074 26270 -1070 26316
rect -1050 26270 -1046 26316
rect -1026 26270 -1022 26316
rect -1002 26270 -998 26316
rect -978 26270 -974 26316
rect -954 26270 -950 26316
rect -930 26270 -926 26316
rect -906 26270 -902 26316
rect -882 26270 -878 26316
rect -858 26270 -854 26316
rect -834 26270 -830 26316
rect -810 26270 -806 26316
rect -786 26270 -782 26316
rect -762 26270 -758 26316
rect -738 26270 -734 26316
rect -714 26270 -710 26316
rect -690 26270 -686 26316
rect -666 26270 -662 26316
rect -642 26270 -638 26316
rect -618 26270 -614 26316
rect -594 26270 -590 26316
rect -570 26270 -566 26316
rect -546 26270 -542 26316
rect -522 26270 -518 26316
rect -498 26270 -494 26316
rect -474 26270 -470 26316
rect -450 26270 -446 26316
rect -426 26270 -422 26316
rect -402 26270 -398 26316
rect -378 26270 -374 26316
rect -354 26270 -350 26316
rect -330 26270 -326 26316
rect -306 26270 -302 26316
rect -282 26270 -278 26316
rect -258 26270 -254 26316
rect -234 26270 -230 26316
rect -210 26270 -206 26316
rect -186 26270 -182 26316
rect -162 26270 -158 26316
rect -138 26270 -134 26316
rect -114 26270 -110 26316
rect -90 26270 -86 26316
rect -77 26285 -72 26295
rect -66 26285 -62 26316
rect -67 26271 -62 26285
rect -77 26270 -43 26271
rect -2393 26268 -43 26270
rect -2371 26246 -2366 26268
rect -2348 26246 -2343 26268
rect -2325 26264 -2317 26268
rect -2325 26248 -2320 26264
rect -2309 26252 -2301 26264
rect -2095 26262 -2084 26268
rect -2054 26267 -1906 26268
rect -2054 26266 -2036 26267
rect -2084 26260 -2079 26262
rect -2317 26248 -2309 26252
rect -2092 26251 -2079 26258
rect -2000 26254 -1992 26267
rect -1920 26266 -1906 26267
rect -1671 26264 -1663 26268
rect -1846 26260 -1806 26262
rect -1854 26254 -1806 26258
rect -2054 26251 -1982 26254
rect -1966 26251 -1806 26254
rect -1655 26252 -1647 26264
rect -2003 26248 -1992 26251
rect -1904 26249 -1902 26251
rect -1854 26249 -1846 26251
rect -2325 26246 -2317 26248
rect -2033 26246 -1992 26248
rect -1854 26247 -1806 26249
rect -1663 26248 -1655 26252
rect -1864 26246 -1796 26247
rect -1671 26246 -1663 26248
rect -1642 26246 -1637 26268
rect -1619 26246 -1614 26268
rect -1530 26246 -1526 26268
rect -1506 26246 -1502 26268
rect -1482 26246 -1478 26268
rect -1458 26246 -1454 26268
rect -1434 26246 -1430 26268
rect -1410 26246 -1406 26268
rect -1386 26246 -1382 26268
rect -1362 26246 -1358 26268
rect -1338 26246 -1334 26268
rect -1314 26246 -1310 26268
rect -1290 26246 -1286 26268
rect -1266 26246 -1262 26268
rect -1242 26246 -1238 26268
rect -1218 26246 -1214 26268
rect -1194 26246 -1190 26268
rect -1170 26246 -1166 26268
rect -1146 26246 -1142 26268
rect -1122 26246 -1118 26268
rect -1098 26246 -1094 26268
rect -1074 26246 -1070 26268
rect -1050 26246 -1046 26268
rect -1026 26246 -1022 26268
rect -1002 26246 -998 26268
rect -978 26246 -974 26268
rect -954 26246 -950 26268
rect -930 26246 -926 26268
rect -906 26246 -902 26268
rect -882 26246 -878 26268
rect -858 26246 -854 26268
rect -834 26246 -830 26268
rect -810 26246 -806 26268
rect -786 26246 -782 26268
rect -762 26246 -758 26268
rect -738 26246 -734 26268
rect -714 26267 -710 26268
rect -2393 26244 -717 26246
rect -2371 26222 -2366 26244
rect -2348 26222 -2343 26244
rect -2325 26236 -2317 26244
rect -2079 26241 -2018 26244
rect -2003 26243 -1966 26244
rect -2000 26242 -1982 26243
rect -2000 26241 -1992 26242
rect -2084 26237 -2009 26241
rect -2028 26236 -2009 26237
rect -2000 26237 -1854 26241
rect -1846 26237 -1798 26244
rect -2325 26222 -2320 26236
rect -2309 26224 -2301 26236
rect -2028 26234 -2018 26236
rect -2092 26224 -2084 26231
rect -2023 26227 -2014 26234
rect -2000 26227 -1992 26237
rect -1671 26236 -1663 26244
rect -1846 26233 -1806 26235
rect -1854 26227 -1806 26231
rect -2054 26224 -1806 26227
rect -1655 26224 -1647 26236
rect -2317 26222 -2309 26224
rect -2054 26222 -2024 26224
rect -2000 26222 -1992 26224
rect -1663 26222 -1655 26224
rect -1642 26222 -1637 26244
rect -1619 26222 -1614 26244
rect -1530 26222 -1526 26244
rect -1506 26222 -1502 26244
rect -1482 26222 -1478 26244
rect -1458 26222 -1454 26244
rect -1434 26222 -1430 26244
rect -1410 26222 -1406 26244
rect -1386 26222 -1382 26244
rect -1362 26222 -1358 26244
rect -1338 26222 -1334 26244
rect -1314 26222 -1310 26244
rect -1290 26222 -1286 26244
rect -1266 26222 -1262 26244
rect -1242 26222 -1238 26244
rect -1218 26222 -1214 26244
rect -1194 26222 -1190 26244
rect -1170 26222 -1166 26244
rect -1146 26222 -1142 26244
rect -1122 26222 -1118 26244
rect -1098 26222 -1094 26244
rect -1074 26222 -1070 26244
rect -1050 26222 -1046 26244
rect -1026 26222 -1022 26244
rect -1002 26222 -998 26244
rect -978 26222 -974 26244
rect -954 26222 -950 26244
rect -930 26222 -926 26244
rect -906 26222 -902 26244
rect -882 26222 -878 26244
rect -858 26222 -854 26244
rect -834 26222 -830 26244
rect -810 26222 -806 26244
rect -786 26222 -782 26244
rect -762 26222 -758 26244
rect -738 26222 -734 26244
rect -731 26243 -717 26244
rect -714 26243 -707 26267
rect -714 26222 -710 26243
rect -690 26222 -686 26268
rect -666 26222 -662 26268
rect -642 26222 -638 26268
rect -618 26222 -614 26268
rect -594 26222 -590 26268
rect -570 26222 -566 26268
rect -557 26237 -552 26247
rect -546 26237 -542 26268
rect -547 26223 -542 26237
rect -546 26222 -542 26223
rect -522 26222 -518 26268
rect -498 26222 -494 26268
rect -474 26222 -470 26268
rect -450 26222 -446 26268
rect -426 26222 -422 26268
rect -402 26222 -398 26268
rect -378 26222 -374 26268
rect -354 26222 -350 26268
rect -330 26222 -326 26268
rect -306 26222 -302 26268
rect -282 26222 -278 26268
rect -258 26222 -254 26268
rect -234 26222 -230 26268
rect -210 26222 -206 26268
rect -186 26222 -182 26268
rect -162 26222 -158 26268
rect -138 26222 -134 26268
rect -114 26222 -110 26268
rect -90 26222 -86 26268
rect -77 26261 -72 26268
rect -67 26247 -62 26261
rect -66 26222 -62 26247
rect -42 26222 -38 26316
rect -18 26222 -14 26316
rect 6 26222 10 26316
rect 30 26222 34 26316
rect 54 26222 58 26316
rect 78 26222 82 26316
rect 102 26222 106 26316
rect 126 26222 130 26316
rect 150 26222 154 26316
rect 174 26222 178 26316
rect 198 26222 202 26316
rect 222 26222 226 26316
rect 246 26222 250 26316
rect 270 26222 274 26316
rect 294 26222 298 26316
rect 318 26222 322 26316
rect 342 26222 346 26316
rect 366 26222 370 26316
rect 390 26222 394 26316
rect 414 26222 418 26316
rect 438 26222 442 26316
rect 462 26222 466 26316
rect 486 26222 490 26316
rect 510 26222 514 26316
rect 534 26222 538 26316
rect 558 26222 562 26316
rect 582 26222 586 26316
rect 606 26222 610 26316
rect 630 26222 634 26316
rect 654 26222 658 26316
rect 678 26222 682 26316
rect 702 26222 706 26316
rect 726 26222 730 26316
rect 750 26222 754 26316
rect 774 26222 778 26316
rect 798 26222 802 26316
rect 822 26222 826 26316
rect 846 26222 850 26316
rect 870 26222 874 26316
rect 894 26222 898 26316
rect 918 26222 922 26316
rect 942 26222 946 26316
rect 966 26222 970 26316
rect 990 26222 994 26316
rect 1014 26222 1018 26316
rect 1038 26222 1042 26316
rect 1062 26223 1066 26316
rect 1051 26222 1085 26223
rect -2393 26220 -2064 26222
rect -2060 26220 1085 26222
rect -2371 26174 -2366 26220
rect -2348 26174 -2343 26220
rect -2325 26208 -2317 26220
rect -2060 26217 -2054 26220
rect -2084 26210 -2054 26217
rect -2050 26214 -2044 26216
rect -2325 26188 -2320 26208
rect -2064 26206 -2054 26210
rect -2325 26180 -2317 26188
rect -2101 26183 -2071 26186
rect -2325 26174 -2320 26180
rect -2317 26174 -2309 26180
rect -2000 26178 -1992 26220
rect -1846 26219 -1806 26220
rect -1846 26210 -1798 26217
rect -1671 26208 -1663 26220
rect -1846 26206 -1806 26208
rect -1854 26192 -1680 26196
rect -1846 26183 -1798 26186
rect -2079 26177 -2043 26178
rect -2007 26177 -1991 26178
rect -2079 26176 -2071 26177
rect -2079 26174 -2029 26176
rect -2011 26174 -1991 26177
rect -1846 26175 -1806 26181
rect -1671 26180 -1663 26188
rect -1864 26174 -1796 26175
rect -1663 26174 -1655 26180
rect -1642 26174 -1637 26220
rect -1619 26174 -1614 26220
rect -1530 26174 -1526 26220
rect -1506 26174 -1502 26220
rect -1482 26174 -1478 26220
rect -1458 26174 -1454 26220
rect -1434 26174 -1430 26220
rect -1410 26174 -1406 26220
rect -1386 26174 -1382 26220
rect -1362 26174 -1358 26220
rect -1338 26174 -1334 26220
rect -1314 26174 -1310 26220
rect -1290 26174 -1286 26220
rect -1266 26174 -1262 26220
rect -1242 26174 -1238 26220
rect -1218 26174 -1214 26220
rect -1194 26174 -1190 26220
rect -1170 26174 -1166 26220
rect -1146 26174 -1142 26220
rect -1122 26174 -1118 26220
rect -1098 26174 -1094 26220
rect -1074 26174 -1070 26220
rect -1050 26174 -1046 26220
rect -1026 26174 -1022 26220
rect -1002 26174 -998 26220
rect -978 26174 -974 26220
rect -954 26174 -950 26220
rect -930 26174 -926 26220
rect -906 26174 -902 26220
rect -882 26174 -878 26220
rect -858 26174 -854 26220
rect -834 26174 -830 26220
rect -810 26174 -806 26220
rect -786 26174 -782 26220
rect -762 26174 -758 26220
rect -738 26174 -734 26220
rect -714 26174 -710 26220
rect -690 26174 -686 26220
rect -666 26174 -662 26220
rect -642 26174 -638 26220
rect -618 26174 -614 26220
rect -594 26174 -590 26220
rect -570 26174 -566 26220
rect -546 26174 -542 26220
rect -522 26174 -518 26220
rect -498 26174 -494 26220
rect -474 26174 -470 26220
rect -461 26189 -456 26199
rect -450 26189 -446 26220
rect -451 26175 -446 26189
rect -450 26174 -446 26175
rect -426 26174 -422 26220
rect -402 26174 -398 26220
rect -378 26174 -374 26220
rect -354 26174 -350 26220
rect -330 26174 -326 26220
rect -306 26174 -302 26220
rect -282 26174 -278 26220
rect -258 26174 -254 26220
rect -234 26174 -230 26220
rect -210 26174 -206 26220
rect -186 26174 -182 26220
rect -162 26174 -158 26220
rect -138 26174 -134 26220
rect -114 26174 -110 26220
rect -90 26174 -86 26220
rect -66 26174 -62 26220
rect -42 26219 -38 26220
rect -2393 26172 -45 26174
rect -2371 26126 -2366 26172
rect -2348 26126 -2343 26172
rect -2325 26160 -2320 26172
rect -2079 26170 -2071 26172
rect -2072 26168 -2071 26170
rect -2109 26163 -2101 26168
rect -2101 26161 -2079 26163
rect -2069 26161 -2068 26168
rect -2325 26152 -2317 26160
rect -2079 26156 -2071 26161
rect -2325 26132 -2320 26152
rect -2317 26144 -2309 26152
rect -2074 26147 -2071 26156
rect -2069 26152 -2068 26156
rect -2109 26138 -2079 26141
rect -2325 26126 -2317 26132
rect -2000 26126 -1992 26172
rect -1846 26170 -1806 26172
rect -1854 26165 -1806 26169
rect -1854 26163 -1846 26165
rect -1846 26161 -1806 26163
rect -1806 26159 -1798 26161
rect -1846 26156 -1798 26159
rect -1846 26143 -1806 26154
rect -1671 26152 -1663 26160
rect -1663 26144 -1655 26152
rect -1854 26138 -1680 26142
rect -1671 26126 -1663 26132
rect -1642 26126 -1637 26172
rect -1619 26126 -1614 26172
rect -1530 26126 -1526 26172
rect -1506 26126 -1502 26172
rect -1482 26126 -1478 26172
rect -1458 26126 -1454 26172
rect -1434 26126 -1430 26172
rect -1410 26126 -1406 26172
rect -1386 26126 -1382 26172
rect -1362 26126 -1358 26172
rect -1338 26126 -1334 26172
rect -1314 26126 -1310 26172
rect -1290 26126 -1286 26172
rect -1266 26126 -1262 26172
rect -1242 26126 -1238 26172
rect -1218 26126 -1214 26172
rect -1194 26126 -1190 26172
rect -1170 26126 -1166 26172
rect -1146 26126 -1142 26172
rect -1122 26126 -1118 26172
rect -1098 26126 -1094 26172
rect -1074 26126 -1070 26172
rect -1050 26126 -1046 26172
rect -1026 26126 -1022 26172
rect -1002 26126 -998 26172
rect -978 26126 -974 26172
rect -954 26126 -950 26172
rect -930 26126 -926 26172
rect -906 26126 -902 26172
rect -882 26126 -878 26172
rect -858 26126 -854 26172
rect -834 26126 -830 26172
rect -810 26126 -806 26172
rect -786 26126 -782 26172
rect -762 26126 -758 26172
rect -738 26126 -734 26172
rect -714 26126 -710 26172
rect -690 26126 -686 26172
rect -666 26126 -662 26172
rect -642 26126 -638 26172
rect -618 26126 -614 26172
rect -594 26126 -590 26172
rect -570 26126 -566 26172
rect -546 26126 -542 26172
rect -522 26171 -518 26172
rect -522 26147 -515 26171
rect -522 26126 -518 26147
rect -498 26126 -494 26172
rect -474 26126 -470 26172
rect -450 26126 -446 26172
rect -426 26126 -422 26172
rect -402 26126 -398 26172
rect -378 26126 -374 26172
rect -354 26126 -350 26172
rect -330 26126 -326 26172
rect -306 26126 -302 26172
rect -282 26126 -278 26172
rect -258 26126 -254 26172
rect -234 26126 -230 26172
rect -210 26126 -206 26172
rect -186 26126 -182 26172
rect -162 26126 -158 26172
rect -138 26126 -134 26172
rect -114 26126 -110 26172
rect -90 26126 -86 26172
rect -66 26126 -62 26172
rect -59 26171 -45 26172
rect -42 26171 -35 26219
rect -42 26126 -38 26171
rect -18 26126 -14 26220
rect 6 26126 10 26220
rect 30 26126 34 26220
rect 54 26126 58 26220
rect 78 26126 82 26220
rect 102 26126 106 26220
rect 126 26126 130 26220
rect 150 26126 154 26220
rect 174 26126 178 26220
rect 198 26126 202 26220
rect 222 26126 226 26220
rect 246 26126 250 26220
rect 270 26126 274 26220
rect 294 26126 298 26220
rect 318 26126 322 26220
rect 342 26126 346 26220
rect 366 26126 370 26220
rect 390 26126 394 26220
rect 414 26126 418 26220
rect 438 26126 442 26220
rect 462 26126 466 26220
rect 486 26126 490 26220
rect 510 26126 514 26220
rect 534 26126 538 26220
rect 558 26126 562 26220
rect 582 26126 586 26220
rect 606 26126 610 26220
rect 630 26126 634 26220
rect 654 26126 658 26220
rect 678 26126 682 26220
rect 702 26126 706 26220
rect 726 26126 730 26220
rect 750 26126 754 26220
rect 774 26126 778 26220
rect 798 26126 802 26220
rect 822 26126 826 26220
rect 846 26126 850 26220
rect 870 26126 874 26220
rect 894 26126 898 26220
rect 918 26126 922 26220
rect 942 26126 946 26220
rect 966 26126 970 26220
rect 990 26126 994 26220
rect 1003 26141 1008 26151
rect 1014 26141 1018 26220
rect 1013 26127 1018 26141
rect 1003 26126 1037 26127
rect -2393 26124 1037 26126
rect -2371 26102 -2366 26124
rect -2348 26102 -2343 26124
rect -2325 26116 -2317 26124
rect -2325 26102 -2320 26116
rect -2309 26104 -2301 26116
rect -2092 26107 -2062 26112
rect -2000 26104 -1992 26124
rect -2317 26102 -2309 26104
rect -2000 26102 -1983 26104
rect -1906 26102 -1904 26124
rect -1806 26116 -1680 26122
rect -1671 26116 -1663 26124
rect -1854 26107 -1806 26112
rect -1846 26102 -1806 26105
rect -1655 26104 -1647 26116
rect -1663 26102 -1655 26104
rect -1642 26102 -1637 26124
rect -1619 26102 -1614 26124
rect -1530 26102 -1526 26124
rect -1506 26102 -1502 26124
rect -1482 26102 -1478 26124
rect -1458 26102 -1454 26124
rect -1434 26102 -1430 26124
rect -1410 26102 -1406 26124
rect -1386 26102 -1382 26124
rect -1362 26102 -1358 26124
rect -1338 26102 -1334 26124
rect -1314 26102 -1310 26124
rect -1290 26102 -1286 26124
rect -1266 26102 -1262 26124
rect -1242 26102 -1238 26124
rect -1218 26102 -1214 26124
rect -1194 26102 -1190 26124
rect -1170 26102 -1166 26124
rect -1146 26102 -1142 26124
rect -1122 26102 -1118 26124
rect -1098 26102 -1094 26124
rect -1074 26102 -1070 26124
rect -1050 26102 -1046 26124
rect -1026 26102 -1022 26124
rect -1002 26102 -998 26124
rect -978 26102 -974 26124
rect -954 26103 -950 26124
rect -965 26102 -931 26103
rect -2393 26100 -931 26102
rect -2371 26078 -2366 26100
rect -2348 26078 -2343 26100
rect -2325 26088 -2317 26100
rect -2071 26096 -2062 26100
rect -2013 26098 -1983 26100
rect -2000 26097 -1983 26098
rect -2325 26078 -2320 26088
rect -2309 26078 -2301 26088
rect -2100 26087 -2092 26094
rect -2064 26092 -2062 26095
rect -2061 26087 -2059 26092
rect -2071 26082 -2062 26087
rect -2071 26080 -2026 26082
rect -2066 26078 -2012 26080
rect -2000 26078 -1992 26097
rect -1906 26095 -1904 26100
rect -1846 26096 -1806 26100
rect -1846 26089 -1798 26094
rect -1806 26087 -1798 26089
rect -1671 26088 -1663 26100
rect -1854 26085 -1846 26087
rect -1854 26080 -1806 26085
rect -1864 26078 -1796 26079
rect -1655 26078 -1647 26088
rect -1642 26078 -1637 26100
rect -1619 26078 -1614 26100
rect -1530 26078 -1526 26100
rect -1506 26078 -1502 26100
rect -1482 26078 -1478 26100
rect -1458 26078 -1454 26100
rect -1434 26078 -1430 26100
rect -1410 26078 -1406 26100
rect -1386 26078 -1382 26100
rect -1362 26078 -1358 26100
rect -1338 26078 -1334 26100
rect -1314 26078 -1310 26100
rect -1290 26078 -1286 26100
rect -1266 26078 -1262 26100
rect -1242 26078 -1238 26100
rect -1218 26078 -1214 26100
rect -1194 26078 -1190 26100
rect -1170 26079 -1166 26100
rect -1181 26078 -1147 26079
rect -2393 26076 -1147 26078
rect -2371 26030 -2366 26076
rect -2348 26030 -2343 26076
rect -2325 26072 -2320 26076
rect -2317 26072 -2309 26076
rect -2325 26060 -2317 26072
rect -2066 26071 -2062 26076
rect -2147 26068 -2134 26070
rect -2292 26062 -2071 26068
rect -2325 26030 -2320 26060
rect -2092 26046 -2062 26048
rect -2094 26042 -2062 26046
rect -2000 26030 -1992 26076
rect -1846 26069 -1806 26076
rect -1663 26072 -1655 26076
rect -1846 26062 -1680 26068
rect -1671 26060 -1663 26072
rect -1854 26046 -1806 26048
rect -1854 26042 -1680 26046
rect -1642 26030 -1637 26076
rect -1619 26030 -1614 26076
rect -1530 26030 -1526 26076
rect -1506 26030 -1502 26076
rect -1482 26030 -1478 26076
rect -1458 26030 -1454 26076
rect -1434 26030 -1430 26076
rect -1410 26030 -1406 26076
rect -1386 26030 -1382 26076
rect -1362 26030 -1358 26076
rect -1338 26030 -1334 26076
rect -1314 26030 -1310 26076
rect -1290 26030 -1286 26076
rect -1266 26030 -1262 26076
rect -1242 26030 -1238 26076
rect -1218 26030 -1214 26076
rect -1194 26030 -1190 26076
rect -1181 26069 -1176 26076
rect -1170 26069 -1166 26076
rect -1171 26055 -1166 26069
rect -1170 26030 -1166 26055
rect -1146 26030 -1142 26100
rect -1122 26030 -1118 26100
rect -1098 26030 -1094 26100
rect -1074 26030 -1070 26100
rect -1050 26030 -1046 26100
rect -1026 26030 -1022 26100
rect -1002 26030 -998 26100
rect -978 26030 -974 26100
rect -965 26093 -960 26100
rect -954 26093 -950 26100
rect -955 26079 -950 26093
rect -954 26030 -950 26079
rect -930 26030 -926 26124
rect -906 26030 -902 26124
rect -882 26030 -878 26124
rect -858 26030 -854 26124
rect -834 26030 -830 26124
rect -810 26030 -806 26124
rect -786 26030 -782 26124
rect -762 26030 -758 26124
rect -738 26030 -734 26124
rect -714 26030 -710 26124
rect -690 26030 -686 26124
rect -666 26030 -662 26124
rect -642 26030 -638 26124
rect -618 26030 -614 26124
rect -594 26030 -590 26124
rect -570 26030 -566 26124
rect -546 26030 -542 26124
rect -522 26030 -518 26124
rect -498 26030 -494 26124
rect -474 26030 -470 26124
rect -450 26030 -446 26124
rect -426 26123 -422 26124
rect -426 26099 -419 26123
rect -426 26030 -422 26099
rect -402 26030 -398 26124
rect -378 26030 -374 26124
rect -354 26030 -350 26124
rect -330 26030 -326 26124
rect -306 26030 -302 26124
rect -282 26030 -278 26124
rect -258 26030 -254 26124
rect -234 26030 -230 26124
rect -210 26030 -206 26124
rect -186 26030 -182 26124
rect -162 26030 -158 26124
rect -138 26030 -134 26124
rect -114 26030 -110 26124
rect -90 26030 -86 26124
rect -66 26030 -62 26124
rect -42 26030 -38 26124
rect -18 26030 -14 26124
rect 6 26030 10 26124
rect 30 26030 34 26124
rect 54 26030 58 26124
rect 78 26030 82 26124
rect 102 26030 106 26124
rect 126 26030 130 26124
rect 150 26030 154 26124
rect 174 26030 178 26124
rect 198 26030 202 26124
rect 222 26030 226 26124
rect 235 26045 240 26055
rect 246 26045 250 26124
rect 245 26031 250 26045
rect 235 26030 269 26031
rect -2393 26028 269 26030
rect -2371 26006 -2366 26028
rect -2348 26006 -2343 26028
rect -2325 26006 -2320 26028
rect -2072 26026 -2036 26027
rect -2072 26020 -2054 26026
rect -2309 26012 -2301 26020
rect -2317 26006 -2309 26012
rect -2092 26011 -2062 26016
rect -2000 26007 -1992 26028
rect -1938 26027 -1906 26028
rect -1920 26026 -1906 26027
rect -1806 26020 -1680 26026
rect -1854 26011 -1806 26016
rect -1655 26012 -1647 26020
rect -1982 26007 -1966 26008
rect -2000 26006 -1966 26007
rect -1846 26006 -1806 26009
rect -1663 26006 -1655 26012
rect -1642 26006 -1637 26028
rect -1619 26006 -1614 26028
rect -1530 26006 -1526 26028
rect -1506 26006 -1502 26028
rect -1482 26006 -1478 26028
rect -1458 26006 -1454 26028
rect -1434 26006 -1430 26028
rect -1410 26006 -1406 26028
rect -1386 26006 -1382 26028
rect -1362 26006 -1358 26028
rect -1338 26006 -1334 26028
rect -1314 26006 -1310 26028
rect -1290 26006 -1286 26028
rect -1266 26006 -1262 26028
rect -1242 26006 -1238 26028
rect -1218 26006 -1214 26028
rect -1194 26006 -1190 26028
rect -1170 26006 -1166 26028
rect -1146 26006 -1142 26028
rect -1122 26006 -1118 26028
rect -1098 26006 -1094 26028
rect -1074 26006 -1070 26028
rect -1050 26006 -1046 26028
rect -1026 26006 -1022 26028
rect -1002 26006 -998 26028
rect -978 26006 -974 26028
rect -954 26006 -950 26028
rect -930 26027 -926 26028
rect -2393 26004 -933 26006
rect -2371 25982 -2366 26004
rect -2348 25982 -2343 26004
rect -2325 25982 -2320 26004
rect -2000 26002 -1966 26004
rect -2309 25984 -2301 25992
rect -2062 25991 -2054 25998
rect -2092 25984 -2084 25991
rect -2062 25984 -2026 25986
rect -2317 25982 -2309 25984
rect -2062 25982 -2012 25984
rect -2000 25982 -1992 26002
rect -1982 26001 -1966 26002
rect -1846 26000 -1806 26004
rect -1846 25993 -1798 25998
rect -1806 25991 -1798 25993
rect -1854 25989 -1846 25991
rect -1854 25984 -1806 25989
rect -1655 25984 -1647 25992
rect -1864 25982 -1796 25983
rect -1663 25982 -1655 25984
rect -1642 25982 -1637 26004
rect -1619 25982 -1614 26004
rect -1530 25982 -1526 26004
rect -1506 25982 -1502 26004
rect -1482 25982 -1478 26004
rect -1458 25982 -1454 26004
rect -1434 25982 -1430 26004
rect -1410 25982 -1406 26004
rect -1386 25982 -1382 26004
rect -1362 25982 -1358 26004
rect -1338 25982 -1334 26004
rect -1314 25982 -1310 26004
rect -1290 25982 -1286 26004
rect -1266 25982 -1262 26004
rect -1242 25982 -1238 26004
rect -1218 25982 -1214 26004
rect -1194 25982 -1190 26004
rect -1170 25983 -1166 26004
rect -1146 26003 -1142 26004
rect -1181 25982 -1149 25983
rect -2393 25980 -1149 25982
rect -2371 25910 -2366 25980
rect -2348 25910 -2343 25980
rect -2325 25910 -2320 25980
rect -2317 25976 -2309 25980
rect -2062 25976 -2054 25980
rect -2154 25972 -2138 25974
rect -2057 25972 -2054 25976
rect -2292 25966 -2054 25972
rect -2052 25966 -2044 25976
rect -2092 25950 -2062 25952
rect -2094 25946 -2062 25950
rect -2309 25916 -2301 25922
rect -2317 25910 -2309 25916
rect -2000 25910 -1992 25980
rect -1846 25973 -1806 25980
rect -1663 25976 -1655 25980
rect -1846 25966 -1680 25972
rect -1854 25950 -1806 25952
rect -1854 25946 -1680 25950
rect -1655 25916 -1647 25922
rect -1663 25910 -1655 25916
rect -1642 25910 -1637 25980
rect -1619 25910 -1614 25980
rect -1530 25910 -1526 25980
rect -1506 25910 -1502 25980
rect -1482 25910 -1478 25980
rect -1458 25910 -1454 25980
rect -1434 25910 -1430 25980
rect -1410 25910 -1406 25980
rect -1386 25910 -1382 25980
rect -1362 25910 -1358 25980
rect -1338 25910 -1334 25980
rect -1314 25910 -1310 25980
rect -1290 25910 -1286 25980
rect -1266 25910 -1262 25980
rect -1242 25910 -1238 25980
rect -1218 25910 -1214 25980
rect -1194 25910 -1190 25980
rect -1181 25973 -1176 25980
rect -1170 25973 -1166 25980
rect -1163 25979 -1149 25980
rect -1146 25979 -1139 26003
rect -1171 25959 -1166 25973
rect -1170 25910 -1166 25959
rect -1146 25910 -1142 25979
rect -1122 25910 -1118 26004
rect -1098 25910 -1094 26004
rect -1074 25910 -1070 26004
rect -1050 25910 -1046 26004
rect -1026 25910 -1022 26004
rect -1002 25910 -998 26004
rect -978 25910 -974 26004
rect -954 25910 -950 26004
rect -947 26003 -933 26004
rect -930 26003 -923 26027
rect -930 25910 -926 26003
rect -906 25910 -902 26028
rect -882 25910 -878 26028
rect -858 25910 -854 26028
rect -834 25910 -830 26028
rect -810 25910 -806 26028
rect -786 25910 -782 26028
rect -762 25910 -758 26028
rect -738 25910 -734 26028
rect -714 25910 -710 26028
rect -690 25910 -686 26028
rect -666 25910 -662 26028
rect -642 25910 -638 26028
rect -618 25910 -614 26028
rect -594 25910 -590 26028
rect -570 25910 -566 26028
rect -546 25910 -542 26028
rect -522 25910 -518 26028
rect -498 25910 -494 26028
rect -474 25910 -470 26028
rect -450 25910 -446 26028
rect -426 25910 -422 26028
rect -402 25910 -398 26028
rect -378 25910 -374 26028
rect -354 25910 -350 26028
rect -330 25910 -326 26028
rect -306 25910 -302 26028
rect -282 25910 -278 26028
rect -258 25910 -254 26028
rect -234 25910 -230 26028
rect -210 25910 -206 26028
rect -186 25910 -182 26028
rect -173 25997 -168 26007
rect -162 25997 -158 26028
rect -163 25983 -158 25997
rect -162 25910 -158 25983
rect -138 25931 -134 26028
rect -2393 25908 -141 25910
rect -2371 25694 -2366 25908
rect -2348 25694 -2343 25908
rect -2325 25846 -2320 25908
rect -2317 25906 -2309 25908
rect -2000 25907 -1966 25908
rect -2000 25906 -1982 25907
rect -1663 25906 -1655 25908
rect -2028 25898 -2018 25900
rect -2309 25888 -2301 25894
rect -2091 25888 -2061 25895
rect -2317 25878 -2309 25888
rect -2044 25886 -2028 25888
rect -2026 25886 -2014 25898
rect -2084 25880 -2061 25886
rect -2044 25884 -2014 25886
rect -2292 25870 -2054 25879
rect -2325 25838 -2317 25846
rect -2325 25818 -2320 25838
rect -2317 25830 -2309 25838
rect -2325 25802 -2317 25818
rect -2325 25786 -2320 25802
rect -2309 25790 -2301 25802
rect -2317 25786 -2309 25790
rect -2103 25786 -2096 25788
rect -2083 25786 -2053 25788
rect -2325 25774 -2317 25786
rect -2103 25777 -2053 25786
rect -2018 25784 -2017 25790
rect -2003 25784 -2002 25786
rect -2026 25780 -2017 25784
rect -2325 25758 -2320 25774
rect -2309 25762 -2301 25774
rect -2017 25770 -2012 25780
rect -2317 25758 -2309 25762
rect -2325 25746 -2317 25758
rect -2325 25726 -2320 25746
rect -2325 25718 -2317 25726
rect -2325 25698 -2320 25718
rect -2317 25710 -2309 25718
rect -2325 25694 -2317 25698
rect -2000 25694 -1992 25906
rect -1982 25905 -1966 25906
rect -1980 25888 -1932 25895
rect -1655 25888 -1647 25894
rect -1846 25870 -1680 25879
rect -1663 25878 -1655 25888
rect -1671 25838 -1663 25846
rect -1663 25830 -1655 25838
rect -1671 25802 -1663 25818
rect -1655 25790 -1647 25802
rect -1972 25786 -1924 25788
rect -1663 25786 -1655 25790
rect -1972 25777 -1922 25786
rect -1671 25774 -1663 25786
rect -1655 25762 -1647 25774
rect -1663 25758 -1655 25762
rect -1671 25746 -1663 25758
rect -1671 25718 -1663 25726
rect -1663 25710 -1655 25718
rect -1671 25694 -1663 25698
rect -1642 25694 -1637 25908
rect -1619 25694 -1614 25908
rect -1530 25694 -1526 25908
rect -1506 25694 -1502 25908
rect -1482 25694 -1478 25908
rect -1458 25694 -1454 25908
rect -1434 25694 -1430 25908
rect -1410 25694 -1406 25908
rect -1386 25694 -1382 25908
rect -1362 25694 -1358 25908
rect -1338 25694 -1334 25908
rect -1314 25694 -1310 25908
rect -1290 25694 -1286 25908
rect -1266 25694 -1262 25908
rect -1242 25694 -1238 25908
rect -1218 25694 -1214 25908
rect -1194 25694 -1190 25908
rect -1170 25694 -1166 25908
rect -1146 25907 -1142 25908
rect -1146 25883 -1139 25907
rect -1146 25694 -1142 25883
rect -1122 25694 -1118 25908
rect -1098 25694 -1094 25908
rect -1074 25694 -1070 25908
rect -1050 25694 -1046 25908
rect -1026 25694 -1022 25908
rect -1002 25694 -998 25908
rect -978 25694 -974 25908
rect -954 25694 -950 25908
rect -930 25694 -926 25908
rect -906 25694 -902 25908
rect -882 25694 -878 25908
rect -858 25694 -854 25908
rect -834 25694 -830 25908
rect -810 25694 -806 25908
rect -786 25694 -782 25908
rect -762 25694 -758 25908
rect -738 25694 -734 25908
rect -725 25853 -720 25863
rect -714 25853 -710 25908
rect -715 25839 -710 25853
rect -714 25694 -710 25839
rect -690 25787 -686 25908
rect -690 25763 -683 25787
rect -690 25694 -686 25763
rect -666 25694 -662 25908
rect -642 25694 -638 25908
rect -618 25694 -614 25908
rect -594 25694 -590 25908
rect -570 25694 -566 25908
rect -546 25694 -542 25908
rect -522 25694 -518 25908
rect -498 25694 -494 25908
rect -474 25694 -470 25908
rect -450 25694 -446 25908
rect -426 25694 -422 25908
rect -402 25694 -398 25908
rect -378 25694 -374 25908
rect -354 25694 -350 25908
rect -330 25694 -326 25908
rect -306 25694 -302 25908
rect -293 25733 -288 25743
rect -282 25733 -278 25908
rect -283 25719 -278 25733
rect -282 25694 -278 25719
rect -258 25694 -254 25908
rect -234 25694 -230 25908
rect -210 25694 -206 25908
rect -186 25694 -182 25908
rect -162 25694 -158 25908
rect -155 25907 -141 25908
rect -138 25907 -131 25931
rect -138 25694 -134 25907
rect -114 25694 -110 26028
rect -90 25694 -86 26028
rect -66 25694 -62 26028
rect -42 25694 -38 26028
rect -18 25694 -14 26028
rect 6 25694 10 26028
rect 30 25694 34 26028
rect 54 25694 58 26028
rect 67 25709 72 25719
rect 78 25709 82 26028
rect 77 25695 82 25709
rect 67 25694 101 25695
rect -2393 25692 101 25694
rect -2371 25646 -2366 25692
rect -2348 25646 -2343 25692
rect -2325 25684 -2317 25692
rect -2018 25691 -2004 25692
rect -2000 25691 -1992 25692
rect -2072 25690 -1928 25691
rect -2072 25684 -2053 25690
rect -2325 25668 -2320 25684
rect -2317 25682 -2309 25684
rect -2309 25670 -2301 25682
rect -2092 25675 -2062 25680
rect -2317 25668 -2309 25670
rect -2325 25656 -2317 25668
rect -2098 25662 -2096 25673
rect -2092 25662 -2084 25675
rect -2000 25674 -1992 25690
rect -1972 25684 -1928 25690
rect -1924 25684 -1918 25692
rect -1671 25684 -1663 25692
rect -1663 25682 -1655 25684
rect -2083 25664 -2062 25673
rect -2027 25672 -1992 25674
rect -2018 25664 -2002 25672
rect -2000 25664 -1992 25672
rect -2100 25657 -2096 25662
rect -2083 25657 -2053 25662
rect -2003 25660 -1990 25664
rect -1972 25662 -1964 25671
rect -1928 25670 -1924 25673
rect -1655 25670 -1647 25682
rect -1663 25668 -1655 25670
rect -2325 25646 -2320 25656
rect -2317 25654 -2309 25656
rect -2309 25646 -2301 25654
rect -2004 25650 -2003 25660
rect -2062 25646 -2012 25648
rect -2000 25646 -1992 25660
rect -1972 25657 -1924 25662
rect -1864 25657 -1796 25663
rect -1671 25656 -1663 25668
rect -1663 25654 -1655 25656
rect -1864 25646 -1796 25647
rect -1655 25646 -1647 25654
rect -1642 25646 -1637 25692
rect -1619 25646 -1614 25692
rect -1530 25646 -1526 25692
rect -1506 25646 -1502 25692
rect -1482 25646 -1478 25692
rect -1458 25646 -1454 25692
rect -1434 25646 -1430 25692
rect -1410 25646 -1406 25692
rect -1386 25646 -1382 25692
rect -1362 25646 -1358 25692
rect -1338 25646 -1334 25692
rect -1314 25646 -1310 25692
rect -1290 25646 -1286 25692
rect -1266 25646 -1262 25692
rect -1242 25646 -1238 25692
rect -1218 25646 -1214 25692
rect -1194 25646 -1190 25692
rect -1170 25647 -1166 25692
rect -1181 25646 -1147 25647
rect -2393 25644 -1147 25646
rect -2371 25598 -2366 25644
rect -2348 25598 -2343 25644
rect -2325 25640 -2320 25644
rect -2309 25642 -2301 25644
rect -2317 25640 -2309 25642
rect -2325 25628 -2317 25640
rect -2325 25598 -2320 25628
rect -2317 25626 -2309 25628
rect -2092 25614 -2062 25616
rect -2094 25610 -2062 25614
rect -2000 25598 -1992 25644
rect -1655 25642 -1647 25644
rect -1663 25640 -1655 25642
rect -1671 25628 -1663 25640
rect -1663 25626 -1655 25628
rect -1854 25614 -1806 25616
rect -1854 25610 -1680 25614
rect -1642 25598 -1637 25644
rect -1619 25598 -1614 25644
rect -1530 25598 -1526 25644
rect -1506 25598 -1502 25644
rect -1482 25598 -1478 25644
rect -1458 25598 -1454 25644
rect -1434 25598 -1430 25644
rect -1410 25598 -1406 25644
rect -1386 25598 -1382 25644
rect -1362 25598 -1358 25644
rect -1338 25598 -1334 25644
rect -1314 25598 -1310 25644
rect -1290 25598 -1286 25644
rect -1266 25598 -1262 25644
rect -1242 25598 -1238 25644
rect -1218 25598 -1214 25644
rect -1194 25598 -1190 25644
rect -1181 25637 -1176 25644
rect -1170 25637 -1166 25644
rect -1171 25623 -1166 25637
rect -1181 25613 -1176 25623
rect -1170 25613 -1166 25623
rect -1171 25599 -1166 25613
rect -1181 25598 -1147 25599
rect -2393 25596 -1147 25598
rect -2371 25574 -2366 25596
rect -2348 25574 -2343 25596
rect -2325 25574 -2320 25596
rect -2072 25594 -2036 25595
rect -2072 25588 -2054 25594
rect -2309 25580 -2301 25588
rect -2317 25574 -2309 25580
rect -2092 25579 -2062 25584
rect -2000 25575 -1992 25596
rect -1938 25595 -1906 25596
rect -1920 25594 -1906 25595
rect -1806 25588 -1680 25594
rect -1854 25579 -1806 25584
rect -1655 25580 -1647 25588
rect -1982 25575 -1966 25576
rect -2000 25574 -1966 25575
rect -1846 25574 -1806 25577
rect -1663 25574 -1655 25580
rect -1642 25574 -1637 25596
rect -1619 25574 -1614 25596
rect -1530 25574 -1526 25596
rect -1506 25574 -1502 25596
rect -1482 25574 -1478 25596
rect -1458 25574 -1454 25596
rect -1434 25574 -1430 25596
rect -1410 25574 -1406 25596
rect -1386 25574 -1382 25596
rect -1362 25574 -1358 25596
rect -1338 25574 -1334 25596
rect -1314 25574 -1310 25596
rect -1290 25574 -1286 25596
rect -1266 25574 -1262 25596
rect -1242 25574 -1238 25596
rect -1218 25574 -1214 25596
rect -1194 25574 -1190 25596
rect -1181 25589 -1176 25596
rect -1171 25575 -1166 25589
rect -1170 25574 -1166 25575
rect -1146 25574 -1142 25692
rect -1122 25574 -1118 25692
rect -1098 25574 -1094 25692
rect -1074 25574 -1070 25692
rect -1050 25574 -1046 25692
rect -1026 25574 -1022 25692
rect -1002 25574 -998 25692
rect -978 25574 -974 25692
rect -954 25574 -950 25692
rect -930 25574 -926 25692
rect -906 25574 -902 25692
rect -882 25574 -878 25692
rect -858 25574 -854 25692
rect -834 25574 -830 25692
rect -810 25574 -806 25692
rect -786 25574 -782 25692
rect -762 25574 -758 25692
rect -738 25574 -734 25692
rect -714 25574 -710 25692
rect -690 25574 -686 25692
rect -666 25574 -662 25692
rect -642 25574 -638 25692
rect -618 25574 -614 25692
rect -594 25574 -590 25692
rect -570 25574 -566 25692
rect -546 25574 -542 25692
rect -522 25574 -518 25692
rect -498 25574 -494 25692
rect -474 25574 -470 25692
rect -450 25575 -446 25692
rect -461 25574 -427 25575
rect -2393 25572 -427 25574
rect -2371 25550 -2366 25572
rect -2348 25550 -2343 25572
rect -2325 25550 -2320 25572
rect -2000 25570 -1966 25572
rect -2309 25552 -2301 25560
rect -2062 25559 -2054 25566
rect -2092 25552 -2084 25559
rect -2062 25552 -2026 25554
rect -2317 25550 -2309 25552
rect -2062 25550 -2012 25552
rect -2000 25550 -1992 25570
rect -1982 25569 -1966 25570
rect -1846 25568 -1806 25572
rect -1846 25561 -1798 25566
rect -1806 25559 -1798 25561
rect -1854 25557 -1846 25559
rect -1854 25552 -1806 25557
rect -1655 25552 -1647 25560
rect -1864 25550 -1796 25551
rect -1663 25550 -1655 25552
rect -1642 25550 -1637 25572
rect -1619 25550 -1614 25572
rect -1530 25550 -1526 25572
rect -1506 25550 -1502 25572
rect -1482 25550 -1478 25572
rect -1458 25550 -1454 25572
rect -1434 25550 -1430 25572
rect -1410 25550 -1406 25572
rect -1386 25550 -1382 25572
rect -1362 25550 -1358 25572
rect -1338 25550 -1334 25572
rect -1314 25550 -1310 25572
rect -1290 25550 -1286 25572
rect -1266 25550 -1262 25572
rect -1242 25550 -1238 25572
rect -1218 25550 -1214 25572
rect -1194 25550 -1190 25572
rect -1170 25550 -1166 25572
rect -1146 25571 -1142 25572
rect -2393 25548 -1149 25550
rect -2371 25502 -2366 25548
rect -2348 25502 -2343 25548
rect -2325 25502 -2320 25548
rect -2317 25544 -2309 25548
rect -2062 25544 -2054 25548
rect -2154 25540 -2138 25542
rect -2057 25540 -2054 25544
rect -2292 25534 -2054 25540
rect -2052 25534 -2044 25544
rect -2092 25518 -2062 25520
rect -2094 25514 -2062 25518
rect -2000 25502 -1992 25548
rect -1846 25541 -1806 25548
rect -1663 25544 -1655 25548
rect -1846 25534 -1680 25540
rect -1854 25518 -1806 25520
rect -1854 25514 -1680 25518
rect -1642 25502 -1637 25548
rect -1619 25502 -1614 25548
rect -1530 25502 -1526 25548
rect -1506 25502 -1502 25548
rect -1482 25502 -1478 25548
rect -1458 25502 -1454 25548
rect -1434 25502 -1430 25548
rect -1410 25502 -1406 25548
rect -1386 25502 -1382 25548
rect -1362 25502 -1358 25548
rect -1338 25502 -1334 25548
rect -1314 25502 -1310 25548
rect -1290 25502 -1286 25548
rect -1266 25502 -1262 25548
rect -1242 25502 -1238 25548
rect -1218 25502 -1214 25548
rect -1194 25502 -1190 25548
rect -1170 25502 -1166 25548
rect -1163 25547 -1149 25548
rect -2393 25500 -1149 25502
rect -2371 25478 -2366 25500
rect -2348 25478 -2343 25500
rect -2325 25478 -2320 25500
rect -2072 25498 -2036 25499
rect -2072 25492 -2054 25498
rect -2309 25484 -2301 25492
rect -2317 25478 -2309 25484
rect -2092 25483 -2062 25488
rect -2000 25479 -1992 25500
rect -1938 25499 -1906 25500
rect -1920 25498 -1906 25499
rect -1806 25492 -1680 25498
rect -1854 25483 -1806 25488
rect -1655 25484 -1647 25492
rect -1982 25479 -1966 25480
rect -2000 25478 -1966 25479
rect -1846 25478 -1806 25481
rect -1663 25478 -1655 25484
rect -1642 25478 -1637 25500
rect -1619 25478 -1614 25500
rect -1530 25478 -1526 25500
rect -1506 25478 -1502 25500
rect -1482 25478 -1478 25500
rect -1458 25478 -1454 25500
rect -1434 25478 -1430 25500
rect -1410 25478 -1406 25500
rect -1386 25478 -1382 25500
rect -1362 25478 -1358 25500
rect -1338 25478 -1334 25500
rect -1314 25478 -1310 25500
rect -1290 25478 -1286 25500
rect -1266 25478 -1262 25500
rect -1242 25478 -1238 25500
rect -1218 25478 -1214 25500
rect -1194 25478 -1190 25500
rect -1170 25478 -1166 25500
rect -1163 25499 -1149 25500
rect -1146 25499 -1139 25571
rect -1146 25478 -1142 25499
rect -1122 25478 -1118 25572
rect -1098 25478 -1094 25572
rect -1074 25478 -1070 25572
rect -1050 25478 -1046 25572
rect -1026 25478 -1022 25572
rect -1002 25478 -998 25572
rect -978 25478 -974 25572
rect -954 25478 -950 25572
rect -930 25478 -926 25572
rect -906 25478 -902 25572
rect -882 25478 -878 25572
rect -858 25478 -854 25572
rect -834 25478 -830 25572
rect -810 25478 -806 25572
rect -786 25478 -782 25572
rect -762 25478 -758 25572
rect -738 25478 -734 25572
rect -714 25478 -710 25572
rect -690 25478 -686 25572
rect -666 25478 -662 25572
rect -642 25478 -638 25572
rect -618 25478 -614 25572
rect -594 25478 -590 25572
rect -570 25478 -566 25572
rect -546 25478 -542 25572
rect -522 25478 -518 25572
rect -498 25478 -494 25572
rect -474 25478 -470 25572
rect -461 25565 -456 25572
rect -450 25565 -446 25572
rect -451 25551 -446 25565
rect -450 25478 -446 25551
rect -426 25499 -422 25692
rect -402 25527 -398 25692
rect -413 25526 -379 25527
rect -378 25526 -374 25692
rect -354 25526 -350 25692
rect -330 25526 -326 25692
rect -306 25526 -302 25692
rect -282 25526 -278 25692
rect -258 25667 -254 25692
rect -258 25643 -251 25667
rect -258 25526 -254 25643
rect -234 25526 -230 25692
rect -210 25526 -206 25692
rect -186 25526 -182 25692
rect -162 25526 -158 25692
rect -138 25526 -134 25692
rect -114 25526 -110 25692
rect -90 25526 -86 25692
rect -66 25526 -62 25692
rect -42 25526 -38 25692
rect -18 25526 -14 25692
rect 6 25526 10 25692
rect 30 25526 34 25692
rect 54 25526 58 25692
rect 67 25685 72 25692
rect 77 25671 82 25685
rect 78 25526 82 25671
rect 102 25643 106 26028
rect 102 25622 109 25643
rect 126 25622 130 26028
rect 150 25622 154 26028
rect 174 25622 178 26028
rect 198 25622 202 26028
rect 222 25622 226 26028
rect 235 26021 240 26028
rect 245 26007 250 26021
rect 246 25622 250 26007
rect 270 25979 274 26124
rect 270 25931 277 25979
rect 270 25622 274 25931
rect 294 25622 298 26124
rect 318 25622 322 26124
rect 342 25622 346 26124
rect 366 25622 370 26124
rect 390 25622 394 26124
rect 414 25622 418 26124
rect 438 25622 442 26124
rect 462 25622 466 26124
rect 486 25622 490 26124
rect 510 25622 514 26124
rect 534 25622 538 26124
rect 558 25622 562 26124
rect 582 25622 586 26124
rect 606 25622 610 26124
rect 630 25622 634 26124
rect 654 25622 658 26124
rect 678 25622 682 26124
rect 702 25622 706 26124
rect 726 25622 730 26124
rect 750 25622 754 26124
rect 774 25622 778 26124
rect 798 25622 802 26124
rect 822 25622 826 26124
rect 846 25622 850 26124
rect 870 25622 874 26124
rect 894 25622 898 26124
rect 918 25622 922 26124
rect 942 25622 946 26124
rect 955 25925 960 25935
rect 966 25925 970 26124
rect 965 25911 970 25925
rect 955 25901 960 25911
rect 965 25887 970 25901
rect 966 25622 970 25887
rect 990 25859 994 26124
rect 1003 26117 1008 26124
rect 1013 26103 1018 26117
rect 990 25811 997 25859
rect 990 25622 994 25811
rect 1014 25622 1018 26103
rect 1038 26075 1042 26220
rect 1051 26213 1056 26220
rect 1062 26213 1066 26220
rect 1061 26199 1066 26213
rect 1038 26054 1045 26075
rect 1062 26054 1066 26199
rect 1086 26147 1090 26316
rect 1086 26123 1093 26147
rect 1086 26054 1090 26123
rect 1110 26054 1114 26316
rect 1134 26054 1138 26316
rect 1158 26054 1162 26316
rect 1182 26054 1186 26316
rect 1206 26054 1210 26316
rect 1230 26054 1234 26316
rect 1254 26054 1258 26316
rect 1278 26054 1282 26316
rect 1302 26054 1306 26316
rect 1326 26054 1330 26316
rect 1350 26054 1354 26316
rect 1374 26054 1378 26316
rect 1398 26054 1402 26316
rect 1422 26054 1426 26316
rect 1446 26054 1450 26316
rect 1470 26054 1474 26316
rect 1494 26054 1498 26316
rect 1518 26054 1522 26316
rect 1542 26054 1546 26316
rect 1566 26054 1570 26316
rect 1590 26054 1594 26316
rect 1614 26054 1618 26316
rect 1638 26054 1642 26316
rect 1662 26054 1666 26316
rect 1686 26054 1690 26316
rect 1710 26054 1714 26316
rect 1734 26054 1738 26316
rect 1758 26054 1762 26316
rect 1782 26054 1786 26316
rect 1806 26054 1810 26316
rect 1830 26315 1834 26316
rect 1830 26294 1837 26315
rect 1854 26294 1858 26316
rect 1878 26294 1882 26316
rect 1902 26294 1906 26316
rect 1926 26294 1930 26316
rect 1950 26294 1954 26316
rect 1974 26294 1978 26316
rect 1998 26294 2002 26316
rect 2022 26294 2026 26316
rect 2046 26294 2050 26316
rect 2070 26294 2074 26316
rect 2094 26294 2098 26316
rect 2118 26294 2122 26316
rect 2142 26294 2146 26316
rect 2166 26294 2170 26316
rect 2190 26294 2194 26316
rect 2214 26294 2218 26316
rect 2238 26294 2242 26316
rect 2262 26294 2266 26316
rect 2275 26309 2280 26316
rect 2286 26309 2290 26316
rect 2293 26315 2307 26316
rect 2285 26295 2290 26309
rect 2299 26305 2307 26309
rect 2293 26295 2299 26305
rect 2275 26294 2307 26295
rect 1813 26292 2307 26294
rect 1813 26291 1827 26292
rect 1830 26267 1837 26292
rect 1830 26054 1834 26267
rect 1854 26054 1858 26292
rect 1878 26054 1882 26292
rect 1902 26054 1906 26292
rect 1926 26054 1930 26292
rect 1950 26054 1954 26292
rect 1974 26054 1978 26292
rect 1998 26054 2002 26292
rect 2022 26054 2026 26292
rect 2046 26054 2050 26292
rect 2070 26054 2074 26292
rect 2094 26054 2098 26292
rect 2118 26054 2122 26292
rect 2142 26054 2146 26292
rect 2166 26054 2170 26292
rect 2190 26054 2194 26292
rect 2214 26054 2218 26292
rect 2238 26054 2242 26292
rect 2262 26054 2266 26292
rect 2275 26285 2280 26292
rect 2293 26291 2307 26292
rect 2285 26271 2290 26285
rect 2275 26165 2280 26175
rect 2286 26165 2290 26271
rect 2285 26151 2290 26165
rect 2275 26141 2280 26151
rect 2285 26127 2290 26141
rect 2286 26054 2290 26127
rect 2299 26054 2307 26055
rect 1021 26052 2307 26054
rect 1021 26051 1035 26052
rect 1038 26027 1045 26052
rect 1038 25622 1042 26027
rect 1062 25622 1066 26052
rect 1086 25622 1090 26052
rect 1110 25622 1114 26052
rect 1134 25622 1138 26052
rect 1158 25622 1162 26052
rect 1182 25622 1186 26052
rect 1195 25661 1200 25671
rect 1206 25661 1210 26052
rect 1205 25647 1210 25661
rect 1206 25622 1210 25647
rect 1230 25622 1234 26052
rect 1254 25622 1258 26052
rect 1278 25622 1282 26052
rect 1302 25622 1306 26052
rect 1326 25622 1330 26052
rect 1350 25622 1354 26052
rect 1374 25622 1378 26052
rect 1398 25622 1402 26052
rect 1422 25622 1426 26052
rect 1446 25622 1450 26052
rect 1470 25622 1474 26052
rect 1494 25622 1498 26052
rect 1518 25622 1522 26052
rect 1531 25805 1536 25815
rect 1542 25805 1546 26052
rect 1541 25791 1546 25805
rect 1531 25781 1536 25791
rect 1541 25767 1546 25781
rect 1542 25622 1546 25767
rect 1566 25739 1570 26052
rect 1566 25718 1573 25739
rect 1590 25718 1594 26052
rect 1614 25718 1618 26052
rect 1638 25718 1642 26052
rect 1662 25718 1666 26052
rect 1686 25718 1690 26052
rect 1710 25718 1714 26052
rect 1734 25718 1738 26052
rect 1758 25718 1762 26052
rect 1782 25718 1786 26052
rect 1806 25718 1810 26052
rect 1830 25718 1834 26052
rect 1854 25718 1858 26052
rect 1878 25718 1882 26052
rect 1902 25718 1906 26052
rect 1926 25718 1930 26052
rect 1950 25718 1954 26052
rect 1974 25718 1978 26052
rect 1998 25718 2002 26052
rect 2022 25718 2026 26052
rect 2046 25718 2050 26052
rect 2070 25718 2074 26052
rect 2094 25718 2098 26052
rect 2118 25718 2122 26052
rect 2142 25718 2146 26052
rect 2166 25718 2170 26052
rect 2190 25718 2194 26052
rect 2214 25718 2218 26052
rect 2238 25718 2242 26052
rect 2262 25718 2266 26052
rect 2286 25718 2290 26052
rect 2293 26051 2307 26052
rect 2299 26045 2304 26051
rect 2309 26031 2314 26045
rect 2310 25718 2314 26031
rect 2323 25925 2328 25935
rect 2333 25911 2338 25925
rect 2334 25718 2338 25911
rect 2347 25805 2352 25815
rect 2357 25791 2362 25805
rect 2358 25718 2362 25791
rect 2371 25718 2379 25719
rect 1549 25716 2379 25718
rect 1549 25715 1563 25716
rect 1566 25691 1573 25716
rect 1566 25622 1570 25691
rect 1590 25622 1594 25716
rect 1614 25622 1618 25716
rect 1638 25622 1642 25716
rect 1662 25622 1666 25716
rect 1686 25622 1690 25716
rect 1710 25622 1714 25716
rect 1734 25622 1738 25716
rect 1758 25622 1762 25716
rect 1782 25622 1786 25716
rect 1806 25622 1810 25716
rect 1830 25622 1834 25716
rect 1854 25622 1858 25716
rect 1878 25622 1882 25716
rect 1902 25622 1906 25716
rect 1926 25622 1930 25716
rect 1950 25622 1954 25716
rect 1974 25622 1978 25716
rect 1998 25622 2002 25716
rect 2022 25622 2026 25716
rect 2046 25622 2050 25716
rect 2070 25622 2074 25716
rect 2094 25622 2098 25716
rect 2118 25622 2122 25716
rect 2142 25622 2146 25716
rect 2166 25622 2170 25716
rect 2190 25622 2194 25716
rect 2214 25622 2218 25716
rect 2238 25622 2242 25716
rect 2262 25622 2266 25716
rect 2286 25622 2290 25716
rect 2310 25622 2314 25716
rect 2334 25622 2338 25716
rect 2358 25622 2362 25716
rect 2365 25715 2379 25716
rect 2371 25709 2376 25715
rect 2381 25695 2386 25709
rect 2382 25622 2386 25695
rect 85 25620 2403 25622
rect 85 25619 99 25620
rect 102 25595 109 25620
rect 102 25526 106 25595
rect 126 25526 130 25620
rect 150 25526 154 25620
rect 174 25526 178 25620
rect 198 25526 202 25620
rect 222 25526 226 25620
rect 246 25526 250 25620
rect 270 25526 274 25620
rect 294 25526 298 25620
rect 318 25526 322 25620
rect 342 25526 346 25620
rect 366 25526 370 25620
rect 390 25526 394 25620
rect 414 25526 418 25620
rect 438 25526 442 25620
rect 462 25526 466 25620
rect 486 25526 490 25620
rect 510 25526 514 25620
rect 534 25526 538 25620
rect 558 25526 562 25620
rect 582 25526 586 25620
rect 606 25526 610 25620
rect 630 25526 634 25620
rect 654 25526 658 25620
rect 678 25526 682 25620
rect 702 25526 706 25620
rect 726 25526 730 25620
rect 750 25526 754 25620
rect 774 25526 778 25620
rect 798 25526 802 25620
rect 822 25526 826 25620
rect 846 25526 850 25620
rect 870 25526 874 25620
rect 894 25526 898 25620
rect 918 25526 922 25620
rect 942 25526 946 25620
rect 966 25526 970 25620
rect 990 25526 994 25620
rect 1014 25526 1018 25620
rect 1038 25526 1042 25620
rect 1062 25526 1066 25620
rect 1086 25526 1090 25620
rect 1110 25526 1114 25620
rect 1134 25526 1138 25620
rect 1158 25526 1162 25620
rect 1182 25526 1186 25620
rect 1206 25526 1210 25620
rect 1230 25595 1234 25620
rect 1230 25571 1237 25595
rect 1230 25526 1234 25571
rect 1254 25526 1258 25620
rect 1278 25526 1282 25620
rect 1302 25526 1306 25620
rect 1326 25526 1330 25620
rect 1350 25526 1354 25620
rect 1374 25526 1378 25620
rect 1398 25526 1402 25620
rect 1422 25526 1426 25620
rect 1446 25526 1450 25620
rect 1470 25526 1474 25620
rect 1494 25526 1498 25620
rect 1518 25526 1522 25620
rect 1542 25526 1546 25620
rect 1566 25526 1570 25620
rect 1590 25526 1594 25620
rect 1614 25526 1618 25620
rect 1638 25526 1642 25620
rect 1662 25526 1666 25620
rect 1686 25526 1690 25620
rect 1710 25526 1714 25620
rect 1734 25526 1738 25620
rect 1758 25526 1762 25620
rect 1782 25526 1786 25620
rect 1806 25526 1810 25620
rect 1830 25526 1834 25620
rect 1854 25526 1858 25620
rect 1878 25526 1882 25620
rect 1902 25526 1906 25620
rect 1926 25526 1930 25620
rect 1950 25526 1954 25620
rect 1974 25526 1978 25620
rect 1998 25526 2002 25620
rect 2022 25526 2026 25620
rect 2046 25526 2050 25620
rect 2070 25526 2074 25620
rect 2094 25526 2098 25620
rect 2118 25526 2122 25620
rect 2142 25526 2146 25620
rect 2166 25526 2170 25620
rect 2190 25526 2194 25620
rect 2214 25526 2218 25620
rect 2238 25526 2242 25620
rect 2262 25526 2266 25620
rect 2286 25526 2290 25620
rect 2310 25526 2314 25620
rect 2334 25526 2338 25620
rect 2358 25526 2362 25620
rect 2382 25526 2386 25620
rect 2389 25619 2403 25620
rect 2406 25619 2413 25643
rect 2406 25526 2410 25619
rect 2419 25613 2424 25623
rect 2429 25599 2434 25613
rect 2419 25541 2424 25551
rect 2430 25541 2434 25599
rect 2429 25527 2434 25541
rect 2443 25537 2451 25541
rect 2437 25527 2443 25537
rect 2419 25526 2451 25527
rect -413 25524 2451 25526
rect -413 25517 -408 25524
rect -402 25517 -398 25524
rect -403 25503 -398 25517
rect -2393 25476 -429 25478
rect -2371 25454 -2366 25476
rect -2348 25454 -2343 25476
rect -2325 25454 -2320 25476
rect -2000 25474 -1966 25476
rect -2309 25456 -2301 25464
rect -2062 25463 -2054 25470
rect -2092 25456 -2084 25463
rect -2062 25456 -2026 25458
rect -2317 25454 -2309 25456
rect -2062 25454 -2012 25456
rect -2000 25454 -1992 25474
rect -1982 25473 -1966 25474
rect -1846 25472 -1806 25476
rect -1846 25465 -1798 25470
rect -1806 25463 -1798 25465
rect -1854 25461 -1846 25463
rect -1854 25456 -1806 25461
rect -1655 25456 -1647 25464
rect -1864 25454 -1796 25455
rect -1663 25454 -1655 25456
rect -1642 25454 -1637 25476
rect -1619 25454 -1614 25476
rect -1530 25454 -1526 25476
rect -1506 25454 -1502 25476
rect -1482 25454 -1478 25476
rect -1458 25454 -1454 25476
rect -1434 25454 -1430 25476
rect -1410 25454 -1406 25476
rect -1386 25454 -1382 25476
rect -1362 25454 -1358 25476
rect -1338 25454 -1334 25476
rect -1314 25454 -1310 25476
rect -1290 25454 -1286 25476
rect -1266 25454 -1262 25476
rect -1242 25454 -1238 25476
rect -1218 25454 -1214 25476
rect -1194 25454 -1190 25476
rect -1170 25454 -1166 25476
rect -1146 25454 -1142 25476
rect -1122 25454 -1118 25476
rect -1098 25454 -1094 25476
rect -1074 25454 -1070 25476
rect -1050 25454 -1046 25476
rect -1026 25454 -1022 25476
rect -1002 25454 -998 25476
rect -978 25454 -974 25476
rect -954 25454 -950 25476
rect -930 25454 -926 25476
rect -906 25454 -902 25476
rect -882 25454 -878 25476
rect -858 25455 -854 25476
rect -869 25454 -835 25455
rect -2393 25452 -835 25454
rect -2371 25382 -2366 25452
rect -2348 25382 -2343 25452
rect -2325 25382 -2320 25452
rect -2317 25448 -2309 25452
rect -2062 25448 -2054 25452
rect -2154 25444 -2138 25446
rect -2057 25444 -2054 25448
rect -2292 25438 -2054 25444
rect -2052 25438 -2044 25448
rect -2092 25422 -2062 25424
rect -2094 25418 -2062 25422
rect -2309 25388 -2301 25394
rect -2317 25382 -2309 25388
rect -2000 25382 -1992 25452
rect -1846 25445 -1806 25452
rect -1663 25448 -1655 25452
rect -1846 25438 -1680 25444
rect -1854 25422 -1806 25424
rect -1854 25418 -1680 25422
rect -1655 25388 -1647 25394
rect -1663 25382 -1655 25388
rect -1642 25382 -1637 25452
rect -1619 25382 -1614 25452
rect -1530 25382 -1526 25452
rect -1506 25382 -1502 25452
rect -1482 25382 -1478 25452
rect -1458 25382 -1454 25452
rect -1434 25382 -1430 25452
rect -1410 25382 -1406 25452
rect -1386 25382 -1382 25452
rect -1362 25382 -1358 25452
rect -1338 25382 -1334 25452
rect -1314 25382 -1310 25452
rect -1290 25382 -1286 25452
rect -1266 25382 -1262 25452
rect -1242 25382 -1238 25452
rect -1218 25382 -1214 25452
rect -1194 25382 -1190 25452
rect -1170 25382 -1166 25452
rect -1146 25382 -1142 25452
rect -1122 25382 -1118 25452
rect -1098 25382 -1094 25452
rect -1074 25382 -1070 25452
rect -1050 25382 -1046 25452
rect -1026 25382 -1022 25452
rect -1002 25382 -998 25452
rect -978 25382 -974 25452
rect -954 25382 -950 25452
rect -930 25382 -926 25452
rect -906 25382 -902 25452
rect -882 25382 -878 25452
rect -869 25445 -864 25452
rect -858 25445 -854 25452
rect -859 25431 -854 25445
rect -858 25382 -854 25431
rect -834 25382 -830 25476
rect -810 25382 -806 25476
rect -786 25382 -782 25476
rect -762 25382 -758 25476
rect -738 25382 -734 25476
rect -714 25382 -710 25476
rect -690 25382 -686 25476
rect -666 25382 -662 25476
rect -642 25382 -638 25476
rect -618 25382 -614 25476
rect -594 25382 -590 25476
rect -570 25382 -566 25476
rect -546 25382 -542 25476
rect -522 25382 -518 25476
rect -498 25382 -494 25476
rect -474 25382 -470 25476
rect -450 25382 -446 25476
rect -443 25475 -429 25476
rect -426 25475 -419 25499
rect -413 25493 -408 25503
rect -403 25479 -398 25493
rect -426 25382 -422 25475
rect -402 25382 -398 25479
rect -378 25451 -374 25524
rect -378 25403 -371 25451
rect -378 25382 -374 25403
rect -354 25382 -350 25524
rect -330 25382 -326 25524
rect -306 25382 -302 25524
rect -282 25382 -278 25524
rect -258 25382 -254 25524
rect -234 25382 -230 25524
rect -210 25382 -206 25524
rect -186 25382 -182 25524
rect -162 25382 -158 25524
rect -138 25382 -134 25524
rect -114 25382 -110 25524
rect -90 25382 -86 25524
rect -66 25382 -62 25524
rect -42 25382 -38 25524
rect -18 25382 -14 25524
rect 6 25382 10 25524
rect 30 25382 34 25524
rect 54 25382 58 25524
rect 78 25382 82 25524
rect 102 25382 106 25524
rect 115 25469 120 25479
rect 126 25469 130 25524
rect 125 25455 130 25469
rect 126 25382 130 25455
rect 150 25403 154 25524
rect -2393 25380 147 25382
rect -2371 25286 -2366 25380
rect -2348 25286 -2343 25380
rect -2325 25318 -2320 25380
rect -2317 25378 -2309 25380
rect -2000 25379 -1966 25380
rect -2000 25378 -1982 25379
rect -1663 25378 -1655 25380
rect -2028 25370 -2018 25372
rect -2309 25360 -2301 25366
rect -2091 25360 -2061 25367
rect -2317 25350 -2309 25360
rect -2044 25358 -2028 25360
rect -2026 25358 -2014 25370
rect -2084 25352 -2061 25358
rect -2044 25356 -2014 25358
rect -2292 25342 -2054 25351
rect -2325 25310 -2317 25318
rect -2325 25290 -2320 25310
rect -2317 25302 -2309 25310
rect -2325 25286 -2317 25290
rect -2000 25286 -1992 25378
rect -1982 25377 -1966 25378
rect -1980 25360 -1932 25367
rect -1655 25360 -1647 25366
rect -1846 25342 -1680 25351
rect -1663 25350 -1655 25360
rect -1671 25310 -1663 25318
rect -1663 25302 -1655 25310
rect -1671 25286 -1663 25290
rect -1642 25286 -1637 25380
rect -1619 25286 -1614 25380
rect -1530 25286 -1526 25380
rect -1506 25286 -1502 25380
rect -1482 25286 -1478 25380
rect -1469 25325 -1464 25335
rect -1458 25325 -1454 25380
rect -1459 25311 -1454 25325
rect -1458 25286 -1454 25311
rect -1434 25286 -1430 25380
rect -1410 25286 -1406 25380
rect -1386 25286 -1382 25380
rect -1362 25286 -1358 25380
rect -1338 25286 -1334 25380
rect -1314 25286 -1310 25380
rect -1290 25286 -1286 25380
rect -1266 25286 -1262 25380
rect -1242 25286 -1238 25380
rect -1218 25286 -1214 25380
rect -1194 25286 -1190 25380
rect -1170 25286 -1166 25380
rect -1146 25286 -1142 25380
rect -1122 25286 -1118 25380
rect -1098 25286 -1094 25380
rect -1074 25286 -1070 25380
rect -1050 25286 -1046 25380
rect -1026 25286 -1022 25380
rect -1002 25286 -998 25380
rect -978 25286 -974 25380
rect -954 25286 -950 25380
rect -930 25286 -926 25380
rect -906 25286 -902 25380
rect -882 25286 -878 25380
rect -858 25286 -854 25380
rect -834 25379 -830 25380
rect -834 25355 -827 25379
rect -834 25286 -830 25355
rect -810 25286 -806 25380
rect -786 25286 -782 25380
rect -762 25286 -758 25380
rect -738 25286 -734 25380
rect -714 25286 -710 25380
rect -690 25286 -686 25380
rect -666 25286 -662 25380
rect -642 25286 -638 25380
rect -618 25286 -614 25380
rect -594 25286 -590 25380
rect -570 25286 -566 25380
rect -546 25286 -542 25380
rect -522 25286 -518 25380
rect -498 25286 -494 25380
rect -474 25286 -470 25380
rect -450 25286 -446 25380
rect -426 25286 -422 25380
rect -402 25286 -398 25380
rect -378 25286 -374 25380
rect -354 25286 -350 25380
rect -330 25286 -326 25380
rect -306 25286 -302 25380
rect -282 25286 -278 25380
rect -258 25286 -254 25380
rect -234 25286 -230 25380
rect -210 25286 -206 25380
rect -186 25286 -182 25380
rect -162 25286 -158 25380
rect -138 25286 -134 25380
rect -114 25286 -110 25380
rect -90 25286 -86 25380
rect -66 25286 -62 25380
rect -42 25286 -38 25380
rect -18 25286 -14 25380
rect 6 25286 10 25380
rect 30 25286 34 25380
rect 54 25286 58 25380
rect 78 25286 82 25380
rect 102 25286 106 25380
rect 126 25286 130 25380
rect 133 25379 147 25380
rect 150 25379 157 25403
rect 150 25286 154 25379
rect 174 25286 178 25524
rect 198 25286 202 25524
rect 211 25301 216 25311
rect 222 25301 226 25524
rect 221 25287 226 25301
rect 211 25286 245 25287
rect -2393 25284 245 25286
rect -2371 25238 -2366 25284
rect -2348 25238 -2343 25284
rect -2325 25276 -2317 25284
rect -2018 25283 -2004 25284
rect -2000 25283 -1992 25284
rect -2072 25282 -1928 25283
rect -2072 25276 -2053 25282
rect -2325 25260 -2320 25276
rect -2317 25274 -2309 25276
rect -2309 25262 -2301 25274
rect -2092 25267 -2062 25272
rect -2317 25260 -2309 25262
rect -2325 25248 -2317 25260
rect -2098 25254 -2096 25265
rect -2092 25254 -2084 25267
rect -2000 25266 -1992 25282
rect -1972 25276 -1928 25282
rect -1924 25276 -1918 25284
rect -1671 25276 -1663 25284
rect -1663 25274 -1655 25276
rect -2083 25256 -2062 25265
rect -2027 25264 -1992 25266
rect -2018 25256 -2002 25264
rect -2000 25256 -1992 25264
rect -2100 25249 -2096 25254
rect -2083 25249 -2053 25254
rect -2003 25252 -1990 25256
rect -1972 25254 -1964 25263
rect -1928 25262 -1924 25265
rect -1655 25262 -1647 25274
rect -1663 25260 -1655 25262
rect -2325 25238 -2320 25248
rect -2317 25246 -2309 25248
rect -2309 25238 -2301 25246
rect -2004 25242 -2003 25252
rect -2062 25238 -2012 25240
rect -2000 25238 -1992 25252
rect -1972 25249 -1924 25254
rect -1864 25249 -1796 25255
rect -1671 25248 -1663 25260
rect -1663 25246 -1655 25248
rect -1864 25238 -1796 25239
rect -1655 25238 -1647 25246
rect -1642 25238 -1637 25284
rect -1619 25238 -1614 25284
rect -1530 25238 -1526 25284
rect -1506 25238 -1502 25284
rect -1482 25238 -1478 25284
rect -1458 25238 -1454 25284
rect -1434 25259 -1430 25284
rect -2393 25236 -1437 25238
rect -2371 25190 -2366 25236
rect -2348 25190 -2343 25236
rect -2325 25232 -2320 25236
rect -2309 25234 -2301 25236
rect -2317 25232 -2309 25234
rect -2325 25220 -2317 25232
rect -2325 25190 -2320 25220
rect -2317 25218 -2309 25220
rect -2092 25206 -2062 25208
rect -2094 25202 -2062 25206
rect -2000 25190 -1992 25236
rect -1655 25234 -1647 25236
rect -1663 25232 -1655 25234
rect -1671 25220 -1663 25232
rect -1663 25218 -1655 25220
rect -1854 25206 -1806 25208
rect -1854 25202 -1680 25206
rect -1642 25190 -1637 25236
rect -1619 25190 -1614 25236
rect -1530 25190 -1526 25236
rect -1506 25190 -1502 25236
rect -1482 25190 -1478 25236
rect -1458 25190 -1454 25236
rect -1451 25235 -1437 25236
rect -1434 25235 -1427 25259
rect -1434 25190 -1430 25235
rect -1410 25190 -1406 25284
rect -1386 25190 -1382 25284
rect -1373 25253 -1368 25263
rect -1362 25253 -1358 25284
rect -1363 25239 -1358 25253
rect -1362 25190 -1358 25239
rect -1338 25190 -1334 25284
rect -1314 25190 -1310 25284
rect -1290 25190 -1286 25284
rect -1266 25190 -1262 25284
rect -1242 25190 -1238 25284
rect -1218 25190 -1214 25284
rect -1194 25190 -1190 25284
rect -1170 25190 -1166 25284
rect -1146 25190 -1142 25284
rect -1122 25190 -1118 25284
rect -1098 25190 -1094 25284
rect -1074 25190 -1070 25284
rect -1050 25190 -1046 25284
rect -1026 25190 -1022 25284
rect -1002 25190 -998 25284
rect -978 25190 -974 25284
rect -954 25190 -950 25284
rect -930 25190 -926 25284
rect -906 25190 -902 25284
rect -882 25190 -878 25284
rect -858 25190 -854 25284
rect -834 25190 -830 25284
rect -810 25190 -806 25284
rect -786 25190 -782 25284
rect -762 25190 -758 25284
rect -738 25190 -734 25284
rect -714 25190 -710 25284
rect -690 25190 -686 25284
rect -666 25190 -662 25284
rect -642 25190 -638 25284
rect -618 25190 -614 25284
rect -594 25190 -590 25284
rect -570 25190 -566 25284
rect -546 25190 -542 25284
rect -522 25190 -518 25284
rect -498 25190 -494 25284
rect -474 25190 -470 25284
rect -450 25190 -446 25284
rect -426 25190 -422 25284
rect -402 25190 -398 25284
rect -378 25190 -374 25284
rect -354 25190 -350 25284
rect -330 25190 -326 25284
rect -306 25190 -302 25284
rect -282 25190 -278 25284
rect -258 25190 -254 25284
rect -234 25190 -230 25284
rect -210 25190 -206 25284
rect -186 25190 -182 25284
rect -162 25190 -158 25284
rect -138 25190 -134 25284
rect -114 25190 -110 25284
rect -90 25190 -86 25284
rect -66 25190 -62 25284
rect -42 25190 -38 25284
rect -18 25190 -14 25284
rect 6 25190 10 25284
rect 30 25190 34 25284
rect 54 25190 58 25284
rect 78 25190 82 25284
rect 102 25190 106 25284
rect 126 25190 130 25284
rect 150 25190 154 25284
rect 174 25190 178 25284
rect 198 25190 202 25284
rect 211 25277 216 25284
rect 221 25263 226 25277
rect 222 25190 226 25263
rect 246 25235 250 25524
rect -2393 25188 243 25190
rect -2371 25166 -2366 25188
rect -2348 25166 -2343 25188
rect -2325 25166 -2320 25188
rect -2072 25186 -2036 25187
rect -2072 25180 -2054 25186
rect -2309 25172 -2301 25180
rect -2317 25166 -2309 25172
rect -2092 25171 -2062 25176
rect -2000 25167 -1992 25188
rect -1938 25187 -1906 25188
rect -1920 25186 -1906 25187
rect -1806 25180 -1680 25186
rect -1854 25171 -1806 25176
rect -1655 25172 -1647 25180
rect -1982 25167 -1966 25168
rect -2000 25166 -1966 25167
rect -1846 25166 -1806 25169
rect -1663 25166 -1655 25172
rect -1642 25166 -1637 25188
rect -1619 25166 -1614 25188
rect -1530 25166 -1526 25188
rect -1506 25166 -1502 25188
rect -1482 25166 -1478 25188
rect -1458 25166 -1454 25188
rect -1434 25166 -1430 25188
rect -1410 25166 -1406 25188
rect -1386 25166 -1382 25188
rect -1362 25166 -1358 25188
rect -1338 25187 -1334 25188
rect -2393 25164 -1341 25166
rect -2371 25142 -2366 25164
rect -2348 25142 -2343 25164
rect -2325 25142 -2320 25164
rect -2000 25162 -1966 25164
rect -2309 25144 -2301 25152
rect -2062 25151 -2054 25158
rect -2092 25144 -2084 25151
rect -2062 25144 -2026 25146
rect -2317 25142 -2309 25144
rect -2062 25142 -2012 25144
rect -2000 25142 -1992 25162
rect -1982 25161 -1966 25162
rect -1846 25160 -1806 25164
rect -1846 25153 -1798 25158
rect -1806 25151 -1798 25153
rect -1854 25149 -1846 25151
rect -1854 25144 -1806 25149
rect -1655 25144 -1647 25152
rect -1864 25142 -1796 25143
rect -1663 25142 -1655 25144
rect -1642 25142 -1637 25164
rect -1619 25142 -1614 25164
rect -1530 25142 -1526 25164
rect -1506 25142 -1502 25164
rect -1482 25142 -1478 25164
rect -1458 25142 -1454 25164
rect -1434 25142 -1430 25164
rect -1410 25142 -1406 25164
rect -1386 25142 -1382 25164
rect -1362 25142 -1358 25164
rect -1355 25163 -1341 25164
rect -1338 25163 -1331 25187
rect -1338 25142 -1334 25163
rect -1314 25142 -1310 25188
rect -1290 25142 -1286 25188
rect -1277 25157 -1272 25167
rect -1266 25157 -1262 25188
rect -1267 25143 -1262 25157
rect -1266 25142 -1262 25143
rect -1242 25142 -1238 25188
rect -1218 25142 -1214 25188
rect -1194 25142 -1190 25188
rect -1170 25142 -1166 25188
rect -1146 25142 -1142 25188
rect -1122 25142 -1118 25188
rect -1098 25142 -1094 25188
rect -1074 25142 -1070 25188
rect -1050 25142 -1046 25188
rect -1026 25142 -1022 25188
rect -1002 25142 -998 25188
rect -978 25142 -974 25188
rect -954 25142 -950 25188
rect -930 25142 -926 25188
rect -906 25142 -902 25188
rect -882 25142 -878 25188
rect -858 25142 -854 25188
rect -834 25142 -830 25188
rect -810 25142 -806 25188
rect -786 25142 -782 25188
rect -762 25142 -758 25188
rect -738 25142 -734 25188
rect -714 25143 -710 25188
rect -725 25142 -691 25143
rect -2393 25140 -691 25142
rect -2371 25094 -2366 25140
rect -2348 25094 -2343 25140
rect -2325 25094 -2320 25140
rect -2317 25136 -2309 25140
rect -2062 25136 -2054 25140
rect -2154 25132 -2138 25134
rect -2057 25132 -2054 25136
rect -2292 25126 -2054 25132
rect -2052 25126 -2044 25136
rect -2092 25110 -2062 25112
rect -2094 25106 -2062 25110
rect -2000 25094 -1992 25140
rect -1846 25133 -1806 25140
rect -1663 25136 -1655 25140
rect -1846 25126 -1680 25132
rect -1854 25110 -1806 25112
rect -1854 25106 -1680 25110
rect -1642 25094 -1637 25140
rect -1619 25094 -1614 25140
rect -1530 25094 -1526 25140
rect -1506 25094 -1502 25140
rect -1482 25094 -1478 25140
rect -1458 25094 -1454 25140
rect -1434 25094 -1430 25140
rect -1410 25094 -1406 25140
rect -1386 25094 -1382 25140
rect -1362 25094 -1358 25140
rect -1338 25094 -1334 25140
rect -1314 25094 -1310 25140
rect -1290 25094 -1286 25140
rect -1266 25094 -1262 25140
rect -1242 25094 -1238 25140
rect -1218 25094 -1214 25140
rect -1194 25094 -1190 25140
rect -1170 25094 -1166 25140
rect -1146 25094 -1142 25140
rect -1122 25094 -1118 25140
rect -1098 25094 -1094 25140
rect -1074 25094 -1070 25140
rect -1050 25094 -1046 25140
rect -1026 25094 -1022 25140
rect -1002 25094 -998 25140
rect -978 25094 -974 25140
rect -954 25094 -950 25140
rect -930 25094 -926 25140
rect -906 25094 -902 25140
rect -882 25094 -878 25140
rect -858 25094 -854 25140
rect -834 25094 -830 25140
rect -810 25094 -806 25140
rect -786 25094 -782 25140
rect -762 25094 -758 25140
rect -738 25094 -734 25140
rect -725 25133 -720 25140
rect -714 25133 -710 25140
rect -715 25119 -710 25133
rect -714 25094 -710 25119
rect -690 25094 -686 25188
rect -666 25094 -662 25188
rect -642 25094 -638 25188
rect -618 25094 -614 25188
rect -594 25094 -590 25188
rect -570 25094 -566 25188
rect -546 25094 -542 25188
rect -522 25094 -518 25188
rect -498 25094 -494 25188
rect -474 25094 -470 25188
rect -450 25094 -446 25188
rect -426 25094 -422 25188
rect -402 25094 -398 25188
rect -378 25094 -374 25188
rect -354 25094 -350 25188
rect -330 25094 -326 25188
rect -306 25094 -302 25188
rect -282 25094 -278 25188
rect -258 25094 -254 25188
rect -234 25094 -230 25188
rect -210 25094 -206 25188
rect -186 25094 -182 25188
rect -162 25094 -158 25188
rect -138 25094 -134 25188
rect -114 25094 -110 25188
rect -90 25094 -86 25188
rect -66 25094 -62 25188
rect -42 25094 -38 25188
rect -18 25094 -14 25188
rect 6 25094 10 25188
rect 30 25094 34 25188
rect 54 25094 58 25188
rect 78 25094 82 25188
rect 102 25094 106 25188
rect 126 25094 130 25188
rect 150 25094 154 25188
rect 174 25094 178 25188
rect 198 25094 202 25188
rect 222 25094 226 25188
rect 229 25187 243 25188
rect 246 25187 253 25235
rect 246 25094 250 25187
rect 270 25094 274 25524
rect 294 25094 298 25524
rect 318 25094 322 25524
rect 342 25094 346 25524
rect 366 25094 370 25524
rect 390 25094 394 25524
rect 414 25094 418 25524
rect 438 25094 442 25524
rect 462 25094 466 25524
rect 486 25094 490 25524
rect 510 25094 514 25524
rect 534 25094 538 25524
rect 558 25094 562 25524
rect 582 25094 586 25524
rect 606 25094 610 25524
rect 630 25094 634 25524
rect 643 25109 648 25119
rect 654 25109 658 25524
rect 653 25095 658 25109
rect 643 25094 677 25095
rect -2393 25092 677 25094
rect -2371 25070 -2366 25092
rect -2348 25070 -2343 25092
rect -2325 25070 -2320 25092
rect -2072 25090 -2036 25091
rect -2072 25084 -2054 25090
rect -2309 25076 -2301 25084
rect -2317 25070 -2309 25076
rect -2092 25075 -2062 25080
rect -2000 25071 -1992 25092
rect -1938 25091 -1906 25092
rect -1920 25090 -1906 25091
rect -1806 25084 -1680 25090
rect -1854 25075 -1806 25080
rect -1655 25076 -1647 25084
rect -1982 25071 -1966 25072
rect -2000 25070 -1966 25071
rect -1846 25070 -1806 25073
rect -1663 25070 -1655 25076
rect -1642 25070 -1637 25092
rect -1619 25070 -1614 25092
rect -1530 25070 -1526 25092
rect -1506 25070 -1502 25092
rect -1482 25070 -1478 25092
rect -1458 25070 -1454 25092
rect -1434 25070 -1430 25092
rect -1410 25070 -1406 25092
rect -1386 25070 -1382 25092
rect -1362 25070 -1358 25092
rect -1338 25070 -1334 25092
rect -1314 25070 -1310 25092
rect -1290 25070 -1286 25092
rect -1266 25070 -1262 25092
rect -1242 25091 -1238 25092
rect -2393 25068 -1245 25070
rect -2371 25046 -2366 25068
rect -2348 25046 -2343 25068
rect -2325 25046 -2320 25068
rect -2000 25066 -1966 25068
rect -2309 25048 -2301 25056
rect -2062 25055 -2054 25062
rect -2092 25048 -2084 25055
rect -2062 25048 -2026 25050
rect -2317 25046 -2309 25048
rect -2062 25046 -2012 25048
rect -2000 25046 -1992 25066
rect -1982 25065 -1966 25066
rect -1846 25064 -1806 25068
rect -1846 25057 -1798 25062
rect -1806 25055 -1798 25057
rect -1854 25053 -1846 25055
rect -1854 25048 -1806 25053
rect -1655 25048 -1647 25056
rect -1864 25046 -1796 25047
rect -1663 25046 -1655 25048
rect -1642 25046 -1637 25068
rect -1619 25046 -1614 25068
rect -1530 25046 -1526 25068
rect -1506 25046 -1502 25068
rect -1482 25046 -1478 25068
rect -1458 25046 -1454 25068
rect -1434 25046 -1430 25068
rect -1410 25046 -1406 25068
rect -1386 25046 -1382 25068
rect -1362 25046 -1358 25068
rect -1338 25046 -1334 25068
rect -1314 25046 -1310 25068
rect -1290 25046 -1286 25068
rect -1266 25046 -1262 25068
rect -1259 25067 -1245 25068
rect -1242 25067 -1235 25091
rect -1242 25046 -1238 25067
rect -1218 25046 -1214 25092
rect -1194 25046 -1190 25092
rect -1170 25046 -1166 25092
rect -1146 25046 -1142 25092
rect -1122 25046 -1118 25092
rect -1098 25046 -1094 25092
rect -1074 25046 -1070 25092
rect -1050 25046 -1046 25092
rect -1026 25046 -1022 25092
rect -1002 25046 -998 25092
rect -978 25046 -974 25092
rect -954 25046 -950 25092
rect -930 25046 -926 25092
rect -906 25046 -902 25092
rect -882 25046 -878 25092
rect -858 25046 -854 25092
rect -834 25046 -830 25092
rect -810 25046 -806 25092
rect -786 25046 -782 25092
rect -762 25046 -758 25092
rect -738 25046 -734 25092
rect -714 25047 -710 25092
rect -690 25067 -686 25092
rect -725 25046 -693 25047
rect -2393 25044 -693 25046
rect -2371 24998 -2366 25044
rect -2348 24998 -2343 25044
rect -2325 24998 -2320 25044
rect -2317 25040 -2309 25044
rect -2062 25040 -2054 25044
rect -2154 25036 -2138 25038
rect -2057 25036 -2054 25040
rect -2292 25030 -2054 25036
rect -2052 25030 -2044 25040
rect -2092 25014 -2062 25016
rect -2094 25010 -2062 25014
rect -2000 24998 -1992 25044
rect -1846 25037 -1806 25044
rect -1663 25040 -1655 25044
rect -1846 25030 -1680 25036
rect -1854 25014 -1806 25016
rect -1854 25010 -1680 25014
rect -1642 24998 -1637 25044
rect -1619 24998 -1614 25044
rect -1530 24998 -1526 25044
rect -1506 24998 -1502 25044
rect -1482 24998 -1478 25044
rect -1458 24998 -1454 25044
rect -1434 24998 -1430 25044
rect -1410 24998 -1406 25044
rect -1386 24998 -1382 25044
rect -1362 24998 -1358 25044
rect -1338 24998 -1334 25044
rect -1314 24998 -1310 25044
rect -1290 24998 -1286 25044
rect -1266 24998 -1262 25044
rect -1242 24998 -1238 25044
rect -1218 24998 -1214 25044
rect -1194 24998 -1190 25044
rect -1170 24998 -1166 25044
rect -1146 24998 -1142 25044
rect -1122 24998 -1118 25044
rect -1098 24998 -1094 25044
rect -1074 24998 -1070 25044
rect -1050 24998 -1046 25044
rect -1026 24998 -1022 25044
rect -1002 24998 -998 25044
rect -978 24998 -974 25044
rect -954 24998 -950 25044
rect -930 24998 -926 25044
rect -906 24998 -902 25044
rect -882 24998 -878 25044
rect -858 24998 -854 25044
rect -834 24998 -830 25044
rect -810 24998 -806 25044
rect -786 24998 -782 25044
rect -762 24998 -758 25044
rect -738 24998 -734 25044
rect -725 25037 -720 25044
rect -714 25037 -710 25044
rect -707 25043 -693 25044
rect -690 25043 -683 25067
rect -715 25023 -710 25037
rect -714 24998 -710 25023
rect -690 24998 -686 25043
rect -666 24998 -662 25092
rect -642 24998 -638 25092
rect -618 24998 -614 25092
rect -594 24998 -590 25092
rect -570 24998 -566 25092
rect -546 24998 -542 25092
rect -522 24998 -518 25092
rect -498 24998 -494 25092
rect -474 24998 -470 25092
rect -450 24998 -446 25092
rect -426 24998 -422 25092
rect -402 24998 -398 25092
rect -378 24998 -374 25092
rect -354 24998 -350 25092
rect -330 24998 -326 25092
rect -306 24998 -302 25092
rect -282 24998 -278 25092
rect -258 24998 -254 25092
rect -234 24998 -230 25092
rect -210 24998 -206 25092
rect -186 24998 -182 25092
rect -162 24998 -158 25092
rect -138 24998 -134 25092
rect -114 24998 -110 25092
rect -90 24998 -86 25092
rect -66 24998 -62 25092
rect -42 24998 -38 25092
rect -18 24998 -14 25092
rect 6 24998 10 25092
rect 30 24998 34 25092
rect 54 24998 58 25092
rect 78 24998 82 25092
rect 102 24998 106 25092
rect 126 24998 130 25092
rect 150 24998 154 25092
rect 174 24998 178 25092
rect 198 24998 202 25092
rect 222 24998 226 25092
rect 246 24998 250 25092
rect 270 24998 274 25092
rect 294 24998 298 25092
rect 318 24998 322 25092
rect 342 24998 346 25092
rect 366 24998 370 25092
rect 390 24998 394 25092
rect 414 24998 418 25092
rect 438 24998 442 25092
rect 462 24998 466 25092
rect 486 24998 490 25092
rect 510 24998 514 25092
rect 534 24998 538 25092
rect 558 24998 562 25092
rect 582 24998 586 25092
rect 606 24998 610 25092
rect 630 24998 634 25092
rect 643 25085 648 25092
rect 653 25071 658 25085
rect 654 24998 658 25071
rect 678 25043 682 25524
rect -2393 24996 675 24998
rect -2371 24974 -2366 24996
rect -2348 24974 -2343 24996
rect -2325 24974 -2320 24996
rect -2072 24994 -2036 24995
rect -2072 24988 -2054 24994
rect -2309 24980 -2301 24988
rect -2317 24974 -2309 24980
rect -2092 24979 -2062 24984
rect -2000 24975 -1992 24996
rect -1938 24995 -1906 24996
rect -1920 24994 -1906 24995
rect -1806 24988 -1680 24994
rect -1854 24979 -1806 24984
rect -1655 24980 -1647 24988
rect -1982 24975 -1966 24976
rect -2000 24974 -1966 24975
rect -1846 24974 -1806 24977
rect -1663 24974 -1655 24980
rect -1642 24974 -1637 24996
rect -1619 24974 -1614 24996
rect -1530 24974 -1526 24996
rect -1506 24974 -1502 24996
rect -1482 24974 -1478 24996
rect -1458 24974 -1454 24996
rect -1434 24974 -1430 24996
rect -1410 24974 -1406 24996
rect -1386 24974 -1382 24996
rect -1362 24974 -1358 24996
rect -1338 24974 -1334 24996
rect -1314 24974 -1310 24996
rect -1290 24974 -1286 24996
rect -1266 24974 -1262 24996
rect -1242 24974 -1238 24996
rect -1218 24974 -1214 24996
rect -1194 24974 -1190 24996
rect -1170 24974 -1166 24996
rect -1146 24974 -1142 24996
rect -1122 24974 -1118 24996
rect -1098 24974 -1094 24996
rect -1074 24974 -1070 24996
rect -1050 24974 -1046 24996
rect -1026 24974 -1022 24996
rect -1002 24974 -998 24996
rect -978 24974 -974 24996
rect -954 24974 -950 24996
rect -930 24974 -926 24996
rect -906 24974 -902 24996
rect -882 24974 -878 24996
rect -858 24974 -854 24996
rect -834 24974 -830 24996
rect -810 24974 -806 24996
rect -786 24974 -782 24996
rect -762 24974 -758 24996
rect -738 24974 -734 24996
rect -714 24974 -710 24996
rect -690 24974 -686 24996
rect -666 24974 -662 24996
rect -642 24974 -638 24996
rect -618 24974 -614 24996
rect -594 24974 -590 24996
rect -570 24974 -566 24996
rect -546 24974 -542 24996
rect -522 24974 -518 24996
rect -498 24974 -494 24996
rect -474 24974 -470 24996
rect -450 24974 -446 24996
rect -426 24974 -422 24996
rect -402 24974 -398 24996
rect -378 24974 -374 24996
rect -354 24974 -350 24996
rect -330 24974 -326 24996
rect -306 24974 -302 24996
rect -282 24974 -278 24996
rect -258 24974 -254 24996
rect -234 24974 -230 24996
rect -210 24974 -206 24996
rect -186 24974 -182 24996
rect -162 24974 -158 24996
rect -138 24974 -134 24996
rect -114 24974 -110 24996
rect -90 24974 -86 24996
rect -66 24974 -62 24996
rect -42 24974 -38 24996
rect -18 24974 -14 24996
rect 6 24974 10 24996
rect 30 24974 34 24996
rect 54 24974 58 24996
rect 78 24974 82 24996
rect 102 24974 106 24996
rect 126 24974 130 24996
rect 150 24974 154 24996
rect 174 24974 178 24996
rect 198 24974 202 24996
rect 222 24974 226 24996
rect 246 24974 250 24996
rect 270 24974 274 24996
rect 294 24974 298 24996
rect 318 24974 322 24996
rect 342 24974 346 24996
rect 366 24974 370 24996
rect 390 24975 394 24996
rect 379 24974 413 24975
rect -2393 24972 413 24974
rect -2371 24950 -2366 24972
rect -2348 24950 -2343 24972
rect -2325 24950 -2320 24972
rect -2000 24970 -1966 24972
rect -2309 24952 -2301 24960
rect -2062 24959 -2054 24966
rect -2092 24952 -2084 24959
rect -2062 24952 -2026 24954
rect -2317 24950 -2309 24952
rect -2062 24950 -2012 24952
rect -2000 24950 -1992 24970
rect -1982 24969 -1966 24970
rect -1846 24968 -1806 24972
rect -1846 24961 -1798 24966
rect -1806 24959 -1798 24961
rect -1854 24957 -1846 24959
rect -1854 24952 -1806 24957
rect -1655 24952 -1647 24960
rect -1864 24950 -1796 24951
rect -1663 24950 -1655 24952
rect -1642 24950 -1637 24972
rect -1619 24950 -1614 24972
rect -1530 24950 -1526 24972
rect -1506 24950 -1502 24972
rect -1482 24950 -1478 24972
rect -1458 24950 -1454 24972
rect -1434 24950 -1430 24972
rect -1410 24950 -1406 24972
rect -1386 24950 -1382 24972
rect -1362 24950 -1358 24972
rect -1338 24950 -1334 24972
rect -1314 24950 -1310 24972
rect -1290 24950 -1286 24972
rect -1266 24950 -1262 24972
rect -1242 24950 -1238 24972
rect -1218 24950 -1214 24972
rect -1194 24950 -1190 24972
rect -1170 24950 -1166 24972
rect -1146 24950 -1142 24972
rect -1122 24950 -1118 24972
rect -1098 24950 -1094 24972
rect -1074 24950 -1070 24972
rect -1050 24950 -1046 24972
rect -1026 24950 -1022 24972
rect -1002 24950 -998 24972
rect -978 24950 -974 24972
rect -954 24950 -950 24972
rect -930 24950 -926 24972
rect -906 24950 -902 24972
rect -882 24950 -878 24972
rect -858 24950 -854 24972
rect -834 24950 -830 24972
rect -810 24950 -806 24972
rect -786 24950 -782 24972
rect -762 24950 -758 24972
rect -738 24950 -734 24972
rect -714 24951 -710 24972
rect -690 24971 -686 24972
rect -725 24950 -693 24951
rect -2393 24948 -693 24950
rect -2371 24902 -2366 24948
rect -2348 24902 -2343 24948
rect -2325 24902 -2320 24948
rect -2317 24944 -2309 24948
rect -2062 24944 -2054 24948
rect -2154 24940 -2138 24942
rect -2057 24940 -2054 24944
rect -2292 24934 -2054 24940
rect -2052 24934 -2044 24944
rect -2092 24918 -2062 24920
rect -2094 24914 -2062 24918
rect -2000 24902 -1992 24948
rect -1846 24941 -1806 24948
rect -1663 24944 -1655 24948
rect -1846 24934 -1680 24940
rect -1854 24918 -1806 24920
rect -1854 24914 -1680 24918
rect -1642 24902 -1637 24948
rect -1619 24902 -1614 24948
rect -1530 24902 -1526 24948
rect -1506 24902 -1502 24948
rect -1482 24902 -1478 24948
rect -1458 24902 -1454 24948
rect -1434 24902 -1430 24948
rect -1410 24902 -1406 24948
rect -1386 24902 -1382 24948
rect -1362 24902 -1358 24948
rect -1338 24902 -1334 24948
rect -1314 24902 -1310 24948
rect -1290 24902 -1286 24948
rect -1266 24902 -1262 24948
rect -1242 24902 -1238 24948
rect -1218 24902 -1214 24948
rect -1194 24902 -1190 24948
rect -1170 24902 -1166 24948
rect -1146 24902 -1142 24948
rect -1122 24902 -1118 24948
rect -1098 24902 -1094 24948
rect -1074 24902 -1070 24948
rect -1050 24902 -1046 24948
rect -1026 24902 -1022 24948
rect -1002 24902 -998 24948
rect -978 24902 -974 24948
rect -954 24902 -950 24948
rect -930 24902 -926 24948
rect -906 24902 -902 24948
rect -882 24902 -878 24948
rect -858 24902 -854 24948
rect -834 24902 -830 24948
rect -810 24902 -806 24948
rect -786 24902 -782 24948
rect -762 24902 -758 24948
rect -738 24902 -734 24948
rect -725 24941 -720 24948
rect -714 24941 -710 24948
rect -707 24947 -693 24948
rect -690 24947 -683 24971
rect -715 24927 -710 24941
rect -714 24902 -710 24927
rect -690 24902 -686 24947
rect -666 24902 -662 24972
rect -642 24902 -638 24972
rect -618 24902 -614 24972
rect -594 24902 -590 24972
rect -570 24902 -566 24972
rect -546 24902 -542 24972
rect -522 24902 -518 24972
rect -498 24902 -494 24972
rect -474 24902 -470 24972
rect -450 24902 -446 24972
rect -426 24902 -422 24972
rect -402 24902 -398 24972
rect -378 24902 -374 24972
rect -354 24902 -350 24972
rect -330 24902 -326 24972
rect -317 24917 -312 24927
rect -306 24917 -302 24972
rect -307 24903 -302 24917
rect -317 24902 -283 24903
rect -2393 24900 -283 24902
rect -2371 24878 -2366 24900
rect -2348 24878 -2343 24900
rect -2325 24878 -2320 24900
rect -2072 24898 -2036 24899
rect -2072 24892 -2054 24898
rect -2309 24884 -2301 24892
rect -2317 24878 -2309 24884
rect -2092 24883 -2062 24888
rect -2000 24879 -1992 24900
rect -1938 24899 -1906 24900
rect -1920 24898 -1906 24899
rect -1806 24892 -1680 24898
rect -1854 24883 -1806 24888
rect -1655 24884 -1647 24892
rect -1982 24879 -1966 24880
rect -2000 24878 -1966 24879
rect -1846 24878 -1806 24881
rect -1663 24878 -1655 24884
rect -1642 24878 -1637 24900
rect -1619 24878 -1614 24900
rect -1530 24878 -1526 24900
rect -1506 24878 -1502 24900
rect -1482 24878 -1478 24900
rect -1458 24878 -1454 24900
rect -1434 24878 -1430 24900
rect -1410 24878 -1406 24900
rect -1386 24878 -1382 24900
rect -1362 24878 -1358 24900
rect -1338 24878 -1334 24900
rect -1314 24878 -1310 24900
rect -1290 24878 -1286 24900
rect -1266 24878 -1262 24900
rect -1242 24878 -1238 24900
rect -1218 24878 -1214 24900
rect -1194 24878 -1190 24900
rect -1170 24878 -1166 24900
rect -1146 24878 -1142 24900
rect -1122 24878 -1118 24900
rect -1098 24878 -1094 24900
rect -1074 24878 -1070 24900
rect -1050 24878 -1046 24900
rect -1026 24878 -1022 24900
rect -1002 24878 -998 24900
rect -978 24878 -974 24900
rect -954 24878 -950 24900
rect -930 24878 -926 24900
rect -906 24878 -902 24900
rect -882 24878 -878 24900
rect -858 24878 -854 24900
rect -834 24878 -830 24900
rect -810 24878 -806 24900
rect -786 24878 -782 24900
rect -762 24878 -758 24900
rect -738 24878 -734 24900
rect -714 24878 -710 24900
rect -690 24878 -686 24900
rect -666 24878 -662 24900
rect -642 24878 -638 24900
rect -618 24878 -614 24900
rect -594 24878 -590 24900
rect -570 24878 -566 24900
rect -546 24878 -542 24900
rect -522 24878 -518 24900
rect -498 24878 -494 24900
rect -474 24878 -470 24900
rect -450 24878 -446 24900
rect -426 24878 -422 24900
rect -402 24878 -398 24900
rect -378 24878 -374 24900
rect -354 24878 -350 24900
rect -330 24878 -326 24900
rect -317 24893 -312 24900
rect -307 24879 -302 24893
rect -306 24878 -302 24879
rect -282 24878 -278 24972
rect -258 24878 -254 24972
rect -234 24878 -230 24972
rect -210 24878 -206 24972
rect -186 24878 -182 24972
rect -162 24878 -158 24972
rect -138 24878 -134 24972
rect -114 24878 -110 24972
rect -90 24878 -86 24972
rect -66 24878 -62 24972
rect -42 24878 -38 24972
rect -18 24878 -14 24972
rect 6 24878 10 24972
rect 30 24878 34 24972
rect 54 24878 58 24972
rect 78 24878 82 24972
rect 102 24878 106 24972
rect 126 24878 130 24972
rect 150 24878 154 24972
rect 174 24878 178 24972
rect 198 24878 202 24972
rect 222 24878 226 24972
rect 246 24878 250 24972
rect 270 24878 274 24972
rect 294 24878 298 24972
rect 318 24879 322 24972
rect 307 24878 341 24879
rect -2393 24876 341 24878
rect -2371 24854 -2366 24876
rect -2348 24854 -2343 24876
rect -2325 24854 -2320 24876
rect -2000 24874 -1966 24876
rect -2309 24856 -2301 24864
rect -2062 24863 -2054 24870
rect -2092 24856 -2084 24863
rect -2062 24856 -2026 24858
rect -2317 24854 -2309 24856
rect -2062 24854 -2012 24856
rect -2000 24854 -1992 24874
rect -1982 24873 -1966 24874
rect -1846 24872 -1806 24876
rect -1846 24865 -1798 24870
rect -1806 24863 -1798 24865
rect -1854 24861 -1846 24863
rect -1854 24856 -1806 24861
rect -1655 24856 -1647 24864
rect -1864 24854 -1796 24855
rect -1663 24854 -1655 24856
rect -1642 24854 -1637 24876
rect -1619 24854 -1614 24876
rect -1530 24854 -1526 24876
rect -1506 24854 -1502 24876
rect -1482 24854 -1478 24876
rect -1458 24854 -1454 24876
rect -1434 24854 -1430 24876
rect -1410 24854 -1406 24876
rect -1386 24854 -1382 24876
rect -1362 24854 -1358 24876
rect -1338 24854 -1334 24876
rect -1314 24854 -1310 24876
rect -1290 24854 -1286 24876
rect -1266 24854 -1262 24876
rect -1242 24854 -1238 24876
rect -1218 24854 -1214 24876
rect -1194 24854 -1190 24876
rect -1170 24854 -1166 24876
rect -1146 24854 -1142 24876
rect -1122 24854 -1118 24876
rect -1098 24854 -1094 24876
rect -1074 24854 -1070 24876
rect -1050 24854 -1046 24876
rect -1026 24854 -1022 24876
rect -1002 24854 -998 24876
rect -978 24854 -974 24876
rect -954 24854 -950 24876
rect -930 24854 -926 24876
rect -906 24854 -902 24876
rect -882 24854 -878 24876
rect -858 24854 -854 24876
rect -834 24854 -830 24876
rect -810 24854 -806 24876
rect -786 24854 -782 24876
rect -762 24854 -758 24876
rect -738 24854 -734 24876
rect -714 24855 -710 24876
rect -690 24875 -686 24876
rect -725 24854 -693 24855
rect -2393 24852 -693 24854
rect -2371 24806 -2366 24852
rect -2348 24806 -2343 24852
rect -2325 24806 -2320 24852
rect -2317 24848 -2309 24852
rect -2062 24848 -2054 24852
rect -2154 24844 -2138 24846
rect -2057 24844 -2054 24848
rect -2292 24838 -2054 24844
rect -2052 24838 -2044 24848
rect -2092 24822 -2062 24824
rect -2094 24818 -2062 24822
rect -2000 24806 -1992 24852
rect -1846 24845 -1806 24852
rect -1663 24848 -1655 24852
rect -1846 24838 -1680 24844
rect -1854 24822 -1806 24824
rect -1854 24818 -1680 24822
rect -1642 24806 -1637 24852
rect -1619 24806 -1614 24852
rect -1530 24806 -1526 24852
rect -1506 24806 -1502 24852
rect -1482 24806 -1478 24852
rect -1458 24806 -1454 24852
rect -1434 24806 -1430 24852
rect -1410 24806 -1406 24852
rect -1386 24806 -1382 24852
rect -1362 24806 -1358 24852
rect -1338 24806 -1334 24852
rect -1314 24806 -1310 24852
rect -1290 24806 -1286 24852
rect -1266 24806 -1262 24852
rect -1242 24806 -1238 24852
rect -1218 24806 -1214 24852
rect -1194 24806 -1190 24852
rect -1170 24806 -1166 24852
rect -1146 24806 -1142 24852
rect -1122 24806 -1118 24852
rect -1098 24806 -1094 24852
rect -1074 24806 -1070 24852
rect -1050 24806 -1046 24852
rect -1026 24806 -1022 24852
rect -1002 24806 -998 24852
rect -978 24806 -974 24852
rect -954 24806 -950 24852
rect -930 24806 -926 24852
rect -906 24806 -902 24852
rect -882 24806 -878 24852
rect -858 24806 -854 24852
rect -834 24806 -830 24852
rect -810 24806 -806 24852
rect -786 24806 -782 24852
rect -762 24806 -758 24852
rect -738 24806 -734 24852
rect -725 24845 -720 24852
rect -714 24845 -710 24852
rect -707 24851 -693 24852
rect -690 24851 -683 24875
rect -715 24831 -710 24845
rect -714 24806 -710 24831
rect -690 24806 -686 24851
rect -666 24806 -662 24876
rect -642 24806 -638 24876
rect -618 24806 -614 24876
rect -594 24806 -590 24876
rect -570 24806 -566 24876
rect -546 24806 -542 24876
rect -522 24806 -518 24876
rect -498 24806 -494 24876
rect -474 24806 -470 24876
rect -450 24806 -446 24876
rect -426 24806 -422 24876
rect -402 24806 -398 24876
rect -378 24806 -374 24876
rect -354 24806 -350 24876
rect -330 24806 -326 24876
rect -306 24806 -302 24876
rect -282 24851 -278 24876
rect -2393 24804 -285 24806
rect -2371 24758 -2366 24804
rect -2348 24758 -2343 24804
rect -2325 24758 -2320 24804
rect -2309 24788 -2301 24798
rect -2317 24782 -2309 24788
rect -2097 24782 -2095 24791
rect -2309 24760 -2301 24770
rect -2097 24768 -2095 24772
rect -2292 24767 -2095 24768
rect -2097 24765 -2095 24767
rect -2084 24760 -2083 24803
rect -2069 24796 -2054 24798
rect -2054 24780 -2018 24782
rect -2054 24778 -2004 24780
rect -2059 24774 -2045 24778
rect -2054 24772 -2049 24774
rect -2317 24758 -2309 24760
rect -2084 24758 -2054 24760
rect -2044 24758 -2039 24772
rect -2025 24762 -2014 24768
rect -2000 24762 -1992 24804
rect -1920 24802 -1906 24804
rect -1977 24787 -1929 24793
rect -1655 24788 -1647 24798
rect -1977 24777 -1966 24787
rect -1663 24782 -1655 24788
rect -1977 24765 -1929 24767
rect -2033 24758 -1992 24762
rect -1655 24760 -1647 24770
rect -1663 24758 -1655 24760
rect -1642 24758 -1637 24804
rect -1619 24758 -1614 24804
rect -1530 24758 -1526 24804
rect -1506 24758 -1502 24804
rect -1482 24758 -1478 24804
rect -1458 24758 -1454 24804
rect -1434 24758 -1430 24804
rect -1410 24758 -1406 24804
rect -1386 24758 -1382 24804
rect -1362 24758 -1358 24804
rect -1338 24758 -1334 24804
rect -1314 24758 -1310 24804
rect -1290 24758 -1286 24804
rect -1266 24758 -1262 24804
rect -1242 24758 -1238 24804
rect -1218 24758 -1214 24804
rect -1194 24758 -1190 24804
rect -1170 24758 -1166 24804
rect -1146 24758 -1142 24804
rect -1122 24758 -1118 24804
rect -1098 24758 -1094 24804
rect -1074 24758 -1070 24804
rect -1050 24758 -1046 24804
rect -1026 24758 -1022 24804
rect -1002 24758 -998 24804
rect -978 24758 -974 24804
rect -954 24758 -950 24804
rect -930 24758 -926 24804
rect -906 24758 -902 24804
rect -882 24758 -878 24804
rect -858 24758 -854 24804
rect -834 24758 -830 24804
rect -810 24758 -806 24804
rect -786 24758 -782 24804
rect -762 24758 -758 24804
rect -738 24758 -734 24804
rect -714 24758 -710 24804
rect -690 24779 -686 24804
rect -2393 24756 -693 24758
rect -2371 24662 -2366 24756
rect -2348 24662 -2343 24756
rect -2325 24722 -2320 24756
rect -2317 24754 -2309 24756
rect -2084 24743 -2083 24756
rect -2084 24742 -2054 24743
rect -2325 24714 -2317 24722
rect -2325 24694 -2320 24714
rect -2317 24706 -2309 24714
rect -2117 24705 -2095 24715
rect -2045 24712 -2037 24726
rect -2325 24678 -2317 24694
rect -2325 24662 -2320 24678
rect -2309 24666 -2301 24678
rect -2317 24662 -2309 24666
rect -2011 24664 -2001 24666
rect -2000 24664 -1992 24756
rect -1663 24754 -1655 24756
rect -1969 24705 -1929 24717
rect -1671 24714 -1663 24722
rect -1663 24706 -1655 24714
rect -1671 24678 -1663 24694
rect -1655 24666 -1647 24678
rect -2025 24663 -1991 24664
rect -2025 24662 -1975 24663
rect -1852 24662 -1804 24663
rect -1663 24662 -1655 24666
rect -1642 24662 -1637 24756
rect -1619 24662 -1614 24756
rect -1530 24662 -1526 24756
rect -1506 24662 -1502 24756
rect -1482 24662 -1478 24756
rect -1458 24662 -1454 24756
rect -1434 24662 -1430 24756
rect -1410 24662 -1406 24756
rect -1386 24662 -1382 24756
rect -1362 24662 -1358 24756
rect -1338 24662 -1334 24756
rect -1314 24662 -1310 24756
rect -1290 24662 -1286 24756
rect -1266 24662 -1262 24756
rect -1242 24662 -1238 24756
rect -1218 24662 -1214 24756
rect -1194 24662 -1190 24756
rect -1170 24662 -1166 24756
rect -1146 24662 -1142 24756
rect -1122 24662 -1118 24756
rect -1098 24662 -1094 24756
rect -1074 24662 -1070 24756
rect -1050 24662 -1046 24756
rect -1026 24662 -1022 24756
rect -1002 24662 -998 24756
rect -978 24662 -974 24756
rect -954 24662 -950 24756
rect -930 24662 -926 24756
rect -906 24662 -902 24756
rect -882 24662 -878 24756
rect -858 24662 -854 24756
rect -834 24662 -830 24756
rect -810 24662 -806 24756
rect -786 24662 -782 24756
rect -762 24662 -758 24756
rect -738 24662 -734 24756
rect -714 24662 -710 24756
rect -707 24755 -693 24756
rect -690 24755 -683 24779
rect -690 24662 -686 24755
rect -666 24662 -662 24804
rect -642 24662 -638 24804
rect -618 24662 -614 24804
rect -594 24662 -590 24804
rect -570 24662 -566 24804
rect -546 24662 -542 24804
rect -522 24662 -518 24804
rect -498 24662 -494 24804
rect -474 24662 -470 24804
rect -450 24662 -446 24804
rect -426 24662 -422 24804
rect -402 24662 -398 24804
rect -378 24662 -374 24804
rect -354 24662 -350 24804
rect -330 24662 -326 24804
rect -306 24662 -302 24804
rect -299 24803 -285 24804
rect -282 24803 -275 24851
rect -282 24662 -278 24803
rect -258 24662 -254 24876
rect -234 24662 -230 24876
rect -210 24662 -206 24876
rect -186 24662 -182 24876
rect -162 24662 -158 24876
rect -138 24662 -134 24876
rect -114 24662 -110 24876
rect -90 24662 -86 24876
rect -66 24662 -62 24876
rect -42 24662 -38 24876
rect -18 24662 -14 24876
rect 6 24662 10 24876
rect 30 24662 34 24876
rect 54 24662 58 24876
rect 78 24662 82 24876
rect 102 24662 106 24876
rect 126 24662 130 24876
rect 150 24662 154 24876
rect 174 24662 178 24876
rect 198 24662 202 24876
rect 222 24662 226 24876
rect 246 24662 250 24876
rect 270 24662 274 24876
rect 294 24662 298 24876
rect 307 24869 312 24876
rect 318 24869 322 24876
rect 317 24855 322 24869
rect 318 24662 322 24855
rect 342 24803 346 24972
rect 342 24779 349 24803
rect 342 24662 346 24779
rect 366 24662 370 24972
rect 379 24965 384 24972
rect 390 24965 394 24972
rect 389 24951 394 24965
rect 390 24662 394 24951
rect 414 24899 418 24996
rect 414 24875 421 24899
rect 414 24662 418 24875
rect 438 24662 442 24996
rect 462 24662 466 24996
rect 486 24662 490 24996
rect 510 24662 514 24996
rect 534 24662 538 24996
rect 558 24662 562 24996
rect 582 24662 586 24996
rect 606 24662 610 24996
rect 630 24662 634 24996
rect 654 24662 658 24996
rect 661 24995 675 24996
rect 678 24995 685 25043
rect 678 24662 682 24995
rect 702 24662 706 25524
rect 726 24662 730 25524
rect 750 24662 754 25524
rect 774 24662 778 25524
rect 798 24662 802 25524
rect 822 24662 826 25524
rect 846 24662 850 25524
rect 870 24662 874 25524
rect 894 24662 898 25524
rect 918 24662 922 25524
rect 942 24662 946 25524
rect 966 24662 970 25524
rect 990 24662 994 25524
rect 1014 24662 1018 25524
rect 1038 24662 1042 25524
rect 1062 24662 1066 25524
rect 1086 24662 1090 25524
rect 1099 24749 1104 24759
rect 1110 24749 1114 25524
rect 1123 25397 1128 25407
rect 1134 25397 1138 25524
rect 1133 25383 1138 25397
rect 1123 25373 1128 25383
rect 1133 25359 1138 25373
rect 1109 24735 1114 24749
rect 1110 24662 1114 24735
rect 1134 24683 1138 25359
rect 1158 25331 1162 25524
rect 1158 25310 1165 25331
rect 1182 25310 1186 25524
rect 1206 25310 1210 25524
rect 1230 25310 1234 25524
rect 1254 25310 1258 25524
rect 1278 25310 1282 25524
rect 1302 25310 1306 25524
rect 1326 25310 1330 25524
rect 1350 25310 1354 25524
rect 1374 25310 1378 25524
rect 1398 25310 1402 25524
rect 1422 25310 1426 25524
rect 1446 25310 1450 25524
rect 1470 25310 1474 25524
rect 1494 25310 1498 25524
rect 1518 25310 1522 25524
rect 1542 25310 1546 25524
rect 1566 25310 1570 25524
rect 1590 25310 1594 25524
rect 1614 25310 1618 25524
rect 1638 25310 1642 25524
rect 1662 25310 1666 25524
rect 1686 25310 1690 25524
rect 1710 25310 1714 25524
rect 1734 25310 1738 25524
rect 1758 25310 1762 25524
rect 1782 25310 1786 25524
rect 1806 25310 1810 25524
rect 1830 25310 1834 25524
rect 1854 25310 1858 25524
rect 1878 25310 1882 25524
rect 1902 25310 1906 25524
rect 1926 25310 1930 25524
rect 1950 25310 1954 25524
rect 1974 25310 1978 25524
rect 1998 25310 2002 25524
rect 2022 25310 2026 25524
rect 2046 25310 2050 25524
rect 2070 25310 2074 25524
rect 2094 25310 2098 25524
rect 2118 25310 2122 25524
rect 2142 25310 2146 25524
rect 2166 25310 2170 25524
rect 2190 25310 2194 25524
rect 2214 25310 2218 25524
rect 2238 25310 2242 25524
rect 2262 25310 2266 25524
rect 2286 25310 2290 25524
rect 2310 25310 2314 25524
rect 2334 25310 2338 25524
rect 2358 25310 2362 25524
rect 2382 25310 2386 25524
rect 2406 25310 2410 25524
rect 2419 25517 2424 25524
rect 2437 25523 2451 25524
rect 2429 25503 2434 25517
rect 2430 25310 2434 25503
rect 2443 25397 2448 25407
rect 2453 25383 2458 25397
rect 2454 25310 2458 25383
rect 2467 25310 2475 25311
rect 1141 25308 2475 25310
rect 1141 25307 1155 25308
rect 1158 25283 1165 25308
rect -2393 24660 1131 24662
rect -2371 24638 -2366 24660
rect -2348 24638 -2343 24660
rect -2325 24650 -2317 24660
rect -2068 24657 -2038 24660
rect -2040 24652 -2038 24655
rect -2325 24638 -2320 24650
rect -2309 24638 -2301 24650
rect -2042 24638 -2038 24650
rect -2037 24640 -2035 24652
rect -2015 24640 -2011 24654
rect -2037 24638 -2021 24640
rect -2000 24638 -1992 24660
rect -1852 24659 -1804 24660
rect -1969 24650 -1921 24655
rect -1671 24650 -1663 24660
rect -1976 24638 -1940 24639
rect -1655 24638 -1647 24650
rect -1642 24638 -1637 24660
rect -1619 24638 -1614 24660
rect -1530 24638 -1526 24660
rect -1506 24638 -1502 24660
rect -1482 24638 -1478 24660
rect -1458 24638 -1454 24660
rect -1434 24638 -1430 24660
rect -1410 24638 -1406 24660
rect -1386 24638 -1382 24660
rect -1362 24638 -1358 24660
rect -1338 24638 -1334 24660
rect -1314 24638 -1310 24660
rect -1290 24638 -1286 24660
rect -1266 24638 -1262 24660
rect -1242 24638 -1238 24660
rect -1218 24638 -1214 24660
rect -1194 24638 -1190 24660
rect -1170 24638 -1166 24660
rect -1146 24638 -1142 24660
rect -1122 24638 -1118 24660
rect -1098 24638 -1094 24660
rect -1074 24638 -1070 24660
rect -1050 24638 -1046 24660
rect -1026 24638 -1022 24660
rect -1002 24638 -998 24660
rect -978 24638 -974 24660
rect -954 24638 -950 24660
rect -930 24638 -926 24660
rect -906 24638 -902 24660
rect -882 24638 -878 24660
rect -858 24638 -854 24660
rect -834 24638 -830 24660
rect -810 24638 -806 24660
rect -786 24638 -782 24660
rect -762 24638 -758 24660
rect -738 24638 -734 24660
rect -714 24638 -710 24660
rect -690 24638 -686 24660
rect -666 24638 -662 24660
rect -642 24638 -638 24660
rect -618 24638 -614 24660
rect -594 24638 -590 24660
rect -570 24638 -566 24660
rect -546 24638 -542 24660
rect -522 24638 -518 24660
rect -498 24638 -494 24660
rect -474 24638 -470 24660
rect -450 24638 -446 24660
rect -426 24638 -422 24660
rect -402 24638 -398 24660
rect -378 24638 -374 24660
rect -354 24638 -350 24660
rect -330 24638 -326 24660
rect -306 24638 -302 24660
rect -282 24638 -278 24660
rect -258 24638 -254 24660
rect -234 24638 -230 24660
rect -210 24638 -206 24660
rect -186 24638 -182 24660
rect -162 24638 -158 24660
rect -138 24638 -134 24660
rect -114 24638 -110 24660
rect -90 24638 -86 24660
rect -66 24638 -62 24660
rect -42 24638 -38 24660
rect -18 24638 -14 24660
rect 6 24638 10 24660
rect 30 24638 34 24660
rect 54 24638 58 24660
rect 78 24638 82 24660
rect 102 24638 106 24660
rect 126 24638 130 24660
rect 150 24638 154 24660
rect 174 24638 178 24660
rect 198 24638 202 24660
rect 222 24638 226 24660
rect 246 24638 250 24660
rect 270 24638 274 24660
rect 294 24638 298 24660
rect 318 24638 322 24660
rect 342 24638 346 24660
rect 366 24638 370 24660
rect 390 24638 394 24660
rect 414 24638 418 24660
rect 438 24638 442 24660
rect 462 24638 466 24660
rect 486 24638 490 24660
rect 510 24638 514 24660
rect 534 24638 538 24660
rect 558 24638 562 24660
rect 582 24638 586 24660
rect 606 24638 610 24660
rect 630 24638 634 24660
rect 654 24638 658 24660
rect 678 24638 682 24660
rect 702 24638 706 24660
rect 726 24638 730 24660
rect 750 24638 754 24660
rect 774 24638 778 24660
rect 798 24638 802 24660
rect 822 24638 826 24660
rect 846 24638 850 24660
rect 870 24638 874 24660
rect 894 24638 898 24660
rect 918 24638 922 24660
rect 942 24638 946 24660
rect 966 24638 970 24660
rect 990 24638 994 24660
rect 1014 24638 1018 24660
rect 1038 24638 1042 24660
rect 1062 24638 1066 24660
rect 1086 24638 1090 24660
rect 1110 24638 1114 24660
rect 1117 24659 1131 24660
rect 1134 24659 1141 24683
rect 1134 24638 1138 24659
rect 1158 24638 1162 25283
rect 1182 24638 1186 25308
rect 1206 24638 1210 25308
rect 1230 24638 1234 25308
rect 1254 24638 1258 25308
rect 1278 25215 1282 25308
rect 1267 25214 1301 25215
rect 1302 25214 1306 25308
rect 1326 25214 1330 25308
rect 1350 25214 1354 25308
rect 1374 25214 1378 25308
rect 1398 25214 1402 25308
rect 1422 25214 1426 25308
rect 1446 25214 1450 25308
rect 1470 25214 1474 25308
rect 1494 25214 1498 25308
rect 1518 25214 1522 25308
rect 1542 25214 1546 25308
rect 1566 25214 1570 25308
rect 1590 25214 1594 25308
rect 1614 25214 1618 25308
rect 1638 25214 1642 25308
rect 1662 25214 1666 25308
rect 1686 25214 1690 25308
rect 1710 25214 1714 25308
rect 1734 25214 1738 25308
rect 1758 25214 1762 25308
rect 1782 25214 1786 25308
rect 1806 25214 1810 25308
rect 1830 25214 1834 25308
rect 1854 25214 1858 25308
rect 1878 25214 1882 25308
rect 1902 25214 1906 25308
rect 1926 25214 1930 25308
rect 1950 25214 1954 25308
rect 1974 25214 1978 25308
rect 1998 25214 2002 25308
rect 2022 25214 2026 25308
rect 2046 25214 2050 25308
rect 2070 25214 2074 25308
rect 2094 25214 2098 25308
rect 2118 25214 2122 25308
rect 2142 25214 2146 25308
rect 2166 25214 2170 25308
rect 2190 25214 2194 25308
rect 2214 25214 2218 25308
rect 2238 25214 2242 25308
rect 2262 25214 2266 25308
rect 2286 25214 2290 25308
rect 2310 25214 2314 25308
rect 2334 25214 2338 25308
rect 2358 25214 2362 25308
rect 2382 25214 2386 25308
rect 2406 25214 2410 25308
rect 2430 25214 2434 25308
rect 2454 25214 2458 25308
rect 2461 25307 2475 25308
rect 2467 25301 2472 25307
rect 2477 25287 2482 25301
rect 2467 25229 2472 25239
rect 2478 25229 2482 25287
rect 2477 25215 2482 25229
rect 2491 25225 2499 25229
rect 2485 25215 2491 25225
rect 2467 25214 2499 25215
rect 1267 25212 2499 25214
rect 1267 25205 1272 25212
rect 1278 25205 1282 25212
rect 1277 25191 1282 25205
rect 1267 25181 1272 25191
rect 1277 25167 1282 25181
rect 1278 24638 1282 25167
rect 1302 25139 1306 25212
rect 1302 25118 1309 25139
rect 1326 25118 1330 25212
rect 1350 25118 1354 25212
rect 1374 25118 1378 25212
rect 1398 25118 1402 25212
rect 1422 25118 1426 25212
rect 1446 25118 1450 25212
rect 1470 25118 1474 25212
rect 1494 25118 1498 25212
rect 1518 25118 1522 25212
rect 1542 25118 1546 25212
rect 1566 25118 1570 25212
rect 1590 25118 1594 25212
rect 1614 25118 1618 25212
rect 1638 25118 1642 25212
rect 1662 25118 1666 25212
rect 1686 25118 1690 25212
rect 1710 25118 1714 25212
rect 1734 25118 1738 25212
rect 1758 25118 1762 25212
rect 1782 25118 1786 25212
rect 1806 25118 1810 25212
rect 1830 25118 1834 25212
rect 1854 25118 1858 25212
rect 1878 25118 1882 25212
rect 1902 25118 1906 25212
rect 1926 25118 1930 25212
rect 1950 25118 1954 25212
rect 1974 25118 1978 25212
rect 1998 25118 2002 25212
rect 2022 25118 2026 25212
rect 2046 25118 2050 25212
rect 2070 25118 2074 25212
rect 2094 25118 2098 25212
rect 2118 25118 2122 25212
rect 2142 25118 2146 25212
rect 2166 25118 2170 25212
rect 2190 25118 2194 25212
rect 2214 25118 2218 25212
rect 2238 25118 2242 25212
rect 2262 25118 2266 25212
rect 2286 25118 2290 25212
rect 2310 25118 2314 25212
rect 2334 25118 2338 25212
rect 2358 25118 2362 25212
rect 2382 25118 2386 25212
rect 2406 25118 2410 25212
rect 2430 25118 2434 25212
rect 2454 25118 2458 25212
rect 2467 25205 2472 25212
rect 2485 25211 2499 25212
rect 2477 25191 2482 25205
rect 2478 25118 2482 25191
rect 2491 25118 2499 25119
rect 1285 25116 2499 25118
rect 1285 25115 1299 25116
rect 1302 25091 1309 25116
rect 1302 24638 1306 25091
rect 1326 24638 1330 25116
rect 1350 24638 1354 25116
rect 1374 24638 1378 25116
rect 1398 24638 1402 25116
rect 1422 24638 1426 25116
rect 1446 24638 1450 25116
rect 1470 24638 1474 25116
rect 1494 24638 1498 25116
rect 1518 24638 1522 25116
rect 1542 24638 1546 25116
rect 1566 24638 1570 25116
rect 1590 24638 1594 25116
rect 1614 24638 1618 25116
rect 1638 24638 1642 25116
rect 1662 24638 1666 25116
rect 1686 24638 1690 25116
rect 1710 24638 1714 25116
rect 1734 25023 1738 25116
rect 1723 25022 1757 25023
rect 1758 25022 1762 25116
rect 1782 25022 1786 25116
rect 1806 25022 1810 25116
rect 1830 25022 1834 25116
rect 1854 25022 1858 25116
rect 1878 25022 1882 25116
rect 1902 25022 1906 25116
rect 1926 25022 1930 25116
rect 1950 25022 1954 25116
rect 1974 25022 1978 25116
rect 1998 25022 2002 25116
rect 2022 25022 2026 25116
rect 2046 25022 2050 25116
rect 2070 25022 2074 25116
rect 2094 25022 2098 25116
rect 2118 25022 2122 25116
rect 2142 25022 2146 25116
rect 2166 25022 2170 25116
rect 2179 25061 2184 25071
rect 2190 25061 2194 25116
rect 2189 25047 2194 25061
rect 2190 25022 2194 25047
rect 2214 25022 2218 25116
rect 2238 25022 2242 25116
rect 2262 25022 2266 25116
rect 2286 25022 2290 25116
rect 2310 25022 2314 25116
rect 2334 25022 2338 25116
rect 2358 25022 2362 25116
rect 2382 25022 2386 25116
rect 2406 25022 2410 25116
rect 2430 25022 2434 25116
rect 2454 25022 2458 25116
rect 2478 25022 2482 25116
rect 2485 25115 2499 25116
rect 2491 25109 2496 25115
rect 2501 25095 2506 25109
rect 2502 25022 2506 25095
rect 2515 25022 2523 25023
rect 1723 25020 2523 25022
rect 1723 25013 1728 25020
rect 1734 25013 1738 25020
rect 1733 24999 1738 25013
rect 1723 24989 1728 24999
rect 1733 24975 1738 24989
rect 1734 24638 1738 24975
rect 1758 24947 1762 25020
rect 1758 24926 1765 24947
rect 1782 24926 1786 25020
rect 1806 24926 1810 25020
rect 1830 24926 1834 25020
rect 1854 24926 1858 25020
rect 1878 24926 1882 25020
rect 1902 24926 1906 25020
rect 1926 24926 1930 25020
rect 1950 24926 1954 25020
rect 1974 24926 1978 25020
rect 1998 24926 2002 25020
rect 2022 24926 2026 25020
rect 2046 24926 2050 25020
rect 2070 24926 2074 25020
rect 2094 24926 2098 25020
rect 2118 24926 2122 25020
rect 2142 24926 2146 25020
rect 2166 24926 2170 25020
rect 2190 24926 2194 25020
rect 2214 24995 2218 25020
rect 2214 24971 2221 24995
rect 2214 24926 2218 24971
rect 2238 24926 2242 25020
rect 2262 24926 2266 25020
rect 2286 24926 2290 25020
rect 2310 24926 2314 25020
rect 2334 24926 2338 25020
rect 2358 24926 2362 25020
rect 2382 24926 2386 25020
rect 2406 24926 2410 25020
rect 2430 24926 2434 25020
rect 2454 24926 2458 25020
rect 2478 24926 2482 25020
rect 2502 24926 2506 25020
rect 2509 25019 2523 25020
rect 2515 25013 2520 25019
rect 2525 24999 2530 25013
rect 2526 24926 2530 24999
rect 2539 24926 2547 24927
rect 1741 24924 2547 24926
rect 1741 24923 1755 24924
rect 1758 24899 1765 24924
rect 1758 24638 1762 24899
rect 1782 24638 1786 24924
rect 1806 24638 1810 24924
rect 1830 24711 1834 24924
rect 1854 24831 1858 24924
rect 1843 24830 1877 24831
rect 1878 24830 1882 24924
rect 1902 24830 1906 24924
rect 1926 24830 1930 24924
rect 1950 24830 1954 24924
rect 1974 24830 1978 24924
rect 1998 24830 2002 24924
rect 2022 24830 2026 24924
rect 2046 24830 2050 24924
rect 2070 24830 2074 24924
rect 2094 24830 2098 24924
rect 2118 24830 2122 24924
rect 2142 24830 2146 24924
rect 2166 24830 2170 24924
rect 2190 24830 2194 24924
rect 2214 24830 2218 24924
rect 2238 24830 2242 24924
rect 2262 24830 2266 24924
rect 2286 24830 2290 24924
rect 2310 24830 2314 24924
rect 2334 24830 2338 24924
rect 2358 24830 2362 24924
rect 2382 24830 2386 24924
rect 2406 24830 2410 24924
rect 2430 24830 2434 24924
rect 2454 24830 2458 24924
rect 2478 24830 2482 24924
rect 2502 24830 2506 24924
rect 2526 24830 2530 24924
rect 2533 24923 2547 24924
rect 2539 24917 2544 24923
rect 2549 24903 2554 24917
rect 2550 24830 2554 24903
rect 2563 24830 2571 24831
rect 1843 24828 2571 24830
rect 1843 24821 1848 24828
rect 1854 24821 1858 24828
rect 1853 24807 1858 24821
rect 1843 24797 1848 24807
rect 1853 24783 1858 24797
rect 1819 24710 1853 24711
rect 1854 24710 1858 24783
rect 1878 24755 1882 24828
rect 1878 24734 1885 24755
rect 1902 24734 1906 24828
rect 1926 24735 1930 24828
rect 1915 24734 1949 24735
rect 1861 24732 1949 24734
rect 1861 24731 1875 24732
rect 1819 24708 1875 24710
rect 1819 24701 1824 24708
rect 1830 24701 1834 24708
rect 1829 24687 1834 24701
rect 1819 24677 1824 24687
rect 1829 24663 1834 24677
rect 1830 24638 1834 24663
rect 1854 24638 1858 24708
rect 1861 24707 1875 24708
rect 1878 24707 1885 24732
rect 1878 24638 1882 24707
rect 1902 24638 1906 24732
rect 1915 24725 1920 24732
rect 1926 24725 1930 24732
rect 1925 24711 1930 24725
rect 1926 24638 1930 24711
rect 1950 24659 1954 24828
rect -2393 24636 1947 24638
rect -2371 24566 -2366 24636
rect -2348 24566 -2343 24636
rect -2325 24634 -2320 24636
rect -2317 24634 -2309 24636
rect -2325 24622 -2317 24634
rect -2042 24631 -2038 24636
rect -2325 24602 -2320 24622
rect -2325 24594 -2317 24602
rect -2060 24596 -2030 24599
rect -2325 24566 -2320 24594
rect -2317 24586 -2309 24594
rect -2060 24583 -2038 24594
rect -2033 24587 -2030 24596
rect -2028 24592 -2027 24596
rect -2068 24578 -2038 24581
rect -2000 24566 -1992 24636
rect -1969 24630 -1966 24636
rect -1663 24634 -1655 24636
rect -1969 24629 -1921 24630
rect -1902 24629 -1794 24631
rect -1671 24622 -1663 24634
rect -1912 24611 -1884 24613
rect -1852 24605 -1804 24609
rect -1844 24596 -1796 24599
rect -1671 24594 -1663 24602
rect -1844 24583 -1804 24594
rect -1663 24586 -1655 24594
rect -1852 24578 -1680 24582
rect -1979 24566 -1945 24568
rect -1642 24566 -1637 24636
rect -1619 24566 -1614 24636
rect -1530 24566 -1526 24636
rect -1506 24566 -1502 24636
rect -1482 24566 -1478 24636
rect -1458 24566 -1454 24636
rect -1434 24566 -1430 24636
rect -1410 24566 -1406 24636
rect -1386 24566 -1382 24636
rect -1362 24566 -1358 24636
rect -1338 24566 -1334 24636
rect -1314 24566 -1310 24636
rect -1290 24566 -1286 24636
rect -1266 24566 -1262 24636
rect -1242 24566 -1238 24636
rect -1218 24566 -1214 24636
rect -1194 24566 -1190 24636
rect -1170 24566 -1166 24636
rect -1146 24566 -1142 24636
rect -1122 24566 -1118 24636
rect -1098 24566 -1094 24636
rect -1074 24566 -1070 24636
rect -1050 24566 -1046 24636
rect -1026 24566 -1022 24636
rect -1002 24566 -998 24636
rect -978 24566 -974 24636
rect -954 24566 -950 24636
rect -930 24566 -926 24636
rect -906 24566 -902 24636
rect -882 24566 -878 24636
rect -858 24566 -854 24636
rect -834 24566 -830 24636
rect -810 24566 -806 24636
rect -786 24566 -782 24636
rect -762 24566 -758 24636
rect -738 24566 -734 24636
rect -714 24566 -710 24636
rect -690 24566 -686 24636
rect -666 24566 -662 24636
rect -642 24566 -638 24636
rect -618 24566 -614 24636
rect -594 24566 -590 24636
rect -570 24566 -566 24636
rect -546 24566 -542 24636
rect -522 24566 -518 24636
rect -498 24566 -494 24636
rect -474 24566 -470 24636
rect -450 24566 -446 24636
rect -426 24566 -422 24636
rect -402 24566 -398 24636
rect -378 24566 -374 24636
rect -354 24566 -350 24636
rect -330 24566 -326 24636
rect -306 24566 -302 24636
rect -282 24566 -278 24636
rect -258 24566 -254 24636
rect -234 24566 -230 24636
rect -210 24566 -206 24636
rect -186 24566 -182 24636
rect -162 24566 -158 24636
rect -138 24566 -134 24636
rect -114 24566 -110 24636
rect -90 24566 -86 24636
rect -66 24566 -62 24636
rect -42 24566 -38 24636
rect -18 24566 -14 24636
rect 6 24566 10 24636
rect 30 24566 34 24636
rect 54 24566 58 24636
rect 78 24566 82 24636
rect 102 24566 106 24636
rect 126 24566 130 24636
rect 150 24566 154 24636
rect 174 24566 178 24636
rect 198 24566 202 24636
rect 222 24566 226 24636
rect 246 24566 250 24636
rect 270 24566 274 24636
rect 294 24566 298 24636
rect 318 24566 322 24636
rect 342 24566 346 24636
rect 366 24566 370 24636
rect 390 24566 394 24636
rect 414 24566 418 24636
rect 438 24566 442 24636
rect 462 24566 466 24636
rect 486 24566 490 24636
rect 510 24566 514 24636
rect 534 24566 538 24636
rect 558 24566 562 24636
rect 582 24566 586 24636
rect 606 24591 610 24636
rect 595 24590 629 24591
rect 630 24590 634 24636
rect 654 24590 658 24636
rect 678 24590 682 24636
rect 702 24590 706 24636
rect 726 24590 730 24636
rect 750 24590 754 24636
rect 774 24590 778 24636
rect 798 24590 802 24636
rect 822 24590 826 24636
rect 846 24590 850 24636
rect 870 24590 874 24636
rect 894 24590 898 24636
rect 918 24590 922 24636
rect 942 24590 946 24636
rect 966 24590 970 24636
rect 990 24590 994 24636
rect 1014 24590 1018 24636
rect 1038 24590 1042 24636
rect 1062 24590 1066 24636
rect 1086 24590 1090 24636
rect 1110 24590 1114 24636
rect 1134 24590 1138 24636
rect 1158 24590 1162 24636
rect 1182 24590 1186 24636
rect 1206 24590 1210 24636
rect 1230 24590 1234 24636
rect 1254 24590 1258 24636
rect 1278 24590 1282 24636
rect 1302 24590 1306 24636
rect 1326 24590 1330 24636
rect 1350 24590 1354 24636
rect 1374 24590 1378 24636
rect 1398 24590 1402 24636
rect 1422 24590 1426 24636
rect 1446 24590 1450 24636
rect 1470 24590 1474 24636
rect 1494 24590 1498 24636
rect 1518 24590 1522 24636
rect 1542 24590 1546 24636
rect 1566 24590 1570 24636
rect 1590 24590 1594 24636
rect 1614 24590 1618 24636
rect 1638 24590 1642 24636
rect 1662 24590 1666 24636
rect 1686 24590 1690 24636
rect 1710 24590 1714 24636
rect 1734 24590 1738 24636
rect 1758 24590 1762 24636
rect 1782 24590 1786 24636
rect 1806 24590 1810 24636
rect 1830 24590 1834 24636
rect 1854 24635 1858 24636
rect 1854 24614 1861 24635
rect 1878 24614 1882 24636
rect 1902 24614 1906 24636
rect 1926 24614 1930 24636
rect 1933 24635 1947 24636
rect 1950 24635 1957 24659
rect 1950 24614 1954 24635
rect 1974 24614 1978 24828
rect 1998 24614 2002 24828
rect 2022 24614 2026 24828
rect 2046 24614 2050 24828
rect 2070 24614 2074 24828
rect 2094 24614 2098 24828
rect 2118 24614 2122 24828
rect 2142 24614 2146 24828
rect 2166 24614 2170 24828
rect 2190 24614 2194 24828
rect 2214 24614 2218 24828
rect 2238 24614 2242 24828
rect 2262 24614 2266 24828
rect 2286 24614 2290 24828
rect 2310 24614 2314 24828
rect 2334 24614 2338 24828
rect 2358 24614 2362 24828
rect 2382 24614 2386 24828
rect 2406 24614 2410 24828
rect 2430 24614 2434 24828
rect 2454 24614 2458 24828
rect 2478 24614 2482 24828
rect 2502 24614 2506 24828
rect 2526 24614 2530 24828
rect 2550 24615 2554 24828
rect 2557 24827 2571 24828
rect 2563 24821 2568 24827
rect 2573 24807 2578 24821
rect 2563 24629 2568 24639
rect 2574 24629 2578 24807
rect 2587 24701 2592 24711
rect 2597 24687 2602 24701
rect 2587 24653 2592 24663
rect 2598 24653 2602 24687
rect 2597 24639 2602 24653
rect 2573 24615 2578 24629
rect 2539 24614 2573 24615
rect 1837 24612 2573 24614
rect 1837 24611 1851 24612
rect 595 24588 1851 24590
rect 595 24581 600 24588
rect 606 24581 610 24588
rect 605 24567 610 24581
rect 595 24566 629 24567
rect -2393 24564 629 24566
rect -2371 24518 -2366 24564
rect -2348 24518 -2343 24564
rect -2325 24518 -2320 24564
rect -2309 24546 -2301 24554
rect -2068 24547 -2040 24554
rect -2317 24538 -2309 24546
rect -2000 24537 -1992 24564
rect -1850 24556 -1844 24564
rect -1840 24556 -1792 24564
rect -1894 24554 -1850 24555
rect -1958 24552 -1955 24553
rect -1969 24546 -1955 24552
rect -1894 24547 -1802 24554
rect -1894 24546 -1850 24547
rect -1655 24546 -1647 24554
rect -1969 24544 -1942 24546
rect -1955 24537 -1942 24544
rect -1844 24539 -1802 24545
rect -1663 24538 -1655 24546
rect -1860 24537 -1796 24538
rect -2040 24530 -2020 24537
rect -2004 24530 -1945 24537
rect -1929 24535 -1794 24537
rect -1929 24530 -1850 24535
rect -1844 24530 -1794 24535
rect -2309 24518 -2301 24526
rect -2136 24518 -2129 24528
rect -2068 24520 -2040 24527
rect -2020 24518 -2004 24520
rect -2000 24518 -1992 24530
rect -1844 24529 -1796 24530
rect -1850 24520 -1802 24527
rect -1978 24518 -1942 24519
rect -1655 24518 -1647 24526
rect -1642 24518 -1637 24564
rect -1619 24518 -1614 24564
rect -1530 24518 -1526 24564
rect -1506 24518 -1502 24564
rect -1482 24518 -1478 24564
rect -1458 24518 -1454 24564
rect -1434 24518 -1430 24564
rect -1410 24518 -1406 24564
rect -1386 24518 -1382 24564
rect -1362 24518 -1358 24564
rect -1338 24518 -1334 24564
rect -1314 24518 -1310 24564
rect -1290 24518 -1286 24564
rect -1266 24518 -1262 24564
rect -1242 24518 -1238 24564
rect -1218 24518 -1214 24564
rect -1194 24518 -1190 24564
rect -1170 24518 -1166 24564
rect -1146 24518 -1142 24564
rect -1122 24518 -1118 24564
rect -1098 24518 -1094 24564
rect -1074 24518 -1070 24564
rect -1050 24518 -1046 24564
rect -1026 24518 -1022 24564
rect -1002 24518 -998 24564
rect -978 24518 -974 24564
rect -954 24518 -950 24564
rect -930 24518 -926 24564
rect -906 24518 -902 24564
rect -882 24518 -878 24564
rect -858 24518 -854 24564
rect -834 24518 -830 24564
rect -810 24518 -806 24564
rect -786 24518 -782 24564
rect -762 24518 -758 24564
rect -738 24518 -734 24564
rect -714 24518 -710 24564
rect -690 24518 -686 24564
rect -666 24518 -662 24564
rect -642 24518 -638 24564
rect -618 24518 -614 24564
rect -594 24518 -590 24564
rect -570 24518 -566 24564
rect -546 24518 -542 24564
rect -522 24518 -518 24564
rect -498 24518 -494 24564
rect -474 24518 -470 24564
rect -450 24518 -446 24564
rect -426 24518 -422 24564
rect -402 24518 -398 24564
rect -378 24518 -374 24564
rect -354 24518 -350 24564
rect -330 24518 -326 24564
rect -306 24518 -302 24564
rect -282 24518 -278 24564
rect -258 24518 -254 24564
rect -234 24518 -230 24564
rect -210 24518 -206 24564
rect -186 24518 -182 24564
rect -162 24518 -158 24564
rect -138 24518 -134 24564
rect -114 24518 -110 24564
rect -90 24518 -86 24564
rect -66 24518 -62 24564
rect -42 24518 -38 24564
rect -18 24518 -14 24564
rect 6 24518 10 24564
rect 30 24518 34 24564
rect 54 24518 58 24564
rect 78 24518 82 24564
rect 102 24518 106 24564
rect 126 24518 130 24564
rect 150 24518 154 24564
rect 174 24518 178 24564
rect 198 24518 202 24564
rect 222 24518 226 24564
rect 246 24518 250 24564
rect 270 24518 274 24564
rect 294 24518 298 24564
rect 318 24518 322 24564
rect 342 24518 346 24564
rect 366 24518 370 24564
rect 390 24518 394 24564
rect 414 24518 418 24564
rect 438 24518 442 24564
rect 462 24518 466 24564
rect 486 24518 490 24564
rect 510 24518 514 24564
rect 534 24518 538 24564
rect 558 24518 562 24564
rect 582 24518 586 24564
rect 595 24557 600 24564
rect 605 24543 610 24557
rect 606 24518 610 24543
rect 630 24518 634 24588
rect 654 24518 658 24588
rect 678 24518 682 24588
rect 702 24518 706 24588
rect 726 24518 730 24588
rect 750 24518 754 24588
rect 774 24518 778 24588
rect 798 24518 802 24588
rect 822 24518 826 24588
rect 846 24518 850 24588
rect 870 24518 874 24588
rect 894 24518 898 24588
rect 918 24518 922 24588
rect 942 24518 946 24588
rect 966 24518 970 24588
rect 990 24518 994 24588
rect 1014 24518 1018 24588
rect 1038 24518 1042 24588
rect 1062 24518 1066 24588
rect 1086 24518 1090 24588
rect 1110 24518 1114 24588
rect 1134 24518 1138 24588
rect 1158 24518 1162 24588
rect 1182 24518 1186 24588
rect 1206 24518 1210 24588
rect 1230 24518 1234 24588
rect 1254 24518 1258 24588
rect 1278 24518 1282 24588
rect 1302 24518 1306 24588
rect 1326 24518 1330 24588
rect 1350 24518 1354 24588
rect 1374 24518 1378 24588
rect 1398 24518 1402 24588
rect 1422 24518 1426 24588
rect 1446 24518 1450 24588
rect 1470 24518 1474 24588
rect 1494 24518 1498 24588
rect 1518 24518 1522 24588
rect 1542 24518 1546 24588
rect 1566 24518 1570 24588
rect 1590 24518 1594 24588
rect 1614 24518 1618 24588
rect 1638 24518 1642 24588
rect 1662 24518 1666 24588
rect 1686 24518 1690 24588
rect 1710 24518 1714 24588
rect 1734 24518 1738 24588
rect 1758 24518 1762 24588
rect 1782 24518 1786 24588
rect 1806 24518 1810 24588
rect 1830 24518 1834 24588
rect 1837 24587 1851 24588
rect 1854 24587 1861 24612
rect 1854 24518 1858 24587
rect 1878 24518 1882 24612
rect 1902 24518 1906 24612
rect 1926 24518 1930 24612
rect 1950 24518 1954 24612
rect 1974 24518 1978 24612
rect 1998 24518 2002 24612
rect 2022 24518 2026 24612
rect 2046 24518 2050 24612
rect 2070 24518 2074 24612
rect 2094 24518 2098 24612
rect 2118 24518 2122 24612
rect 2142 24518 2146 24612
rect 2166 24518 2170 24612
rect 2190 24518 2194 24612
rect 2214 24518 2218 24612
rect 2238 24518 2242 24612
rect 2262 24518 2266 24612
rect 2286 24518 2290 24612
rect 2310 24518 2314 24612
rect 2334 24518 2338 24612
rect 2358 24518 2362 24612
rect 2382 24518 2386 24612
rect 2406 24518 2410 24612
rect 2430 24518 2434 24612
rect 2454 24518 2458 24612
rect 2478 24518 2482 24612
rect 2502 24518 2506 24612
rect 2526 24518 2530 24612
rect 2539 24605 2544 24612
rect 2550 24605 2554 24612
rect 2549 24591 2554 24605
rect 2539 24581 2544 24591
rect 2549 24567 2554 24581
rect 2550 24519 2554 24567
rect 2539 24518 2571 24519
rect -2393 24516 2571 24518
rect -2371 24398 -2366 24516
rect -2348 24398 -2343 24516
rect -2325 24478 -2320 24516
rect -2317 24510 -2309 24516
rect -2124 24512 -2117 24516
rect -2060 24512 -2040 24516
rect -2060 24503 -2030 24510
rect -2062 24478 -2032 24479
rect -2000 24478 -1992 24516
rect -1844 24512 -1802 24516
rect -1844 24502 -1792 24511
rect -1663 24510 -1655 24516
rect -1942 24480 -1937 24492
rect -1850 24489 -1822 24490
rect -1850 24485 -1802 24489
rect -2325 24470 -2317 24478
rect -2062 24476 -1961 24478
rect -2325 24450 -2320 24470
rect -2317 24462 -2309 24470
rect -2062 24463 -2040 24474
rect -2032 24469 -1961 24476
rect -1947 24470 -1942 24478
rect -1842 24476 -1794 24479
rect -2070 24458 -2022 24462
rect -2325 24434 -2317 24450
rect -2080 24436 -2032 24445
rect -2325 24418 -2320 24434
rect -2309 24422 -2301 24434
rect -2070 24427 -2040 24434
rect -2317 24418 -2309 24422
rect -2325 24406 -2317 24418
rect -2000 24417 -1992 24469
rect -1942 24468 -1937 24470
rect -1932 24460 -1927 24468
rect -1912 24465 -1896 24471
rect -1842 24463 -1802 24474
rect -1671 24470 -1663 24478
rect -1663 24462 -1655 24470
rect -1850 24458 -1680 24462
rect -1937 24444 -1934 24446
rect -1924 24444 -1921 24446
rect -1850 24436 -1842 24446
rect -1840 24436 -1792 24445
rect -1924 24434 -1850 24435
rect -1671 24434 -1663 24450
rect -1960 24432 -1955 24433
rect -1969 24426 -1955 24432
rect -1924 24427 -1802 24434
rect -1924 24426 -1850 24427
rect -1969 24424 -1944 24426
rect -1955 24417 -1944 24424
rect -1842 24419 -1802 24425
rect -1655 24422 -1647 24434
rect -1663 24418 -1655 24422
rect -1860 24417 -1794 24418
rect -2040 24410 -1945 24417
rect -1929 24415 -1794 24417
rect -1929 24410 -1850 24415
rect -2325 24398 -2320 24406
rect -2309 24398 -2301 24406
rect -2070 24400 -2040 24407
rect -2000 24398 -1992 24410
rect -1842 24409 -1794 24415
rect -1945 24400 -1942 24402
rect -1850 24400 -1802 24407
rect -1671 24406 -1663 24418
rect -1978 24398 -1942 24399
rect -1655 24398 -1647 24406
rect -1642 24398 -1637 24516
rect -1619 24398 -1614 24516
rect -1530 24398 -1526 24516
rect -1506 24398 -1502 24516
rect -1482 24398 -1478 24516
rect -1458 24398 -1454 24516
rect -1434 24398 -1430 24516
rect -1410 24398 -1406 24516
rect -1386 24398 -1382 24516
rect -1362 24398 -1358 24516
rect -1338 24398 -1334 24516
rect -1314 24398 -1310 24516
rect -1290 24398 -1286 24516
rect -1266 24398 -1262 24516
rect -1242 24398 -1238 24516
rect -1218 24398 -1214 24516
rect -1194 24398 -1190 24516
rect -1170 24398 -1166 24516
rect -1146 24398 -1142 24516
rect -1122 24398 -1118 24516
rect -1098 24398 -1094 24516
rect -1074 24398 -1070 24516
rect -1050 24398 -1046 24516
rect -1026 24398 -1022 24516
rect -1002 24398 -998 24516
rect -978 24398 -974 24516
rect -954 24398 -950 24516
rect -930 24398 -926 24516
rect -906 24398 -902 24516
rect -882 24398 -878 24516
rect -858 24398 -854 24516
rect -834 24398 -830 24516
rect -810 24398 -806 24516
rect -786 24398 -782 24516
rect -762 24398 -758 24516
rect -738 24398 -734 24516
rect -714 24398 -710 24516
rect -690 24398 -686 24516
rect -666 24398 -662 24516
rect -642 24398 -638 24516
rect -618 24398 -614 24516
rect -594 24398 -590 24516
rect -570 24398 -566 24516
rect -546 24398 -542 24516
rect -522 24398 -518 24516
rect -498 24398 -494 24516
rect -474 24398 -470 24516
rect -450 24398 -446 24516
rect -426 24398 -422 24516
rect -402 24398 -398 24516
rect -378 24398 -374 24516
rect -354 24398 -350 24516
rect -330 24398 -326 24516
rect -306 24398 -302 24516
rect -282 24398 -278 24516
rect -258 24398 -254 24516
rect -234 24398 -230 24516
rect -210 24398 -206 24516
rect -186 24398 -182 24516
rect -162 24398 -158 24516
rect -138 24398 -134 24516
rect -114 24398 -110 24516
rect -90 24398 -86 24516
rect -66 24398 -62 24516
rect -42 24398 -38 24516
rect -18 24398 -14 24516
rect 6 24398 10 24516
rect 30 24398 34 24516
rect 54 24398 58 24516
rect 78 24398 82 24516
rect 102 24398 106 24516
rect 126 24398 130 24516
rect 150 24398 154 24516
rect 174 24398 178 24516
rect 198 24398 202 24516
rect 222 24398 226 24516
rect 246 24398 250 24516
rect 270 24398 274 24516
rect 294 24398 298 24516
rect 318 24398 322 24516
rect 342 24398 346 24516
rect 366 24398 370 24516
rect 390 24398 394 24516
rect 414 24398 418 24516
rect 438 24398 442 24516
rect 462 24398 466 24516
rect 486 24398 490 24516
rect 510 24398 514 24516
rect 534 24398 538 24516
rect 558 24398 562 24516
rect 582 24398 586 24516
rect 606 24398 610 24516
rect 630 24515 634 24516
rect 630 24494 637 24515
rect 654 24494 658 24516
rect 678 24494 682 24516
rect 702 24494 706 24516
rect 726 24494 730 24516
rect 750 24494 754 24516
rect 774 24494 778 24516
rect 798 24494 802 24516
rect 822 24494 826 24516
rect 846 24494 850 24516
rect 870 24494 874 24516
rect 894 24494 898 24516
rect 918 24494 922 24516
rect 942 24494 946 24516
rect 966 24494 970 24516
rect 990 24494 994 24516
rect 1014 24494 1018 24516
rect 1038 24494 1042 24516
rect 1062 24494 1066 24516
rect 1086 24494 1090 24516
rect 1110 24494 1114 24516
rect 1134 24494 1138 24516
rect 1158 24494 1162 24516
rect 1182 24494 1186 24516
rect 1206 24494 1210 24516
rect 1230 24494 1234 24516
rect 1254 24494 1258 24516
rect 1278 24494 1282 24516
rect 1302 24494 1306 24516
rect 1326 24494 1330 24516
rect 1350 24494 1354 24516
rect 1374 24494 1378 24516
rect 1398 24494 1402 24516
rect 1422 24494 1426 24516
rect 1446 24494 1450 24516
rect 1470 24494 1474 24516
rect 1494 24494 1498 24516
rect 1518 24494 1522 24516
rect 1542 24494 1546 24516
rect 1566 24494 1570 24516
rect 1590 24494 1594 24516
rect 1614 24494 1618 24516
rect 1638 24494 1642 24516
rect 1662 24494 1666 24516
rect 1686 24494 1690 24516
rect 1710 24494 1714 24516
rect 1734 24494 1738 24516
rect 1758 24494 1762 24516
rect 1782 24494 1786 24516
rect 1806 24494 1810 24516
rect 1830 24494 1834 24516
rect 1854 24494 1858 24516
rect 1878 24494 1882 24516
rect 1902 24494 1906 24516
rect 1926 24494 1930 24516
rect 1950 24494 1954 24516
rect 1974 24494 1978 24516
rect 1998 24494 2002 24516
rect 2022 24494 2026 24516
rect 2046 24494 2050 24516
rect 2070 24494 2074 24516
rect 2094 24494 2098 24516
rect 2118 24494 2122 24516
rect 2142 24494 2146 24516
rect 2166 24494 2170 24516
rect 2190 24494 2194 24516
rect 2214 24494 2218 24516
rect 2238 24494 2242 24516
rect 2262 24494 2266 24516
rect 2286 24494 2290 24516
rect 2310 24494 2314 24516
rect 2334 24494 2338 24516
rect 2358 24494 2362 24516
rect 2382 24494 2386 24516
rect 2406 24494 2410 24516
rect 2430 24494 2434 24516
rect 2454 24494 2458 24516
rect 2478 24494 2482 24516
rect 2502 24494 2506 24516
rect 2526 24495 2530 24516
rect 2539 24509 2544 24516
rect 2550 24509 2554 24516
rect 2557 24515 2571 24516
rect 2549 24495 2554 24509
rect 2563 24505 2571 24509
rect 2557 24495 2563 24505
rect 2515 24494 2549 24495
rect 613 24492 2549 24494
rect 613 24491 627 24492
rect 630 24467 637 24492
rect 630 24398 634 24467
rect 654 24398 658 24492
rect 678 24398 682 24492
rect 702 24398 706 24492
rect 726 24398 730 24492
rect 750 24398 754 24492
rect 774 24398 778 24492
rect 798 24398 802 24492
rect 822 24398 826 24492
rect 846 24398 850 24492
rect 870 24398 874 24492
rect 894 24398 898 24492
rect 918 24398 922 24492
rect 942 24398 946 24492
rect 966 24398 970 24492
rect 990 24398 994 24492
rect 1014 24398 1018 24492
rect 1038 24398 1042 24492
rect 1062 24398 1066 24492
rect 1086 24398 1090 24492
rect 1110 24398 1114 24492
rect 1134 24398 1138 24492
rect 1158 24398 1162 24492
rect 1182 24398 1186 24492
rect 1206 24398 1210 24492
rect 1230 24398 1234 24492
rect 1254 24398 1258 24492
rect 1278 24398 1282 24492
rect 1302 24398 1306 24492
rect 1326 24398 1330 24492
rect 1350 24398 1354 24492
rect 1374 24398 1378 24492
rect 1398 24398 1402 24492
rect 1422 24398 1426 24492
rect 1446 24398 1450 24492
rect 1470 24398 1474 24492
rect 1494 24398 1498 24492
rect 1518 24398 1522 24492
rect 1542 24398 1546 24492
rect 1566 24398 1570 24492
rect 1590 24398 1594 24492
rect 1614 24398 1618 24492
rect 1638 24398 1642 24492
rect 1662 24398 1666 24492
rect 1686 24398 1690 24492
rect 1710 24398 1714 24492
rect 1734 24398 1738 24492
rect 1758 24398 1762 24492
rect 1782 24398 1786 24492
rect 1806 24398 1810 24492
rect 1830 24398 1834 24492
rect 1854 24398 1858 24492
rect 1878 24398 1882 24492
rect 1902 24398 1906 24492
rect 1926 24398 1930 24492
rect 1950 24398 1954 24492
rect 1974 24398 1978 24492
rect 1998 24398 2002 24492
rect 2022 24398 2026 24492
rect 2046 24398 2050 24492
rect 2070 24398 2074 24492
rect 2094 24398 2098 24492
rect 2107 24461 2112 24471
rect 2118 24461 2122 24492
rect 2117 24447 2122 24461
rect 2107 24437 2112 24447
rect 2117 24423 2122 24437
rect 2118 24398 2122 24423
rect 2142 24398 2146 24492
rect 2166 24398 2170 24492
rect 2190 24398 2194 24492
rect 2214 24398 2218 24492
rect 2238 24398 2242 24492
rect 2262 24398 2266 24492
rect 2286 24398 2290 24492
rect 2310 24398 2314 24492
rect 2334 24398 2338 24492
rect 2358 24398 2362 24492
rect 2382 24398 2386 24492
rect 2406 24398 2410 24492
rect 2430 24398 2434 24492
rect 2454 24398 2458 24492
rect 2478 24398 2482 24492
rect 2502 24398 2506 24492
rect 2515 24485 2520 24492
rect 2526 24485 2530 24492
rect 2525 24471 2530 24485
rect 2515 24461 2520 24471
rect 2525 24447 2530 24461
rect 2526 24399 2530 24447
rect 2515 24398 2547 24399
rect -2393 24396 2547 24398
rect -2371 24302 -2366 24396
rect -2348 24302 -2343 24396
rect -2325 24390 -2320 24396
rect -2309 24394 -2301 24396
rect -2317 24390 -2309 24394
rect -2062 24392 -2040 24396
rect -2325 24378 -2317 24390
rect -2062 24383 -2032 24390
rect -2325 24358 -2320 24378
rect -2062 24358 -2032 24359
rect -2000 24358 -1992 24396
rect -1888 24391 -1874 24396
rect -1842 24392 -1802 24396
rect -1655 24394 -1647 24396
rect -1932 24382 -1924 24391
rect -1904 24389 -1874 24391
rect -1842 24382 -1792 24391
rect -1663 24390 -1655 24394
rect -1671 24378 -1663 24390
rect -1942 24360 -1937 24372
rect -1850 24369 -1822 24370
rect -1850 24365 -1802 24369
rect -2325 24350 -2317 24358
rect -2062 24356 -1961 24358
rect -2325 24330 -2320 24350
rect -2317 24342 -2309 24350
rect -2062 24343 -2040 24354
rect -2032 24349 -1961 24356
rect -1947 24350 -1942 24358
rect -1842 24356 -1794 24359
rect -2070 24338 -2022 24342
rect -2325 24316 -2317 24330
rect -2072 24322 -2032 24323
rect -2102 24316 -2032 24322
rect -2325 24302 -2320 24316
rect -2317 24314 -2309 24316
rect -2309 24302 -2301 24314
rect -2070 24307 -2062 24312
rect -2000 24302 -1992 24349
rect -1942 24348 -1937 24350
rect -1932 24340 -1927 24348
rect -1912 24345 -1896 24351
rect -1842 24343 -1802 24354
rect -1671 24350 -1663 24358
rect -1663 24342 -1655 24350
rect -1850 24338 -1680 24342
rect -1924 24324 -1921 24326
rect -1806 24316 -1680 24322
rect -1671 24316 -1663 24330
rect -1663 24314 -1655 24316
rect -1854 24307 -1806 24312
rect -1974 24302 -1964 24303
rect -1960 24302 -1944 24304
rect -1842 24302 -1806 24305
rect -1655 24302 -1647 24314
rect -1642 24302 -1637 24396
rect -1619 24302 -1614 24396
rect -1530 24302 -1526 24396
rect -1506 24302 -1502 24396
rect -1482 24302 -1478 24396
rect -1458 24302 -1454 24396
rect -1434 24302 -1430 24396
rect -1410 24302 -1406 24396
rect -1386 24302 -1382 24396
rect -1362 24302 -1358 24396
rect -1338 24302 -1334 24396
rect -1314 24302 -1310 24396
rect -1290 24302 -1286 24396
rect -1266 24302 -1262 24396
rect -1242 24302 -1238 24396
rect -1218 24302 -1214 24396
rect -1194 24302 -1190 24396
rect -1170 24302 -1166 24396
rect -1146 24302 -1142 24396
rect -1122 24302 -1118 24396
rect -1098 24302 -1094 24396
rect -1074 24302 -1070 24396
rect -1050 24302 -1046 24396
rect -1026 24302 -1022 24396
rect -1002 24302 -998 24396
rect -978 24302 -974 24396
rect -954 24302 -950 24396
rect -930 24302 -926 24396
rect -906 24302 -902 24396
rect -882 24302 -878 24396
rect -858 24302 -854 24396
rect -834 24302 -830 24396
rect -810 24302 -806 24396
rect -786 24302 -782 24396
rect -762 24302 -758 24396
rect -738 24302 -734 24396
rect -714 24302 -710 24396
rect -690 24302 -686 24396
rect -666 24302 -662 24396
rect -642 24302 -638 24396
rect -618 24302 -614 24396
rect -594 24302 -590 24396
rect -570 24302 -566 24396
rect -546 24302 -542 24396
rect -522 24302 -518 24396
rect -498 24302 -494 24396
rect -474 24302 -470 24396
rect -450 24302 -446 24396
rect -426 24302 -422 24396
rect -402 24302 -398 24396
rect -378 24302 -374 24396
rect -354 24302 -350 24396
rect -330 24302 -326 24396
rect -306 24302 -302 24396
rect -282 24302 -278 24396
rect -258 24302 -254 24396
rect -234 24302 -230 24396
rect -210 24302 -206 24396
rect -186 24302 -182 24396
rect -162 24302 -158 24396
rect -138 24302 -134 24396
rect -114 24302 -110 24396
rect -90 24302 -86 24396
rect -66 24302 -62 24396
rect -42 24302 -38 24396
rect -18 24302 -14 24396
rect 6 24302 10 24396
rect 30 24302 34 24396
rect 54 24302 58 24396
rect 78 24302 82 24396
rect 102 24302 106 24396
rect 126 24302 130 24396
rect 150 24302 154 24396
rect 174 24302 178 24396
rect 198 24302 202 24396
rect 222 24302 226 24396
rect 246 24302 250 24396
rect 270 24302 274 24396
rect 294 24302 298 24396
rect 318 24302 322 24396
rect 342 24302 346 24396
rect 366 24302 370 24396
rect 390 24302 394 24396
rect 414 24302 418 24396
rect 438 24302 442 24396
rect 462 24302 466 24396
rect 486 24302 490 24396
rect 510 24302 514 24396
rect 534 24302 538 24396
rect 558 24302 562 24396
rect 582 24302 586 24396
rect 606 24302 610 24396
rect 630 24302 634 24396
rect 654 24302 658 24396
rect 678 24302 682 24396
rect 702 24351 706 24396
rect 691 24350 725 24351
rect 726 24350 730 24396
rect 750 24350 754 24396
rect 774 24350 778 24396
rect 798 24350 802 24396
rect 822 24350 826 24396
rect 846 24350 850 24396
rect 870 24350 874 24396
rect 894 24350 898 24396
rect 918 24350 922 24396
rect 942 24350 946 24396
rect 966 24350 970 24396
rect 990 24350 994 24396
rect 1014 24350 1018 24396
rect 1038 24350 1042 24396
rect 1062 24350 1066 24396
rect 1086 24350 1090 24396
rect 1110 24350 1114 24396
rect 1134 24350 1138 24396
rect 1158 24350 1162 24396
rect 1182 24350 1186 24396
rect 1206 24350 1210 24396
rect 1230 24350 1234 24396
rect 1254 24350 1258 24396
rect 1278 24350 1282 24396
rect 1302 24350 1306 24396
rect 1326 24350 1330 24396
rect 1350 24350 1354 24396
rect 1374 24350 1378 24396
rect 1398 24350 1402 24396
rect 1422 24350 1426 24396
rect 1446 24350 1450 24396
rect 1470 24350 1474 24396
rect 1494 24350 1498 24396
rect 1518 24350 1522 24396
rect 1542 24350 1546 24396
rect 1566 24350 1570 24396
rect 1590 24350 1594 24396
rect 1614 24350 1618 24396
rect 1638 24350 1642 24396
rect 1662 24350 1666 24396
rect 1686 24350 1690 24396
rect 1710 24350 1714 24396
rect 1734 24350 1738 24396
rect 1758 24350 1762 24396
rect 1782 24350 1786 24396
rect 1806 24350 1810 24396
rect 1830 24350 1834 24396
rect 1854 24350 1858 24396
rect 1878 24350 1882 24396
rect 1902 24350 1906 24396
rect 1926 24350 1930 24396
rect 1950 24350 1954 24396
rect 1974 24350 1978 24396
rect 1998 24350 2002 24396
rect 2022 24350 2026 24396
rect 2046 24350 2050 24396
rect 2070 24350 2074 24396
rect 2094 24350 2098 24396
rect 2118 24350 2122 24396
rect 2142 24395 2146 24396
rect 2142 24374 2149 24395
rect 2166 24374 2170 24396
rect 2190 24374 2194 24396
rect 2214 24374 2218 24396
rect 2238 24374 2242 24396
rect 2262 24374 2266 24396
rect 2286 24374 2290 24396
rect 2310 24374 2314 24396
rect 2334 24374 2338 24396
rect 2358 24374 2362 24396
rect 2382 24374 2386 24396
rect 2406 24374 2410 24396
rect 2430 24374 2434 24396
rect 2454 24374 2458 24396
rect 2478 24374 2482 24396
rect 2502 24375 2506 24396
rect 2515 24389 2520 24396
rect 2526 24389 2530 24396
rect 2533 24395 2547 24396
rect 2525 24375 2530 24389
rect 2539 24385 2547 24389
rect 2533 24375 2539 24385
rect 2491 24374 2525 24375
rect 2125 24372 2525 24374
rect 2125 24371 2139 24372
rect 691 24348 2139 24350
rect 691 24341 696 24348
rect 702 24341 706 24348
rect 701 24327 706 24341
rect 691 24317 696 24327
rect 701 24303 706 24317
rect 702 24302 706 24303
rect 726 24302 730 24348
rect 750 24302 754 24348
rect 774 24302 778 24348
rect 798 24302 802 24348
rect 822 24302 826 24348
rect 846 24302 850 24348
rect 870 24302 874 24348
rect 894 24302 898 24348
rect 918 24302 922 24348
rect 942 24302 946 24348
rect 966 24302 970 24348
rect 990 24302 994 24348
rect 1014 24302 1018 24348
rect 1038 24302 1042 24348
rect 1062 24302 1066 24348
rect 1086 24302 1090 24348
rect 1110 24302 1114 24348
rect 1134 24302 1138 24348
rect 1158 24302 1162 24348
rect 1182 24302 1186 24348
rect 1206 24302 1210 24348
rect 1230 24302 1234 24348
rect 1254 24302 1258 24348
rect 1278 24302 1282 24348
rect 1302 24302 1306 24348
rect 1326 24302 1330 24348
rect 1350 24302 1354 24348
rect 1374 24302 1378 24348
rect 1398 24302 1402 24348
rect 1422 24302 1426 24348
rect 1446 24302 1450 24348
rect 1470 24302 1474 24348
rect 1494 24302 1498 24348
rect 1518 24302 1522 24348
rect 1542 24302 1546 24348
rect 1566 24303 1570 24348
rect 1555 24302 1589 24303
rect -2393 24300 1589 24302
rect -2371 24278 -2366 24300
rect -2348 24278 -2343 24300
rect -2325 24288 -2317 24300
rect -2325 24278 -2320 24288
rect -2317 24286 -2309 24288
rect -2062 24287 -2032 24294
rect -2309 24278 -2301 24286
rect -2070 24280 -2062 24287
rect -2000 24282 -1992 24300
rect -1974 24298 -1944 24300
rect -1960 24297 -1944 24298
rect -1842 24296 -1806 24300
rect -1842 24289 -1798 24294
rect -1806 24287 -1798 24289
rect -1671 24288 -1663 24300
rect -1854 24285 -1842 24287
rect -1663 24286 -1655 24288
rect -2062 24278 -2036 24280
rect -2393 24276 -2036 24278
rect -2032 24278 -2012 24280
rect -2004 24278 -1974 24282
rect -1854 24280 -1806 24285
rect -1864 24278 -1796 24279
rect -1655 24278 -1647 24286
rect -1642 24278 -1637 24300
rect -1619 24278 -1614 24300
rect -1530 24278 -1526 24300
rect -1506 24278 -1502 24300
rect -1482 24278 -1478 24300
rect -1458 24278 -1454 24300
rect -1434 24278 -1430 24300
rect -1410 24278 -1406 24300
rect -1386 24278 -1382 24300
rect -1362 24278 -1358 24300
rect -1338 24278 -1334 24300
rect -1314 24278 -1310 24300
rect -1290 24278 -1286 24300
rect -1266 24278 -1262 24300
rect -1242 24278 -1238 24300
rect -1218 24278 -1214 24300
rect -1194 24278 -1190 24300
rect -1170 24278 -1166 24300
rect -1146 24278 -1142 24300
rect -1122 24278 -1118 24300
rect -1098 24278 -1094 24300
rect -1074 24278 -1070 24300
rect -1050 24278 -1046 24300
rect -1026 24278 -1022 24300
rect -1002 24278 -998 24300
rect -978 24278 -974 24300
rect -954 24278 -950 24300
rect -930 24278 -926 24300
rect -906 24278 -902 24300
rect -882 24278 -878 24300
rect -858 24278 -854 24300
rect -834 24278 -830 24300
rect -810 24278 -806 24300
rect -786 24278 -782 24300
rect -762 24278 -758 24300
rect -738 24278 -734 24300
rect -714 24278 -710 24300
rect -690 24278 -686 24300
rect -666 24278 -662 24300
rect -642 24278 -638 24300
rect -618 24278 -614 24300
rect -594 24278 -590 24300
rect -570 24278 -566 24300
rect -546 24278 -542 24300
rect -522 24278 -518 24300
rect -498 24278 -494 24300
rect -474 24278 -470 24300
rect -450 24278 -446 24300
rect -426 24278 -422 24300
rect -402 24278 -398 24300
rect -378 24278 -374 24300
rect -354 24278 -350 24300
rect -330 24278 -326 24300
rect -306 24278 -302 24300
rect -282 24278 -278 24300
rect -258 24278 -254 24300
rect -234 24278 -230 24300
rect -210 24278 -206 24300
rect -186 24278 -182 24300
rect -162 24278 -158 24300
rect -138 24278 -134 24300
rect -114 24278 -110 24300
rect -90 24278 -86 24300
rect -66 24278 -62 24300
rect -42 24278 -38 24300
rect -18 24278 -14 24300
rect 6 24278 10 24300
rect 30 24278 34 24300
rect 54 24278 58 24300
rect 78 24278 82 24300
rect 102 24278 106 24300
rect 126 24278 130 24300
rect 150 24278 154 24300
rect 174 24278 178 24300
rect 198 24278 202 24300
rect 222 24278 226 24300
rect 246 24278 250 24300
rect 270 24278 274 24300
rect 294 24278 298 24300
rect 318 24278 322 24300
rect 342 24278 346 24300
rect 366 24278 370 24300
rect 390 24278 394 24300
rect 414 24278 418 24300
rect 438 24278 442 24300
rect 462 24278 466 24300
rect 486 24278 490 24300
rect 510 24278 514 24300
rect 534 24278 538 24300
rect 558 24278 562 24300
rect 582 24278 586 24300
rect 606 24278 610 24300
rect 630 24278 634 24300
rect 654 24278 658 24300
rect 678 24278 682 24300
rect 702 24278 706 24300
rect 726 24278 730 24300
rect 750 24278 754 24300
rect 774 24278 778 24300
rect 798 24278 802 24300
rect 822 24278 826 24300
rect 846 24278 850 24300
rect 870 24278 874 24300
rect 894 24278 898 24300
rect 918 24278 922 24300
rect 942 24278 946 24300
rect 966 24278 970 24300
rect 990 24278 994 24300
rect 1014 24278 1018 24300
rect 1038 24278 1042 24300
rect 1062 24278 1066 24300
rect 1086 24278 1090 24300
rect 1110 24278 1114 24300
rect 1134 24278 1138 24300
rect 1158 24278 1162 24300
rect 1182 24278 1186 24300
rect 1206 24278 1210 24300
rect 1230 24278 1234 24300
rect 1254 24278 1258 24300
rect 1278 24278 1282 24300
rect 1302 24278 1306 24300
rect 1326 24278 1330 24300
rect 1350 24278 1354 24300
rect 1374 24278 1378 24300
rect 1398 24278 1402 24300
rect 1422 24278 1426 24300
rect 1446 24278 1450 24300
rect 1470 24278 1474 24300
rect 1494 24278 1498 24300
rect 1518 24278 1522 24300
rect 1542 24278 1546 24300
rect 1555 24293 1560 24300
rect 1566 24293 1570 24300
rect 1565 24279 1570 24293
rect 1566 24278 1570 24279
rect 1590 24278 1594 24348
rect 1614 24278 1618 24348
rect 1638 24278 1642 24348
rect 1662 24278 1666 24348
rect 1686 24278 1690 24348
rect 1710 24278 1714 24348
rect 1734 24278 1738 24348
rect 1758 24278 1762 24348
rect 1782 24278 1786 24348
rect 1806 24278 1810 24348
rect 1830 24278 1834 24348
rect 1854 24278 1858 24348
rect 1878 24278 1882 24348
rect 1902 24278 1906 24348
rect 1926 24278 1930 24348
rect 1950 24278 1954 24348
rect 1974 24278 1978 24348
rect 1998 24278 2002 24348
rect 2022 24278 2026 24348
rect 2046 24278 2050 24348
rect 2070 24278 2074 24348
rect 2094 24278 2098 24348
rect 2118 24278 2122 24348
rect 2125 24347 2139 24348
rect 2142 24347 2149 24372
rect 2142 24278 2146 24347
rect 2166 24278 2170 24372
rect 2190 24278 2194 24372
rect 2214 24278 2218 24372
rect 2238 24278 2242 24372
rect 2262 24278 2266 24372
rect 2286 24278 2290 24372
rect 2310 24278 2314 24372
rect 2334 24278 2338 24372
rect 2358 24278 2362 24372
rect 2382 24278 2386 24372
rect 2406 24278 2410 24372
rect 2430 24278 2434 24372
rect 2454 24278 2458 24372
rect 2478 24278 2482 24372
rect 2491 24365 2496 24372
rect 2502 24365 2506 24372
rect 2501 24351 2506 24365
rect 2491 24341 2496 24351
rect 2501 24327 2506 24341
rect 2502 24279 2506 24327
rect 2491 24278 2523 24279
rect -2032 24276 2523 24278
rect -2371 24230 -2366 24276
rect -2348 24230 -2343 24276
rect -2325 24272 -2320 24276
rect -2309 24274 -2301 24276
rect -2317 24272 -2309 24274
rect -2325 24260 -2317 24272
rect -2052 24270 -2036 24272
rect -2052 24268 -2032 24270
rect -2062 24262 -2032 24268
rect -2325 24230 -2320 24260
rect -2317 24258 -2309 24260
rect -2092 24246 -2062 24248
rect -2094 24242 -2062 24246
rect -2000 24230 -1992 24276
rect -1904 24269 -1874 24276
rect -1842 24269 -1806 24276
rect -1655 24274 -1647 24276
rect -1663 24272 -1655 24274
rect -1842 24262 -1680 24268
rect -1671 24260 -1663 24272
rect -1663 24258 -1655 24260
rect -1854 24246 -1806 24248
rect -1854 24242 -1680 24246
rect -1642 24230 -1637 24276
rect -1619 24230 -1614 24276
rect -1530 24230 -1526 24276
rect -1506 24230 -1502 24276
rect -1482 24230 -1478 24276
rect -1458 24230 -1454 24276
rect -1434 24230 -1430 24276
rect -1410 24230 -1406 24276
rect -1386 24230 -1382 24276
rect -1362 24230 -1358 24276
rect -1338 24230 -1334 24276
rect -1314 24230 -1310 24276
rect -1290 24230 -1286 24276
rect -1266 24230 -1262 24276
rect -1242 24230 -1238 24276
rect -1218 24230 -1214 24276
rect -1194 24230 -1190 24276
rect -1170 24230 -1166 24276
rect -1146 24230 -1142 24276
rect -1122 24230 -1118 24276
rect -1098 24230 -1094 24276
rect -1074 24230 -1070 24276
rect -1050 24230 -1046 24276
rect -1026 24230 -1022 24276
rect -1002 24230 -998 24276
rect -978 24230 -974 24276
rect -954 24230 -950 24276
rect -930 24230 -926 24276
rect -906 24230 -902 24276
rect -882 24230 -878 24276
rect -858 24230 -854 24276
rect -834 24230 -830 24276
rect -810 24230 -806 24276
rect -786 24230 -782 24276
rect -762 24230 -758 24276
rect -738 24230 -734 24276
rect -714 24230 -710 24276
rect -690 24230 -686 24276
rect -666 24230 -662 24276
rect -642 24230 -638 24276
rect -618 24230 -614 24276
rect -594 24230 -590 24276
rect -570 24230 -566 24276
rect -546 24230 -542 24276
rect -522 24230 -518 24276
rect -498 24230 -494 24276
rect -474 24230 -470 24276
rect -450 24230 -446 24276
rect -426 24230 -422 24276
rect -402 24230 -398 24276
rect -378 24230 -374 24276
rect -354 24230 -350 24276
rect -330 24230 -326 24276
rect -306 24230 -302 24276
rect -282 24230 -278 24276
rect -258 24230 -254 24276
rect -234 24230 -230 24276
rect -210 24230 -206 24276
rect -186 24230 -182 24276
rect -162 24230 -158 24276
rect -138 24230 -134 24276
rect -114 24230 -110 24276
rect -90 24230 -86 24276
rect -66 24230 -62 24276
rect -42 24230 -38 24276
rect -18 24230 -14 24276
rect 6 24230 10 24276
rect 30 24230 34 24276
rect 54 24230 58 24276
rect 78 24230 82 24276
rect 102 24230 106 24276
rect 126 24230 130 24276
rect 150 24230 154 24276
rect 174 24230 178 24276
rect 198 24230 202 24276
rect 222 24230 226 24276
rect 246 24230 250 24276
rect 270 24230 274 24276
rect 294 24230 298 24276
rect 318 24230 322 24276
rect 342 24230 346 24276
rect 366 24230 370 24276
rect 390 24230 394 24276
rect 414 24230 418 24276
rect 438 24230 442 24276
rect 462 24230 466 24276
rect 486 24230 490 24276
rect 510 24230 514 24276
rect 534 24230 538 24276
rect 558 24230 562 24276
rect 582 24230 586 24276
rect 606 24230 610 24276
rect 630 24230 634 24276
rect 654 24230 658 24276
rect 678 24230 682 24276
rect 702 24230 706 24276
rect 726 24275 730 24276
rect -2393 24228 723 24230
rect -2371 24206 -2366 24228
rect -2348 24206 -2343 24228
rect -2325 24206 -2320 24228
rect -2072 24226 -2036 24227
rect -2072 24220 -2054 24226
rect -2309 24212 -2301 24220
rect -2317 24206 -2309 24212
rect -2092 24211 -2062 24216
rect -2000 24207 -1992 24228
rect -1938 24227 -1906 24228
rect -1920 24226 -1906 24227
rect -1806 24220 -1680 24226
rect -1854 24211 -1806 24216
rect -1655 24212 -1647 24220
rect -1982 24207 -1966 24208
rect -2000 24206 -1966 24207
rect -1846 24206 -1806 24209
rect -1663 24206 -1655 24212
rect -1642 24206 -1637 24228
rect -1619 24206 -1614 24228
rect -1530 24206 -1526 24228
rect -1506 24206 -1502 24228
rect -1482 24206 -1478 24228
rect -1458 24206 -1454 24228
rect -1434 24206 -1430 24228
rect -1410 24206 -1406 24228
rect -1386 24206 -1382 24228
rect -1362 24206 -1358 24228
rect -1338 24206 -1334 24228
rect -1314 24206 -1310 24228
rect -1290 24206 -1286 24228
rect -1266 24206 -1262 24228
rect -1242 24206 -1238 24228
rect -1218 24206 -1214 24228
rect -1194 24206 -1190 24228
rect -1170 24206 -1166 24228
rect -1146 24206 -1142 24228
rect -1122 24206 -1118 24228
rect -1098 24206 -1094 24228
rect -1074 24206 -1070 24228
rect -1050 24206 -1046 24228
rect -1026 24206 -1022 24228
rect -1002 24206 -998 24228
rect -978 24206 -974 24228
rect -954 24206 -950 24228
rect -930 24206 -926 24228
rect -906 24206 -902 24228
rect -882 24206 -878 24228
rect -858 24206 -854 24228
rect -834 24206 -830 24228
rect -810 24206 -806 24228
rect -786 24206 -782 24228
rect -762 24206 -758 24228
rect -738 24206 -734 24228
rect -714 24206 -710 24228
rect -690 24206 -686 24228
rect -666 24206 -662 24228
rect -642 24206 -638 24228
rect -618 24206 -614 24228
rect -594 24206 -590 24228
rect -570 24206 -566 24228
rect -546 24206 -542 24228
rect -522 24206 -518 24228
rect -498 24206 -494 24228
rect -474 24206 -470 24228
rect -450 24206 -446 24228
rect -426 24206 -422 24228
rect -402 24206 -398 24228
rect -378 24206 -374 24228
rect -354 24206 -350 24228
rect -330 24206 -326 24228
rect -306 24206 -302 24228
rect -282 24206 -278 24228
rect -258 24206 -254 24228
rect -234 24206 -230 24228
rect -210 24206 -206 24228
rect -186 24206 -182 24228
rect -162 24206 -158 24228
rect -138 24206 -134 24228
rect -114 24206 -110 24228
rect -90 24206 -86 24228
rect -66 24206 -62 24228
rect -42 24206 -38 24228
rect -18 24206 -14 24228
rect 6 24206 10 24228
rect 30 24206 34 24228
rect 54 24206 58 24228
rect 78 24206 82 24228
rect 102 24206 106 24228
rect 126 24206 130 24228
rect 150 24206 154 24228
rect 174 24206 178 24228
rect 198 24206 202 24228
rect 222 24206 226 24228
rect 246 24206 250 24228
rect 270 24206 274 24228
rect 294 24206 298 24228
rect 318 24206 322 24228
rect 342 24206 346 24228
rect 366 24206 370 24228
rect 390 24206 394 24228
rect 414 24206 418 24228
rect 438 24206 442 24228
rect 462 24206 466 24228
rect 486 24206 490 24228
rect 510 24206 514 24228
rect 534 24206 538 24228
rect 558 24206 562 24228
rect 582 24206 586 24228
rect 606 24206 610 24228
rect 630 24206 634 24228
rect 654 24206 658 24228
rect 678 24206 682 24228
rect 702 24206 706 24228
rect 709 24227 723 24228
rect 726 24227 733 24275
rect 726 24206 730 24227
rect 750 24206 754 24276
rect 774 24206 778 24276
rect 798 24206 802 24276
rect 822 24206 826 24276
rect 846 24206 850 24276
rect 870 24206 874 24276
rect 894 24206 898 24276
rect 918 24206 922 24276
rect 942 24206 946 24276
rect 966 24206 970 24276
rect 990 24206 994 24276
rect 1014 24206 1018 24276
rect 1038 24206 1042 24276
rect 1062 24206 1066 24276
rect 1086 24206 1090 24276
rect 1110 24206 1114 24276
rect 1134 24206 1138 24276
rect 1158 24206 1162 24276
rect 1182 24206 1186 24276
rect 1206 24206 1210 24276
rect 1230 24206 1234 24276
rect 1254 24206 1258 24276
rect 1278 24206 1282 24276
rect 1302 24206 1306 24276
rect 1326 24206 1330 24276
rect 1350 24206 1354 24276
rect 1374 24206 1378 24276
rect 1398 24206 1402 24276
rect 1422 24206 1426 24276
rect 1446 24206 1450 24276
rect 1470 24206 1474 24276
rect 1494 24206 1498 24276
rect 1518 24206 1522 24276
rect 1542 24206 1546 24276
rect 1566 24206 1570 24276
rect 1590 24227 1594 24276
rect -2393 24204 1587 24206
rect -2371 24182 -2366 24204
rect -2348 24182 -2343 24204
rect -2325 24182 -2320 24204
rect -2000 24202 -1966 24204
rect -2309 24184 -2301 24192
rect -2062 24191 -2054 24198
rect -2092 24184 -2084 24191
rect -2062 24184 -2026 24186
rect -2317 24182 -2309 24184
rect -2062 24182 -2012 24184
rect -2000 24182 -1992 24202
rect -1982 24201 -1966 24202
rect -1846 24200 -1806 24204
rect -1846 24193 -1798 24198
rect -1806 24191 -1798 24193
rect -1854 24189 -1846 24191
rect -1854 24184 -1806 24189
rect -1655 24184 -1647 24192
rect -1864 24182 -1796 24183
rect -1663 24182 -1655 24184
rect -1642 24182 -1637 24204
rect -1619 24182 -1614 24204
rect -1530 24182 -1526 24204
rect -1506 24182 -1502 24204
rect -1482 24182 -1478 24204
rect -1458 24182 -1454 24204
rect -1434 24182 -1430 24204
rect -1410 24182 -1406 24204
rect -1386 24182 -1382 24204
rect -1362 24182 -1358 24204
rect -1338 24182 -1334 24204
rect -1314 24182 -1310 24204
rect -1290 24182 -1286 24204
rect -1266 24182 -1262 24204
rect -1242 24182 -1238 24204
rect -1218 24182 -1214 24204
rect -1194 24182 -1190 24204
rect -1170 24182 -1166 24204
rect -1146 24182 -1142 24204
rect -1122 24182 -1118 24204
rect -1098 24182 -1094 24204
rect -1074 24182 -1070 24204
rect -1050 24182 -1046 24204
rect -1026 24182 -1022 24204
rect -1002 24182 -998 24204
rect -978 24182 -974 24204
rect -954 24182 -950 24204
rect -930 24182 -926 24204
rect -906 24182 -902 24204
rect -882 24182 -878 24204
rect -858 24182 -854 24204
rect -834 24182 -830 24204
rect -810 24182 -806 24204
rect -786 24182 -782 24204
rect -762 24182 -758 24204
rect -738 24182 -734 24204
rect -714 24182 -710 24204
rect -690 24182 -686 24204
rect -666 24182 -662 24204
rect -642 24182 -638 24204
rect -618 24182 -614 24204
rect -594 24182 -590 24204
rect -570 24182 -566 24204
rect -546 24182 -542 24204
rect -522 24182 -518 24204
rect -498 24182 -494 24204
rect -474 24182 -470 24204
rect -450 24182 -446 24204
rect -426 24182 -422 24204
rect -402 24182 -398 24204
rect -378 24182 -374 24204
rect -354 24182 -350 24204
rect -330 24182 -326 24204
rect -306 24182 -302 24204
rect -282 24182 -278 24204
rect -258 24182 -254 24204
rect -234 24182 -230 24204
rect -210 24182 -206 24204
rect -186 24182 -182 24204
rect -162 24182 -158 24204
rect -138 24182 -134 24204
rect -114 24182 -110 24204
rect -90 24182 -86 24204
rect -66 24182 -62 24204
rect -42 24182 -38 24204
rect -18 24182 -14 24204
rect 6 24182 10 24204
rect 30 24182 34 24204
rect 54 24182 58 24204
rect 78 24182 82 24204
rect 102 24182 106 24204
rect 126 24182 130 24204
rect 150 24182 154 24204
rect 174 24182 178 24204
rect 198 24182 202 24204
rect 222 24182 226 24204
rect 246 24182 250 24204
rect 270 24182 274 24204
rect 294 24182 298 24204
rect 318 24182 322 24204
rect 342 24182 346 24204
rect 366 24182 370 24204
rect 390 24182 394 24204
rect 414 24182 418 24204
rect 438 24182 442 24204
rect 462 24182 466 24204
rect 486 24182 490 24204
rect 510 24182 514 24204
rect 534 24182 538 24204
rect 558 24182 562 24204
rect 582 24182 586 24204
rect 606 24182 610 24204
rect 630 24182 634 24204
rect 654 24182 658 24204
rect 678 24182 682 24204
rect 702 24182 706 24204
rect 726 24182 730 24204
rect 750 24182 754 24204
rect 774 24182 778 24204
rect 798 24182 802 24204
rect 822 24182 826 24204
rect 846 24182 850 24204
rect 870 24182 874 24204
rect 894 24182 898 24204
rect 918 24182 922 24204
rect 942 24182 946 24204
rect 966 24182 970 24204
rect 990 24182 994 24204
rect 1014 24182 1018 24204
rect 1038 24182 1042 24204
rect 1062 24182 1066 24204
rect 1086 24182 1090 24204
rect 1110 24182 1114 24204
rect 1134 24182 1138 24204
rect 1158 24182 1162 24204
rect 1182 24182 1186 24204
rect 1206 24182 1210 24204
rect 1230 24182 1234 24204
rect 1254 24182 1258 24204
rect 1278 24182 1282 24204
rect 1302 24182 1306 24204
rect 1326 24182 1330 24204
rect 1350 24182 1354 24204
rect 1374 24182 1378 24204
rect 1398 24182 1402 24204
rect 1422 24182 1426 24204
rect 1446 24182 1450 24204
rect 1470 24182 1474 24204
rect 1494 24182 1498 24204
rect 1518 24182 1522 24204
rect 1542 24182 1546 24204
rect 1566 24182 1570 24204
rect 1573 24203 1587 24204
rect 1590 24203 1597 24227
rect 1590 24182 1594 24203
rect 1614 24182 1618 24276
rect 1638 24182 1642 24276
rect 1662 24182 1666 24276
rect 1686 24182 1690 24276
rect 1710 24182 1714 24276
rect 1734 24182 1738 24276
rect 1758 24182 1762 24276
rect 1782 24182 1786 24276
rect 1806 24182 1810 24276
rect 1830 24182 1834 24276
rect 1854 24182 1858 24276
rect 1878 24182 1882 24276
rect 1902 24182 1906 24276
rect 1926 24182 1930 24276
rect 1950 24182 1954 24276
rect 1974 24182 1978 24276
rect 1998 24255 2002 24276
rect 1987 24254 2021 24255
rect 2022 24254 2026 24276
rect 2046 24254 2050 24276
rect 2070 24254 2074 24276
rect 2094 24254 2098 24276
rect 2118 24254 2122 24276
rect 2142 24254 2146 24276
rect 2166 24254 2170 24276
rect 2190 24254 2194 24276
rect 2214 24254 2218 24276
rect 2238 24254 2242 24276
rect 2262 24254 2266 24276
rect 2286 24254 2290 24276
rect 2310 24254 2314 24276
rect 2334 24254 2338 24276
rect 2358 24254 2362 24276
rect 2382 24254 2386 24276
rect 2406 24254 2410 24276
rect 2430 24254 2434 24276
rect 2454 24254 2458 24276
rect 2478 24254 2482 24276
rect 2491 24269 2496 24276
rect 2502 24269 2506 24276
rect 2509 24275 2523 24276
rect 2501 24255 2506 24269
rect 2515 24265 2523 24269
rect 2509 24255 2515 24265
rect 2491 24254 2523 24255
rect 1987 24252 2523 24254
rect 1987 24245 1992 24252
rect 1998 24245 2002 24252
rect 1997 24231 2002 24245
rect 1987 24221 1992 24231
rect 1997 24207 2002 24221
rect 1998 24182 2002 24207
rect 2022 24182 2026 24252
rect 2046 24182 2050 24252
rect 2070 24182 2074 24252
rect 2094 24182 2098 24252
rect 2118 24182 2122 24252
rect 2142 24182 2146 24252
rect 2166 24182 2170 24252
rect 2190 24182 2194 24252
rect 2214 24182 2218 24252
rect 2238 24182 2242 24252
rect 2262 24182 2266 24252
rect 2286 24182 2290 24252
rect 2310 24182 2314 24252
rect 2334 24182 2338 24252
rect 2358 24182 2362 24252
rect 2382 24182 2386 24252
rect 2406 24182 2410 24252
rect 2430 24182 2434 24252
rect 2443 24197 2448 24207
rect 2454 24197 2458 24252
rect 2453 24183 2458 24197
rect 2454 24182 2458 24183
rect 2478 24182 2482 24252
rect 2491 24245 2496 24252
rect 2509 24251 2523 24252
rect 2501 24231 2506 24245
rect 2502 24183 2506 24231
rect 2491 24182 2523 24183
rect -2393 24180 2523 24182
rect -2371 24134 -2366 24180
rect -2348 24134 -2343 24180
rect -2325 24134 -2320 24180
rect -2317 24176 -2309 24180
rect -2062 24176 -2054 24180
rect -2154 24172 -2138 24174
rect -2057 24172 -2054 24176
rect -2292 24166 -2054 24172
rect -2052 24166 -2044 24176
rect -2092 24150 -2062 24152
rect -2094 24146 -2062 24150
rect -2000 24134 -1992 24180
rect -1846 24173 -1806 24180
rect -1663 24176 -1655 24180
rect -1846 24166 -1680 24172
rect -1854 24150 -1806 24152
rect -1854 24146 -1680 24150
rect -1642 24134 -1637 24180
rect -1619 24134 -1614 24180
rect -1530 24134 -1526 24180
rect -1506 24134 -1502 24180
rect -1482 24134 -1478 24180
rect -1458 24134 -1454 24180
rect -1434 24134 -1430 24180
rect -1410 24134 -1406 24180
rect -1386 24134 -1382 24180
rect -1362 24134 -1358 24180
rect -1338 24134 -1334 24180
rect -1314 24134 -1310 24180
rect -1290 24134 -1286 24180
rect -1266 24134 -1262 24180
rect -1242 24134 -1238 24180
rect -1218 24134 -1214 24180
rect -1194 24134 -1190 24180
rect -1170 24134 -1166 24180
rect -1146 24134 -1142 24180
rect -1122 24134 -1118 24180
rect -1098 24134 -1094 24180
rect -1074 24134 -1070 24180
rect -1050 24134 -1046 24180
rect -1026 24134 -1022 24180
rect -1002 24134 -998 24180
rect -978 24134 -974 24180
rect -954 24134 -950 24180
rect -930 24134 -926 24180
rect -906 24134 -902 24180
rect -882 24134 -878 24180
rect -858 24134 -854 24180
rect -834 24134 -830 24180
rect -810 24134 -806 24180
rect -786 24134 -782 24180
rect -762 24134 -758 24180
rect -738 24134 -734 24180
rect -714 24134 -710 24180
rect -690 24134 -686 24180
rect -666 24134 -662 24180
rect -642 24134 -638 24180
rect -618 24134 -614 24180
rect -594 24134 -590 24180
rect -570 24134 -566 24180
rect -546 24134 -542 24180
rect -522 24134 -518 24180
rect -498 24134 -494 24180
rect -474 24134 -470 24180
rect -450 24134 -446 24180
rect -426 24134 -422 24180
rect -402 24134 -398 24180
rect -378 24134 -374 24180
rect -354 24134 -350 24180
rect -330 24134 -326 24180
rect -306 24134 -302 24180
rect -282 24134 -278 24180
rect -258 24134 -254 24180
rect -234 24134 -230 24180
rect -210 24134 -206 24180
rect -186 24134 -182 24180
rect -162 24134 -158 24180
rect -138 24134 -134 24180
rect -114 24134 -110 24180
rect -90 24134 -86 24180
rect -66 24134 -62 24180
rect -42 24134 -38 24180
rect -18 24134 -14 24180
rect 6 24134 10 24180
rect 30 24134 34 24180
rect 54 24134 58 24180
rect 78 24134 82 24180
rect 102 24134 106 24180
rect 126 24134 130 24180
rect 150 24134 154 24180
rect 174 24134 178 24180
rect 198 24134 202 24180
rect 222 24134 226 24180
rect 246 24134 250 24180
rect 270 24134 274 24180
rect 294 24134 298 24180
rect 318 24134 322 24180
rect 342 24134 346 24180
rect 366 24134 370 24180
rect 390 24134 394 24180
rect 414 24134 418 24180
rect 438 24134 442 24180
rect 462 24134 466 24180
rect 486 24134 490 24180
rect 510 24134 514 24180
rect 534 24134 538 24180
rect 558 24134 562 24180
rect 582 24134 586 24180
rect 606 24134 610 24180
rect 630 24134 634 24180
rect 654 24134 658 24180
rect 678 24134 682 24180
rect 702 24134 706 24180
rect 726 24134 730 24180
rect 750 24134 754 24180
rect 774 24134 778 24180
rect 798 24134 802 24180
rect 822 24134 826 24180
rect 846 24134 850 24180
rect 870 24134 874 24180
rect 894 24134 898 24180
rect 918 24134 922 24180
rect 942 24134 946 24180
rect 966 24134 970 24180
rect 990 24134 994 24180
rect 1014 24134 1018 24180
rect 1038 24134 1042 24180
rect 1062 24134 1066 24180
rect 1086 24134 1090 24180
rect 1110 24134 1114 24180
rect 1134 24134 1138 24180
rect 1158 24134 1162 24180
rect 1182 24134 1186 24180
rect 1206 24134 1210 24180
rect 1230 24134 1234 24180
rect 1254 24134 1258 24180
rect 1278 24134 1282 24180
rect 1302 24134 1306 24180
rect 1326 24134 1330 24180
rect 1350 24134 1354 24180
rect 1374 24134 1378 24180
rect 1398 24134 1402 24180
rect 1422 24134 1426 24180
rect 1446 24134 1450 24180
rect 1470 24134 1474 24180
rect 1494 24134 1498 24180
rect 1518 24134 1522 24180
rect 1542 24134 1546 24180
rect 1566 24134 1570 24180
rect 1590 24134 1594 24180
rect 1614 24134 1618 24180
rect 1638 24134 1642 24180
rect 1662 24134 1666 24180
rect 1686 24134 1690 24180
rect 1710 24134 1714 24180
rect 1734 24134 1738 24180
rect 1747 24149 1752 24159
rect 1758 24149 1762 24180
rect 1757 24135 1762 24149
rect 1747 24134 1781 24135
rect -2393 24132 1781 24134
rect -2371 24110 -2366 24132
rect -2348 24110 -2343 24132
rect -2325 24110 -2320 24132
rect -2072 24130 -2036 24131
rect -2072 24124 -2054 24130
rect -2309 24116 -2301 24124
rect -2317 24110 -2309 24116
rect -2092 24115 -2062 24120
rect -2000 24111 -1992 24132
rect -1938 24131 -1906 24132
rect -1920 24130 -1906 24131
rect -1806 24124 -1680 24130
rect -1854 24115 -1806 24120
rect -1655 24116 -1647 24124
rect -1982 24111 -1966 24112
rect -2000 24110 -1966 24111
rect -1846 24110 -1806 24113
rect -1663 24110 -1655 24116
rect -1642 24110 -1637 24132
rect -1619 24110 -1614 24132
rect -1530 24110 -1526 24132
rect -1506 24110 -1502 24132
rect -1482 24110 -1478 24132
rect -1458 24110 -1454 24132
rect -1434 24110 -1430 24132
rect -1410 24110 -1406 24132
rect -1386 24110 -1382 24132
rect -1362 24110 -1358 24132
rect -1338 24110 -1334 24132
rect -1314 24110 -1310 24132
rect -1290 24110 -1286 24132
rect -1266 24110 -1262 24132
rect -1242 24110 -1238 24132
rect -1218 24110 -1214 24132
rect -1194 24110 -1190 24132
rect -1170 24110 -1166 24132
rect -1146 24110 -1142 24132
rect -1122 24110 -1118 24132
rect -1098 24110 -1094 24132
rect -1074 24110 -1070 24132
rect -1050 24110 -1046 24132
rect -1026 24110 -1022 24132
rect -1002 24110 -998 24132
rect -978 24110 -974 24132
rect -954 24110 -950 24132
rect -930 24110 -926 24132
rect -906 24110 -902 24132
rect -882 24110 -878 24132
rect -858 24110 -854 24132
rect -834 24110 -830 24132
rect -810 24110 -806 24132
rect -786 24110 -782 24132
rect -762 24110 -758 24132
rect -738 24110 -734 24132
rect -714 24110 -710 24132
rect -690 24110 -686 24132
rect -666 24110 -662 24132
rect -642 24110 -638 24132
rect -618 24110 -614 24132
rect -594 24110 -590 24132
rect -570 24110 -566 24132
rect -546 24110 -542 24132
rect -522 24110 -518 24132
rect -498 24110 -494 24132
rect -474 24110 -470 24132
rect -450 24110 -446 24132
rect -426 24110 -422 24132
rect -402 24110 -398 24132
rect -378 24110 -374 24132
rect -354 24110 -350 24132
rect -330 24110 -326 24132
rect -306 24110 -302 24132
rect -282 24110 -278 24132
rect -258 24110 -254 24132
rect -234 24110 -230 24132
rect -210 24110 -206 24132
rect -186 24110 -182 24132
rect -162 24110 -158 24132
rect -138 24110 -134 24132
rect -114 24110 -110 24132
rect -90 24110 -86 24132
rect -66 24110 -62 24132
rect -42 24110 -38 24132
rect -18 24110 -14 24132
rect 6 24110 10 24132
rect 30 24110 34 24132
rect 54 24110 58 24132
rect 78 24110 82 24132
rect 102 24110 106 24132
rect 126 24110 130 24132
rect 150 24110 154 24132
rect 174 24110 178 24132
rect 198 24110 202 24132
rect 222 24110 226 24132
rect 246 24110 250 24132
rect 270 24110 274 24132
rect 294 24110 298 24132
rect 318 24110 322 24132
rect 342 24110 346 24132
rect 366 24110 370 24132
rect 390 24110 394 24132
rect 414 24110 418 24132
rect 438 24110 442 24132
rect 462 24110 466 24132
rect 486 24110 490 24132
rect 510 24110 514 24132
rect 534 24110 538 24132
rect 558 24110 562 24132
rect 582 24110 586 24132
rect 606 24110 610 24132
rect 630 24110 634 24132
rect 654 24110 658 24132
rect 678 24110 682 24132
rect 702 24110 706 24132
rect 726 24110 730 24132
rect 750 24110 754 24132
rect 774 24110 778 24132
rect 798 24110 802 24132
rect 822 24110 826 24132
rect 846 24110 850 24132
rect 870 24110 874 24132
rect 894 24110 898 24132
rect 918 24110 922 24132
rect 942 24110 946 24132
rect 966 24110 970 24132
rect 990 24110 994 24132
rect 1014 24110 1018 24132
rect 1038 24110 1042 24132
rect 1062 24110 1066 24132
rect 1086 24110 1090 24132
rect 1110 24110 1114 24132
rect 1134 24110 1138 24132
rect 1158 24110 1162 24132
rect 1182 24110 1186 24132
rect 1206 24110 1210 24132
rect 1230 24110 1234 24132
rect 1254 24110 1258 24132
rect 1278 24110 1282 24132
rect 1302 24110 1306 24132
rect 1326 24110 1330 24132
rect 1350 24110 1354 24132
rect 1374 24110 1378 24132
rect 1398 24110 1402 24132
rect 1422 24110 1426 24132
rect 1446 24110 1450 24132
rect 1470 24110 1474 24132
rect 1494 24110 1498 24132
rect 1518 24110 1522 24132
rect 1542 24110 1546 24132
rect 1566 24110 1570 24132
rect 1590 24110 1594 24132
rect 1614 24110 1618 24132
rect 1638 24110 1642 24132
rect 1662 24110 1666 24132
rect 1686 24110 1690 24132
rect 1710 24110 1714 24132
rect 1734 24110 1738 24132
rect 1747 24125 1752 24132
rect 1757 24111 1762 24125
rect 1758 24110 1762 24111
rect 1782 24110 1786 24180
rect 1806 24110 1810 24180
rect 1830 24110 1834 24180
rect 1854 24110 1858 24180
rect 1878 24110 1882 24180
rect 1902 24110 1906 24180
rect 1926 24110 1930 24180
rect 1950 24110 1954 24180
rect 1974 24110 1978 24180
rect 1998 24110 2002 24180
rect 2022 24179 2026 24180
rect 2022 24158 2029 24179
rect 2046 24158 2050 24180
rect 2070 24158 2074 24180
rect 2094 24158 2098 24180
rect 2118 24158 2122 24180
rect 2142 24158 2146 24180
rect 2166 24158 2170 24180
rect 2190 24158 2194 24180
rect 2214 24158 2218 24180
rect 2238 24158 2242 24180
rect 2262 24158 2266 24180
rect 2286 24158 2290 24180
rect 2310 24158 2314 24180
rect 2334 24158 2338 24180
rect 2358 24158 2362 24180
rect 2382 24158 2386 24180
rect 2406 24158 2410 24180
rect 2430 24158 2434 24180
rect 2454 24158 2458 24180
rect 2478 24158 2482 24180
rect 2491 24173 2496 24180
rect 2502 24173 2506 24180
rect 2509 24179 2523 24180
rect 2501 24159 2506 24173
rect 2515 24169 2523 24173
rect 2509 24159 2515 24169
rect 2491 24158 2523 24159
rect 2005 24156 2523 24158
rect 2005 24155 2019 24156
rect 2022 24131 2029 24156
rect 2022 24110 2026 24131
rect 2046 24110 2050 24156
rect 2070 24110 2074 24156
rect 2094 24110 2098 24156
rect 2118 24110 2122 24156
rect 2142 24110 2146 24156
rect 2166 24110 2170 24156
rect 2190 24110 2194 24156
rect 2214 24110 2218 24156
rect 2238 24110 2242 24156
rect 2262 24110 2266 24156
rect 2286 24110 2290 24156
rect 2310 24110 2314 24156
rect 2334 24110 2338 24156
rect 2358 24110 2362 24156
rect 2382 24110 2386 24156
rect 2406 24110 2410 24156
rect 2430 24110 2434 24156
rect 2454 24110 2458 24156
rect 2478 24131 2482 24156
rect 2491 24149 2496 24156
rect 2509 24155 2523 24156
rect 2501 24135 2506 24149
rect -2393 24108 2475 24110
rect -2371 24086 -2366 24108
rect -2348 24086 -2343 24108
rect -2325 24086 -2320 24108
rect -2000 24106 -1966 24108
rect -2309 24088 -2301 24096
rect -2062 24095 -2054 24102
rect -2092 24088 -2084 24095
rect -2062 24088 -2026 24090
rect -2317 24086 -2309 24088
rect -2062 24086 -2012 24088
rect -2000 24086 -1992 24106
rect -1982 24105 -1966 24106
rect -1846 24104 -1806 24108
rect -1846 24097 -1798 24102
rect -1806 24095 -1798 24097
rect -1854 24093 -1846 24095
rect -1854 24088 -1806 24093
rect -1655 24088 -1647 24096
rect -1864 24086 -1796 24087
rect -1663 24086 -1655 24088
rect -1642 24086 -1637 24108
rect -1619 24086 -1614 24108
rect -1530 24086 -1526 24108
rect -1506 24086 -1502 24108
rect -1482 24086 -1478 24108
rect -1458 24086 -1454 24108
rect -1434 24086 -1430 24108
rect -1410 24086 -1406 24108
rect -1386 24086 -1382 24108
rect -1362 24086 -1358 24108
rect -1338 24086 -1334 24108
rect -1314 24086 -1310 24108
rect -1290 24086 -1286 24108
rect -1266 24086 -1262 24108
rect -1242 24086 -1238 24108
rect -1218 24086 -1214 24108
rect -1194 24086 -1190 24108
rect -1170 24086 -1166 24108
rect -1146 24086 -1142 24108
rect -1122 24086 -1118 24108
rect -1098 24086 -1094 24108
rect -1074 24086 -1070 24108
rect -1050 24086 -1046 24108
rect -1026 24086 -1022 24108
rect -1002 24086 -998 24108
rect -978 24086 -974 24108
rect -954 24086 -950 24108
rect -930 24086 -926 24108
rect -906 24086 -902 24108
rect -882 24086 -878 24108
rect -858 24086 -854 24108
rect -834 24086 -830 24108
rect -810 24086 -806 24108
rect -786 24086 -782 24108
rect -762 24086 -758 24108
rect -738 24086 -734 24108
rect -714 24086 -710 24108
rect -690 24086 -686 24108
rect -666 24086 -662 24108
rect -642 24086 -638 24108
rect -618 24086 -614 24108
rect -594 24086 -590 24108
rect -570 24086 -566 24108
rect -546 24086 -542 24108
rect -522 24086 -518 24108
rect -498 24086 -494 24108
rect -474 24086 -470 24108
rect -450 24086 -446 24108
rect -426 24086 -422 24108
rect -402 24086 -398 24108
rect -378 24086 -374 24108
rect -354 24086 -350 24108
rect -330 24086 -326 24108
rect -306 24086 -302 24108
rect -282 24086 -278 24108
rect -258 24086 -254 24108
rect -234 24086 -230 24108
rect -210 24086 -206 24108
rect -186 24086 -182 24108
rect -162 24086 -158 24108
rect -138 24086 -134 24108
rect -114 24086 -110 24108
rect -90 24086 -86 24108
rect -66 24086 -62 24108
rect -42 24086 -38 24108
rect -18 24086 -14 24108
rect 6 24086 10 24108
rect 30 24086 34 24108
rect 54 24086 58 24108
rect 78 24086 82 24108
rect 102 24086 106 24108
rect 126 24086 130 24108
rect 150 24086 154 24108
rect 174 24086 178 24108
rect 198 24086 202 24108
rect 222 24086 226 24108
rect 246 24086 250 24108
rect 270 24086 274 24108
rect 294 24086 298 24108
rect 318 24086 322 24108
rect 342 24086 346 24108
rect 366 24086 370 24108
rect 390 24086 394 24108
rect 414 24086 418 24108
rect 438 24086 442 24108
rect 462 24086 466 24108
rect 486 24086 490 24108
rect 510 24086 514 24108
rect 534 24086 538 24108
rect 558 24086 562 24108
rect 582 24086 586 24108
rect 606 24086 610 24108
rect 630 24086 634 24108
rect 654 24086 658 24108
rect 678 24086 682 24108
rect 702 24086 706 24108
rect 726 24086 730 24108
rect 750 24086 754 24108
rect 774 24086 778 24108
rect 798 24086 802 24108
rect 822 24086 826 24108
rect 846 24086 850 24108
rect 870 24086 874 24108
rect 894 24086 898 24108
rect 918 24086 922 24108
rect 942 24086 946 24108
rect 966 24086 970 24108
rect 990 24086 994 24108
rect 1014 24086 1018 24108
rect 1038 24086 1042 24108
rect 1062 24086 1066 24108
rect 1086 24086 1090 24108
rect 1110 24086 1114 24108
rect 1134 24086 1138 24108
rect 1158 24086 1162 24108
rect 1182 24086 1186 24108
rect 1206 24086 1210 24108
rect 1230 24086 1234 24108
rect 1254 24086 1258 24108
rect 1278 24086 1282 24108
rect 1302 24086 1306 24108
rect 1326 24086 1330 24108
rect 1350 24086 1354 24108
rect 1374 24086 1378 24108
rect 1398 24086 1402 24108
rect 1422 24086 1426 24108
rect 1446 24086 1450 24108
rect 1470 24086 1474 24108
rect 1494 24086 1498 24108
rect 1518 24086 1522 24108
rect 1542 24086 1546 24108
rect 1566 24086 1570 24108
rect 1590 24086 1594 24108
rect 1614 24086 1618 24108
rect 1638 24086 1642 24108
rect 1662 24086 1666 24108
rect 1686 24086 1690 24108
rect 1710 24086 1714 24108
rect 1734 24086 1738 24108
rect 1758 24086 1762 24108
rect 1782 24086 1786 24108
rect 1806 24086 1810 24108
rect 1830 24086 1834 24108
rect 1854 24086 1858 24108
rect 1878 24086 1882 24108
rect 1902 24086 1906 24108
rect 1926 24086 1930 24108
rect 1950 24086 1954 24108
rect 1974 24086 1978 24108
rect 1998 24086 2002 24108
rect 2022 24086 2026 24108
rect 2046 24086 2050 24108
rect 2070 24086 2074 24108
rect 2094 24086 2098 24108
rect 2118 24086 2122 24108
rect 2142 24086 2146 24108
rect 2166 24086 2170 24108
rect 2190 24086 2194 24108
rect 2214 24086 2218 24108
rect 2238 24086 2242 24108
rect 2262 24086 2266 24108
rect 2286 24086 2290 24108
rect 2310 24086 2314 24108
rect 2334 24086 2338 24108
rect 2358 24086 2362 24108
rect 2382 24086 2386 24108
rect 2406 24086 2410 24108
rect 2430 24086 2434 24108
rect 2454 24086 2458 24108
rect 2461 24107 2475 24108
rect 2478 24107 2485 24131
rect 2478 24087 2482 24107
rect 2491 24101 2496 24111
rect 2502 24101 2506 24135
rect 2501 24087 2506 24101
rect 2515 24097 2523 24101
rect 2509 24087 2515 24097
rect 2467 24086 2501 24087
rect -2393 24084 2501 24086
rect -2371 24038 -2366 24084
rect -2348 24038 -2343 24084
rect -2325 24048 -2320 24084
rect -2317 24080 -2309 24084
rect -2062 24080 -2054 24084
rect -2154 24076 -2138 24078
rect -2057 24076 -2054 24080
rect -2292 24070 -2054 24076
rect -2052 24070 -2044 24080
rect -2092 24054 -2062 24056
rect -2094 24050 -2062 24054
rect -2325 24038 -2317 24048
rect -2095 24040 -2084 24044
rect -2000 24041 -1992 24084
rect -1846 24077 -1806 24084
rect -1663 24080 -1655 24084
rect -1846 24070 -1680 24076
rect -1854 24054 -1806 24056
rect -1854 24050 -1680 24054
rect -2119 24038 -2069 24040
rect -2054 24038 -1892 24041
rect -1671 24038 -1663 24048
rect -1642 24038 -1637 24084
rect -1619 24038 -1614 24084
rect -1530 24038 -1526 24084
rect -1506 24038 -1502 24084
rect -1482 24038 -1478 24084
rect -1458 24038 -1454 24084
rect -1434 24038 -1430 24084
rect -1410 24038 -1406 24084
rect -1386 24038 -1382 24084
rect -1362 24038 -1358 24084
rect -1338 24038 -1334 24084
rect -1314 24038 -1310 24084
rect -1290 24038 -1286 24084
rect -1266 24038 -1262 24084
rect -1242 24038 -1238 24084
rect -1218 24038 -1214 24084
rect -1194 24038 -1190 24084
rect -1170 24038 -1166 24084
rect -1146 24038 -1142 24084
rect -1122 24038 -1118 24084
rect -1098 24038 -1094 24084
rect -1074 24038 -1070 24084
rect -1050 24038 -1046 24084
rect -1026 24038 -1022 24084
rect -1002 24038 -998 24084
rect -978 24038 -974 24084
rect -954 24038 -950 24084
rect -930 24038 -926 24084
rect -906 24038 -902 24084
rect -882 24038 -878 24084
rect -858 24038 -854 24084
rect -834 24038 -830 24084
rect -810 24038 -806 24084
rect -786 24038 -782 24084
rect -762 24038 -758 24084
rect -738 24038 -734 24084
rect -714 24038 -710 24084
rect -690 24038 -686 24084
rect -666 24038 -662 24084
rect -642 24038 -638 24084
rect -618 24038 -614 24084
rect -594 24038 -590 24084
rect -570 24038 -566 24084
rect -546 24038 -542 24084
rect -522 24038 -518 24084
rect -498 24038 -494 24084
rect -474 24038 -470 24084
rect -450 24038 -446 24084
rect -426 24038 -422 24084
rect -402 24038 -398 24084
rect -378 24038 -374 24084
rect -354 24038 -350 24084
rect -330 24038 -326 24084
rect -306 24038 -302 24084
rect -282 24038 -278 24084
rect -258 24038 -254 24084
rect -234 24038 -230 24084
rect -210 24038 -206 24084
rect -186 24038 -182 24084
rect -162 24038 -158 24084
rect -138 24038 -134 24084
rect -114 24038 -110 24084
rect -90 24038 -86 24084
rect -66 24038 -62 24084
rect -42 24038 -38 24084
rect -18 24038 -14 24084
rect 6 24038 10 24084
rect 30 24038 34 24084
rect 54 24038 58 24084
rect 78 24038 82 24084
rect 102 24038 106 24084
rect 126 24038 130 24084
rect 150 24038 154 24084
rect 174 24038 178 24084
rect 198 24038 202 24084
rect 222 24038 226 24084
rect 246 24038 250 24084
rect 270 24038 274 24084
rect 294 24038 298 24084
rect 318 24038 322 24084
rect 342 24038 346 24084
rect 366 24038 370 24084
rect 390 24038 394 24084
rect 414 24038 418 24084
rect 438 24038 442 24084
rect 462 24038 466 24084
rect 486 24038 490 24084
rect 510 24038 514 24084
rect 534 24038 538 24084
rect 558 24038 562 24084
rect 582 24038 586 24084
rect 606 24038 610 24084
rect 630 24038 634 24084
rect 654 24038 658 24084
rect 678 24038 682 24084
rect 702 24038 706 24084
rect 726 24038 730 24084
rect 750 24038 754 24084
rect 774 24038 778 24084
rect 798 24038 802 24084
rect 822 24038 826 24084
rect 846 24038 850 24084
rect 870 24038 874 24084
rect 894 24038 898 24084
rect 918 24038 922 24084
rect 942 24038 946 24084
rect 966 24038 970 24084
rect 990 24038 994 24084
rect 1014 24038 1018 24084
rect 1038 24038 1042 24084
rect 1062 24038 1066 24084
rect 1086 24038 1090 24084
rect 1110 24038 1114 24084
rect 1134 24038 1138 24084
rect 1158 24038 1162 24084
rect 1182 24038 1186 24084
rect 1206 24038 1210 24084
rect 1230 24038 1234 24084
rect 1254 24038 1258 24084
rect 1278 24038 1282 24084
rect 1302 24038 1306 24084
rect 1326 24038 1330 24084
rect 1350 24038 1354 24084
rect 1374 24038 1378 24084
rect 1398 24038 1402 24084
rect 1422 24038 1426 24084
rect 1446 24038 1450 24084
rect 1470 24038 1474 24084
rect 1494 24038 1498 24084
rect 1518 24038 1522 24084
rect 1542 24038 1546 24084
rect 1566 24038 1570 24084
rect 1590 24038 1594 24084
rect 1614 24038 1618 24084
rect 1638 24038 1642 24084
rect 1662 24038 1666 24084
rect 1686 24038 1690 24084
rect 1710 24038 1714 24084
rect 1734 24038 1738 24084
rect 1758 24038 1762 24084
rect 1782 24083 1786 24084
rect -2393 24036 1779 24038
rect -2371 24014 -2366 24036
rect -2348 24014 -2343 24036
rect -2325 24032 -2317 24036
rect -2325 24016 -2320 24032
rect -2309 24020 -2301 24032
rect -2095 24030 -2084 24036
rect -2054 24035 -1906 24036
rect -2054 24034 -2036 24035
rect -2084 24028 -2079 24030
rect -2317 24016 -2309 24020
rect -2092 24019 -2079 24026
rect -2000 24022 -1992 24035
rect -1920 24034 -1906 24035
rect -1671 24032 -1663 24036
rect -1846 24028 -1806 24030
rect -1854 24022 -1806 24026
rect -2054 24019 -1982 24022
rect -1966 24019 -1806 24022
rect -1655 24020 -1647 24032
rect -2003 24016 -1992 24019
rect -1904 24017 -1902 24019
rect -1854 24017 -1846 24019
rect -2325 24014 -2317 24016
rect -2033 24014 -1992 24016
rect -1854 24015 -1806 24017
rect -1663 24016 -1655 24020
rect -1864 24014 -1796 24015
rect -1671 24014 -1663 24016
rect -1642 24014 -1637 24036
rect -1619 24014 -1614 24036
rect -1530 24014 -1526 24036
rect -1506 24014 -1502 24036
rect -1482 24014 -1478 24036
rect -1458 24014 -1454 24036
rect -1434 24014 -1430 24036
rect -1410 24014 -1406 24036
rect -1386 24014 -1382 24036
rect -1362 24014 -1358 24036
rect -1338 24014 -1334 24036
rect -1314 24014 -1310 24036
rect -1290 24014 -1286 24036
rect -1266 24014 -1262 24036
rect -1242 24014 -1238 24036
rect -1218 24014 -1214 24036
rect -1194 24014 -1190 24036
rect -1170 24014 -1166 24036
rect -1146 24014 -1142 24036
rect -1122 24014 -1118 24036
rect -1098 24014 -1094 24036
rect -1074 24014 -1070 24036
rect -1050 24014 -1046 24036
rect -1026 24014 -1022 24036
rect -1002 24014 -998 24036
rect -978 24014 -974 24036
rect -954 24014 -950 24036
rect -930 24014 -926 24036
rect -906 24014 -902 24036
rect -882 24014 -878 24036
rect -858 24014 -854 24036
rect -834 24014 -830 24036
rect -810 24014 -806 24036
rect -786 24014 -782 24036
rect -762 24014 -758 24036
rect -738 24014 -734 24036
rect -714 24014 -710 24036
rect -690 24014 -686 24036
rect -666 24014 -662 24036
rect -642 24014 -638 24036
rect -618 24014 -614 24036
rect -594 24014 -590 24036
rect -570 24014 -566 24036
rect -546 24014 -542 24036
rect -522 24014 -518 24036
rect -498 24014 -494 24036
rect -474 24014 -470 24036
rect -450 24014 -446 24036
rect -426 24014 -422 24036
rect -402 24014 -398 24036
rect -378 24014 -374 24036
rect -354 24014 -350 24036
rect -330 24014 -326 24036
rect -306 24014 -302 24036
rect -282 24014 -278 24036
rect -258 24014 -254 24036
rect -234 24014 -230 24036
rect -210 24014 -206 24036
rect -186 24014 -182 24036
rect -162 24014 -158 24036
rect -138 24014 -134 24036
rect -114 24014 -110 24036
rect -90 24014 -86 24036
rect -66 24014 -62 24036
rect -42 24014 -38 24036
rect -18 24014 -14 24036
rect 6 24014 10 24036
rect 30 24014 34 24036
rect 54 24014 58 24036
rect 78 24014 82 24036
rect 102 24014 106 24036
rect 126 24014 130 24036
rect 150 24014 154 24036
rect 174 24014 178 24036
rect 198 24014 202 24036
rect 222 24014 226 24036
rect 246 24014 250 24036
rect 270 24014 274 24036
rect 294 24014 298 24036
rect 318 24014 322 24036
rect 342 24014 346 24036
rect 366 24014 370 24036
rect 390 24014 394 24036
rect 414 24014 418 24036
rect 438 24014 442 24036
rect 462 24014 466 24036
rect 486 24014 490 24036
rect 510 24014 514 24036
rect 534 24014 538 24036
rect 558 24014 562 24036
rect 582 24014 586 24036
rect 606 24014 610 24036
rect 630 24014 634 24036
rect 654 24014 658 24036
rect 678 24014 682 24036
rect 702 24014 706 24036
rect 726 24014 730 24036
rect 750 24014 754 24036
rect 774 24014 778 24036
rect 798 24014 802 24036
rect 822 24014 826 24036
rect 846 24014 850 24036
rect 870 24014 874 24036
rect 894 24014 898 24036
rect 918 24014 922 24036
rect 942 24014 946 24036
rect 966 24014 970 24036
rect 990 24014 994 24036
rect 1014 24014 1018 24036
rect 1038 24014 1042 24036
rect 1062 24014 1066 24036
rect 1086 24014 1090 24036
rect 1110 24014 1114 24036
rect 1134 24014 1138 24036
rect 1158 24014 1162 24036
rect 1182 24014 1186 24036
rect 1206 24014 1210 24036
rect 1230 24014 1234 24036
rect 1254 24014 1258 24036
rect 1278 24014 1282 24036
rect 1302 24014 1306 24036
rect 1326 24014 1330 24036
rect 1350 24014 1354 24036
rect 1374 24014 1378 24036
rect 1398 24015 1402 24036
rect 1387 24014 1421 24015
rect -2393 24012 1421 24014
rect -2371 23990 -2366 24012
rect -2348 23990 -2343 24012
rect -2325 24004 -2317 24012
rect -2079 24009 -2018 24012
rect -2003 24011 -1966 24012
rect -2000 24010 -1982 24011
rect -2000 24009 -1992 24010
rect -2084 24005 -2009 24009
rect -2028 24004 -2009 24005
rect -2000 24005 -1854 24009
rect -1846 24005 -1798 24012
rect -2325 23990 -2320 24004
rect -2309 23992 -2301 24004
rect -2028 24002 -2018 24004
rect -2092 23992 -2084 23999
rect -2023 23995 -2014 24002
rect -2000 23995 -1992 24005
rect -1671 24004 -1663 24012
rect -1846 24001 -1806 24003
rect -1854 23995 -1806 23999
rect -2054 23992 -1806 23995
rect -1655 23992 -1647 24004
rect -2317 23990 -2309 23992
rect -2054 23990 -2024 23992
rect -2000 23990 -1992 23992
rect -1663 23990 -1655 23992
rect -1642 23990 -1637 24012
rect -1619 23990 -1614 24012
rect -1530 23990 -1526 24012
rect -1506 23990 -1502 24012
rect -1482 23990 -1478 24012
rect -1458 23990 -1454 24012
rect -1434 23990 -1430 24012
rect -1410 23990 -1406 24012
rect -1386 23990 -1382 24012
rect -1362 23990 -1358 24012
rect -1338 23990 -1334 24012
rect -1314 23990 -1310 24012
rect -1290 23990 -1286 24012
rect -1266 23990 -1262 24012
rect -1242 23990 -1238 24012
rect -1218 23990 -1214 24012
rect -1194 23990 -1190 24012
rect -1170 23990 -1166 24012
rect -1146 23990 -1142 24012
rect -1122 23990 -1118 24012
rect -1098 23990 -1094 24012
rect -1074 23990 -1070 24012
rect -1050 23990 -1046 24012
rect -1026 23990 -1022 24012
rect -1002 23990 -998 24012
rect -978 23990 -974 24012
rect -954 23990 -950 24012
rect -930 23990 -926 24012
rect -906 23990 -902 24012
rect -882 23990 -878 24012
rect -858 23990 -854 24012
rect -834 23990 -830 24012
rect -810 23990 -806 24012
rect -786 23990 -782 24012
rect -762 23990 -758 24012
rect -738 23990 -734 24012
rect -714 23990 -710 24012
rect -690 23990 -686 24012
rect -666 23990 -662 24012
rect -642 23990 -638 24012
rect -618 23990 -614 24012
rect -594 23990 -590 24012
rect -570 23990 -566 24012
rect -546 23990 -542 24012
rect -522 23990 -518 24012
rect -498 23990 -494 24012
rect -474 23990 -470 24012
rect -450 23990 -446 24012
rect -426 23990 -422 24012
rect -402 23990 -398 24012
rect -378 23990 -374 24012
rect -354 23990 -350 24012
rect -330 23990 -326 24012
rect -306 23990 -302 24012
rect -282 23990 -278 24012
rect -258 23990 -254 24012
rect -234 23990 -230 24012
rect -210 23990 -206 24012
rect -186 23990 -182 24012
rect -162 23990 -158 24012
rect -138 23990 -134 24012
rect -114 23990 -110 24012
rect -90 23990 -86 24012
rect -66 23990 -62 24012
rect -42 23990 -38 24012
rect -18 23990 -14 24012
rect 6 23990 10 24012
rect 30 23990 34 24012
rect 54 23990 58 24012
rect 78 23990 82 24012
rect 102 23990 106 24012
rect 126 23990 130 24012
rect 150 23990 154 24012
rect 174 23990 178 24012
rect 198 23990 202 24012
rect 222 23990 226 24012
rect 246 23990 250 24012
rect 270 23990 274 24012
rect 294 23990 298 24012
rect 318 23990 322 24012
rect 342 23990 346 24012
rect 366 23990 370 24012
rect 390 23990 394 24012
rect 414 23990 418 24012
rect 438 23990 442 24012
rect 462 23990 466 24012
rect 486 23990 490 24012
rect 510 23990 514 24012
rect 534 23990 538 24012
rect 558 23990 562 24012
rect 582 23990 586 24012
rect 606 23990 610 24012
rect 630 23990 634 24012
rect 654 23990 658 24012
rect 678 23990 682 24012
rect 702 23990 706 24012
rect 726 23990 730 24012
rect 750 23990 754 24012
rect 774 23990 778 24012
rect 798 23990 802 24012
rect 822 23990 826 24012
rect 846 23990 850 24012
rect 870 23990 874 24012
rect 894 23990 898 24012
rect 918 23990 922 24012
rect 942 23990 946 24012
rect 966 23990 970 24012
rect 990 23990 994 24012
rect 1014 23990 1018 24012
rect 1038 23990 1042 24012
rect 1062 23990 1066 24012
rect 1086 23990 1090 24012
rect 1110 23990 1114 24012
rect 1134 23990 1138 24012
rect 1158 23990 1162 24012
rect 1182 23990 1186 24012
rect 1206 23990 1210 24012
rect 1230 23990 1234 24012
rect 1254 23990 1258 24012
rect 1278 23990 1282 24012
rect 1302 23990 1306 24012
rect 1326 23990 1330 24012
rect 1350 23990 1354 24012
rect 1374 23990 1378 24012
rect 1387 24005 1392 24012
rect 1398 24005 1402 24012
rect 1397 23991 1402 24005
rect 1398 23990 1402 23991
rect 1422 23990 1426 24036
rect 1446 23990 1450 24036
rect 1470 23990 1474 24036
rect 1494 23990 1498 24036
rect 1518 23990 1522 24036
rect 1542 23990 1546 24036
rect 1566 23990 1570 24036
rect 1590 23990 1594 24036
rect 1614 23990 1618 24036
rect 1638 23990 1642 24036
rect 1662 23990 1666 24036
rect 1686 23990 1690 24036
rect 1710 23990 1714 24036
rect 1734 23990 1738 24036
rect 1758 23990 1762 24036
rect 1765 24035 1779 24036
rect 1782 24035 1789 24083
rect 1782 23990 1786 24035
rect 1806 23990 1810 24084
rect 1830 23990 1834 24084
rect 1854 23990 1858 24084
rect 1878 23990 1882 24084
rect 1902 23990 1906 24084
rect 1926 23990 1930 24084
rect 1950 23990 1954 24084
rect 1974 23990 1978 24084
rect 1998 23990 2002 24084
rect 2022 23990 2026 24084
rect 2046 23990 2050 24084
rect 2070 23990 2074 24084
rect 2094 23990 2098 24084
rect 2118 23990 2122 24084
rect 2142 23990 2146 24084
rect 2166 23990 2170 24084
rect 2190 23990 2194 24084
rect 2214 23990 2218 24084
rect 2238 23990 2242 24084
rect 2262 23990 2266 24084
rect 2286 23990 2290 24084
rect 2310 23990 2314 24084
rect 2334 23990 2338 24084
rect 2358 23990 2362 24084
rect 2382 23990 2386 24084
rect 2406 23990 2410 24084
rect 2430 24063 2434 24084
rect 2419 24062 2453 24063
rect 2454 24062 2458 24084
rect 2467 24077 2472 24084
rect 2478 24077 2482 24084
rect 2477 24063 2482 24077
rect 2467 24062 2501 24063
rect 2419 24060 2501 24062
rect 2419 24053 2424 24060
rect 2430 24053 2434 24060
rect 2429 24039 2434 24053
rect 2419 24029 2424 24039
rect 2429 24015 2434 24029
rect 2430 23990 2434 24015
rect 2454 23990 2458 24060
rect 2467 24053 2472 24060
rect 2477 24039 2482 24053
rect 2478 23991 2482 24039
rect 2467 23990 2499 23991
rect -2393 23988 -2064 23990
rect -2060 23988 2499 23990
rect -2371 23942 -2366 23988
rect -2348 23942 -2343 23988
rect -2325 23976 -2317 23988
rect -2060 23985 -2054 23988
rect -2084 23978 -2054 23985
rect -2050 23982 -2044 23984
rect -2325 23956 -2320 23976
rect -2064 23974 -2054 23978
rect -2325 23948 -2317 23956
rect -2101 23951 -2071 23954
rect -2325 23942 -2320 23948
rect -2317 23942 -2309 23948
rect -2000 23946 -1992 23988
rect -1846 23987 -1806 23988
rect -1846 23978 -1798 23985
rect -1671 23976 -1663 23988
rect -1846 23974 -1806 23976
rect -1854 23960 -1680 23964
rect -1846 23951 -1798 23954
rect -2079 23945 -2043 23946
rect -2007 23945 -1991 23946
rect -2079 23944 -2071 23945
rect -2079 23942 -2029 23944
rect -2011 23942 -1991 23945
rect -1846 23943 -1806 23949
rect -1671 23948 -1663 23956
rect -1864 23942 -1796 23943
rect -1663 23942 -1655 23948
rect -1642 23942 -1637 23988
rect -1619 23942 -1614 23988
rect -1530 23942 -1526 23988
rect -1506 23942 -1502 23988
rect -1482 23942 -1478 23988
rect -1458 23942 -1454 23988
rect -1434 23942 -1430 23988
rect -1410 23942 -1406 23988
rect -1386 23942 -1382 23988
rect -1362 23942 -1358 23988
rect -1338 23942 -1334 23988
rect -1314 23942 -1310 23988
rect -1290 23942 -1286 23988
rect -1266 23942 -1262 23988
rect -1242 23942 -1238 23988
rect -1218 23942 -1214 23988
rect -1194 23942 -1190 23988
rect -1170 23942 -1166 23988
rect -1146 23942 -1142 23988
rect -1122 23942 -1118 23988
rect -1098 23942 -1094 23988
rect -1074 23942 -1070 23988
rect -1050 23942 -1046 23988
rect -1026 23942 -1022 23988
rect -1002 23942 -998 23988
rect -978 23942 -974 23988
rect -954 23942 -950 23988
rect -930 23942 -926 23988
rect -906 23942 -902 23988
rect -882 23942 -878 23988
rect -869 23957 -864 23967
rect -858 23957 -854 23988
rect -859 23943 -854 23957
rect -858 23942 -854 23943
rect -834 23942 -830 23988
rect -810 23942 -806 23988
rect -786 23942 -782 23988
rect -762 23942 -758 23988
rect -738 23942 -734 23988
rect -714 23942 -710 23988
rect -690 23942 -686 23988
rect -666 23942 -662 23988
rect -642 23942 -638 23988
rect -618 23942 -614 23988
rect -594 23942 -590 23988
rect -570 23942 -566 23988
rect -546 23942 -542 23988
rect -522 23942 -518 23988
rect -498 23942 -494 23988
rect -474 23942 -470 23988
rect -450 23942 -446 23988
rect -426 23942 -422 23988
rect -402 23942 -398 23988
rect -378 23942 -374 23988
rect -354 23942 -350 23988
rect -330 23942 -326 23988
rect -306 23942 -302 23988
rect -282 23942 -278 23988
rect -258 23942 -254 23988
rect -234 23942 -230 23988
rect -210 23942 -206 23988
rect -186 23942 -182 23988
rect -162 23942 -158 23988
rect -138 23942 -134 23988
rect -114 23942 -110 23988
rect -90 23942 -86 23988
rect -66 23942 -62 23988
rect -42 23942 -38 23988
rect -18 23942 -14 23988
rect 6 23942 10 23988
rect 30 23942 34 23988
rect 54 23942 58 23988
rect 78 23942 82 23988
rect 102 23942 106 23988
rect 126 23942 130 23988
rect 150 23942 154 23988
rect 174 23942 178 23988
rect 198 23942 202 23988
rect 222 23942 226 23988
rect 246 23942 250 23988
rect 270 23942 274 23988
rect 294 23942 298 23988
rect 318 23942 322 23988
rect 342 23942 346 23988
rect 366 23942 370 23988
rect 390 23942 394 23988
rect 414 23942 418 23988
rect 438 23942 442 23988
rect 462 23942 466 23988
rect 486 23942 490 23988
rect 510 23942 514 23988
rect 534 23942 538 23988
rect 558 23942 562 23988
rect 582 23942 586 23988
rect 606 23942 610 23988
rect 630 23942 634 23988
rect 654 23942 658 23988
rect 678 23942 682 23988
rect 702 23942 706 23988
rect 726 23942 730 23988
rect 750 23942 754 23988
rect 774 23942 778 23988
rect 798 23942 802 23988
rect 822 23942 826 23988
rect 846 23942 850 23988
rect 870 23942 874 23988
rect 894 23942 898 23988
rect 918 23942 922 23988
rect 942 23942 946 23988
rect 966 23942 970 23988
rect 990 23942 994 23988
rect 1014 23942 1018 23988
rect 1038 23942 1042 23988
rect 1062 23942 1066 23988
rect 1086 23942 1090 23988
rect 1110 23942 1114 23988
rect 1134 23942 1138 23988
rect 1158 23942 1162 23988
rect 1182 23942 1186 23988
rect 1206 23942 1210 23988
rect 1230 23942 1234 23988
rect 1254 23942 1258 23988
rect 1278 23942 1282 23988
rect 1302 23942 1306 23988
rect 1326 23942 1330 23988
rect 1350 23942 1354 23988
rect 1374 23942 1378 23988
rect 1398 23942 1402 23988
rect 1422 23942 1426 23988
rect 1446 23942 1450 23988
rect 1470 23942 1474 23988
rect 1494 23942 1498 23988
rect 1518 23942 1522 23988
rect 1542 23942 1546 23988
rect 1566 23942 1570 23988
rect 1590 23942 1594 23988
rect 1614 23942 1618 23988
rect 1638 23942 1642 23988
rect 1662 23942 1666 23988
rect 1686 23942 1690 23988
rect 1710 23942 1714 23988
rect 1734 23942 1738 23988
rect 1758 23942 1762 23988
rect 1782 23942 1786 23988
rect 1806 23942 1810 23988
rect 1830 23942 1834 23988
rect 1854 23942 1858 23988
rect 1878 23942 1882 23988
rect 1902 23942 1906 23988
rect 1926 23942 1930 23988
rect 1950 23942 1954 23988
rect 1974 23942 1978 23988
rect 1998 23942 2002 23988
rect 2022 23942 2026 23988
rect 2046 23942 2050 23988
rect 2070 23942 2074 23988
rect 2094 23942 2098 23988
rect 2118 23942 2122 23988
rect 2142 23942 2146 23988
rect 2166 23942 2170 23988
rect 2190 23942 2194 23988
rect 2214 23942 2218 23988
rect 2238 23942 2242 23988
rect 2262 23942 2266 23988
rect 2286 23942 2290 23988
rect 2310 23942 2314 23988
rect 2334 23942 2338 23988
rect 2358 23942 2362 23988
rect 2382 23942 2386 23988
rect 2406 23942 2410 23988
rect 2430 23942 2434 23988
rect 2454 23987 2458 23988
rect 2443 23942 2451 23943
rect -2393 23940 2451 23942
rect -2371 23870 -2366 23940
rect -2348 23870 -2343 23940
rect -2325 23928 -2320 23940
rect -2079 23938 -2071 23940
rect -2072 23936 -2071 23938
rect -2109 23931 -2101 23936
rect -2101 23929 -2079 23931
rect -2069 23929 -2068 23936
rect -2325 23920 -2317 23928
rect -2079 23924 -2071 23929
rect -2325 23870 -2320 23920
rect -2317 23912 -2309 23920
rect -2074 23915 -2071 23924
rect -2069 23920 -2068 23924
rect -2109 23906 -2079 23909
rect -2309 23872 -2301 23882
rect -2317 23870 -2309 23872
rect -2000 23870 -1992 23940
rect -1846 23938 -1806 23940
rect -1854 23933 -1806 23937
rect -1854 23931 -1846 23933
rect -1846 23929 -1806 23931
rect -1806 23927 -1798 23929
rect -1846 23924 -1798 23927
rect -1846 23911 -1806 23922
rect -1671 23920 -1663 23928
rect -1663 23912 -1655 23920
rect -1854 23906 -1680 23910
rect -1655 23872 -1647 23882
rect -1663 23870 -1655 23872
rect -1642 23870 -1637 23940
rect -1619 23870 -1614 23940
rect -1530 23870 -1526 23940
rect -1506 23870 -1502 23940
rect -1482 23870 -1478 23940
rect -1458 23870 -1454 23940
rect -1434 23870 -1430 23940
rect -1410 23870 -1406 23940
rect -1386 23870 -1382 23940
rect -1362 23870 -1358 23940
rect -1338 23870 -1334 23940
rect -1314 23870 -1310 23940
rect -1290 23870 -1286 23940
rect -1266 23870 -1262 23940
rect -1242 23870 -1238 23940
rect -1218 23870 -1214 23940
rect -1194 23870 -1190 23940
rect -1170 23870 -1166 23940
rect -1146 23870 -1142 23940
rect -1122 23870 -1118 23940
rect -1098 23870 -1094 23940
rect -1074 23870 -1070 23940
rect -1050 23870 -1046 23940
rect -1026 23870 -1022 23940
rect -1002 23870 -998 23940
rect -978 23870 -974 23940
rect -954 23870 -950 23940
rect -930 23870 -926 23940
rect -906 23870 -902 23940
rect -882 23870 -878 23940
rect -858 23870 -854 23940
rect -834 23891 -830 23940
rect -2393 23868 -837 23870
rect -2371 23774 -2366 23868
rect -2348 23774 -2343 23868
rect -2325 23806 -2320 23868
rect -2317 23866 -2309 23868
rect -2013 23866 -1992 23868
rect -1663 23866 -1655 23868
rect -2000 23865 -1983 23866
rect -2026 23856 -2021 23860
rect -2062 23855 -2061 23856
rect -2309 23844 -2301 23854
rect -2091 23848 -2061 23855
rect -2317 23838 -2309 23844
rect -2132 23839 -2131 23841
rect -2101 23839 -2092 23841
rect -2091 23840 -2071 23846
rect -2062 23844 -2045 23848
rect -2036 23844 -2031 23846
rect -2292 23830 -2071 23839
rect -2107 23825 -2104 23829
rect -2325 23798 -2317 23806
rect -2325 23778 -2320 23798
rect -2317 23790 -2309 23798
rect -2325 23774 -2317 23778
rect -2000 23774 -1992 23865
rect -1980 23848 -1932 23855
rect -1655 23844 -1647 23854
rect -1846 23830 -1680 23839
rect -1663 23838 -1655 23844
rect -1671 23798 -1663 23806
rect -1663 23790 -1655 23798
rect -1671 23774 -1663 23778
rect -1642 23774 -1637 23868
rect -1619 23774 -1614 23868
rect -1530 23774 -1526 23868
rect -1506 23774 -1502 23868
rect -1482 23774 -1478 23868
rect -1458 23774 -1454 23868
rect -1434 23774 -1430 23868
rect -1410 23774 -1406 23868
rect -1386 23774 -1382 23868
rect -1362 23774 -1358 23868
rect -1338 23774 -1334 23868
rect -1314 23774 -1310 23868
rect -1290 23774 -1286 23868
rect -1266 23774 -1262 23868
rect -1242 23774 -1238 23868
rect -1218 23774 -1214 23868
rect -1194 23774 -1190 23868
rect -1170 23774 -1166 23868
rect -1146 23774 -1142 23868
rect -1122 23774 -1118 23868
rect -1098 23774 -1094 23868
rect -1074 23774 -1070 23868
rect -1050 23774 -1046 23868
rect -1026 23774 -1022 23868
rect -1002 23774 -998 23868
rect -978 23774 -974 23868
rect -954 23774 -950 23868
rect -930 23774 -926 23868
rect -906 23774 -902 23868
rect -882 23774 -878 23868
rect -858 23774 -854 23868
rect -851 23867 -837 23868
rect -834 23867 -827 23891
rect -834 23774 -830 23867
rect -810 23774 -806 23940
rect -786 23774 -782 23940
rect -762 23774 -758 23940
rect -738 23774 -734 23940
rect -714 23774 -710 23940
rect -690 23774 -686 23940
rect -666 23774 -662 23940
rect -642 23774 -638 23940
rect -618 23774 -614 23940
rect -594 23774 -590 23940
rect -570 23774 -566 23940
rect -546 23774 -542 23940
rect -522 23774 -518 23940
rect -498 23774 -494 23940
rect -474 23774 -470 23940
rect -450 23774 -446 23940
rect -426 23774 -422 23940
rect -413 23813 -408 23823
rect -402 23813 -398 23940
rect -403 23799 -398 23813
rect -402 23774 -398 23799
rect -378 23774 -374 23940
rect -354 23774 -350 23940
rect -330 23774 -326 23940
rect -306 23774 -302 23940
rect -282 23895 -278 23940
rect -293 23894 -259 23895
rect -258 23894 -254 23940
rect -234 23894 -230 23940
rect -210 23894 -206 23940
rect -186 23894 -182 23940
rect -162 23894 -158 23940
rect -138 23894 -134 23940
rect -114 23894 -110 23940
rect -90 23894 -86 23940
rect -66 23894 -62 23940
rect -42 23894 -38 23940
rect -18 23894 -14 23940
rect 6 23894 10 23940
rect 30 23894 34 23940
rect 54 23894 58 23940
rect 78 23894 82 23940
rect 102 23894 106 23940
rect 126 23894 130 23940
rect 150 23894 154 23940
rect 174 23894 178 23940
rect 198 23894 202 23940
rect 222 23894 226 23940
rect 246 23894 250 23940
rect 270 23894 274 23940
rect 294 23894 298 23940
rect 318 23894 322 23940
rect 342 23894 346 23940
rect 366 23894 370 23940
rect 390 23894 394 23940
rect 414 23894 418 23940
rect 438 23894 442 23940
rect 462 23894 466 23940
rect 486 23894 490 23940
rect 510 23894 514 23940
rect 534 23894 538 23940
rect 558 23894 562 23940
rect 582 23894 586 23940
rect 606 23894 610 23940
rect 630 23894 634 23940
rect 654 23894 658 23940
rect 678 23894 682 23940
rect 702 23894 706 23940
rect 726 23894 730 23940
rect 750 23894 754 23940
rect 774 23894 778 23940
rect 798 23894 802 23940
rect 822 23894 826 23940
rect 846 23894 850 23940
rect 870 23894 874 23940
rect 894 23894 898 23940
rect 918 23894 922 23940
rect 942 23894 946 23940
rect 966 23894 970 23940
rect 990 23894 994 23940
rect 1014 23894 1018 23940
rect 1038 23894 1042 23940
rect 1062 23894 1066 23940
rect 1086 23894 1090 23940
rect 1110 23894 1114 23940
rect 1134 23894 1138 23940
rect 1158 23894 1162 23940
rect 1182 23894 1186 23940
rect 1206 23894 1210 23940
rect 1230 23894 1234 23940
rect 1254 23894 1258 23940
rect 1278 23894 1282 23940
rect 1302 23894 1306 23940
rect 1326 23894 1330 23940
rect 1350 23894 1354 23940
rect 1374 23894 1378 23940
rect 1398 23894 1402 23940
rect 1422 23939 1426 23940
rect 1422 23915 1429 23939
rect 1422 23894 1426 23915
rect 1446 23894 1450 23940
rect 1470 23894 1474 23940
rect 1494 23894 1498 23940
rect 1518 23894 1522 23940
rect 1542 23894 1546 23940
rect 1566 23894 1570 23940
rect 1590 23894 1594 23940
rect 1614 23894 1618 23940
rect 1638 23894 1642 23940
rect 1662 23894 1666 23940
rect 1686 23894 1690 23940
rect 1710 23894 1714 23940
rect 1734 23894 1738 23940
rect 1758 23894 1762 23940
rect 1782 23894 1786 23940
rect 1806 23894 1810 23940
rect 1830 23894 1834 23940
rect 1854 23894 1858 23940
rect 1878 23894 1882 23940
rect 1902 23894 1906 23940
rect 1926 23894 1930 23940
rect 1950 23894 1954 23940
rect 1974 23894 1978 23940
rect 1998 23894 2002 23940
rect 2022 23894 2026 23940
rect 2046 23894 2050 23940
rect 2070 23894 2074 23940
rect 2094 23894 2098 23940
rect 2118 23894 2122 23940
rect 2142 23894 2146 23940
rect 2166 23894 2170 23940
rect 2190 23894 2194 23940
rect 2214 23894 2218 23940
rect 2238 23894 2242 23940
rect 2262 23894 2266 23940
rect 2286 23894 2290 23940
rect 2310 23894 2314 23940
rect 2334 23894 2338 23940
rect 2358 23894 2362 23940
rect 2382 23894 2386 23940
rect 2406 23894 2410 23940
rect 2430 23894 2434 23940
rect 2437 23939 2451 23940
rect 2454 23939 2461 23987
rect 2467 23981 2472 23988
rect 2478 23981 2482 23988
rect 2485 23987 2499 23988
rect 2477 23967 2482 23981
rect 2491 23977 2499 23981
rect 2485 23967 2491 23977
rect 2443 23933 2448 23939
rect 2454 23933 2458 23939
rect 2453 23919 2458 23933
rect 2443 23894 2477 23895
rect -293 23892 2477 23894
rect -293 23885 -288 23892
rect -282 23885 -278 23892
rect -283 23871 -278 23885
rect -293 23861 -288 23871
rect -283 23847 -278 23861
rect -282 23774 -278 23847
rect -258 23819 -254 23892
rect -2393 23772 -261 23774
rect -2371 23726 -2366 23772
rect -2348 23726 -2343 23772
rect -2325 23764 -2317 23772
rect -2018 23771 -2004 23772
rect -2000 23771 -1992 23772
rect -2072 23770 -1928 23771
rect -2072 23764 -2053 23770
rect -2325 23748 -2320 23764
rect -2317 23762 -2309 23764
rect -2309 23750 -2301 23762
rect -2092 23755 -2062 23760
rect -2317 23748 -2309 23750
rect -2325 23736 -2317 23748
rect -2098 23742 -2096 23753
rect -2092 23742 -2084 23755
rect -2000 23754 -1992 23770
rect -1972 23764 -1928 23770
rect -1924 23764 -1918 23772
rect -1671 23764 -1663 23772
rect -1663 23762 -1655 23764
rect -2083 23744 -2062 23753
rect -2027 23752 -1992 23754
rect -2018 23744 -2002 23752
rect -2000 23744 -1992 23752
rect -2100 23737 -2096 23742
rect -2083 23737 -2053 23742
rect -2003 23740 -1990 23744
rect -1972 23742 -1964 23751
rect -1928 23750 -1924 23753
rect -1655 23750 -1647 23762
rect -1663 23748 -1655 23750
rect -2325 23726 -2320 23736
rect -2317 23734 -2309 23736
rect -2309 23726 -2301 23734
rect -2004 23730 -2003 23740
rect -2062 23726 -2012 23728
rect -2000 23726 -1992 23740
rect -1972 23737 -1924 23742
rect -1864 23737 -1796 23743
rect -1671 23736 -1663 23748
rect -1663 23734 -1655 23736
rect -1864 23726 -1796 23727
rect -1655 23726 -1647 23734
rect -1642 23726 -1637 23772
rect -1619 23726 -1614 23772
rect -1530 23726 -1526 23772
rect -1506 23726 -1502 23772
rect -1482 23726 -1478 23772
rect -1458 23726 -1454 23772
rect -1434 23726 -1430 23772
rect -1410 23726 -1406 23772
rect -1386 23726 -1382 23772
rect -1362 23726 -1358 23772
rect -1338 23726 -1334 23772
rect -1314 23726 -1310 23772
rect -1290 23726 -1286 23772
rect -1266 23726 -1262 23772
rect -1242 23726 -1238 23772
rect -1218 23726 -1214 23772
rect -1194 23726 -1190 23772
rect -1170 23726 -1166 23772
rect -1146 23726 -1142 23772
rect -1122 23726 -1118 23772
rect -1098 23726 -1094 23772
rect -1074 23726 -1070 23772
rect -1050 23726 -1046 23772
rect -1026 23726 -1022 23772
rect -1002 23726 -998 23772
rect -978 23726 -974 23772
rect -954 23726 -950 23772
rect -930 23726 -926 23772
rect -906 23726 -902 23772
rect -882 23726 -878 23772
rect -858 23726 -854 23772
rect -834 23726 -830 23772
rect -810 23726 -806 23772
rect -786 23726 -782 23772
rect -762 23726 -758 23772
rect -738 23726 -734 23772
rect -714 23726 -710 23772
rect -690 23726 -686 23772
rect -666 23726 -662 23772
rect -642 23726 -638 23772
rect -618 23726 -614 23772
rect -594 23726 -590 23772
rect -570 23726 -566 23772
rect -546 23726 -542 23772
rect -522 23726 -518 23772
rect -498 23726 -494 23772
rect -474 23726 -470 23772
rect -450 23726 -446 23772
rect -426 23726 -422 23772
rect -413 23741 -408 23751
rect -402 23741 -398 23772
rect -378 23747 -374 23772
rect -403 23727 -398 23741
rect -389 23737 -381 23741
rect -395 23727 -389 23737
rect -402 23726 -398 23727
rect -2393 23724 -381 23726
rect -2371 23678 -2366 23724
rect -2348 23678 -2343 23724
rect -2325 23720 -2320 23724
rect -2309 23722 -2301 23724
rect -2317 23720 -2309 23722
rect -2325 23708 -2317 23720
rect -2325 23678 -2320 23708
rect -2317 23706 -2309 23708
rect -2092 23694 -2062 23696
rect -2094 23690 -2062 23694
rect -2000 23678 -1992 23724
rect -1655 23722 -1647 23724
rect -1663 23720 -1655 23722
rect -1671 23708 -1663 23720
rect -1663 23706 -1655 23708
rect -1854 23694 -1806 23696
rect -1854 23690 -1680 23694
rect -1642 23678 -1637 23724
rect -1619 23678 -1614 23724
rect -1530 23678 -1526 23724
rect -1506 23678 -1502 23724
rect -1482 23678 -1478 23724
rect -1458 23678 -1454 23724
rect -1434 23678 -1430 23724
rect -1410 23678 -1406 23724
rect -1386 23678 -1382 23724
rect -1362 23678 -1358 23724
rect -1338 23678 -1334 23724
rect -1314 23678 -1310 23724
rect -1290 23678 -1286 23724
rect -1266 23678 -1262 23724
rect -1242 23678 -1238 23724
rect -1218 23678 -1214 23724
rect -1194 23678 -1190 23724
rect -1170 23678 -1166 23724
rect -1146 23678 -1142 23724
rect -1122 23678 -1118 23724
rect -1098 23678 -1094 23724
rect -1074 23678 -1070 23724
rect -1050 23678 -1046 23724
rect -1026 23678 -1022 23724
rect -1002 23678 -998 23724
rect -978 23678 -974 23724
rect -954 23678 -950 23724
rect -930 23678 -926 23724
rect -906 23678 -902 23724
rect -882 23678 -878 23724
rect -858 23678 -854 23724
rect -834 23678 -830 23724
rect -810 23678 -806 23724
rect -786 23678 -782 23724
rect -762 23678 -758 23724
rect -738 23678 -734 23724
rect -714 23678 -710 23724
rect -690 23678 -686 23724
rect -666 23678 -662 23724
rect -642 23678 -638 23724
rect -618 23678 -614 23724
rect -594 23678 -590 23724
rect -570 23678 -566 23724
rect -546 23678 -542 23724
rect -522 23678 -518 23724
rect -498 23678 -494 23724
rect -474 23678 -470 23724
rect -450 23678 -446 23724
rect -426 23678 -422 23724
rect -402 23678 -398 23724
rect -395 23723 -381 23724
rect -378 23723 -371 23747
rect -378 23678 -374 23723
rect -354 23678 -350 23772
rect -330 23678 -326 23772
rect -306 23678 -302 23772
rect -282 23678 -278 23772
rect -275 23771 -261 23772
rect -258 23771 -251 23819
rect -258 23678 -254 23771
rect -234 23678 -230 23892
rect -210 23678 -206 23892
rect -186 23678 -182 23892
rect -162 23678 -158 23892
rect -138 23678 -134 23892
rect -114 23678 -110 23892
rect -90 23678 -86 23892
rect -66 23678 -62 23892
rect -42 23678 -38 23892
rect -18 23678 -14 23892
rect 6 23678 10 23892
rect 30 23678 34 23892
rect 54 23678 58 23892
rect 78 23678 82 23892
rect 102 23678 106 23892
rect 126 23678 130 23892
rect 150 23678 154 23892
rect 174 23678 178 23892
rect 198 23678 202 23892
rect 222 23678 226 23892
rect 246 23678 250 23892
rect 270 23678 274 23892
rect 294 23678 298 23892
rect 318 23678 322 23892
rect 342 23678 346 23892
rect 366 23678 370 23892
rect 390 23678 394 23892
rect 414 23678 418 23892
rect 438 23678 442 23892
rect 462 23678 466 23892
rect 486 23678 490 23892
rect 510 23678 514 23892
rect 534 23678 538 23892
rect 558 23678 562 23892
rect 582 23678 586 23892
rect 606 23678 610 23892
rect 630 23678 634 23892
rect 654 23678 658 23892
rect 678 23678 682 23892
rect 702 23678 706 23892
rect 726 23678 730 23892
rect 750 23678 754 23892
rect 774 23678 778 23892
rect 798 23678 802 23892
rect 822 23678 826 23892
rect 846 23678 850 23892
rect 870 23678 874 23892
rect 894 23678 898 23892
rect 918 23678 922 23892
rect 942 23678 946 23892
rect 966 23678 970 23892
rect 990 23678 994 23892
rect 1014 23678 1018 23892
rect 1038 23678 1042 23892
rect 1062 23678 1066 23892
rect 1086 23678 1090 23892
rect 1110 23678 1114 23892
rect 1134 23678 1138 23892
rect 1158 23678 1162 23892
rect 1182 23678 1186 23892
rect 1206 23678 1210 23892
rect 1230 23678 1234 23892
rect 1254 23678 1258 23892
rect 1278 23678 1282 23892
rect 1302 23678 1306 23892
rect 1326 23678 1330 23892
rect 1350 23678 1354 23892
rect 1374 23678 1378 23892
rect 1398 23678 1402 23892
rect 1422 23678 1426 23892
rect 1435 23693 1440 23703
rect 1446 23693 1450 23892
rect 1445 23679 1450 23693
rect 1435 23678 1469 23679
rect -2393 23676 1469 23678
rect -2371 23654 -2366 23676
rect -2348 23654 -2343 23676
rect -2325 23654 -2320 23676
rect -2072 23674 -2036 23675
rect -2072 23668 -2054 23674
rect -2309 23660 -2301 23668
rect -2317 23654 -2309 23660
rect -2092 23659 -2062 23664
rect -2000 23655 -1992 23676
rect -1938 23675 -1906 23676
rect -1920 23674 -1906 23675
rect -1806 23668 -1680 23674
rect -1854 23659 -1806 23664
rect -1655 23660 -1647 23668
rect -1982 23655 -1966 23656
rect -2000 23654 -1966 23655
rect -1846 23654 -1806 23657
rect -1663 23654 -1655 23660
rect -1642 23654 -1637 23676
rect -1619 23654 -1614 23676
rect -1530 23654 -1526 23676
rect -1506 23654 -1502 23676
rect -1482 23654 -1478 23676
rect -1458 23654 -1454 23676
rect -1434 23654 -1430 23676
rect -1410 23654 -1406 23676
rect -1386 23654 -1382 23676
rect -1362 23654 -1358 23676
rect -1338 23654 -1334 23676
rect -1314 23654 -1310 23676
rect -1290 23654 -1286 23676
rect -1266 23654 -1262 23676
rect -1242 23654 -1238 23676
rect -1218 23654 -1214 23676
rect -1194 23654 -1190 23676
rect -1170 23654 -1166 23676
rect -1146 23654 -1142 23676
rect -1122 23654 -1118 23676
rect -1098 23654 -1094 23676
rect -1074 23654 -1070 23676
rect -1050 23654 -1046 23676
rect -1026 23654 -1022 23676
rect -1002 23654 -998 23676
rect -978 23654 -974 23676
rect -954 23654 -950 23676
rect -930 23654 -926 23676
rect -906 23654 -902 23676
rect -882 23654 -878 23676
rect -858 23654 -854 23676
rect -834 23654 -830 23676
rect -810 23654 -806 23676
rect -786 23654 -782 23676
rect -762 23654 -758 23676
rect -738 23654 -734 23676
rect -714 23654 -710 23676
rect -690 23654 -686 23676
rect -666 23654 -662 23676
rect -642 23654 -638 23676
rect -618 23654 -614 23676
rect -594 23654 -590 23676
rect -570 23654 -566 23676
rect -546 23654 -542 23676
rect -522 23654 -518 23676
rect -498 23654 -494 23676
rect -474 23654 -470 23676
rect -450 23654 -446 23676
rect -426 23654 -422 23676
rect -402 23654 -398 23676
rect -378 23675 -374 23676
rect -2393 23652 -381 23654
rect -2371 23630 -2366 23652
rect -2348 23630 -2343 23652
rect -2325 23630 -2320 23652
rect -2000 23650 -1966 23652
rect -2309 23632 -2301 23640
rect -2062 23639 -2054 23646
rect -2092 23632 -2084 23639
rect -2062 23632 -2026 23634
rect -2317 23630 -2309 23632
rect -2062 23630 -2012 23632
rect -2000 23630 -1992 23650
rect -1982 23649 -1966 23650
rect -1846 23648 -1806 23652
rect -1846 23641 -1798 23646
rect -1806 23639 -1798 23641
rect -1854 23637 -1846 23639
rect -1854 23632 -1806 23637
rect -1655 23632 -1647 23640
rect -1864 23630 -1796 23631
rect -1663 23630 -1655 23632
rect -1642 23630 -1637 23652
rect -1619 23630 -1614 23652
rect -1530 23630 -1526 23652
rect -1506 23630 -1502 23652
rect -1482 23630 -1478 23652
rect -1458 23630 -1454 23652
rect -1434 23630 -1430 23652
rect -1410 23630 -1406 23652
rect -1386 23630 -1382 23652
rect -1362 23630 -1358 23652
rect -1338 23630 -1334 23652
rect -1314 23630 -1310 23652
rect -1290 23630 -1286 23652
rect -1266 23630 -1262 23652
rect -1242 23630 -1238 23652
rect -1218 23630 -1214 23652
rect -1194 23630 -1190 23652
rect -1170 23630 -1166 23652
rect -1146 23630 -1142 23652
rect -1122 23630 -1118 23652
rect -1098 23630 -1094 23652
rect -1074 23630 -1070 23652
rect -1050 23630 -1046 23652
rect -1026 23630 -1022 23652
rect -1002 23631 -998 23652
rect -1013 23630 -979 23631
rect -2393 23628 -979 23630
rect -2371 23582 -2366 23628
rect -2348 23582 -2343 23628
rect -2325 23582 -2320 23628
rect -2317 23624 -2309 23628
rect -2062 23624 -2054 23628
rect -2154 23620 -2138 23622
rect -2057 23620 -2054 23624
rect -2292 23614 -2054 23620
rect -2052 23614 -2044 23624
rect -2092 23598 -2062 23600
rect -2094 23594 -2062 23598
rect -2000 23582 -1992 23628
rect -1846 23621 -1806 23628
rect -1663 23624 -1655 23628
rect -1846 23614 -1680 23620
rect -1854 23598 -1806 23600
rect -1854 23594 -1680 23598
rect -1979 23582 -1945 23584
rect -1642 23582 -1637 23628
rect -1619 23582 -1614 23628
rect -1530 23582 -1526 23628
rect -1506 23582 -1502 23628
rect -1482 23582 -1478 23628
rect -1458 23582 -1454 23628
rect -1434 23582 -1430 23628
rect -1410 23582 -1406 23628
rect -1386 23582 -1382 23628
rect -1362 23582 -1358 23628
rect -1338 23582 -1334 23628
rect -1314 23582 -1310 23628
rect -1290 23582 -1286 23628
rect -1266 23582 -1262 23628
rect -1242 23582 -1238 23628
rect -1218 23582 -1214 23628
rect -1194 23582 -1190 23628
rect -1170 23582 -1166 23628
rect -1146 23582 -1142 23628
rect -1122 23582 -1118 23628
rect -1098 23582 -1094 23628
rect -1074 23582 -1070 23628
rect -1050 23582 -1046 23628
rect -1026 23582 -1022 23628
rect -1013 23621 -1008 23628
rect -1002 23621 -998 23628
rect -1003 23607 -998 23621
rect -1002 23582 -998 23607
rect -978 23582 -974 23652
rect -954 23582 -950 23652
rect -930 23582 -926 23652
rect -906 23582 -902 23652
rect -882 23582 -878 23652
rect -858 23582 -854 23652
rect -834 23582 -830 23652
rect -810 23582 -806 23652
rect -786 23582 -782 23652
rect -762 23582 -758 23652
rect -738 23582 -734 23652
rect -714 23582 -710 23652
rect -690 23582 -686 23652
rect -666 23582 -662 23652
rect -642 23582 -638 23652
rect -618 23582 -614 23652
rect -594 23582 -590 23652
rect -570 23582 -566 23652
rect -546 23582 -542 23652
rect -522 23582 -518 23652
rect -498 23582 -494 23652
rect -474 23582 -470 23652
rect -450 23582 -446 23652
rect -426 23582 -422 23652
rect -402 23582 -398 23652
rect -395 23651 -381 23652
rect -378 23651 -371 23675
rect -378 23582 -374 23651
rect -354 23582 -350 23676
rect -330 23582 -326 23676
rect -306 23582 -302 23676
rect -282 23582 -278 23676
rect -258 23582 -254 23676
rect -245 23597 -240 23607
rect -234 23597 -230 23676
rect -235 23583 -230 23597
rect -245 23582 -211 23583
rect -2393 23580 -211 23582
rect -2371 23534 -2366 23580
rect -2348 23534 -2343 23580
rect -2325 23534 -2320 23580
rect -2080 23579 -1906 23580
rect -2080 23578 -2036 23579
rect -2080 23572 -2054 23578
rect -2309 23564 -2301 23570
rect -2317 23554 -2309 23564
rect -2070 23563 -2040 23570
rect -2054 23555 -2040 23558
rect -2000 23553 -1992 23579
rect -1920 23578 -1906 23579
rect -1850 23572 -1846 23580
rect -1840 23572 -1792 23580
rect -1969 23560 -1966 23569
rect -1850 23565 -1802 23570
rect -1906 23563 -1802 23565
rect -1655 23564 -1647 23570
rect -1906 23562 -1850 23563
rect -1846 23555 -1802 23561
rect -1663 23554 -1655 23564
rect -1860 23553 -1798 23554
rect -2078 23546 -2070 23553
rect -2309 23536 -2301 23542
rect -2317 23534 -2309 23536
rect -2154 23534 -2145 23544
rect -2044 23543 -2040 23548
rect -2028 23546 -1945 23553
rect -1929 23546 -1794 23553
rect -2070 23536 -2040 23543
rect -2044 23534 -2028 23536
rect -2000 23534 -1992 23546
rect -1860 23545 -1798 23546
rect -1850 23536 -1802 23543
rect -1655 23536 -1647 23542
rect -1978 23534 -1942 23535
rect -1663 23534 -1655 23536
rect -1642 23534 -1637 23580
rect -1619 23534 -1614 23580
rect -1589 23534 -1555 23535
rect -2393 23532 -1555 23534
rect -2371 23438 -2366 23532
rect -2348 23438 -2343 23532
rect -2325 23494 -2320 23532
rect -2317 23526 -2309 23532
rect -2145 23528 -2138 23532
rect -2070 23528 -2054 23532
rect -2078 23519 -2054 23526
rect -2062 23494 -2032 23495
rect -2000 23494 -1992 23532
rect -1846 23528 -1802 23532
rect -1846 23518 -1792 23527
rect -1663 23526 -1655 23532
rect -1942 23496 -1937 23508
rect -1850 23505 -1822 23506
rect -1850 23501 -1802 23505
rect -2325 23486 -2317 23494
rect -2062 23492 -1961 23494
rect -2325 23466 -2320 23486
rect -2317 23478 -2309 23486
rect -2062 23479 -2040 23490
rect -2032 23485 -1961 23492
rect -1947 23486 -1942 23494
rect -1842 23492 -1794 23495
rect -2070 23474 -2022 23478
rect -2325 23452 -2317 23466
rect -2072 23458 -2032 23459
rect -2102 23452 -2032 23458
rect -2325 23438 -2320 23452
rect -2317 23450 -2309 23452
rect -2309 23438 -2301 23450
rect -2070 23443 -2062 23448
rect -2000 23438 -1992 23485
rect -1942 23484 -1937 23486
rect -1932 23476 -1927 23484
rect -1912 23481 -1896 23487
rect -1842 23479 -1802 23490
rect -1671 23486 -1663 23494
rect -1663 23478 -1655 23486
rect -1850 23474 -1680 23478
rect -1924 23460 -1921 23462
rect -1806 23452 -1680 23458
rect -1671 23452 -1663 23466
rect -1663 23450 -1655 23452
rect -1854 23443 -1806 23448
rect -1974 23438 -1964 23439
rect -1960 23438 -1944 23440
rect -1842 23438 -1806 23441
rect -1655 23438 -1647 23450
rect -1642 23438 -1637 23532
rect -1619 23438 -1614 23532
rect -1554 23446 -1547 23459
rect -2393 23436 -1557 23438
rect -2371 23414 -2366 23436
rect -2348 23414 -2343 23436
rect -2325 23424 -2317 23436
rect -2325 23414 -2320 23424
rect -2317 23422 -2309 23424
rect -2062 23423 -2032 23430
rect -2309 23414 -2301 23422
rect -2070 23416 -2062 23423
rect -2000 23418 -1992 23436
rect -1974 23434 -1944 23436
rect -1960 23433 -1944 23434
rect -1842 23432 -1806 23436
rect -1842 23425 -1798 23430
rect -1806 23423 -1798 23425
rect -1671 23424 -1663 23436
rect -1854 23421 -1842 23423
rect -1663 23422 -1655 23424
rect -2062 23414 -2036 23416
rect -2393 23412 -2036 23414
rect -2032 23414 -2012 23416
rect -2004 23414 -1974 23418
rect -1854 23416 -1806 23421
rect -1864 23414 -1796 23415
rect -1655 23414 -1647 23422
rect -1642 23414 -1637 23436
rect -1619 23414 -1614 23436
rect -1571 23435 -1557 23436
rect -1554 23435 -1547 23436
rect -1530 23414 -1526 23580
rect -1517 23501 -1512 23511
rect -1506 23501 -1502 23580
rect -1507 23487 -1502 23501
rect -1506 23414 -1502 23487
rect -1482 23435 -1478 23580
rect -2032 23412 -1485 23414
rect -2371 23366 -2366 23412
rect -2348 23366 -2343 23412
rect -2325 23408 -2320 23412
rect -2309 23410 -2301 23412
rect -2317 23408 -2309 23410
rect -2325 23396 -2317 23408
rect -2052 23406 -2036 23408
rect -2052 23404 -2032 23406
rect -2062 23398 -2032 23404
rect -2325 23366 -2320 23396
rect -2317 23394 -2309 23396
rect -2092 23382 -2062 23384
rect -2094 23378 -2062 23382
rect -2000 23366 -1992 23412
rect -1904 23405 -1874 23412
rect -1842 23405 -1806 23412
rect -1655 23410 -1647 23412
rect -1663 23408 -1655 23410
rect -1842 23398 -1680 23404
rect -1671 23396 -1663 23408
rect -1663 23394 -1655 23396
rect -1854 23382 -1806 23384
rect -1854 23378 -1680 23382
rect -1642 23366 -1637 23412
rect -1619 23366 -1614 23412
rect -1530 23366 -1526 23412
rect -1506 23366 -1502 23412
rect -1499 23411 -1485 23412
rect -1482 23411 -1475 23435
rect -1482 23366 -1478 23411
rect -1469 23381 -1464 23391
rect -1458 23381 -1454 23580
rect -1459 23367 -1454 23381
rect -1469 23366 -1435 23367
rect -2393 23364 -1435 23366
rect -2371 23342 -2366 23364
rect -2348 23342 -2343 23364
rect -2325 23342 -2320 23364
rect -2072 23362 -2036 23363
rect -2072 23356 -2054 23362
rect -2309 23348 -2301 23356
rect -2317 23342 -2309 23348
rect -2092 23347 -2062 23352
rect -2000 23343 -1992 23364
rect -1938 23363 -1906 23364
rect -1920 23362 -1906 23363
rect -1806 23356 -1680 23362
rect -1854 23347 -1806 23352
rect -1655 23348 -1647 23356
rect -1982 23343 -1966 23344
rect -2000 23342 -1966 23343
rect -1846 23342 -1806 23345
rect -1663 23342 -1655 23348
rect -1642 23342 -1637 23364
rect -1619 23342 -1614 23364
rect -1530 23342 -1526 23364
rect -1506 23342 -1502 23364
rect -1482 23342 -1478 23364
rect -1469 23357 -1464 23364
rect -1459 23343 -1454 23357
rect -1458 23342 -1454 23343
rect -1434 23342 -1430 23580
rect -1410 23342 -1406 23580
rect -1386 23342 -1382 23580
rect -1362 23342 -1358 23580
rect -1338 23342 -1334 23580
rect -1314 23342 -1310 23580
rect -1290 23342 -1286 23580
rect -1266 23342 -1262 23580
rect -1242 23342 -1238 23580
rect -1218 23342 -1214 23580
rect -1194 23342 -1190 23580
rect -1170 23342 -1166 23580
rect -1146 23342 -1142 23580
rect -1122 23342 -1118 23580
rect -1098 23342 -1094 23580
rect -1074 23342 -1070 23580
rect -1050 23342 -1046 23580
rect -1026 23342 -1022 23580
rect -1002 23342 -998 23580
rect -978 23555 -974 23580
rect -978 23531 -971 23555
rect -978 23342 -974 23531
rect -954 23342 -950 23580
rect -930 23342 -926 23580
rect -906 23342 -902 23580
rect -882 23342 -878 23580
rect -858 23342 -854 23580
rect -834 23342 -830 23580
rect -810 23342 -806 23580
rect -786 23342 -782 23580
rect -762 23342 -758 23580
rect -738 23342 -734 23580
rect -714 23342 -710 23580
rect -690 23342 -686 23580
rect -666 23342 -662 23580
rect -642 23342 -638 23580
rect -618 23342 -614 23580
rect -594 23342 -590 23580
rect -570 23342 -566 23580
rect -546 23342 -542 23580
rect -522 23342 -518 23580
rect -498 23342 -494 23580
rect -474 23342 -470 23580
rect -450 23342 -446 23580
rect -426 23342 -422 23580
rect -413 23429 -408 23439
rect -402 23429 -398 23580
rect -403 23415 -398 23429
rect -402 23342 -398 23415
rect -378 23363 -374 23580
rect -2393 23340 -381 23342
rect -2371 23318 -2366 23340
rect -2348 23318 -2343 23340
rect -2325 23318 -2320 23340
rect -2000 23338 -1966 23340
rect -2309 23320 -2301 23328
rect -2062 23327 -2054 23334
rect -2092 23320 -2084 23327
rect -2062 23320 -2026 23322
rect -2317 23318 -2309 23320
rect -2062 23318 -2012 23320
rect -2000 23318 -1992 23338
rect -1982 23337 -1966 23338
rect -1846 23336 -1806 23340
rect -1846 23329 -1798 23334
rect -1806 23327 -1798 23329
rect -1854 23325 -1846 23327
rect -1854 23320 -1806 23325
rect -1655 23320 -1647 23328
rect -1864 23318 -1796 23319
rect -1663 23318 -1655 23320
rect -1642 23318 -1637 23340
rect -1619 23318 -1614 23340
rect -1530 23318 -1526 23340
rect -1506 23318 -1502 23340
rect -1482 23318 -1478 23340
rect -1458 23318 -1454 23340
rect -1434 23318 -1430 23340
rect -1410 23318 -1406 23340
rect -1386 23318 -1382 23340
rect -1362 23318 -1358 23340
rect -1338 23318 -1334 23340
rect -1314 23318 -1310 23340
rect -1290 23318 -1286 23340
rect -1266 23318 -1262 23340
rect -1242 23318 -1238 23340
rect -1218 23318 -1214 23340
rect -1194 23318 -1190 23340
rect -1170 23318 -1166 23340
rect -1146 23318 -1142 23340
rect -1122 23318 -1118 23340
rect -1098 23318 -1094 23340
rect -1074 23318 -1070 23340
rect -1050 23318 -1046 23340
rect -1026 23318 -1022 23340
rect -1002 23318 -998 23340
rect -978 23318 -974 23340
rect -954 23318 -950 23340
rect -930 23318 -926 23340
rect -906 23318 -902 23340
rect -882 23318 -878 23340
rect -858 23318 -854 23340
rect -834 23318 -830 23340
rect -810 23318 -806 23340
rect -786 23318 -782 23340
rect -762 23318 -758 23340
rect -738 23318 -734 23340
rect -714 23318 -710 23340
rect -690 23318 -686 23340
rect -666 23318 -662 23340
rect -642 23318 -638 23340
rect -618 23318 -614 23340
rect -594 23318 -590 23340
rect -570 23318 -566 23340
rect -546 23318 -542 23340
rect -522 23318 -518 23340
rect -498 23318 -494 23340
rect -474 23318 -470 23340
rect -450 23318 -446 23340
rect -426 23318 -422 23340
rect -402 23318 -398 23340
rect -395 23339 -381 23340
rect -378 23339 -371 23363
rect -378 23318 -374 23339
rect -354 23318 -350 23580
rect -330 23318 -326 23580
rect -306 23318 -302 23580
rect -282 23318 -278 23580
rect -258 23318 -254 23580
rect -245 23573 -240 23580
rect -235 23559 -230 23573
rect -234 23318 -230 23559
rect -210 23531 -206 23676
rect -210 23483 -203 23531
rect -210 23318 -206 23483
rect -186 23318 -182 23676
rect -162 23318 -158 23676
rect -138 23318 -134 23676
rect -114 23318 -110 23676
rect -90 23318 -86 23676
rect -66 23318 -62 23676
rect -42 23318 -38 23676
rect -18 23318 -14 23676
rect 6 23318 10 23676
rect 30 23318 34 23676
rect 54 23318 58 23676
rect 78 23318 82 23676
rect 102 23318 106 23676
rect 126 23318 130 23676
rect 150 23318 154 23676
rect 174 23318 178 23676
rect 198 23318 202 23676
rect 222 23318 226 23676
rect 246 23318 250 23676
rect 270 23318 274 23676
rect 294 23318 298 23676
rect 318 23318 322 23676
rect 342 23318 346 23676
rect 366 23318 370 23676
rect 390 23318 394 23676
rect 414 23318 418 23676
rect 438 23318 442 23676
rect 462 23318 466 23676
rect 486 23318 490 23676
rect 499 23645 504 23655
rect 510 23645 514 23676
rect 509 23631 514 23645
rect 510 23318 514 23631
rect 534 23579 538 23676
rect 534 23555 541 23579
rect 534 23318 538 23555
rect 558 23318 562 23676
rect 582 23318 586 23676
rect 606 23318 610 23676
rect 630 23318 634 23676
rect 654 23318 658 23676
rect 678 23318 682 23676
rect 702 23318 706 23676
rect 726 23318 730 23676
rect 750 23318 754 23676
rect 774 23318 778 23676
rect 798 23318 802 23676
rect 822 23318 826 23676
rect 846 23318 850 23676
rect 870 23318 874 23676
rect 894 23318 898 23676
rect 918 23318 922 23676
rect 942 23318 946 23676
rect 966 23318 970 23676
rect 990 23318 994 23676
rect 1014 23318 1018 23676
rect 1038 23318 1042 23676
rect 1062 23318 1066 23676
rect 1086 23318 1090 23676
rect 1110 23318 1114 23676
rect 1134 23318 1138 23676
rect 1158 23318 1162 23676
rect 1182 23318 1186 23676
rect 1206 23318 1210 23676
rect 1230 23318 1234 23676
rect 1254 23318 1258 23676
rect 1278 23318 1282 23676
rect 1302 23318 1306 23676
rect 1326 23318 1330 23676
rect 1350 23318 1354 23676
rect 1374 23318 1378 23676
rect 1398 23318 1402 23676
rect 1422 23318 1426 23676
rect 1435 23669 1440 23676
rect 1445 23655 1450 23669
rect 1446 23318 1450 23655
rect 1470 23627 1474 23892
rect 1470 23606 1477 23627
rect 1494 23606 1498 23892
rect 1518 23606 1522 23892
rect 1542 23606 1546 23892
rect 1566 23606 1570 23892
rect 1590 23606 1594 23892
rect 1614 23606 1618 23892
rect 1638 23606 1642 23892
rect 1662 23606 1666 23892
rect 1686 23606 1690 23892
rect 1710 23606 1714 23892
rect 1734 23606 1738 23892
rect 1758 23606 1762 23892
rect 1782 23606 1786 23892
rect 1806 23606 1810 23892
rect 1830 23606 1834 23892
rect 1854 23606 1858 23892
rect 1878 23606 1882 23892
rect 1902 23606 1906 23892
rect 1926 23799 1930 23892
rect 1915 23798 1949 23799
rect 1950 23798 1954 23892
rect 1974 23798 1978 23892
rect 1998 23798 2002 23892
rect 2022 23798 2026 23892
rect 2046 23798 2050 23892
rect 2070 23798 2074 23892
rect 2094 23798 2098 23892
rect 2118 23798 2122 23892
rect 2142 23798 2146 23892
rect 2166 23798 2170 23892
rect 2190 23798 2194 23892
rect 2214 23798 2218 23892
rect 2238 23798 2242 23892
rect 2262 23798 2266 23892
rect 2286 23798 2290 23892
rect 2310 23798 2314 23892
rect 2334 23798 2338 23892
rect 2358 23798 2362 23892
rect 2382 23798 2386 23892
rect 2406 23798 2410 23892
rect 2430 23798 2434 23892
rect 2443 23885 2448 23892
rect 2453 23871 2458 23885
rect 2454 23798 2458 23871
rect 2467 23798 2475 23799
rect 1915 23796 2475 23798
rect 1915 23789 1920 23796
rect 1926 23789 1930 23796
rect 1925 23775 1930 23789
rect 1915 23765 1920 23775
rect 1925 23751 1930 23765
rect 1926 23606 1930 23751
rect 1950 23723 1954 23796
rect 1950 23702 1957 23723
rect 1974 23702 1978 23796
rect 1998 23702 2002 23796
rect 2022 23702 2026 23796
rect 2046 23702 2050 23796
rect 2070 23702 2074 23796
rect 2094 23702 2098 23796
rect 2118 23702 2122 23796
rect 2142 23702 2146 23796
rect 2166 23702 2170 23796
rect 2190 23702 2194 23796
rect 2214 23702 2218 23796
rect 2238 23702 2242 23796
rect 2262 23702 2266 23796
rect 2286 23702 2290 23796
rect 2310 23702 2314 23796
rect 2334 23702 2338 23796
rect 2358 23702 2362 23796
rect 2382 23702 2386 23796
rect 2406 23702 2410 23796
rect 2430 23702 2434 23796
rect 2454 23702 2458 23796
rect 2461 23795 2475 23796
rect 2467 23789 2472 23795
rect 2477 23775 2482 23789
rect 2467 23717 2472 23727
rect 2478 23717 2482 23775
rect 2477 23703 2482 23717
rect 2491 23713 2499 23717
rect 2485 23703 2491 23713
rect 2467 23702 2499 23703
rect 1933 23700 2499 23702
rect 1933 23699 1947 23700
rect 1950 23675 1957 23700
rect 1950 23606 1954 23675
rect 1974 23606 1978 23700
rect 1998 23606 2002 23700
rect 2022 23606 2026 23700
rect 2046 23606 2050 23700
rect 2070 23606 2074 23700
rect 2094 23606 2098 23700
rect 2118 23606 2122 23700
rect 2142 23606 2146 23700
rect 2166 23606 2170 23700
rect 2190 23606 2194 23700
rect 2214 23606 2218 23700
rect 2238 23606 2242 23700
rect 2262 23606 2266 23700
rect 2286 23606 2290 23700
rect 2310 23606 2314 23700
rect 2334 23606 2338 23700
rect 2358 23606 2362 23700
rect 2382 23606 2386 23700
rect 2406 23606 2410 23700
rect 2430 23606 2434 23700
rect 2454 23606 2458 23700
rect 2467 23693 2472 23700
rect 2485 23699 2499 23700
rect 2477 23679 2482 23693
rect 2478 23606 2482 23679
rect 2491 23606 2499 23607
rect 1453 23604 2499 23606
rect 1453 23603 1467 23604
rect 1470 23579 1477 23604
rect 1470 23318 1474 23579
rect 1494 23318 1498 23604
rect 1518 23318 1522 23604
rect 1542 23318 1546 23604
rect 1566 23318 1570 23604
rect 1590 23318 1594 23604
rect 1614 23318 1618 23604
rect 1638 23318 1642 23604
rect 1662 23318 1666 23604
rect 1686 23318 1690 23604
rect 1710 23318 1714 23604
rect 1734 23318 1738 23604
rect 1758 23318 1762 23604
rect 1782 23318 1786 23604
rect 1806 23318 1810 23604
rect 1830 23318 1834 23604
rect 1854 23318 1858 23604
rect 1867 23333 1872 23343
rect 1878 23333 1882 23604
rect 1877 23319 1882 23333
rect 1878 23318 1882 23319
rect 1902 23318 1906 23604
rect 1926 23318 1930 23604
rect 1950 23318 1954 23604
rect 1974 23318 1978 23604
rect 1998 23318 2002 23604
rect 2022 23318 2026 23604
rect 2046 23318 2050 23604
rect 2070 23318 2074 23604
rect 2094 23318 2098 23604
rect 2118 23318 2122 23604
rect 2142 23318 2146 23604
rect 2166 23318 2170 23604
rect 2190 23318 2194 23604
rect 2214 23318 2218 23604
rect 2238 23318 2242 23604
rect 2262 23318 2266 23604
rect 2286 23318 2290 23604
rect 2310 23318 2314 23604
rect 2334 23318 2338 23604
rect 2358 23318 2362 23604
rect 2382 23318 2386 23604
rect 2406 23318 2410 23604
rect 2430 23318 2434 23604
rect 2443 23477 2448 23487
rect 2454 23477 2458 23604
rect 2453 23463 2458 23477
rect 2443 23453 2448 23463
rect 2453 23439 2458 23453
rect 2454 23318 2458 23439
rect 2478 23411 2482 23604
rect 2485 23603 2499 23604
rect 2491 23597 2496 23603
rect 2501 23583 2506 23597
rect 2478 23390 2485 23411
rect 2502 23390 2506 23583
rect 2515 23477 2520 23487
rect 2525 23463 2530 23477
rect 2515 23405 2520 23415
rect 2526 23405 2530 23463
rect 2525 23391 2530 23405
rect 2539 23401 2547 23405
rect 2533 23391 2539 23401
rect 2515 23390 2547 23391
rect 2461 23388 2547 23390
rect 2461 23387 2475 23388
rect 2478 23363 2485 23388
rect 2478 23318 2482 23363
rect 2502 23318 2506 23388
rect 2515 23381 2520 23388
rect 2533 23387 2547 23388
rect 2525 23367 2530 23381
rect 2526 23319 2530 23367
rect 2515 23318 2547 23319
rect -2393 23316 2547 23318
rect -2371 23270 -2366 23316
rect -2348 23270 -2343 23316
rect -2325 23270 -2320 23316
rect -2317 23312 -2309 23316
rect -2062 23312 -2054 23316
rect -2154 23308 -2138 23310
rect -2057 23308 -2054 23312
rect -2292 23302 -2054 23308
rect -2052 23302 -2044 23312
rect -2092 23286 -2062 23288
rect -2094 23282 -2062 23286
rect -2000 23270 -1992 23316
rect -1846 23309 -1806 23316
rect -1663 23312 -1655 23316
rect -1846 23302 -1680 23308
rect -1854 23286 -1806 23288
rect -1854 23282 -1680 23286
rect -1642 23270 -1637 23316
rect -1619 23270 -1614 23316
rect -1530 23270 -1526 23316
rect -1506 23270 -1502 23316
rect -1482 23270 -1478 23316
rect -1458 23270 -1454 23316
rect -1434 23315 -1430 23316
rect -2393 23268 -1437 23270
rect -2371 23246 -2366 23268
rect -2348 23246 -2343 23268
rect -2325 23246 -2320 23268
rect -2072 23266 -2036 23267
rect -2072 23260 -2054 23266
rect -2309 23252 -2301 23260
rect -2317 23246 -2309 23252
rect -2092 23251 -2062 23256
rect -2000 23247 -1992 23268
rect -1938 23267 -1906 23268
rect -1920 23266 -1906 23267
rect -1806 23260 -1680 23266
rect -1854 23251 -1806 23256
rect -1655 23252 -1647 23260
rect -1982 23247 -1966 23248
rect -2000 23246 -1966 23247
rect -1846 23246 -1806 23249
rect -1663 23246 -1655 23252
rect -1642 23246 -1637 23268
rect -1619 23246 -1614 23268
rect -1530 23246 -1526 23268
rect -1506 23246 -1502 23268
rect -1482 23246 -1478 23268
rect -1458 23246 -1454 23268
rect -1451 23267 -1437 23268
rect -1434 23267 -1427 23315
rect -1434 23246 -1430 23267
rect -1410 23246 -1406 23316
rect -1386 23246 -1382 23316
rect -1362 23246 -1358 23316
rect -1338 23246 -1334 23316
rect -1314 23246 -1310 23316
rect -1290 23246 -1286 23316
rect -1266 23246 -1262 23316
rect -1242 23246 -1238 23316
rect -1218 23246 -1214 23316
rect -1194 23246 -1190 23316
rect -1170 23246 -1166 23316
rect -1146 23246 -1142 23316
rect -1122 23246 -1118 23316
rect -1098 23246 -1094 23316
rect -1074 23246 -1070 23316
rect -1050 23246 -1046 23316
rect -1026 23246 -1022 23316
rect -1002 23246 -998 23316
rect -978 23246 -974 23316
rect -954 23246 -950 23316
rect -930 23246 -926 23316
rect -906 23246 -902 23316
rect -882 23246 -878 23316
rect -858 23246 -854 23316
rect -834 23246 -830 23316
rect -810 23246 -806 23316
rect -786 23246 -782 23316
rect -762 23246 -758 23316
rect -738 23246 -734 23316
rect -714 23246 -710 23316
rect -690 23246 -686 23316
rect -666 23246 -662 23316
rect -642 23246 -638 23316
rect -618 23246 -614 23316
rect -594 23246 -590 23316
rect -570 23246 -566 23316
rect -546 23246 -542 23316
rect -522 23246 -518 23316
rect -498 23246 -494 23316
rect -474 23246 -470 23316
rect -450 23246 -446 23316
rect -426 23246 -422 23316
rect -402 23246 -398 23316
rect -378 23246 -374 23316
rect -354 23246 -350 23316
rect -330 23246 -326 23316
rect -306 23246 -302 23316
rect -282 23246 -278 23316
rect -258 23246 -254 23316
rect -234 23246 -230 23316
rect -210 23246 -206 23316
rect -186 23246 -182 23316
rect -162 23246 -158 23316
rect -138 23246 -134 23316
rect -114 23246 -110 23316
rect -90 23246 -86 23316
rect -66 23246 -62 23316
rect -42 23246 -38 23316
rect -18 23246 -14 23316
rect 6 23246 10 23316
rect 30 23246 34 23316
rect 54 23246 58 23316
rect 78 23246 82 23316
rect 102 23246 106 23316
rect 126 23246 130 23316
rect 150 23246 154 23316
rect 174 23247 178 23316
rect 163 23246 197 23247
rect -2393 23244 197 23246
rect -2371 23222 -2366 23244
rect -2348 23222 -2343 23244
rect -2325 23222 -2320 23244
rect -2000 23242 -1966 23244
rect -2309 23224 -2301 23232
rect -2062 23231 -2054 23238
rect -2092 23224 -2084 23231
rect -2062 23224 -2026 23226
rect -2317 23222 -2309 23224
rect -2062 23222 -2012 23224
rect -2000 23222 -1992 23242
rect -1982 23241 -1966 23242
rect -1846 23240 -1806 23244
rect -1846 23233 -1798 23238
rect -1806 23231 -1798 23233
rect -1854 23229 -1846 23231
rect -1854 23224 -1806 23229
rect -1655 23224 -1647 23232
rect -1864 23222 -1796 23223
rect -1663 23222 -1655 23224
rect -1642 23222 -1637 23244
rect -1619 23222 -1614 23244
rect -1530 23222 -1526 23244
rect -1506 23222 -1502 23244
rect -1482 23222 -1478 23244
rect -1458 23222 -1454 23244
rect -1434 23222 -1430 23244
rect -1410 23222 -1406 23244
rect -1386 23222 -1382 23244
rect -1362 23222 -1358 23244
rect -1338 23222 -1334 23244
rect -1314 23222 -1310 23244
rect -1290 23222 -1286 23244
rect -1266 23222 -1262 23244
rect -1242 23222 -1238 23244
rect -1218 23222 -1214 23244
rect -1194 23222 -1190 23244
rect -1170 23222 -1166 23244
rect -1146 23222 -1142 23244
rect -1122 23222 -1118 23244
rect -1098 23222 -1094 23244
rect -1074 23222 -1070 23244
rect -1050 23222 -1046 23244
rect -1026 23222 -1022 23244
rect -1002 23222 -998 23244
rect -978 23222 -974 23244
rect -954 23222 -950 23244
rect -930 23222 -926 23244
rect -906 23222 -902 23244
rect -882 23222 -878 23244
rect -858 23222 -854 23244
rect -834 23222 -830 23244
rect -810 23222 -806 23244
rect -786 23222 -782 23244
rect -762 23222 -758 23244
rect -738 23222 -734 23244
rect -714 23222 -710 23244
rect -690 23222 -686 23244
rect -666 23222 -662 23244
rect -642 23222 -638 23244
rect -618 23222 -614 23244
rect -594 23222 -590 23244
rect -570 23222 -566 23244
rect -546 23222 -542 23244
rect -522 23222 -518 23244
rect -498 23222 -494 23244
rect -474 23222 -470 23244
rect -450 23222 -446 23244
rect -426 23222 -422 23244
rect -402 23222 -398 23244
rect -378 23222 -374 23244
rect -354 23222 -350 23244
rect -330 23222 -326 23244
rect -306 23222 -302 23244
rect -282 23222 -278 23244
rect -258 23222 -254 23244
rect -234 23222 -230 23244
rect -210 23222 -206 23244
rect -186 23222 -182 23244
rect -162 23222 -158 23244
rect -138 23222 -134 23244
rect -114 23222 -110 23244
rect -90 23222 -86 23244
rect -66 23222 -62 23244
rect -42 23222 -38 23244
rect -18 23222 -14 23244
rect 6 23222 10 23244
rect 30 23222 34 23244
rect 54 23222 58 23244
rect 78 23222 82 23244
rect 102 23222 106 23244
rect 126 23222 130 23244
rect 150 23222 154 23244
rect 163 23237 168 23244
rect 174 23237 178 23244
rect 173 23223 178 23237
rect 174 23222 178 23223
rect 198 23222 202 23316
rect 222 23222 226 23316
rect 246 23222 250 23316
rect 270 23222 274 23316
rect 294 23222 298 23316
rect 318 23222 322 23316
rect 342 23222 346 23316
rect 366 23222 370 23316
rect 390 23222 394 23316
rect 414 23222 418 23316
rect 438 23222 442 23316
rect 462 23222 466 23316
rect 486 23222 490 23316
rect 510 23222 514 23316
rect 534 23222 538 23316
rect 558 23222 562 23316
rect 582 23222 586 23316
rect 606 23222 610 23316
rect 630 23222 634 23316
rect 654 23222 658 23316
rect 678 23222 682 23316
rect 702 23222 706 23316
rect 726 23222 730 23316
rect 750 23222 754 23316
rect 774 23222 778 23316
rect 798 23222 802 23316
rect 822 23222 826 23316
rect 846 23222 850 23316
rect 870 23222 874 23316
rect 894 23222 898 23316
rect 918 23222 922 23316
rect 942 23222 946 23316
rect 966 23295 970 23316
rect 955 23294 989 23295
rect 990 23294 994 23316
rect 1014 23294 1018 23316
rect 1038 23294 1042 23316
rect 1062 23294 1066 23316
rect 1086 23294 1090 23316
rect 1110 23294 1114 23316
rect 1134 23294 1138 23316
rect 1158 23294 1162 23316
rect 1182 23294 1186 23316
rect 1206 23294 1210 23316
rect 1230 23294 1234 23316
rect 1254 23294 1258 23316
rect 1278 23294 1282 23316
rect 1302 23294 1306 23316
rect 1326 23294 1330 23316
rect 1350 23294 1354 23316
rect 1374 23294 1378 23316
rect 1398 23294 1402 23316
rect 1422 23294 1426 23316
rect 1446 23294 1450 23316
rect 1470 23294 1474 23316
rect 1494 23294 1498 23316
rect 1518 23294 1522 23316
rect 1542 23294 1546 23316
rect 1566 23294 1570 23316
rect 1590 23294 1594 23316
rect 1614 23294 1618 23316
rect 1638 23294 1642 23316
rect 1662 23294 1666 23316
rect 1686 23294 1690 23316
rect 1710 23294 1714 23316
rect 1734 23294 1738 23316
rect 1758 23294 1762 23316
rect 1782 23294 1786 23316
rect 1806 23294 1810 23316
rect 1830 23294 1834 23316
rect 1854 23294 1858 23316
rect 1878 23294 1882 23316
rect 1902 23294 1906 23316
rect 1926 23294 1930 23316
rect 1950 23294 1954 23316
rect 1974 23294 1978 23316
rect 1998 23294 2002 23316
rect 2022 23294 2026 23316
rect 2046 23294 2050 23316
rect 2070 23294 2074 23316
rect 2094 23294 2098 23316
rect 2118 23294 2122 23316
rect 2142 23294 2146 23316
rect 2166 23294 2170 23316
rect 2190 23294 2194 23316
rect 2214 23294 2218 23316
rect 2238 23294 2242 23316
rect 2262 23294 2266 23316
rect 2286 23294 2290 23316
rect 2310 23294 2314 23316
rect 2334 23294 2338 23316
rect 2358 23294 2362 23316
rect 2382 23294 2386 23316
rect 2406 23294 2410 23316
rect 2430 23294 2434 23316
rect 2454 23294 2458 23316
rect 2478 23294 2482 23316
rect 2502 23294 2506 23316
rect 2515 23309 2520 23316
rect 2526 23309 2530 23316
rect 2533 23315 2547 23316
rect 2525 23295 2530 23309
rect 2539 23305 2547 23309
rect 2533 23295 2539 23305
rect 2515 23294 2547 23295
rect 955 23292 2547 23294
rect 955 23285 960 23292
rect 966 23285 970 23292
rect 965 23271 970 23285
rect 955 23261 960 23271
rect 965 23247 970 23261
rect 966 23222 970 23247
rect 990 23222 994 23292
rect 1014 23222 1018 23292
rect 1038 23222 1042 23292
rect 1062 23222 1066 23292
rect 1086 23222 1090 23292
rect 1110 23222 1114 23292
rect 1134 23222 1138 23292
rect 1158 23222 1162 23292
rect 1182 23222 1186 23292
rect 1206 23222 1210 23292
rect 1230 23222 1234 23292
rect 1254 23222 1258 23292
rect 1278 23222 1282 23292
rect 1302 23222 1306 23292
rect 1326 23222 1330 23292
rect 1350 23222 1354 23292
rect 1374 23222 1378 23292
rect 1398 23222 1402 23292
rect 1422 23222 1426 23292
rect 1446 23222 1450 23292
rect 1470 23222 1474 23292
rect 1494 23222 1498 23292
rect 1518 23222 1522 23292
rect 1542 23222 1546 23292
rect 1566 23222 1570 23292
rect 1590 23222 1594 23292
rect 1614 23222 1618 23292
rect 1638 23222 1642 23292
rect 1662 23222 1666 23292
rect 1686 23222 1690 23292
rect 1710 23222 1714 23292
rect 1734 23222 1738 23292
rect 1758 23222 1762 23292
rect 1782 23222 1786 23292
rect 1806 23222 1810 23292
rect 1830 23222 1834 23292
rect 1854 23222 1858 23292
rect 1878 23222 1882 23292
rect 1902 23267 1906 23292
rect 1902 23243 1909 23267
rect 1902 23222 1906 23243
rect 1926 23222 1930 23292
rect 1950 23222 1954 23292
rect 1974 23222 1978 23292
rect 1998 23222 2002 23292
rect 2022 23222 2026 23292
rect 2046 23222 2050 23292
rect 2070 23222 2074 23292
rect 2094 23222 2098 23292
rect 2118 23222 2122 23292
rect 2142 23222 2146 23292
rect 2166 23222 2170 23292
rect 2190 23222 2194 23292
rect 2214 23222 2218 23292
rect 2238 23222 2242 23292
rect 2262 23222 2266 23292
rect 2286 23222 2290 23292
rect 2310 23222 2314 23292
rect 2334 23222 2338 23292
rect 2358 23222 2362 23292
rect 2382 23222 2386 23292
rect 2406 23222 2410 23292
rect 2430 23222 2434 23292
rect 2454 23222 2458 23292
rect 2478 23222 2482 23292
rect 2502 23222 2506 23292
rect 2515 23285 2520 23292
rect 2533 23291 2547 23292
rect 2525 23271 2530 23285
rect 2526 23223 2530 23271
rect 2515 23222 2547 23223
rect -2393 23220 2547 23222
rect -2371 23174 -2366 23220
rect -2348 23174 -2343 23220
rect -2325 23174 -2320 23220
rect -2317 23216 -2309 23220
rect -2062 23216 -2054 23220
rect -2154 23212 -2138 23214
rect -2057 23212 -2054 23216
rect -2292 23206 -2054 23212
rect -2052 23206 -2044 23216
rect -2092 23190 -2062 23192
rect -2094 23186 -2062 23190
rect -2000 23174 -1992 23220
rect -1846 23213 -1806 23220
rect -1663 23216 -1655 23220
rect -1846 23206 -1680 23212
rect -1854 23190 -1806 23192
rect -1854 23186 -1680 23190
rect -1979 23174 -1945 23176
rect -1642 23174 -1637 23220
rect -1619 23174 -1614 23220
rect -1530 23174 -1526 23220
rect -1506 23174 -1502 23220
rect -1482 23174 -1478 23220
rect -1458 23174 -1454 23220
rect -1434 23174 -1430 23220
rect -1410 23174 -1406 23220
rect -1386 23174 -1382 23220
rect -1362 23174 -1358 23220
rect -1338 23174 -1334 23220
rect -1314 23174 -1310 23220
rect -1290 23174 -1286 23220
rect -1266 23174 -1262 23220
rect -1242 23174 -1238 23220
rect -1218 23174 -1214 23220
rect -1194 23174 -1190 23220
rect -1170 23174 -1166 23220
rect -1146 23174 -1142 23220
rect -1122 23174 -1118 23220
rect -1098 23174 -1094 23220
rect -1074 23174 -1070 23220
rect -1050 23174 -1046 23220
rect -1026 23174 -1022 23220
rect -1002 23174 -998 23220
rect -978 23174 -974 23220
rect -954 23174 -950 23220
rect -930 23174 -926 23220
rect -906 23174 -902 23220
rect -882 23174 -878 23220
rect -858 23174 -854 23220
rect -845 23189 -840 23199
rect -834 23189 -830 23220
rect -835 23175 -830 23189
rect -845 23174 -811 23175
rect -2393 23172 -811 23174
rect -2371 23126 -2366 23172
rect -2348 23126 -2343 23172
rect -2325 23126 -2320 23172
rect -2080 23171 -1906 23172
rect -2080 23170 -2036 23171
rect -2080 23164 -2054 23170
rect -2309 23156 -2301 23162
rect -2317 23146 -2309 23156
rect -2070 23155 -2040 23162
rect -2054 23147 -2040 23150
rect -2000 23145 -1992 23171
rect -1920 23170 -1906 23171
rect -1850 23164 -1846 23172
rect -1840 23164 -1792 23172
rect -1969 23152 -1966 23161
rect -1850 23157 -1802 23162
rect -1906 23155 -1802 23157
rect -1655 23156 -1647 23162
rect -1906 23154 -1850 23155
rect -1846 23147 -1802 23153
rect -1663 23146 -1655 23156
rect -1860 23145 -1798 23146
rect -2078 23138 -2070 23145
rect -2309 23128 -2301 23134
rect -2317 23126 -2309 23128
rect -2154 23126 -2145 23136
rect -2044 23135 -2040 23140
rect -2028 23138 -1945 23145
rect -1929 23138 -1794 23145
rect -2070 23128 -2040 23135
rect -2044 23126 -2028 23128
rect -2000 23126 -1992 23138
rect -1860 23137 -1798 23138
rect -1850 23128 -1802 23135
rect -1655 23128 -1647 23134
rect -1978 23126 -1942 23127
rect -1663 23126 -1655 23128
rect -1642 23126 -1637 23172
rect -1619 23126 -1614 23172
rect -1530 23126 -1526 23172
rect -1506 23126 -1502 23172
rect -1482 23126 -1478 23172
rect -1458 23126 -1454 23172
rect -1434 23126 -1430 23172
rect -1410 23126 -1406 23172
rect -1386 23126 -1382 23172
rect -1362 23126 -1358 23172
rect -1338 23126 -1334 23172
rect -1314 23126 -1310 23172
rect -1290 23126 -1286 23172
rect -1266 23126 -1262 23172
rect -1242 23126 -1238 23172
rect -1218 23126 -1214 23172
rect -1194 23126 -1190 23172
rect -1170 23126 -1166 23172
rect -1146 23126 -1142 23172
rect -1122 23126 -1118 23172
rect -1098 23126 -1094 23172
rect -1074 23126 -1070 23172
rect -1050 23126 -1046 23172
rect -1026 23126 -1022 23172
rect -1002 23126 -998 23172
rect -978 23126 -974 23172
rect -954 23126 -950 23172
rect -930 23126 -926 23172
rect -906 23126 -902 23172
rect -882 23126 -878 23172
rect -858 23126 -854 23172
rect -845 23165 -840 23172
rect -835 23151 -830 23165
rect -834 23126 -830 23151
rect -810 23126 -806 23220
rect -786 23126 -782 23220
rect -762 23126 -758 23220
rect -738 23126 -734 23220
rect -714 23126 -710 23220
rect -690 23126 -686 23220
rect -666 23126 -662 23220
rect -642 23126 -638 23220
rect -618 23126 -614 23220
rect -594 23126 -590 23220
rect -570 23126 -566 23220
rect -546 23126 -542 23220
rect -522 23126 -518 23220
rect -498 23126 -494 23220
rect -474 23126 -470 23220
rect -450 23126 -446 23220
rect -426 23126 -422 23220
rect -402 23126 -398 23220
rect -378 23126 -374 23220
rect -354 23126 -350 23220
rect -330 23126 -326 23220
rect -306 23126 -302 23220
rect -282 23126 -278 23220
rect -258 23126 -254 23220
rect -234 23126 -230 23220
rect -210 23126 -206 23220
rect -186 23126 -182 23220
rect -162 23126 -158 23220
rect -138 23126 -134 23220
rect -114 23126 -110 23220
rect -90 23126 -86 23220
rect -66 23126 -62 23220
rect -42 23126 -38 23220
rect -18 23126 -14 23220
rect 6 23126 10 23220
rect 30 23126 34 23220
rect 54 23126 58 23220
rect 78 23126 82 23220
rect 102 23126 106 23220
rect 126 23126 130 23220
rect 150 23126 154 23220
rect 174 23126 178 23220
rect 198 23171 202 23220
rect 198 23147 205 23171
rect 198 23126 202 23147
rect 222 23126 226 23220
rect 246 23126 250 23220
rect 270 23126 274 23220
rect 294 23126 298 23220
rect 318 23126 322 23220
rect 342 23126 346 23220
rect 366 23126 370 23220
rect 390 23126 394 23220
rect 414 23126 418 23220
rect 438 23126 442 23220
rect 462 23126 466 23220
rect 486 23126 490 23220
rect 510 23126 514 23220
rect 534 23126 538 23220
rect 558 23126 562 23220
rect 582 23126 586 23220
rect 606 23126 610 23220
rect 630 23126 634 23220
rect 654 23126 658 23220
rect 678 23126 682 23220
rect 702 23126 706 23220
rect 726 23126 730 23220
rect 750 23126 754 23220
rect 774 23126 778 23220
rect 798 23126 802 23220
rect 822 23126 826 23220
rect 846 23126 850 23220
rect 870 23126 874 23220
rect 894 23126 898 23220
rect 918 23126 922 23220
rect 942 23126 946 23220
rect 966 23126 970 23220
rect 990 23219 994 23220
rect 990 23198 997 23219
rect 1014 23198 1018 23220
rect 1038 23198 1042 23220
rect 1062 23198 1066 23220
rect 1086 23198 1090 23220
rect 1110 23198 1114 23220
rect 1134 23198 1138 23220
rect 1158 23198 1162 23220
rect 1182 23198 1186 23220
rect 1206 23198 1210 23220
rect 1230 23198 1234 23220
rect 1254 23198 1258 23220
rect 1278 23198 1282 23220
rect 1302 23198 1306 23220
rect 1326 23198 1330 23220
rect 1350 23198 1354 23220
rect 1374 23198 1378 23220
rect 1398 23198 1402 23220
rect 1422 23198 1426 23220
rect 1446 23198 1450 23220
rect 1470 23198 1474 23220
rect 1494 23198 1498 23220
rect 1518 23198 1522 23220
rect 1542 23198 1546 23220
rect 1566 23198 1570 23220
rect 1590 23198 1594 23220
rect 1614 23198 1618 23220
rect 1638 23198 1642 23220
rect 1662 23198 1666 23220
rect 1686 23198 1690 23220
rect 1710 23198 1714 23220
rect 1734 23198 1738 23220
rect 1758 23198 1762 23220
rect 1782 23198 1786 23220
rect 1806 23198 1810 23220
rect 1830 23198 1834 23220
rect 1854 23198 1858 23220
rect 1878 23198 1882 23220
rect 1902 23198 1906 23220
rect 1926 23198 1930 23220
rect 1950 23198 1954 23220
rect 1974 23198 1978 23220
rect 1998 23198 2002 23220
rect 2022 23198 2026 23220
rect 2046 23198 2050 23220
rect 2070 23198 2074 23220
rect 2094 23198 2098 23220
rect 2118 23198 2122 23220
rect 2142 23198 2146 23220
rect 2166 23198 2170 23220
rect 2190 23198 2194 23220
rect 2214 23198 2218 23220
rect 2238 23198 2242 23220
rect 2262 23198 2266 23220
rect 2286 23198 2290 23220
rect 2310 23198 2314 23220
rect 2334 23198 2338 23220
rect 2358 23198 2362 23220
rect 2382 23198 2386 23220
rect 2406 23198 2410 23220
rect 2430 23198 2434 23220
rect 2454 23198 2458 23220
rect 2478 23198 2482 23220
rect 2502 23198 2506 23220
rect 2515 23213 2520 23220
rect 2526 23213 2530 23220
rect 2533 23219 2547 23220
rect 2525 23199 2530 23213
rect 2539 23209 2547 23213
rect 2533 23199 2539 23209
rect 2515 23198 2547 23199
rect 973 23196 2547 23198
rect 973 23195 987 23196
rect 990 23171 997 23196
rect 990 23126 994 23171
rect 1014 23126 1018 23196
rect 1038 23126 1042 23196
rect 1062 23126 1066 23196
rect 1086 23126 1090 23196
rect 1110 23126 1114 23196
rect 1134 23126 1138 23196
rect 1158 23126 1162 23196
rect 1182 23126 1186 23196
rect 1206 23126 1210 23196
rect 1230 23126 1234 23196
rect 1254 23126 1258 23196
rect 1278 23126 1282 23196
rect 1302 23126 1306 23196
rect 1326 23126 1330 23196
rect 1350 23126 1354 23196
rect 1374 23126 1378 23196
rect 1398 23127 1402 23196
rect 1387 23126 1421 23127
rect -2393 23124 1421 23126
rect -2371 23030 -2366 23124
rect -2348 23030 -2343 23124
rect -2325 23086 -2320 23124
rect -2317 23118 -2309 23124
rect -2145 23120 -2138 23124
rect -2070 23120 -2054 23124
rect -2078 23111 -2054 23118
rect -2062 23086 -2032 23087
rect -2000 23086 -1992 23124
rect -1846 23120 -1802 23124
rect -1846 23110 -1792 23119
rect -1663 23118 -1655 23124
rect -1942 23088 -1937 23100
rect -1850 23097 -1822 23098
rect -1850 23093 -1802 23097
rect -2325 23078 -2317 23086
rect -2062 23084 -1961 23086
rect -2325 23058 -2320 23078
rect -2317 23070 -2309 23078
rect -2062 23071 -2040 23082
rect -2032 23077 -1961 23084
rect -1947 23078 -1942 23086
rect -1842 23084 -1794 23087
rect -2070 23066 -2022 23070
rect -2325 23044 -2317 23058
rect -2072 23050 -2032 23051
rect -2102 23044 -2032 23050
rect -2325 23030 -2320 23044
rect -2317 23042 -2309 23044
rect -2309 23030 -2301 23042
rect -2070 23035 -2062 23040
rect -2000 23030 -1992 23077
rect -1942 23076 -1937 23078
rect -1932 23068 -1927 23076
rect -1912 23073 -1896 23079
rect -1842 23071 -1802 23082
rect -1671 23078 -1663 23086
rect -1663 23070 -1655 23078
rect -1850 23066 -1680 23070
rect -1924 23052 -1921 23054
rect -1806 23044 -1680 23050
rect -1671 23044 -1663 23058
rect -1663 23042 -1655 23044
rect -1854 23035 -1806 23040
rect -1974 23030 -1964 23031
rect -1960 23030 -1944 23032
rect -1842 23030 -1806 23033
rect -1655 23030 -1647 23042
rect -1642 23030 -1637 23124
rect -1619 23030 -1614 23124
rect -1530 23030 -1526 23124
rect -1517 23093 -1512 23103
rect -1506 23093 -1502 23124
rect -1507 23079 -1502 23093
rect -1506 23030 -1502 23079
rect -1482 23030 -1478 23124
rect -1458 23030 -1454 23124
rect -1434 23030 -1430 23124
rect -1410 23030 -1406 23124
rect -1386 23030 -1382 23124
rect -1362 23030 -1358 23124
rect -1338 23030 -1334 23124
rect -1314 23030 -1310 23124
rect -1290 23030 -1286 23124
rect -1266 23030 -1262 23124
rect -1242 23030 -1238 23124
rect -1218 23030 -1214 23124
rect -1194 23030 -1190 23124
rect -1170 23030 -1166 23124
rect -1146 23030 -1142 23124
rect -1122 23030 -1118 23124
rect -1098 23030 -1094 23124
rect -1074 23030 -1070 23124
rect -1050 23031 -1046 23124
rect -1061 23030 -1027 23031
rect -2393 23028 -1027 23030
rect -2371 23006 -2366 23028
rect -2348 23006 -2343 23028
rect -2325 23016 -2317 23028
rect -2325 23006 -2320 23016
rect -2317 23014 -2309 23016
rect -2062 23015 -2032 23022
rect -2309 23006 -2301 23014
rect -2070 23008 -2062 23015
rect -2000 23010 -1992 23028
rect -1974 23026 -1944 23028
rect -1960 23025 -1944 23026
rect -1842 23024 -1806 23028
rect -1842 23017 -1798 23022
rect -1806 23015 -1798 23017
rect -1671 23016 -1663 23028
rect -1854 23013 -1842 23015
rect -1663 23014 -1655 23016
rect -2062 23006 -2036 23008
rect -2393 23004 -2036 23006
rect -2032 23006 -2012 23008
rect -2004 23006 -1974 23010
rect -1854 23008 -1806 23013
rect -1864 23006 -1796 23007
rect -1655 23006 -1647 23014
rect -1642 23006 -1637 23028
rect -1619 23006 -1614 23028
rect -1530 23006 -1526 23028
rect -1506 23007 -1502 23028
rect -1482 23027 -1478 23028
rect -1517 23006 -1485 23007
rect -2032 23004 -1485 23006
rect -2371 22934 -2366 23004
rect -2348 22934 -2343 23004
rect -2325 23000 -2320 23004
rect -2309 23002 -2301 23004
rect -2317 23000 -2309 23002
rect -2325 22988 -2317 23000
rect -2052 22998 -2036 23000
rect -2052 22996 -2032 22998
rect -2062 22990 -2032 22996
rect -2325 22934 -2320 22988
rect -2317 22986 -2309 22988
rect -2092 22974 -2062 22976
rect -2094 22970 -2062 22974
rect -2309 22940 -2301 22946
rect -2317 22934 -2309 22940
rect -2000 22934 -1992 23004
rect -1904 22997 -1874 23004
rect -1842 22997 -1806 23004
rect -1655 23002 -1647 23004
rect -1663 23000 -1655 23002
rect -1842 22990 -1680 22996
rect -1671 22988 -1663 23000
rect -1663 22986 -1655 22988
rect -1854 22974 -1806 22976
rect -1854 22970 -1680 22974
rect -1655 22940 -1647 22946
rect -1663 22934 -1655 22940
rect -1642 22934 -1637 23004
rect -1619 22934 -1614 23004
rect -1530 22934 -1526 23004
rect -1517 22997 -1512 23004
rect -1506 22997 -1502 23004
rect -1499 23003 -1485 23004
rect -1482 23003 -1475 23027
rect -1507 22983 -1502 22997
rect -1506 22934 -1502 22983
rect -1482 22934 -1478 23003
rect -1458 22934 -1454 23028
rect -1434 22934 -1430 23028
rect -1410 22934 -1406 23028
rect -1386 22934 -1382 23028
rect -1362 22934 -1358 23028
rect -1338 22934 -1334 23028
rect -1314 22934 -1310 23028
rect -1290 22934 -1286 23028
rect -1266 22934 -1262 23028
rect -1242 22934 -1238 23028
rect -1218 22934 -1214 23028
rect -1194 22934 -1190 23028
rect -1170 22934 -1166 23028
rect -1146 22934 -1142 23028
rect -1122 22934 -1118 23028
rect -1098 22934 -1094 23028
rect -1074 22934 -1070 23028
rect -1061 23021 -1056 23028
rect -1050 23021 -1046 23028
rect -1051 23007 -1046 23021
rect -1050 22934 -1046 23007
rect -1026 22955 -1022 23124
rect -2393 22932 -1029 22934
rect -2371 22838 -2366 22932
rect -2348 22838 -2343 22932
rect -2325 22870 -2320 22932
rect -2317 22930 -2309 22932
rect -2000 22931 -1966 22932
rect -2000 22930 -1982 22931
rect -1663 22930 -1655 22932
rect -2028 22922 -2018 22924
rect -2309 22912 -2301 22918
rect -2091 22912 -2061 22919
rect -2317 22902 -2309 22912
rect -2044 22910 -2028 22912
rect -2026 22910 -2014 22922
rect -2084 22904 -2061 22910
rect -2044 22908 -2014 22910
rect -2292 22894 -2054 22903
rect -2325 22862 -2317 22870
rect -2325 22842 -2320 22862
rect -2317 22854 -2309 22862
rect -2325 22838 -2317 22842
rect -2000 22838 -1992 22930
rect -1982 22929 -1966 22930
rect -1980 22912 -1932 22919
rect -1655 22912 -1647 22918
rect -1846 22894 -1680 22903
rect -1663 22902 -1655 22912
rect -1671 22862 -1663 22870
rect -1663 22854 -1655 22862
rect -1671 22838 -1663 22842
rect -1642 22838 -1637 22932
rect -1619 22838 -1614 22932
rect -1530 22838 -1526 22932
rect -1506 22838 -1502 22932
rect -1482 22931 -1478 22932
rect -1482 22907 -1475 22931
rect -1482 22838 -1478 22907
rect -1458 22838 -1454 22932
rect -1434 22838 -1430 22932
rect -1410 22838 -1406 22932
rect -1386 22838 -1382 22932
rect -1362 22838 -1358 22932
rect -1338 22838 -1334 22932
rect -1314 22838 -1310 22932
rect -1290 22838 -1286 22932
rect -1266 22838 -1262 22932
rect -1242 22838 -1238 22932
rect -1218 22838 -1214 22932
rect -1194 22838 -1190 22932
rect -1170 22838 -1166 22932
rect -1146 22838 -1142 22932
rect -1122 22838 -1118 22932
rect -1098 22838 -1094 22932
rect -1074 22838 -1070 22932
rect -1050 22838 -1046 22932
rect -1043 22931 -1029 22932
rect -1026 22931 -1019 22955
rect -1026 22838 -1022 22931
rect -1002 22838 -998 23124
rect -978 22838 -974 23124
rect -954 22838 -950 23124
rect -930 22838 -926 23124
rect -906 22838 -902 23124
rect -882 22838 -878 23124
rect -858 22838 -854 23124
rect -834 22838 -830 23124
rect -810 23123 -806 23124
rect -810 23075 -803 23123
rect -810 22838 -806 23075
rect -786 22838 -782 23124
rect -762 22838 -758 23124
rect -738 22838 -734 23124
rect -714 22838 -710 23124
rect -690 22838 -686 23124
rect -666 22838 -662 23124
rect -642 22838 -638 23124
rect -618 22838 -614 23124
rect -594 22838 -590 23124
rect -570 22838 -566 23124
rect -546 22838 -542 23124
rect -522 22838 -518 23124
rect -498 22838 -494 23124
rect -474 22838 -470 23124
rect -450 22838 -446 23124
rect -426 22838 -422 23124
rect -402 22838 -398 23124
rect -378 22838 -374 23124
rect -354 22838 -350 23124
rect -330 22838 -326 23124
rect -306 22838 -302 23124
rect -282 22838 -278 23124
rect -258 22838 -254 23124
rect -234 22838 -230 23124
rect -210 22838 -206 23124
rect -186 22838 -182 23124
rect -162 22838 -158 23124
rect -138 22838 -134 23124
rect -114 22838 -110 23124
rect -90 22838 -86 23124
rect -66 22838 -62 23124
rect -42 22838 -38 23124
rect -18 22838 -14 23124
rect 6 22838 10 23124
rect 30 22838 34 23124
rect 54 22838 58 23124
rect 78 22838 82 23124
rect 102 22838 106 23124
rect 126 22838 130 23124
rect 150 22838 154 23124
rect 174 22838 178 23124
rect 198 22838 202 23124
rect 222 22838 226 23124
rect 246 22838 250 23124
rect 270 22838 274 23124
rect 294 22838 298 23124
rect 318 22838 322 23124
rect 342 22838 346 23124
rect 366 22838 370 23124
rect 390 22838 394 23124
rect 414 22838 418 23124
rect 438 22838 442 23124
rect 462 22838 466 23124
rect 486 22838 490 23124
rect 510 22838 514 23124
rect 534 22838 538 23124
rect 558 22838 562 23124
rect 582 22838 586 23124
rect 606 22838 610 23124
rect 630 22838 634 23124
rect 654 22838 658 23124
rect 678 22838 682 23124
rect 702 22838 706 23124
rect 726 22838 730 23124
rect 750 22838 754 23124
rect 774 22838 778 23124
rect 798 22838 802 23124
rect 822 22838 826 23124
rect 846 22838 850 23124
rect 870 22838 874 23124
rect 894 22838 898 23124
rect 918 22838 922 23124
rect 942 22838 946 23124
rect 966 22838 970 23124
rect 990 22838 994 23124
rect 1014 22838 1018 23124
rect 1038 22838 1042 23124
rect 1062 22838 1066 23124
rect 1086 22838 1090 23124
rect 1110 22838 1114 23124
rect 1134 22838 1138 23124
rect 1158 22838 1162 23124
rect 1182 22838 1186 23124
rect 1206 22838 1210 23124
rect 1230 22838 1234 23124
rect 1254 22838 1258 23124
rect 1267 22877 1272 22887
rect 1278 22877 1282 23124
rect 1277 22863 1282 22877
rect 1278 22838 1282 22863
rect 1302 22838 1306 23124
rect 1326 22838 1330 23124
rect 1350 22838 1354 23124
rect 1374 22838 1378 23124
rect 1387 23117 1392 23124
rect 1398 23117 1402 23124
rect 1397 23103 1402 23117
rect 1398 22838 1402 23103
rect 1422 23051 1426 23196
rect 1422 23027 1429 23051
rect 1422 22838 1426 23027
rect 1446 22838 1450 23196
rect 1459 23069 1464 23079
rect 1470 23069 1474 23196
rect 1469 23055 1474 23069
rect 1459 23045 1464 23055
rect 1469 23031 1474 23045
rect 1470 22838 1474 23031
rect 1494 23003 1498 23196
rect 1483 22955 1491 22959
rect 1494 22955 1501 23003
rect 1483 22949 1488 22955
rect 1494 22949 1498 22955
rect 1493 22935 1498 22949
rect 1483 22925 1488 22935
rect 1493 22911 1498 22925
rect 1494 22838 1498 22911
rect 1518 22883 1522 23196
rect -2393 22836 1515 22838
rect -2371 22790 -2366 22836
rect -2348 22790 -2343 22836
rect -2325 22828 -2317 22836
rect -2018 22835 -2004 22836
rect -2000 22835 -1992 22836
rect -2072 22834 -1928 22835
rect -2072 22828 -2053 22834
rect -2325 22812 -2320 22828
rect -2317 22826 -2309 22828
rect -2309 22814 -2301 22826
rect -2092 22819 -2062 22824
rect -2317 22812 -2309 22814
rect -2325 22800 -2317 22812
rect -2098 22806 -2096 22817
rect -2092 22806 -2084 22819
rect -2000 22818 -1992 22834
rect -1972 22828 -1928 22834
rect -1924 22828 -1918 22836
rect -1671 22828 -1663 22836
rect -1663 22826 -1655 22828
rect -2083 22808 -2062 22817
rect -2027 22816 -1992 22818
rect -2018 22808 -2002 22816
rect -2000 22808 -1992 22816
rect -2100 22801 -2096 22806
rect -2083 22801 -2053 22806
rect -2003 22804 -1990 22808
rect -1972 22806 -1964 22815
rect -1928 22814 -1924 22817
rect -1655 22814 -1647 22826
rect -1663 22812 -1655 22814
rect -2325 22790 -2320 22800
rect -2317 22798 -2309 22800
rect -2309 22790 -2301 22798
rect -2004 22794 -2003 22804
rect -2062 22790 -2012 22792
rect -2000 22790 -1992 22804
rect -1972 22801 -1924 22806
rect -1864 22801 -1796 22807
rect -1671 22800 -1663 22812
rect -1663 22798 -1655 22800
rect -1864 22790 -1796 22791
rect -1655 22790 -1647 22798
rect -1642 22790 -1637 22836
rect -1619 22790 -1614 22836
rect -1530 22790 -1526 22836
rect -1506 22790 -1502 22836
rect -1482 22790 -1478 22836
rect -1458 22790 -1454 22836
rect -1434 22790 -1430 22836
rect -1410 22790 -1406 22836
rect -1386 22790 -1382 22836
rect -1362 22790 -1358 22836
rect -1338 22790 -1334 22836
rect -1314 22790 -1310 22836
rect -1290 22790 -1286 22836
rect -1266 22790 -1262 22836
rect -1242 22790 -1238 22836
rect -1218 22790 -1214 22836
rect -1194 22790 -1190 22836
rect -1170 22790 -1166 22836
rect -1146 22790 -1142 22836
rect -1122 22790 -1118 22836
rect -1098 22790 -1094 22836
rect -1074 22790 -1070 22836
rect -1050 22790 -1046 22836
rect -1026 22790 -1022 22836
rect -1002 22790 -998 22836
rect -978 22790 -974 22836
rect -954 22790 -950 22836
rect -930 22790 -926 22836
rect -906 22790 -902 22836
rect -882 22790 -878 22836
rect -858 22790 -854 22836
rect -834 22790 -830 22836
rect -810 22790 -806 22836
rect -786 22790 -782 22836
rect -762 22790 -758 22836
rect -738 22790 -734 22836
rect -714 22790 -710 22836
rect -690 22790 -686 22836
rect -666 22790 -662 22836
rect -642 22790 -638 22836
rect -618 22790 -614 22836
rect -594 22790 -590 22836
rect -570 22790 -566 22836
rect -546 22790 -542 22836
rect -522 22790 -518 22836
rect -498 22790 -494 22836
rect -474 22790 -470 22836
rect -450 22790 -446 22836
rect -426 22790 -422 22836
rect -402 22791 -398 22836
rect -413 22790 -379 22791
rect -2393 22788 -379 22790
rect -2371 22742 -2366 22788
rect -2348 22742 -2343 22788
rect -2325 22784 -2320 22788
rect -2309 22786 -2301 22788
rect -2317 22784 -2309 22786
rect -2325 22772 -2317 22784
rect -2325 22742 -2320 22772
rect -2317 22770 -2309 22772
rect -2092 22758 -2062 22760
rect -2094 22754 -2062 22758
rect -2000 22742 -1992 22788
rect -1655 22786 -1647 22788
rect -1663 22784 -1655 22786
rect -1671 22772 -1663 22784
rect -1663 22770 -1655 22772
rect -1854 22758 -1806 22760
rect -1854 22754 -1680 22758
rect -1642 22742 -1637 22788
rect -1619 22742 -1614 22788
rect -1530 22742 -1526 22788
rect -1506 22742 -1502 22788
rect -1482 22742 -1478 22788
rect -1458 22742 -1454 22788
rect -1434 22742 -1430 22788
rect -1410 22742 -1406 22788
rect -1386 22742 -1382 22788
rect -1362 22742 -1358 22788
rect -1338 22742 -1334 22788
rect -1314 22742 -1310 22788
rect -1290 22742 -1286 22788
rect -1266 22742 -1262 22788
rect -1242 22742 -1238 22788
rect -1218 22742 -1214 22788
rect -1194 22742 -1190 22788
rect -1170 22742 -1166 22788
rect -1146 22742 -1142 22788
rect -1122 22742 -1118 22788
rect -1098 22742 -1094 22788
rect -1074 22742 -1070 22788
rect -1050 22742 -1046 22788
rect -1026 22742 -1022 22788
rect -1002 22742 -998 22788
rect -978 22742 -974 22788
rect -954 22742 -950 22788
rect -930 22742 -926 22788
rect -906 22742 -902 22788
rect -882 22742 -878 22788
rect -858 22742 -854 22788
rect -834 22742 -830 22788
rect -810 22742 -806 22788
rect -786 22742 -782 22788
rect -762 22742 -758 22788
rect -738 22742 -734 22788
rect -714 22742 -710 22788
rect -690 22742 -686 22788
rect -666 22742 -662 22788
rect -642 22742 -638 22788
rect -618 22742 -614 22788
rect -594 22742 -590 22788
rect -570 22742 -566 22788
rect -546 22742 -542 22788
rect -522 22742 -518 22788
rect -498 22742 -494 22788
rect -474 22742 -470 22788
rect -450 22742 -446 22788
rect -426 22742 -422 22788
rect -413 22781 -408 22788
rect -402 22781 -398 22788
rect -403 22767 -398 22781
rect -402 22742 -398 22767
rect -378 22742 -374 22836
rect -354 22742 -350 22836
rect -330 22742 -326 22836
rect -306 22742 -302 22836
rect -282 22742 -278 22836
rect -258 22742 -254 22836
rect -234 22742 -230 22836
rect -210 22742 -206 22836
rect -186 22742 -182 22836
rect -162 22742 -158 22836
rect -138 22742 -134 22836
rect -114 22742 -110 22836
rect -90 22742 -86 22836
rect -66 22742 -62 22836
rect -42 22742 -38 22836
rect -18 22742 -14 22836
rect 6 22742 10 22836
rect 30 22742 34 22836
rect 54 22742 58 22836
rect 78 22742 82 22836
rect 102 22742 106 22836
rect 126 22742 130 22836
rect 150 22742 154 22836
rect 174 22742 178 22836
rect 198 22742 202 22836
rect 222 22742 226 22836
rect 246 22742 250 22836
rect 270 22742 274 22836
rect 294 22742 298 22836
rect 318 22742 322 22836
rect 342 22742 346 22836
rect 366 22742 370 22836
rect 390 22742 394 22836
rect 414 22742 418 22836
rect 438 22742 442 22836
rect 462 22742 466 22836
rect 486 22742 490 22836
rect 510 22742 514 22836
rect 534 22742 538 22836
rect 558 22742 562 22836
rect 582 22742 586 22836
rect 606 22742 610 22836
rect 630 22742 634 22836
rect 654 22742 658 22836
rect 678 22742 682 22836
rect 702 22742 706 22836
rect 726 22742 730 22836
rect 750 22742 754 22836
rect 774 22742 778 22836
rect 798 22742 802 22836
rect 822 22742 826 22836
rect 846 22742 850 22836
rect 870 22742 874 22836
rect 894 22742 898 22836
rect 918 22742 922 22836
rect 942 22742 946 22836
rect 966 22742 970 22836
rect 990 22742 994 22836
rect 1014 22742 1018 22836
rect 1038 22742 1042 22836
rect 1062 22742 1066 22836
rect 1086 22742 1090 22836
rect 1099 22757 1104 22767
rect 1110 22757 1114 22836
rect 1109 22743 1114 22757
rect 1099 22742 1133 22743
rect -2393 22740 1133 22742
rect -2371 22718 -2366 22740
rect -2348 22718 -2343 22740
rect -2325 22718 -2320 22740
rect -2072 22738 -2036 22739
rect -2072 22732 -2054 22738
rect -2309 22724 -2301 22732
rect -2317 22718 -2309 22724
rect -2092 22723 -2062 22728
rect -2000 22719 -1992 22740
rect -1938 22739 -1906 22740
rect -1920 22738 -1906 22739
rect -1806 22732 -1680 22738
rect -1854 22723 -1806 22728
rect -1655 22724 -1647 22732
rect -1982 22719 -1966 22720
rect -2000 22718 -1966 22719
rect -1846 22718 -1806 22721
rect -1663 22718 -1655 22724
rect -1642 22718 -1637 22740
rect -1619 22718 -1614 22740
rect -1530 22718 -1526 22740
rect -1506 22718 -1502 22740
rect -1482 22718 -1478 22740
rect -1458 22718 -1454 22740
rect -1434 22718 -1430 22740
rect -1410 22718 -1406 22740
rect -1386 22718 -1382 22740
rect -1362 22718 -1358 22740
rect -1338 22718 -1334 22740
rect -1314 22718 -1310 22740
rect -1290 22718 -1286 22740
rect -1266 22718 -1262 22740
rect -1242 22718 -1238 22740
rect -1218 22718 -1214 22740
rect -1194 22718 -1190 22740
rect -1170 22718 -1166 22740
rect -1146 22718 -1142 22740
rect -1122 22718 -1118 22740
rect -1098 22718 -1094 22740
rect -1074 22718 -1070 22740
rect -1050 22718 -1046 22740
rect -1026 22718 -1022 22740
rect -1002 22718 -998 22740
rect -978 22718 -974 22740
rect -954 22718 -950 22740
rect -930 22718 -926 22740
rect -906 22718 -902 22740
rect -882 22718 -878 22740
rect -858 22718 -854 22740
rect -834 22718 -830 22740
rect -810 22718 -806 22740
rect -786 22718 -782 22740
rect -762 22718 -758 22740
rect -738 22718 -734 22740
rect -714 22718 -710 22740
rect -690 22718 -686 22740
rect -666 22718 -662 22740
rect -642 22718 -638 22740
rect -618 22718 -614 22740
rect -594 22718 -590 22740
rect -570 22718 -566 22740
rect -546 22718 -542 22740
rect -522 22718 -518 22740
rect -498 22718 -494 22740
rect -474 22718 -470 22740
rect -450 22718 -446 22740
rect -426 22718 -422 22740
rect -402 22718 -398 22740
rect -378 22718 -374 22740
rect -354 22718 -350 22740
rect -330 22718 -326 22740
rect -306 22718 -302 22740
rect -282 22718 -278 22740
rect -258 22718 -254 22740
rect -234 22718 -230 22740
rect -210 22718 -206 22740
rect -186 22718 -182 22740
rect -162 22718 -158 22740
rect -138 22718 -134 22740
rect -114 22718 -110 22740
rect -90 22718 -86 22740
rect -66 22718 -62 22740
rect -42 22718 -38 22740
rect -18 22718 -14 22740
rect 6 22718 10 22740
rect 30 22718 34 22740
rect 54 22718 58 22740
rect 78 22718 82 22740
rect 102 22718 106 22740
rect 126 22718 130 22740
rect 150 22718 154 22740
rect 174 22718 178 22740
rect 198 22718 202 22740
rect 222 22718 226 22740
rect 246 22718 250 22740
rect 270 22718 274 22740
rect 294 22718 298 22740
rect 318 22718 322 22740
rect 342 22718 346 22740
rect 366 22718 370 22740
rect 390 22718 394 22740
rect 414 22718 418 22740
rect 438 22718 442 22740
rect 462 22718 466 22740
rect 486 22718 490 22740
rect 510 22718 514 22740
rect 534 22718 538 22740
rect 558 22718 562 22740
rect 582 22718 586 22740
rect 606 22718 610 22740
rect 630 22718 634 22740
rect 654 22718 658 22740
rect 678 22718 682 22740
rect 702 22718 706 22740
rect 726 22718 730 22740
rect 750 22718 754 22740
rect 774 22718 778 22740
rect 798 22718 802 22740
rect 822 22718 826 22740
rect 846 22718 850 22740
rect 870 22718 874 22740
rect 894 22718 898 22740
rect 918 22718 922 22740
rect 942 22718 946 22740
rect 966 22718 970 22740
rect 990 22718 994 22740
rect 1014 22718 1018 22740
rect 1038 22718 1042 22740
rect 1062 22718 1066 22740
rect 1086 22718 1090 22740
rect 1099 22733 1104 22740
rect 1109 22719 1114 22733
rect 1110 22718 1114 22719
rect 1134 22718 1138 22836
rect 1158 22718 1162 22836
rect 1182 22718 1186 22836
rect 1206 22718 1210 22836
rect 1230 22718 1234 22836
rect 1254 22718 1258 22836
rect 1278 22718 1282 22836
rect 1302 22811 1306 22836
rect 1302 22787 1309 22811
rect 1302 22718 1306 22787
rect 1326 22718 1330 22836
rect 1350 22718 1354 22836
rect 1374 22718 1378 22836
rect 1398 22718 1402 22836
rect 1422 22718 1426 22836
rect 1446 22718 1450 22836
rect 1470 22718 1474 22836
rect 1494 22718 1498 22836
rect 1501 22835 1515 22836
rect 1518 22835 1525 22883
rect 1518 22718 1522 22835
rect 1542 22718 1546 23196
rect 1566 22718 1570 23196
rect 1590 22718 1594 23196
rect 1614 22718 1618 23196
rect 1638 22718 1642 23196
rect 1662 22718 1666 23196
rect 1686 22718 1690 23196
rect 1710 22718 1714 23196
rect 1734 22718 1738 23196
rect 1758 22718 1762 23196
rect 1782 22863 1786 23196
rect 1771 22862 1805 22863
rect 1806 22862 1810 23196
rect 1830 22862 1834 23196
rect 1854 22862 1858 23196
rect 1878 22862 1882 23196
rect 1902 22862 1906 23196
rect 1926 22862 1930 23196
rect 1950 22862 1954 23196
rect 1974 22862 1978 23196
rect 1998 22862 2002 23196
rect 2022 22862 2026 23196
rect 2046 22862 2050 23196
rect 2070 22862 2074 23196
rect 2094 22862 2098 23196
rect 2118 22862 2122 23196
rect 2142 22862 2146 23196
rect 2166 22862 2170 23196
rect 2190 22862 2194 23196
rect 2214 22862 2218 23196
rect 2238 22862 2242 23196
rect 2262 22862 2266 23196
rect 2286 22862 2290 23196
rect 2310 22862 2314 23196
rect 2334 22862 2338 23196
rect 2358 22862 2362 23196
rect 2382 22862 2386 23196
rect 2406 22862 2410 23196
rect 2430 22862 2434 23196
rect 2454 22862 2458 23196
rect 2478 22862 2482 23196
rect 2502 22862 2506 23196
rect 2515 23189 2520 23196
rect 2533 23195 2547 23196
rect 2525 23175 2530 23189
rect 2526 22862 2530 23175
rect 2539 23069 2544 23079
rect 2549 23055 2554 23069
rect 2550 22862 2554 23055
rect 2563 22949 2568 22959
rect 2573 22935 2578 22949
rect 2574 22862 2578 22935
rect 2587 22862 2595 22863
rect 1771 22860 2595 22862
rect 1771 22853 1776 22860
rect 1782 22853 1786 22860
rect 1781 22839 1786 22853
rect 1771 22829 1776 22839
rect 1781 22815 1786 22829
rect 1782 22718 1786 22815
rect 1806 22787 1810 22860
rect 1806 22766 1813 22787
rect 1830 22766 1834 22860
rect 1854 22766 1858 22860
rect 1878 22766 1882 22860
rect 1902 22766 1906 22860
rect 1926 22766 1930 22860
rect 1950 22766 1954 22860
rect 1974 22766 1978 22860
rect 1998 22766 2002 22860
rect 2022 22766 2026 22860
rect 2046 22766 2050 22860
rect 2070 22766 2074 22860
rect 2094 22766 2098 22860
rect 2118 22766 2122 22860
rect 2142 22766 2146 22860
rect 2166 22766 2170 22860
rect 2190 22766 2194 22860
rect 2214 22766 2218 22860
rect 2238 22766 2242 22860
rect 2262 22766 2266 22860
rect 2286 22766 2290 22860
rect 2310 22766 2314 22860
rect 2334 22766 2338 22860
rect 2358 22766 2362 22860
rect 2382 22766 2386 22860
rect 2406 22766 2410 22860
rect 2430 22766 2434 22860
rect 2454 22766 2458 22860
rect 2467 22781 2472 22791
rect 2478 22781 2482 22860
rect 2477 22767 2482 22781
rect 2502 22766 2506 22860
rect 2526 22766 2530 22860
rect 2550 22766 2554 22860
rect 2574 22766 2578 22860
rect 2581 22859 2595 22860
rect 2587 22853 2592 22859
rect 2597 22839 2602 22853
rect 2587 22805 2592 22815
rect 2598 22805 2602 22839
rect 2597 22791 2602 22805
rect 2587 22781 2592 22791
rect 2597 22767 2602 22781
rect 2611 22777 2619 22781
rect 2605 22767 2611 22777
rect 2598 22766 2602 22767
rect 2611 22766 2619 22767
rect 1789 22764 2619 22766
rect 1789 22763 1803 22764
rect 1806 22739 1813 22764
rect 1806 22718 1810 22739
rect 1830 22718 1834 22764
rect 1854 22718 1858 22764
rect 1878 22718 1882 22764
rect 1902 22718 1906 22764
rect 1926 22718 1930 22764
rect 1950 22718 1954 22764
rect 1974 22718 1978 22764
rect 1998 22718 2002 22764
rect 2022 22718 2026 22764
rect 2046 22718 2050 22764
rect 2070 22718 2074 22764
rect 2094 22718 2098 22764
rect 2118 22718 2122 22764
rect 2142 22718 2146 22764
rect 2166 22718 2170 22764
rect 2190 22718 2194 22764
rect 2214 22718 2218 22764
rect 2238 22718 2242 22764
rect 2262 22718 2266 22764
rect 2286 22718 2290 22764
rect 2310 22718 2314 22764
rect 2334 22718 2338 22764
rect 2358 22718 2362 22764
rect 2382 22718 2386 22764
rect 2406 22718 2410 22764
rect 2430 22718 2434 22764
rect 2454 22718 2458 22764
rect 2467 22733 2472 22743
rect 2477 22719 2482 22733
rect 2478 22718 2482 22719
rect 2502 22718 2506 22764
rect 2526 22718 2530 22764
rect 2550 22718 2554 22764
rect 2574 22718 2578 22764
rect 2598 22718 2602 22764
rect 2605 22763 2619 22764
rect 2611 22757 2616 22763
rect 2621 22743 2626 22757
rect 2622 22739 2626 22743
rect 2611 22718 2619 22719
rect -2393 22716 2619 22718
rect -2371 22694 -2366 22716
rect -2348 22694 -2343 22716
rect -2325 22694 -2320 22716
rect -2000 22714 -1966 22716
rect -2309 22696 -2301 22704
rect -2062 22703 -2054 22710
rect -2092 22696 -2084 22703
rect -2062 22696 -2026 22698
rect -2317 22694 -2309 22696
rect -2062 22694 -2012 22696
rect -2000 22694 -1992 22714
rect -1982 22713 -1966 22714
rect -1846 22712 -1806 22716
rect -1846 22705 -1798 22710
rect -1806 22703 -1798 22705
rect -1854 22701 -1846 22703
rect -1854 22696 -1806 22701
rect -1655 22696 -1647 22704
rect -1864 22694 -1796 22695
rect -1663 22694 -1655 22696
rect -1642 22694 -1637 22716
rect -1619 22694 -1614 22716
rect -1530 22694 -1526 22716
rect -1506 22694 -1502 22716
rect -1482 22694 -1478 22716
rect -1458 22694 -1454 22716
rect -1434 22694 -1430 22716
rect -1410 22694 -1406 22716
rect -1386 22694 -1382 22716
rect -1362 22694 -1358 22716
rect -1338 22694 -1334 22716
rect -1314 22694 -1310 22716
rect -1290 22694 -1286 22716
rect -1266 22694 -1262 22716
rect -1242 22694 -1238 22716
rect -1218 22694 -1214 22716
rect -1194 22694 -1190 22716
rect -1170 22694 -1166 22716
rect -1146 22694 -1142 22716
rect -1122 22694 -1118 22716
rect -1098 22694 -1094 22716
rect -1074 22694 -1070 22716
rect -1050 22694 -1046 22716
rect -1026 22694 -1022 22716
rect -1002 22694 -998 22716
rect -978 22694 -974 22716
rect -954 22694 -950 22716
rect -930 22694 -926 22716
rect -906 22694 -902 22716
rect -882 22694 -878 22716
rect -858 22694 -854 22716
rect -834 22694 -830 22716
rect -810 22694 -806 22716
rect -786 22694 -782 22716
rect -762 22694 -758 22716
rect -738 22694 -734 22716
rect -714 22694 -710 22716
rect -690 22694 -686 22716
rect -666 22694 -662 22716
rect -642 22694 -638 22716
rect -618 22694 -614 22716
rect -594 22694 -590 22716
rect -570 22694 -566 22716
rect -546 22694 -542 22716
rect -522 22694 -518 22716
rect -498 22694 -494 22716
rect -474 22694 -470 22716
rect -450 22694 -446 22716
rect -426 22694 -422 22716
rect -402 22694 -398 22716
rect -378 22715 -374 22716
rect -2393 22692 -381 22694
rect -2371 22646 -2366 22692
rect -2348 22646 -2343 22692
rect -2325 22646 -2320 22692
rect -2317 22688 -2309 22692
rect -2062 22688 -2054 22692
rect -2154 22684 -2138 22686
rect -2057 22684 -2054 22688
rect -2292 22678 -2054 22684
rect -2052 22678 -2044 22688
rect -2092 22662 -2062 22664
rect -2094 22658 -2062 22662
rect -2000 22646 -1992 22692
rect -1846 22685 -1806 22692
rect -1663 22688 -1655 22692
rect -1846 22678 -1680 22684
rect -1854 22662 -1806 22664
rect -1854 22658 -1680 22662
rect -1979 22646 -1945 22648
rect -1642 22646 -1637 22692
rect -1619 22646 -1614 22692
rect -1530 22646 -1526 22692
rect -1506 22646 -1502 22692
rect -1482 22646 -1478 22692
rect -1458 22646 -1454 22692
rect -1434 22646 -1430 22692
rect -1410 22646 -1406 22692
rect -1386 22646 -1382 22692
rect -1362 22646 -1358 22692
rect -1338 22646 -1334 22692
rect -1314 22646 -1310 22692
rect -1290 22646 -1286 22692
rect -1266 22646 -1262 22692
rect -1242 22646 -1238 22692
rect -1218 22646 -1214 22692
rect -1194 22646 -1190 22692
rect -1170 22646 -1166 22692
rect -1146 22646 -1142 22692
rect -1122 22646 -1118 22692
rect -1098 22646 -1094 22692
rect -1074 22646 -1070 22692
rect -1050 22646 -1046 22692
rect -1026 22646 -1022 22692
rect -1002 22646 -998 22692
rect -978 22646 -974 22692
rect -954 22646 -950 22692
rect -930 22646 -926 22692
rect -906 22646 -902 22692
rect -882 22646 -878 22692
rect -858 22646 -854 22692
rect -834 22646 -830 22692
rect -810 22646 -806 22692
rect -786 22646 -782 22692
rect -762 22646 -758 22692
rect -738 22646 -734 22692
rect -714 22646 -710 22692
rect -690 22646 -686 22692
rect -666 22646 -662 22692
rect -642 22646 -638 22692
rect -618 22646 -614 22692
rect -594 22646 -590 22692
rect -570 22646 -566 22692
rect -546 22646 -542 22692
rect -522 22646 -518 22692
rect -498 22646 -494 22692
rect -474 22646 -470 22692
rect -450 22646 -446 22692
rect -426 22646 -422 22692
rect -402 22646 -398 22692
rect -395 22691 -381 22692
rect -378 22691 -371 22715
rect -378 22646 -374 22691
rect -354 22646 -350 22716
rect -330 22646 -326 22716
rect -306 22646 -302 22716
rect -282 22646 -278 22716
rect -258 22646 -254 22716
rect -234 22646 -230 22716
rect -210 22646 -206 22716
rect -186 22646 -182 22716
rect -162 22646 -158 22716
rect -138 22646 -134 22716
rect -114 22646 -110 22716
rect -90 22646 -86 22716
rect -66 22646 -62 22716
rect -42 22646 -38 22716
rect -18 22646 -14 22716
rect 6 22646 10 22716
rect 30 22646 34 22716
rect 54 22646 58 22716
rect 78 22646 82 22716
rect 102 22646 106 22716
rect 126 22646 130 22716
rect 150 22646 154 22716
rect 174 22646 178 22716
rect 198 22646 202 22716
rect 222 22646 226 22716
rect 246 22646 250 22716
rect 270 22646 274 22716
rect 294 22646 298 22716
rect 318 22646 322 22716
rect 342 22646 346 22716
rect 366 22646 370 22716
rect 390 22646 394 22716
rect 414 22646 418 22716
rect 438 22646 442 22716
rect 462 22646 466 22716
rect 486 22646 490 22716
rect 510 22646 514 22716
rect 534 22646 538 22716
rect 558 22646 562 22716
rect 582 22646 586 22716
rect 606 22646 610 22716
rect 630 22646 634 22716
rect 654 22646 658 22716
rect 678 22646 682 22716
rect 702 22646 706 22716
rect 726 22646 730 22716
rect 750 22646 754 22716
rect 774 22646 778 22716
rect 798 22646 802 22716
rect 822 22646 826 22716
rect 846 22646 850 22716
rect 870 22646 874 22716
rect 894 22646 898 22716
rect 918 22646 922 22716
rect 942 22646 946 22716
rect 966 22646 970 22716
rect 990 22646 994 22716
rect 1014 22646 1018 22716
rect 1038 22646 1042 22716
rect 1062 22646 1066 22716
rect 1086 22646 1090 22716
rect 1110 22646 1114 22716
rect 1134 22691 1138 22716
rect -2393 22644 1131 22646
rect -2371 22598 -2366 22644
rect -2348 22598 -2343 22644
rect -2325 22598 -2320 22644
rect -2080 22643 -1906 22644
rect -2080 22642 -2036 22643
rect -2080 22636 -2054 22642
rect -2309 22628 -2301 22634
rect -2317 22618 -2309 22628
rect -2070 22627 -2040 22634
rect -2054 22619 -2040 22622
rect -2000 22617 -1992 22643
rect -1920 22642 -1906 22643
rect -1850 22636 -1846 22644
rect -1840 22636 -1792 22644
rect -1969 22624 -1966 22633
rect -1850 22629 -1802 22634
rect -1906 22627 -1802 22629
rect -1655 22628 -1647 22634
rect -1906 22626 -1850 22627
rect -1846 22619 -1802 22625
rect -1663 22618 -1655 22628
rect -1860 22617 -1798 22618
rect -2078 22610 -2070 22617
rect -2309 22600 -2301 22606
rect -2317 22598 -2309 22600
rect -2154 22598 -2145 22608
rect -2044 22607 -2040 22612
rect -2028 22610 -1945 22617
rect -1929 22610 -1794 22617
rect -2070 22600 -2040 22607
rect -2044 22598 -2028 22600
rect -2000 22598 -1992 22610
rect -1860 22609 -1798 22610
rect -1850 22600 -1802 22607
rect -1655 22600 -1647 22606
rect -1978 22598 -1942 22599
rect -1663 22598 -1655 22600
rect -1642 22598 -1637 22644
rect -1619 22598 -1614 22644
rect -1530 22598 -1526 22644
rect -1506 22598 -1502 22644
rect -1482 22598 -1478 22644
rect -1458 22598 -1454 22644
rect -1434 22598 -1430 22644
rect -1410 22598 -1406 22644
rect -1386 22598 -1382 22644
rect -1362 22598 -1358 22644
rect -1338 22598 -1334 22644
rect -1314 22598 -1310 22644
rect -1290 22598 -1286 22644
rect -1266 22598 -1262 22644
rect -1242 22598 -1238 22644
rect -1218 22598 -1214 22644
rect -1194 22598 -1190 22644
rect -1170 22598 -1166 22644
rect -1146 22598 -1142 22644
rect -1122 22598 -1118 22644
rect -1098 22598 -1094 22644
rect -1074 22598 -1070 22644
rect -1050 22598 -1046 22644
rect -1026 22598 -1022 22644
rect -1002 22598 -998 22644
rect -978 22598 -974 22644
rect -954 22598 -950 22644
rect -930 22598 -926 22644
rect -906 22598 -902 22644
rect -882 22598 -878 22644
rect -858 22598 -854 22644
rect -834 22598 -830 22644
rect -810 22598 -806 22644
rect -786 22598 -782 22644
rect -762 22598 -758 22644
rect -738 22598 -734 22644
rect -714 22598 -710 22644
rect -690 22598 -686 22644
rect -666 22598 -662 22644
rect -642 22598 -638 22644
rect -618 22598 -614 22644
rect -594 22598 -590 22644
rect -570 22598 -566 22644
rect -546 22598 -542 22644
rect -522 22598 -518 22644
rect -498 22598 -494 22644
rect -474 22598 -470 22644
rect -450 22598 -446 22644
rect -426 22598 -422 22644
rect -402 22598 -398 22644
rect -378 22598 -374 22644
rect -354 22598 -350 22644
rect -330 22598 -326 22644
rect -306 22598 -302 22644
rect -282 22598 -278 22644
rect -258 22598 -254 22644
rect -234 22598 -230 22644
rect -210 22598 -206 22644
rect -186 22598 -182 22644
rect -162 22598 -158 22644
rect -138 22598 -134 22644
rect -114 22598 -110 22644
rect -90 22598 -86 22644
rect -66 22598 -62 22644
rect -42 22598 -38 22644
rect -18 22598 -14 22644
rect 6 22598 10 22644
rect 30 22598 34 22644
rect 54 22598 58 22644
rect 78 22598 82 22644
rect 102 22598 106 22644
rect 126 22598 130 22644
rect 150 22598 154 22644
rect 174 22598 178 22644
rect 198 22598 202 22644
rect 222 22598 226 22644
rect 246 22598 250 22644
rect 270 22598 274 22644
rect 294 22599 298 22644
rect 283 22598 317 22599
rect -2393 22596 317 22598
rect -2371 22502 -2366 22596
rect -2348 22502 -2343 22596
rect -2325 22558 -2320 22596
rect -2317 22590 -2309 22596
rect -2145 22592 -2138 22596
rect -2070 22592 -2054 22596
rect -2078 22583 -2054 22590
rect -2062 22558 -2032 22559
rect -2000 22558 -1992 22596
rect -1846 22592 -1802 22596
rect -1846 22582 -1792 22591
rect -1663 22590 -1655 22596
rect -1942 22560 -1937 22572
rect -1850 22569 -1822 22570
rect -1850 22565 -1802 22569
rect -2325 22550 -2317 22558
rect -2062 22556 -1961 22558
rect -2325 22530 -2320 22550
rect -2317 22542 -2309 22550
rect -2062 22543 -2040 22554
rect -2032 22549 -1961 22556
rect -1947 22550 -1942 22558
rect -1842 22556 -1794 22559
rect -2070 22538 -2022 22542
rect -2325 22518 -2317 22530
rect -2325 22502 -2320 22518
rect -2317 22514 -2309 22518
rect -2309 22502 -2301 22514
rect -2068 22507 -2038 22514
rect -2000 22504 -1992 22549
rect -1942 22548 -1937 22550
rect -1932 22540 -1927 22548
rect -1912 22545 -1896 22551
rect -1842 22543 -1802 22554
rect -1671 22550 -1663 22558
rect -1663 22542 -1655 22550
rect -1850 22538 -1680 22542
rect -1937 22524 -1934 22526
rect -1926 22524 -1921 22529
rect -1926 22519 -1924 22524
rect -1916 22516 -1914 22519
rect -1842 22516 -1794 22525
rect -1671 22518 -1663 22530
rect -1924 22506 -1916 22515
rect -1663 22514 -1655 22518
rect -1852 22507 -1804 22514
rect -1916 22505 -1914 22506
rect -2025 22503 -1991 22504
rect -2025 22502 -1975 22503
rect -1842 22502 -1804 22505
rect -1655 22502 -1647 22514
rect -1642 22502 -1637 22596
rect -1619 22502 -1614 22596
rect -1530 22502 -1526 22596
rect -1517 22565 -1512 22575
rect -1506 22565 -1502 22596
rect -1507 22551 -1502 22565
rect -1506 22502 -1502 22551
rect -1482 22502 -1478 22596
rect -1458 22502 -1454 22596
rect -1434 22502 -1430 22596
rect -1410 22502 -1406 22596
rect -1386 22502 -1382 22596
rect -1362 22502 -1358 22596
rect -1338 22502 -1334 22596
rect -1314 22502 -1310 22596
rect -1290 22502 -1286 22596
rect -1266 22502 -1262 22596
rect -1242 22502 -1238 22596
rect -1218 22502 -1214 22596
rect -1194 22502 -1190 22596
rect -1170 22502 -1166 22596
rect -1146 22502 -1142 22596
rect -1122 22502 -1118 22596
rect -1098 22502 -1094 22596
rect -1074 22502 -1070 22596
rect -1050 22502 -1046 22596
rect -1026 22502 -1022 22596
rect -1002 22502 -998 22596
rect -978 22551 -974 22596
rect -989 22550 -955 22551
rect -954 22550 -950 22596
rect -930 22550 -926 22596
rect -906 22550 -902 22596
rect -882 22550 -878 22596
rect -858 22550 -854 22596
rect -834 22550 -830 22596
rect -810 22550 -806 22596
rect -786 22550 -782 22596
rect -762 22550 -758 22596
rect -738 22550 -734 22596
rect -714 22550 -710 22596
rect -690 22550 -686 22596
rect -666 22550 -662 22596
rect -642 22550 -638 22596
rect -618 22550 -614 22596
rect -594 22550 -590 22596
rect -570 22550 -566 22596
rect -546 22550 -542 22596
rect -522 22550 -518 22596
rect -498 22550 -494 22596
rect -474 22550 -470 22596
rect -450 22550 -446 22596
rect -426 22550 -422 22596
rect -402 22550 -398 22596
rect -378 22550 -374 22596
rect -354 22550 -350 22596
rect -330 22550 -326 22596
rect -306 22550 -302 22596
rect -282 22550 -278 22596
rect -258 22550 -254 22596
rect -234 22550 -230 22596
rect -210 22550 -206 22596
rect -186 22550 -182 22596
rect -162 22550 -158 22596
rect -138 22550 -134 22596
rect -114 22550 -110 22596
rect -90 22550 -86 22596
rect -66 22550 -62 22596
rect -42 22550 -38 22596
rect -18 22550 -14 22596
rect 6 22550 10 22596
rect 30 22550 34 22596
rect 54 22550 58 22596
rect 78 22550 82 22596
rect 102 22550 106 22596
rect 126 22550 130 22596
rect 150 22550 154 22596
rect 174 22550 178 22596
rect 198 22550 202 22596
rect 222 22550 226 22596
rect 246 22550 250 22596
rect 270 22550 274 22596
rect 283 22589 288 22596
rect 294 22589 298 22596
rect 293 22575 298 22589
rect 294 22550 298 22575
rect 318 22550 322 22644
rect 342 22550 346 22644
rect 366 22550 370 22644
rect 390 22550 394 22644
rect 414 22550 418 22644
rect 438 22550 442 22644
rect 462 22550 466 22644
rect 486 22550 490 22644
rect 510 22550 514 22644
rect 534 22550 538 22644
rect 558 22550 562 22644
rect 582 22550 586 22644
rect 606 22550 610 22644
rect 630 22550 634 22644
rect 654 22550 658 22644
rect 678 22550 682 22644
rect 702 22550 706 22644
rect 726 22550 730 22644
rect 750 22550 754 22644
rect 774 22550 778 22644
rect 798 22550 802 22644
rect 822 22550 826 22644
rect 846 22550 850 22644
rect 870 22550 874 22644
rect 894 22550 898 22644
rect 918 22550 922 22644
rect 942 22550 946 22644
rect 966 22550 970 22644
rect 990 22550 994 22644
rect 1014 22550 1018 22644
rect 1038 22550 1042 22644
rect 1062 22550 1066 22644
rect 1086 22550 1090 22644
rect 1110 22550 1114 22644
rect 1117 22643 1131 22644
rect 1134 22643 1141 22691
rect 1134 22550 1138 22643
rect 1158 22550 1162 22716
rect 1182 22550 1186 22716
rect 1206 22550 1210 22716
rect 1230 22550 1234 22716
rect 1254 22550 1258 22716
rect 1278 22550 1282 22716
rect 1302 22550 1306 22716
rect 1326 22671 1330 22716
rect 1315 22670 1349 22671
rect 1350 22670 1354 22716
rect 1374 22670 1378 22716
rect 1398 22670 1402 22716
rect 1422 22670 1426 22716
rect 1446 22670 1450 22716
rect 1470 22670 1474 22716
rect 1494 22670 1498 22716
rect 1518 22670 1522 22716
rect 1531 22685 1536 22695
rect 1542 22685 1546 22716
rect 1541 22671 1546 22685
rect 1542 22670 1546 22671
rect 1566 22670 1570 22716
rect 1590 22670 1594 22716
rect 1614 22670 1618 22716
rect 1638 22670 1642 22716
rect 1662 22670 1666 22716
rect 1686 22670 1690 22716
rect 1710 22670 1714 22716
rect 1734 22670 1738 22716
rect 1758 22670 1762 22716
rect 1782 22670 1786 22716
rect 1806 22670 1810 22716
rect 1830 22670 1834 22716
rect 1854 22670 1858 22716
rect 1878 22670 1882 22716
rect 1891 22685 1896 22695
rect 1902 22685 1906 22716
rect 1901 22671 1906 22685
rect 1926 22670 1930 22716
rect 1950 22670 1954 22716
rect 1974 22670 1978 22716
rect 1998 22670 2002 22716
rect 2022 22670 2026 22716
rect 2046 22670 2050 22716
rect 2070 22670 2074 22716
rect 2094 22670 2098 22716
rect 2118 22670 2122 22716
rect 2142 22670 2146 22716
rect 2166 22670 2170 22716
rect 2190 22670 2194 22716
rect 2214 22670 2218 22716
rect 2238 22670 2242 22716
rect 2262 22670 2266 22716
rect 2286 22670 2290 22716
rect 2310 22670 2314 22716
rect 2334 22670 2338 22716
rect 2358 22670 2362 22716
rect 2382 22670 2386 22716
rect 2406 22670 2410 22716
rect 2430 22670 2434 22716
rect 2454 22670 2458 22716
rect 2478 22670 2482 22716
rect 2502 22715 2506 22716
rect 2502 22694 2509 22715
rect 2526 22694 2530 22716
rect 2550 22694 2554 22716
rect 2574 22694 2578 22716
rect 2598 22694 2602 22716
rect 2605 22715 2619 22716
rect 2622 22709 2629 22739
rect 2659 22733 2664 22743
rect 2669 22719 2674 22733
rect 2621 22695 2629 22709
rect 2611 22694 2619 22695
rect 2485 22692 2619 22694
rect 2485 22691 2499 22692
rect 2502 22691 2509 22692
rect 2526 22670 2530 22692
rect 2550 22670 2554 22692
rect 2574 22670 2578 22692
rect 2598 22670 2602 22692
rect 2605 22691 2619 22692
rect 2611 22685 2616 22691
rect 2621 22671 2626 22685
rect 2635 22681 2643 22685
rect 2629 22671 2635 22681
rect 2622 22670 2626 22671
rect 1315 22668 2643 22670
rect 1315 22661 1320 22668
rect 1326 22661 1330 22668
rect 1325 22647 1330 22661
rect 1315 22637 1320 22647
rect 1325 22623 1330 22637
rect 1350 22623 1354 22668
rect 1326 22550 1330 22623
rect 1339 22622 1373 22623
rect 1374 22622 1378 22668
rect 1398 22622 1402 22668
rect 1422 22622 1426 22668
rect 1446 22622 1450 22668
rect 1470 22622 1474 22668
rect 1494 22622 1498 22668
rect 1518 22622 1522 22668
rect 1542 22622 1546 22668
rect 1566 22622 1570 22668
rect 1590 22622 1594 22668
rect 1614 22622 1618 22668
rect 1638 22622 1642 22668
rect 1662 22622 1666 22668
rect 1686 22622 1690 22668
rect 1710 22622 1714 22668
rect 1734 22622 1738 22668
rect 1758 22622 1762 22668
rect 1782 22622 1786 22668
rect 1806 22622 1810 22668
rect 1830 22622 1834 22668
rect 1854 22622 1858 22668
rect 1878 22622 1882 22668
rect 1891 22637 1896 22647
rect 1901 22623 1906 22637
rect 1902 22622 1906 22623
rect 1926 22622 1930 22668
rect 1950 22622 1954 22668
rect 1974 22622 1978 22668
rect 1998 22622 2002 22668
rect 2022 22622 2026 22668
rect 2046 22622 2050 22668
rect 2070 22622 2074 22668
rect 2094 22622 2098 22668
rect 2118 22622 2122 22668
rect 2142 22622 2146 22668
rect 2166 22622 2170 22668
rect 2190 22622 2194 22668
rect 2214 22622 2218 22668
rect 2238 22622 2242 22668
rect 2262 22622 2266 22668
rect 2286 22622 2290 22668
rect 2310 22622 2314 22668
rect 2334 22622 2338 22668
rect 2358 22622 2362 22668
rect 2382 22622 2386 22668
rect 2406 22622 2410 22668
rect 2430 22622 2434 22668
rect 2454 22622 2458 22668
rect 2478 22622 2482 22668
rect 2502 22646 2509 22667
rect 2526 22646 2530 22668
rect 2550 22646 2554 22668
rect 2574 22646 2578 22668
rect 2598 22646 2602 22668
rect 2622 22646 2626 22668
rect 2629 22667 2643 22668
rect 2646 22667 2653 22691
rect 2646 22646 2650 22667
rect 2659 22661 2664 22671
rect 2669 22647 2674 22661
rect 2683 22657 2691 22661
rect 2677 22647 2683 22657
rect 2670 22646 2674 22647
rect 2683 22646 2717 22647
rect 2485 22644 2717 22646
rect 2485 22643 2499 22644
rect 2502 22643 2509 22644
rect 2502 22622 2506 22643
rect 2526 22622 2530 22644
rect 2550 22622 2554 22644
rect 2574 22622 2578 22644
rect 2598 22622 2602 22644
rect 2622 22622 2626 22644
rect 2646 22643 2650 22644
rect 1339 22620 2643 22622
rect 1339 22613 1344 22620
rect 1350 22613 1354 22620
rect 1349 22599 1354 22613
rect 1339 22598 1373 22599
rect 1374 22598 1378 22620
rect 1398 22598 1402 22620
rect 1422 22598 1426 22620
rect 1446 22598 1450 22620
rect 1470 22598 1474 22620
rect 1494 22598 1498 22620
rect 1518 22598 1522 22620
rect 1542 22598 1546 22620
rect 1566 22619 1570 22620
rect 1339 22596 1563 22598
rect 1339 22589 1344 22596
rect 1349 22575 1357 22589
rect 1374 22575 1378 22596
rect -989 22548 1347 22550
rect -989 22541 -984 22548
rect -978 22541 -974 22548
rect -979 22527 -974 22541
rect -989 22517 -984 22527
rect -979 22503 -974 22517
rect -978 22502 -974 22503
rect -954 22502 -950 22548
rect -930 22502 -926 22548
rect -906 22502 -902 22548
rect -882 22502 -878 22548
rect -858 22502 -854 22548
rect -834 22502 -830 22548
rect -810 22502 -806 22548
rect -786 22502 -782 22548
rect -762 22502 -758 22548
rect -738 22502 -734 22548
rect -714 22502 -710 22548
rect -690 22502 -686 22548
rect -666 22502 -662 22548
rect -642 22502 -638 22548
rect -618 22502 -614 22548
rect -594 22502 -590 22548
rect -570 22502 -566 22548
rect -546 22503 -542 22548
rect -557 22502 -523 22503
rect -2393 22500 -523 22502
rect -2371 22478 -2366 22500
rect -2348 22478 -2343 22500
rect -2325 22490 -2317 22500
rect -2076 22490 -2068 22497
rect -2062 22490 -2001 22497
rect -2325 22478 -2320 22490
rect -2317 22486 -2309 22490
rect -2015 22489 -2001 22490
rect -2309 22478 -2301 22486
rect -2068 22480 -2062 22487
rect -2000 22482 -1992 22500
rect -1974 22498 -1960 22500
rect -1842 22499 -1804 22500
rect -1862 22497 -1794 22498
rect -1985 22495 -1794 22497
rect -1985 22490 -1852 22495
rect -1842 22489 -1794 22495
rect -1671 22490 -1663 22500
rect -2015 22480 -1985 22482
rect -1852 22480 -1804 22487
rect -1663 22486 -1655 22490
rect -2000 22478 -1992 22480
rect -1976 22478 -1940 22479
rect -1655 22478 -1647 22486
rect -1642 22478 -1637 22500
rect -1619 22478 -1614 22500
rect -1530 22478 -1526 22500
rect -1506 22478 -1502 22500
rect -1482 22499 -1478 22500
rect -2393 22476 -1485 22478
rect -2371 22382 -2366 22476
rect -2348 22382 -2343 22476
rect -2325 22474 -2320 22476
rect -2309 22474 -2301 22476
rect -2325 22462 -2317 22474
rect -2062 22463 -2032 22470
rect -2325 22442 -2320 22462
rect -2317 22458 -2309 22462
rect -2325 22434 -2317 22442
rect -2060 22436 -2030 22439
rect -2325 22382 -2320 22434
rect -2317 22426 -2309 22434
rect -2060 22423 -2038 22434
rect -2033 22427 -2030 22436
rect -2028 22432 -2027 22436
rect -2068 22418 -2038 22421
rect -2309 22386 -2301 22394
rect -2317 22382 -2309 22386
rect -2000 22382 -1992 22476
rect -1888 22471 -1874 22476
rect -1842 22472 -1804 22476
rect -1655 22474 -1647 22476
rect -1902 22469 -1874 22471
rect -1842 22462 -1794 22471
rect -1671 22462 -1663 22474
rect -1663 22458 -1655 22462
rect -1912 22451 -1884 22453
rect -1852 22445 -1804 22449
rect -1844 22436 -1796 22439
rect -1671 22434 -1663 22442
rect -1844 22423 -1804 22434
rect -1663 22426 -1655 22434
rect -1852 22418 -1680 22422
rect -1655 22386 -1647 22394
rect -1663 22382 -1655 22386
rect -1642 22382 -1637 22476
rect -1619 22382 -1614 22476
rect -1530 22382 -1526 22476
rect -1506 22382 -1502 22476
rect -1499 22475 -1485 22476
rect -1482 22475 -1475 22499
rect -1482 22382 -1478 22475
rect -1458 22382 -1454 22500
rect -1434 22382 -1430 22500
rect -1410 22382 -1406 22500
rect -1386 22382 -1382 22500
rect -1362 22382 -1358 22500
rect -1338 22382 -1334 22500
rect -1314 22382 -1310 22500
rect -1290 22382 -1286 22500
rect -1266 22382 -1262 22500
rect -1242 22382 -1238 22500
rect -1218 22382 -1214 22500
rect -1194 22382 -1190 22500
rect -1170 22382 -1166 22500
rect -1157 22469 -1152 22479
rect -1146 22469 -1142 22500
rect -1147 22455 -1142 22469
rect -1146 22382 -1142 22455
rect -1122 22403 -1118 22500
rect -2393 22380 -2020 22382
rect -2012 22380 -1125 22382
rect -2371 22286 -2366 22380
rect -2348 22286 -2343 22380
rect -2325 22318 -2320 22380
rect -2317 22378 -2309 22380
rect -2062 22367 -2061 22368
rect -2060 22367 -2049 22380
rect -2309 22358 -2301 22366
rect -2068 22360 -2061 22367
rect -2020 22360 -2012 22372
rect -2317 22350 -2309 22358
rect -2124 22351 -2108 22353
rect -2060 22351 -2049 22360
rect -2020 22358 -2004 22360
rect -2000 22358 -1992 22380
rect -1972 22378 -1958 22380
rect -1663 22378 -1655 22380
rect -1958 22377 -1942 22378
rect -1980 22360 -1932 22367
rect -1655 22358 -1647 22366
rect -2292 22350 -2049 22351
rect -2036 22350 -2030 22358
rect -2020 22356 -1992 22358
rect -2292 22343 -2030 22350
rect -2292 22342 -2049 22343
rect -2031 22342 -2030 22343
rect -2026 22342 -2020 22348
rect -2325 22310 -2317 22318
rect -2325 22290 -2320 22310
rect -2317 22302 -2309 22310
rect -2325 22286 -2317 22290
rect -2000 22286 -1992 22356
rect -1844 22342 -1680 22351
rect -1663 22350 -1655 22358
rect -1671 22310 -1663 22318
rect -1663 22302 -1655 22310
rect -1926 22286 -1892 22289
rect -1671 22286 -1663 22290
rect -1642 22286 -1637 22380
rect -1619 22286 -1614 22380
rect -1530 22286 -1526 22380
rect -1506 22286 -1502 22380
rect -1482 22286 -1478 22380
rect -1458 22286 -1454 22380
rect -1434 22286 -1430 22380
rect -1410 22286 -1406 22380
rect -1386 22286 -1382 22380
rect -1362 22286 -1358 22380
rect -1338 22286 -1334 22380
rect -1314 22286 -1310 22380
rect -1290 22286 -1286 22380
rect -1266 22286 -1262 22380
rect -1242 22286 -1238 22380
rect -1218 22286 -1214 22380
rect -1194 22286 -1190 22380
rect -1170 22286 -1166 22380
rect -1146 22286 -1142 22380
rect -1139 22379 -1125 22380
rect -1122 22379 -1115 22403
rect -1122 22286 -1118 22379
rect -1098 22286 -1094 22500
rect -1074 22286 -1070 22500
rect -1050 22286 -1046 22500
rect -1026 22286 -1022 22500
rect -1002 22286 -998 22500
rect -978 22286 -974 22500
rect -954 22475 -950 22500
rect -954 22454 -947 22475
rect -930 22454 -926 22500
rect -906 22454 -902 22500
rect -882 22454 -878 22500
rect -858 22454 -854 22500
rect -834 22454 -830 22500
rect -810 22454 -806 22500
rect -786 22454 -782 22500
rect -762 22454 -758 22500
rect -738 22454 -734 22500
rect -714 22454 -710 22500
rect -690 22454 -686 22500
rect -666 22454 -662 22500
rect -642 22454 -638 22500
rect -618 22454 -614 22500
rect -594 22454 -590 22500
rect -570 22454 -566 22500
rect -557 22493 -552 22500
rect -546 22493 -542 22500
rect -547 22479 -542 22493
rect -546 22454 -542 22479
rect -522 22454 -518 22548
rect -498 22454 -494 22548
rect -474 22454 -470 22548
rect -450 22454 -446 22548
rect -426 22454 -422 22548
rect -402 22454 -398 22548
rect -378 22454 -374 22548
rect -354 22454 -350 22548
rect -330 22454 -326 22548
rect -306 22454 -302 22548
rect -282 22454 -278 22548
rect -258 22454 -254 22548
rect -234 22454 -230 22548
rect -210 22454 -206 22548
rect -186 22454 -182 22548
rect -162 22454 -158 22548
rect -138 22454 -134 22548
rect -114 22454 -110 22548
rect -90 22454 -86 22548
rect -66 22454 -62 22548
rect -42 22454 -38 22548
rect -18 22454 -14 22548
rect 6 22454 10 22548
rect 30 22454 34 22548
rect 54 22454 58 22548
rect 78 22454 82 22548
rect 102 22454 106 22548
rect 126 22454 130 22548
rect 150 22454 154 22548
rect 174 22454 178 22548
rect 198 22454 202 22548
rect 222 22454 226 22548
rect 246 22454 250 22548
rect 270 22454 274 22548
rect 294 22454 298 22548
rect 318 22523 322 22548
rect 318 22499 325 22523
rect 318 22454 322 22499
rect 342 22454 346 22548
rect 366 22454 370 22548
rect 390 22454 394 22548
rect 414 22454 418 22548
rect 438 22454 442 22548
rect 462 22454 466 22548
rect 486 22454 490 22548
rect 510 22454 514 22548
rect 534 22454 538 22548
rect 558 22454 562 22548
rect 582 22454 586 22548
rect 606 22454 610 22548
rect 630 22454 634 22548
rect 654 22454 658 22548
rect 678 22454 682 22548
rect 702 22454 706 22548
rect 726 22454 730 22548
rect 750 22454 754 22548
rect 774 22454 778 22548
rect 798 22454 802 22548
rect 822 22454 826 22548
rect 846 22454 850 22548
rect 870 22454 874 22548
rect 894 22454 898 22548
rect 918 22454 922 22548
rect 942 22454 946 22548
rect 966 22454 970 22548
rect 990 22454 994 22548
rect 1014 22454 1018 22548
rect 1038 22454 1042 22548
rect 1062 22454 1066 22548
rect 1086 22454 1090 22548
rect 1110 22454 1114 22548
rect 1134 22454 1138 22548
rect 1158 22454 1162 22548
rect 1182 22454 1186 22548
rect 1206 22454 1210 22548
rect 1230 22454 1234 22548
rect 1254 22454 1258 22548
rect 1278 22454 1282 22548
rect 1302 22454 1306 22548
rect 1326 22454 1330 22548
rect 1333 22547 1347 22548
rect 1350 22547 1357 22575
rect 1363 22574 1397 22575
rect 1398 22574 1402 22596
rect 1422 22574 1426 22596
rect 1446 22574 1450 22596
rect 1470 22574 1474 22596
rect 1494 22574 1498 22596
rect 1518 22574 1522 22596
rect 1542 22574 1546 22596
rect 1549 22595 1563 22596
rect 1566 22595 1573 22619
rect 1566 22574 1570 22595
rect 1590 22574 1594 22620
rect 1614 22574 1618 22620
rect 1638 22574 1642 22620
rect 1662 22574 1666 22620
rect 1686 22574 1690 22620
rect 1710 22574 1714 22620
rect 1734 22574 1738 22620
rect 1758 22574 1762 22620
rect 1782 22574 1786 22620
rect 1806 22574 1810 22620
rect 1830 22574 1834 22620
rect 1854 22574 1858 22620
rect 1878 22574 1882 22620
rect 1902 22574 1906 22620
rect 1926 22619 1930 22620
rect 1926 22598 1933 22619
rect 1950 22598 1954 22620
rect 1974 22598 1978 22620
rect 1998 22598 2002 22620
rect 2022 22598 2026 22620
rect 2046 22598 2050 22620
rect 2070 22598 2074 22620
rect 2094 22598 2098 22620
rect 2118 22598 2122 22620
rect 2142 22598 2146 22620
rect 2166 22598 2170 22620
rect 2190 22598 2194 22620
rect 2214 22598 2218 22620
rect 2238 22598 2242 22620
rect 2262 22598 2266 22620
rect 2286 22598 2290 22620
rect 2310 22598 2314 22620
rect 2334 22598 2338 22620
rect 2358 22598 2362 22620
rect 2382 22598 2386 22620
rect 2406 22598 2410 22620
rect 2430 22598 2434 22620
rect 2454 22598 2458 22620
rect 2478 22598 2482 22620
rect 2502 22598 2506 22620
rect 2526 22598 2530 22620
rect 2550 22598 2554 22620
rect 2574 22598 2578 22620
rect 2598 22598 2602 22620
rect 2622 22598 2626 22620
rect 2629 22619 2643 22620
rect 1909 22596 2643 22598
rect 1909 22595 1923 22596
rect 1926 22595 1933 22596
rect 1950 22574 1954 22596
rect 1974 22574 1978 22596
rect 1998 22574 2002 22596
rect 2022 22574 2026 22596
rect 2046 22574 2050 22596
rect 2070 22574 2074 22596
rect 2094 22574 2098 22596
rect 2118 22574 2122 22596
rect 2142 22574 2146 22596
rect 2166 22574 2170 22596
rect 2190 22574 2194 22596
rect 2214 22574 2218 22596
rect 2238 22574 2242 22596
rect 2262 22574 2266 22596
rect 2286 22574 2290 22596
rect 2310 22574 2314 22596
rect 2334 22574 2338 22596
rect 2358 22574 2362 22596
rect 2382 22574 2386 22596
rect 2406 22574 2410 22596
rect 2430 22574 2434 22596
rect 2454 22574 2458 22596
rect 2478 22574 2482 22596
rect 2502 22574 2506 22596
rect 2526 22574 2530 22596
rect 2550 22574 2554 22596
rect 2574 22574 2578 22596
rect 2598 22574 2602 22596
rect 2622 22574 2626 22596
rect 2629 22595 2643 22596
rect 2646 22595 2653 22643
rect 2646 22574 2650 22595
rect 2670 22574 2674 22644
rect 2677 22643 2691 22644
rect 3139 22637 3144 22647
rect 3859 22637 3864 22647
rect 3149 22623 3154 22637
rect 3869 22623 3874 22637
rect 1363 22572 2691 22574
rect 1363 22565 1368 22572
rect 1374 22565 1378 22572
rect 1373 22551 1378 22565
rect 1350 22454 1354 22547
rect 1363 22526 1397 22527
rect 1398 22526 1402 22572
rect 1422 22526 1426 22572
rect 1446 22526 1450 22572
rect 1470 22526 1474 22572
rect 1494 22526 1498 22572
rect 1518 22526 1522 22572
rect 1542 22526 1546 22572
rect 1566 22526 1570 22572
rect 1590 22526 1594 22572
rect 1614 22526 1618 22572
rect 1638 22526 1642 22572
rect 1662 22526 1666 22572
rect 1686 22526 1690 22572
rect 1710 22526 1714 22572
rect 1734 22526 1738 22572
rect 1758 22526 1762 22572
rect 1782 22526 1786 22572
rect 1806 22526 1810 22572
rect 1830 22526 1834 22572
rect 1854 22526 1858 22572
rect 1878 22526 1882 22572
rect 1902 22526 1906 22572
rect 1926 22550 1933 22571
rect 1950 22550 1954 22572
rect 1974 22550 1978 22572
rect 1998 22550 2002 22572
rect 2022 22550 2026 22572
rect 2046 22550 2050 22572
rect 2070 22550 2074 22572
rect 2094 22550 2098 22572
rect 2118 22550 2122 22572
rect 2142 22550 2146 22572
rect 2166 22550 2170 22572
rect 2190 22550 2194 22572
rect 2214 22550 2218 22572
rect 2238 22550 2242 22572
rect 2262 22550 2266 22572
rect 2286 22550 2290 22572
rect 2310 22550 2314 22572
rect 2334 22550 2338 22572
rect 2358 22550 2362 22572
rect 2382 22550 2386 22572
rect 2406 22550 2410 22572
rect 2430 22550 2434 22572
rect 2454 22550 2458 22572
rect 2478 22550 2482 22572
rect 2502 22550 2506 22572
rect 2526 22550 2530 22572
rect 2550 22550 2554 22572
rect 2574 22550 2578 22572
rect 2598 22550 2602 22572
rect 2622 22550 2626 22572
rect 2646 22550 2650 22572
rect 2670 22550 2674 22572
rect 2677 22571 2691 22572
rect 2694 22571 2701 22595
rect 3139 22589 3144 22599
rect 3859 22589 3864 22599
rect 3149 22575 3154 22589
rect 3869 22575 3874 22589
rect 2694 22550 2698 22571
rect 2717 22558 2725 22565
rect 2717 22552 2719 22558
rect 2717 22551 2725 22552
rect 1909 22548 2715 22550
rect 2755 22548 2789 22551
rect 1909 22547 1923 22548
rect 1926 22547 1933 22548
rect 1926 22526 1930 22547
rect 1950 22526 1954 22548
rect 1974 22526 1978 22548
rect 1998 22526 2002 22548
rect 2022 22526 2026 22548
rect 2046 22526 2050 22548
rect 2070 22526 2074 22548
rect 2094 22526 2098 22548
rect 2118 22526 2122 22548
rect 2142 22526 2146 22548
rect 2166 22526 2170 22548
rect 2190 22526 2194 22548
rect 2214 22526 2218 22548
rect 2238 22526 2242 22548
rect 2262 22526 2266 22548
rect 2286 22526 2290 22548
rect 2310 22526 2314 22548
rect 2334 22526 2338 22548
rect 2358 22526 2362 22548
rect 2382 22526 2386 22548
rect 2406 22527 2410 22548
rect 2395 22526 2429 22527
rect 1363 22524 2429 22526
rect 1363 22523 1371 22524
rect 1373 22503 1381 22517
rect 1374 22499 1381 22503
rect 1398 22499 1402 22524
rect 1374 22454 1378 22499
rect 1398 22475 1405 22499
rect 1387 22454 1421 22455
rect -971 22452 1421 22454
rect -971 22451 -957 22452
rect -954 22427 -947 22452
rect -954 22286 -950 22427
rect -930 22286 -926 22452
rect -906 22286 -902 22452
rect -882 22286 -878 22452
rect -858 22286 -854 22452
rect -834 22286 -830 22452
rect -810 22286 -806 22452
rect -786 22286 -782 22452
rect -762 22286 -758 22452
rect -738 22286 -734 22452
rect -714 22286 -710 22452
rect -690 22286 -686 22452
rect -666 22286 -662 22452
rect -642 22286 -638 22452
rect -618 22286 -614 22452
rect -594 22286 -590 22452
rect -570 22286 -566 22452
rect -546 22286 -542 22452
rect -522 22427 -518 22452
rect -522 22403 -515 22427
rect -522 22286 -518 22403
rect -498 22286 -494 22452
rect -474 22286 -470 22452
rect -450 22286 -446 22452
rect -426 22286 -422 22452
rect -402 22286 -398 22452
rect -378 22286 -374 22452
rect -354 22286 -350 22452
rect -330 22286 -326 22452
rect -306 22286 -302 22452
rect -282 22286 -278 22452
rect -258 22286 -254 22452
rect -234 22286 -230 22452
rect -210 22286 -206 22452
rect -186 22286 -182 22452
rect -162 22286 -158 22452
rect -138 22286 -134 22452
rect -114 22286 -110 22452
rect -90 22286 -86 22452
rect -66 22286 -62 22452
rect -42 22286 -38 22452
rect -18 22286 -14 22452
rect 6 22286 10 22452
rect 30 22286 34 22452
rect 54 22286 58 22452
rect 78 22286 82 22452
rect 91 22397 96 22407
rect 102 22397 106 22452
rect 101 22383 106 22397
rect 91 22373 96 22383
rect 101 22359 106 22373
rect 102 22286 106 22359
rect 126 22331 130 22452
rect -2393 22284 123 22286
rect -2371 22238 -2366 22284
rect -2348 22238 -2343 22284
rect -2325 22278 -2317 22284
rect -2053 22282 -1972 22284
rect -2325 22262 -2320 22278
rect -2317 22274 -2309 22278
rect -2069 22274 -2068 22275
rect -2309 22262 -2301 22274
rect -2069 22267 -2038 22274
rect -2069 22265 -2068 22267
rect -2000 22266 -1992 22282
rect -1926 22279 -1924 22284
rect -1916 22276 -1914 22279
rect -1671 22278 -1663 22284
rect -1982 22266 -1916 22275
rect -1663 22274 -1655 22278
rect -2325 22250 -2317 22262
rect -2068 22259 -2053 22265
rect -2027 22264 -1992 22266
rect -2076 22250 -2053 22257
rect -2011 22256 -2002 22264
rect -2000 22256 -1992 22264
rect -1655 22262 -1647 22274
rect -2003 22254 -1992 22256
rect -2325 22238 -2320 22250
rect -2317 22246 -2309 22250
rect -2309 22238 -2301 22246
rect -2015 22242 -2003 22254
rect -2000 22238 -1992 22254
rect -1972 22250 -1924 22257
rect -1862 22249 -1680 22258
rect -1671 22250 -1663 22262
rect -1663 22246 -1655 22250
rect -1976 22238 -1940 22239
rect -1655 22238 -1647 22246
rect -1642 22238 -1637 22284
rect -1619 22238 -1614 22284
rect -1530 22238 -1526 22284
rect -1506 22238 -1502 22284
rect -1482 22238 -1478 22284
rect -1458 22238 -1454 22284
rect -1434 22238 -1430 22284
rect -1410 22238 -1406 22284
rect -1386 22238 -1382 22284
rect -1362 22238 -1358 22284
rect -1338 22238 -1334 22284
rect -1314 22238 -1310 22284
rect -1290 22238 -1286 22284
rect -1266 22238 -1262 22284
rect -1242 22238 -1238 22284
rect -1218 22238 -1214 22284
rect -1194 22238 -1190 22284
rect -1170 22238 -1166 22284
rect -1146 22238 -1142 22284
rect -1122 22238 -1118 22284
rect -1098 22238 -1094 22284
rect -1074 22238 -1070 22284
rect -1050 22238 -1046 22284
rect -1026 22238 -1022 22284
rect -1002 22238 -998 22284
rect -978 22238 -974 22284
rect -954 22238 -950 22284
rect -930 22238 -926 22284
rect -906 22238 -902 22284
rect -882 22238 -878 22284
rect -858 22238 -854 22284
rect -834 22238 -830 22284
rect -810 22238 -806 22284
rect -786 22238 -782 22284
rect -762 22238 -758 22284
rect -738 22238 -734 22284
rect -714 22238 -710 22284
rect -690 22238 -686 22284
rect -666 22238 -662 22284
rect -642 22238 -638 22284
rect -618 22238 -614 22284
rect -594 22238 -590 22284
rect -570 22238 -566 22284
rect -546 22238 -542 22284
rect -522 22238 -518 22284
rect -498 22238 -494 22284
rect -474 22238 -470 22284
rect -450 22238 -446 22284
rect -426 22238 -422 22284
rect -402 22238 -398 22284
rect -378 22238 -374 22284
rect -354 22238 -350 22284
rect -330 22238 -326 22284
rect -306 22238 -302 22284
rect -282 22238 -278 22284
rect -258 22238 -254 22284
rect -234 22238 -230 22284
rect -210 22238 -206 22284
rect -186 22238 -182 22284
rect -162 22238 -158 22284
rect -138 22238 -134 22284
rect -114 22238 -110 22284
rect -90 22238 -86 22284
rect -66 22238 -62 22284
rect -42 22238 -38 22284
rect -18 22238 -14 22284
rect 6 22238 10 22284
rect 30 22238 34 22284
rect 54 22238 58 22284
rect 78 22238 82 22284
rect 102 22238 106 22284
rect 109 22283 123 22284
rect 126 22283 133 22331
rect 126 22238 130 22283
rect 150 22238 154 22452
rect 174 22238 178 22452
rect 198 22238 202 22452
rect 222 22238 226 22452
rect 246 22238 250 22452
rect 270 22238 274 22452
rect 294 22238 298 22452
rect 318 22238 322 22452
rect 342 22238 346 22452
rect 366 22238 370 22452
rect 390 22238 394 22452
rect 414 22238 418 22452
rect 438 22238 442 22452
rect 462 22238 466 22452
rect 486 22238 490 22452
rect 510 22238 514 22452
rect 534 22238 538 22452
rect 558 22238 562 22452
rect 582 22238 586 22452
rect 606 22238 610 22452
rect 630 22238 634 22452
rect 654 22238 658 22452
rect 678 22238 682 22452
rect 702 22238 706 22452
rect 726 22238 730 22452
rect 750 22238 754 22452
rect 774 22238 778 22452
rect 798 22238 802 22452
rect 822 22238 826 22452
rect 846 22238 850 22452
rect 870 22239 874 22452
rect 894 22239 898 22452
rect 859 22238 917 22239
rect 918 22238 922 22452
rect 931 22253 936 22263
rect 942 22253 946 22452
rect 941 22239 946 22253
rect 942 22238 946 22239
rect 966 22238 970 22452
rect 990 22238 994 22452
rect 1014 22238 1018 22452
rect 1038 22238 1042 22452
rect 1062 22238 1066 22452
rect 1086 22238 1090 22452
rect 1110 22238 1114 22452
rect 1134 22238 1138 22452
rect 1158 22238 1162 22452
rect 1182 22238 1186 22452
rect 1206 22238 1210 22452
rect 1230 22238 1234 22452
rect 1254 22238 1258 22452
rect 1278 22238 1282 22452
rect 1302 22238 1306 22452
rect 1315 22253 1320 22263
rect 1326 22253 1330 22452
rect 1325 22239 1330 22253
rect 1350 22238 1354 22452
rect 1374 22238 1378 22452
rect 1398 22445 1405 22451
rect 1397 22431 1405 22445
rect 1398 22427 1405 22431
rect 1398 22311 1402 22427
rect 1422 22379 1426 22524
rect 1422 22355 1429 22379
rect 1387 22310 1421 22311
rect 1422 22310 1426 22355
rect 1446 22310 1450 22524
rect 1470 22310 1474 22524
rect 1494 22310 1498 22524
rect 1518 22310 1522 22524
rect 1542 22310 1546 22524
rect 1566 22310 1570 22524
rect 1590 22310 1594 22524
rect 1614 22310 1618 22524
rect 1638 22310 1642 22524
rect 1662 22310 1666 22524
rect 1686 22310 1690 22524
rect 1710 22310 1714 22524
rect 1734 22310 1738 22524
rect 1758 22310 1762 22524
rect 1782 22310 1786 22524
rect 1806 22310 1810 22524
rect 1819 22325 1824 22335
rect 1830 22325 1834 22524
rect 1829 22311 1834 22325
rect 1854 22310 1858 22524
rect 1878 22310 1882 22524
rect 1902 22310 1906 22524
rect 1926 22310 1930 22524
rect 1950 22312 1954 22524
rect 1963 22349 1968 22359
rect 1974 22349 1978 22524
rect 1973 22335 1978 22349
rect 1963 22325 1968 22335
rect 1973 22322 1978 22325
rect 1973 22311 1978 22312
rect 1998 22310 2002 22524
rect 2022 22310 2026 22524
rect 2046 22310 2050 22524
rect 2070 22310 2074 22524
rect 2094 22310 2098 22524
rect 2118 22310 2122 22524
rect 2131 22373 2136 22383
rect 2142 22373 2146 22524
rect 2141 22359 2146 22373
rect 2166 22310 2170 22524
rect 2190 22408 2194 22524
rect 2214 22455 2218 22524
rect 2203 22454 2237 22455
rect 2238 22454 2242 22524
rect 2262 22454 2266 22524
rect 2286 22454 2290 22524
rect 2310 22454 2314 22524
rect 2334 22456 2338 22524
rect 2358 22503 2362 22524
rect 2347 22502 2381 22503
rect 2382 22502 2386 22524
rect 2395 22517 2400 22524
rect 2406 22517 2410 22524
rect 2405 22503 2410 22517
rect 2430 22502 2434 22548
rect 2454 22527 2458 22548
rect 2443 22526 2477 22527
rect 2478 22526 2482 22548
rect 2502 22526 2506 22548
rect 2526 22526 2530 22548
rect 2550 22526 2554 22548
rect 2574 22526 2578 22548
rect 2598 22526 2602 22548
rect 2622 22526 2626 22548
rect 2646 22526 2650 22548
rect 2670 22526 2674 22548
rect 2694 22526 2698 22548
rect 2701 22547 2715 22548
rect 3126 22547 3133 22571
rect 3846 22547 3853 22571
rect 7219 22565 7224 22575
rect 7229 22551 7234 22565
rect 7219 22541 7224 22551
rect 7229 22527 7234 22541
rect 2443 22524 2715 22526
rect 2443 22517 2448 22524
rect 2454 22517 2458 22524
rect 2453 22503 2458 22517
rect 2478 22502 2482 22524
rect 2502 22502 2506 22524
rect 2526 22502 2530 22524
rect 2550 22502 2554 22524
rect 2574 22502 2578 22524
rect 2598 22502 2602 22524
rect 2622 22502 2626 22524
rect 2646 22502 2650 22524
rect 2670 22502 2674 22524
rect 2694 22502 2698 22524
rect 2701 22523 2715 22524
rect 2742 22510 2749 22523
rect 2347 22500 2739 22502
rect 2803 22500 2837 22503
rect 2347 22493 2352 22500
rect 2358 22493 2362 22500
rect 2357 22479 2362 22493
rect 2347 22478 2381 22479
rect 2382 22478 2386 22500
rect 2430 22478 2434 22500
rect 2478 22478 2482 22500
rect 2502 22478 2506 22500
rect 2526 22478 2530 22500
rect 2550 22478 2554 22500
rect 2574 22478 2578 22500
rect 2598 22478 2602 22500
rect 2622 22478 2626 22500
rect 2646 22478 2650 22500
rect 2670 22478 2674 22500
rect 2694 22478 2698 22500
rect 2725 22499 2739 22500
rect 2742 22486 2749 22500
rect 3126 22499 3133 22523
rect 3846 22499 3853 22523
rect 7219 22517 7224 22527
rect 10579 22517 10584 22527
rect 7229 22503 7234 22517
rect 10589 22503 10594 22517
rect 2347 22476 2739 22478
rect 2347 22469 2352 22476
rect 2357 22466 2362 22469
rect 2357 22455 2362 22456
rect 2382 22454 2386 22476
rect 2430 22454 2434 22476
rect 2478 22454 2482 22476
rect 2502 22454 2506 22476
rect 2526 22454 2530 22476
rect 2550 22454 2554 22476
rect 2574 22454 2578 22476
rect 2598 22454 2602 22476
rect 2622 22454 2626 22476
rect 2646 22454 2650 22476
rect 2670 22454 2674 22476
rect 2694 22454 2698 22476
rect 2725 22475 2739 22476
rect 2742 22475 2749 22476
rect 2766 22454 2770 22496
rect 7195 22489 7203 22493
rect 7189 22479 7195 22489
rect 2203 22452 2787 22454
rect 2203 22445 2208 22452
rect 2214 22445 2218 22452
rect 2213 22431 2218 22445
rect 2203 22430 2237 22431
rect 2238 22430 2242 22452
rect 2262 22430 2266 22452
rect 2286 22430 2290 22452
rect 2310 22430 2314 22452
rect 2382 22430 2386 22452
rect 2430 22451 2434 22452
rect 2478 22451 2482 22452
rect 2203 22428 2427 22430
rect 2203 22421 2208 22428
rect 2213 22418 2218 22421
rect 2213 22407 2218 22408
rect 2238 22379 2242 22428
rect 2238 22358 2245 22379
rect 2262 22358 2266 22428
rect 2286 22358 2290 22428
rect 2310 22358 2314 22428
rect 2382 22427 2386 22428
rect 2413 22427 2427 22428
rect 2430 22427 2437 22451
rect 2478 22430 2485 22451
rect 2502 22430 2506 22452
rect 2526 22430 2530 22452
rect 2550 22430 2554 22452
rect 2574 22430 2578 22452
rect 2598 22430 2602 22452
rect 2622 22430 2626 22452
rect 2646 22430 2650 22452
rect 2670 22430 2674 22452
rect 2694 22430 2698 22452
rect 2766 22430 2770 22452
rect 2773 22451 2787 22452
rect 2790 22451 2797 22475
rect 3139 22469 3144 22479
rect 3859 22469 3864 22479
rect 4579 22469 4584 22479
rect 4819 22469 4824 22479
rect 6979 22476 7013 22479
rect 7189 22475 7203 22476
rect 7206 22475 7213 22499
rect 7219 22493 7224 22503
rect 10579 22493 10584 22503
rect 7229 22479 7234 22493
rect 7243 22489 7251 22493
rect 7237 22479 7243 22489
rect 10589 22479 10594 22493
rect 3149 22455 3154 22469
rect 3869 22455 3874 22469
rect 4589 22455 4594 22469
rect 4829 22455 4834 22469
rect 6907 22452 6912 22455
rect 2790 22430 2794 22451
rect 2461 22428 2811 22430
rect 2461 22427 2475 22428
rect 2478 22427 2485 22428
rect 2382 22406 2389 22427
rect 2502 22406 2506 22428
rect 2526 22406 2530 22428
rect 2550 22406 2554 22428
rect 2574 22406 2578 22428
rect 2598 22406 2602 22428
rect 2622 22406 2626 22428
rect 2646 22406 2650 22428
rect 2670 22406 2674 22428
rect 2694 22406 2698 22428
rect 2766 22406 2770 22428
rect 2790 22406 2794 22428
rect 2797 22427 2811 22428
rect 2814 22427 2821 22451
rect 6859 22438 6864 22441
rect 6894 22428 6898 22452
rect 7189 22451 7203 22452
rect 7237 22451 7251 22452
rect 10555 22441 10563 22445
rect 10549 22431 10555 22441
rect 6907 22428 6936 22431
rect 10531 22430 10565 22431
rect 10566 22430 10573 22451
rect 10579 22445 10584 22455
rect 10589 22431 10594 22445
rect 10603 22441 10611 22445
rect 10597 22431 10603 22441
rect 10579 22430 10613 22431
rect 10531 22428 10613 22430
rect 2814 22406 2818 22427
rect 2365 22404 2835 22406
rect 2365 22403 2379 22404
rect 2382 22382 2389 22404
rect 2502 22382 2506 22404
rect 2526 22382 2530 22404
rect 2550 22382 2554 22404
rect 2574 22382 2578 22404
rect 2598 22382 2602 22404
rect 2622 22382 2626 22404
rect 2646 22382 2650 22404
rect 2670 22382 2674 22404
rect 2694 22382 2698 22404
rect 2766 22382 2770 22404
rect 2790 22382 2794 22404
rect 2814 22382 2818 22404
rect 2821 22403 2835 22404
rect 2838 22403 2845 22427
rect 6835 22404 6864 22407
rect 6870 22404 6874 22428
rect 6894 22406 6901 22427
rect 6907 22421 6912 22428
rect 7189 22427 7203 22428
rect 7237 22427 7251 22428
rect 10549 22427 10563 22428
rect 6917 22407 6922 22421
rect 6931 22417 6939 22421
rect 10555 22417 10563 22421
rect 6925 22407 6931 22417
rect 10549 22407 10555 22417
rect 6907 22406 6941 22407
rect 6877 22404 6941 22406
rect 6979 22404 7013 22407
rect 7027 22404 7061 22407
rect 10531 22406 10565 22407
rect 10566 22406 10573 22428
rect 10579 22421 10584 22428
rect 10597 22427 10611 22428
rect 10589 22407 10594 22421
rect 10603 22417 10611 22421
rect 10597 22407 10603 22417
rect 10579 22406 10613 22407
rect 10531 22404 10613 22406
rect 2838 22382 2842 22403
rect 2365 22380 2859 22382
rect 2365 22379 2379 22380
rect 2382 22379 2389 22380
rect 2502 22358 2506 22380
rect 2526 22358 2530 22380
rect 2550 22358 2554 22380
rect 2574 22358 2578 22380
rect 2598 22358 2602 22380
rect 2622 22358 2626 22380
rect 2646 22358 2650 22380
rect 2670 22358 2674 22380
rect 2694 22358 2698 22380
rect 2766 22358 2770 22380
rect 2790 22358 2794 22380
rect 2814 22358 2818 22380
rect 2838 22358 2842 22380
rect 2845 22379 2859 22380
rect 2862 22379 2869 22403
rect 3019 22380 3053 22383
rect 3126 22379 3133 22403
rect 3846 22379 3853 22403
rect 4566 22379 4573 22403
rect 4806 22379 4813 22403
rect 6764 22394 6768 22404
rect 6877 22403 6891 22404
rect 6894 22403 6901 22404
rect 6733 22379 6747 22380
rect 2862 22358 2866 22379
rect 2910 22366 2917 22379
rect 6774 22370 6778 22394
rect 6859 22393 6867 22397
rect 6853 22383 6859 22393
rect 6835 22382 6869 22383
rect 6870 22382 6877 22403
rect 6894 22382 6898 22403
rect 6907 22397 6912 22404
rect 6925 22403 6939 22404
rect 6979 22397 6984 22404
rect 7189 22403 7203 22404
rect 7237 22403 7251 22404
rect 10549 22403 10563 22404
rect 10566 22403 10573 22404
rect 6917 22383 6922 22397
rect 6989 22394 6994 22397
rect 7003 22393 7011 22397
rect 6989 22383 6994 22384
rect 6997 22383 7003 22393
rect 7014 22390 7021 22403
rect 10579 22397 10584 22404
rect 10597 22403 10611 22404
rect 12019 22397 12024 22407
rect 10589 22383 10594 22397
rect 12029 22383 12034 22397
rect 6907 22382 6941 22383
rect 6835 22380 6941 22382
rect 6979 22380 7013 22383
rect 7027 22380 7061 22383
rect 6788 22379 6795 22380
rect 6853 22379 6867 22380
rect 6784 22366 6792 22370
rect 6859 22369 6867 22373
rect 6853 22359 6859 22369
rect 2221 22356 2907 22358
rect 2221 22355 2235 22356
rect 2238 22334 2245 22356
rect 2262 22334 2266 22356
rect 2286 22334 2290 22356
rect 2310 22334 2314 22356
rect 2502 22334 2506 22356
rect 2526 22334 2530 22356
rect 2550 22334 2554 22356
rect 2574 22334 2578 22356
rect 2598 22334 2602 22356
rect 2622 22334 2626 22356
rect 2646 22334 2650 22356
rect 2670 22334 2674 22356
rect 2694 22334 2698 22356
rect 2766 22334 2770 22356
rect 2790 22334 2794 22356
rect 2814 22334 2818 22356
rect 2838 22334 2842 22356
rect 2862 22334 2866 22356
rect 2893 22355 2907 22356
rect 2910 22355 2917 22356
rect 2221 22332 2955 22334
rect 2221 22331 2235 22332
rect 2238 22331 2245 22332
rect 2262 22310 2266 22332
rect 2286 22310 2290 22332
rect 2310 22310 2314 22332
rect 2502 22310 2506 22332
rect 2526 22310 2530 22332
rect 2550 22310 2554 22332
rect 2574 22310 2578 22332
rect 2598 22310 2602 22332
rect 2622 22310 2626 22332
rect 2646 22310 2650 22332
rect 2670 22310 2674 22332
rect 2694 22310 2698 22332
rect 2766 22310 2770 22332
rect 2790 22310 2794 22332
rect 2814 22310 2818 22332
rect 2838 22310 2842 22332
rect 2862 22310 2866 22332
rect 2941 22331 2955 22332
rect 3006 22310 3010 22352
rect 6740 22346 6744 22356
rect 6798 22346 6802 22356
rect 6688 22342 6696 22346
rect 6750 22332 6754 22346
rect 6808 22342 6816 22346
rect 6787 22332 6792 22335
rect 6870 22334 6877 22380
rect 6894 22334 6898 22380
rect 6907 22373 6912 22380
rect 6979 22373 6984 22380
rect 6997 22379 7011 22380
rect 7014 22379 7021 22380
rect 6917 22359 6922 22373
rect 6931 22369 6939 22373
rect 6989 22370 6994 22373
rect 10555 22369 10563 22373
rect 6925 22359 6931 22369
rect 7003 22366 7008 22369
rect 6989 22359 6994 22360
rect 10549 22359 10555 22369
rect 6979 22356 6984 22359
rect 7027 22356 7061 22359
rect 10531 22358 10565 22359
rect 10566 22358 10573 22379
rect 10579 22373 10584 22383
rect 12019 22373 12024 22383
rect 12499 22373 12504 22383
rect 12739 22373 12744 22383
rect 10589 22359 10594 22373
rect 10603 22369 10611 22373
rect 10597 22359 10603 22369
rect 12029 22359 12034 22373
rect 12509 22359 12514 22373
rect 12749 22359 12754 22373
rect 10579 22358 10613 22359
rect 10531 22356 10613 22358
rect 6908 22346 6912 22356
rect 6925 22355 6939 22356
rect 6918 22335 6922 22346
rect 6907 22334 6941 22335
rect 6853 22332 6941 22334
rect 6979 22332 7008 22335
rect 7014 22332 7018 22356
rect 10549 22355 10563 22356
rect 10555 22345 10563 22349
rect 10549 22335 10555 22345
rect 7027 22332 7061 22335
rect 10531 22334 10565 22335
rect 10566 22334 10573 22356
rect 10579 22349 10584 22356
rect 10597 22355 10611 22356
rect 12019 22349 12024 22359
rect 12499 22349 12504 22359
rect 12739 22349 12744 22359
rect 10589 22335 10594 22349
rect 10603 22345 10611 22349
rect 10597 22335 10603 22345
rect 12029 22335 12034 22349
rect 12509 22335 12514 22349
rect 12749 22335 12754 22349
rect 10579 22334 10613 22335
rect 10531 22332 10613 22334
rect 1387 22308 3027 22310
rect 1387 22301 1392 22308
rect 1398 22301 1402 22308
rect 1397 22287 1402 22301
rect 1422 22238 1426 22308
rect 1446 22238 1450 22308
rect 1470 22238 1474 22308
rect 1494 22238 1498 22308
rect 1518 22238 1522 22308
rect 1542 22238 1546 22308
rect 1566 22238 1570 22308
rect 1590 22238 1594 22308
rect 1614 22238 1618 22308
rect 1638 22238 1642 22308
rect 1662 22238 1666 22308
rect 1686 22238 1690 22308
rect 1710 22238 1714 22308
rect 1734 22238 1738 22308
rect 1758 22238 1762 22308
rect 1782 22238 1786 22308
rect 1806 22238 1810 22308
rect 1854 22259 1858 22308
rect -2393 22236 1851 22238
rect -2371 22166 -2366 22236
rect -2348 22166 -2343 22236
rect -2325 22234 -2320 22236
rect -2309 22234 -2301 22236
rect -2325 22222 -2317 22234
rect -2325 22202 -2320 22222
rect -2317 22218 -2309 22222
rect -2325 22194 -2317 22202
rect -2060 22196 -2030 22199
rect -2325 22174 -2320 22194
rect -2317 22186 -2309 22194
rect -2060 22183 -2038 22194
rect -2033 22187 -2030 22196
rect -2028 22192 -2027 22196
rect -2068 22178 -2038 22181
rect -2325 22166 -2317 22174
rect -2000 22166 -1992 22236
rect -1655 22234 -1647 22236
rect -1671 22222 -1663 22234
rect -1663 22218 -1655 22222
rect -1912 22211 -1884 22213
rect -1852 22205 -1804 22209
rect -1844 22196 -1796 22199
rect -1671 22194 -1663 22202
rect -1844 22183 -1804 22194
rect -1663 22186 -1655 22194
rect -1852 22178 -1680 22182
rect -1926 22166 -1892 22169
rect -1671 22166 -1663 22174
rect -1642 22166 -1637 22236
rect -1619 22166 -1614 22236
rect -1530 22166 -1526 22236
rect -1506 22166 -1502 22236
rect -1482 22166 -1478 22236
rect -1458 22166 -1454 22236
rect -1434 22166 -1430 22236
rect -1410 22166 -1406 22236
rect -1386 22166 -1382 22236
rect -1362 22166 -1358 22236
rect -1338 22166 -1334 22236
rect -1314 22166 -1310 22236
rect -1290 22166 -1286 22236
rect -1266 22166 -1262 22236
rect -1242 22166 -1238 22236
rect -1218 22166 -1214 22236
rect -1194 22166 -1190 22236
rect -1170 22166 -1166 22236
rect -1146 22166 -1142 22236
rect -1122 22166 -1118 22236
rect -1098 22166 -1094 22236
rect -1074 22166 -1070 22236
rect -1050 22166 -1046 22236
rect -1026 22166 -1022 22236
rect -1002 22166 -998 22236
rect -978 22166 -974 22236
rect -954 22166 -950 22236
rect -930 22166 -926 22236
rect -906 22166 -902 22236
rect -882 22166 -878 22236
rect -858 22166 -854 22236
rect -834 22166 -830 22236
rect -810 22166 -806 22236
rect -786 22166 -782 22236
rect -762 22166 -758 22236
rect -738 22166 -734 22236
rect -714 22166 -710 22236
rect -690 22166 -686 22236
rect -666 22166 -662 22236
rect -642 22166 -638 22236
rect -618 22166 -614 22236
rect -594 22166 -590 22236
rect -570 22166 -566 22236
rect -546 22166 -542 22236
rect -522 22166 -518 22236
rect -498 22166 -494 22236
rect -474 22166 -470 22236
rect -450 22166 -446 22236
rect -426 22166 -422 22236
rect -402 22166 -398 22236
rect -378 22166 -374 22236
rect -354 22166 -350 22236
rect -330 22166 -326 22236
rect -306 22166 -302 22236
rect -282 22166 -278 22236
rect -258 22166 -254 22236
rect -234 22166 -230 22236
rect -210 22166 -206 22236
rect -186 22166 -182 22236
rect -162 22166 -158 22236
rect -138 22166 -134 22236
rect -114 22166 -110 22236
rect -90 22166 -86 22236
rect -66 22166 -62 22236
rect -42 22166 -38 22236
rect -18 22166 -14 22236
rect 6 22166 10 22236
rect 30 22166 34 22236
rect 54 22166 58 22236
rect 78 22166 82 22236
rect 102 22166 106 22236
rect 126 22166 130 22236
rect 150 22166 154 22236
rect 174 22166 178 22236
rect 198 22166 202 22236
rect 222 22166 226 22236
rect 246 22166 250 22236
rect 270 22166 274 22236
rect 294 22166 298 22236
rect 318 22166 322 22236
rect 342 22166 346 22236
rect 366 22166 370 22236
rect 390 22166 394 22236
rect 414 22191 418 22236
rect 403 22190 437 22191
rect 438 22190 442 22236
rect 462 22190 466 22236
rect 486 22190 490 22236
rect 499 22205 504 22215
rect 510 22205 514 22236
rect 509 22191 514 22205
rect 534 22190 538 22236
rect 558 22190 562 22236
rect 582 22190 586 22236
rect 606 22190 610 22236
rect 630 22190 634 22236
rect 654 22190 658 22236
rect 678 22190 682 22236
rect 702 22190 706 22236
rect 726 22190 730 22236
rect 750 22190 754 22236
rect 774 22190 778 22236
rect 798 22190 802 22236
rect 822 22190 826 22236
rect 846 22190 850 22236
rect 859 22229 864 22236
rect 870 22229 874 22236
rect 883 22229 888 22236
rect 894 22229 898 22236
rect 869 22215 874 22229
rect 893 22215 898 22229
rect 918 22190 922 22236
rect 942 22190 946 22236
rect 966 22190 970 22236
rect 990 22190 994 22236
rect 1014 22190 1018 22236
rect 1038 22190 1042 22236
rect 1062 22190 1066 22236
rect 1086 22190 1090 22236
rect 1110 22190 1114 22236
rect 1134 22190 1138 22236
rect 1158 22190 1162 22236
rect 1182 22190 1186 22236
rect 1206 22190 1210 22236
rect 1230 22190 1234 22236
rect 1254 22190 1258 22236
rect 1278 22190 1282 22236
rect 1302 22190 1306 22236
rect 1350 22190 1354 22236
rect 1374 22190 1378 22236
rect 1422 22235 1426 22236
rect 1422 22214 1429 22235
rect 1446 22214 1450 22236
rect 1470 22214 1474 22236
rect 1494 22214 1498 22236
rect 1518 22214 1522 22236
rect 1542 22214 1546 22236
rect 1566 22214 1570 22236
rect 1590 22214 1594 22236
rect 1614 22214 1618 22236
rect 1638 22214 1642 22236
rect 1662 22214 1666 22236
rect 1686 22214 1690 22236
rect 1710 22214 1714 22236
rect 1734 22214 1738 22236
rect 1758 22214 1762 22236
rect 1782 22214 1786 22236
rect 1806 22214 1810 22236
rect 1837 22235 1851 22236
rect 1854 22235 1861 22259
rect 1878 22214 1882 22308
rect 1902 22214 1906 22308
rect 1926 22214 1930 22308
rect 1998 22283 2002 22308
rect 1998 22262 2005 22283
rect 2022 22262 2026 22308
rect 2046 22262 2050 22308
rect 2070 22262 2074 22308
rect 2094 22262 2098 22308
rect 2118 22262 2122 22308
rect 2166 22307 2170 22308
rect 2166 22286 2173 22307
rect 2262 22286 2266 22308
rect 2286 22286 2290 22308
rect 2310 22286 2314 22308
rect 2502 22286 2506 22308
rect 2526 22286 2530 22308
rect 2550 22286 2554 22308
rect 2574 22286 2578 22308
rect 2598 22286 2602 22308
rect 2622 22286 2626 22308
rect 2646 22286 2650 22308
rect 2670 22286 2674 22308
rect 2694 22286 2698 22308
rect 2707 22286 2741 22287
rect 2149 22284 2741 22286
rect 2149 22283 2163 22284
rect 2166 22283 2173 22284
rect 2262 22262 2266 22284
rect 2286 22262 2290 22284
rect 2310 22262 2314 22284
rect 2502 22262 2506 22284
rect 2526 22262 2530 22284
rect 2550 22262 2554 22284
rect 2574 22262 2578 22284
rect 2598 22262 2602 22284
rect 2622 22262 2626 22284
rect 2646 22262 2650 22284
rect 2670 22262 2674 22284
rect 2694 22262 2698 22284
rect 2707 22277 2712 22284
rect 2717 22263 2722 22277
rect 2718 22262 2722 22263
rect 2766 22262 2770 22308
rect 2790 22262 2794 22308
rect 2814 22287 2818 22308
rect 2803 22286 2837 22287
rect 2838 22286 2842 22308
rect 2862 22286 2866 22308
rect 3006 22286 3010 22308
rect 3013 22307 3027 22308
rect 3030 22307 3037 22331
rect 6702 22322 6706 22332
rect 6764 22322 6768 22332
rect 6712 22318 6720 22322
rect 3030 22286 3034 22307
rect 2803 22284 3051 22286
rect 2803 22277 2808 22284
rect 2814 22277 2818 22284
rect 2813 22263 2818 22277
rect 2838 22262 2842 22284
rect 2862 22262 2866 22284
rect 3006 22262 3010 22284
rect 3030 22262 3034 22284
rect 3037 22283 3051 22284
rect 3054 22283 3061 22307
rect 3139 22301 3144 22311
rect 6774 22308 6778 22322
rect 6787 22308 6816 22311
rect 6822 22308 6826 22332
rect 6853 22331 6867 22332
rect 6870 22310 6877 22332
rect 6894 22310 6898 22332
rect 6907 22325 6912 22332
rect 6918 22325 6922 22332
rect 6925 22331 6939 22332
rect 6917 22311 6922 22325
rect 6931 22321 6939 22325
rect 6925 22311 6931 22321
rect 6942 22318 6949 22322
rect 7003 22321 7011 22325
rect 6997 22311 7003 22321
rect 7014 22310 7021 22331
rect 7027 22325 7032 22332
rect 10549 22331 10563 22332
rect 7037 22311 7042 22325
rect 7051 22321 7059 22325
rect 10555 22321 10563 22325
rect 7045 22311 7051 22321
rect 10549 22311 10555 22321
rect 7027 22310 7061 22311
rect 6853 22308 6939 22310
rect 6997 22308 7061 22310
rect 10531 22310 10565 22311
rect 10566 22310 10573 22332
rect 10579 22325 10584 22332
rect 10597 22331 10611 22332
rect 10589 22311 10594 22325
rect 10603 22321 10611 22325
rect 11995 22321 12003 22325
rect 10597 22311 10603 22321
rect 11989 22311 11995 22321
rect 10579 22310 10613 22311
rect 10531 22308 10613 22310
rect 11971 22310 12005 22311
rect 12006 22310 12013 22331
rect 12019 22325 12024 22335
rect 12499 22325 12504 22335
rect 12739 22325 12744 22335
rect 12029 22311 12034 22325
rect 12043 22321 12051 22325
rect 12037 22311 12043 22321
rect 12509 22311 12514 22325
rect 12749 22311 12754 22325
rect 12019 22310 12053 22311
rect 11971 22308 12053 22310
rect 3149 22287 3154 22301
rect 6726 22298 6730 22308
rect 6787 22301 6792 22308
rect 6853 22307 6867 22308
rect 6736 22294 6744 22298
rect 6797 22287 6802 22301
rect 3054 22262 3058 22283
rect 1981 22260 3075 22262
rect 1981 22259 1995 22260
rect 1998 22238 2005 22260
rect 2022 22238 2026 22260
rect 2046 22238 2050 22260
rect 2070 22238 2074 22260
rect 2094 22238 2098 22260
rect 2118 22238 2122 22260
rect 2262 22238 2266 22260
rect 2286 22238 2290 22260
rect 2310 22238 2314 22260
rect 2502 22238 2506 22260
rect 2526 22238 2530 22260
rect 2550 22238 2554 22260
rect 2574 22238 2578 22260
rect 2598 22238 2602 22260
rect 2622 22238 2626 22260
rect 2646 22238 2650 22260
rect 2670 22238 2674 22260
rect 2694 22238 2698 22260
rect 2718 22238 2722 22260
rect 2766 22238 2770 22260
rect 2790 22238 2794 22260
rect 2838 22238 2842 22260
rect 2862 22238 2866 22260
rect 3006 22238 3010 22260
rect 3030 22238 3034 22260
rect 3054 22238 3058 22260
rect 3061 22259 3075 22260
rect 3078 22259 3085 22283
rect 3078 22238 3082 22259
rect 1981 22236 3099 22238
rect 1981 22235 1995 22236
rect 1998 22235 2005 22236
rect 2022 22214 2026 22236
rect 2046 22214 2050 22236
rect 2070 22214 2074 22236
rect 2094 22214 2098 22236
rect 2118 22214 2122 22236
rect 2262 22214 2266 22236
rect 2286 22214 2290 22236
rect 2310 22214 2314 22236
rect 2502 22214 2506 22236
rect 2526 22214 2530 22236
rect 2550 22214 2554 22236
rect 2574 22214 2578 22236
rect 2598 22214 2602 22236
rect 2622 22214 2626 22236
rect 2646 22214 2650 22236
rect 2670 22214 2674 22236
rect 2694 22214 2698 22236
rect 2718 22214 2722 22236
rect 2766 22214 2770 22236
rect 2790 22214 2794 22236
rect 2838 22215 2842 22236
rect 2803 22214 2861 22215
rect 2862 22214 2866 22236
rect 3006 22214 3010 22236
rect 3030 22214 3034 22236
rect 3054 22214 3058 22236
rect 3078 22214 3082 22236
rect 3085 22235 3099 22236
rect 3150 22214 3154 22287
rect 6715 22277 6720 22287
rect 6787 22284 6792 22287
rect 6798 22284 6802 22287
rect 6835 22284 6840 22287
rect 6853 22286 6869 22287
rect 6870 22286 6877 22308
rect 6894 22286 6898 22308
rect 6925 22307 6939 22308
rect 6942 22294 6949 22308
rect 6997 22307 7011 22308
rect 7014 22286 7021 22308
rect 7027 22301 7032 22308
rect 7045 22307 7059 22308
rect 10549 22307 10563 22308
rect 7037 22287 7042 22301
rect 7051 22297 7059 22301
rect 10555 22297 10563 22301
rect 7045 22287 7051 22297
rect 10549 22287 10555 22297
rect 7027 22286 7061 22287
rect 6853 22284 6939 22286
rect 6997 22284 7061 22286
rect 10531 22286 10565 22287
rect 10566 22286 10573 22308
rect 10579 22301 10584 22308
rect 10597 22307 10611 22308
rect 11989 22307 12003 22308
rect 10589 22287 10594 22301
rect 10603 22297 10611 22301
rect 11995 22297 12003 22301
rect 10597 22287 10603 22297
rect 11989 22287 11995 22297
rect 10579 22286 10613 22287
rect 10531 22284 10613 22286
rect 11971 22286 12005 22287
rect 12006 22286 12013 22308
rect 12019 22301 12024 22308
rect 12037 22307 12051 22308
rect 12029 22287 12034 22301
rect 12043 22297 12051 22301
rect 12475 22297 12483 22301
rect 12037 22287 12043 22297
rect 12469 22287 12475 22297
rect 12019 22286 12053 22287
rect 11971 22284 12053 22286
rect 12451 22286 12485 22287
rect 12486 22286 12493 22307
rect 12499 22301 12504 22311
rect 12509 22287 12514 22301
rect 12523 22297 12531 22301
rect 12715 22297 12723 22301
rect 12517 22287 12523 22297
rect 12709 22287 12715 22297
rect 12499 22286 12533 22287
rect 12451 22284 12533 22286
rect 12691 22286 12725 22287
rect 12726 22286 12733 22307
rect 12739 22301 12744 22311
rect 12749 22287 12754 22301
rect 12763 22297 12771 22301
rect 12757 22287 12763 22297
rect 12739 22286 12773 22287
rect 12691 22284 12773 22286
rect 6725 22274 6730 22277
rect 6725 22263 6730 22264
rect 6630 22236 6634 22260
rect 6715 22253 6720 22263
rect 6725 22250 6730 22253
rect 6725 22239 6730 22240
rect 6715 22236 6720 22239
rect 1405 22212 3171 22214
rect 1405 22211 1419 22212
rect 1422 22211 1429 22212
rect 1446 22190 1450 22212
rect 1470 22190 1474 22212
rect 1494 22190 1498 22212
rect 1518 22190 1522 22212
rect 1542 22190 1546 22212
rect 1566 22190 1570 22212
rect 1590 22190 1594 22212
rect 1614 22190 1618 22212
rect 1638 22190 1642 22212
rect 1662 22190 1666 22212
rect 1686 22190 1690 22212
rect 1710 22190 1714 22212
rect 1734 22190 1738 22212
rect 1758 22190 1762 22212
rect 1782 22190 1786 22212
rect 1806 22190 1810 22212
rect 1878 22190 1882 22212
rect 1902 22190 1906 22212
rect 1926 22190 1930 22212
rect 2022 22190 2026 22212
rect 2046 22190 2050 22212
rect 2070 22190 2074 22212
rect 2094 22190 2098 22212
rect 2118 22190 2122 22212
rect 2262 22190 2266 22212
rect 2286 22190 2290 22212
rect 2310 22190 2314 22212
rect 2502 22190 2506 22212
rect 2526 22190 2530 22212
rect 2550 22190 2554 22212
rect 2574 22190 2578 22212
rect 2598 22190 2602 22212
rect 2622 22190 2626 22212
rect 2646 22190 2650 22212
rect 2670 22190 2674 22212
rect 2694 22190 2698 22212
rect 2718 22190 2722 22212
rect 403 22188 2739 22190
rect 403 22181 408 22188
rect 414 22181 418 22188
rect 413 22167 418 22181
rect 438 22166 442 22188
rect 462 22166 466 22188
rect 486 22166 490 22188
rect 499 22166 533 22167
rect -2393 22164 533 22166
rect -2371 22142 -2366 22164
rect -2348 22142 -2343 22164
rect -2325 22158 -2317 22164
rect -2325 22142 -2320 22158
rect -2309 22146 -2301 22158
rect -2068 22147 -2038 22154
rect -2317 22142 -2309 22146
rect -2000 22144 -1992 22164
rect -1844 22156 -1794 22164
rect -1671 22158 -1663 22164
rect -1852 22147 -1804 22154
rect -1655 22146 -1647 22158
rect -2025 22143 -1991 22144
rect -2025 22142 -1975 22143
rect -1844 22142 -1804 22145
rect -1663 22142 -1655 22146
rect -1642 22142 -1637 22164
rect -1619 22142 -1614 22164
rect -1530 22142 -1526 22164
rect -1506 22142 -1502 22164
rect -1482 22142 -1478 22164
rect -1458 22142 -1454 22164
rect -1434 22142 -1430 22164
rect -1410 22142 -1406 22164
rect -1386 22142 -1382 22164
rect -1362 22142 -1358 22164
rect -1338 22142 -1334 22164
rect -1314 22142 -1310 22164
rect -1290 22142 -1286 22164
rect -1266 22142 -1262 22164
rect -1242 22142 -1238 22164
rect -1218 22142 -1214 22164
rect -1194 22142 -1190 22164
rect -1170 22142 -1166 22164
rect -1146 22142 -1142 22164
rect -1122 22142 -1118 22164
rect -1098 22142 -1094 22164
rect -1074 22142 -1070 22164
rect -1050 22142 -1046 22164
rect -1026 22142 -1022 22164
rect -1002 22142 -998 22164
rect -978 22142 -974 22164
rect -954 22142 -950 22164
rect -930 22142 -926 22164
rect -906 22142 -902 22164
rect -882 22142 -878 22164
rect -858 22142 -854 22164
rect -834 22142 -830 22164
rect -810 22142 -806 22164
rect -786 22142 -782 22164
rect -762 22142 -758 22164
rect -738 22142 -734 22164
rect -714 22142 -710 22164
rect -690 22142 -686 22164
rect -666 22142 -662 22164
rect -642 22142 -638 22164
rect -618 22142 -614 22164
rect -594 22142 -590 22164
rect -570 22142 -566 22164
rect -546 22142 -542 22164
rect -522 22142 -518 22164
rect -498 22142 -494 22164
rect -474 22142 -470 22164
rect -450 22142 -446 22164
rect -426 22142 -422 22164
rect -402 22142 -398 22164
rect -378 22142 -374 22164
rect -354 22142 -350 22164
rect -330 22142 -326 22164
rect -306 22142 -302 22164
rect -282 22142 -278 22164
rect -258 22142 -254 22164
rect -234 22142 -230 22164
rect -210 22142 -206 22164
rect -186 22142 -182 22164
rect -162 22142 -158 22164
rect -138 22142 -134 22164
rect -114 22142 -110 22164
rect -90 22142 -86 22164
rect -66 22142 -62 22164
rect -42 22142 -38 22164
rect -18 22142 -14 22164
rect 6 22142 10 22164
rect 30 22142 34 22164
rect 54 22142 58 22164
rect 78 22142 82 22164
rect 102 22142 106 22164
rect 126 22142 130 22164
rect 150 22142 154 22164
rect 174 22142 178 22164
rect 198 22142 202 22164
rect 222 22142 226 22164
rect 246 22142 250 22164
rect 270 22142 274 22164
rect 294 22142 298 22164
rect 318 22142 322 22164
rect 342 22142 346 22164
rect 366 22142 370 22164
rect 390 22143 394 22164
rect 379 22142 437 22143
rect 438 22142 442 22164
rect 462 22142 466 22164
rect 486 22142 490 22164
rect 499 22157 504 22164
rect 509 22143 514 22157
rect 510 22142 514 22143
rect 534 22142 538 22188
rect 558 22142 562 22188
rect 582 22142 586 22188
rect 606 22142 610 22188
rect 630 22142 634 22188
rect 654 22142 658 22188
rect 678 22167 682 22188
rect 667 22166 701 22167
rect 702 22166 706 22188
rect 726 22166 730 22188
rect 750 22166 754 22188
rect 774 22166 778 22188
rect 798 22166 802 22188
rect 822 22166 826 22188
rect 846 22166 850 22188
rect 918 22166 922 22188
rect 942 22166 946 22188
rect 966 22187 970 22188
rect 667 22164 963 22166
rect 667 22157 672 22164
rect 678 22157 682 22164
rect 677 22143 682 22157
rect 702 22142 706 22164
rect 726 22142 730 22164
rect 750 22142 754 22164
rect 774 22142 778 22164
rect 798 22142 802 22164
rect 822 22142 826 22164
rect 846 22142 850 22164
rect 918 22163 922 22164
rect 918 22142 925 22163
rect 942 22142 946 22164
rect 949 22163 963 22164
rect 966 22163 973 22187
rect 966 22142 970 22163
rect 990 22142 994 22188
rect 1014 22142 1018 22188
rect 1038 22142 1042 22188
rect 1062 22142 1066 22188
rect 1086 22142 1090 22188
rect 1110 22142 1114 22188
rect 1134 22142 1138 22188
rect 1158 22142 1162 22188
rect 1182 22142 1186 22188
rect 1206 22142 1210 22188
rect 1230 22142 1234 22188
rect 1254 22142 1258 22188
rect 1278 22142 1282 22188
rect 1302 22142 1306 22188
rect 1350 22187 1354 22188
rect 1350 22166 1357 22187
rect 1374 22166 1378 22188
rect 1446 22166 1450 22188
rect 1470 22166 1474 22188
rect 1494 22166 1498 22188
rect 1518 22166 1522 22188
rect 1542 22166 1546 22188
rect 1566 22166 1570 22188
rect 1590 22166 1594 22188
rect 1614 22166 1618 22188
rect 1638 22166 1642 22188
rect 1662 22166 1666 22188
rect 1686 22166 1690 22188
rect 1710 22166 1714 22188
rect 1734 22166 1738 22188
rect 1758 22166 1762 22188
rect 1782 22166 1786 22188
rect 1806 22166 1810 22188
rect 1878 22166 1882 22188
rect 1902 22166 1906 22188
rect 1926 22166 1930 22188
rect 2022 22166 2026 22188
rect 2046 22166 2050 22188
rect 2070 22166 2074 22188
rect 2094 22166 2098 22188
rect 2118 22166 2122 22188
rect 2179 22166 2237 22167
rect 2262 22166 2266 22188
rect 2286 22166 2290 22188
rect 2310 22166 2314 22188
rect 2502 22166 2506 22188
rect 2526 22166 2530 22188
rect 2550 22166 2554 22188
rect 2574 22166 2578 22188
rect 2598 22166 2602 22188
rect 2622 22166 2626 22188
rect 2646 22166 2650 22188
rect 2670 22166 2674 22188
rect 2694 22166 2698 22188
rect 2718 22166 2722 22188
rect 2725 22187 2739 22188
rect 2742 22187 2749 22211
rect 2742 22166 2746 22187
rect 2766 22166 2770 22212
rect 2790 22166 2794 22212
rect 2803 22205 2808 22212
rect 2827 22205 2832 22212
rect 2838 22211 2842 22212
rect 2838 22205 2845 22211
rect 2813 22191 2818 22205
rect 2827 22201 2835 22205
rect 2821 22191 2827 22201
rect 2837 22191 2845 22205
rect 2814 22166 2818 22191
rect 2862 22190 2866 22212
rect 3006 22190 3010 22212
rect 3030 22190 3034 22212
rect 3054 22190 3058 22212
rect 3078 22190 3082 22212
rect 3150 22190 3154 22212
rect 3157 22211 3171 22212
rect 3174 22211 3181 22235
rect 6596 22226 6600 22236
rect 3174 22190 3178 22211
rect 6568 22198 6576 22202
rect 2821 22188 3195 22190
rect 6606 22188 6610 22226
rect 6619 22212 6648 22215
rect 6654 22212 6658 22236
rect 6691 22212 6725 22215
rect 6750 22212 6754 22284
rect 6822 22260 6826 22284
rect 6853 22283 6867 22284
rect 6870 22283 6877 22284
rect 6870 22260 6874 22283
rect 6619 22205 6624 22212
rect 6629 22191 6634 22205
rect 2821 22187 2835 22188
rect 2862 22166 2866 22188
rect 3006 22166 3010 22188
rect 3030 22166 3034 22188
rect 3054 22166 3058 22188
rect 3078 22166 3082 22188
rect 3150 22166 3154 22188
rect 3174 22166 3178 22188
rect 3181 22187 3195 22188
rect 3222 22174 3229 22187
rect 1333 22164 3219 22166
rect 1333 22163 1347 22164
rect 1350 22163 1357 22164
rect 1374 22142 1378 22164
rect 1446 22142 1450 22164
rect 1470 22142 1474 22164
rect 1494 22142 1498 22164
rect 1518 22142 1522 22164
rect 1542 22142 1546 22164
rect 1566 22142 1570 22164
rect 1590 22142 1594 22164
rect 1614 22142 1618 22164
rect 1638 22142 1642 22164
rect 1662 22142 1666 22164
rect 1686 22142 1690 22164
rect 1710 22142 1714 22164
rect 1734 22142 1738 22164
rect 1758 22142 1762 22164
rect 1782 22142 1786 22164
rect 1806 22142 1810 22164
rect 1878 22142 1882 22164
rect 1902 22142 1906 22164
rect 1926 22142 1930 22164
rect 2022 22142 2026 22164
rect 2046 22142 2050 22164
rect 2070 22142 2074 22164
rect 2094 22142 2098 22164
rect 2118 22142 2122 22164
rect 2179 22157 2184 22164
rect 2189 22143 2194 22157
rect 2190 22142 2194 22143
rect 2262 22142 2266 22164
rect 2286 22142 2290 22164
rect 2310 22142 2314 22164
rect 2502 22142 2506 22164
rect 2526 22142 2530 22164
rect 2550 22142 2554 22164
rect 2574 22142 2578 22164
rect 2598 22142 2602 22164
rect 2622 22142 2626 22164
rect 2646 22142 2650 22164
rect 2670 22142 2674 22164
rect 2694 22142 2698 22164
rect 2718 22142 2722 22164
rect 2742 22142 2746 22164
rect 2766 22142 2770 22164
rect 2790 22142 2794 22164
rect 2814 22142 2818 22164
rect 2862 22142 2866 22164
rect 3006 22142 3010 22164
rect 3030 22142 3034 22164
rect 3054 22142 3058 22164
rect 3078 22142 3082 22164
rect 3091 22142 3149 22143
rect 3150 22142 3154 22164
rect 3174 22142 3178 22164
rect 3205 22163 3219 22164
rect 3222 22163 3229 22164
rect 3187 22142 3221 22143
rect -2393 22140 891 22142
rect -2371 22118 -2366 22140
rect -2348 22118 -2343 22140
rect -2325 22130 -2317 22140
rect -2060 22130 -2020 22137
rect -2004 22132 -2001 22137
rect -2015 22130 -2001 22132
rect -2000 22130 -1992 22140
rect -1972 22138 -1958 22140
rect -1844 22139 -1804 22140
rect -1862 22137 -1796 22138
rect -1985 22135 -1796 22137
rect -1985 22130 -1852 22135
rect -2325 22118 -2320 22130
rect -2309 22118 -2301 22130
rect -2068 22120 -2060 22127
rect -2015 22120 -1990 22130
rect -1844 22129 -1796 22135
rect -1671 22130 -1663 22140
rect -1852 22120 -1804 22127
rect -2020 22118 -2004 22120
rect -2000 22118 -1992 22120
rect -1976 22118 -1940 22119
rect -1655 22118 -1647 22130
rect -1642 22118 -1637 22140
rect -1619 22118 -1614 22140
rect -1530 22118 -1526 22140
rect -1506 22118 -1502 22140
rect -1482 22118 -1478 22140
rect -1458 22118 -1454 22140
rect -1434 22118 -1430 22140
rect -1410 22118 -1406 22140
rect -1386 22118 -1382 22140
rect -1362 22118 -1358 22140
rect -1338 22118 -1334 22140
rect -1314 22118 -1310 22140
rect -1290 22118 -1286 22140
rect -1266 22118 -1262 22140
rect -1242 22118 -1238 22140
rect -1218 22118 -1214 22140
rect -1194 22118 -1190 22140
rect -1170 22118 -1166 22140
rect -1146 22118 -1142 22140
rect -1122 22118 -1118 22140
rect -1098 22118 -1094 22140
rect -1074 22118 -1070 22140
rect -1050 22118 -1046 22140
rect -1026 22118 -1022 22140
rect -1002 22118 -998 22140
rect -978 22118 -974 22140
rect -954 22118 -950 22140
rect -930 22118 -926 22140
rect -906 22118 -902 22140
rect -882 22118 -878 22140
rect -858 22118 -854 22140
rect -834 22118 -830 22140
rect -810 22118 -806 22140
rect -786 22118 -782 22140
rect -762 22118 -758 22140
rect -738 22118 -734 22140
rect -714 22119 -710 22140
rect -725 22118 -691 22119
rect -2393 22116 -691 22118
rect -2371 22046 -2366 22116
rect -2348 22046 -2343 22116
rect -2325 22114 -2320 22116
rect -2317 22114 -2309 22116
rect -2325 22102 -2317 22114
rect -2060 22103 -2030 22110
rect -2325 22082 -2320 22102
rect -2325 22074 -2317 22082
rect -2060 22076 -2030 22079
rect -2325 22046 -2320 22074
rect -2317 22066 -2309 22074
rect -2060 22063 -2038 22074
rect -2033 22067 -2030 22076
rect -2028 22072 -2027 22076
rect -2068 22058 -2038 22061
rect -2000 22046 -1992 22116
rect -1844 22112 -1804 22116
rect -1663 22114 -1655 22116
rect -1844 22102 -1794 22111
rect -1671 22102 -1663 22114
rect -1912 22091 -1884 22093
rect -1852 22085 -1804 22089
rect -1844 22076 -1796 22079
rect -1671 22074 -1663 22082
rect -1844 22063 -1804 22074
rect -1663 22066 -1655 22074
rect -1852 22058 -1680 22062
rect -1642 22046 -1637 22116
rect -1619 22046 -1614 22116
rect -1530 22046 -1526 22116
rect -1506 22046 -1502 22116
rect -1482 22046 -1478 22116
rect -1458 22046 -1454 22116
rect -1434 22046 -1430 22116
rect -1410 22046 -1406 22116
rect -1386 22046 -1382 22116
rect -1362 22046 -1358 22116
rect -1338 22046 -1334 22116
rect -1314 22046 -1310 22116
rect -1290 22046 -1286 22116
rect -1266 22046 -1262 22116
rect -1242 22046 -1238 22116
rect -1218 22046 -1214 22116
rect -1194 22046 -1190 22116
rect -1170 22046 -1166 22116
rect -1146 22046 -1142 22116
rect -1122 22046 -1118 22116
rect -1098 22046 -1094 22116
rect -1074 22046 -1070 22116
rect -1050 22046 -1046 22116
rect -1026 22046 -1022 22116
rect -1002 22071 -998 22116
rect -1013 22070 -979 22071
rect -978 22070 -974 22116
rect -954 22070 -950 22116
rect -930 22070 -926 22116
rect -906 22070 -902 22116
rect -882 22070 -878 22116
rect -858 22070 -854 22116
rect -834 22070 -830 22116
rect -810 22070 -806 22116
rect -797 22085 -792 22095
rect -786 22085 -782 22116
rect -787 22071 -782 22085
rect -762 22070 -758 22116
rect -738 22070 -734 22116
rect -725 22109 -720 22116
rect -714 22109 -710 22116
rect -715 22095 -710 22109
rect -725 22085 -720 22095
rect -715 22071 -710 22085
rect -714 22070 -710 22071
rect -690 22070 -686 22140
rect -666 22070 -662 22140
rect -642 22070 -638 22140
rect -618 22072 -614 22140
rect -594 22119 -590 22140
rect -605 22118 -571 22119
rect -570 22118 -566 22140
rect -546 22118 -542 22140
rect -522 22118 -518 22140
rect -498 22118 -494 22140
rect -474 22118 -470 22140
rect -450 22118 -446 22140
rect -426 22118 -422 22140
rect -402 22118 -398 22140
rect -378 22118 -374 22140
rect -354 22118 -350 22140
rect -330 22118 -326 22140
rect -306 22118 -302 22140
rect -282 22118 -278 22140
rect -258 22118 -254 22140
rect -234 22118 -230 22140
rect -210 22118 -206 22140
rect -186 22118 -182 22140
rect -162 22118 -158 22140
rect -138 22118 -134 22140
rect -114 22118 -110 22140
rect -90 22118 -86 22140
rect -66 22118 -62 22140
rect -42 22118 -38 22140
rect -18 22118 -14 22140
rect 6 22118 10 22140
rect 30 22118 34 22140
rect 54 22118 58 22140
rect 78 22118 82 22140
rect 102 22118 106 22140
rect 126 22118 130 22140
rect 150 22118 154 22140
rect 174 22118 178 22140
rect 198 22118 202 22140
rect 222 22118 226 22140
rect 246 22118 250 22140
rect 270 22118 274 22140
rect 294 22118 298 22140
rect 318 22118 322 22140
rect 342 22118 346 22140
rect 366 22118 370 22140
rect 379 22133 384 22140
rect 390 22133 394 22140
rect 403 22133 408 22140
rect 389 22119 394 22133
rect 413 22130 418 22133
rect 413 22119 418 22120
rect 438 22118 442 22140
rect 462 22118 466 22140
rect 486 22118 490 22140
rect 510 22118 514 22140
rect 534 22139 538 22140
rect 534 22118 541 22139
rect 558 22118 562 22140
rect 582 22118 586 22140
rect 606 22118 610 22140
rect 630 22118 634 22140
rect 654 22118 658 22140
rect 702 22118 706 22140
rect 726 22118 730 22140
rect 750 22118 754 22140
rect 774 22118 778 22140
rect 798 22118 802 22140
rect 822 22118 826 22140
rect 846 22118 850 22140
rect 877 22139 891 22140
rect 901 22140 3221 22142
rect 901 22139 915 22140
rect 918 22139 925 22140
rect 942 22118 946 22140
rect 966 22118 970 22140
rect 990 22118 994 22140
rect 1014 22118 1018 22140
rect 1038 22118 1042 22140
rect 1062 22118 1066 22140
rect 1086 22118 1090 22140
rect 1110 22118 1114 22140
rect 1134 22118 1138 22140
rect 1158 22118 1162 22140
rect 1182 22118 1186 22140
rect 1206 22118 1210 22140
rect 1230 22118 1234 22140
rect 1254 22118 1258 22140
rect 1278 22118 1282 22140
rect 1302 22118 1306 22140
rect 1374 22118 1378 22140
rect 1446 22118 1450 22140
rect 1470 22118 1474 22140
rect 1494 22118 1498 22140
rect 1518 22118 1522 22140
rect 1542 22118 1546 22140
rect 1566 22118 1570 22140
rect 1590 22118 1594 22140
rect 1614 22118 1618 22140
rect 1638 22118 1642 22140
rect 1662 22118 1666 22140
rect 1686 22118 1690 22140
rect 1710 22118 1714 22140
rect 1734 22118 1738 22140
rect 1758 22118 1762 22140
rect 1782 22118 1786 22140
rect 1806 22118 1810 22140
rect 1878 22118 1882 22140
rect 1902 22118 1906 22140
rect 1926 22118 1930 22140
rect 2022 22118 2026 22140
rect 2046 22118 2050 22140
rect 2070 22118 2074 22140
rect 2094 22118 2098 22140
rect 2118 22118 2122 22140
rect 2190 22118 2194 22140
rect 2262 22118 2266 22140
rect 2286 22118 2290 22140
rect 2310 22118 2314 22140
rect 2323 22118 2381 22119
rect 2502 22118 2506 22140
rect 2526 22118 2530 22140
rect 2550 22118 2554 22140
rect 2574 22118 2578 22140
rect 2598 22118 2602 22140
rect 2622 22118 2626 22140
rect 2646 22118 2650 22140
rect 2670 22118 2674 22140
rect 2694 22118 2698 22140
rect 2718 22118 2722 22140
rect 2742 22118 2746 22140
rect 2766 22118 2770 22140
rect 2790 22118 2794 22140
rect 2814 22118 2818 22140
rect 2862 22139 2866 22140
rect 2862 22118 2869 22139
rect 3006 22118 3010 22140
rect 3030 22118 3034 22140
rect 3054 22118 3058 22140
rect 3078 22118 3082 22140
rect 3091 22133 3096 22140
rect 3101 22119 3106 22133
rect 3102 22118 3106 22119
rect 3150 22118 3154 22140
rect 3174 22118 3178 22140
rect 3187 22133 3192 22140
rect 3197 22119 3202 22133
rect 3198 22118 3202 22119
rect 3246 22118 3250 22184
rect 6582 22178 6586 22188
rect 6592 22174 6600 22178
rect 3270 22139 3277 22163
rect 3859 22157 3864 22167
rect 4579 22157 4584 22167
rect 4819 22157 4824 22167
rect 6571 22157 6576 22167
rect 6619 22164 6624 22167
rect 6630 22164 6634 22191
rect 6678 22188 6682 22212
rect 6715 22190 6749 22191
rect 6750 22190 6757 22211
rect 6774 22190 6778 22260
rect 6822 22238 6829 22259
rect 6846 22238 6850 22260
rect 6894 22238 6898 22284
rect 6925 22283 6939 22284
rect 6942 22283 6949 22284
rect 6997 22283 7011 22284
rect 7014 22262 7021 22284
rect 7027 22277 7032 22284
rect 7045 22283 7059 22284
rect 10549 22283 10563 22284
rect 7037 22263 7042 22277
rect 7051 22273 7059 22277
rect 10555 22273 10563 22277
rect 7045 22263 7051 22273
rect 10549 22263 10555 22273
rect 7027 22262 7061 22263
rect 6997 22260 7061 22262
rect 10531 22262 10565 22263
rect 10566 22262 10573 22284
rect 10579 22277 10584 22284
rect 10597 22283 10611 22284
rect 11989 22283 12003 22284
rect 10589 22263 10594 22277
rect 10603 22273 10611 22277
rect 11995 22273 12003 22277
rect 10597 22263 10603 22273
rect 11989 22263 11995 22273
rect 10579 22262 10613 22263
rect 10531 22260 10613 22262
rect 11971 22262 12005 22263
rect 12006 22262 12013 22284
rect 12019 22277 12024 22284
rect 12037 22283 12051 22284
rect 12469 22283 12483 22284
rect 12029 22263 12034 22277
rect 12043 22273 12051 22277
rect 12475 22273 12483 22277
rect 12037 22263 12043 22273
rect 12469 22263 12475 22273
rect 12019 22262 12053 22263
rect 11971 22260 12053 22262
rect 12451 22262 12485 22263
rect 12486 22262 12493 22284
rect 12499 22277 12504 22284
rect 12517 22283 12531 22284
rect 12709 22283 12723 22284
rect 12509 22263 12514 22277
rect 12523 22273 12531 22277
rect 12715 22273 12723 22277
rect 12517 22263 12523 22273
rect 12709 22263 12715 22273
rect 12499 22262 12533 22263
rect 12451 22260 12533 22262
rect 12691 22262 12725 22263
rect 12726 22262 12733 22284
rect 12739 22277 12744 22284
rect 12757 22283 12771 22284
rect 13939 22277 13944 22287
rect 12749 22263 12754 22277
rect 12763 22273 12771 22277
rect 12757 22263 12763 22273
rect 13949 22263 13954 22277
rect 12739 22262 12773 22263
rect 12691 22260 12773 22262
rect 6942 22259 6946 22260
rect 6997 22259 7011 22260
rect 6805 22236 6939 22238
rect 6805 22235 6819 22236
rect 6787 22205 6792 22215
rect 6805 22214 6821 22215
rect 6822 22214 6829 22236
rect 6846 22214 6850 22236
rect 6894 22214 6898 22236
rect 6925 22235 6939 22236
rect 6942 22235 6949 22259
rect 7014 22238 7021 22260
rect 7027 22253 7032 22260
rect 7045 22259 7059 22260
rect 10549 22259 10563 22260
rect 7037 22239 7042 22253
rect 7051 22249 7059 22253
rect 10555 22249 10563 22253
rect 7045 22239 7051 22249
rect 10549 22239 10555 22249
rect 7027 22238 7061 22239
rect 6997 22236 7061 22238
rect 10531 22238 10565 22239
rect 10566 22238 10573 22260
rect 10579 22253 10584 22260
rect 10597 22259 10611 22260
rect 11989 22259 12003 22260
rect 10589 22239 10594 22253
rect 10603 22249 10611 22253
rect 11995 22249 12003 22253
rect 10597 22239 10603 22249
rect 11989 22239 11995 22249
rect 10579 22238 10613 22239
rect 10531 22236 10613 22238
rect 11971 22238 12005 22239
rect 12006 22238 12013 22260
rect 12019 22253 12024 22260
rect 12037 22259 12051 22260
rect 12469 22259 12483 22260
rect 12029 22239 12034 22253
rect 12043 22249 12051 22253
rect 12475 22249 12483 22253
rect 12037 22239 12043 22249
rect 12469 22239 12475 22249
rect 12019 22238 12053 22239
rect 11971 22236 12053 22238
rect 12451 22238 12485 22239
rect 12486 22238 12493 22260
rect 12499 22253 12504 22260
rect 12517 22259 12531 22260
rect 12709 22259 12723 22260
rect 12509 22239 12514 22253
rect 12523 22249 12531 22253
rect 12715 22249 12723 22253
rect 12517 22239 12523 22249
rect 12709 22239 12715 22249
rect 12499 22238 12533 22239
rect 12451 22236 12533 22238
rect 12691 22238 12725 22239
rect 12726 22238 12733 22260
rect 12739 22253 12744 22260
rect 12757 22259 12771 22260
rect 13939 22253 13944 22263
rect 12749 22239 12754 22253
rect 12763 22249 12771 22253
rect 12757 22239 12763 22249
rect 13949 22239 13954 22253
rect 12739 22238 12773 22239
rect 12691 22236 12773 22238
rect 6997 22235 7011 22236
rect 7014 22235 7021 22236
rect 7027 22229 7032 22236
rect 7045 22235 7059 22236
rect 10549 22235 10563 22236
rect 7037 22215 7042 22229
rect 7051 22225 7059 22229
rect 10555 22225 10563 22229
rect 7045 22215 7051 22225
rect 10549 22215 10555 22225
rect 7027 22214 7061 22215
rect 6805 22212 7061 22214
rect 10531 22214 10565 22215
rect 10566 22214 10573 22236
rect 10579 22229 10584 22236
rect 10597 22235 10611 22236
rect 11989 22235 12003 22236
rect 10589 22215 10594 22229
rect 10603 22225 10611 22229
rect 11995 22225 12003 22229
rect 10597 22215 10603 22225
rect 11989 22215 11995 22225
rect 10579 22214 10613 22215
rect 10531 22212 10613 22214
rect 11971 22214 12005 22215
rect 12006 22214 12013 22236
rect 12019 22229 12024 22236
rect 12037 22235 12051 22236
rect 12469 22235 12483 22236
rect 12029 22215 12034 22229
rect 12043 22225 12051 22229
rect 12475 22225 12483 22229
rect 12037 22215 12043 22225
rect 12469 22215 12475 22225
rect 12019 22214 12053 22215
rect 11971 22212 12053 22214
rect 12451 22214 12485 22215
rect 12486 22214 12493 22236
rect 12499 22229 12504 22236
rect 12517 22235 12531 22236
rect 12709 22235 12723 22236
rect 12509 22215 12514 22229
rect 12523 22225 12531 22229
rect 12715 22225 12723 22229
rect 12517 22215 12523 22225
rect 12709 22215 12715 22225
rect 12499 22214 12533 22215
rect 12451 22212 12533 22214
rect 12691 22214 12725 22215
rect 12726 22214 12733 22236
rect 12739 22229 12744 22236
rect 12757 22235 12771 22236
rect 13939 22229 13944 22239
rect 12749 22215 12754 22229
rect 12763 22225 12771 22229
rect 12757 22215 12763 22225
rect 13949 22215 13954 22229
rect 12739 22214 12773 22215
rect 12691 22212 12773 22214
rect 6805 22211 6819 22212
rect 6797 22191 6802 22205
rect 6811 22201 6819 22205
rect 6805 22191 6811 22201
rect 6787 22190 6819 22191
rect 6715 22188 6819 22190
rect 3869 22143 3874 22157
rect 4589 22143 4594 22157
rect 4829 22143 4834 22157
rect 6581 22143 6586 22157
rect 3270 22118 3274 22139
rect 3294 22120 3301 22139
rect 3859 22133 3864 22143
rect 4579 22133 4584 22143
rect 4819 22133 4824 22143
rect 3869 22119 3874 22133
rect 4589 22119 4594 22133
rect 4829 22119 4834 22133
rect 6547 22126 6552 22129
rect 3283 22118 3291 22119
rect -605 22116 2835 22118
rect -605 22109 -600 22116
rect -594 22109 -590 22116
rect -595 22095 -590 22109
rect -605 22085 -600 22095
rect -595 22082 -590 22085
rect -595 22071 -590 22072
rect -629 22070 -571 22071
rect -570 22070 -566 22116
rect -546 22070 -542 22116
rect -522 22070 -518 22116
rect -498 22070 -494 22116
rect -474 22070 -470 22116
rect -450 22070 -446 22116
rect -426 22070 -422 22116
rect -402 22070 -398 22116
rect -378 22070 -374 22116
rect -354 22070 -350 22116
rect -330 22070 -326 22116
rect -306 22070 -302 22116
rect -282 22070 -278 22116
rect -258 22070 -254 22116
rect -234 22070 -230 22116
rect -210 22070 -206 22116
rect -186 22070 -182 22116
rect -162 22070 -158 22116
rect -138 22070 -134 22116
rect -114 22070 -110 22116
rect -90 22070 -86 22116
rect -66 22070 -62 22116
rect -42 22070 -38 22116
rect -18 22070 -14 22116
rect 6 22070 10 22116
rect 30 22070 34 22116
rect 54 22070 58 22116
rect 78 22070 82 22116
rect 102 22070 106 22116
rect 126 22070 130 22116
rect 150 22070 154 22116
rect 174 22070 178 22116
rect 198 22070 202 22116
rect 222 22070 226 22116
rect 246 22070 250 22116
rect 270 22070 274 22116
rect 294 22070 298 22116
rect 318 22070 322 22116
rect 342 22070 346 22116
rect 366 22070 370 22116
rect 438 22115 442 22116
rect 438 22094 445 22115
rect 462 22094 466 22116
rect 486 22094 490 22116
rect 510 22094 514 22116
rect 517 22115 531 22116
rect 534 22115 541 22116
rect 558 22094 562 22116
rect 582 22094 586 22116
rect 606 22094 610 22116
rect 630 22094 634 22116
rect 654 22094 658 22116
rect 702 22094 706 22116
rect 726 22094 730 22116
rect 750 22094 754 22116
rect 774 22094 778 22116
rect 798 22094 802 22116
rect 822 22094 826 22116
rect 846 22094 850 22116
rect 942 22094 946 22116
rect 966 22094 970 22116
rect 990 22094 994 22116
rect 1014 22094 1018 22116
rect 1038 22094 1042 22116
rect 1062 22094 1066 22116
rect 1086 22094 1090 22116
rect 1110 22094 1114 22116
rect 1134 22094 1138 22116
rect 1158 22094 1162 22116
rect 1182 22094 1186 22116
rect 1206 22094 1210 22116
rect 1230 22094 1234 22116
rect 1254 22094 1258 22116
rect 1278 22094 1282 22116
rect 1302 22094 1306 22116
rect 1374 22094 1378 22116
rect 1446 22094 1450 22116
rect 1470 22094 1474 22116
rect 1494 22094 1498 22116
rect 1518 22094 1522 22116
rect 1542 22094 1546 22116
rect 1566 22094 1570 22116
rect 1590 22094 1594 22116
rect 1614 22094 1618 22116
rect 1638 22094 1642 22116
rect 1662 22094 1666 22116
rect 1686 22094 1690 22116
rect 1710 22094 1714 22116
rect 1734 22094 1738 22116
rect 1758 22094 1762 22116
rect 1782 22094 1786 22116
rect 1806 22094 1810 22116
rect 1878 22094 1882 22116
rect 1902 22094 1906 22116
rect 1926 22094 1930 22116
rect 1939 22094 1997 22095
rect 2022 22094 2026 22116
rect 2046 22094 2050 22116
rect 2070 22094 2074 22116
rect 2094 22094 2098 22116
rect 2118 22094 2122 22116
rect 2190 22094 2194 22116
rect 2203 22094 2237 22095
rect 421 22092 2237 22094
rect 421 22091 435 22092
rect 438 22091 445 22092
rect 462 22070 466 22092
rect 486 22070 490 22092
rect 510 22070 514 22092
rect -1013 22068 531 22070
rect -1013 22061 -1008 22068
rect -1002 22061 -998 22068
rect -1003 22047 -998 22061
rect -1013 22046 -979 22047
rect -2393 22044 -979 22046
rect -2371 22022 -2366 22044
rect -2348 22022 -2343 22044
rect -2325 22022 -2320 22044
rect -2309 22026 -2301 22036
rect -2068 22027 -2062 22032
rect -2317 22022 -2309 22026
rect -2060 22022 -2050 22027
rect -2000 22022 -1992 22044
rect -1806 22036 -1680 22042
rect -1854 22027 -1806 22032
rect -1655 22026 -1647 22036
rect -1972 22022 -1964 22023
rect -1958 22022 -1942 22024
rect -1844 22022 -1806 22025
rect -1663 22022 -1655 22026
rect -1642 22022 -1637 22044
rect -1619 22022 -1614 22044
rect -1530 22022 -1526 22044
rect -1506 22022 -1502 22044
rect -1482 22022 -1478 22044
rect -1458 22022 -1454 22044
rect -1434 22022 -1430 22044
rect -1410 22022 -1406 22044
rect -1386 22022 -1382 22044
rect -1362 22022 -1358 22044
rect -1338 22022 -1334 22044
rect -1314 22022 -1310 22044
rect -1290 22022 -1286 22044
rect -1266 22022 -1262 22044
rect -1242 22022 -1238 22044
rect -1218 22022 -1214 22044
rect -1194 22022 -1190 22044
rect -1170 22022 -1166 22044
rect -1146 22022 -1142 22044
rect -1122 22022 -1118 22044
rect -1098 22022 -1094 22044
rect -1074 22022 -1070 22044
rect -1050 22022 -1046 22044
rect -1026 22022 -1022 22044
rect -1013 22037 -1008 22044
rect -1003 22023 -998 22037
rect -1002 22022 -998 22023
rect -978 22022 -974 22068
rect -954 22022 -950 22068
rect -930 22022 -926 22068
rect -906 22022 -902 22068
rect -882 22022 -878 22068
rect -858 22022 -854 22068
rect -834 22022 -830 22068
rect -810 22022 -806 22068
rect -797 22046 -763 22047
rect -762 22046 -758 22068
rect -738 22046 -734 22068
rect -714 22046 -710 22068
rect -690 22046 -686 22068
rect -666 22046 -662 22068
rect -642 22046 -638 22068
rect -629 22061 -624 22068
rect -605 22061 -600 22068
rect -619 22047 -614 22061
rect -595 22047 -590 22061
rect -618 22046 -614 22047
rect -594 22046 -590 22047
rect -570 22046 -566 22068
rect -546 22046 -542 22068
rect -522 22046 -518 22068
rect -498 22046 -494 22068
rect -474 22046 -470 22068
rect -450 22046 -446 22068
rect -426 22046 -422 22068
rect -402 22046 -398 22068
rect -378 22046 -374 22068
rect -354 22046 -350 22068
rect -330 22046 -326 22068
rect -306 22046 -302 22068
rect -282 22046 -278 22068
rect -258 22046 -254 22068
rect -234 22046 -230 22068
rect -210 22046 -206 22068
rect -186 22046 -182 22068
rect -162 22046 -158 22068
rect -138 22046 -134 22068
rect -114 22046 -110 22068
rect -90 22046 -86 22068
rect -66 22046 -62 22068
rect -42 22046 -38 22068
rect -18 22046 -14 22068
rect 6 22046 10 22068
rect 30 22046 34 22068
rect 54 22046 58 22068
rect 78 22046 82 22068
rect 102 22046 106 22068
rect 126 22046 130 22068
rect 150 22046 154 22068
rect 174 22046 178 22068
rect 198 22046 202 22068
rect 222 22046 226 22068
rect 246 22046 250 22068
rect 270 22046 274 22068
rect 294 22046 298 22068
rect 318 22046 322 22068
rect 342 22046 346 22068
rect 366 22046 370 22068
rect 438 22046 445 22067
rect 462 22046 466 22068
rect 486 22046 490 22068
rect 510 22046 514 22068
rect 517 22067 531 22068
rect 534 22067 541 22091
rect 534 22046 538 22067
rect 558 22046 562 22092
rect 582 22046 586 22092
rect 606 22046 610 22092
rect 630 22046 634 22092
rect 654 22046 658 22092
rect 702 22091 706 22092
rect 702 22070 709 22091
rect 726 22070 730 22092
rect 750 22070 754 22092
rect 774 22070 778 22092
rect 798 22070 802 22092
rect 822 22070 826 22092
rect 846 22070 850 22092
rect 942 22070 946 22092
rect 966 22070 970 22092
rect 990 22070 994 22092
rect 1014 22070 1018 22092
rect 1038 22070 1042 22092
rect 1062 22070 1066 22092
rect 1086 22070 1090 22092
rect 1110 22070 1114 22092
rect 1134 22070 1138 22092
rect 1158 22070 1162 22092
rect 1182 22070 1186 22092
rect 1206 22070 1210 22092
rect 1230 22070 1234 22092
rect 1254 22070 1258 22092
rect 1278 22070 1282 22092
rect 1302 22070 1306 22092
rect 1374 22071 1378 22092
rect 1363 22070 1421 22071
rect 1446 22070 1450 22092
rect 1470 22070 1474 22092
rect 1494 22070 1498 22092
rect 1518 22070 1522 22092
rect 1542 22070 1546 22092
rect 1566 22070 1570 22092
rect 1590 22070 1594 22092
rect 1614 22070 1618 22092
rect 1638 22070 1642 22092
rect 1662 22070 1666 22092
rect 1686 22070 1690 22092
rect 1710 22070 1714 22092
rect 1734 22070 1738 22092
rect 1758 22070 1762 22092
rect 1782 22070 1786 22092
rect 1806 22070 1810 22092
rect 1878 22070 1882 22092
rect 1902 22070 1906 22092
rect 1926 22070 1930 22092
rect 1939 22085 1944 22092
rect 1949 22071 1954 22085
rect 1950 22070 1954 22071
rect 1963 22070 1997 22071
rect 685 22068 1997 22070
rect 685 22067 699 22068
rect 702 22067 709 22068
rect 726 22046 730 22068
rect 750 22046 754 22068
rect 774 22046 778 22068
rect 798 22046 802 22068
rect 822 22046 826 22068
rect 846 22046 850 22068
rect 942 22046 946 22068
rect 966 22046 970 22068
rect 990 22046 994 22068
rect 1014 22046 1018 22068
rect 1038 22046 1042 22068
rect 1062 22046 1066 22068
rect 1086 22046 1090 22068
rect 1110 22046 1114 22068
rect 1134 22046 1138 22068
rect 1158 22046 1162 22068
rect 1182 22046 1186 22068
rect 1206 22046 1210 22068
rect 1230 22046 1234 22068
rect 1254 22046 1258 22068
rect 1278 22046 1282 22068
rect 1302 22046 1306 22068
rect 1363 22061 1368 22068
rect 1374 22061 1378 22068
rect 1387 22061 1392 22068
rect 1373 22047 1378 22061
rect 1397 22047 1402 22061
rect 1398 22046 1402 22047
rect 1446 22046 1450 22068
rect 1470 22046 1474 22068
rect 1494 22046 1498 22068
rect 1518 22046 1522 22068
rect 1542 22046 1546 22068
rect 1566 22046 1570 22068
rect 1590 22046 1594 22068
rect 1614 22046 1618 22068
rect 1638 22046 1642 22068
rect 1662 22046 1666 22068
rect 1686 22046 1690 22068
rect 1710 22046 1714 22068
rect 1734 22046 1738 22068
rect 1758 22046 1762 22068
rect 1782 22046 1786 22068
rect 1806 22046 1810 22068
rect 1878 22046 1882 22068
rect 1902 22046 1906 22068
rect 1926 22046 1930 22068
rect 1950 22046 1954 22068
rect 2022 22046 2026 22092
rect 2046 22046 2050 22092
rect 2070 22046 2074 22092
rect 2094 22046 2098 22092
rect 2118 22046 2122 22092
rect 2131 22070 2165 22071
rect 2190 22070 2194 22092
rect 2214 22085 2221 22091
rect 2213 22081 2221 22085
rect 2227 22081 2235 22085
rect 2213 22071 2227 22081
rect 2238 22070 2245 22091
rect 2262 22070 2266 22116
rect 2286 22070 2290 22116
rect 2310 22070 2314 22116
rect 2323 22109 2328 22116
rect 2333 22095 2338 22109
rect 2334 22070 2338 22095
rect 2443 22094 2477 22095
rect 2502 22094 2506 22116
rect 2526 22094 2530 22116
rect 2550 22094 2554 22116
rect 2574 22094 2578 22116
rect 2598 22094 2602 22116
rect 2622 22094 2626 22116
rect 2646 22094 2650 22116
rect 2670 22094 2674 22116
rect 2694 22094 2698 22116
rect 2718 22094 2722 22116
rect 2742 22094 2746 22116
rect 2766 22094 2770 22116
rect 2790 22094 2794 22116
rect 2814 22094 2818 22116
rect 2821 22115 2835 22116
rect 2845 22116 3291 22118
rect 2845 22115 2859 22116
rect 2862 22115 2869 22116
rect 3006 22094 3010 22116
rect 3030 22094 3034 22116
rect 3054 22094 3058 22116
rect 3078 22094 3082 22116
rect 3102 22094 3106 22116
rect 3150 22094 3154 22116
rect 3174 22094 3178 22116
rect 3198 22094 3202 22116
rect 3246 22094 3250 22116
rect 3270 22094 3274 22116
rect 3277 22115 3291 22116
rect 3283 22109 3288 22115
rect 3859 22109 3864 22119
rect 4579 22109 4584 22119
rect 4819 22109 4824 22119
rect 6582 22116 6586 22143
rect 3293 22095 3298 22109
rect 3307 22105 3315 22109
rect 3301 22095 3307 22105
rect 3869 22095 3874 22109
rect 4589 22095 4594 22109
rect 4829 22095 4834 22109
rect 6558 22106 6562 22116
rect 6568 22102 6576 22106
rect 3283 22094 3315 22095
rect 2443 22092 3315 22094
rect 2443 22085 2448 22092
rect 2453 22071 2458 22085
rect 2347 22070 2381 22071
rect 2131 22068 2211 22070
rect 2131 22061 2136 22068
rect 2141 22047 2146 22061
rect 2142 22046 2146 22047
rect 2190 22046 2194 22068
rect 2197 22067 2211 22068
rect 2221 22068 2381 22070
rect 2221 22067 2235 22068
rect 2238 22067 2245 22068
rect 2238 22046 2242 22067
rect 2262 22046 2266 22068
rect 2286 22046 2290 22068
rect 2310 22046 2314 22068
rect 2334 22046 2338 22068
rect 2454 22046 2458 22071
rect 2502 22046 2506 22092
rect 2526 22046 2530 22092
rect 2550 22046 2554 22092
rect 2574 22046 2578 22092
rect 2598 22046 2602 22092
rect 2622 22046 2626 22092
rect 2646 22046 2650 22092
rect 2670 22046 2674 22092
rect 2694 22046 2698 22092
rect 2718 22046 2722 22092
rect 2742 22046 2746 22092
rect 2766 22046 2770 22092
rect 2790 22046 2794 22092
rect 2814 22046 2818 22092
rect 2827 22070 2861 22071
rect 3006 22070 3010 22092
rect 3030 22070 3034 22092
rect 3054 22070 3058 22092
rect 3078 22070 3082 22092
rect 3102 22070 3106 22092
rect 3150 22070 3154 22092
rect 3174 22070 3178 22092
rect 3198 22070 3202 22092
rect 3246 22070 3250 22092
rect 3270 22070 3274 22092
rect 3283 22085 3288 22092
rect 3301 22091 3315 22092
rect 3293 22071 3298 22085
rect 3835 22081 3843 22085
rect 3829 22071 3835 22081
rect 3283 22070 3317 22071
rect 2827 22068 3317 22070
rect 3811 22070 3845 22071
rect 3846 22070 3853 22091
rect 3859 22085 3864 22095
rect 3869 22071 3874 22085
rect 3883 22081 3891 22085
rect 4555 22081 4563 22085
rect 3877 22071 3883 22081
rect 4549 22071 4555 22081
rect 3859 22070 3893 22071
rect 3811 22068 3893 22070
rect 4531 22070 4565 22071
rect 4566 22070 4573 22091
rect 4579 22085 4584 22095
rect 4589 22071 4594 22085
rect 4603 22081 4611 22085
rect 4795 22081 4803 22085
rect 4597 22071 4603 22081
rect 4789 22071 4795 22081
rect 4579 22070 4613 22071
rect 4531 22068 4613 22070
rect 4771 22070 4805 22071
rect 4806 22070 4813 22091
rect 4819 22085 4824 22095
rect 6547 22085 6552 22095
rect 6606 22092 6610 22164
rect 6654 22140 6658 22188
rect 6692 22178 6696 22188
rect 6733 22187 6747 22188
rect 6702 22164 6706 22178
rect 6739 22177 6747 22181
rect 6733 22167 6739 22177
rect 6715 22166 6749 22167
rect 6750 22166 6757 22188
rect 6774 22166 6778 22188
rect 6787 22181 6792 22188
rect 6798 22181 6802 22188
rect 6805 22187 6819 22188
rect 6822 22187 6829 22212
rect 6797 22167 6802 22181
rect 6846 22166 6850 22212
rect 6870 22187 6877 22211
rect 6870 22166 6874 22187
rect 6894 22166 6898 22212
rect 7027 22205 7032 22212
rect 7045 22211 7059 22212
rect 10549 22211 10563 22212
rect 7037 22191 7042 22205
rect 7051 22201 7059 22205
rect 10555 22201 10563 22205
rect 7045 22191 7051 22201
rect 10549 22191 10555 22201
rect 6907 22190 6941 22191
rect 7027 22190 7061 22191
rect 6907 22188 7061 22190
rect 10531 22190 10565 22191
rect 10566 22190 10573 22212
rect 10579 22205 10584 22212
rect 10597 22211 10611 22212
rect 11989 22211 12003 22212
rect 10589 22191 10594 22205
rect 10603 22201 10611 22205
rect 11995 22201 12003 22205
rect 10597 22191 10603 22201
rect 11989 22191 11995 22201
rect 10579 22190 10613 22191
rect 10531 22188 10613 22190
rect 11971 22190 12005 22191
rect 12006 22190 12013 22212
rect 12019 22205 12024 22212
rect 12037 22211 12051 22212
rect 12469 22211 12483 22212
rect 12029 22191 12034 22205
rect 12043 22201 12051 22205
rect 12475 22201 12483 22205
rect 12037 22191 12043 22201
rect 12469 22191 12475 22201
rect 12019 22190 12053 22191
rect 11971 22188 12053 22190
rect 12451 22190 12485 22191
rect 12486 22190 12493 22212
rect 12499 22205 12504 22212
rect 12517 22211 12531 22212
rect 12709 22211 12723 22212
rect 12509 22191 12514 22205
rect 12523 22201 12531 22205
rect 12715 22201 12723 22205
rect 12517 22191 12523 22201
rect 12709 22191 12715 22201
rect 12499 22190 12533 22191
rect 12451 22188 12533 22190
rect 12691 22190 12725 22191
rect 12726 22190 12733 22212
rect 12739 22205 12744 22212
rect 12757 22211 12771 22212
rect 12749 22191 12754 22205
rect 12763 22201 12771 22205
rect 13915 22201 13923 22205
rect 12757 22191 12763 22201
rect 13909 22191 13915 22201
rect 12739 22190 12773 22191
rect 12691 22188 12773 22190
rect 13891 22190 13925 22191
rect 13926 22190 13933 22211
rect 13939 22205 13944 22215
rect 13949 22191 13954 22205
rect 13963 22201 13971 22205
rect 13957 22191 13963 22201
rect 13939 22190 13973 22191
rect 13891 22188 13973 22190
rect 6907 22181 6912 22188
rect 7027 22181 7032 22188
rect 7045 22187 7059 22188
rect 10549 22187 10563 22188
rect 6917 22167 6922 22181
rect 7037 22167 7042 22181
rect 7051 22177 7059 22181
rect 10555 22177 10563 22181
rect 7045 22167 7051 22177
rect 10549 22167 10555 22177
rect 6918 22166 6922 22167
rect 7027 22166 7061 22167
rect 6715 22164 7061 22166
rect 10531 22166 10565 22167
rect 10566 22166 10573 22188
rect 10579 22181 10584 22188
rect 10597 22187 10611 22188
rect 11989 22187 12003 22188
rect 10589 22167 10594 22181
rect 10603 22177 10611 22181
rect 11995 22177 12003 22181
rect 10597 22167 10603 22177
rect 11989 22167 11995 22177
rect 10579 22166 10613 22167
rect 10531 22164 10613 22166
rect 11971 22166 12005 22167
rect 12006 22166 12013 22188
rect 12019 22181 12024 22188
rect 12037 22187 12051 22188
rect 12469 22187 12483 22188
rect 12029 22167 12034 22181
rect 12043 22177 12051 22181
rect 12475 22177 12483 22181
rect 12037 22167 12043 22177
rect 12469 22167 12475 22177
rect 12019 22166 12053 22167
rect 11971 22164 12053 22166
rect 12451 22166 12485 22167
rect 12486 22166 12493 22188
rect 12499 22181 12504 22188
rect 12517 22187 12531 22188
rect 12709 22187 12723 22188
rect 12509 22167 12514 22181
rect 12523 22177 12531 22181
rect 12715 22177 12723 22181
rect 12517 22167 12523 22177
rect 12709 22167 12715 22177
rect 12499 22166 12533 22167
rect 12451 22164 12533 22166
rect 12691 22166 12725 22167
rect 12726 22166 12733 22188
rect 12739 22181 12744 22188
rect 12757 22187 12771 22188
rect 13909 22187 13923 22188
rect 12749 22167 12754 22181
rect 12763 22177 12771 22181
rect 13915 22177 13923 22181
rect 12757 22167 12763 22177
rect 13909 22167 13915 22177
rect 12739 22166 12773 22167
rect 12691 22164 12773 22166
rect 13891 22166 13925 22167
rect 13926 22166 13933 22188
rect 13939 22181 13944 22188
rect 13957 22187 13971 22188
rect 13949 22167 13954 22181
rect 13963 22177 13971 22181
rect 13957 22167 13963 22177
rect 13939 22166 13973 22167
rect 13891 22164 13973 22166
rect 6619 22109 6624 22119
rect 6637 22118 6653 22119
rect 6654 22118 6661 22139
rect 6678 22118 6682 22164
rect 6715 22157 6720 22164
rect 6733 22163 6747 22164
rect 6725 22143 6730 22157
rect 6739 22153 6747 22157
rect 6733 22143 6739 22153
rect 6726 22140 6730 22143
rect 6750 22142 6757 22164
rect 6774 22142 6778 22164
rect 6846 22142 6850 22164
rect 6870 22142 6874 22164
rect 6894 22142 6898 22164
rect 6918 22142 6922 22164
rect 7027 22157 7032 22164
rect 7045 22163 7059 22164
rect 10549 22163 10563 22164
rect 7037 22143 7042 22157
rect 7051 22153 7059 22157
rect 10555 22153 10563 22157
rect 7045 22143 7051 22153
rect 10549 22143 10555 22153
rect 7027 22142 7061 22143
rect 6733 22140 7061 22142
rect 6702 22118 6706 22140
rect 6733 22139 6747 22140
rect 6750 22139 6757 22140
rect 6726 22126 6733 22139
rect 6637 22116 6723 22118
rect 6750 22116 6754 22139
rect 6637 22115 6651 22116
rect 6654 22115 6661 22116
rect 6629 22095 6634 22109
rect 4829 22071 4834 22085
rect 4843 22081 4851 22085
rect 6557 22082 6562 22085
rect 4837 22071 4843 22081
rect 6557 22071 6562 22072
rect 4819 22070 4853 22071
rect 4771 22068 4853 22070
rect 6547 22068 6552 22071
rect 2827 22061 2832 22068
rect 2837 22047 2842 22061
rect 2838 22046 2842 22047
rect 3006 22046 3010 22068
rect 3030 22046 3034 22068
rect 3054 22046 3058 22068
rect 3078 22046 3082 22068
rect 3102 22046 3106 22068
rect 3150 22067 3154 22068
rect 3150 22046 3157 22067
rect 3174 22046 3178 22068
rect 3198 22046 3202 22068
rect -797 22044 411 22046
rect -797 22037 -792 22044
rect -787 22023 -782 22037
rect -786 22022 -782 22023
rect -762 22022 -758 22044
rect -738 22022 -734 22044
rect -714 22022 -710 22044
rect -690 22043 -686 22044
rect -2393 22020 -693 22022
rect -2371 21998 -2366 22020
rect -2348 21998 -2343 22020
rect -2325 21998 -2320 22020
rect -2060 22014 -2050 22020
rect -2309 21998 -2301 22008
rect -2060 22007 -2030 22014
rect -2000 22010 -1992 22020
rect -1972 22018 -1942 22020
rect -1958 22017 -1942 22018
rect -1844 22016 -1806 22020
rect -2068 22000 -2062 22007
rect -2062 21998 -2036 22000
rect -2393 21996 -2036 21998
rect -2030 21998 -2012 22000
rect -2004 21998 -1990 22010
rect -1844 22009 -1798 22014
rect -1806 22007 -1798 22009
rect -1854 22005 -1844 22007
rect -1854 22000 -1806 22005
rect -1864 21998 -1796 21999
rect -1655 21998 -1647 22008
rect -1642 21998 -1637 22020
rect -1619 21998 -1614 22020
rect -1530 21998 -1526 22020
rect -1506 21998 -1502 22020
rect -1482 21998 -1478 22020
rect -1458 21998 -1454 22020
rect -1434 21998 -1430 22020
rect -1410 21998 -1406 22020
rect -1386 21998 -1382 22020
rect -1362 21998 -1358 22020
rect -1338 21998 -1334 22020
rect -1314 21998 -1310 22020
rect -1290 21998 -1286 22020
rect -1266 21998 -1262 22020
rect -1242 21998 -1238 22020
rect -1218 21998 -1214 22020
rect -1194 21998 -1190 22020
rect -1170 21998 -1166 22020
rect -1146 21998 -1142 22020
rect -1122 21998 -1118 22020
rect -1098 21998 -1094 22020
rect -1074 21998 -1070 22020
rect -1050 21998 -1046 22020
rect -1026 21998 -1022 22020
rect -1002 21998 -998 22020
rect -978 21998 -974 22020
rect -954 21998 -950 22020
rect -930 21998 -926 22020
rect -906 21998 -902 22020
rect -882 21998 -878 22020
rect -858 21998 -854 22020
rect -834 21998 -830 22020
rect -810 21998 -806 22020
rect -786 21998 -782 22020
rect -762 22019 -758 22020
rect -762 21998 -755 22019
rect -738 21998 -734 22020
rect -714 21998 -710 22020
rect -707 22019 -693 22020
rect -701 21998 -693 21999
rect -2030 21996 -693 21998
rect -2371 21950 -2366 21996
rect -2348 21950 -2343 21996
rect -2325 21950 -2320 21996
rect -2317 21992 -2309 21996
rect -2060 21992 -2050 21996
rect -2060 21990 -2036 21992
rect -2060 21988 -2030 21990
rect -2292 21982 -2030 21988
rect -2092 21966 -2062 21968
rect -2094 21962 -2062 21966
rect -2000 21950 -1992 21996
rect -1844 21989 -1806 21996
rect -1663 21992 -1655 21996
rect -1844 21982 -1680 21988
rect -1854 21966 -1806 21968
rect -1854 21962 -1680 21966
rect -1642 21950 -1637 21996
rect -1619 21950 -1614 21996
rect -1530 21950 -1526 21996
rect -1506 21950 -1502 21996
rect -1482 21950 -1478 21996
rect -1458 21950 -1454 21996
rect -1434 21950 -1430 21996
rect -1410 21950 -1406 21996
rect -1386 21950 -1382 21996
rect -1362 21950 -1358 21996
rect -1338 21950 -1334 21996
rect -1314 21950 -1310 21996
rect -1290 21950 -1286 21996
rect -1266 21950 -1262 21996
rect -1242 21950 -1238 21996
rect -1218 21950 -1214 21996
rect -1194 21950 -1190 21996
rect -1170 21950 -1166 21996
rect -1146 21950 -1142 21996
rect -1122 21950 -1118 21996
rect -1098 21950 -1094 21996
rect -1074 21950 -1070 21996
rect -1050 21950 -1046 21996
rect -1026 21950 -1022 21996
rect -1002 21950 -998 21996
rect -978 21995 -974 21996
rect -2393 21948 -981 21950
rect -2371 21926 -2366 21948
rect -2348 21926 -2343 21948
rect -2325 21926 -2320 21948
rect -2072 21946 -2036 21947
rect -2072 21940 -2054 21946
rect -2309 21932 -2301 21940
rect -2317 21926 -2309 21932
rect -2092 21931 -2062 21936
rect -2000 21927 -1992 21948
rect -1938 21947 -1906 21948
rect -1920 21946 -1906 21947
rect -1806 21940 -1680 21946
rect -1854 21931 -1806 21936
rect -1655 21932 -1647 21940
rect -1982 21927 -1966 21928
rect -2000 21926 -1966 21927
rect -1846 21926 -1806 21929
rect -1663 21926 -1655 21932
rect -1642 21926 -1637 21948
rect -1619 21926 -1614 21948
rect -1530 21926 -1526 21948
rect -1506 21926 -1502 21948
rect -1482 21926 -1478 21948
rect -1458 21926 -1454 21948
rect -1434 21926 -1430 21948
rect -1410 21926 -1406 21948
rect -1386 21926 -1382 21948
rect -1362 21926 -1358 21948
rect -1338 21926 -1334 21948
rect -1314 21926 -1310 21948
rect -1290 21926 -1286 21948
rect -1266 21926 -1262 21948
rect -1242 21926 -1238 21948
rect -1218 21926 -1214 21948
rect -1194 21926 -1190 21948
rect -1170 21926 -1166 21948
rect -1146 21926 -1142 21948
rect -1122 21926 -1118 21948
rect -1098 21926 -1094 21948
rect -1074 21926 -1070 21948
rect -1050 21926 -1046 21948
rect -1026 21926 -1022 21948
rect -1002 21926 -998 21948
rect -995 21947 -981 21948
rect -978 21947 -971 21995
rect -978 21926 -974 21947
rect -954 21926 -950 21996
rect -930 21926 -926 21996
rect -906 21926 -902 21996
rect -882 21926 -878 21996
rect -858 21926 -854 21996
rect -834 21926 -830 21996
rect -810 21926 -806 21996
rect -786 21926 -782 21996
rect -779 21995 -765 21996
rect -762 21995 -755 21996
rect -762 21950 -755 21971
rect -738 21950 -734 21996
rect -714 21950 -710 21996
rect -707 21995 -693 21996
rect -690 21995 -683 22043
rect -701 21989 -696 21995
rect -690 21989 -686 21995
rect -691 21975 -686 21989
rect -701 21974 -667 21975
rect -666 21974 -662 22044
rect -642 21974 -638 22044
rect -618 21974 -614 22044
rect -594 22006 -590 22044
rect -570 22043 -566 22044
rect -570 22022 -563 22043
rect -546 22022 -542 22044
rect -522 22022 -518 22044
rect -498 22022 -494 22044
rect -474 22022 -470 22044
rect -450 22022 -446 22044
rect -426 22022 -422 22044
rect -402 22022 -398 22044
rect -378 22022 -374 22044
rect -354 22022 -350 22044
rect -330 22022 -326 22044
rect -306 22022 -302 22044
rect -282 22022 -278 22044
rect -258 22022 -254 22044
rect -234 22022 -230 22044
rect -210 22023 -206 22044
rect -221 22022 -187 22023
rect -587 22020 -187 22022
rect -587 22019 -573 22020
rect -594 21974 -587 21995
rect -570 21974 -563 22020
rect -546 21974 -542 22020
rect -522 21974 -518 22020
rect -498 21974 -494 22020
rect -474 21974 -470 22020
rect -450 21974 -446 22020
rect -426 21974 -422 22020
rect -402 21974 -398 22020
rect -378 21974 -374 22020
rect -354 21974 -350 22020
rect -330 21974 -326 22020
rect -306 21974 -302 22020
rect -282 21974 -278 22020
rect -258 21974 -254 22020
rect -234 21974 -230 22020
rect -221 22013 -216 22020
rect -210 22013 -206 22020
rect -211 21999 -206 22013
rect -221 21998 -187 21999
rect -186 21998 -182 22044
rect -162 21998 -158 22044
rect -138 21998 -134 22044
rect -114 21998 -110 22044
rect -90 21998 -86 22044
rect -66 21998 -62 22044
rect -42 21998 -38 22044
rect -18 21998 -14 22044
rect 6 21998 10 22044
rect 30 21998 34 22044
rect 54 21998 58 22044
rect 78 21998 82 22044
rect 102 21998 106 22044
rect 126 21998 130 22044
rect 150 21998 154 22044
rect 174 21998 178 22044
rect 198 22023 202 22044
rect 187 22022 221 22023
rect 222 22022 226 22044
rect 246 22022 250 22044
rect 270 22022 274 22044
rect 294 22022 298 22044
rect 318 22022 322 22044
rect 342 22022 346 22044
rect 366 22022 370 22044
rect 397 22043 411 22044
rect 421 22044 3123 22046
rect 421 22043 435 22044
rect 438 22043 445 22044
rect 462 22022 466 22044
rect 486 22022 490 22044
rect 510 22022 514 22044
rect 534 22022 538 22044
rect 558 22022 562 22044
rect 582 22022 586 22044
rect 606 22022 610 22044
rect 630 22022 634 22044
rect 654 22022 658 22044
rect 726 22022 730 22044
rect 750 22022 754 22044
rect 774 22022 778 22044
rect 798 22022 802 22044
rect 822 22022 826 22044
rect 846 22022 850 22044
rect 859 22022 917 22023
rect 942 22022 946 22044
rect 966 22022 970 22044
rect 990 22022 994 22044
rect 1014 22022 1018 22044
rect 1038 22022 1042 22044
rect 1062 22022 1066 22044
rect 1086 22022 1090 22044
rect 1110 22022 1114 22044
rect 1134 22022 1138 22044
rect 1158 22022 1162 22044
rect 1182 22022 1186 22044
rect 1206 22022 1210 22044
rect 1230 22022 1234 22044
rect 1254 22022 1258 22044
rect 1278 22022 1282 22044
rect 1302 22022 1306 22044
rect 1315 22022 1349 22023
rect 187 22020 1349 22022
rect 187 22013 192 22020
rect 198 22013 202 22020
rect 197 21999 202 22013
rect 222 21998 226 22020
rect 246 21998 250 22020
rect 270 21998 274 22020
rect 294 21998 298 22020
rect 318 21998 322 22020
rect 342 21998 346 22020
rect 366 21998 370 22020
rect 462 21998 466 22020
rect 486 21998 490 22020
rect 510 21998 514 22020
rect 534 21998 538 22020
rect 558 21998 562 22020
rect 582 21998 586 22020
rect 606 21998 610 22020
rect 630 21998 634 22020
rect 654 21998 658 22020
rect 726 21998 730 22020
rect 750 21998 754 22020
rect 774 21998 778 22020
rect 798 21998 802 22020
rect 822 21998 826 22020
rect 846 21998 850 22020
rect 859 22013 864 22020
rect 869 21999 874 22013
rect 870 21998 874 21999
rect 883 21998 917 21999
rect -221 21996 917 21998
rect -221 21989 -216 21996
rect -211 21975 -206 21989
rect -210 21974 -206 21975
rect -186 21974 -182 21996
rect -162 21974 -158 21996
rect -138 21974 -134 21996
rect -114 21974 -110 21996
rect -90 21974 -86 21996
rect -66 21974 -62 21996
rect -42 21974 -38 21996
rect -18 21974 -14 21996
rect 6 21974 10 21996
rect 30 21974 34 21996
rect 54 21974 58 21996
rect 78 21974 82 21996
rect 102 21974 106 21996
rect 126 21974 130 21996
rect 150 21974 154 21996
rect 174 21974 178 21996
rect 222 21974 226 21996
rect 246 21974 250 21996
rect 270 21974 274 21996
rect 294 21974 298 21996
rect 318 21974 322 21996
rect 342 21974 346 21996
rect 366 21974 370 21996
rect 462 21974 466 21996
rect 486 21974 490 21996
rect 510 21974 514 21996
rect 534 21974 538 21996
rect 558 21974 562 21996
rect 582 21974 586 21996
rect 606 21974 610 21996
rect 630 21974 634 21996
rect 654 21974 658 21996
rect 726 21974 730 21996
rect 750 21974 754 21996
rect 774 21974 778 21996
rect 798 21974 802 21996
rect 822 21974 826 21996
rect 846 21974 850 21996
rect 870 21974 874 21996
rect 942 21974 946 22020
rect 966 21974 970 22020
rect 990 21974 994 22020
rect 1014 21974 1018 22020
rect 1038 21974 1042 22020
rect 1062 21974 1066 22020
rect 1086 21974 1090 22020
rect 1110 21974 1114 22020
rect 1134 21974 1138 22020
rect 1158 21974 1162 22020
rect 1182 21974 1186 22020
rect 1206 21974 1210 22020
rect 1230 21974 1234 22020
rect 1254 21974 1258 22020
rect 1278 21974 1282 22020
rect 1302 21974 1306 22020
rect 1315 22013 1320 22020
rect 1325 21999 1330 22013
rect 1364 22010 1368 22020
rect 1398 22010 1402 22044
rect 1316 21986 1320 21996
rect 1374 21986 1378 22010
rect 1387 21998 1421 21999
rect 1446 21998 1450 22044
rect 1470 21998 1474 22044
rect 1494 21998 1498 22044
rect 1518 21998 1522 22044
rect 1542 21998 1546 22044
rect 1566 21998 1570 22044
rect 1590 21998 1594 22044
rect 1614 21998 1618 22044
rect 1638 21998 1642 22044
rect 1662 21998 1666 22044
rect 1686 21998 1690 22044
rect 1710 21998 1714 22044
rect 1734 21998 1738 22044
rect 1758 21998 1762 22044
rect 1782 21998 1786 22044
rect 1806 21998 1810 22044
rect 1819 22022 1853 22023
rect 1878 22022 1882 22044
rect 1902 22022 1906 22044
rect 1926 22022 1930 22044
rect 1950 22022 1954 22044
rect 2022 22022 2026 22044
rect 2046 22022 2050 22044
rect 2070 22022 2074 22044
rect 2094 22022 2098 22044
rect 2118 22022 2122 22044
rect 2142 22023 2146 22044
rect 2131 22022 2165 22023
rect 1819 22020 2165 22022
rect 1819 22013 1824 22020
rect 1829 21999 1834 22013
rect 1830 21998 1834 21999
rect 1878 21998 1882 22020
rect 1902 21998 1906 22020
rect 1926 21998 1930 22020
rect 1950 21998 1954 22020
rect 1998 21998 2005 22019
rect 2022 21998 2026 22020
rect 2046 21998 2050 22020
rect 2070 21998 2074 22020
rect 2094 21998 2098 22020
rect 2118 21998 2122 22020
rect 2131 22013 2136 22020
rect 2142 22013 2146 22020
rect 2141 21999 2146 22013
rect 2190 21998 2194 22044
rect 2203 22022 2237 22023
rect 2238 22022 2242 22044
rect 2262 22022 2266 22044
rect 2286 22022 2290 22044
rect 2310 22022 2314 22044
rect 2334 22022 2338 22044
rect 2382 22022 2389 22043
rect 2454 22023 2458 22044
rect 2443 22022 2477 22023
rect 2203 22020 2355 22022
rect 2203 22013 2208 22020
rect 2238 22019 2242 22020
rect 2213 21999 2218 22013
rect 2227 22009 2235 22013
rect 2221 21999 2227 22009
rect 2214 21998 2218 21999
rect 1387 21996 1971 21998
rect 1387 21989 1392 21996
rect 1326 21974 1330 21986
rect 1397 21985 1405 21989
rect 1411 21985 1419 21989
rect 1397 21975 1411 21985
rect 1398 21974 1405 21975
rect 1422 21974 1429 21995
rect 1446 21974 1450 21996
rect 1470 21974 1474 21996
rect 1494 21974 1498 21996
rect 1518 21974 1522 21996
rect 1542 21974 1546 21996
rect 1566 21974 1570 21996
rect 1590 21974 1594 21996
rect 1614 21974 1618 21996
rect 1638 21974 1642 21996
rect 1662 21974 1666 21996
rect 1686 21974 1690 21996
rect 1710 21974 1714 21996
rect 1734 21974 1738 21996
rect 1758 21974 1762 21996
rect 1782 21974 1786 21996
rect 1806 21974 1810 21996
rect 1830 21974 1834 21996
rect 1878 21974 1882 21996
rect 1902 21974 1906 21996
rect 1926 21974 1930 21996
rect 1950 21974 1954 21996
rect 1957 21995 1971 21996
rect 1981 21996 2235 21998
rect 1981 21995 1995 21996
rect -701 21972 -597 21974
rect -701 21965 -696 21972
rect -691 21951 -686 21965
rect -690 21950 -686 21951
rect -666 21950 -662 21972
rect -642 21950 -638 21972
rect -618 21950 -614 21972
rect -611 21971 -597 21972
rect -594 21972 1395 21974
rect -594 21971 -573 21972
rect -570 21971 -563 21972
rect -594 21950 -590 21971
rect -570 21950 -566 21971
rect -546 21950 -542 21972
rect -522 21950 -518 21972
rect -498 21950 -494 21972
rect -474 21950 -470 21972
rect -450 21950 -446 21972
rect -426 21950 -422 21972
rect -402 21950 -398 21972
rect -378 21950 -374 21972
rect -354 21950 -350 21972
rect -330 21950 -326 21972
rect -306 21950 -302 21972
rect -282 21950 -278 21972
rect -258 21950 -254 21972
rect -234 21950 -230 21972
rect -210 21950 -206 21972
rect -186 21950 -182 21972
rect -162 21950 -158 21972
rect -138 21950 -134 21972
rect -114 21950 -110 21972
rect -90 21950 -86 21972
rect -66 21950 -62 21972
rect -42 21950 -38 21972
rect -18 21950 -14 21972
rect 6 21950 10 21972
rect 30 21950 34 21972
rect 54 21950 58 21972
rect 78 21950 82 21972
rect 102 21950 106 21972
rect 126 21950 130 21972
rect 150 21950 154 21972
rect 174 21950 178 21972
rect 222 21950 226 21972
rect 246 21950 250 21972
rect 270 21950 274 21972
rect 294 21950 298 21972
rect 318 21950 322 21972
rect 342 21950 346 21972
rect 366 21950 370 21972
rect 462 21950 466 21972
rect 486 21950 490 21972
rect 510 21950 514 21972
rect 534 21950 538 21972
rect 558 21950 562 21972
rect 582 21950 586 21972
rect 606 21950 610 21972
rect 630 21950 634 21972
rect 654 21950 658 21972
rect 726 21950 730 21972
rect 750 21950 754 21972
rect 774 21950 778 21972
rect 798 21950 802 21972
rect 822 21950 826 21972
rect 846 21950 850 21972
rect 870 21950 874 21972
rect 942 21950 946 21972
rect 966 21950 970 21972
rect 990 21950 994 21972
rect 1014 21950 1018 21972
rect 1038 21950 1042 21972
rect 1062 21950 1066 21972
rect 1086 21950 1090 21972
rect 1110 21950 1114 21972
rect 1134 21950 1138 21972
rect 1158 21950 1162 21972
rect 1182 21950 1186 21972
rect 1206 21950 1210 21972
rect 1230 21950 1234 21972
rect 1254 21950 1258 21972
rect 1278 21950 1282 21972
rect 1302 21950 1306 21972
rect 1326 21950 1330 21972
rect 1381 21971 1395 21972
rect 1398 21972 1995 21974
rect 1398 21971 1419 21972
rect 1422 21971 1429 21972
rect 1422 21950 1426 21971
rect 1446 21950 1450 21972
rect 1470 21950 1474 21972
rect 1494 21950 1498 21972
rect 1518 21950 1522 21972
rect 1542 21950 1546 21972
rect 1566 21950 1570 21972
rect 1590 21950 1594 21972
rect 1614 21950 1618 21972
rect 1638 21950 1642 21972
rect 1662 21950 1666 21972
rect 1686 21950 1690 21972
rect 1710 21950 1714 21972
rect 1734 21950 1738 21972
rect 1758 21950 1762 21972
rect 1782 21950 1786 21972
rect 1806 21950 1810 21972
rect 1830 21950 1834 21972
rect 1878 21950 1882 21972
rect 1902 21950 1906 21972
rect 1926 21950 1930 21972
rect 1950 21950 1954 21972
rect 1981 21971 1995 21972
rect 1998 21971 2005 21996
rect 1963 21950 1997 21951
rect -779 21948 1997 21950
rect -779 21947 -765 21948
rect -762 21947 -755 21948
rect -762 21926 -758 21947
rect -738 21926 -734 21948
rect -714 21926 -710 21948
rect -690 21926 -686 21948
rect -666 21926 -662 21948
rect -642 21926 -638 21948
rect -618 21926 -614 21948
rect -594 21926 -590 21948
rect -570 21926 -566 21948
rect -546 21926 -542 21948
rect -522 21926 -518 21948
rect -498 21926 -494 21948
rect -474 21926 -470 21948
rect -450 21926 -446 21948
rect -426 21926 -422 21948
rect -402 21926 -398 21948
rect -378 21926 -374 21948
rect -354 21926 -350 21948
rect -330 21926 -326 21948
rect -306 21926 -302 21948
rect -282 21926 -278 21948
rect -258 21926 -254 21948
rect -234 21926 -230 21948
rect -210 21926 -206 21948
rect -186 21947 -182 21948
rect -2393 21924 -189 21926
rect -2371 21902 -2366 21924
rect -2348 21902 -2343 21924
rect -2325 21902 -2320 21924
rect -2000 21922 -1966 21924
rect -2309 21904 -2301 21912
rect -2062 21911 -2054 21918
rect -2092 21904 -2084 21911
rect -2062 21904 -2026 21906
rect -2317 21902 -2309 21904
rect -2062 21902 -2012 21904
rect -2000 21902 -1992 21922
rect -1982 21921 -1966 21922
rect -1846 21920 -1806 21924
rect -1846 21913 -1798 21918
rect -1806 21911 -1798 21913
rect -1854 21909 -1846 21911
rect -1854 21904 -1806 21909
rect -1655 21904 -1647 21912
rect -1864 21902 -1796 21903
rect -1663 21902 -1655 21904
rect -1642 21902 -1637 21924
rect -1619 21902 -1614 21924
rect -1530 21902 -1526 21924
rect -1506 21902 -1502 21924
rect -1482 21902 -1478 21924
rect -1458 21902 -1454 21924
rect -1434 21902 -1430 21924
rect -1410 21902 -1406 21924
rect -1386 21902 -1382 21924
rect -1362 21902 -1358 21924
rect -1338 21902 -1334 21924
rect -1314 21902 -1310 21924
rect -1290 21902 -1286 21924
rect -1266 21902 -1262 21924
rect -1242 21902 -1238 21924
rect -1218 21902 -1214 21924
rect -1194 21902 -1190 21924
rect -1170 21902 -1166 21924
rect -1146 21902 -1142 21924
rect -1122 21902 -1118 21924
rect -1098 21902 -1094 21924
rect -1074 21902 -1070 21924
rect -1050 21902 -1046 21924
rect -1026 21903 -1022 21924
rect -1037 21902 -1003 21903
rect -1002 21902 -998 21924
rect -978 21902 -974 21924
rect -954 21902 -950 21924
rect -930 21902 -926 21924
rect -906 21902 -902 21924
rect -882 21902 -878 21924
rect -858 21902 -854 21924
rect -834 21902 -830 21924
rect -810 21902 -806 21924
rect -786 21902 -782 21924
rect -762 21902 -758 21924
rect -738 21902 -734 21924
rect -714 21902 -710 21924
rect -690 21902 -686 21924
rect -666 21923 -662 21924
rect -2393 21900 -669 21902
rect -2371 21854 -2366 21900
rect -2348 21854 -2343 21900
rect -2325 21854 -2320 21900
rect -2317 21896 -2309 21900
rect -2062 21896 -2054 21900
rect -2154 21892 -2138 21894
rect -2057 21892 -2054 21896
rect -2292 21886 -2054 21892
rect -2052 21886 -2044 21896
rect -2092 21870 -2062 21872
rect -2094 21866 -2062 21870
rect -2000 21854 -1992 21900
rect -1846 21893 -1806 21900
rect -1663 21896 -1655 21900
rect -1846 21886 -1680 21892
rect -1854 21870 -1806 21872
rect -1854 21866 -1680 21870
rect -1642 21854 -1637 21900
rect -1619 21854 -1614 21900
rect -1530 21854 -1526 21900
rect -1506 21854 -1502 21900
rect -1482 21854 -1478 21900
rect -1458 21854 -1454 21900
rect -1434 21854 -1430 21900
rect -1410 21854 -1406 21900
rect -1386 21854 -1382 21900
rect -1362 21854 -1358 21900
rect -1338 21854 -1334 21900
rect -1314 21854 -1310 21900
rect -1290 21854 -1286 21900
rect -1266 21854 -1262 21900
rect -1242 21854 -1238 21900
rect -1218 21854 -1214 21900
rect -1194 21854 -1190 21900
rect -1170 21854 -1166 21900
rect -1146 21854 -1142 21900
rect -1122 21854 -1118 21900
rect -1098 21854 -1094 21900
rect -1074 21854 -1070 21900
rect -1050 21854 -1046 21900
rect -1037 21893 -1032 21900
rect -1026 21893 -1022 21900
rect -1027 21879 -1022 21893
rect -1037 21869 -1032 21879
rect -1027 21855 -1022 21869
rect -1026 21854 -1022 21855
rect -1002 21854 -998 21900
rect -978 21854 -974 21900
rect -954 21854 -950 21900
rect -930 21854 -926 21900
rect -906 21854 -902 21900
rect -882 21854 -878 21900
rect -858 21854 -854 21900
rect -834 21854 -830 21900
rect -810 21854 -806 21900
rect -786 21854 -782 21900
rect -762 21854 -758 21900
rect -738 21854 -734 21900
rect -714 21854 -710 21900
rect -690 21854 -686 21900
rect -683 21899 -669 21900
rect -666 21878 -659 21923
rect -642 21878 -638 21924
rect -618 21878 -614 21924
rect -594 21878 -590 21924
rect -570 21878 -566 21924
rect -546 21878 -542 21924
rect -522 21878 -518 21924
rect -498 21878 -494 21924
rect -474 21878 -470 21924
rect -450 21878 -446 21924
rect -426 21878 -422 21924
rect -402 21878 -398 21924
rect -378 21878 -374 21924
rect -354 21878 -350 21924
rect -330 21878 -326 21924
rect -306 21878 -302 21924
rect -282 21878 -278 21924
rect -258 21878 -254 21924
rect -234 21878 -230 21924
rect -210 21878 -206 21924
rect -203 21923 -189 21924
rect -186 21902 -179 21947
rect -162 21902 -158 21948
rect -149 21917 -144 21927
rect -138 21917 -134 21948
rect -139 21903 -134 21917
rect -114 21902 -110 21948
rect -90 21902 -86 21948
rect -66 21902 -62 21948
rect -42 21902 -38 21948
rect -18 21902 -14 21948
rect -5 21917 0 21927
rect 6 21917 10 21948
rect 5 21903 10 21917
rect 30 21902 34 21948
rect 54 21902 58 21948
rect 78 21902 82 21948
rect 102 21902 106 21948
rect 126 21902 130 21948
rect 150 21902 154 21948
rect 174 21902 178 21948
rect 222 21947 226 21948
rect 222 21926 229 21947
rect 246 21926 250 21948
rect 270 21926 274 21948
rect 294 21926 298 21948
rect 318 21926 322 21948
rect 342 21926 346 21948
rect 366 21926 370 21948
rect 379 21926 437 21927
rect 462 21926 466 21948
rect 486 21926 490 21948
rect 510 21926 514 21948
rect 534 21926 538 21948
rect 558 21926 562 21948
rect 582 21926 586 21948
rect 606 21926 610 21948
rect 630 21926 634 21948
rect 654 21926 658 21948
rect 726 21926 730 21948
rect 750 21926 754 21948
rect 774 21926 778 21948
rect 798 21926 802 21948
rect 822 21926 826 21948
rect 846 21926 850 21948
rect 870 21926 874 21948
rect 918 21926 925 21947
rect 942 21926 946 21948
rect 966 21926 970 21948
rect 990 21926 994 21948
rect 1014 21926 1018 21948
rect 1038 21926 1042 21948
rect 1062 21926 1066 21948
rect 1086 21926 1090 21948
rect 1110 21926 1114 21948
rect 1134 21926 1138 21948
rect 1158 21926 1162 21948
rect 1182 21926 1186 21948
rect 1206 21926 1210 21948
rect 1230 21926 1234 21948
rect 1254 21926 1258 21948
rect 1278 21926 1282 21948
rect 1302 21926 1306 21948
rect 1326 21927 1330 21948
rect 1315 21926 1349 21927
rect 205 21924 891 21926
rect 205 21923 219 21924
rect 222 21923 229 21924
rect 246 21902 250 21924
rect 270 21902 274 21924
rect 294 21902 298 21924
rect 318 21902 322 21924
rect 342 21902 346 21924
rect 366 21902 370 21924
rect 379 21917 384 21924
rect 389 21903 394 21917
rect 390 21902 394 21903
rect 462 21902 466 21924
rect 486 21902 490 21924
rect 510 21902 514 21924
rect 534 21902 538 21924
rect 558 21902 562 21924
rect 582 21902 586 21924
rect 606 21902 610 21924
rect 630 21902 634 21924
rect 654 21902 658 21924
rect 726 21902 730 21924
rect 750 21902 754 21924
rect 774 21902 778 21924
rect 798 21902 802 21924
rect 822 21902 826 21924
rect 846 21902 850 21924
rect 870 21902 874 21924
rect 877 21923 891 21924
rect 901 21924 1349 21926
rect 1422 21924 1426 21948
rect 901 21923 915 21924
rect 883 21902 915 21903
rect -203 21900 915 21902
rect -203 21899 -189 21900
rect -186 21899 -179 21900
rect -186 21878 -182 21899
rect -162 21878 -158 21900
rect -114 21878 -110 21900
rect -90 21878 -86 21900
rect -66 21878 -62 21900
rect -42 21878 -38 21900
rect -18 21878 -14 21900
rect 30 21878 34 21900
rect 54 21878 58 21900
rect 78 21878 82 21900
rect 102 21878 106 21900
rect 126 21878 130 21900
rect 150 21878 154 21900
rect 174 21878 178 21900
rect 246 21878 250 21900
rect 270 21878 274 21900
rect 294 21878 298 21900
rect 318 21878 322 21900
rect 342 21878 346 21900
rect 366 21878 370 21900
rect 390 21878 394 21900
rect 462 21878 466 21900
rect 486 21878 490 21900
rect 510 21878 514 21900
rect 534 21878 538 21900
rect 558 21878 562 21900
rect 582 21878 586 21900
rect 606 21878 610 21900
rect 630 21878 634 21900
rect 654 21878 658 21900
rect 726 21878 730 21900
rect 750 21878 754 21900
rect 774 21878 778 21900
rect 798 21878 802 21900
rect 822 21878 826 21900
rect 846 21878 850 21900
rect 870 21878 874 21900
rect 883 21893 888 21900
rect 901 21899 915 21900
rect 918 21899 925 21924
rect 893 21879 898 21893
rect 894 21878 898 21879
rect 942 21878 946 21924
rect 966 21878 970 21924
rect 990 21878 994 21924
rect 1014 21878 1018 21924
rect 1038 21878 1042 21924
rect 1062 21878 1066 21924
rect 1086 21878 1090 21924
rect 1110 21878 1114 21924
rect 1134 21878 1138 21924
rect 1158 21878 1162 21924
rect 1182 21878 1186 21924
rect 1206 21878 1210 21924
rect 1219 21893 1224 21903
rect 1230 21893 1234 21924
rect 1229 21879 1234 21893
rect 1254 21878 1258 21924
rect 1278 21878 1282 21924
rect 1302 21878 1306 21924
rect 1315 21917 1320 21924
rect 1326 21917 1330 21924
rect 1333 21923 1347 21924
rect 1325 21903 1330 21917
rect 1398 21914 1402 21924
rect 1408 21913 1415 21914
rect 1339 21910 1344 21913
rect 1315 21893 1320 21903
rect 1387 21900 1392 21903
rect 1405 21902 1421 21903
rect 1422 21902 1429 21923
rect 1446 21902 1450 21948
rect 1470 21902 1474 21948
rect 1494 21902 1498 21948
rect 1518 21902 1522 21948
rect 1542 21902 1546 21948
rect 1566 21902 1570 21948
rect 1590 21902 1594 21948
rect 1614 21902 1618 21948
rect 1638 21902 1642 21948
rect 1662 21902 1666 21948
rect 1686 21902 1690 21948
rect 1710 21902 1714 21948
rect 1734 21902 1738 21948
rect 1758 21902 1762 21948
rect 1782 21902 1786 21948
rect 1806 21902 1810 21948
rect 1830 21902 1834 21948
rect 1854 21923 1861 21947
rect 1854 21902 1858 21923
rect 1878 21902 1882 21948
rect 1902 21902 1906 21948
rect 1926 21902 1930 21948
rect 1950 21902 1954 21948
rect 1963 21941 1968 21948
rect 1973 21927 1978 21941
rect 1974 21902 1978 21927
rect 2022 21902 2026 21996
rect 2046 21902 2050 21996
rect 2070 21902 2074 21996
rect 2094 21902 2098 21996
rect 2118 21902 2122 21996
rect 2166 21974 2173 21995
rect 2190 21974 2194 21996
rect 2214 21974 2218 21996
rect 2221 21995 2235 21996
rect 2238 21995 2245 22019
rect 2262 21974 2266 22020
rect 2286 21974 2290 22020
rect 2310 21974 2314 22020
rect 2334 21974 2338 22020
rect 2341 22019 2355 22020
rect 2365 22020 2477 22022
rect 2365 22019 2379 22020
rect 2382 22019 2389 22020
rect 2382 21995 2386 22019
rect 2443 22013 2448 22020
rect 2454 22013 2458 22020
rect 2453 21999 2458 22013
rect 2467 22009 2475 22013
rect 2461 21999 2467 22009
rect 2478 21998 2485 22019
rect 2502 21998 2506 22044
rect 2526 21998 2530 22044
rect 2550 21998 2554 22044
rect 2574 21998 2578 22044
rect 2598 21998 2602 22044
rect 2622 21998 2626 22044
rect 2646 21998 2650 22044
rect 2670 21998 2674 22044
rect 2694 21998 2698 22044
rect 2718 21998 2722 22044
rect 2742 21998 2746 22044
rect 2766 21998 2770 22044
rect 2790 21998 2794 22044
rect 2814 21998 2818 22044
rect 2838 21998 2842 22044
rect 2875 22022 2909 22023
rect 3006 22022 3010 22044
rect 3030 22022 3034 22044
rect 3054 22022 3058 22044
rect 3078 22022 3082 22044
rect 3102 22022 3106 22044
rect 3109 22043 3123 22044
rect 3133 22044 3219 22046
rect 3133 22043 3147 22044
rect 3150 22043 3157 22044
rect 3174 22022 3178 22044
rect 3198 22022 3202 22044
rect 3205 22043 3219 22044
rect 3222 22043 3229 22067
rect 3222 22022 3226 22043
rect 3246 22022 3250 22068
rect 3270 22022 3274 22068
rect 3283 22061 3288 22068
rect 3325 22067 3339 22068
rect 3829 22067 3843 22068
rect 3293 22047 3298 22061
rect 3835 22057 3843 22061
rect 3829 22047 3835 22057
rect 3283 22037 3288 22047
rect 3302 22044 3317 22047
rect 3811 22046 3845 22047
rect 3846 22046 3853 22068
rect 3859 22061 3864 22068
rect 3877 22067 3891 22068
rect 4549 22067 4563 22068
rect 3869 22047 3874 22061
rect 3883 22057 3891 22061
rect 4555 22057 4563 22061
rect 3877 22047 3883 22057
rect 4549 22047 4555 22057
rect 3859 22046 3893 22047
rect 3811 22044 3893 22046
rect 4531 22046 4565 22047
rect 4566 22046 4573 22068
rect 4579 22061 4584 22068
rect 4597 22067 4611 22068
rect 4789 22067 4803 22068
rect 4589 22047 4594 22061
rect 4603 22057 4611 22061
rect 4795 22057 4803 22061
rect 4597 22047 4603 22057
rect 4789 22047 4795 22057
rect 4579 22046 4613 22047
rect 4531 22044 4613 22046
rect 4771 22046 4805 22047
rect 4806 22046 4813 22068
rect 4819 22061 4824 22068
rect 4837 22067 4851 22068
rect 4829 22047 4834 22061
rect 4843 22057 4851 22061
rect 4837 22047 4843 22057
rect 6557 22056 6565 22061
rect 6557 22048 6559 22056
rect 6557 22047 6565 22048
rect 4819 22046 4853 22047
rect 4771 22044 4853 22046
rect 6547 22046 6581 22047
rect 6582 22046 6586 22092
rect 6606 22070 6613 22091
rect 6630 22070 6634 22095
rect 6654 22091 6658 22115
rect 6589 22068 6651 22070
rect 6589 22067 6603 22068
rect 6606 22067 6613 22068
rect 6606 22046 6610 22067
rect 6630 22046 6634 22068
rect 6637 22067 6651 22068
rect 6654 22067 6661 22091
rect 6678 22046 6682 22116
rect 6702 22046 6706 22116
rect 6709 22115 6723 22116
rect 6726 22115 6733 22116
rect 6750 22094 6757 22115
rect 6774 22094 6778 22140
rect 6822 22118 6829 22139
rect 6846 22118 6850 22140
rect 6870 22118 6874 22140
rect 6894 22118 6898 22140
rect 6918 22118 6922 22140
rect 7027 22133 7032 22140
rect 7045 22139 7059 22140
rect 7037 22119 7042 22133
rect 7051 22129 7059 22133
rect 7045 22119 7051 22129
rect 7027 22118 7061 22119
rect 6805 22116 7061 22118
rect 7099 22116 7133 22119
rect 7147 22116 7181 22119
rect 10531 22118 10565 22119
rect 10566 22118 10573 22164
rect 10579 22157 10584 22164
rect 10597 22163 10611 22164
rect 11989 22163 12003 22164
rect 10589 22143 10594 22157
rect 10603 22153 10611 22157
rect 11995 22153 12003 22157
rect 10597 22143 10603 22153
rect 11989 22143 11995 22153
rect 10579 22118 10613 22119
rect 10531 22116 10613 22118
rect 11971 22118 12005 22119
rect 12006 22118 12013 22164
rect 12019 22157 12024 22164
rect 12037 22163 12051 22164
rect 12469 22163 12483 22164
rect 12029 22143 12034 22157
rect 12043 22153 12051 22157
rect 12475 22153 12483 22157
rect 12037 22143 12043 22153
rect 12469 22143 12475 22153
rect 12019 22118 12053 22119
rect 11971 22116 12053 22118
rect 12451 22118 12485 22119
rect 12486 22118 12493 22164
rect 12499 22157 12504 22164
rect 12517 22163 12531 22164
rect 12709 22163 12723 22164
rect 12509 22143 12514 22157
rect 12523 22153 12531 22157
rect 12715 22153 12723 22157
rect 12517 22143 12523 22153
rect 12709 22143 12715 22153
rect 12499 22118 12533 22119
rect 12451 22116 12533 22118
rect 12691 22118 12725 22119
rect 12726 22118 12733 22164
rect 12739 22157 12744 22164
rect 12757 22163 12771 22164
rect 13909 22163 13923 22164
rect 12749 22143 12754 22157
rect 12763 22153 12771 22157
rect 13915 22153 13923 22157
rect 12757 22143 12763 22153
rect 13909 22143 13915 22153
rect 12739 22118 12773 22119
rect 12691 22116 12773 22118
rect 13891 22118 13925 22119
rect 13926 22118 13933 22164
rect 13939 22157 13944 22164
rect 13957 22163 13971 22164
rect 13949 22143 13954 22157
rect 13963 22153 13971 22157
rect 13957 22143 13963 22153
rect 13939 22118 13973 22119
rect 13891 22116 13973 22118
rect 6805 22115 6819 22116
rect 6733 22092 6819 22094
rect 6726 22046 6730 22092
rect 6733 22091 6747 22092
rect 6750 22070 6757 22092
rect 6774 22070 6778 22092
rect 6805 22091 6819 22092
rect 6822 22091 6829 22116
rect 6846 22070 6850 22116
rect 6870 22070 6874 22116
rect 6894 22070 6898 22116
rect 6918 22070 6922 22116
rect 6942 22094 6949 22115
rect 7027 22109 7032 22116
rect 7045 22115 7059 22116
rect 10549 22115 10563 22116
rect 7037 22095 7042 22109
rect 7051 22105 7059 22109
rect 10555 22105 10563 22109
rect 7045 22095 7051 22105
rect 10549 22095 10555 22105
rect 7027 22094 7061 22095
rect 6925 22092 7061 22094
rect 7099 22092 7133 22095
rect 7147 22092 7181 22095
rect 10531 22094 10565 22095
rect 10566 22094 10573 22116
rect 10579 22109 10584 22116
rect 10597 22115 10611 22116
rect 11989 22115 12003 22116
rect 10589 22095 10594 22109
rect 10603 22105 10611 22109
rect 11995 22105 12003 22109
rect 10597 22095 10603 22105
rect 11989 22095 11995 22105
rect 10579 22094 10613 22095
rect 10531 22092 10613 22094
rect 6925 22091 6939 22092
rect 6942 22091 6949 22092
rect 6942 22070 6946 22091
rect 7027 22085 7032 22092
rect 7045 22091 7059 22092
rect 10549 22091 10563 22092
rect 7037 22071 7042 22085
rect 7051 22081 7059 22085
rect 10555 22081 10563 22085
rect 7045 22071 7051 22081
rect 10549 22071 10555 22081
rect 7027 22070 7061 22071
rect 6733 22068 7061 22070
rect 7099 22068 7133 22071
rect 7147 22068 7181 22071
rect 10531 22070 10565 22071
rect 10566 22070 10573 22092
rect 10579 22085 10584 22092
rect 10597 22091 10611 22092
rect 11989 22091 12003 22092
rect 12006 22091 12013 22116
rect 12019 22109 12024 22116
rect 12037 22115 12051 22116
rect 12469 22115 12483 22116
rect 12029 22095 12034 22109
rect 12043 22105 12051 22109
rect 12475 22105 12483 22109
rect 12037 22095 12043 22105
rect 12469 22095 12475 22105
rect 10589 22071 10594 22085
rect 10603 22081 10611 22085
rect 10597 22071 10603 22081
rect 10579 22070 10613 22071
rect 10531 22068 10613 22070
rect 6733 22067 6747 22068
rect 6750 22067 6757 22068
rect 6750 22046 6754 22067
rect 6774 22046 6778 22068
rect 6846 22046 6850 22068
rect 6870 22046 6874 22068
rect 6894 22046 6898 22068
rect 6918 22046 6922 22068
rect 6942 22046 6946 22068
rect 7027 22061 7032 22068
rect 7045 22067 7059 22068
rect 10549 22067 10563 22068
rect 10566 22067 10573 22068
rect 10579 22061 10584 22068
rect 10597 22067 10611 22068
rect 11989 22067 12003 22068
rect 12037 22067 12051 22068
rect 12469 22067 12483 22068
rect 12486 22067 12493 22116
rect 12499 22109 12504 22116
rect 12517 22115 12531 22116
rect 12709 22115 12723 22116
rect 12509 22095 12514 22109
rect 12523 22105 12531 22109
rect 12715 22105 12723 22109
rect 12517 22095 12523 22105
rect 12709 22095 12715 22105
rect 12726 22067 12733 22116
rect 12739 22109 12744 22116
rect 12757 22115 12771 22116
rect 13909 22115 13923 22116
rect 12749 22095 12754 22109
rect 12763 22105 12771 22109
rect 13915 22105 13923 22109
rect 12757 22095 12763 22105
rect 13909 22095 13915 22105
rect 13926 22067 13933 22116
rect 13939 22109 13944 22116
rect 13957 22115 13971 22116
rect 15619 22109 15624 22119
rect 13949 22095 13954 22109
rect 13963 22105 13971 22109
rect 13957 22095 13963 22105
rect 15629 22095 15634 22109
rect 7037 22047 7042 22061
rect 7051 22057 7059 22061
rect 7045 22047 7051 22057
rect 7157 22047 7162 22061
rect 10589 22047 10594 22061
rect 7027 22046 7061 22047
rect 6547 22044 7061 22046
rect 7099 22044 7133 22047
rect 3829 22043 3843 22044
rect 3293 22023 3298 22037
rect 3307 22033 3315 22037
rect 3835 22033 3843 22037
rect 3301 22023 3307 22033
rect 3829 22023 3835 22033
rect 3283 22022 3317 22023
rect 2875 22020 3317 22022
rect 3811 22022 3845 22023
rect 3846 22022 3853 22044
rect 3859 22037 3864 22044
rect 3877 22043 3891 22044
rect 4549 22043 4563 22044
rect 3869 22023 3874 22037
rect 3883 22033 3891 22037
rect 4555 22033 4563 22037
rect 3877 22023 3883 22033
rect 4549 22023 4555 22033
rect 3859 22022 3893 22023
rect 3811 22020 3893 22022
rect 4531 22022 4565 22023
rect 4566 22022 4573 22044
rect 4579 22037 4584 22044
rect 4597 22043 4611 22044
rect 4789 22043 4803 22044
rect 4589 22023 4594 22037
rect 4603 22033 4611 22037
rect 4795 22033 4803 22037
rect 4597 22023 4603 22033
rect 4789 22023 4795 22033
rect 4579 22022 4613 22023
rect 4531 22020 4613 22022
rect 4771 22022 4805 22023
rect 4806 22022 4813 22044
rect 4819 22037 4824 22044
rect 4837 22043 4851 22044
rect 6541 22043 6555 22044
rect 4829 22023 4834 22037
rect 4843 22033 4851 22037
rect 4837 22023 4843 22033
rect 4819 22022 4853 22023
rect 4771 22020 4853 22022
rect 6547 22020 6576 22023
rect 6582 22020 6586 22044
rect 2875 22013 2880 22020
rect 2885 21999 2890 22013
rect 2886 21998 2890 21999
rect 3006 21998 3010 22020
rect 3030 21998 3034 22020
rect 3054 21998 3058 22020
rect 3078 21998 3082 22020
rect 3102 21998 3106 22020
rect 3174 21998 3178 22020
rect 3198 21998 3202 22020
rect 3222 21998 3226 22020
rect 3246 21998 3250 22020
rect 3270 21998 3274 22020
rect 3283 22013 3288 22020
rect 3301 22019 3315 22020
rect 3829 22019 3843 22020
rect 3293 21999 3298 22013
rect 3307 22009 3315 22013
rect 3835 22009 3843 22013
rect 3301 21999 3307 22009
rect 3829 21999 3835 22009
rect 3283 21998 3317 21999
rect 2461 21996 3317 21998
rect 3811 21998 3845 21999
rect 3846 21998 3853 22020
rect 3859 22013 3864 22020
rect 3877 22019 3891 22020
rect 4549 22019 4563 22020
rect 3869 21999 3874 22013
rect 3883 22009 3891 22013
rect 4555 22009 4563 22013
rect 3877 21999 3883 22009
rect 4549 21999 4555 22009
rect 3859 21998 3893 21999
rect 3811 21996 3893 21998
rect 4531 21998 4565 21999
rect 4566 21998 4573 22020
rect 4579 22013 4584 22020
rect 4597 22019 4611 22020
rect 4789 22019 4803 22020
rect 4589 21999 4594 22013
rect 4603 22009 4611 22013
rect 4795 22009 4803 22013
rect 4597 21999 4603 22009
rect 4789 21999 4795 22009
rect 4579 21998 4613 21999
rect 4531 21996 4613 21998
rect 4771 21998 4805 21999
rect 4806 21998 4813 22020
rect 4819 22013 4824 22020
rect 4837 22019 4851 22020
rect 4829 21999 4834 22013
rect 4843 22009 4851 22013
rect 6571 22009 6579 22013
rect 4837 21999 4843 22009
rect 6565 21999 6571 22009
rect 4819 21998 4853 21999
rect 4771 21996 4853 21998
rect 6547 21998 6581 21999
rect 6582 21998 6589 22019
rect 6606 21998 6610 22044
rect 6630 21998 6634 22044
rect 6654 22022 6661 22043
rect 6678 22022 6682 22044
rect 6702 22022 6706 22044
rect 6726 22022 6730 22044
rect 6750 22022 6754 22044
rect 6774 22022 6778 22044
rect 6846 22022 6850 22044
rect 6870 22022 6874 22044
rect 6894 22022 6898 22044
rect 6918 22022 6922 22044
rect 6942 22022 6946 22044
rect 7027 22037 7032 22044
rect 7045 22043 7059 22044
rect 7037 22023 7042 22037
rect 7051 22033 7059 22037
rect 7123 22033 7131 22037
rect 7045 22023 7051 22033
rect 7117 22023 7123 22033
rect 7027 22022 7061 22023
rect 6637 22020 7061 22022
rect 7099 22022 7133 22023
rect 7134 22022 7141 22043
rect 7147 22037 7152 22047
rect 7157 22023 7162 22037
rect 7171 22033 7179 22037
rect 7165 22023 7171 22033
rect 7147 22022 7181 22023
rect 7099 22020 7181 22022
rect 12691 22022 12725 22023
rect 12726 22022 12733 22043
rect 12739 22022 12773 22023
rect 12691 22020 12773 22022
rect 6637 22019 6651 22020
rect 6654 22019 6661 22020
rect 6654 21998 6658 22019
rect 6678 21998 6682 22020
rect 6702 21998 6706 22020
rect 6726 21998 6730 22020
rect 6750 21998 6754 22020
rect 6774 21998 6778 22020
rect 6846 21998 6850 22020
rect 6870 21998 6874 22020
rect 6894 21998 6898 22020
rect 6918 21998 6922 22020
rect 6942 21998 6946 22020
rect 7027 22013 7032 22020
rect 7045 22019 7059 22020
rect 7117 22019 7131 22020
rect 7037 21999 7042 22013
rect 7051 22009 7059 22013
rect 7123 22009 7131 22013
rect 7045 21999 7051 22009
rect 7117 21999 7123 22009
rect 7027 21998 7061 21999
rect 6547 21996 7061 21998
rect 7099 21998 7133 21999
rect 7134 21998 7141 22020
rect 7147 22013 7152 22020
rect 7165 22019 7179 22020
rect 10549 22019 10563 22020
rect 10597 22019 10611 22020
rect 11989 22019 12003 22020
rect 12037 22019 12051 22020
rect 12469 22019 12483 22020
rect 12517 22019 12531 22020
rect 12709 22019 12723 22020
rect 12726 22019 12733 22020
rect 12739 22013 12744 22020
rect 12757 22019 12771 22020
rect 13909 22019 13923 22020
rect 13926 22019 13933 22043
rect 15606 22019 15613 22043
rect 7157 21999 7162 22013
rect 7171 22009 7179 22013
rect 7165 21999 7171 22009
rect 12749 21999 12754 22013
rect 7147 21998 7181 21999
rect 7099 21996 7181 21998
rect 2461 21995 2475 21996
rect 2478 21995 2485 21996
rect 2149 21972 2379 21974
rect 2149 21971 2163 21972
rect 2166 21971 2173 21972
rect 2131 21950 2165 21951
rect 2166 21950 2170 21971
rect 2190 21950 2194 21972
rect 2214 21950 2218 21972
rect 2262 21950 2266 21972
rect 2286 21950 2290 21972
rect 2310 21950 2314 21972
rect 2334 21950 2338 21972
rect 2365 21971 2379 21972
rect 2382 21971 2389 21995
rect 2478 21950 2482 21995
rect 2502 21950 2506 21996
rect 2526 21950 2530 21996
rect 2550 21950 2554 21996
rect 2574 21950 2578 21996
rect 2598 21950 2602 21996
rect 2622 21950 2626 21996
rect 2646 21950 2650 21996
rect 2670 21950 2674 21996
rect 2694 21950 2698 21996
rect 2718 21950 2722 21996
rect 2742 21950 2746 21996
rect 2766 21950 2770 21996
rect 2790 21950 2794 21996
rect 2814 21950 2818 21996
rect 2838 21950 2842 21996
rect 2862 21974 2869 21995
rect 2886 21974 2890 21996
rect 3006 21974 3010 21996
rect 3030 21974 3034 21996
rect 3054 21974 3058 21996
rect 3078 21974 3082 21996
rect 3102 21974 3106 21996
rect 3174 21974 3178 21996
rect 3198 21974 3202 21996
rect 3222 21974 3226 21996
rect 3246 21974 3250 21996
rect 3270 21974 3274 21996
rect 3283 21989 3288 21996
rect 3301 21995 3315 21996
rect 3829 21995 3843 21996
rect 3293 21975 3298 21989
rect 3307 21985 3315 21989
rect 3835 21985 3843 21989
rect 3301 21975 3307 21985
rect 3829 21975 3835 21985
rect 3283 21974 3317 21975
rect 2845 21972 3317 21974
rect 3811 21974 3845 21975
rect 3846 21974 3853 21996
rect 3859 21989 3864 21996
rect 3877 21995 3891 21996
rect 4549 21995 4563 21996
rect 3869 21975 3874 21989
rect 3883 21985 3891 21989
rect 4555 21985 4563 21989
rect 3877 21975 3883 21985
rect 4549 21975 4555 21985
rect 3859 21974 3893 21975
rect 3811 21972 3893 21974
rect 4531 21974 4565 21975
rect 4566 21974 4573 21996
rect 4579 21989 4584 21996
rect 4597 21995 4611 21996
rect 4789 21995 4803 21996
rect 4589 21975 4594 21989
rect 4603 21985 4611 21989
rect 4795 21985 4803 21989
rect 4597 21975 4603 21985
rect 4789 21975 4795 21985
rect 4579 21974 4613 21975
rect 4531 21972 4613 21974
rect 4771 21974 4805 21975
rect 4806 21974 4813 21996
rect 4819 21989 4824 21996
rect 4837 21995 4851 21996
rect 6565 21995 6579 21996
rect 4829 21975 4834 21989
rect 4843 21985 4851 21989
rect 6571 21985 6579 21989
rect 4837 21975 4843 21985
rect 6565 21975 6571 21985
rect 4819 21974 4853 21975
rect 4771 21972 4853 21974
rect 6547 21974 6581 21975
rect 6582 21974 6589 21996
rect 6606 21974 6610 21996
rect 6630 21974 6634 21996
rect 6654 21974 6658 21996
rect 6678 21974 6682 21996
rect 6702 21974 6706 21996
rect 6726 21974 6730 21996
rect 6750 21974 6754 21996
rect 6774 21974 6778 21996
rect 6846 21974 6850 21996
rect 6870 21974 6874 21996
rect 6894 21974 6898 21996
rect 6918 21974 6922 21996
rect 6942 21974 6946 21996
rect 7027 21989 7032 21996
rect 7045 21995 7059 21996
rect 7117 21995 7131 21996
rect 7037 21975 7042 21989
rect 7051 21985 7059 21989
rect 7123 21985 7131 21989
rect 7045 21975 7051 21985
rect 7117 21975 7123 21985
rect 7027 21974 7061 21975
rect 6547 21972 7061 21974
rect 7099 21974 7133 21975
rect 7134 21974 7141 21996
rect 7147 21989 7152 21996
rect 7165 21995 7179 21996
rect 10549 21995 10563 21996
rect 10597 21995 10611 21996
rect 7157 21975 7162 21989
rect 7171 21985 7179 21989
rect 7165 21975 7171 21985
rect 7147 21974 7181 21975
rect 7099 21972 7181 21974
rect 2845 21971 2859 21972
rect 2862 21971 2869 21972
rect 2862 21950 2866 21971
rect 2886 21950 2890 21972
rect 3006 21950 3010 21972
rect 3030 21950 3034 21972
rect 3054 21950 3058 21972
rect 3078 21950 3082 21972
rect 3102 21950 3106 21972
rect 3174 21950 3178 21972
rect 3198 21950 3202 21972
rect 3222 21950 3226 21972
rect 3246 21950 3250 21972
rect 3270 21950 3274 21972
rect 3283 21965 3288 21972
rect 3301 21971 3315 21972
rect 3829 21971 3843 21972
rect 3293 21951 3298 21965
rect 3307 21961 3315 21965
rect 3835 21961 3843 21965
rect 3301 21951 3307 21961
rect 3829 21951 3835 21961
rect 3283 21950 3317 21951
rect 2131 21948 3317 21950
rect 3811 21950 3845 21951
rect 3846 21950 3853 21972
rect 3859 21965 3864 21972
rect 3877 21971 3891 21972
rect 4549 21971 4563 21972
rect 3869 21951 3874 21965
rect 3883 21961 3891 21965
rect 4555 21961 4563 21965
rect 3877 21951 3883 21961
rect 4549 21951 4555 21961
rect 3859 21950 3893 21951
rect 3811 21948 3893 21950
rect 4531 21950 4565 21951
rect 4566 21950 4573 21972
rect 4579 21965 4584 21972
rect 4597 21971 4611 21972
rect 4789 21971 4803 21972
rect 4589 21951 4594 21965
rect 4603 21961 4611 21965
rect 4795 21961 4803 21965
rect 4597 21951 4603 21961
rect 4789 21951 4795 21961
rect 4579 21950 4613 21951
rect 4531 21948 4613 21950
rect 4771 21950 4805 21951
rect 4806 21950 4813 21972
rect 4819 21965 4824 21972
rect 4837 21971 4851 21972
rect 6565 21971 6579 21972
rect 4829 21951 4834 21965
rect 4843 21961 4851 21965
rect 6571 21961 6579 21965
rect 4837 21951 4843 21961
rect 6565 21951 6571 21961
rect 4819 21950 4853 21951
rect 4771 21948 4853 21950
rect 6547 21950 6581 21951
rect 6582 21950 6589 21972
rect 6606 21950 6610 21972
rect 6630 21950 6634 21972
rect 6654 21950 6658 21972
rect 6678 21950 6682 21972
rect 6702 21950 6706 21972
rect 6726 21950 6730 21972
rect 6750 21950 6754 21972
rect 6774 21950 6778 21972
rect 6846 21950 6850 21972
rect 6870 21950 6874 21972
rect 6894 21950 6898 21972
rect 6918 21950 6922 21972
rect 6942 21951 6946 21972
rect 7027 21965 7032 21972
rect 7045 21971 7059 21972
rect 7117 21971 7131 21972
rect 7037 21951 7042 21965
rect 7051 21961 7059 21965
rect 7123 21961 7131 21965
rect 7045 21951 7051 21961
rect 7117 21951 7123 21961
rect 6931 21950 6965 21951
rect 6547 21948 6965 21950
rect 6979 21950 7013 21951
rect 7027 21950 7061 21951
rect 6979 21948 7061 21950
rect 7099 21950 7133 21951
rect 7134 21950 7141 21972
rect 7147 21965 7152 21972
rect 7165 21971 7179 21972
rect 10549 21971 10563 21972
rect 10597 21971 10611 21972
rect 7157 21951 7162 21965
rect 7171 21961 7179 21965
rect 7165 21951 7171 21961
rect 7147 21950 7181 21951
rect 7099 21948 7181 21950
rect 2131 21941 2136 21948
rect 2166 21947 2170 21948
rect 2141 21927 2146 21941
rect 2155 21937 2163 21941
rect 2149 21927 2155 21937
rect 2142 21902 2146 21927
rect 2166 21923 2173 21947
rect 2190 21902 2194 21948
rect 2214 21902 2218 21948
rect 2238 21923 2245 21947
rect 2238 21902 2242 21923
rect 2262 21902 2266 21948
rect 2286 21902 2290 21948
rect 2310 21902 2314 21948
rect 2334 21902 2338 21948
rect 2478 21947 2482 21948
rect 2347 21926 2381 21927
rect 2347 21924 2475 21926
rect 2347 21917 2352 21924
rect 2461 21923 2475 21924
rect 2478 21923 2485 21947
rect 2357 21903 2362 21917
rect 2358 21902 2362 21903
rect 2502 21902 2506 21948
rect 2526 21902 2530 21948
rect 2550 21902 2554 21948
rect 2574 21902 2578 21948
rect 2598 21902 2602 21948
rect 2622 21902 2626 21948
rect 2646 21902 2650 21948
rect 2670 21902 2674 21948
rect 2694 21902 2698 21948
rect 2718 21902 2722 21948
rect 2742 21902 2746 21948
rect 2766 21902 2770 21948
rect 2790 21902 2794 21948
rect 2814 21902 2818 21948
rect 2838 21902 2842 21948
rect 2862 21902 2866 21948
rect 2886 21902 2890 21948
rect 2910 21926 2917 21947
rect 3006 21926 3010 21948
rect 3030 21926 3034 21948
rect 3054 21926 3058 21948
rect 3078 21926 3082 21948
rect 3102 21926 3106 21948
rect 3174 21926 3178 21948
rect 3198 21926 3202 21948
rect 3222 21926 3226 21948
rect 3246 21926 3250 21948
rect 3270 21926 3274 21948
rect 3283 21941 3288 21948
rect 3301 21947 3315 21948
rect 3829 21947 3843 21948
rect 3293 21927 3298 21941
rect 3307 21937 3315 21941
rect 3835 21937 3843 21941
rect 3301 21927 3307 21937
rect 3829 21927 3835 21937
rect 3283 21926 3317 21927
rect 2893 21924 3317 21926
rect 3811 21926 3845 21927
rect 3846 21926 3853 21948
rect 3859 21941 3864 21948
rect 3877 21947 3891 21948
rect 4549 21947 4563 21948
rect 3869 21927 3874 21941
rect 3883 21937 3891 21941
rect 4555 21937 4563 21941
rect 3877 21927 3883 21937
rect 4549 21927 4555 21937
rect 3859 21926 3893 21927
rect 3811 21924 3893 21926
rect 4531 21926 4565 21927
rect 4566 21926 4573 21948
rect 4579 21941 4584 21948
rect 4597 21947 4611 21948
rect 4789 21947 4803 21948
rect 4589 21927 4594 21941
rect 4603 21937 4611 21941
rect 4795 21937 4803 21941
rect 4597 21927 4603 21937
rect 4789 21927 4795 21937
rect 4579 21926 4613 21927
rect 4531 21924 4613 21926
rect 4771 21926 4805 21927
rect 4806 21926 4813 21948
rect 4819 21941 4824 21948
rect 4837 21947 4851 21948
rect 6565 21947 6579 21948
rect 4829 21927 4834 21941
rect 4843 21937 4851 21941
rect 6571 21937 6579 21941
rect 4837 21927 4843 21937
rect 6565 21927 6571 21937
rect 4819 21926 4853 21927
rect 4771 21924 4853 21926
rect 6547 21926 6581 21927
rect 6582 21926 6589 21948
rect 6606 21926 6610 21948
rect 6630 21926 6634 21948
rect 6654 21926 6658 21948
rect 6678 21927 6682 21948
rect 6667 21926 6701 21927
rect 6547 21924 6701 21926
rect 2893 21923 2907 21924
rect 2910 21923 2917 21924
rect 2910 21902 2914 21923
rect 3006 21902 3010 21924
rect 3030 21902 3034 21924
rect 3054 21902 3058 21924
rect 3078 21902 3082 21924
rect 3102 21902 3106 21924
rect 3174 21902 3178 21924
rect 3198 21902 3202 21924
rect 3222 21902 3226 21924
rect 3246 21902 3250 21924
rect 3270 21902 3274 21924
rect 3283 21917 3288 21924
rect 3301 21923 3315 21924
rect 3829 21923 3843 21924
rect 3293 21903 3298 21917
rect 3307 21913 3315 21917
rect 3835 21913 3843 21917
rect 3301 21903 3307 21913
rect 3829 21903 3835 21913
rect 3283 21902 3317 21903
rect 1405 21900 3317 21902
rect 3811 21902 3845 21903
rect 3846 21902 3853 21924
rect 3859 21917 3864 21924
rect 3877 21923 3891 21924
rect 4549 21923 4563 21924
rect 3869 21903 3874 21917
rect 3883 21913 3891 21917
rect 4555 21913 4563 21917
rect 3877 21903 3883 21913
rect 4549 21903 4555 21913
rect 3859 21902 3893 21903
rect 3811 21900 3893 21902
rect 4531 21902 4565 21903
rect 4566 21902 4573 21924
rect 4579 21917 4584 21924
rect 4597 21923 4611 21924
rect 4789 21923 4803 21924
rect 4589 21903 4594 21917
rect 4603 21913 4611 21917
rect 4795 21913 4803 21917
rect 4597 21903 4603 21913
rect 4789 21903 4795 21913
rect 4579 21902 4613 21903
rect 4531 21900 4613 21902
rect 4771 21902 4805 21903
rect 4806 21902 4813 21924
rect 4819 21917 4824 21924
rect 4837 21923 4851 21924
rect 6565 21923 6579 21924
rect 4829 21903 4834 21917
rect 4843 21913 4851 21917
rect 6571 21913 6579 21917
rect 4837 21903 4843 21913
rect 6565 21903 6571 21913
rect 4819 21902 4853 21903
rect 4771 21900 4853 21902
rect 6547 21902 6581 21903
rect 6582 21902 6589 21924
rect 6606 21902 6610 21924
rect 6630 21902 6634 21924
rect 6654 21903 6658 21924
rect 6667 21917 6672 21924
rect 6678 21917 6682 21924
rect 6677 21903 6682 21917
rect 6643 21902 6701 21903
rect 6702 21902 6706 21948
rect 6726 21902 6730 21948
rect 6750 21902 6754 21948
rect 6774 21902 6778 21948
rect 6787 21926 6821 21927
rect 6846 21926 6850 21948
rect 6870 21926 6874 21948
rect 6894 21926 6898 21948
rect 6918 21926 6922 21948
rect 6931 21941 6936 21948
rect 6942 21941 6946 21948
rect 6941 21927 6946 21941
rect 6956 21938 6960 21948
rect 7027 21941 7032 21948
rect 7045 21947 7059 21948
rect 7117 21947 7131 21948
rect 6931 21926 6965 21927
rect 6787 21924 6965 21926
rect 6787 21917 6792 21924
rect 6797 21903 6802 21917
rect 6787 21902 6821 21903
rect 6547 21900 6821 21902
rect 1325 21879 1330 21893
rect 1326 21878 1330 21879
rect 1350 21878 1354 21900
rect 1405 21899 1419 21900
rect 1422 21899 1429 21900
rect 1422 21878 1426 21899
rect 1446 21878 1450 21900
rect 1470 21878 1474 21900
rect 1494 21878 1498 21900
rect 1518 21878 1522 21900
rect 1542 21878 1546 21900
rect 1566 21878 1570 21900
rect 1590 21878 1594 21900
rect 1614 21878 1618 21900
rect 1638 21878 1642 21900
rect 1662 21878 1666 21900
rect 1686 21878 1690 21900
rect 1710 21878 1714 21900
rect 1734 21878 1738 21900
rect 1758 21878 1762 21900
rect 1782 21878 1786 21900
rect 1806 21878 1810 21900
rect 1830 21878 1834 21900
rect 1854 21878 1858 21900
rect 1878 21878 1882 21900
rect 1902 21878 1906 21900
rect 1926 21878 1930 21900
rect 1950 21878 1954 21900
rect 1974 21878 1978 21900
rect 2022 21878 2026 21900
rect 2046 21878 2050 21900
rect 2070 21878 2074 21900
rect 2094 21878 2098 21900
rect 2118 21878 2122 21900
rect 2142 21878 2146 21900
rect 2190 21878 2194 21900
rect 2214 21878 2218 21900
rect 2238 21878 2242 21900
rect 2262 21878 2266 21900
rect 2286 21878 2290 21900
rect 2310 21878 2314 21900
rect 2334 21878 2338 21900
rect 2358 21878 2362 21900
rect 2502 21878 2506 21900
rect 2526 21878 2530 21900
rect 2550 21878 2554 21900
rect 2574 21878 2578 21900
rect 2598 21878 2602 21900
rect 2622 21878 2626 21900
rect 2646 21878 2650 21900
rect 2670 21878 2674 21900
rect 2694 21878 2698 21900
rect 2718 21878 2722 21900
rect 2742 21878 2746 21900
rect 2766 21878 2770 21900
rect 2790 21878 2794 21900
rect 2814 21878 2818 21900
rect 2838 21878 2842 21900
rect 2862 21878 2866 21900
rect 2886 21878 2890 21900
rect 2910 21878 2914 21900
rect 3006 21878 3010 21900
rect 3030 21878 3034 21900
rect 3054 21878 3058 21900
rect 3078 21878 3082 21900
rect 3102 21878 3106 21900
rect 3174 21878 3178 21900
rect 3198 21878 3202 21900
rect 3222 21878 3226 21900
rect 3246 21878 3250 21900
rect 3270 21878 3274 21900
rect 3283 21893 3288 21900
rect 3301 21899 3315 21900
rect 3829 21899 3843 21900
rect 3293 21879 3298 21893
rect 3307 21889 3315 21893
rect 3835 21889 3843 21893
rect 3301 21879 3307 21889
rect 3829 21879 3835 21889
rect 3283 21878 3317 21879
rect -683 21876 3317 21878
rect 3811 21878 3845 21879
rect 3846 21878 3853 21900
rect 3859 21893 3864 21900
rect 3877 21899 3891 21900
rect 4549 21899 4563 21900
rect 3869 21879 3874 21893
rect 3883 21889 3891 21893
rect 4555 21889 4563 21893
rect 3877 21879 3883 21889
rect 4549 21879 4555 21889
rect 3859 21878 3893 21879
rect 3811 21876 3893 21878
rect 4531 21878 4565 21879
rect 4566 21878 4573 21900
rect 4579 21893 4584 21900
rect 4597 21899 4611 21900
rect 4789 21899 4803 21900
rect 4589 21879 4594 21893
rect 4603 21889 4611 21893
rect 4795 21889 4803 21893
rect 4597 21879 4603 21889
rect 4789 21879 4795 21889
rect 4579 21878 4613 21879
rect 4531 21876 4613 21878
rect 4771 21878 4805 21879
rect 4806 21878 4813 21900
rect 4819 21893 4824 21900
rect 4837 21899 4851 21900
rect 6565 21899 6579 21900
rect 4829 21879 4834 21893
rect 4843 21889 4851 21893
rect 6571 21889 6579 21893
rect 4837 21879 4843 21889
rect 6565 21879 6571 21889
rect 4819 21878 4853 21879
rect 4771 21876 4853 21878
rect 6547 21878 6581 21879
rect 6582 21878 6589 21900
rect 6606 21878 6610 21900
rect 6630 21878 6634 21900
rect 6643 21893 6648 21900
rect 6654 21893 6658 21900
rect 6667 21893 6672 21900
rect 6653 21879 6658 21893
rect 6677 21879 6682 21893
rect 6678 21878 6682 21879
rect 6702 21878 6706 21900
rect 6726 21879 6730 21900
rect 6715 21878 6749 21879
rect 6547 21876 6749 21878
rect -683 21875 -669 21876
rect -666 21875 -659 21876
rect -666 21854 -662 21875
rect -642 21854 -638 21876
rect -618 21854 -614 21876
rect -594 21854 -590 21876
rect -570 21854 -566 21876
rect -546 21854 -542 21876
rect -522 21854 -518 21876
rect -498 21854 -494 21876
rect -474 21854 -470 21876
rect -450 21854 -446 21876
rect -426 21854 -422 21876
rect -402 21854 -398 21876
rect -378 21854 -374 21876
rect -354 21854 -350 21876
rect -330 21854 -326 21876
rect -306 21854 -302 21876
rect -282 21854 -278 21876
rect -258 21854 -254 21876
rect -234 21854 -230 21876
rect -210 21854 -206 21876
rect -186 21854 -182 21876
rect -162 21854 -158 21876
rect -114 21854 -110 21876
rect -90 21854 -86 21876
rect -66 21854 -62 21876
rect -42 21854 -38 21876
rect -18 21854 -14 21876
rect -5 21854 29 21855
rect -2393 21852 29 21854
rect -2371 21830 -2366 21852
rect -2348 21830 -2343 21852
rect -2325 21830 -2320 21852
rect -2072 21850 -2036 21851
rect -2072 21844 -2054 21850
rect -2309 21836 -2301 21844
rect -2317 21830 -2309 21836
rect -2092 21835 -2062 21840
rect -2000 21831 -1992 21852
rect -1938 21851 -1906 21852
rect -1920 21850 -1906 21851
rect -1806 21844 -1680 21850
rect -1854 21835 -1806 21840
rect -1655 21836 -1647 21844
rect -1982 21831 -1966 21832
rect -2000 21830 -1966 21831
rect -1846 21830 -1806 21833
rect -1663 21830 -1655 21836
rect -1642 21830 -1637 21852
rect -1619 21830 -1614 21852
rect -1530 21830 -1526 21852
rect -1506 21830 -1502 21852
rect -1482 21830 -1478 21852
rect -1458 21830 -1454 21852
rect -1434 21830 -1430 21852
rect -1410 21830 -1406 21852
rect -1386 21830 -1382 21852
rect -1362 21830 -1358 21852
rect -1338 21830 -1334 21852
rect -1314 21830 -1310 21852
rect -1290 21830 -1286 21852
rect -1266 21830 -1262 21852
rect -1242 21830 -1238 21852
rect -1218 21830 -1214 21852
rect -1194 21830 -1190 21852
rect -1170 21830 -1166 21852
rect -1146 21830 -1142 21852
rect -1122 21830 -1118 21852
rect -1098 21830 -1094 21852
rect -1074 21830 -1070 21852
rect -1050 21830 -1046 21852
rect -1026 21830 -1022 21852
rect -1002 21830 -998 21852
rect -978 21830 -974 21852
rect -954 21830 -950 21852
rect -930 21830 -926 21852
rect -906 21830 -902 21852
rect -882 21831 -878 21852
rect -893 21830 -859 21831
rect -2393 21828 -859 21830
rect -2371 21806 -2366 21828
rect -2348 21806 -2343 21828
rect -2325 21806 -2320 21828
rect -2000 21826 -1966 21828
rect -2309 21808 -2301 21816
rect -2062 21815 -2054 21822
rect -2092 21808 -2084 21815
rect -2062 21808 -2026 21810
rect -2317 21806 -2309 21808
rect -2062 21806 -2012 21808
rect -2000 21806 -1992 21826
rect -1982 21825 -1966 21826
rect -1846 21824 -1806 21828
rect -1846 21817 -1798 21822
rect -1806 21815 -1798 21817
rect -1854 21813 -1846 21815
rect -1854 21808 -1806 21813
rect -1655 21808 -1647 21816
rect -1864 21806 -1796 21807
rect -1663 21806 -1655 21808
rect -1642 21806 -1637 21828
rect -1619 21806 -1614 21828
rect -1530 21806 -1526 21828
rect -1506 21806 -1502 21828
rect -1482 21806 -1478 21828
rect -1458 21806 -1454 21828
rect -1434 21806 -1430 21828
rect -1410 21806 -1406 21828
rect -1386 21806 -1382 21828
rect -1362 21806 -1358 21828
rect -1338 21806 -1334 21828
rect -1314 21806 -1310 21828
rect -1290 21806 -1286 21828
rect -1266 21806 -1262 21828
rect -1242 21806 -1238 21828
rect -1218 21806 -1214 21828
rect -1194 21807 -1190 21828
rect -1205 21806 -1171 21807
rect -1170 21806 -1166 21828
rect -1146 21806 -1142 21828
rect -1122 21806 -1118 21828
rect -1098 21806 -1094 21828
rect -1074 21806 -1070 21828
rect -1050 21806 -1046 21828
rect -1026 21806 -1022 21828
rect -1002 21827 -998 21828
rect -1002 21806 -995 21827
rect -978 21806 -974 21828
rect -954 21806 -950 21828
rect -930 21806 -926 21828
rect -906 21806 -902 21828
rect -893 21821 -888 21828
rect -882 21821 -878 21828
rect -883 21807 -878 21821
rect -882 21806 -878 21807
rect -858 21806 -854 21852
rect -834 21806 -830 21852
rect -810 21806 -806 21852
rect -786 21806 -782 21852
rect -762 21806 -758 21852
rect -738 21806 -734 21852
rect -714 21806 -710 21852
rect -690 21806 -686 21852
rect -666 21806 -662 21852
rect -642 21806 -638 21852
rect -618 21806 -614 21852
rect -594 21806 -590 21852
rect -570 21806 -566 21852
rect -546 21806 -542 21852
rect -522 21806 -518 21852
rect -498 21806 -494 21852
rect -474 21806 -470 21852
rect -450 21806 -446 21852
rect -426 21806 -422 21852
rect -402 21806 -398 21852
rect -378 21806 -374 21852
rect -354 21806 -350 21852
rect -330 21806 -326 21852
rect -306 21806 -302 21852
rect -282 21806 -278 21852
rect -258 21806 -254 21852
rect -234 21806 -230 21852
rect -210 21806 -206 21852
rect -186 21806 -182 21852
rect -162 21806 -158 21852
rect -114 21851 -110 21852
rect -149 21828 -117 21831
rect -149 21821 -144 21828
rect -131 21827 -117 21828
rect -114 21827 -107 21851
rect -139 21807 -134 21821
rect -138 21806 -134 21807
rect -90 21806 -86 21852
rect -66 21806 -62 21852
rect -42 21806 -38 21852
rect -18 21806 -14 21852
rect -5 21845 0 21852
rect 30 21851 34 21876
rect 5 21831 10 21845
rect 19 21841 27 21845
rect 13 21831 19 21841
rect 6 21806 10 21831
rect 30 21830 37 21851
rect 54 21830 58 21876
rect 78 21830 82 21876
rect 102 21830 106 21876
rect 126 21830 130 21876
rect 150 21830 154 21876
rect 174 21830 178 21876
rect 187 21854 221 21855
rect 246 21854 250 21876
rect 270 21854 274 21876
rect 294 21854 298 21876
rect 318 21854 322 21876
rect 342 21854 346 21876
rect 366 21854 370 21876
rect 390 21854 394 21876
rect 403 21854 437 21855
rect 187 21852 437 21854
rect 187 21845 192 21852
rect 197 21831 202 21845
rect 198 21830 202 21831
rect 246 21830 250 21852
rect 270 21830 274 21852
rect 294 21830 298 21852
rect 318 21830 322 21852
rect 342 21830 346 21852
rect 366 21830 370 21852
rect 390 21830 394 21852
rect 414 21845 421 21851
rect 413 21841 421 21845
rect 427 21841 435 21845
rect 413 21831 427 21841
rect 438 21830 445 21851
rect 462 21830 466 21876
rect 486 21830 490 21876
rect 510 21830 514 21876
rect 534 21830 538 21876
rect 558 21830 562 21876
rect 582 21830 586 21876
rect 606 21830 610 21876
rect 630 21830 634 21876
rect 654 21830 658 21876
rect 667 21854 701 21855
rect 726 21854 730 21876
rect 750 21854 754 21876
rect 774 21854 778 21876
rect 798 21854 802 21876
rect 822 21854 826 21876
rect 846 21854 850 21876
rect 870 21854 874 21876
rect 894 21854 898 21876
rect 942 21854 946 21876
rect 966 21854 970 21876
rect 990 21854 994 21876
rect 1014 21854 1018 21876
rect 1038 21854 1042 21876
rect 1062 21854 1066 21876
rect 1086 21854 1090 21876
rect 1110 21854 1114 21876
rect 1134 21854 1138 21876
rect 1158 21854 1162 21876
rect 1182 21854 1186 21876
rect 1206 21854 1210 21876
rect 1254 21854 1258 21876
rect 1278 21854 1282 21876
rect 1302 21854 1306 21876
rect 1326 21854 1330 21876
rect 1350 21854 1354 21876
rect 1422 21854 1426 21876
rect 1446 21854 1450 21876
rect 1470 21854 1474 21876
rect 1494 21854 1498 21876
rect 1518 21854 1522 21876
rect 1542 21854 1546 21876
rect 1566 21854 1570 21876
rect 1590 21854 1594 21876
rect 1614 21854 1618 21876
rect 1638 21854 1642 21876
rect 1662 21854 1666 21876
rect 1686 21854 1690 21876
rect 1710 21854 1714 21876
rect 1734 21854 1738 21876
rect 1758 21854 1762 21876
rect 1782 21854 1786 21876
rect 1806 21854 1810 21876
rect 1830 21854 1834 21876
rect 1854 21854 1858 21876
rect 1878 21854 1882 21876
rect 1902 21854 1906 21876
rect 1926 21854 1930 21876
rect 1950 21854 1954 21876
rect 1974 21854 1978 21876
rect 667 21852 1995 21854
rect 667 21845 672 21852
rect 677 21831 682 21845
rect 678 21830 682 21831
rect 726 21830 730 21852
rect 750 21830 754 21852
rect 774 21830 778 21852
rect 798 21830 802 21852
rect 822 21830 826 21852
rect 846 21830 850 21852
rect 870 21830 874 21852
rect 894 21830 898 21852
rect 942 21830 946 21852
rect 966 21830 970 21852
rect 990 21830 994 21852
rect 1014 21830 1018 21852
rect 1038 21830 1042 21852
rect 1062 21830 1066 21852
rect 1086 21830 1090 21852
rect 1110 21830 1114 21852
rect 1134 21830 1138 21852
rect 1158 21830 1162 21852
rect 1182 21830 1186 21852
rect 1206 21830 1210 21852
rect 1254 21830 1258 21852
rect 1278 21830 1282 21852
rect 1302 21830 1306 21852
rect 1326 21830 1330 21852
rect 1350 21851 1354 21852
rect 13 21828 411 21830
rect 13 21827 27 21828
rect 30 21827 37 21828
rect 54 21806 58 21828
rect 78 21806 82 21828
rect 102 21806 106 21828
rect 126 21806 130 21828
rect 150 21806 154 21828
rect 174 21806 178 21828
rect 198 21806 202 21828
rect 246 21806 250 21828
rect 270 21806 274 21828
rect 294 21806 298 21828
rect 318 21806 322 21828
rect 342 21806 346 21828
rect 366 21806 370 21828
rect 390 21806 394 21828
rect 397 21827 411 21828
rect 421 21828 1347 21830
rect 421 21827 435 21828
rect 438 21827 445 21828
rect 438 21806 442 21827
rect 462 21806 466 21828
rect 486 21806 490 21828
rect 510 21806 514 21828
rect 534 21806 538 21828
rect 558 21806 562 21828
rect 582 21806 586 21828
rect 606 21806 610 21828
rect 630 21806 634 21828
rect 654 21806 658 21828
rect 678 21806 682 21828
rect 726 21806 730 21828
rect 750 21806 754 21828
rect 774 21806 778 21828
rect 798 21806 802 21828
rect 822 21806 826 21828
rect 846 21806 850 21828
rect 870 21806 874 21828
rect 894 21806 898 21828
rect -2393 21804 915 21806
rect -2371 21758 -2366 21804
rect -2348 21758 -2343 21804
rect -2325 21758 -2320 21804
rect -2317 21800 -2309 21804
rect -2062 21800 -2054 21804
rect -2154 21796 -2138 21798
rect -2057 21796 -2054 21800
rect -2292 21790 -2054 21796
rect -2052 21790 -2044 21800
rect -2092 21774 -2062 21776
rect -2094 21770 -2062 21774
rect -2000 21758 -1992 21804
rect -1846 21797 -1806 21804
rect -1663 21800 -1655 21804
rect -1846 21790 -1680 21796
rect -1854 21774 -1806 21776
rect -1854 21770 -1680 21774
rect -1642 21758 -1637 21804
rect -1619 21758 -1614 21804
rect -1530 21758 -1526 21804
rect -1506 21758 -1502 21804
rect -1482 21758 -1478 21804
rect -1458 21758 -1454 21804
rect -1434 21758 -1430 21804
rect -1410 21758 -1406 21804
rect -1386 21758 -1382 21804
rect -1362 21758 -1358 21804
rect -1338 21758 -1334 21804
rect -1314 21758 -1310 21804
rect -1290 21758 -1286 21804
rect -1266 21758 -1262 21804
rect -1242 21758 -1238 21804
rect -1218 21758 -1214 21804
rect -1205 21797 -1200 21804
rect -1194 21797 -1190 21804
rect -1195 21783 -1190 21797
rect -1205 21773 -1200 21783
rect -1195 21759 -1190 21773
rect -1194 21758 -1190 21759
rect -1170 21758 -1166 21804
rect -1146 21758 -1142 21804
rect -1122 21758 -1118 21804
rect -1098 21758 -1094 21804
rect -1074 21758 -1070 21804
rect -1050 21758 -1046 21804
rect -1026 21758 -1022 21804
rect -1019 21803 -1005 21804
rect -1002 21782 -995 21804
rect -978 21782 -974 21804
rect -954 21782 -950 21804
rect -930 21782 -926 21804
rect -906 21782 -902 21804
rect -882 21782 -878 21804
rect -858 21782 -854 21804
rect -834 21782 -830 21804
rect -810 21782 -806 21804
rect -786 21782 -782 21804
rect -762 21782 -758 21804
rect -738 21782 -734 21804
rect -714 21782 -710 21804
rect -690 21782 -686 21804
rect -666 21782 -662 21804
rect -642 21782 -638 21804
rect -618 21782 -614 21804
rect -594 21782 -590 21804
rect -570 21782 -566 21804
rect -546 21782 -542 21804
rect -522 21782 -518 21804
rect -498 21782 -494 21804
rect -474 21782 -470 21804
rect -450 21782 -446 21804
rect -426 21782 -422 21804
rect -402 21782 -398 21804
rect -378 21782 -374 21804
rect -354 21782 -350 21804
rect -330 21782 -326 21804
rect -306 21782 -302 21804
rect -282 21782 -278 21804
rect -258 21782 -254 21804
rect -234 21782 -230 21804
rect -210 21782 -206 21804
rect -186 21782 -182 21804
rect -162 21782 -158 21804
rect -138 21782 -134 21804
rect -90 21782 -86 21804
rect -66 21782 -62 21804
rect -42 21782 -38 21804
rect -18 21782 -14 21804
rect 6 21782 10 21804
rect 54 21782 58 21804
rect 78 21782 82 21804
rect 102 21782 106 21804
rect 126 21782 130 21804
rect 150 21782 154 21804
rect 174 21782 178 21804
rect 198 21782 202 21804
rect 246 21782 250 21804
rect 270 21782 274 21804
rect 294 21782 298 21804
rect 318 21782 322 21804
rect 342 21782 346 21804
rect 366 21782 370 21804
rect 390 21782 394 21804
rect 438 21782 442 21804
rect 462 21782 466 21804
rect 486 21782 490 21804
rect 510 21782 514 21804
rect 534 21782 538 21804
rect 558 21782 562 21804
rect 582 21782 586 21804
rect 606 21782 610 21804
rect 630 21782 634 21804
rect 654 21782 658 21804
rect 678 21782 682 21804
rect 726 21782 730 21804
rect 750 21782 754 21804
rect 774 21782 778 21804
rect 798 21782 802 21804
rect 822 21782 826 21804
rect 846 21782 850 21804
rect 870 21782 874 21804
rect 894 21782 898 21804
rect 901 21803 915 21804
rect 918 21803 925 21827
rect 918 21782 922 21803
rect 942 21782 946 21828
rect 966 21782 970 21828
rect 990 21782 994 21828
rect 1014 21782 1018 21828
rect 1038 21782 1042 21828
rect 1062 21782 1066 21828
rect 1086 21782 1090 21828
rect 1110 21782 1114 21828
rect 1134 21782 1138 21828
rect 1158 21782 1162 21828
rect 1182 21782 1186 21828
rect 1206 21782 1210 21828
rect 1254 21827 1258 21828
rect 1254 21806 1261 21827
rect 1278 21806 1282 21828
rect 1302 21806 1306 21828
rect 1326 21806 1330 21828
rect 1333 21827 1347 21828
rect 1237 21804 1347 21806
rect 1237 21803 1251 21804
rect 1254 21803 1261 21804
rect 1278 21782 1282 21804
rect 1302 21782 1306 21804
rect 1326 21782 1330 21804
rect 1333 21803 1347 21804
rect 1350 21803 1357 21851
rect 1422 21828 1426 21852
rect 1350 21782 1354 21803
rect 1374 21782 1378 21828
rect 1422 21806 1429 21827
rect 1446 21806 1450 21852
rect 1470 21806 1474 21852
rect 1494 21806 1498 21852
rect 1518 21806 1522 21852
rect 1542 21806 1546 21852
rect 1566 21806 1570 21852
rect 1590 21806 1594 21852
rect 1614 21806 1618 21852
rect 1638 21806 1642 21852
rect 1662 21806 1666 21852
rect 1686 21806 1690 21852
rect 1710 21806 1714 21852
rect 1734 21806 1738 21852
rect 1758 21806 1762 21852
rect 1782 21806 1786 21852
rect 1806 21806 1810 21852
rect 1830 21806 1834 21852
rect 1854 21806 1858 21852
rect 1878 21806 1882 21852
rect 1902 21806 1906 21852
rect 1926 21806 1930 21852
rect 1950 21806 1954 21852
rect 1974 21806 1978 21852
rect 1981 21851 1995 21852
rect 1998 21851 2005 21875
rect 1998 21806 2002 21851
rect 2022 21806 2026 21876
rect 2046 21806 2050 21876
rect 2070 21806 2074 21876
rect 2094 21806 2098 21876
rect 2118 21806 2122 21876
rect 2142 21806 2146 21876
rect 2166 21854 2173 21875
rect 2190 21854 2194 21876
rect 2214 21854 2218 21876
rect 2238 21854 2242 21876
rect 2262 21854 2266 21876
rect 2286 21854 2290 21876
rect 2310 21854 2314 21876
rect 2334 21854 2338 21876
rect 2358 21854 2362 21876
rect 2502 21854 2506 21876
rect 2526 21854 2530 21876
rect 2550 21854 2554 21876
rect 2574 21854 2578 21876
rect 2598 21854 2602 21876
rect 2622 21854 2626 21876
rect 2646 21854 2650 21876
rect 2670 21854 2674 21876
rect 2694 21854 2698 21876
rect 2718 21854 2722 21876
rect 2742 21854 2746 21876
rect 2766 21854 2770 21876
rect 2790 21854 2794 21876
rect 2814 21854 2818 21876
rect 2838 21854 2842 21876
rect 2862 21854 2866 21876
rect 2886 21854 2890 21876
rect 2910 21854 2914 21876
rect 3006 21854 3010 21876
rect 3030 21854 3034 21876
rect 3054 21854 3058 21876
rect 3078 21854 3082 21876
rect 3102 21854 3106 21876
rect 3174 21854 3178 21876
rect 3198 21854 3202 21876
rect 3222 21854 3226 21876
rect 3246 21854 3250 21876
rect 3270 21854 3274 21876
rect 3283 21869 3288 21876
rect 3301 21875 3315 21876
rect 3829 21875 3843 21876
rect 3293 21855 3298 21869
rect 3307 21865 3315 21869
rect 3835 21865 3843 21869
rect 3301 21855 3307 21865
rect 3829 21855 3835 21865
rect 3283 21854 3317 21855
rect 2149 21852 3317 21854
rect 3811 21854 3845 21855
rect 3846 21854 3853 21876
rect 3859 21869 3864 21876
rect 3877 21875 3891 21876
rect 4549 21875 4563 21876
rect 3869 21855 3874 21869
rect 3883 21865 3891 21869
rect 4555 21865 4563 21869
rect 3877 21855 3883 21865
rect 4549 21855 4555 21865
rect 3859 21854 3893 21855
rect 3811 21852 3893 21854
rect 4531 21854 4565 21855
rect 4566 21854 4573 21876
rect 4579 21869 4584 21876
rect 4597 21875 4611 21876
rect 4789 21875 4803 21876
rect 4589 21855 4594 21869
rect 4603 21865 4611 21869
rect 4795 21865 4803 21869
rect 4597 21855 4603 21865
rect 4789 21855 4795 21865
rect 4579 21854 4613 21855
rect 4531 21852 4613 21854
rect 4771 21854 4805 21855
rect 4806 21854 4813 21876
rect 4819 21869 4824 21876
rect 4837 21875 4851 21876
rect 6565 21875 6579 21876
rect 4829 21855 4834 21869
rect 4843 21865 4851 21869
rect 6571 21865 6579 21869
rect 4837 21855 4843 21865
rect 6565 21855 6571 21865
rect 4819 21854 4853 21855
rect 4771 21852 4853 21854
rect 2149 21851 2163 21852
rect 2166 21851 2173 21852
rect 2166 21806 2170 21851
rect 2190 21806 2194 21852
rect 2214 21806 2218 21852
rect 2238 21806 2242 21852
rect 2262 21806 2266 21852
rect 2286 21806 2290 21852
rect 2310 21806 2314 21852
rect 2334 21806 2338 21852
rect 2358 21806 2362 21852
rect 2382 21830 2389 21851
rect 2502 21830 2506 21852
rect 2526 21830 2530 21852
rect 2550 21830 2554 21852
rect 2574 21830 2578 21852
rect 2598 21830 2602 21852
rect 2622 21830 2626 21852
rect 2646 21830 2650 21852
rect 2670 21830 2674 21852
rect 2694 21830 2698 21852
rect 2718 21830 2722 21852
rect 2742 21830 2746 21852
rect 2766 21830 2770 21852
rect 2790 21830 2794 21852
rect 2814 21830 2818 21852
rect 2838 21830 2842 21852
rect 2862 21830 2866 21852
rect 2886 21830 2890 21852
rect 2910 21830 2914 21852
rect 3006 21830 3010 21852
rect 3030 21830 3034 21852
rect 3054 21830 3058 21852
rect 3078 21830 3082 21852
rect 3102 21830 3106 21852
rect 3174 21830 3178 21852
rect 3198 21830 3202 21852
rect 3222 21830 3226 21852
rect 3246 21830 3250 21852
rect 3270 21830 3274 21852
rect 3283 21845 3288 21852
rect 3301 21851 3315 21852
rect 3829 21851 3843 21852
rect 3293 21831 3298 21845
rect 3307 21841 3315 21845
rect 3835 21841 3843 21845
rect 3301 21831 3307 21841
rect 3829 21831 3835 21841
rect 3283 21830 3317 21831
rect 2365 21828 3317 21830
rect 3811 21830 3845 21831
rect 3846 21830 3853 21852
rect 3859 21845 3864 21852
rect 3877 21851 3891 21852
rect 4549 21851 4563 21852
rect 3869 21831 3874 21845
rect 3883 21841 3891 21845
rect 4555 21841 4563 21845
rect 3877 21831 3883 21841
rect 4549 21831 4555 21841
rect 3859 21830 3893 21831
rect 3811 21828 3893 21830
rect 4531 21830 4565 21831
rect 4566 21830 4573 21852
rect 4579 21845 4584 21852
rect 4597 21851 4611 21852
rect 4789 21851 4803 21852
rect 4589 21831 4594 21845
rect 4603 21841 4611 21845
rect 4795 21841 4803 21845
rect 4597 21831 4603 21841
rect 4789 21831 4795 21841
rect 4579 21830 4613 21831
rect 4531 21828 4613 21830
rect 4771 21830 4805 21831
rect 4806 21830 4813 21852
rect 4819 21845 4824 21852
rect 4837 21851 4851 21852
rect 6565 21851 6579 21852
rect 6582 21851 6589 21876
rect 4829 21831 4834 21845
rect 4843 21841 4851 21845
rect 4837 21831 4843 21841
rect 4819 21830 4853 21831
rect 4771 21828 4853 21830
rect 6571 21830 6605 21831
rect 6606 21830 6610 21876
rect 6630 21830 6634 21876
rect 6644 21842 6648 21852
rect 6678 21842 6682 21876
rect 6702 21851 6706 21876
rect 6715 21869 6720 21876
rect 6726 21869 6730 21876
rect 6725 21855 6730 21869
rect 6715 21854 6749 21855
rect 6750 21854 6754 21900
rect 6774 21854 6778 21900
rect 6787 21893 6792 21900
rect 6798 21893 6802 21900
rect 6797 21879 6802 21893
rect 6787 21878 6821 21879
rect 6846 21878 6850 21924
rect 6870 21878 6874 21924
rect 6894 21878 6898 21924
rect 6918 21878 6922 21924
rect 6931 21917 6936 21924
rect 6941 21903 6946 21917
rect 6966 21914 6970 21938
rect 7037 21927 7042 21941
rect 7051 21937 7059 21941
rect 7123 21937 7131 21941
rect 7045 21927 7051 21937
rect 7117 21927 7123 21937
rect 6979 21926 7013 21927
rect 7027 21926 7061 21927
rect 6979 21924 7061 21926
rect 7027 21917 7032 21924
rect 7045 21923 7059 21924
rect 7117 21923 7130 21924
rect 7037 21903 7042 21917
rect 7051 21913 7059 21917
rect 7045 21903 7051 21913
rect 7134 21904 7141 21948
rect 7147 21941 7152 21948
rect 7165 21947 7179 21948
rect 7157 21927 7162 21941
rect 7171 21937 7179 21941
rect 7165 21927 7171 21937
rect 7165 21923 7179 21924
rect 6932 21890 6936 21900
rect 7028 21890 7032 21900
rect 7045 21899 7059 21900
rect 7120 21899 7131 21900
rect 7165 21899 7179 21900
rect 6942 21879 6946 21890
rect 6931 21878 6965 21879
rect 6787 21876 6965 21878
rect 6979 21878 7013 21879
rect 7038 21878 7042 21890
rect 6979 21876 7059 21878
rect 7099 21876 7133 21879
rect 7555 21876 7589 21879
rect 7603 21876 7637 21879
rect 6787 21869 6792 21876
rect 6797 21855 6802 21869
rect 6787 21854 6821 21855
rect 6715 21852 6821 21854
rect 6654 21831 6658 21842
rect 6643 21830 6699 21831
rect 6571 21828 6699 21830
rect 2365 21827 2379 21828
rect 2382 21827 2389 21828
rect 2382 21806 2386 21827
rect 2443 21806 2477 21807
rect 1405 21804 2477 21806
rect 1405 21803 1419 21804
rect 1422 21803 1429 21804
rect 1446 21782 1450 21804
rect 1470 21782 1474 21804
rect 1494 21782 1498 21804
rect 1518 21782 1522 21804
rect 1542 21782 1546 21804
rect 1566 21782 1570 21804
rect 1590 21782 1594 21804
rect 1614 21782 1618 21804
rect 1638 21782 1642 21804
rect 1662 21782 1666 21804
rect 1686 21782 1690 21804
rect 1710 21782 1714 21804
rect 1734 21782 1738 21804
rect 1758 21782 1762 21804
rect 1782 21782 1786 21804
rect 1806 21782 1810 21804
rect 1830 21782 1834 21804
rect 1854 21782 1858 21804
rect 1878 21782 1882 21804
rect 1902 21782 1906 21804
rect 1926 21782 1930 21804
rect 1950 21782 1954 21804
rect 1974 21782 1978 21804
rect 1998 21782 2002 21804
rect 2022 21782 2026 21804
rect 2046 21782 2050 21804
rect 2070 21782 2074 21804
rect 2094 21782 2098 21804
rect 2118 21782 2122 21804
rect 2142 21782 2146 21804
rect 2166 21782 2170 21804
rect 2190 21782 2194 21804
rect 2214 21782 2218 21804
rect 2238 21782 2242 21804
rect 2262 21782 2266 21804
rect 2286 21782 2290 21804
rect 2310 21782 2314 21804
rect 2334 21782 2338 21804
rect 2358 21782 2362 21804
rect 2382 21782 2386 21804
rect 2443 21797 2448 21804
rect 2453 21783 2458 21797
rect 2454 21782 2458 21783
rect 2502 21782 2506 21828
rect 2526 21782 2530 21828
rect 2550 21782 2554 21828
rect 2574 21782 2578 21828
rect 2598 21782 2602 21828
rect 2622 21782 2626 21828
rect 2646 21782 2650 21828
rect 2670 21782 2674 21828
rect 2694 21807 2698 21828
rect 2683 21806 2717 21807
rect 2718 21806 2722 21828
rect 2742 21806 2746 21828
rect 2766 21806 2770 21828
rect 2790 21806 2794 21828
rect 2814 21806 2818 21828
rect 2838 21806 2842 21828
rect 2862 21806 2866 21828
rect 2886 21806 2890 21828
rect 2910 21806 2914 21828
rect 2923 21806 2981 21807
rect 3006 21806 3010 21828
rect 3030 21806 3034 21828
rect 3054 21806 3058 21828
rect 3078 21806 3082 21828
rect 3102 21806 3106 21828
rect 3174 21806 3178 21828
rect 3198 21806 3202 21828
rect 3222 21806 3226 21828
rect 3246 21806 3250 21828
rect 3270 21806 3274 21828
rect 3283 21821 3288 21828
rect 3301 21827 3315 21828
rect 3829 21827 3843 21828
rect 3293 21807 3298 21821
rect 3307 21817 3315 21821
rect 3835 21817 3843 21821
rect 3301 21807 3307 21817
rect 3829 21807 3835 21817
rect 3283 21806 3317 21807
rect 2683 21804 3317 21806
rect 3811 21806 3845 21807
rect 3846 21806 3853 21828
rect 3859 21821 3864 21828
rect 3877 21827 3891 21828
rect 4549 21827 4563 21828
rect 3869 21807 3874 21821
rect 3883 21817 3891 21821
rect 4555 21817 4563 21821
rect 3877 21807 3883 21817
rect 4549 21807 4555 21817
rect 3859 21806 3893 21807
rect 3811 21804 3893 21806
rect 4531 21806 4565 21807
rect 4566 21806 4573 21828
rect 4579 21821 4584 21828
rect 4597 21827 4611 21828
rect 4789 21827 4803 21828
rect 4589 21807 4594 21821
rect 4603 21817 4611 21821
rect 4795 21817 4803 21821
rect 4597 21807 4603 21817
rect 4789 21807 4795 21817
rect 4579 21806 4613 21807
rect 4531 21804 4613 21806
rect 4771 21806 4805 21807
rect 4806 21806 4813 21828
rect 4819 21821 4824 21828
rect 4837 21827 4851 21828
rect 6565 21827 6579 21828
rect 4829 21807 4834 21821
rect 4843 21817 4851 21821
rect 4837 21807 4843 21817
rect 6581 21816 6589 21821
rect 6581 21808 6583 21816
rect 6581 21807 6589 21808
rect 4819 21806 4853 21807
rect 4771 21804 4853 21806
rect 6571 21806 6605 21807
rect 6606 21806 6610 21828
rect 6630 21807 6634 21828
rect 6643 21821 6648 21828
rect 6654 21821 6658 21828
rect 6653 21807 6658 21821
rect 6667 21821 6672 21828
rect 6685 21827 6699 21828
rect 6667 21817 6675 21821
rect 6677 21817 6685 21821
rect 6691 21817 6699 21821
rect 6661 21807 6667 21817
rect 6677 21807 6691 21817
rect 6619 21806 6653 21807
rect 6571 21804 6653 21806
rect 2683 21797 2688 21804
rect 2694 21797 2698 21804
rect 2693 21783 2698 21797
rect 2718 21782 2722 21804
rect 2742 21782 2746 21804
rect 2766 21782 2770 21804
rect 2790 21782 2794 21804
rect 2814 21782 2818 21804
rect 2838 21782 2842 21804
rect 2862 21782 2866 21804
rect 2886 21782 2890 21804
rect 2910 21782 2914 21804
rect 2923 21797 2928 21804
rect 2933 21783 2938 21797
rect 2934 21782 2938 21783
rect 3006 21782 3010 21804
rect 3030 21782 3034 21804
rect 3054 21782 3058 21804
rect 3078 21782 3082 21804
rect 3102 21782 3106 21804
rect 3174 21782 3178 21804
rect 3198 21782 3202 21804
rect 3222 21782 3226 21804
rect 3246 21782 3250 21804
rect 3270 21782 3274 21804
rect 3283 21797 3288 21804
rect 3301 21803 3315 21804
rect 3829 21803 3843 21804
rect 3293 21783 3298 21797
rect 3307 21793 3315 21797
rect 3835 21793 3843 21797
rect 3301 21783 3307 21793
rect 3829 21783 3835 21793
rect 3283 21782 3317 21783
rect -1019 21780 3317 21782
rect 3811 21782 3845 21783
rect 3846 21782 3853 21804
rect 3859 21797 3864 21804
rect 3877 21803 3891 21804
rect 4549 21803 4563 21804
rect 3869 21783 3874 21797
rect 3883 21793 3891 21797
rect 4555 21793 4563 21797
rect 3877 21783 3883 21793
rect 4549 21783 4555 21793
rect 3859 21782 3893 21783
rect 3811 21780 3893 21782
rect 4531 21782 4565 21783
rect 4566 21782 4573 21804
rect 4579 21797 4584 21804
rect 4597 21803 4611 21804
rect 4789 21803 4803 21804
rect 4589 21783 4594 21797
rect 4603 21793 4611 21797
rect 4795 21793 4803 21797
rect 4597 21783 4603 21793
rect 4789 21783 4795 21793
rect 4579 21782 4613 21783
rect 4531 21780 4613 21782
rect 4771 21782 4805 21783
rect 4806 21782 4813 21804
rect 4819 21797 4824 21804
rect 4837 21803 4851 21804
rect 6565 21803 6579 21804
rect 4829 21783 4834 21797
rect 4843 21793 4851 21797
rect 4837 21783 4843 21793
rect 6581 21792 6589 21797
rect 6581 21784 6583 21792
rect 6581 21783 6589 21784
rect 4819 21782 4853 21783
rect 4771 21780 4853 21782
rect 6571 21782 6605 21783
rect 6606 21782 6610 21804
rect 6619 21797 6624 21804
rect 6630 21797 6634 21804
rect 6629 21783 6634 21797
rect 6644 21794 6648 21804
rect 6661 21803 6675 21804
rect 6678 21803 6685 21807
rect 6702 21803 6709 21851
rect 6715 21845 6720 21852
rect 6725 21831 6730 21845
rect 6715 21821 6720 21831
rect 6726 21821 6730 21831
rect 6725 21807 6730 21821
rect 6715 21806 6749 21807
rect 6750 21806 6754 21852
rect 6774 21806 6778 21852
rect 6787 21845 6792 21852
rect 6798 21845 6802 21852
rect 6797 21831 6802 21845
rect 6811 21841 6819 21845
rect 6805 21831 6811 21841
rect 6787 21821 6792 21831
rect 6805 21830 6821 21831
rect 6822 21830 6829 21851
rect 6846 21830 6850 21876
rect 6870 21830 6874 21876
rect 6894 21830 6898 21876
rect 6918 21830 6922 21876
rect 6931 21869 6936 21876
rect 6942 21869 6946 21876
rect 6956 21869 6960 21876
rect 6941 21855 6946 21869
rect 6955 21865 6963 21869
rect 6949 21855 6955 21865
rect 6931 21852 6963 21855
rect 6931 21845 6936 21852
rect 6949 21851 6963 21852
rect 6941 21831 6946 21845
rect 6955 21841 6963 21845
rect 6949 21831 6955 21841
rect 6966 21838 6973 21866
rect 7003 21865 7011 21869
rect 6997 21855 7003 21865
rect 7014 21854 7021 21875
rect 7038 21854 7042 21876
rect 7045 21875 7059 21876
rect 7117 21875 7131 21876
rect 7165 21875 7179 21876
rect 7123 21865 7131 21869
rect 7117 21855 7123 21865
rect 6997 21852 7059 21854
rect 7099 21852 7133 21855
rect 8251 21852 8285 21855
rect 8299 21852 8333 21855
rect 6997 21851 7011 21852
rect 6942 21830 6946 21831
rect 7014 21830 7021 21852
rect 7038 21830 7042 21852
rect 7045 21851 7059 21852
rect 7117 21851 7131 21852
rect 7165 21851 7179 21852
rect 6805 21828 6963 21830
rect 6997 21828 7059 21830
rect 7099 21828 7118 21831
rect 6805 21827 6819 21828
rect 6797 21807 6802 21821
rect 6811 21817 6819 21821
rect 6805 21807 6811 21817
rect 6798 21806 6802 21807
rect 6715 21804 6819 21806
rect 6619 21782 6653 21783
rect 6571 21780 6653 21782
rect -1019 21779 -1005 21780
rect -1002 21779 -995 21780
rect -1002 21758 -998 21779
rect -978 21758 -974 21780
rect -954 21758 -950 21780
rect -930 21758 -926 21780
rect -906 21758 -902 21780
rect -882 21758 -878 21780
rect -858 21758 -854 21780
rect -834 21758 -830 21780
rect -810 21758 -806 21780
rect -786 21758 -782 21780
rect -762 21758 -758 21780
rect -738 21758 -734 21780
rect -714 21758 -710 21780
rect -690 21758 -686 21780
rect -666 21758 -662 21780
rect -642 21758 -638 21780
rect -618 21758 -614 21780
rect -594 21758 -590 21780
rect -570 21758 -566 21780
rect -546 21758 -542 21780
rect -522 21758 -518 21780
rect -498 21758 -494 21780
rect -474 21758 -470 21780
rect -450 21758 -446 21780
rect -426 21758 -422 21780
rect -402 21758 -398 21780
rect -378 21758 -374 21780
rect -354 21758 -350 21780
rect -330 21758 -326 21780
rect -306 21758 -302 21780
rect -282 21758 -278 21780
rect -258 21758 -254 21780
rect -234 21758 -230 21780
rect -210 21758 -206 21780
rect -186 21758 -182 21780
rect -162 21758 -158 21780
rect -138 21758 -134 21780
rect -90 21758 -86 21780
rect -66 21758 -62 21780
rect -42 21758 -38 21780
rect -18 21758 -14 21780
rect 6 21758 10 21780
rect -2393 21756 27 21758
rect -2371 21710 -2366 21756
rect -2348 21710 -2343 21756
rect -2325 21710 -2320 21756
rect -2309 21740 -2301 21750
rect -2317 21734 -2309 21740
rect -2097 21734 -2095 21743
rect -2309 21712 -2301 21722
rect -2097 21720 -2095 21724
rect -2292 21719 -2095 21720
rect -2097 21717 -2095 21719
rect -2084 21712 -2083 21755
rect -2069 21748 -2054 21750
rect -2054 21732 -2018 21734
rect -2054 21730 -2004 21732
rect -2059 21726 -2045 21730
rect -2054 21724 -2049 21726
rect -2317 21710 -2309 21712
rect -2084 21710 -2054 21712
rect -2044 21710 -2039 21724
rect -2025 21714 -2014 21720
rect -2000 21714 -1992 21756
rect -1920 21754 -1906 21756
rect -1977 21739 -1929 21745
rect -1655 21740 -1647 21750
rect -1977 21729 -1966 21739
rect -1663 21734 -1655 21740
rect -1977 21717 -1929 21719
rect -2033 21710 -1992 21714
rect -1655 21712 -1647 21722
rect -1663 21710 -1655 21712
rect -1642 21710 -1637 21756
rect -1619 21710 -1614 21756
rect -1530 21710 -1526 21756
rect -1506 21710 -1502 21756
rect -1482 21710 -1478 21756
rect -1458 21710 -1454 21756
rect -1434 21710 -1430 21756
rect -1410 21710 -1406 21756
rect -1386 21710 -1382 21756
rect -1362 21710 -1358 21756
rect -1338 21710 -1334 21756
rect -1314 21710 -1310 21756
rect -1290 21710 -1286 21756
rect -1266 21710 -1262 21756
rect -1242 21710 -1238 21756
rect -1218 21710 -1214 21756
rect -1194 21710 -1190 21756
rect -1170 21731 -1166 21756
rect -1170 21710 -1163 21731
rect -1146 21710 -1142 21756
rect -1122 21710 -1118 21756
rect -1098 21710 -1094 21756
rect -1074 21710 -1070 21756
rect -1050 21710 -1046 21756
rect -1026 21710 -1022 21756
rect -1002 21710 -998 21756
rect -978 21710 -974 21756
rect -954 21710 -950 21756
rect -930 21710 -926 21756
rect -906 21710 -902 21756
rect -882 21710 -878 21756
rect -858 21755 -854 21756
rect -858 21731 -851 21755
rect -858 21710 -854 21731
rect -834 21710 -830 21756
rect -810 21710 -806 21756
rect -786 21710 -782 21756
rect -762 21710 -758 21756
rect -738 21710 -734 21756
rect -714 21710 -710 21756
rect -690 21710 -686 21756
rect -666 21710 -662 21756
rect -642 21710 -638 21756
rect -618 21710 -614 21756
rect -594 21710 -590 21756
rect -570 21710 -566 21756
rect -546 21710 -542 21756
rect -522 21710 -518 21756
rect -498 21710 -494 21756
rect -474 21710 -470 21756
rect -450 21710 -446 21756
rect -426 21710 -422 21756
rect -402 21710 -398 21756
rect -378 21711 -374 21756
rect -389 21710 -355 21711
rect -2393 21708 -355 21710
rect -2371 21614 -2366 21708
rect -2348 21614 -2343 21708
rect -2325 21674 -2320 21708
rect -2317 21706 -2309 21708
rect -2084 21695 -2083 21708
rect -2084 21694 -2054 21695
rect -2325 21666 -2317 21674
rect -2325 21646 -2320 21666
rect -2317 21658 -2309 21666
rect -2117 21657 -2095 21667
rect -2045 21664 -2037 21678
rect -2325 21632 -2317 21646
rect -2325 21616 -2320 21632
rect -2317 21630 -2309 21632
rect -2309 21618 -2301 21630
rect -2109 21629 -2079 21630
rect -2317 21616 -2309 21618
rect -2325 21614 -2317 21616
rect -2109 21615 -2087 21629
rect -2015 21616 -2001 21621
rect -2000 21616 -1992 21708
rect -1663 21706 -1655 21708
rect -1969 21657 -1929 21669
rect -1671 21666 -1663 21674
rect -1663 21658 -1655 21666
rect -1671 21632 -1663 21646
rect -1663 21630 -1655 21632
rect -1655 21618 -1647 21630
rect -1663 21616 -1655 21618
rect -2109 21614 -2079 21615
rect -2033 21614 -1992 21616
rect -1864 21614 -1680 21615
rect -1671 21614 -1663 21616
rect -1642 21614 -1637 21708
rect -1619 21614 -1614 21708
rect -1530 21614 -1526 21708
rect -1506 21614 -1502 21708
rect -1482 21614 -1478 21708
rect -1458 21614 -1454 21708
rect -1434 21614 -1430 21708
rect -1410 21614 -1406 21708
rect -1386 21614 -1382 21708
rect -1362 21614 -1358 21708
rect -1338 21614 -1334 21708
rect -1314 21614 -1310 21708
rect -1290 21614 -1286 21708
rect -1266 21614 -1262 21708
rect -1242 21614 -1238 21708
rect -1218 21614 -1214 21708
rect -1194 21614 -1190 21708
rect -1187 21707 -1173 21708
rect -1170 21686 -1163 21708
rect -1146 21686 -1142 21708
rect -1122 21686 -1118 21708
rect -1098 21687 -1094 21708
rect -1109 21686 -1075 21687
rect -1187 21684 -1075 21686
rect -1187 21683 -1173 21684
rect -1170 21683 -1163 21684
rect -1170 21614 -1166 21683
rect -1146 21614 -1142 21684
rect -1122 21614 -1118 21684
rect -1109 21677 -1104 21684
rect -1098 21677 -1094 21684
rect -1099 21663 -1094 21677
rect -1109 21662 -1075 21663
rect -1074 21662 -1070 21708
rect -1050 21662 -1046 21708
rect -1026 21662 -1022 21708
rect -1002 21662 -998 21708
rect -978 21662 -974 21708
rect -954 21662 -950 21708
rect -930 21662 -926 21708
rect -906 21662 -902 21708
rect -882 21662 -878 21708
rect -858 21662 -854 21708
rect -834 21662 -830 21708
rect -810 21662 -806 21708
rect -786 21662 -782 21708
rect -762 21662 -758 21708
rect -738 21662 -734 21708
rect -714 21662 -710 21708
rect -690 21662 -686 21708
rect -666 21662 -662 21708
rect -642 21662 -638 21708
rect -618 21662 -614 21708
rect -594 21662 -590 21708
rect -570 21662 -566 21708
rect -546 21662 -542 21708
rect -522 21662 -518 21708
rect -498 21662 -494 21708
rect -474 21662 -470 21708
rect -450 21662 -446 21708
rect -426 21662 -422 21708
rect -402 21662 -398 21708
rect -389 21701 -384 21708
rect -378 21701 -374 21708
rect -379 21687 -374 21701
rect -389 21686 -355 21687
rect -354 21686 -350 21756
rect -330 21686 -326 21756
rect -306 21686 -302 21756
rect -282 21686 -278 21756
rect -258 21686 -254 21756
rect -234 21686 -230 21756
rect -210 21686 -206 21756
rect -186 21686 -182 21756
rect -162 21686 -158 21756
rect -138 21686 -134 21756
rect -114 21731 -107 21755
rect -114 21686 -110 21731
rect -90 21686 -86 21756
rect -66 21686 -62 21756
rect -42 21686 -38 21756
rect -18 21686 -14 21756
rect 6 21686 10 21756
rect 13 21755 27 21756
rect 30 21755 37 21779
rect 30 21686 34 21755
rect 54 21686 58 21780
rect 78 21686 82 21780
rect 102 21686 106 21780
rect 126 21686 130 21780
rect 150 21686 154 21780
rect 174 21686 178 21780
rect 198 21686 202 21780
rect 222 21758 229 21779
rect 246 21758 250 21780
rect 270 21758 274 21780
rect 294 21758 298 21780
rect 318 21758 322 21780
rect 342 21758 346 21780
rect 366 21758 370 21780
rect 390 21758 394 21780
rect 438 21779 442 21780
rect 205 21756 435 21758
rect 205 21755 219 21756
rect 222 21755 229 21756
rect 222 21686 226 21755
rect 246 21686 250 21756
rect 270 21686 274 21756
rect 294 21686 298 21756
rect 318 21686 322 21756
rect 342 21686 346 21756
rect 366 21686 370 21756
rect 390 21686 394 21756
rect 421 21755 435 21756
rect 438 21755 445 21779
rect 403 21734 437 21735
rect 462 21734 466 21780
rect 486 21734 490 21780
rect 510 21734 514 21780
rect 534 21734 538 21780
rect 558 21734 562 21780
rect 582 21734 586 21780
rect 606 21734 610 21780
rect 630 21734 634 21780
rect 654 21734 658 21780
rect 678 21734 682 21780
rect 702 21758 709 21779
rect 726 21758 730 21780
rect 750 21758 754 21780
rect 774 21758 778 21780
rect 798 21758 802 21780
rect 822 21758 826 21780
rect 846 21758 850 21780
rect 870 21758 874 21780
rect 894 21758 898 21780
rect 918 21758 922 21780
rect 942 21758 946 21780
rect 966 21758 970 21780
rect 990 21758 994 21780
rect 1014 21758 1018 21780
rect 1038 21758 1042 21780
rect 1062 21758 1066 21780
rect 1086 21758 1090 21780
rect 1110 21758 1114 21780
rect 1134 21758 1138 21780
rect 1158 21758 1162 21780
rect 1182 21758 1186 21780
rect 1206 21758 1210 21780
rect 1278 21758 1282 21780
rect 1302 21758 1306 21780
rect 1326 21758 1330 21780
rect 1350 21758 1354 21780
rect 1374 21758 1378 21780
rect 1446 21758 1450 21780
rect 1470 21758 1474 21780
rect 1494 21758 1498 21780
rect 1518 21758 1522 21780
rect 1542 21758 1546 21780
rect 1566 21758 1570 21780
rect 1590 21758 1594 21780
rect 1614 21758 1618 21780
rect 1638 21758 1642 21780
rect 1662 21758 1666 21780
rect 1686 21758 1690 21780
rect 1710 21758 1714 21780
rect 1734 21758 1738 21780
rect 1758 21758 1762 21780
rect 1782 21758 1786 21780
rect 1806 21758 1810 21780
rect 1830 21758 1834 21780
rect 1854 21758 1858 21780
rect 1878 21758 1882 21780
rect 1902 21758 1906 21780
rect 1926 21758 1930 21780
rect 1950 21758 1954 21780
rect 1974 21758 1978 21780
rect 1998 21758 2002 21780
rect 2022 21758 2026 21780
rect 2046 21758 2050 21780
rect 2070 21758 2074 21780
rect 2094 21758 2098 21780
rect 2118 21758 2122 21780
rect 2142 21758 2146 21780
rect 2166 21758 2170 21780
rect 2190 21758 2194 21780
rect 2214 21758 2218 21780
rect 2238 21758 2242 21780
rect 2262 21758 2266 21780
rect 2286 21758 2290 21780
rect 2310 21758 2314 21780
rect 2334 21758 2338 21780
rect 2358 21758 2362 21780
rect 2382 21758 2386 21780
rect 2395 21758 2429 21759
rect 685 21756 2429 21758
rect 685 21755 699 21756
rect 702 21755 709 21756
rect 702 21734 706 21755
rect 726 21734 730 21756
rect 750 21734 754 21756
rect 774 21734 778 21756
rect 798 21734 802 21756
rect 822 21734 826 21756
rect 846 21734 850 21756
rect 870 21734 874 21756
rect 894 21734 898 21756
rect 918 21734 922 21756
rect 942 21734 946 21756
rect 966 21734 970 21756
rect 990 21734 994 21756
rect 1014 21734 1018 21756
rect 1038 21734 1042 21756
rect 1062 21734 1066 21756
rect 1086 21734 1090 21756
rect 1110 21734 1114 21756
rect 1134 21734 1138 21756
rect 1158 21734 1162 21756
rect 1182 21734 1186 21756
rect 1206 21734 1210 21756
rect 1278 21734 1282 21756
rect 1302 21734 1306 21756
rect 1326 21734 1330 21756
rect 1350 21734 1354 21756
rect 1374 21734 1378 21756
rect 1446 21734 1450 21756
rect 1470 21734 1474 21756
rect 1494 21734 1498 21756
rect 1518 21734 1522 21756
rect 1542 21734 1546 21756
rect 1566 21734 1570 21756
rect 1590 21734 1594 21756
rect 1614 21734 1618 21756
rect 1638 21734 1642 21756
rect 1662 21734 1666 21756
rect 1686 21734 1690 21756
rect 1710 21734 1714 21756
rect 1734 21734 1738 21756
rect 1758 21734 1762 21756
rect 1782 21734 1786 21756
rect 1806 21734 1810 21756
rect 1830 21734 1834 21756
rect 1854 21734 1858 21756
rect 1878 21734 1882 21756
rect 1902 21734 1906 21756
rect 1926 21734 1930 21756
rect 1950 21734 1954 21756
rect 1974 21734 1978 21756
rect 1998 21734 2002 21756
rect 2022 21734 2026 21756
rect 2046 21734 2050 21756
rect 2070 21734 2074 21756
rect 2094 21734 2098 21756
rect 2118 21734 2122 21756
rect 2142 21734 2146 21756
rect 2166 21734 2170 21756
rect 2190 21734 2194 21756
rect 2214 21734 2218 21756
rect 2238 21734 2242 21756
rect 2262 21734 2266 21756
rect 2286 21734 2290 21756
rect 2310 21734 2314 21756
rect 2334 21734 2338 21756
rect 2358 21734 2362 21756
rect 2382 21734 2386 21756
rect 2395 21749 2400 21756
rect 2405 21735 2410 21749
rect 2406 21734 2410 21735
rect 2454 21734 2458 21780
rect 2502 21734 2506 21780
rect 2526 21734 2530 21780
rect 2550 21734 2554 21780
rect 2574 21734 2578 21780
rect 2598 21734 2602 21780
rect 2622 21734 2626 21780
rect 2646 21734 2650 21780
rect 2670 21734 2674 21780
rect 2683 21758 2717 21759
rect 2718 21758 2722 21780
rect 2742 21758 2746 21780
rect 2766 21758 2770 21780
rect 2790 21758 2794 21780
rect 2814 21758 2818 21780
rect 2838 21759 2842 21780
rect 2827 21758 2861 21759
rect 2683 21756 2861 21758
rect 2683 21749 2688 21756
rect 2693 21735 2698 21749
rect 2694 21734 2698 21735
rect 2718 21734 2722 21756
rect 2742 21734 2746 21756
rect 2766 21734 2770 21756
rect 2790 21734 2794 21756
rect 2814 21734 2818 21756
rect 2827 21749 2832 21756
rect 2838 21749 2842 21756
rect 2837 21735 2842 21749
rect 2862 21734 2866 21780
rect 2886 21734 2890 21780
rect 2910 21734 2914 21780
rect 2934 21734 2938 21780
rect 3006 21734 3010 21780
rect 3030 21734 3034 21780
rect 3054 21759 3058 21780
rect 3043 21758 3077 21759
rect 3078 21758 3082 21780
rect 3102 21758 3106 21780
rect 3115 21758 3149 21759
rect 3043 21756 3149 21758
rect 3043 21749 3048 21756
rect 3054 21749 3058 21756
rect 3053 21735 3058 21749
rect 3078 21734 3082 21756
rect 3102 21734 3106 21756
rect 3115 21749 3120 21756
rect 3125 21735 3130 21749
rect 3126 21734 3130 21735
rect 3174 21734 3178 21780
rect 3198 21734 3202 21780
rect 3222 21734 3226 21780
rect 3246 21759 3250 21780
rect 3235 21758 3269 21759
rect 3270 21758 3274 21780
rect 3283 21773 3288 21780
rect 3301 21779 3315 21780
rect 3829 21779 3843 21780
rect 3293 21759 3298 21773
rect 3307 21769 3315 21773
rect 3835 21769 3843 21773
rect 3301 21759 3307 21769
rect 3829 21759 3835 21769
rect 3283 21758 3317 21759
rect 3235 21756 3317 21758
rect 3235 21749 3240 21756
rect 3246 21749 3250 21756
rect 3245 21735 3250 21749
rect 3270 21734 3274 21756
rect 3283 21749 3288 21756
rect 3301 21755 3315 21756
rect 3293 21735 3298 21749
rect 3307 21745 3315 21749
rect 3301 21735 3307 21745
rect 3283 21734 3317 21735
rect 403 21732 3317 21734
rect 3331 21732 3365 21735
rect 3379 21732 3413 21735
rect 3811 21734 3845 21735
rect 3846 21734 3853 21780
rect 3859 21773 3864 21780
rect 3877 21779 3891 21780
rect 4549 21779 4563 21780
rect 3869 21759 3874 21773
rect 3883 21769 3891 21773
rect 4555 21769 4563 21773
rect 3877 21759 3883 21769
rect 4549 21759 4555 21769
rect 3859 21734 3893 21735
rect 3811 21732 3893 21734
rect 4531 21734 4565 21735
rect 4566 21734 4573 21780
rect 4579 21773 4584 21780
rect 4597 21779 4611 21780
rect 4789 21779 4803 21780
rect 4589 21759 4594 21773
rect 4603 21769 4611 21773
rect 4795 21769 4803 21773
rect 4597 21759 4603 21769
rect 4789 21759 4795 21769
rect 4579 21734 4613 21735
rect 4531 21732 4613 21734
rect 4771 21734 4805 21735
rect 4806 21734 4813 21780
rect 4819 21773 4824 21780
rect 4837 21779 4851 21780
rect 6565 21779 6579 21780
rect 4829 21759 4834 21773
rect 4843 21769 4851 21773
rect 4837 21759 4843 21769
rect 6606 21756 6610 21780
rect 6619 21773 6624 21780
rect 6629 21759 6634 21773
rect 6654 21770 6658 21794
rect 6667 21782 6701 21783
rect 6702 21782 6706 21803
rect 6715 21797 6720 21804
rect 6750 21803 6754 21804
rect 6725 21783 6730 21797
rect 6739 21793 6747 21797
rect 6733 21783 6739 21793
rect 6726 21782 6730 21783
rect 6667 21780 6747 21782
rect 6664 21766 6672 21770
rect 4819 21734 4853 21735
rect 4771 21732 4853 21734
rect 6571 21734 6605 21735
rect 6606 21734 6613 21755
rect 6620 21746 6624 21756
rect 6643 21749 6648 21759
rect 6702 21756 6706 21780
rect 6678 21755 6682 21756
rect 6653 21746 6658 21749
rect 6630 21734 6634 21746
rect 6667 21745 6675 21749
rect 6653 21735 6658 21736
rect 6661 21735 6667 21745
rect 6678 21734 6685 21755
rect 6702 21734 6709 21755
rect 6726 21734 6730 21780
rect 6733 21779 6747 21780
rect 6750 21758 6757 21803
rect 6774 21758 6778 21804
rect 6798 21758 6802 21804
rect 6805 21803 6819 21804
rect 6822 21782 6829 21828
rect 6846 21782 6850 21828
rect 6870 21782 6874 21828
rect 6894 21782 6898 21828
rect 6918 21782 6922 21828
rect 6942 21782 6946 21828
rect 6949 21827 6963 21828
rect 6966 21827 6973 21828
rect 6997 21827 7011 21828
rect 7014 21827 7021 21828
rect 7014 21804 7018 21827
rect 6966 21803 6970 21804
rect 6805 21780 6963 21782
rect 6805 21779 6819 21780
rect 6733 21756 6819 21758
rect 6733 21755 6747 21756
rect 6571 21732 6675 21734
rect 403 21725 408 21732
rect 413 21711 418 21725
rect 414 21686 418 21711
rect 462 21686 466 21732
rect 486 21686 490 21732
rect 510 21686 514 21732
rect 534 21686 538 21732
rect 558 21686 562 21732
rect 582 21686 586 21732
rect 606 21686 610 21732
rect 630 21686 634 21732
rect 654 21686 658 21732
rect 678 21686 682 21732
rect 702 21686 706 21732
rect 726 21686 730 21732
rect 750 21686 754 21732
rect 774 21686 778 21732
rect 798 21686 802 21732
rect 822 21686 826 21732
rect 846 21686 850 21732
rect 870 21686 874 21732
rect 894 21686 898 21732
rect 918 21686 922 21732
rect 942 21686 946 21732
rect 966 21686 970 21732
rect 990 21686 994 21732
rect 1014 21686 1018 21732
rect 1038 21686 1042 21732
rect 1062 21686 1066 21732
rect 1086 21686 1090 21732
rect 1110 21686 1114 21732
rect 1134 21686 1138 21732
rect 1158 21686 1162 21732
rect 1182 21686 1186 21732
rect 1206 21686 1210 21732
rect 1219 21710 1253 21711
rect 1278 21710 1282 21732
rect 1302 21710 1306 21732
rect 1326 21710 1330 21732
rect 1350 21710 1354 21732
rect 1374 21710 1378 21732
rect 1446 21710 1450 21732
rect 1470 21710 1474 21732
rect 1494 21710 1498 21732
rect 1518 21710 1522 21732
rect 1542 21710 1546 21732
rect 1566 21710 1570 21732
rect 1590 21710 1594 21732
rect 1614 21710 1618 21732
rect 1638 21710 1642 21732
rect 1662 21710 1666 21732
rect 1686 21710 1690 21732
rect 1710 21710 1714 21732
rect 1734 21710 1738 21732
rect 1758 21710 1762 21732
rect 1782 21710 1786 21732
rect 1806 21710 1810 21732
rect 1830 21710 1834 21732
rect 1854 21710 1858 21732
rect 1878 21710 1882 21732
rect 1902 21710 1906 21732
rect 1926 21710 1930 21732
rect 1950 21710 1954 21732
rect 1974 21710 1978 21732
rect 1998 21710 2002 21732
rect 2022 21710 2026 21732
rect 2046 21710 2050 21732
rect 2070 21710 2074 21732
rect 2094 21710 2098 21732
rect 2118 21710 2122 21732
rect 2142 21710 2146 21732
rect 2166 21710 2170 21732
rect 2190 21710 2194 21732
rect 2214 21710 2218 21732
rect 2238 21710 2242 21732
rect 2262 21710 2266 21732
rect 2286 21710 2290 21732
rect 2310 21710 2314 21732
rect 2334 21710 2338 21732
rect 2358 21710 2362 21732
rect 2382 21710 2386 21732
rect 2406 21710 2410 21732
rect 2454 21710 2458 21732
rect 1219 21708 2475 21710
rect 1219 21701 1224 21708
rect 1229 21687 1234 21701
rect 1230 21686 1234 21687
rect 1278 21686 1282 21708
rect 1302 21686 1306 21708
rect 1326 21686 1330 21708
rect 1350 21686 1354 21708
rect 1374 21686 1378 21708
rect 1446 21686 1450 21708
rect 1470 21686 1474 21708
rect 1494 21686 1498 21708
rect 1518 21686 1522 21708
rect 1542 21686 1546 21708
rect 1566 21686 1570 21708
rect 1590 21686 1594 21708
rect 1614 21686 1618 21708
rect 1638 21686 1642 21708
rect 1662 21686 1666 21708
rect 1686 21686 1690 21708
rect 1710 21686 1714 21708
rect 1734 21686 1738 21708
rect 1758 21686 1762 21708
rect 1782 21686 1786 21708
rect 1806 21686 1810 21708
rect 1830 21686 1834 21708
rect 1854 21686 1858 21708
rect 1878 21686 1882 21708
rect 1902 21686 1906 21708
rect 1926 21686 1930 21708
rect 1950 21686 1954 21708
rect 1974 21686 1978 21708
rect 1998 21686 2002 21708
rect 2022 21686 2026 21708
rect 2046 21686 2050 21708
rect 2070 21686 2074 21708
rect 2094 21686 2098 21708
rect 2118 21686 2122 21708
rect 2142 21686 2146 21708
rect 2166 21686 2170 21708
rect 2190 21686 2194 21708
rect 2214 21686 2218 21708
rect 2238 21686 2242 21708
rect 2262 21686 2266 21708
rect 2286 21686 2290 21708
rect 2310 21686 2314 21708
rect 2334 21686 2338 21708
rect 2358 21686 2362 21708
rect 2382 21686 2386 21708
rect 2406 21686 2410 21708
rect 2454 21686 2458 21708
rect 2461 21707 2475 21708
rect 2478 21707 2485 21731
rect 2478 21686 2482 21707
rect 2502 21686 2506 21732
rect 2526 21686 2530 21732
rect 2550 21686 2554 21732
rect 2574 21686 2578 21732
rect 2598 21686 2602 21732
rect 2622 21686 2626 21732
rect 2646 21686 2650 21732
rect 2670 21686 2674 21732
rect 2694 21686 2698 21732
rect 2718 21731 2722 21732
rect 2718 21710 2725 21731
rect 2742 21710 2746 21732
rect 2766 21710 2770 21732
rect 2790 21710 2794 21732
rect 2814 21710 2818 21732
rect 2862 21710 2866 21732
rect 2886 21710 2890 21732
rect 2910 21710 2914 21732
rect 2934 21710 2938 21732
rect 2958 21710 2965 21731
rect 2982 21710 2989 21731
rect 3006 21710 3010 21732
rect 3030 21710 3034 21732
rect 3078 21710 3082 21732
rect 3102 21710 3106 21732
rect 3126 21710 3130 21732
rect 3174 21710 3178 21732
rect 3198 21710 3202 21732
rect 3222 21710 3226 21732
rect 3270 21710 3274 21732
rect 3283 21725 3288 21732
rect 3301 21731 3315 21732
rect 3829 21731 3843 21732
rect 3293 21711 3298 21725
rect 3307 21721 3315 21725
rect 3835 21721 3843 21725
rect 3301 21711 3307 21721
rect 3829 21711 3835 21721
rect 3283 21710 3317 21711
rect 2701 21708 2955 21710
rect 2701 21707 2715 21708
rect 2718 21707 2725 21708
rect 2742 21686 2746 21708
rect 2766 21686 2770 21708
rect 2790 21686 2794 21708
rect 2814 21686 2818 21708
rect 2862 21686 2866 21708
rect 2886 21686 2890 21708
rect 2910 21686 2914 21708
rect 2934 21686 2938 21708
rect 2941 21707 2955 21708
rect 2958 21708 3317 21710
rect 3331 21708 3365 21711
rect 3379 21708 3413 21711
rect 3811 21710 3845 21711
rect 3846 21710 3853 21732
rect 3859 21725 3864 21732
rect 3877 21731 3891 21732
rect 4549 21731 4563 21732
rect 3869 21711 3874 21725
rect 3883 21721 3891 21725
rect 4555 21721 4563 21725
rect 3877 21711 3883 21721
rect 4549 21711 4555 21721
rect 3859 21710 3893 21711
rect 3811 21708 3893 21710
rect 4531 21710 4565 21711
rect 4566 21710 4573 21732
rect 4579 21725 4584 21732
rect 4597 21731 4611 21732
rect 4789 21731 4803 21732
rect 4589 21711 4594 21725
rect 4603 21721 4611 21725
rect 4795 21721 4803 21725
rect 4597 21711 4603 21721
rect 4789 21711 4795 21721
rect 4579 21710 4613 21711
rect 4531 21708 4613 21710
rect 4771 21710 4805 21711
rect 4806 21710 4813 21732
rect 4819 21725 4824 21732
rect 4837 21731 4851 21732
rect 6589 21731 6603 21732
rect 4829 21711 4834 21725
rect 4843 21721 4851 21725
rect 6595 21721 6603 21725
rect 4837 21711 4843 21721
rect 6589 21711 6595 21721
rect 4819 21710 4853 21711
rect 4771 21708 4853 21710
rect 6571 21710 6605 21711
rect 6606 21710 6613 21732
rect 6630 21710 6634 21732
rect 6661 21731 6675 21732
rect 6678 21732 6747 21734
rect 6678 21731 6699 21732
rect 6702 21731 6709 21732
rect 6571 21708 6651 21710
rect 6702 21708 6706 21731
rect 2958 21707 2979 21708
rect 2982 21707 2989 21708
rect 2958 21686 2962 21707
rect 2982 21686 2986 21707
rect 3006 21686 3010 21708
rect 3030 21686 3034 21708
rect 3078 21686 3082 21708
rect 3102 21686 3106 21708
rect 3126 21686 3130 21708
rect 3174 21686 3178 21708
rect 3198 21686 3202 21708
rect 3222 21686 3226 21708
rect 3270 21686 3274 21708
rect 3283 21701 3288 21708
rect 3301 21707 3315 21708
rect 3829 21707 3843 21708
rect 3293 21687 3298 21701
rect 3307 21697 3315 21701
rect 3835 21697 3843 21701
rect 3301 21687 3307 21697
rect 3829 21687 3835 21697
rect 3283 21686 3317 21687
rect -389 21684 3317 21686
rect 3331 21684 3365 21687
rect 3379 21684 3413 21687
rect 3811 21686 3845 21687
rect 3846 21686 3853 21708
rect 3859 21701 3864 21708
rect 3877 21707 3891 21708
rect 4549 21707 4563 21708
rect 3869 21687 3874 21701
rect 3883 21697 3891 21701
rect 4555 21697 4563 21701
rect 3877 21687 3883 21697
rect 4549 21687 4555 21697
rect 3859 21686 3893 21687
rect 3811 21684 3893 21686
rect 4531 21686 4565 21687
rect 4566 21686 4573 21708
rect 4579 21701 4584 21708
rect 4597 21707 4611 21708
rect 4789 21707 4803 21708
rect 4589 21687 4594 21701
rect 4603 21697 4611 21701
rect 4795 21697 4803 21701
rect 4597 21687 4603 21697
rect 4789 21687 4795 21697
rect 4579 21686 4613 21687
rect 4531 21684 4613 21686
rect 4771 21686 4805 21687
rect 4806 21686 4813 21708
rect 4819 21701 4824 21708
rect 4837 21707 4851 21708
rect 6589 21707 6603 21708
rect 4829 21687 4834 21701
rect 4843 21697 4851 21701
rect 6595 21697 6603 21701
rect 4837 21687 4843 21697
rect 6589 21687 6595 21697
rect 4819 21686 4853 21687
rect 4771 21684 4853 21686
rect 6571 21686 6605 21687
rect 6606 21686 6613 21708
rect 6630 21686 6634 21708
rect 6637 21707 6651 21708
rect 6571 21684 6651 21686
rect 6678 21684 6682 21708
rect 6702 21686 6709 21707
rect 6726 21686 6730 21732
rect 6733 21731 6747 21732
rect 6750 21710 6757 21756
rect 6774 21710 6778 21756
rect 6798 21710 6802 21756
rect 6805 21755 6819 21756
rect 6822 21734 6829 21780
rect 6846 21734 6850 21780
rect 6870 21734 6874 21780
rect 6894 21734 6898 21780
rect 6918 21734 6922 21780
rect 6942 21734 6946 21780
rect 6949 21779 6963 21780
rect 6966 21758 6973 21803
rect 7014 21782 7021 21803
rect 7038 21782 7042 21828
rect 7045 21827 7059 21828
rect 7109 21807 7114 21821
rect 7099 21797 7104 21807
rect 7118 21804 7133 21807
rect 7507 21804 7541 21807
rect 7555 21804 7589 21807
rect 8251 21804 8285 21807
rect 8299 21804 8318 21807
rect 7109 21783 7114 21797
rect 7123 21793 7131 21797
rect 7579 21793 7587 21797
rect 7117 21783 7123 21793
rect 7573 21783 7579 21793
rect 8309 21783 8314 21797
rect 7099 21782 7133 21783
rect 6997 21780 7133 21782
rect 7507 21780 7541 21783
rect 7555 21780 7589 21783
rect 14515 21780 14549 21783
rect 14563 21780 14582 21783
rect 6997 21779 7011 21780
rect 7014 21779 7021 21780
rect 7038 21758 7042 21780
rect 7099 21773 7104 21780
rect 7117 21779 7131 21780
rect 7573 21779 7587 21780
rect 7621 21779 7635 21780
rect 7109 21759 7114 21773
rect 7123 21769 7131 21773
rect 7117 21759 7123 21769
rect 8286 21760 8293 21779
rect 14573 21759 14578 21773
rect 7099 21758 7133 21759
rect 6949 21756 7133 21758
rect 7507 21756 7541 21759
rect 7555 21756 7574 21759
rect 8227 21756 8261 21759
rect 8275 21758 8309 21759
rect 8269 21756 8309 21758
rect 14515 21756 14549 21759
rect 6949 21755 6963 21756
rect 6966 21755 6973 21756
rect 6966 21734 6970 21755
rect 7038 21734 7042 21756
rect 7099 21749 7104 21756
rect 7117 21755 7131 21756
rect 8269 21755 8283 21756
rect 8317 21755 8331 21756
rect 7109 21735 7114 21749
rect 7123 21745 7131 21749
rect 7117 21735 7123 21745
rect 7565 21735 7570 21749
rect 8285 21735 8293 21749
rect 14539 21745 14547 21749
rect 14533 21735 14539 21745
rect 7099 21734 7133 21735
rect 6805 21732 7133 21734
rect 7507 21732 7541 21735
rect 6805 21731 6819 21732
rect 6822 21731 6829 21732
rect 6822 21710 6826 21731
rect 6846 21710 6850 21732
rect 6870 21710 6874 21732
rect 6894 21710 6898 21732
rect 6918 21710 6922 21732
rect 6942 21710 6946 21732
rect 6966 21710 6970 21732
rect 7038 21710 7042 21732
rect 7099 21725 7104 21732
rect 7117 21731 7131 21732
rect 7109 21711 7114 21725
rect 7123 21721 7131 21725
rect 7531 21721 7539 21725
rect 7117 21711 7123 21721
rect 7525 21711 7531 21721
rect 7099 21710 7133 21711
rect 6733 21708 7133 21710
rect 7507 21710 7541 21711
rect 7542 21710 7549 21731
rect 7555 21725 7560 21735
rect 7574 21732 7589 21735
rect 8227 21732 8261 21735
rect 8275 21734 8309 21735
rect 8269 21732 8309 21734
rect 14515 21734 14549 21735
rect 14550 21734 14557 21755
rect 14563 21749 14568 21759
rect 14582 21756 14597 21759
rect 14573 21735 14578 21749
rect 14587 21745 14595 21749
rect 14581 21735 14587 21745
rect 14563 21734 14597 21735
rect 14515 21732 14597 21734
rect 14731 21732 14765 21735
rect 14779 21732 14798 21735
rect 14971 21732 15005 21735
rect 15019 21732 15038 21735
rect 8269 21731 8283 21732
rect 8317 21731 8331 21732
rect 14533 21731 14547 21732
rect 7565 21711 7570 21725
rect 7579 21721 7587 21725
rect 7573 21711 7579 21721
rect 8285 21711 8293 21725
rect 14539 21721 14547 21725
rect 14533 21711 14539 21721
rect 7555 21710 7589 21711
rect 7507 21708 7589 21710
rect 8227 21708 8261 21711
rect 8275 21710 8309 21711
rect 8269 21708 8309 21710
rect 14515 21710 14549 21711
rect 14550 21710 14557 21732
rect 14563 21725 14568 21732
rect 14581 21731 14595 21732
rect 14573 21711 14578 21725
rect 14587 21721 14595 21725
rect 14581 21711 14587 21721
rect 14789 21711 14797 21725
rect 15029 21711 15034 21725
rect 14563 21710 14597 21711
rect 14515 21708 14597 21710
rect 14731 21708 14765 21711
rect 14779 21710 14813 21711
rect 14773 21708 14813 21710
rect 14971 21708 15005 21711
rect 6733 21707 6747 21708
rect 6750 21707 6757 21708
rect 6750 21686 6754 21707
rect 6774 21686 6778 21708
rect 6798 21686 6802 21708
rect 6822 21686 6826 21708
rect 6846 21686 6850 21708
rect 6870 21686 6874 21708
rect 6894 21686 6898 21708
rect 6918 21686 6922 21708
rect 6942 21686 6946 21708
rect 6966 21686 6970 21708
rect 7038 21686 7042 21708
rect 7099 21701 7104 21708
rect 7117 21707 7131 21708
rect 7525 21707 7539 21708
rect 7109 21687 7114 21701
rect 7123 21697 7131 21701
rect 7531 21697 7539 21701
rect 7117 21687 7123 21697
rect 7525 21687 7531 21697
rect 7099 21686 7133 21687
rect 6685 21684 7133 21686
rect -389 21677 -384 21684
rect -379 21663 -374 21677
rect -378 21662 -374 21663
rect -354 21662 -350 21684
rect -330 21662 -326 21684
rect -306 21662 -302 21684
rect -282 21662 -278 21684
rect -258 21662 -254 21684
rect -234 21662 -230 21684
rect -210 21662 -206 21684
rect -186 21662 -182 21684
rect -162 21662 -158 21684
rect -138 21662 -134 21684
rect -114 21662 -110 21684
rect -90 21662 -86 21684
rect -66 21662 -62 21684
rect -42 21662 -38 21684
rect -18 21662 -14 21684
rect 6 21662 10 21684
rect 30 21662 34 21684
rect 54 21662 58 21684
rect 78 21662 82 21684
rect 102 21662 106 21684
rect 126 21662 130 21684
rect 150 21662 154 21684
rect 174 21662 178 21684
rect 198 21662 202 21684
rect 222 21662 226 21684
rect 246 21662 250 21684
rect 270 21662 274 21684
rect 294 21662 298 21684
rect 318 21662 322 21684
rect 342 21662 346 21684
rect 366 21662 370 21684
rect 390 21662 394 21684
rect 414 21662 418 21684
rect 462 21662 466 21684
rect 486 21662 490 21684
rect 510 21662 514 21684
rect 534 21662 538 21684
rect 558 21662 562 21684
rect 582 21662 586 21684
rect 606 21662 610 21684
rect 630 21662 634 21684
rect 654 21662 658 21684
rect 678 21662 682 21684
rect 702 21662 706 21684
rect 726 21662 730 21684
rect 750 21662 754 21684
rect 774 21662 778 21684
rect 798 21662 802 21684
rect 822 21662 826 21684
rect 846 21662 850 21684
rect 870 21662 874 21684
rect 894 21662 898 21684
rect 918 21662 922 21684
rect 942 21662 946 21684
rect 966 21662 970 21684
rect 990 21662 994 21684
rect 1014 21662 1018 21684
rect 1038 21662 1042 21684
rect 1062 21662 1066 21684
rect 1086 21662 1090 21684
rect 1110 21662 1114 21684
rect 1134 21662 1138 21684
rect 1158 21662 1162 21684
rect 1182 21662 1186 21684
rect 1206 21662 1210 21684
rect 1230 21662 1234 21684
rect 1278 21662 1282 21684
rect 1302 21662 1306 21684
rect 1326 21662 1330 21684
rect 1350 21662 1354 21684
rect 1374 21662 1378 21684
rect 1446 21662 1450 21684
rect 1470 21662 1474 21684
rect 1494 21662 1498 21684
rect 1518 21662 1522 21684
rect 1542 21662 1546 21684
rect 1566 21662 1570 21684
rect 1590 21662 1594 21684
rect 1614 21662 1618 21684
rect 1638 21662 1642 21684
rect 1662 21662 1666 21684
rect 1686 21662 1690 21684
rect 1710 21662 1714 21684
rect 1734 21662 1738 21684
rect 1758 21662 1762 21684
rect 1782 21662 1786 21684
rect 1806 21662 1810 21684
rect 1830 21662 1834 21684
rect 1854 21662 1858 21684
rect 1878 21662 1882 21684
rect 1902 21662 1906 21684
rect 1926 21662 1930 21684
rect 1950 21662 1954 21684
rect 1974 21662 1978 21684
rect 1998 21662 2002 21684
rect 2022 21662 2026 21684
rect 2046 21662 2050 21684
rect 2070 21662 2074 21684
rect 2094 21662 2098 21684
rect 2118 21662 2122 21684
rect 2142 21662 2146 21684
rect 2166 21662 2170 21684
rect 2190 21662 2194 21684
rect 2214 21662 2218 21684
rect 2238 21662 2242 21684
rect 2262 21662 2266 21684
rect 2286 21662 2290 21684
rect 2310 21662 2314 21684
rect 2334 21662 2338 21684
rect 2358 21662 2362 21684
rect 2382 21662 2386 21684
rect 2406 21662 2410 21684
rect -1109 21660 2427 21662
rect -1109 21653 -1104 21660
rect -1099 21639 -1094 21653
rect -1098 21614 -1094 21639
rect -1074 21614 -1070 21660
rect -1050 21614 -1046 21660
rect -1026 21614 -1022 21660
rect -1002 21614 -998 21660
rect -978 21614 -974 21660
rect -954 21614 -950 21660
rect -930 21614 -926 21660
rect -906 21614 -902 21660
rect -882 21614 -878 21660
rect -858 21614 -854 21660
rect -834 21614 -830 21660
rect -810 21614 -806 21660
rect -786 21614 -782 21660
rect -762 21614 -758 21660
rect -738 21614 -734 21660
rect -714 21614 -710 21660
rect -690 21614 -686 21660
rect -666 21614 -662 21660
rect -642 21614 -638 21660
rect -618 21614 -614 21660
rect -594 21614 -590 21660
rect -570 21614 -566 21660
rect -546 21614 -542 21660
rect -522 21614 -518 21660
rect -498 21614 -494 21660
rect -474 21614 -470 21660
rect -450 21614 -446 21660
rect -426 21614 -422 21660
rect -402 21614 -398 21660
rect -378 21614 -374 21660
rect -354 21635 -350 21660
rect -2393 21612 -357 21614
rect -2371 21590 -2366 21612
rect -2348 21590 -2343 21612
rect -2325 21604 -2317 21612
rect -2109 21607 -2087 21612
rect -2117 21605 -2085 21607
rect -2325 21590 -2320 21604
rect -2317 21602 -2309 21604
rect -2309 21590 -2301 21602
rect -2023 21595 -2021 21604
rect -2037 21594 -2021 21595
rect -2051 21592 -2021 21594
rect -2074 21590 -2021 21592
rect -2000 21590 -1992 21612
rect -1969 21605 -1921 21607
rect -1671 21604 -1663 21612
rect -1663 21602 -1655 21604
rect -1655 21590 -1647 21602
rect -1642 21590 -1637 21612
rect -1619 21590 -1614 21612
rect -1530 21590 -1526 21612
rect -1506 21590 -1502 21612
rect -1482 21590 -1478 21612
rect -1458 21590 -1454 21612
rect -1434 21590 -1430 21612
rect -1410 21590 -1406 21612
rect -1386 21590 -1382 21612
rect -1362 21590 -1358 21612
rect -1338 21590 -1334 21612
rect -1314 21590 -1310 21612
rect -1290 21590 -1286 21612
rect -1266 21590 -1262 21612
rect -1242 21590 -1238 21612
rect -1218 21590 -1214 21612
rect -1194 21590 -1190 21612
rect -1170 21590 -1166 21612
rect -1146 21590 -1142 21612
rect -1122 21590 -1118 21612
rect -1098 21590 -1094 21612
rect -1074 21611 -1070 21612
rect -2393 21588 -1077 21590
rect -2371 21542 -2366 21588
rect -2348 21542 -2343 21588
rect -2325 21576 -2317 21588
rect -2117 21581 -2087 21585
rect -2325 21556 -2320 21576
rect -2317 21574 -2309 21576
rect -2325 21548 -2317 21556
rect -2101 21551 -2071 21554
rect -2325 21542 -2320 21548
rect -2317 21542 -2309 21548
rect -2000 21546 -1992 21588
rect -1969 21581 -1921 21585
rect -1864 21581 -1680 21586
rect -1671 21576 -1663 21588
rect -1663 21574 -1655 21576
rect -1854 21560 -1680 21564
rect -1846 21551 -1798 21554
rect -2079 21545 -2043 21546
rect -2007 21545 -1991 21546
rect -2079 21544 -2071 21545
rect -2079 21542 -2029 21544
rect -2011 21542 -1991 21545
rect -1846 21543 -1806 21549
rect -1671 21548 -1663 21556
rect -1864 21542 -1796 21543
rect -1663 21542 -1655 21548
rect -1642 21542 -1637 21588
rect -1619 21542 -1614 21588
rect -1530 21542 -1526 21588
rect -1506 21542 -1502 21588
rect -1482 21542 -1478 21588
rect -1458 21542 -1454 21588
rect -1434 21542 -1430 21588
rect -1410 21542 -1406 21588
rect -1386 21542 -1382 21588
rect -1362 21542 -1358 21588
rect -1338 21542 -1334 21588
rect -1314 21542 -1310 21588
rect -1290 21542 -1286 21588
rect -1266 21542 -1262 21588
rect -1242 21542 -1238 21588
rect -1218 21542 -1214 21588
rect -1194 21542 -1190 21588
rect -1170 21542 -1166 21588
rect -1146 21542 -1142 21588
rect -1122 21542 -1118 21588
rect -1098 21542 -1094 21588
rect -1091 21587 -1077 21588
rect -1074 21566 -1067 21611
rect -1050 21566 -1046 21612
rect -1026 21566 -1022 21612
rect -1002 21566 -998 21612
rect -978 21566 -974 21612
rect -954 21566 -950 21612
rect -930 21566 -926 21612
rect -906 21566 -902 21612
rect -882 21566 -878 21612
rect -858 21566 -854 21612
rect -834 21566 -830 21612
rect -810 21566 -806 21612
rect -786 21566 -782 21612
rect -762 21566 -758 21612
rect -738 21566 -734 21612
rect -714 21566 -710 21612
rect -690 21566 -686 21612
rect -666 21566 -662 21612
rect -642 21566 -638 21612
rect -618 21566 -614 21612
rect -594 21566 -590 21612
rect -570 21566 -566 21612
rect -546 21566 -542 21612
rect -522 21566 -518 21612
rect -498 21566 -494 21612
rect -474 21566 -470 21612
rect -450 21566 -446 21612
rect -426 21566 -422 21612
rect -402 21566 -398 21612
rect -378 21566 -374 21612
rect -371 21611 -357 21612
rect -354 21590 -347 21635
rect -330 21590 -326 21660
rect -306 21590 -302 21660
rect -282 21590 -278 21660
rect -258 21590 -254 21660
rect -234 21590 -230 21660
rect -210 21590 -206 21660
rect -186 21590 -182 21660
rect -162 21590 -158 21660
rect -138 21590 -134 21660
rect -114 21590 -110 21660
rect -90 21590 -86 21660
rect -66 21590 -62 21660
rect -42 21590 -38 21660
rect -18 21590 -14 21660
rect 6 21590 10 21660
rect 30 21590 34 21660
rect 54 21590 58 21660
rect 78 21590 82 21660
rect 102 21590 106 21660
rect 126 21590 130 21660
rect 150 21590 154 21660
rect 174 21590 178 21660
rect 198 21590 202 21660
rect 222 21590 226 21660
rect 246 21590 250 21660
rect 270 21590 274 21660
rect 294 21590 298 21660
rect 318 21590 322 21660
rect 342 21590 346 21660
rect 366 21590 370 21660
rect 390 21590 394 21660
rect 414 21590 418 21660
rect 438 21638 445 21659
rect 462 21638 466 21660
rect 486 21638 490 21660
rect 510 21638 514 21660
rect 534 21638 538 21660
rect 558 21638 562 21660
rect 582 21638 586 21660
rect 606 21638 610 21660
rect 630 21638 634 21660
rect 654 21638 658 21660
rect 678 21638 682 21660
rect 702 21638 706 21660
rect 726 21638 730 21660
rect 750 21638 754 21660
rect 774 21638 778 21660
rect 798 21638 802 21660
rect 822 21638 826 21660
rect 846 21638 850 21660
rect 870 21638 874 21660
rect 894 21638 898 21660
rect 918 21638 922 21660
rect 942 21638 946 21660
rect 966 21638 970 21660
rect 990 21638 994 21660
rect 1014 21638 1018 21660
rect 1038 21638 1042 21660
rect 1062 21638 1066 21660
rect 1086 21638 1090 21660
rect 1110 21638 1114 21660
rect 1134 21638 1138 21660
rect 1158 21638 1162 21660
rect 1182 21638 1186 21660
rect 1206 21638 1210 21660
rect 1230 21638 1234 21660
rect 1278 21638 1282 21660
rect 1302 21638 1306 21660
rect 1326 21638 1330 21660
rect 1350 21638 1354 21660
rect 1374 21638 1378 21660
rect 1387 21638 1421 21639
rect 421 21636 1421 21638
rect 421 21635 435 21636
rect 438 21635 445 21636
rect 438 21590 442 21635
rect 462 21590 466 21636
rect 486 21590 490 21636
rect 510 21590 514 21636
rect 534 21590 538 21636
rect 558 21590 562 21636
rect 582 21590 586 21636
rect 606 21590 610 21636
rect 630 21590 634 21636
rect 654 21590 658 21636
rect 678 21590 682 21636
rect 702 21590 706 21636
rect 726 21590 730 21636
rect 750 21590 754 21636
rect 774 21590 778 21636
rect 798 21590 802 21636
rect 822 21590 826 21636
rect 846 21590 850 21636
rect 870 21590 874 21636
rect 894 21590 898 21636
rect 918 21590 922 21636
rect 942 21590 946 21636
rect 966 21590 970 21636
rect 990 21590 994 21636
rect 1014 21590 1018 21636
rect 1038 21590 1042 21636
rect 1062 21590 1066 21636
rect 1086 21590 1090 21636
rect 1110 21590 1114 21636
rect 1134 21590 1138 21636
rect 1158 21590 1162 21636
rect 1182 21590 1186 21636
rect 1206 21590 1210 21636
rect 1230 21590 1234 21636
rect 1254 21614 1261 21635
rect 1278 21614 1282 21636
rect 1302 21614 1306 21636
rect 1326 21614 1330 21636
rect 1350 21614 1354 21636
rect 1374 21614 1378 21636
rect 1387 21629 1392 21636
rect 1397 21615 1402 21629
rect 1398 21614 1402 21615
rect 1446 21614 1450 21660
rect 1470 21614 1474 21660
rect 1494 21614 1498 21660
rect 1518 21614 1522 21660
rect 1542 21614 1546 21660
rect 1566 21614 1570 21660
rect 1590 21614 1594 21660
rect 1614 21614 1618 21660
rect 1638 21614 1642 21660
rect 1662 21614 1666 21660
rect 1686 21614 1690 21660
rect 1710 21614 1714 21660
rect 1734 21614 1738 21660
rect 1758 21614 1762 21660
rect 1782 21614 1786 21660
rect 1806 21614 1810 21660
rect 1830 21614 1834 21660
rect 1854 21614 1858 21660
rect 1878 21614 1882 21660
rect 1902 21614 1906 21660
rect 1926 21614 1930 21660
rect 1950 21614 1954 21660
rect 1974 21614 1978 21660
rect 1998 21614 2002 21660
rect 2022 21614 2026 21660
rect 2046 21614 2050 21660
rect 2070 21614 2074 21660
rect 2094 21614 2098 21660
rect 2118 21614 2122 21660
rect 2142 21614 2146 21660
rect 2166 21614 2170 21660
rect 2190 21614 2194 21660
rect 2214 21614 2218 21660
rect 2238 21614 2242 21660
rect 2262 21614 2266 21660
rect 2286 21614 2290 21660
rect 2310 21614 2314 21660
rect 2334 21614 2338 21660
rect 2358 21614 2362 21660
rect 2382 21615 2386 21660
rect 2371 21614 2405 21615
rect 1237 21612 2405 21614
rect 1237 21611 1251 21612
rect 1254 21611 1261 21612
rect 1254 21590 1258 21611
rect 1278 21590 1282 21612
rect 1302 21590 1306 21612
rect 1326 21590 1330 21612
rect 1350 21590 1354 21612
rect 1374 21590 1378 21612
rect 1398 21590 1402 21612
rect 1446 21590 1450 21612
rect 1470 21590 1474 21612
rect 1494 21590 1498 21612
rect 1518 21590 1522 21612
rect 1542 21590 1546 21612
rect 1566 21590 1570 21612
rect 1590 21590 1594 21612
rect 1614 21590 1618 21612
rect 1638 21590 1642 21612
rect 1662 21590 1666 21612
rect 1686 21590 1690 21612
rect 1710 21590 1714 21612
rect 1734 21590 1738 21612
rect 1758 21590 1762 21612
rect 1782 21590 1786 21612
rect 1806 21590 1810 21612
rect 1830 21590 1834 21612
rect 1854 21590 1858 21612
rect 1878 21590 1882 21612
rect 1902 21590 1906 21612
rect 1926 21590 1930 21612
rect 1950 21590 1954 21612
rect 1974 21590 1978 21612
rect 1998 21590 2002 21612
rect 2022 21590 2026 21612
rect 2046 21590 2050 21612
rect 2070 21590 2074 21612
rect 2094 21590 2098 21612
rect 2118 21590 2122 21612
rect 2142 21590 2146 21612
rect 2166 21590 2170 21612
rect 2190 21590 2194 21612
rect 2214 21590 2218 21612
rect 2238 21590 2242 21612
rect 2262 21590 2266 21612
rect 2286 21590 2290 21612
rect 2310 21590 2314 21612
rect 2334 21591 2338 21612
rect 2323 21590 2357 21591
rect -371 21588 2357 21590
rect -371 21587 -357 21588
rect -354 21587 -347 21588
rect -354 21566 -350 21587
rect -330 21566 -326 21588
rect -306 21566 -302 21588
rect -282 21566 -278 21588
rect -258 21566 -254 21588
rect -234 21566 -230 21588
rect -210 21566 -206 21588
rect -186 21566 -182 21588
rect -162 21566 -158 21588
rect -138 21566 -134 21588
rect -114 21566 -110 21588
rect -90 21566 -86 21588
rect -66 21566 -62 21588
rect -42 21566 -38 21588
rect -18 21566 -14 21588
rect 6 21566 10 21588
rect 30 21566 34 21588
rect 54 21566 58 21588
rect 78 21566 82 21588
rect 102 21566 106 21588
rect 126 21566 130 21588
rect 150 21566 154 21588
rect 174 21566 178 21588
rect 198 21566 202 21588
rect 222 21566 226 21588
rect 246 21566 250 21588
rect 270 21566 274 21588
rect 294 21566 298 21588
rect 318 21566 322 21588
rect 342 21566 346 21588
rect 366 21566 370 21588
rect 390 21566 394 21588
rect 414 21566 418 21588
rect 438 21566 442 21588
rect 462 21566 466 21588
rect 486 21566 490 21588
rect 510 21566 514 21588
rect 534 21566 538 21588
rect 558 21566 562 21588
rect 582 21566 586 21588
rect 606 21566 610 21588
rect 630 21566 634 21588
rect 654 21566 658 21588
rect 678 21566 682 21588
rect 702 21566 706 21588
rect 726 21566 730 21588
rect 750 21566 754 21588
rect 774 21566 778 21588
rect 798 21566 802 21588
rect 822 21566 826 21588
rect 846 21566 850 21588
rect 870 21566 874 21588
rect 894 21566 898 21588
rect 918 21566 922 21588
rect 942 21566 946 21588
rect 966 21566 970 21588
rect 990 21566 994 21588
rect 1014 21566 1018 21588
rect 1038 21566 1042 21588
rect 1062 21566 1066 21588
rect 1086 21566 1090 21588
rect 1110 21566 1114 21588
rect 1134 21566 1138 21588
rect 1158 21566 1162 21588
rect 1182 21566 1186 21588
rect 1206 21566 1210 21588
rect 1230 21566 1234 21588
rect 1254 21566 1258 21588
rect 1278 21566 1282 21588
rect 1302 21566 1306 21588
rect 1326 21567 1330 21588
rect 1315 21566 1349 21567
rect -1091 21564 1349 21566
rect -1091 21563 -1077 21564
rect -1074 21563 -1067 21564
rect -1074 21542 -1070 21563
rect -1050 21542 -1046 21564
rect -1026 21542 -1022 21564
rect -1002 21542 -998 21564
rect -978 21542 -974 21564
rect -954 21542 -950 21564
rect -930 21542 -926 21564
rect -906 21542 -902 21564
rect -882 21542 -878 21564
rect -858 21542 -854 21564
rect -834 21542 -830 21564
rect -810 21542 -806 21564
rect -786 21542 -782 21564
rect -762 21542 -758 21564
rect -738 21542 -734 21564
rect -714 21542 -710 21564
rect -690 21542 -686 21564
rect -666 21542 -662 21564
rect -642 21542 -638 21564
rect -618 21542 -614 21564
rect -594 21542 -590 21564
rect -570 21542 -566 21564
rect -546 21542 -542 21564
rect -522 21542 -518 21564
rect -498 21542 -494 21564
rect -474 21542 -470 21564
rect -450 21542 -446 21564
rect -426 21542 -422 21564
rect -402 21542 -398 21564
rect -378 21542 -374 21564
rect -354 21542 -350 21564
rect -330 21542 -326 21564
rect -306 21542 -302 21564
rect -282 21542 -278 21564
rect -258 21542 -254 21564
rect -234 21542 -230 21564
rect -210 21542 -206 21564
rect -186 21542 -182 21564
rect -162 21542 -158 21564
rect -138 21542 -134 21564
rect -114 21542 -110 21564
rect -90 21542 -86 21564
rect -66 21542 -62 21564
rect -42 21542 -38 21564
rect -18 21542 -14 21564
rect 6 21542 10 21564
rect 30 21542 34 21564
rect 54 21542 58 21564
rect 78 21542 82 21564
rect 102 21542 106 21564
rect 126 21542 130 21564
rect 150 21542 154 21564
rect 174 21542 178 21564
rect 198 21542 202 21564
rect 222 21542 226 21564
rect 246 21542 250 21564
rect 270 21542 274 21564
rect 294 21542 298 21564
rect 318 21542 322 21564
rect 342 21542 346 21564
rect 366 21542 370 21564
rect 390 21542 394 21564
rect 414 21542 418 21564
rect 438 21542 442 21564
rect 462 21542 466 21564
rect 486 21542 490 21564
rect 510 21542 514 21564
rect 534 21542 538 21564
rect 558 21542 562 21564
rect 582 21542 586 21564
rect 606 21542 610 21564
rect 630 21542 634 21564
rect 654 21542 658 21564
rect 678 21542 682 21564
rect 702 21542 706 21564
rect 726 21542 730 21564
rect 750 21542 754 21564
rect 774 21542 778 21564
rect 798 21542 802 21564
rect 822 21542 826 21564
rect 846 21542 850 21564
rect 870 21542 874 21564
rect 894 21542 898 21564
rect 918 21542 922 21564
rect 942 21542 946 21564
rect 966 21542 970 21564
rect 990 21542 994 21564
rect 1014 21542 1018 21564
rect 1038 21542 1042 21564
rect 1062 21542 1066 21564
rect 1086 21542 1090 21564
rect 1110 21542 1114 21564
rect 1134 21542 1138 21564
rect 1158 21542 1162 21564
rect 1182 21542 1186 21564
rect 1206 21542 1210 21564
rect 1230 21542 1234 21564
rect 1254 21542 1258 21564
rect 1278 21542 1282 21564
rect 1302 21543 1306 21564
rect 1315 21557 1320 21564
rect 1326 21557 1330 21564
rect 1325 21543 1330 21557
rect 1291 21542 1349 21543
rect 1350 21542 1354 21588
rect 1374 21542 1378 21588
rect 1398 21542 1402 21588
rect -2393 21540 1419 21542
rect -2371 21470 -2366 21540
rect -2348 21470 -2343 21540
rect -2325 21528 -2320 21540
rect -2079 21538 -2071 21540
rect -2072 21536 -2071 21538
rect -2109 21531 -2101 21536
rect -2101 21529 -2079 21531
rect -2069 21529 -2068 21536
rect -2325 21520 -2317 21528
rect -2079 21524 -2071 21529
rect -2325 21470 -2320 21520
rect -2317 21512 -2309 21520
rect -2074 21515 -2071 21524
rect -2069 21520 -2068 21524
rect -2109 21506 -2079 21509
rect -2309 21472 -2301 21482
rect -2317 21470 -2309 21472
rect -2000 21470 -1992 21540
rect -1846 21538 -1806 21540
rect -1854 21533 -1806 21537
rect -1854 21531 -1846 21533
rect -1846 21529 -1806 21531
rect -1806 21527 -1798 21529
rect -1846 21524 -1798 21527
rect -1846 21511 -1806 21522
rect -1671 21520 -1663 21528
rect -1663 21512 -1655 21520
rect -1854 21506 -1680 21510
rect -1655 21472 -1647 21482
rect -1663 21470 -1655 21472
rect -1642 21470 -1637 21540
rect -1619 21470 -1614 21540
rect -1530 21470 -1526 21540
rect -1506 21470 -1502 21540
rect -1482 21470 -1478 21540
rect -1458 21470 -1454 21540
rect -1434 21470 -1430 21540
rect -1410 21470 -1406 21540
rect -1386 21470 -1382 21540
rect -1362 21470 -1358 21540
rect -1338 21470 -1334 21540
rect -1314 21470 -1310 21540
rect -1290 21470 -1286 21540
rect -1266 21470 -1262 21540
rect -1242 21470 -1238 21540
rect -1218 21470 -1214 21540
rect -1194 21470 -1190 21540
rect -1170 21470 -1166 21540
rect -1146 21470 -1142 21540
rect -1122 21470 -1118 21540
rect -1098 21470 -1094 21540
rect -1074 21470 -1070 21540
rect -1050 21470 -1046 21540
rect -1026 21470 -1022 21540
rect -1002 21470 -998 21540
rect -978 21470 -974 21540
rect -954 21470 -950 21540
rect -930 21470 -926 21540
rect -906 21470 -902 21540
rect -882 21470 -878 21540
rect -858 21470 -854 21540
rect -834 21470 -830 21540
rect -810 21470 -806 21540
rect -786 21470 -782 21540
rect -762 21470 -758 21540
rect -738 21470 -734 21540
rect -714 21470 -710 21540
rect -690 21470 -686 21540
rect -666 21470 -662 21540
rect -642 21470 -638 21540
rect -618 21470 -614 21540
rect -594 21470 -590 21540
rect -570 21470 -566 21540
rect -546 21470 -542 21540
rect -522 21470 -518 21540
rect -498 21470 -494 21540
rect -474 21470 -470 21540
rect -450 21470 -446 21540
rect -426 21470 -422 21540
rect -402 21470 -398 21540
rect -378 21470 -374 21540
rect -354 21470 -350 21540
rect -330 21470 -326 21540
rect -306 21470 -302 21540
rect -282 21470 -278 21540
rect -258 21470 -254 21540
rect -234 21470 -230 21540
rect -210 21470 -206 21540
rect -186 21470 -182 21540
rect -162 21470 -158 21540
rect -138 21470 -134 21540
rect -114 21470 -110 21540
rect -90 21470 -86 21540
rect -66 21470 -62 21540
rect -42 21470 -38 21540
rect -18 21470 -14 21540
rect 6 21470 10 21540
rect 30 21470 34 21540
rect 54 21470 58 21540
rect 78 21470 82 21540
rect 102 21470 106 21540
rect 126 21470 130 21540
rect 150 21470 154 21540
rect 174 21470 178 21540
rect 198 21470 202 21540
rect 222 21470 226 21540
rect 246 21470 250 21540
rect 270 21470 274 21540
rect 294 21470 298 21540
rect 318 21470 322 21540
rect 342 21470 346 21540
rect 366 21470 370 21540
rect 390 21470 394 21540
rect 414 21470 418 21540
rect 438 21470 442 21540
rect 462 21470 466 21540
rect 486 21470 490 21540
rect 510 21470 514 21540
rect 534 21470 538 21540
rect 558 21495 562 21540
rect 547 21494 581 21495
rect 582 21494 586 21540
rect 606 21494 610 21540
rect 630 21494 634 21540
rect 654 21494 658 21540
rect 678 21494 682 21540
rect 702 21494 706 21540
rect 726 21494 730 21540
rect 750 21494 754 21540
rect 774 21494 778 21540
rect 798 21494 802 21540
rect 822 21494 826 21540
rect 846 21494 850 21540
rect 870 21494 874 21540
rect 894 21494 898 21540
rect 918 21494 922 21540
rect 942 21494 946 21540
rect 966 21494 970 21540
rect 990 21494 994 21540
rect 1014 21494 1018 21540
rect 1038 21494 1042 21540
rect 1062 21494 1066 21540
rect 1086 21494 1090 21540
rect 1110 21494 1114 21540
rect 1134 21494 1138 21540
rect 1158 21494 1162 21540
rect 1182 21494 1186 21540
rect 1206 21494 1210 21540
rect 1230 21494 1234 21540
rect 1254 21494 1258 21540
rect 1278 21494 1282 21540
rect 1291 21533 1296 21540
rect 1302 21533 1306 21540
rect 1315 21533 1320 21540
rect 1301 21519 1306 21533
rect 1325 21519 1330 21533
rect 1291 21518 1325 21519
rect 1326 21518 1330 21519
rect 1350 21518 1354 21540
rect 1374 21518 1378 21540
rect 1398 21518 1402 21540
rect 1405 21539 1419 21540
rect 1422 21539 1429 21563
rect 1422 21518 1426 21539
rect 1446 21518 1450 21588
rect 1470 21518 1474 21588
rect 1494 21518 1498 21588
rect 1518 21518 1522 21588
rect 1542 21518 1546 21588
rect 1566 21518 1570 21588
rect 1590 21518 1594 21588
rect 1614 21518 1618 21588
rect 1638 21518 1642 21588
rect 1662 21518 1666 21588
rect 1686 21518 1690 21588
rect 1710 21518 1714 21588
rect 1734 21518 1738 21588
rect 1758 21518 1762 21588
rect 1782 21518 1786 21588
rect 1806 21518 1810 21588
rect 1830 21518 1834 21588
rect 1854 21518 1858 21588
rect 1878 21518 1882 21588
rect 1902 21518 1906 21588
rect 1926 21518 1930 21588
rect 1950 21518 1954 21588
rect 1974 21518 1978 21588
rect 1998 21518 2002 21588
rect 2022 21518 2026 21588
rect 2046 21518 2050 21588
rect 2070 21518 2074 21588
rect 2094 21518 2098 21588
rect 2118 21518 2122 21588
rect 2142 21518 2146 21588
rect 2166 21518 2170 21588
rect 2190 21518 2194 21588
rect 2214 21518 2218 21588
rect 2238 21518 2242 21588
rect 2262 21518 2266 21588
rect 2286 21518 2290 21588
rect 2310 21518 2314 21588
rect 2323 21581 2328 21588
rect 2334 21581 2338 21588
rect 2333 21567 2338 21581
rect 2323 21566 2357 21567
rect 2358 21566 2362 21612
rect 2371 21605 2376 21612
rect 2382 21605 2386 21612
rect 2381 21591 2386 21605
rect 2371 21590 2405 21591
rect 2406 21590 2410 21660
rect 2413 21659 2427 21660
rect 2430 21659 2437 21683
rect 2430 21590 2434 21659
rect 2454 21590 2458 21684
rect 2478 21590 2482 21684
rect 2502 21590 2506 21684
rect 2526 21590 2530 21684
rect 2550 21590 2554 21684
rect 2574 21590 2578 21684
rect 2598 21590 2602 21684
rect 2622 21590 2626 21684
rect 2646 21590 2650 21684
rect 2670 21590 2674 21684
rect 2694 21590 2698 21684
rect 2718 21662 2725 21683
rect 2742 21662 2746 21684
rect 2766 21662 2770 21684
rect 2790 21662 2794 21684
rect 2814 21662 2818 21684
rect 2862 21683 2866 21684
rect 2701 21660 2859 21662
rect 2701 21659 2715 21660
rect 2718 21659 2725 21660
rect 2718 21590 2722 21659
rect 2742 21590 2746 21660
rect 2766 21590 2770 21660
rect 2790 21590 2794 21660
rect 2814 21590 2818 21660
rect 2845 21659 2859 21660
rect 2862 21659 2869 21683
rect 2827 21638 2861 21639
rect 2886 21638 2890 21684
rect 2910 21638 2914 21684
rect 2934 21638 2938 21684
rect 2958 21639 2962 21684
rect 2947 21638 2981 21639
rect 2827 21636 2981 21638
rect 2827 21629 2832 21636
rect 2837 21615 2842 21629
rect 2838 21590 2842 21615
rect 2886 21590 2890 21636
rect 2910 21590 2914 21636
rect 2934 21590 2938 21636
rect 2947 21629 2952 21636
rect 2958 21629 2962 21636
rect 2957 21615 2962 21629
rect 2947 21614 2981 21615
rect 2982 21614 2986 21684
rect 3006 21614 3010 21684
rect 3030 21614 3034 21684
rect 3078 21683 3082 21684
rect 3078 21662 3085 21683
rect 3102 21662 3106 21684
rect 3126 21662 3130 21684
rect 3061 21660 3147 21662
rect 3061 21659 3075 21660
rect 3078 21659 3085 21660
rect 3043 21638 3077 21639
rect 3102 21638 3106 21660
rect 3126 21638 3130 21660
rect 3133 21659 3147 21660
rect 3150 21659 3157 21683
rect 3150 21638 3154 21659
rect 3174 21638 3178 21684
rect 3198 21638 3202 21684
rect 3222 21638 3226 21684
rect 3270 21683 3274 21684
rect 3270 21662 3277 21683
rect 3283 21677 3288 21684
rect 3301 21683 3315 21684
rect 3829 21683 3843 21684
rect 3846 21683 3853 21684
rect 3859 21677 3864 21684
rect 3877 21683 3891 21684
rect 4549 21683 4563 21684
rect 4566 21683 4573 21684
rect 4579 21677 4584 21684
rect 4597 21683 4611 21684
rect 4789 21683 4803 21684
rect 4806 21683 4813 21684
rect 4819 21677 4824 21684
rect 4837 21683 4851 21684
rect 6589 21683 6603 21684
rect 6606 21683 6613 21684
rect 3293 21663 3298 21677
rect 3307 21673 3315 21677
rect 3301 21663 3307 21673
rect 3389 21663 3394 21677
rect 3869 21663 3874 21677
rect 4589 21663 4594 21677
rect 4829 21663 4834 21677
rect 3283 21662 3317 21663
rect 3253 21660 3317 21662
rect 3331 21660 3365 21663
rect 3253 21659 3267 21660
rect 3270 21659 3277 21660
rect 3283 21653 3288 21660
rect 3301 21659 3315 21660
rect 3293 21639 3298 21653
rect 3307 21649 3315 21653
rect 3355 21649 3363 21653
rect 3301 21639 3307 21649
rect 3349 21639 3355 21649
rect 3283 21638 3317 21639
rect 3043 21636 3317 21638
rect 3331 21638 3365 21639
rect 3366 21638 3373 21659
rect 3379 21653 3384 21663
rect 3389 21639 3394 21653
rect 3403 21649 3411 21653
rect 3835 21649 3843 21653
rect 3397 21639 3403 21649
rect 3829 21639 3835 21649
rect 3379 21638 3413 21639
rect 3331 21636 3413 21638
rect 3811 21638 3845 21639
rect 3846 21638 3853 21659
rect 3859 21653 3864 21663
rect 3869 21639 3874 21653
rect 3883 21649 3891 21653
rect 4555 21649 4563 21653
rect 3877 21639 3883 21649
rect 4549 21639 4555 21649
rect 3859 21638 3893 21639
rect 3811 21636 3893 21638
rect 4531 21638 4565 21639
rect 4566 21638 4573 21659
rect 4579 21653 4584 21663
rect 4589 21639 4594 21653
rect 4603 21649 4611 21653
rect 4795 21649 4803 21653
rect 4597 21639 4603 21649
rect 4789 21639 4795 21649
rect 4579 21638 4613 21639
rect 4531 21636 4613 21638
rect 4771 21638 4805 21639
rect 4806 21638 4813 21659
rect 4819 21653 4824 21663
rect 4829 21639 4834 21653
rect 4843 21649 4851 21653
rect 6595 21649 6603 21653
rect 4837 21639 4843 21649
rect 6589 21639 6595 21649
rect 4819 21638 4853 21639
rect 4771 21636 4853 21638
rect 6571 21638 6605 21639
rect 6606 21638 6613 21659
rect 6630 21638 6634 21684
rect 6637 21683 6651 21684
rect 6685 21683 6699 21684
rect 6702 21683 6709 21684
rect 6678 21662 6685 21683
rect 6702 21662 6706 21683
rect 6726 21662 6730 21684
rect 6750 21662 6754 21684
rect 6774 21662 6778 21684
rect 6798 21662 6802 21684
rect 6822 21662 6826 21684
rect 6846 21662 6850 21684
rect 6870 21662 6874 21684
rect 6894 21662 6898 21684
rect 6918 21662 6922 21684
rect 6942 21662 6946 21684
rect 6966 21662 6970 21684
rect 7038 21662 7042 21684
rect 7099 21677 7104 21684
rect 7117 21683 7131 21684
rect 7525 21683 7538 21684
rect 7109 21663 7114 21677
rect 7123 21673 7131 21677
rect 7117 21663 7123 21673
rect 7542 21664 7549 21708
rect 7555 21701 7560 21708
rect 7573 21707 7587 21708
rect 8269 21707 8283 21708
rect 8317 21707 8331 21708
rect 14533 21707 14547 21708
rect 7565 21687 7570 21701
rect 7579 21697 7587 21701
rect 7573 21687 7579 21697
rect 8285 21687 8290 21701
rect 14539 21697 14547 21701
rect 14533 21687 14539 21697
rect 8227 21684 8261 21687
rect 7573 21683 7587 21684
rect 8251 21673 8259 21677
rect 8245 21663 8251 21673
rect 7099 21662 7133 21663
rect 6661 21660 7133 21662
rect 7483 21660 7517 21663
rect 7531 21662 7565 21663
rect 7525 21660 7565 21662
rect 8227 21662 8261 21663
rect 8262 21662 8269 21683
rect 8275 21677 8280 21687
rect 8294 21684 8309 21687
rect 14515 21686 14549 21687
rect 14550 21686 14557 21708
rect 14563 21701 14568 21708
rect 14581 21707 14595 21708
rect 14773 21707 14787 21708
rect 14821 21707 14835 21708
rect 14573 21687 14578 21701
rect 14587 21697 14595 21701
rect 14581 21687 14587 21697
rect 14789 21687 14797 21701
rect 14995 21697 15003 21701
rect 14989 21687 14995 21697
rect 14563 21686 14597 21687
rect 14515 21684 14597 21686
rect 14731 21684 14765 21687
rect 14779 21686 14813 21687
rect 14773 21684 14813 21686
rect 14971 21686 15005 21687
rect 15006 21686 15013 21707
rect 15019 21701 15024 21711
rect 15038 21708 15053 21711
rect 15211 21708 15245 21711
rect 15259 21708 15278 21711
rect 15029 21687 15034 21701
rect 15043 21697 15051 21701
rect 15037 21687 15043 21697
rect 15269 21687 15274 21701
rect 15019 21686 15053 21687
rect 14971 21684 15053 21686
rect 15211 21684 15245 21687
rect 14533 21683 14547 21684
rect 8285 21663 8290 21677
rect 8299 21673 8307 21677
rect 14539 21673 14547 21677
rect 8293 21663 8299 21673
rect 14533 21663 14539 21673
rect 8275 21662 8309 21663
rect 8227 21660 8309 21662
rect 14515 21662 14549 21663
rect 14550 21662 14557 21684
rect 14563 21677 14568 21684
rect 14581 21683 14595 21684
rect 14773 21683 14787 21684
rect 14821 21683 14835 21684
rect 14989 21683 15003 21684
rect 14573 21663 14578 21677
rect 14587 21673 14595 21677
rect 14581 21663 14587 21673
rect 14789 21663 14794 21677
rect 14995 21673 15003 21677
rect 14989 21663 14995 21673
rect 14563 21662 14597 21663
rect 14515 21660 14597 21662
rect 14731 21660 14765 21663
rect 6661 21659 6675 21660
rect 6678 21659 6685 21660
rect 6702 21638 6706 21660
rect 6726 21638 6730 21660
rect 6750 21638 6754 21660
rect 6774 21638 6778 21660
rect 6798 21638 6802 21660
rect 6822 21638 6826 21660
rect 6846 21638 6850 21660
rect 6870 21638 6874 21660
rect 6894 21638 6898 21660
rect 6918 21638 6922 21660
rect 6942 21638 6946 21660
rect 6966 21638 6970 21660
rect 7038 21638 7042 21660
rect 7099 21653 7104 21660
rect 7117 21659 7131 21660
rect 7525 21659 7539 21660
rect 7573 21659 7587 21660
rect 8245 21659 8259 21660
rect 7109 21639 7114 21653
rect 7123 21649 7131 21653
rect 7117 21639 7123 21649
rect 7541 21639 7549 21653
rect 8251 21649 8259 21653
rect 8245 21639 8251 21649
rect 7099 21638 7133 21639
rect 6571 21636 7133 21638
rect 7483 21636 7517 21639
rect 7531 21638 7565 21639
rect 7525 21636 7565 21638
rect 8227 21638 8261 21639
rect 8262 21638 8269 21660
rect 8275 21653 8280 21660
rect 8293 21659 8307 21660
rect 14533 21659 14547 21660
rect 8285 21639 8290 21653
rect 8299 21649 8307 21653
rect 14539 21649 14547 21653
rect 8293 21639 8299 21649
rect 14533 21639 14539 21649
rect 8275 21638 8309 21639
rect 8227 21636 8309 21638
rect 3043 21629 3048 21636
rect 3053 21615 3058 21629
rect 3054 21614 3058 21615
rect 3102 21614 3106 21636
rect 3126 21614 3130 21636
rect 3150 21614 3154 21636
rect 3174 21614 3178 21636
rect 3198 21614 3202 21636
rect 3222 21614 3226 21636
rect 3283 21629 3288 21636
rect 3301 21635 3315 21636
rect 3349 21635 3363 21636
rect 3293 21615 3298 21629
rect 3307 21625 3315 21629
rect 3355 21625 3363 21629
rect 3301 21615 3307 21625
rect 3349 21615 3355 21625
rect 3283 21614 3317 21615
rect 2947 21612 3317 21614
rect 3331 21614 3365 21615
rect 3366 21614 3373 21636
rect 3379 21629 3384 21636
rect 3397 21635 3411 21636
rect 3829 21635 3843 21636
rect 3389 21615 3394 21629
rect 3403 21625 3411 21629
rect 3835 21625 3843 21629
rect 3397 21615 3403 21625
rect 3829 21615 3835 21625
rect 3379 21614 3413 21615
rect 3331 21612 3413 21614
rect 3811 21614 3845 21615
rect 3846 21614 3853 21636
rect 3859 21629 3864 21636
rect 3877 21635 3891 21636
rect 4549 21635 4563 21636
rect 3869 21615 3874 21629
rect 3883 21625 3891 21629
rect 4555 21625 4563 21629
rect 3877 21615 3883 21625
rect 4549 21615 4555 21625
rect 3859 21614 3893 21615
rect 3811 21612 3893 21614
rect 4531 21614 4565 21615
rect 4566 21614 4573 21636
rect 4579 21629 4584 21636
rect 4597 21635 4611 21636
rect 4789 21635 4803 21636
rect 4589 21615 4594 21629
rect 4603 21625 4611 21629
rect 4795 21625 4803 21629
rect 4597 21615 4603 21625
rect 4789 21615 4795 21625
rect 4579 21614 4613 21615
rect 4531 21612 4613 21614
rect 4771 21614 4805 21615
rect 4806 21614 4813 21636
rect 4819 21629 4824 21636
rect 4837 21635 4851 21636
rect 6589 21635 6603 21636
rect 4829 21615 4834 21629
rect 4843 21625 4851 21629
rect 6595 21625 6603 21629
rect 4837 21615 4843 21625
rect 6589 21615 6595 21625
rect 4819 21614 4853 21615
rect 4771 21612 4853 21614
rect 6571 21614 6605 21615
rect 6606 21614 6613 21636
rect 6630 21614 6634 21636
rect 6643 21614 6677 21615
rect 6571 21612 6677 21614
rect 2947 21605 2952 21612
rect 2957 21591 2962 21605
rect 2958 21590 2962 21591
rect 2982 21590 2986 21612
rect 3006 21590 3010 21612
rect 3030 21590 3034 21612
rect 3054 21590 3058 21612
rect 3102 21590 3106 21612
rect 3126 21590 3130 21612
rect 3150 21590 3154 21612
rect 3174 21590 3178 21612
rect 3198 21590 3202 21612
rect 3222 21590 3226 21612
rect 3283 21605 3288 21612
rect 3301 21611 3315 21612
rect 3349 21611 3363 21612
rect 3293 21591 3298 21605
rect 3307 21601 3315 21605
rect 3355 21601 3363 21605
rect 3301 21591 3307 21601
rect 3349 21591 3355 21601
rect 3283 21590 3317 21591
rect 2371 21588 3317 21590
rect 3331 21590 3365 21591
rect 3366 21590 3373 21612
rect 3379 21605 3384 21612
rect 3397 21611 3411 21612
rect 3829 21611 3843 21612
rect 3389 21591 3394 21605
rect 3403 21601 3411 21605
rect 3835 21601 3843 21605
rect 3397 21591 3403 21601
rect 3829 21591 3835 21601
rect 3379 21590 3413 21591
rect 3331 21588 3413 21590
rect 3811 21590 3845 21591
rect 3846 21590 3853 21612
rect 3859 21605 3864 21612
rect 3877 21611 3891 21612
rect 4549 21611 4563 21612
rect 3869 21591 3874 21605
rect 3883 21601 3891 21605
rect 4555 21601 4563 21605
rect 3877 21591 3883 21601
rect 4549 21591 4555 21601
rect 3859 21590 3893 21591
rect 3811 21588 3893 21590
rect 4531 21590 4565 21591
rect 4566 21590 4573 21612
rect 4579 21605 4584 21612
rect 4597 21611 4611 21612
rect 4789 21611 4803 21612
rect 4589 21591 4594 21605
rect 4603 21601 4611 21605
rect 4795 21601 4803 21605
rect 4597 21591 4603 21601
rect 4789 21591 4795 21601
rect 4579 21590 4613 21591
rect 4531 21588 4613 21590
rect 4771 21590 4805 21591
rect 4806 21590 4813 21612
rect 4819 21605 4824 21612
rect 4837 21611 4851 21612
rect 6589 21611 6603 21612
rect 4829 21591 4834 21605
rect 4843 21601 4851 21605
rect 6595 21601 6603 21605
rect 4837 21591 4843 21601
rect 6589 21591 6595 21601
rect 4819 21590 4853 21591
rect 4771 21588 4853 21590
rect 6571 21590 6605 21591
rect 6606 21590 6613 21612
rect 6630 21591 6634 21612
rect 6643 21605 6648 21612
rect 6653 21591 6658 21605
rect 6619 21590 6653 21591
rect 6571 21588 6653 21590
rect 6667 21590 6701 21591
rect 6702 21590 6706 21636
rect 6726 21590 6730 21636
rect 6750 21590 6754 21636
rect 6774 21590 6778 21636
rect 6798 21590 6802 21636
rect 6822 21590 6826 21636
rect 6846 21590 6850 21636
rect 6870 21590 6874 21636
rect 6894 21590 6898 21636
rect 6918 21590 6922 21636
rect 6942 21590 6946 21636
rect 6966 21590 6970 21636
rect 6979 21614 7013 21615
rect 7038 21614 7042 21636
rect 7099 21629 7104 21636
rect 7117 21635 7131 21636
rect 7525 21635 7539 21636
rect 7573 21635 7587 21636
rect 8245 21635 8259 21636
rect 7109 21615 7114 21629
rect 7123 21625 7131 21629
rect 7117 21615 7123 21625
rect 7541 21615 7549 21629
rect 8251 21625 8259 21629
rect 8245 21615 8251 21625
rect 7099 21614 7133 21615
rect 6979 21612 7133 21614
rect 7483 21612 7517 21615
rect 7531 21614 7565 21615
rect 7525 21612 7565 21614
rect 8227 21614 8261 21615
rect 8262 21614 8269 21636
rect 8275 21629 8280 21636
rect 8293 21635 8307 21636
rect 14533 21635 14546 21636
rect 8285 21615 8290 21629
rect 8299 21625 8307 21629
rect 8293 21615 8299 21625
rect 14550 21616 14557 21660
rect 14563 21653 14568 21660
rect 14581 21659 14595 21660
rect 14573 21639 14578 21653
rect 14587 21649 14595 21653
rect 14755 21649 14763 21653
rect 14581 21639 14587 21649
rect 14749 21639 14755 21649
rect 14731 21638 14765 21639
rect 14766 21638 14773 21659
rect 14779 21653 14784 21663
rect 14798 21660 14813 21663
rect 14971 21662 15005 21663
rect 15006 21662 15013 21684
rect 15019 21677 15024 21684
rect 15037 21683 15051 21684
rect 15029 21663 15034 21677
rect 15043 21673 15051 21677
rect 15235 21673 15243 21677
rect 15037 21663 15043 21673
rect 15229 21663 15235 21673
rect 15019 21662 15053 21663
rect 14971 21660 15053 21662
rect 15211 21662 15245 21663
rect 15246 21662 15253 21683
rect 15259 21677 15264 21687
rect 15278 21684 15293 21687
rect 15691 21684 15725 21687
rect 15739 21684 15773 21687
rect 15269 21663 15274 21677
rect 15283 21673 15291 21677
rect 15277 21663 15283 21673
rect 15259 21662 15293 21663
rect 15211 21660 15293 21662
rect 15691 21660 15725 21663
rect 15739 21660 15758 21663
rect 15931 21660 15965 21663
rect 15979 21660 16013 21663
rect 14989 21659 15003 21660
rect 14789 21639 14794 21653
rect 14803 21649 14811 21653
rect 14995 21649 15003 21653
rect 14797 21639 14803 21649
rect 14989 21639 14995 21649
rect 14779 21638 14813 21639
rect 14731 21636 14813 21638
rect 14971 21638 15005 21639
rect 15006 21638 15013 21660
rect 15019 21653 15024 21660
rect 15037 21659 15051 21660
rect 15229 21659 15243 21660
rect 15029 21639 15034 21653
rect 15043 21649 15051 21653
rect 15235 21649 15243 21653
rect 15037 21639 15043 21649
rect 15229 21639 15235 21649
rect 15019 21638 15053 21639
rect 14971 21636 15053 21638
rect 15211 21638 15245 21639
rect 15246 21638 15253 21660
rect 15259 21653 15264 21660
rect 15277 21659 15291 21660
rect 15269 21639 15274 21653
rect 15283 21649 15291 21653
rect 15277 21639 15283 21649
rect 15749 21639 15754 21653
rect 15259 21638 15293 21639
rect 15211 21636 15293 21638
rect 15691 21636 15725 21639
rect 14581 21635 14595 21636
rect 14749 21635 14763 21636
rect 14755 21625 14763 21629
rect 14749 21615 14755 21625
rect 8275 21614 8309 21615
rect 8227 21612 8309 21614
rect 14491 21612 14525 21615
rect 14539 21614 14573 21615
rect 14533 21612 14573 21614
rect 14731 21614 14765 21615
rect 14766 21614 14773 21636
rect 14779 21629 14784 21636
rect 14797 21635 14811 21636
rect 14989 21635 15003 21636
rect 14789 21615 14794 21629
rect 14803 21625 14811 21629
rect 14995 21625 15003 21629
rect 14797 21615 14803 21625
rect 14989 21615 14995 21625
rect 14779 21614 14813 21615
rect 14731 21612 14813 21614
rect 14971 21614 15005 21615
rect 15006 21614 15013 21636
rect 15019 21629 15024 21636
rect 15037 21635 15051 21636
rect 15229 21635 15243 21636
rect 15029 21615 15034 21629
rect 15043 21625 15051 21629
rect 15235 21625 15243 21629
rect 15037 21615 15043 21625
rect 15229 21615 15235 21625
rect 15019 21614 15053 21615
rect 14971 21612 15053 21614
rect 15211 21614 15245 21615
rect 15246 21614 15253 21636
rect 15259 21629 15264 21636
rect 15277 21635 15291 21636
rect 15269 21615 15274 21629
rect 15283 21625 15291 21629
rect 15715 21625 15723 21629
rect 15277 21615 15283 21625
rect 15709 21615 15715 21625
rect 15259 21614 15293 21615
rect 15211 21612 15293 21614
rect 15691 21614 15725 21615
rect 15726 21614 15733 21635
rect 15739 21629 15744 21639
rect 15758 21636 15773 21639
rect 15931 21636 15965 21639
rect 15979 21636 15998 21639
rect 16171 21636 16205 21639
rect 16219 21636 16238 21639
rect 15749 21615 15754 21629
rect 15763 21625 15771 21629
rect 15757 21615 15763 21625
rect 15989 21615 15994 21629
rect 16229 21615 16234 21629
rect 15739 21614 15773 21615
rect 15691 21612 15773 21614
rect 15931 21612 15965 21615
rect 6979 21605 6984 21612
rect 6989 21591 6994 21605
rect 6990 21590 6994 21591
rect 7038 21590 7042 21612
rect 7099 21605 7104 21612
rect 7117 21611 7131 21612
rect 7525 21611 7539 21612
rect 7573 21611 7587 21612
rect 8245 21611 8259 21612
rect 7109 21591 7114 21605
rect 7123 21601 7131 21605
rect 7117 21591 7123 21601
rect 7541 21591 7546 21605
rect 8251 21601 8259 21605
rect 8245 21591 8251 21601
rect 7099 21590 7133 21591
rect 6667 21588 7133 21590
rect 7483 21588 7517 21591
rect 2371 21581 2376 21588
rect 2381 21567 2386 21581
rect 2382 21566 2386 21567
rect 2406 21566 2410 21588
rect 2430 21566 2434 21588
rect 2454 21566 2458 21588
rect 2478 21566 2482 21588
rect 2502 21566 2506 21588
rect 2526 21566 2530 21588
rect 2550 21566 2554 21588
rect 2574 21566 2578 21588
rect 2598 21566 2602 21588
rect 2622 21566 2626 21588
rect 2646 21566 2650 21588
rect 2670 21566 2674 21588
rect 2694 21566 2698 21588
rect 2718 21566 2722 21588
rect 2742 21566 2746 21588
rect 2766 21566 2770 21588
rect 2790 21566 2794 21588
rect 2814 21566 2818 21588
rect 2838 21566 2842 21588
rect 2886 21566 2890 21588
rect 2910 21566 2914 21588
rect 2934 21566 2938 21588
rect 2958 21566 2962 21588
rect 2982 21566 2986 21588
rect 3006 21566 3010 21588
rect 3030 21566 3034 21588
rect 3054 21566 3058 21588
rect 3102 21566 3106 21588
rect 3126 21566 3130 21588
rect 3150 21566 3154 21588
rect 3174 21566 3178 21588
rect 3198 21566 3202 21588
rect 3222 21566 3226 21588
rect 3283 21581 3288 21588
rect 3301 21587 3315 21588
rect 3349 21587 3363 21588
rect 3293 21567 3298 21581
rect 3307 21577 3315 21581
rect 3355 21577 3363 21581
rect 3301 21567 3307 21577
rect 3349 21567 3355 21577
rect 3283 21566 3317 21567
rect 2323 21564 3317 21566
rect 3331 21566 3365 21567
rect 3366 21566 3373 21588
rect 3379 21581 3384 21588
rect 3397 21587 3411 21588
rect 3829 21587 3843 21588
rect 3389 21567 3394 21581
rect 3403 21577 3411 21581
rect 3835 21577 3843 21581
rect 3397 21567 3403 21577
rect 3829 21567 3835 21577
rect 3379 21566 3413 21567
rect 3331 21564 3413 21566
rect 3811 21566 3845 21567
rect 3846 21566 3853 21588
rect 3859 21581 3864 21588
rect 3877 21587 3891 21588
rect 4549 21587 4563 21588
rect 3869 21567 3874 21581
rect 3883 21577 3891 21581
rect 4555 21577 4563 21581
rect 3877 21567 3883 21577
rect 4549 21567 4555 21577
rect 3859 21566 3893 21567
rect 3811 21564 3893 21566
rect 4531 21566 4565 21567
rect 4566 21566 4573 21588
rect 4579 21581 4584 21588
rect 4597 21587 4611 21588
rect 4789 21587 4803 21588
rect 4589 21567 4594 21581
rect 4603 21577 4611 21581
rect 4795 21577 4803 21581
rect 4597 21567 4603 21577
rect 4789 21567 4795 21577
rect 4579 21566 4613 21567
rect 4531 21564 4613 21566
rect 4771 21566 4805 21567
rect 4806 21566 4813 21588
rect 4819 21581 4824 21588
rect 4837 21587 4851 21588
rect 6589 21587 6603 21588
rect 4829 21567 4834 21581
rect 4843 21577 4851 21581
rect 6595 21577 6603 21581
rect 4837 21567 4843 21577
rect 6589 21567 6595 21577
rect 4819 21566 4853 21567
rect 4771 21564 4853 21566
rect 6571 21566 6605 21567
rect 6606 21566 6613 21588
rect 6619 21581 6624 21588
rect 6630 21581 6634 21588
rect 6629 21567 6634 21581
rect 6644 21578 6648 21588
rect 6654 21566 6658 21578
rect 6702 21566 6706 21588
rect 6726 21566 6730 21588
rect 6750 21566 6754 21588
rect 6774 21566 6778 21588
rect 6798 21566 6802 21588
rect 6822 21566 6826 21588
rect 6846 21566 6850 21588
rect 6870 21566 6874 21588
rect 6894 21566 6898 21588
rect 6918 21566 6922 21588
rect 6942 21566 6946 21588
rect 6966 21566 6970 21588
rect 6990 21566 6994 21588
rect 7038 21566 7042 21588
rect 7099 21581 7104 21588
rect 7117 21587 7131 21588
rect 7109 21567 7114 21581
rect 7123 21577 7131 21581
rect 7507 21577 7515 21581
rect 7117 21567 7123 21577
rect 7501 21567 7507 21577
rect 7099 21566 7133 21567
rect 6571 21564 7133 21566
rect 7483 21566 7517 21567
rect 7518 21566 7525 21587
rect 7531 21581 7536 21591
rect 7550 21588 7565 21591
rect 8227 21590 8261 21591
rect 8262 21590 8269 21612
rect 8275 21605 8280 21612
rect 8293 21611 8307 21612
rect 14533 21611 14547 21612
rect 14581 21611 14595 21612
rect 14749 21611 14763 21612
rect 8285 21591 8290 21605
rect 8299 21601 8307 21605
rect 8293 21591 8299 21601
rect 14549 21591 14557 21605
rect 14755 21601 14763 21605
rect 14749 21591 14755 21601
rect 8275 21590 8309 21591
rect 8227 21588 8309 21590
rect 14491 21588 14525 21591
rect 14539 21590 14573 21591
rect 14533 21588 14573 21590
rect 14731 21590 14765 21591
rect 14766 21590 14773 21612
rect 14779 21605 14784 21612
rect 14797 21611 14811 21612
rect 14989 21611 15003 21612
rect 14789 21591 14794 21605
rect 14803 21601 14811 21605
rect 14995 21601 15003 21605
rect 14797 21591 14803 21601
rect 14989 21591 14995 21601
rect 14779 21590 14813 21591
rect 14731 21588 14813 21590
rect 14971 21590 15005 21591
rect 15006 21590 15013 21612
rect 15019 21605 15024 21612
rect 15037 21611 15051 21612
rect 15229 21611 15243 21612
rect 15029 21591 15034 21605
rect 15043 21601 15051 21605
rect 15235 21601 15243 21605
rect 15037 21591 15043 21601
rect 15229 21591 15235 21601
rect 15019 21590 15053 21591
rect 14971 21588 15053 21590
rect 15211 21590 15245 21591
rect 15246 21590 15253 21612
rect 15259 21605 15264 21612
rect 15277 21611 15291 21612
rect 15709 21611 15723 21612
rect 15269 21591 15274 21605
rect 15283 21601 15291 21605
rect 15715 21601 15723 21605
rect 15277 21591 15283 21601
rect 15709 21591 15715 21601
rect 15259 21590 15293 21591
rect 15211 21588 15293 21590
rect 15691 21590 15725 21591
rect 15726 21590 15733 21612
rect 15739 21605 15744 21612
rect 15757 21611 15771 21612
rect 15749 21591 15754 21605
rect 15763 21601 15771 21605
rect 15955 21601 15963 21605
rect 15757 21591 15763 21601
rect 15949 21591 15955 21601
rect 15739 21590 15773 21591
rect 15691 21588 15773 21590
rect 15931 21590 15965 21591
rect 15966 21590 15973 21611
rect 15979 21605 15984 21615
rect 15998 21612 16013 21615
rect 16171 21612 16205 21615
rect 15989 21591 15994 21605
rect 16003 21601 16011 21605
rect 16195 21601 16203 21605
rect 15997 21591 16003 21601
rect 16189 21591 16195 21601
rect 15979 21590 16013 21591
rect 15931 21588 16013 21590
rect 16171 21590 16205 21591
rect 16206 21590 16213 21611
rect 16219 21605 16224 21615
rect 16238 21612 16253 21615
rect 16363 21612 16397 21615
rect 16411 21612 16430 21615
rect 16229 21591 16234 21605
rect 16243 21601 16251 21605
rect 16237 21591 16243 21601
rect 16421 21591 16426 21605
rect 16219 21590 16253 21591
rect 16171 21588 16253 21590
rect 16363 21588 16397 21591
rect 8245 21587 8259 21588
rect 7541 21567 7546 21581
rect 7555 21577 7563 21581
rect 8251 21577 8259 21581
rect 7549 21567 7555 21577
rect 8245 21567 8251 21577
rect 7531 21566 7565 21567
rect 7483 21564 7565 21566
rect 8227 21566 8261 21567
rect 8262 21566 8269 21588
rect 8275 21581 8280 21588
rect 8293 21587 8307 21588
rect 14533 21587 14547 21588
rect 14581 21587 14595 21588
rect 14749 21587 14763 21588
rect 8285 21567 8290 21581
rect 8299 21577 8307 21581
rect 8293 21567 8299 21577
rect 14549 21567 14557 21581
rect 14755 21577 14763 21581
rect 14749 21567 14755 21577
rect 8275 21566 8309 21567
rect 8227 21564 8309 21566
rect 14491 21564 14525 21567
rect 14539 21566 14573 21567
rect 14533 21564 14573 21566
rect 14731 21566 14765 21567
rect 14766 21566 14773 21588
rect 14779 21581 14784 21588
rect 14797 21587 14811 21588
rect 14989 21587 15003 21588
rect 14789 21567 14794 21581
rect 14803 21577 14811 21581
rect 14995 21577 15003 21581
rect 14797 21567 14803 21577
rect 14989 21567 14995 21577
rect 14779 21566 14813 21567
rect 14731 21564 14813 21566
rect 14971 21566 15005 21567
rect 15006 21566 15013 21588
rect 15019 21581 15024 21588
rect 15037 21587 15051 21588
rect 15229 21587 15243 21588
rect 15029 21567 15034 21581
rect 15043 21577 15051 21581
rect 15235 21577 15243 21581
rect 15037 21567 15043 21577
rect 15229 21567 15235 21577
rect 15019 21566 15053 21567
rect 14971 21564 15053 21566
rect 15211 21566 15245 21567
rect 15246 21566 15253 21588
rect 15259 21581 15264 21588
rect 15277 21587 15291 21588
rect 15709 21587 15723 21588
rect 15269 21567 15274 21581
rect 15283 21577 15291 21581
rect 15715 21577 15723 21581
rect 15277 21567 15283 21577
rect 15709 21567 15715 21577
rect 15259 21566 15293 21567
rect 15211 21564 15293 21566
rect 15691 21566 15725 21567
rect 15726 21566 15733 21588
rect 15739 21581 15744 21588
rect 15757 21587 15771 21588
rect 15949 21587 15963 21588
rect 15749 21567 15754 21581
rect 15763 21577 15771 21581
rect 15955 21577 15963 21581
rect 15757 21567 15763 21577
rect 15949 21567 15955 21577
rect 15739 21566 15773 21567
rect 15691 21564 15773 21566
rect 15931 21566 15965 21567
rect 15966 21566 15973 21588
rect 15979 21581 15984 21588
rect 15997 21587 16011 21588
rect 16189 21587 16203 21588
rect 15989 21567 15994 21581
rect 16003 21577 16011 21581
rect 16195 21577 16203 21581
rect 15997 21567 16003 21577
rect 16189 21567 16195 21577
rect 15979 21566 16013 21567
rect 15931 21564 16013 21566
rect 16171 21566 16205 21567
rect 16206 21566 16213 21588
rect 16219 21581 16224 21588
rect 16237 21587 16251 21588
rect 16229 21567 16234 21581
rect 16243 21577 16251 21581
rect 16387 21577 16395 21581
rect 16237 21567 16243 21577
rect 16381 21567 16387 21577
rect 16219 21566 16253 21567
rect 16171 21564 16253 21566
rect 16363 21566 16397 21567
rect 16398 21566 16405 21587
rect 16411 21581 16416 21591
rect 16430 21588 16445 21591
rect 25771 21588 25805 21591
rect 25819 21588 25838 21591
rect 16421 21567 16426 21581
rect 16435 21577 16443 21581
rect 16429 21567 16435 21577
rect 25829 21567 25834 21581
rect 16411 21566 16445 21567
rect 16363 21564 16445 21566
rect 25771 21564 25805 21567
rect 2323 21557 2328 21564
rect 2333 21543 2338 21557
rect 2334 21518 2338 21543
rect 2358 21518 2362 21564
rect 2382 21518 2386 21564
rect 2406 21539 2410 21564
rect 1291 21516 2403 21518
rect 1291 21509 1296 21516
rect 1301 21495 1306 21509
rect 1302 21494 1306 21495
rect 1326 21494 1330 21516
rect 1350 21494 1354 21516
rect 1374 21494 1378 21516
rect 1398 21494 1402 21516
rect 1422 21494 1426 21516
rect 1446 21494 1450 21516
rect 1470 21494 1474 21516
rect 1494 21494 1498 21516
rect 1518 21494 1522 21516
rect 1542 21494 1546 21516
rect 1566 21494 1570 21516
rect 1590 21494 1594 21516
rect 1614 21494 1618 21516
rect 1638 21494 1642 21516
rect 1662 21494 1666 21516
rect 1686 21494 1690 21516
rect 1710 21494 1714 21516
rect 1734 21494 1738 21516
rect 1758 21494 1762 21516
rect 1782 21494 1786 21516
rect 1806 21494 1810 21516
rect 1830 21494 1834 21516
rect 1854 21494 1858 21516
rect 1878 21494 1882 21516
rect 1902 21494 1906 21516
rect 1926 21494 1930 21516
rect 1950 21494 1954 21516
rect 1974 21494 1978 21516
rect 1998 21494 2002 21516
rect 2022 21494 2026 21516
rect 2046 21494 2050 21516
rect 2070 21494 2074 21516
rect 2094 21494 2098 21516
rect 2118 21494 2122 21516
rect 2142 21494 2146 21516
rect 2166 21494 2170 21516
rect 2190 21494 2194 21516
rect 2214 21494 2218 21516
rect 2238 21494 2242 21516
rect 2262 21494 2266 21516
rect 2286 21494 2290 21516
rect 2310 21494 2314 21516
rect 2334 21494 2338 21516
rect 2358 21515 2362 21516
rect 547 21492 2355 21494
rect 547 21485 552 21492
rect 558 21485 562 21492
rect 557 21471 562 21485
rect 547 21470 581 21471
rect -2393 21468 581 21470
rect -2371 21374 -2366 21468
rect -2348 21374 -2343 21468
rect -2325 21406 -2320 21468
rect -2317 21466 -2309 21468
rect -2013 21466 -1992 21468
rect -1663 21466 -1655 21468
rect -2000 21465 -1983 21466
rect -2026 21456 -2021 21460
rect -2062 21455 -2061 21456
rect -2309 21444 -2301 21454
rect -2091 21448 -2061 21455
rect -2317 21438 -2309 21444
rect -2132 21439 -2131 21441
rect -2101 21439 -2092 21441
rect -2091 21440 -2071 21446
rect -2062 21444 -2045 21448
rect -2036 21444 -2031 21446
rect -2292 21430 -2071 21439
rect -2107 21425 -2104 21429
rect -2325 21398 -2317 21406
rect -2325 21378 -2320 21398
rect -2317 21390 -2309 21398
rect -2325 21374 -2317 21378
rect -2000 21374 -1992 21465
rect -1980 21448 -1932 21455
rect -1655 21444 -1647 21454
rect -1846 21430 -1680 21439
rect -1663 21438 -1655 21444
rect -1671 21398 -1663 21406
rect -1663 21390 -1655 21398
rect -1671 21374 -1663 21378
rect -1642 21374 -1637 21468
rect -1619 21374 -1614 21468
rect -1530 21374 -1526 21468
rect -1506 21374 -1502 21468
rect -1482 21374 -1478 21468
rect -1458 21374 -1454 21468
rect -1434 21374 -1430 21468
rect -1410 21374 -1406 21468
rect -1386 21374 -1382 21468
rect -1362 21374 -1358 21468
rect -1338 21374 -1334 21468
rect -1314 21374 -1310 21468
rect -1290 21374 -1286 21468
rect -1266 21374 -1262 21468
rect -1242 21374 -1238 21468
rect -1218 21374 -1214 21468
rect -1194 21374 -1190 21468
rect -1170 21374 -1166 21468
rect -1146 21374 -1142 21468
rect -1122 21374 -1118 21468
rect -1098 21374 -1094 21468
rect -1074 21374 -1070 21468
rect -1050 21374 -1046 21468
rect -1026 21374 -1022 21468
rect -1002 21374 -998 21468
rect -978 21374 -974 21468
rect -954 21374 -950 21468
rect -930 21374 -926 21468
rect -906 21374 -902 21468
rect -882 21374 -878 21468
rect -858 21374 -854 21468
rect -834 21374 -830 21468
rect -810 21374 -806 21468
rect -786 21374 -782 21468
rect -762 21374 -758 21468
rect -738 21374 -734 21468
rect -714 21374 -710 21468
rect -690 21374 -686 21468
rect -666 21374 -662 21468
rect -642 21374 -638 21468
rect -618 21374 -614 21468
rect -594 21374 -590 21468
rect -570 21374 -566 21468
rect -546 21374 -542 21468
rect -522 21374 -518 21468
rect -498 21374 -494 21468
rect -474 21374 -470 21468
rect -450 21374 -446 21468
rect -426 21374 -422 21468
rect -402 21374 -398 21468
rect -378 21374 -374 21468
rect -354 21374 -350 21468
rect -330 21374 -326 21468
rect -306 21374 -302 21468
rect -282 21374 -278 21468
rect -258 21374 -254 21468
rect -234 21374 -230 21468
rect -210 21374 -206 21468
rect -186 21374 -182 21468
rect -162 21374 -158 21468
rect -138 21374 -134 21468
rect -114 21374 -110 21468
rect -90 21374 -86 21468
rect -66 21374 -62 21468
rect -42 21374 -38 21468
rect -18 21374 -14 21468
rect 6 21374 10 21468
rect 30 21374 34 21468
rect 54 21374 58 21468
rect 78 21374 82 21468
rect 102 21374 106 21468
rect 126 21374 130 21468
rect 150 21374 154 21468
rect 174 21374 178 21468
rect 198 21374 202 21468
rect 222 21374 226 21468
rect 246 21374 250 21468
rect 270 21374 274 21468
rect 294 21374 298 21468
rect 318 21374 322 21468
rect 342 21374 346 21468
rect 366 21374 370 21468
rect 390 21374 394 21468
rect 414 21374 418 21468
rect 438 21374 442 21468
rect 462 21374 466 21468
rect 486 21374 490 21468
rect 510 21374 514 21468
rect 534 21374 538 21468
rect 547 21461 552 21468
rect 557 21447 562 21461
rect 558 21374 562 21447
rect 582 21419 586 21492
rect -2393 21372 579 21374
rect -2371 21326 -2366 21372
rect -2348 21326 -2343 21372
rect -2325 21364 -2317 21372
rect -2018 21371 -2004 21372
rect -2000 21371 -1992 21372
rect -2072 21370 -1928 21371
rect -2072 21364 -2053 21370
rect -2325 21348 -2320 21364
rect -2317 21362 -2309 21364
rect -2309 21350 -2301 21362
rect -2092 21355 -2062 21360
rect -2317 21348 -2309 21350
rect -2325 21336 -2317 21348
rect -2098 21342 -2096 21353
rect -2092 21342 -2084 21355
rect -2000 21354 -1992 21370
rect -1972 21364 -1928 21370
rect -1924 21364 -1918 21372
rect -1671 21364 -1663 21372
rect -1663 21362 -1655 21364
rect -2083 21344 -2062 21353
rect -2027 21352 -1992 21354
rect -2018 21344 -2002 21352
rect -2000 21344 -1992 21352
rect -2100 21337 -2096 21342
rect -2083 21337 -2053 21342
rect -2003 21340 -1990 21344
rect -1972 21342 -1964 21351
rect -1928 21350 -1924 21353
rect -1655 21350 -1647 21362
rect -1663 21348 -1655 21350
rect -2325 21326 -2320 21336
rect -2317 21334 -2309 21336
rect -2309 21326 -2301 21334
rect -2004 21330 -2003 21340
rect -2062 21326 -2012 21328
rect -2000 21326 -1992 21340
rect -1972 21337 -1924 21342
rect -1864 21337 -1796 21343
rect -1671 21336 -1663 21348
rect -1663 21334 -1655 21336
rect -1864 21326 -1796 21327
rect -1655 21326 -1647 21334
rect -1642 21326 -1637 21372
rect -1619 21326 -1614 21372
rect -1530 21326 -1526 21372
rect -1506 21327 -1502 21372
rect -1517 21326 -1483 21327
rect -2393 21324 -1483 21326
rect -2371 21278 -2366 21324
rect -2348 21278 -2343 21324
rect -2325 21320 -2320 21324
rect -2309 21322 -2301 21324
rect -2317 21320 -2309 21322
rect -2325 21308 -2317 21320
rect -2325 21278 -2320 21308
rect -2317 21306 -2309 21308
rect -2092 21294 -2062 21296
rect -2094 21290 -2062 21294
rect -2000 21278 -1992 21324
rect -1655 21322 -1647 21324
rect -1663 21320 -1655 21322
rect -1671 21308 -1663 21320
rect -1663 21306 -1655 21308
rect -1854 21294 -1806 21296
rect -1854 21290 -1680 21294
rect -1926 21278 -1892 21281
rect -1642 21278 -1637 21324
rect -1619 21278 -1614 21324
rect -1530 21278 -1526 21324
rect -1517 21317 -1512 21324
rect -1506 21317 -1502 21324
rect -1507 21303 -1502 21317
rect -1506 21278 -1502 21303
rect -1482 21278 -1478 21372
rect -1458 21278 -1454 21372
rect -1434 21278 -1430 21372
rect -1410 21278 -1406 21372
rect -1386 21278 -1382 21372
rect -1362 21278 -1358 21372
rect -1338 21278 -1334 21372
rect -1314 21278 -1310 21372
rect -1290 21278 -1286 21372
rect -1266 21278 -1262 21372
rect -1242 21278 -1238 21372
rect -1218 21278 -1214 21372
rect -1194 21278 -1190 21372
rect -1170 21278 -1166 21372
rect -1146 21278 -1142 21372
rect -1122 21278 -1118 21372
rect -1098 21278 -1094 21372
rect -1074 21278 -1070 21372
rect -1050 21278 -1046 21372
rect -1026 21278 -1022 21372
rect -1002 21278 -998 21372
rect -978 21278 -974 21372
rect -954 21278 -950 21372
rect -930 21278 -926 21372
rect -906 21278 -902 21372
rect -882 21278 -878 21372
rect -858 21278 -854 21372
rect -834 21278 -830 21372
rect -810 21278 -806 21372
rect -786 21278 -782 21372
rect -762 21278 -758 21372
rect -738 21278 -734 21372
rect -714 21278 -710 21372
rect -690 21278 -686 21372
rect -666 21278 -662 21372
rect -642 21278 -638 21372
rect -618 21278 -614 21372
rect -594 21278 -590 21372
rect -570 21278 -566 21372
rect -546 21278 -542 21372
rect -522 21278 -518 21372
rect -498 21278 -494 21372
rect -474 21278 -470 21372
rect -450 21278 -446 21372
rect -426 21278 -422 21372
rect -402 21278 -398 21372
rect -378 21278 -374 21372
rect -354 21278 -350 21372
rect -330 21278 -326 21372
rect -306 21278 -302 21372
rect -282 21278 -278 21372
rect -258 21278 -254 21372
rect -234 21278 -230 21372
rect -210 21278 -206 21372
rect -186 21278 -182 21372
rect -162 21278 -158 21372
rect -138 21278 -134 21372
rect -114 21278 -110 21372
rect -90 21278 -86 21372
rect -66 21278 -62 21372
rect -42 21278 -38 21372
rect -18 21278 -14 21372
rect 6 21278 10 21372
rect 30 21278 34 21372
rect 54 21278 58 21372
rect 78 21278 82 21372
rect 102 21278 106 21372
rect 126 21278 130 21372
rect 150 21278 154 21372
rect 174 21278 178 21372
rect 198 21278 202 21372
rect 222 21278 226 21372
rect 246 21278 250 21372
rect 270 21278 274 21372
rect 294 21278 298 21372
rect 318 21278 322 21372
rect 342 21278 346 21372
rect 366 21278 370 21372
rect 390 21278 394 21372
rect 414 21278 418 21372
rect 438 21278 442 21372
rect 462 21278 466 21372
rect 486 21278 490 21372
rect 510 21278 514 21372
rect 534 21278 538 21372
rect 558 21278 562 21372
rect 565 21371 579 21372
rect 582 21371 589 21419
rect 582 21278 586 21371
rect 606 21278 610 21492
rect 630 21278 634 21492
rect 654 21471 658 21492
rect 643 21470 677 21471
rect 678 21470 682 21492
rect 702 21470 706 21492
rect 726 21470 730 21492
rect 750 21470 754 21492
rect 774 21484 778 21492
rect 763 21470 797 21471
rect 643 21468 797 21470
rect 643 21461 648 21468
rect 654 21461 658 21468
rect 653 21447 658 21461
rect 643 21446 677 21447
rect 678 21446 682 21468
rect 702 21446 706 21468
rect 726 21446 730 21468
rect 750 21446 754 21468
rect 763 21461 768 21468
rect 773 21447 778 21461
rect 774 21446 778 21447
rect 798 21446 802 21492
rect 822 21471 826 21492
rect 811 21470 845 21471
rect 846 21470 850 21492
rect 870 21470 874 21492
rect 894 21470 898 21492
rect 918 21484 922 21492
rect 907 21470 941 21471
rect 811 21468 941 21470
rect 811 21461 816 21468
rect 822 21461 826 21468
rect 821 21447 826 21461
rect 846 21446 850 21468
rect 870 21446 874 21468
rect 894 21446 898 21468
rect 907 21461 912 21468
rect 917 21447 922 21461
rect 918 21446 922 21447
rect 942 21446 946 21492
rect 966 21446 970 21492
rect 990 21446 994 21492
rect 1014 21471 1018 21492
rect 1003 21470 1037 21471
rect 1038 21470 1042 21492
rect 1062 21484 1066 21492
rect 1051 21470 1085 21471
rect 1003 21468 1085 21470
rect 1003 21461 1008 21468
rect 1014 21461 1018 21468
rect 1013 21447 1018 21461
rect 1038 21446 1042 21468
rect 1051 21461 1056 21468
rect 1061 21447 1066 21461
rect 1062 21446 1066 21447
rect 1086 21446 1090 21492
rect 1110 21471 1114 21492
rect 1099 21470 1133 21471
rect 1134 21470 1138 21492
rect 1158 21484 1162 21492
rect 1147 21470 1181 21471
rect 1099 21468 1181 21470
rect 1099 21461 1104 21468
rect 1110 21461 1114 21468
rect 1109 21447 1114 21461
rect 1134 21446 1138 21468
rect 1147 21461 1152 21468
rect 1157 21447 1162 21461
rect 1158 21446 1162 21447
rect 1182 21446 1186 21492
rect 1206 21446 1210 21492
rect 1230 21446 1234 21492
rect 1254 21448 1258 21492
rect 1278 21484 1282 21492
rect 1278 21446 1282 21448
rect 1302 21446 1306 21492
rect 1326 21467 1330 21492
rect 1350 21491 1354 21492
rect 1326 21446 1333 21467
rect 1350 21446 1357 21491
rect 1374 21446 1378 21492
rect 1398 21446 1402 21492
rect 1411 21461 1416 21471
rect 1422 21461 1426 21492
rect 1421 21447 1426 21461
rect 1446 21446 1450 21492
rect 1470 21484 1474 21492
rect 1459 21461 1464 21471
rect 1469 21447 1474 21461
rect 1470 21446 1474 21447
rect 1494 21446 1498 21492
rect 1518 21446 1522 21492
rect 1542 21446 1546 21492
rect 1555 21461 1560 21471
rect 1566 21461 1570 21492
rect 1565 21447 1570 21461
rect 1590 21446 1594 21492
rect 1614 21446 1618 21492
rect 1638 21446 1642 21492
rect 1662 21446 1666 21492
rect 1686 21446 1690 21492
rect 1710 21446 1714 21492
rect 1734 21484 1738 21492
rect 1723 21461 1728 21471
rect 1733 21447 1738 21461
rect 1734 21446 1738 21447
rect 1758 21446 1762 21492
rect 1782 21448 1786 21492
rect 1806 21484 1810 21492
rect 1806 21446 1810 21448
rect 1830 21446 1834 21492
rect 1843 21461 1848 21471
rect 1854 21461 1858 21492
rect 1853 21447 1858 21461
rect 1878 21446 1882 21492
rect 1902 21446 1906 21492
rect 1926 21446 1930 21492
rect 1950 21446 1954 21492
rect 1974 21484 1978 21492
rect 1963 21461 1968 21471
rect 1973 21447 1978 21461
rect 1974 21446 1978 21447
rect 1998 21446 2002 21492
rect 2022 21446 2026 21492
rect 2046 21446 2050 21492
rect 2059 21461 2064 21471
rect 2070 21461 2074 21492
rect 2069 21447 2074 21461
rect 2094 21446 2098 21492
rect 2118 21484 2122 21492
rect 2107 21461 2112 21471
rect 2117 21447 2122 21461
rect 2118 21446 2122 21447
rect 2142 21446 2146 21492
rect 2166 21446 2170 21492
rect 2179 21461 2184 21471
rect 2190 21461 2194 21492
rect 2189 21447 2194 21461
rect 2214 21446 2218 21492
rect 2238 21446 2242 21492
rect 2262 21446 2266 21492
rect 2286 21446 2290 21492
rect 2310 21484 2314 21492
rect 2299 21461 2304 21471
rect 2309 21447 2314 21461
rect 2310 21446 2314 21447
rect 2334 21446 2338 21492
rect 2341 21491 2355 21492
rect 2358 21467 2365 21515
rect 2358 21446 2362 21467
rect 2382 21446 2386 21516
rect 2389 21515 2403 21516
rect 2406 21494 2413 21539
rect 2430 21494 2434 21564
rect 2454 21494 2458 21564
rect 2478 21494 2482 21564
rect 2502 21494 2506 21564
rect 2526 21495 2530 21564
rect 2515 21494 2549 21495
rect 2389 21492 2549 21494
rect 2389 21491 2403 21492
rect 2406 21491 2413 21492
rect 2406 21446 2410 21491
rect 2430 21446 2434 21492
rect 2454 21446 2458 21492
rect 2478 21446 2482 21492
rect 2502 21471 2506 21492
rect 2515 21485 2520 21492
rect 2526 21485 2530 21492
rect 2525 21471 2530 21485
rect 2550 21472 2554 21564
rect 2491 21470 2525 21471
rect 2526 21470 2530 21471
rect 2539 21470 2573 21471
rect 2491 21468 2573 21470
rect 2491 21461 2496 21468
rect 2502 21461 2506 21468
rect 2501 21447 2506 21461
rect 2491 21446 2525 21447
rect 643 21444 1323 21446
rect 643 21437 648 21444
rect 653 21423 658 21437
rect 654 21278 658 21423
rect 678 21395 682 21444
rect 678 21374 685 21395
rect 702 21374 706 21444
rect 726 21374 730 21444
rect 750 21374 754 21444
rect 774 21374 778 21444
rect 798 21408 802 21444
rect 812 21412 816 21422
rect 661 21372 795 21374
rect 661 21371 675 21372
rect 678 21350 685 21372
rect 702 21350 706 21372
rect 726 21350 730 21372
rect 750 21350 754 21372
rect 774 21350 778 21372
rect 781 21371 795 21372
rect 798 21371 805 21395
rect 798 21350 802 21371
rect 822 21350 826 21412
rect 846 21395 850 21444
rect 846 21374 853 21395
rect 870 21374 874 21444
rect 894 21374 898 21444
rect 918 21374 922 21444
rect 942 21408 946 21444
rect 829 21372 939 21374
rect 829 21371 843 21372
rect 846 21371 853 21372
rect 870 21350 874 21372
rect 894 21350 898 21372
rect 918 21350 922 21372
rect 925 21371 939 21372
rect 942 21371 949 21395
rect 942 21350 946 21371
rect 966 21350 970 21444
rect 990 21350 994 21444
rect 1004 21412 1008 21422
rect 1014 21350 1018 21412
rect 1038 21395 1042 21444
rect 1038 21374 1045 21395
rect 1062 21374 1066 21444
rect 1086 21408 1090 21444
rect 1100 21412 1104 21422
rect 1021 21372 1083 21374
rect 1021 21371 1035 21372
rect 1038 21371 1045 21372
rect 1062 21350 1066 21372
rect 1069 21371 1083 21372
rect 1086 21371 1093 21395
rect 1086 21350 1090 21371
rect 1110 21350 1114 21412
rect 1134 21395 1138 21444
rect 1134 21374 1141 21395
rect 1158 21374 1162 21444
rect 1182 21408 1186 21444
rect 1117 21372 1179 21374
rect 1117 21371 1131 21372
rect 1134 21371 1141 21372
rect 1158 21350 1162 21372
rect 1165 21371 1179 21372
rect 1182 21371 1189 21395
rect 1182 21350 1186 21371
rect 1206 21350 1210 21444
rect 1230 21350 1234 21444
rect 1244 21412 1248 21422
rect 1254 21350 1258 21412
rect 1278 21382 1282 21444
rect 1302 21408 1306 21444
rect 1309 21443 1323 21444
rect 1326 21444 2525 21446
rect 1326 21443 1347 21444
rect 1350 21443 1357 21444
rect 1326 21422 1333 21443
rect 1350 21422 1354 21443
rect 1374 21422 1378 21444
rect 1398 21422 1402 21444
rect 1446 21422 1450 21444
rect 1470 21422 1474 21444
rect 1494 21422 1498 21444
rect 1518 21422 1522 21444
rect 1542 21422 1546 21444
rect 1590 21422 1594 21444
rect 1614 21422 1618 21444
rect 1638 21422 1642 21444
rect 1662 21422 1666 21444
rect 1686 21422 1690 21444
rect 1710 21422 1714 21444
rect 1734 21422 1738 21444
rect 1758 21422 1762 21444
rect 1806 21422 1810 21444
rect 1830 21422 1834 21444
rect 1878 21422 1882 21444
rect 1902 21422 1906 21444
rect 1926 21422 1930 21444
rect 1950 21422 1954 21444
rect 1974 21422 1978 21444
rect 1998 21422 2002 21444
rect 2022 21422 2026 21444
rect 2046 21422 2050 21444
rect 2094 21422 2098 21444
rect 2118 21422 2122 21444
rect 2142 21422 2146 21444
rect 2166 21422 2170 21444
rect 2214 21422 2218 21444
rect 2238 21422 2242 21444
rect 2262 21422 2266 21444
rect 2286 21422 2290 21444
rect 2310 21422 2314 21444
rect 2334 21422 2338 21444
rect 2358 21422 2362 21444
rect 2382 21422 2386 21444
rect 2406 21422 2410 21444
rect 2430 21423 2434 21444
rect 2419 21422 2453 21423
rect 1309 21420 2453 21422
rect 1309 21419 1323 21420
rect 1326 21419 1333 21420
rect 1302 21350 1306 21392
rect 1326 21350 1330 21419
rect 1350 21350 1354 21420
rect 1374 21350 1378 21420
rect 1398 21350 1402 21420
rect 1412 21412 1416 21420
rect 1422 21350 1426 21412
rect 1446 21395 1450 21420
rect 1446 21374 1453 21395
rect 1470 21374 1474 21420
rect 1494 21408 1498 21420
rect 1429 21372 1491 21374
rect 1429 21371 1443 21372
rect 1446 21371 1453 21372
rect 1470 21350 1474 21372
rect 1477 21371 1491 21372
rect 1494 21371 1501 21395
rect 1494 21350 1498 21371
rect 1518 21350 1522 21420
rect 1542 21350 1546 21420
rect 1556 21412 1560 21420
rect 1566 21350 1570 21412
rect 1590 21395 1594 21420
rect 1590 21374 1597 21395
rect 1614 21374 1618 21420
rect 1638 21374 1642 21420
rect 1662 21374 1666 21420
rect 1686 21374 1690 21420
rect 1710 21374 1714 21420
rect 1734 21374 1738 21420
rect 1758 21408 1762 21420
rect 1772 21412 1776 21420
rect 1573 21372 1755 21374
rect 1573 21371 1587 21372
rect 1590 21371 1597 21372
rect 1614 21350 1618 21372
rect 1638 21350 1642 21372
rect 1662 21350 1666 21372
rect 1686 21350 1690 21372
rect 1710 21350 1714 21372
rect 1734 21350 1738 21372
rect 1741 21371 1755 21372
rect 1758 21371 1765 21395
rect 1758 21350 1762 21371
rect 1782 21350 1786 21412
rect 1806 21382 1810 21420
rect 1830 21408 1834 21420
rect 1844 21412 1848 21420
rect 1830 21350 1834 21392
rect 1854 21350 1858 21412
rect 1878 21395 1882 21420
rect 1878 21374 1885 21395
rect 1902 21374 1906 21420
rect 1926 21374 1930 21420
rect 1950 21374 1954 21420
rect 1974 21374 1978 21420
rect 1998 21408 2002 21420
rect 1861 21372 1995 21374
rect 1861 21371 1875 21372
rect 1878 21371 1885 21372
rect 1902 21350 1906 21372
rect 1926 21350 1930 21372
rect 1950 21350 1954 21372
rect 1974 21350 1978 21372
rect 1981 21371 1995 21372
rect 1998 21371 2005 21395
rect 1998 21350 2002 21371
rect 2022 21350 2026 21420
rect 2046 21350 2050 21420
rect 2060 21412 2064 21420
rect 2070 21350 2074 21412
rect 2094 21395 2098 21420
rect 2094 21374 2101 21395
rect 2118 21374 2122 21420
rect 2142 21408 2146 21420
rect 2077 21372 2139 21374
rect 2077 21371 2091 21372
rect 2094 21371 2101 21372
rect 2118 21350 2122 21372
rect 2125 21371 2139 21372
rect 2142 21371 2149 21395
rect 2142 21350 2146 21371
rect 2166 21350 2170 21420
rect 2180 21412 2184 21420
rect 2190 21350 2194 21412
rect 2214 21395 2218 21420
rect 2214 21374 2221 21395
rect 2238 21374 2242 21420
rect 2262 21374 2266 21420
rect 2286 21374 2290 21420
rect 2310 21374 2314 21420
rect 2334 21408 2338 21420
rect 2197 21372 2331 21374
rect 2197 21371 2211 21372
rect 2214 21371 2221 21372
rect 2238 21350 2242 21372
rect 2262 21350 2266 21372
rect 2286 21350 2290 21372
rect 2310 21350 2314 21372
rect 2317 21371 2331 21372
rect 2334 21371 2341 21395
rect 2334 21350 2338 21371
rect 2358 21350 2362 21420
rect 2382 21350 2386 21420
rect 2406 21350 2410 21420
rect 2419 21413 2424 21420
rect 2430 21413 2434 21420
rect 2429 21399 2434 21413
rect 2419 21398 2453 21399
rect 2454 21398 2458 21444
rect 2478 21398 2482 21444
rect 2491 21437 2496 21444
rect 2501 21423 2506 21437
rect 2526 21434 2530 21468
rect 2539 21461 2544 21468
rect 2549 21447 2554 21461
rect 2492 21412 2496 21422
rect 2516 21412 2520 21422
rect 2550 21419 2554 21447
rect 2502 21398 2506 21412
rect 2526 21398 2530 21412
rect 2419 21396 2547 21398
rect 2419 21389 2424 21396
rect 2429 21375 2434 21389
rect 2430 21350 2434 21375
rect 2454 21350 2458 21396
rect 2478 21350 2482 21396
rect 2502 21350 2506 21396
rect 2526 21395 2530 21396
rect 2533 21395 2547 21396
rect 2550 21395 2557 21419
rect 2574 21396 2578 21564
rect 2526 21374 2533 21395
rect 2550 21374 2554 21395
rect 2509 21372 2571 21374
rect 2509 21371 2523 21372
rect 2526 21358 2533 21372
rect 661 21348 2523 21350
rect 2550 21348 2554 21372
rect 2557 21371 2571 21372
rect 2574 21371 2581 21395
rect 661 21347 675 21348
rect 678 21347 685 21348
rect 678 21278 682 21347
rect 702 21278 706 21348
rect 726 21278 730 21348
rect 750 21278 754 21348
rect 774 21278 778 21348
rect 798 21278 802 21348
rect 822 21278 826 21348
rect 846 21278 850 21346
rect 870 21278 874 21348
rect 894 21278 898 21348
rect 918 21278 922 21348
rect 942 21278 946 21348
rect 966 21278 970 21348
rect 990 21278 994 21348
rect 1014 21278 1018 21348
rect 1038 21278 1042 21346
rect 1062 21278 1066 21348
rect 1086 21278 1090 21348
rect 1110 21278 1114 21348
rect 1134 21278 1138 21346
rect 1158 21278 1162 21348
rect 1182 21278 1186 21348
rect 1206 21278 1210 21348
rect 1230 21278 1234 21348
rect 1254 21278 1258 21348
rect 1278 21278 1282 21346
rect 1302 21278 1306 21348
rect 1326 21278 1330 21348
rect 1350 21278 1354 21348
rect 1374 21278 1378 21348
rect 1398 21278 1402 21348
rect 1422 21278 1426 21348
rect 1446 21278 1450 21346
rect 1470 21278 1474 21348
rect 1494 21278 1498 21348
rect 1518 21278 1522 21348
rect 1542 21278 1546 21348
rect 1566 21278 1570 21348
rect 1590 21278 1594 21346
rect 1614 21278 1618 21348
rect 1638 21278 1642 21348
rect 1662 21278 1666 21348
rect 1686 21278 1690 21348
rect 1710 21278 1714 21348
rect 1734 21278 1738 21348
rect 1758 21278 1762 21348
rect 1782 21278 1786 21348
rect 1806 21278 1810 21346
rect 1830 21278 1834 21348
rect 1854 21278 1858 21348
rect 1878 21278 1882 21346
rect 1902 21278 1906 21348
rect 1926 21278 1930 21348
rect 1950 21278 1954 21348
rect 1974 21278 1978 21348
rect 1998 21278 2002 21348
rect 2022 21278 2026 21348
rect 2046 21278 2050 21348
rect 2070 21278 2074 21348
rect 2094 21278 2098 21346
rect 2118 21278 2122 21348
rect 2142 21278 2146 21348
rect 2166 21278 2170 21348
rect 2190 21278 2194 21348
rect 2214 21278 2218 21346
rect 2238 21278 2242 21348
rect 2262 21278 2266 21348
rect 2286 21278 2290 21348
rect 2310 21278 2314 21348
rect 2334 21278 2338 21348
rect 2358 21278 2362 21348
rect 2382 21278 2386 21348
rect 2406 21278 2410 21348
rect 2430 21278 2434 21348
rect 2454 21347 2458 21348
rect 2454 21299 2461 21347
rect 2454 21278 2458 21299
rect 2478 21278 2482 21348
rect 2502 21278 2506 21348
rect 2509 21347 2523 21348
rect 2526 21347 2533 21348
rect 2526 21278 2530 21346
rect 2550 21278 2554 21346
rect 2574 21278 2578 21371
rect 2598 21278 2602 21564
rect 2622 21471 2626 21564
rect 2611 21470 2645 21471
rect 2646 21470 2650 21564
rect 2670 21495 2674 21564
rect 2659 21494 2693 21495
rect 2694 21494 2698 21564
rect 2718 21494 2722 21564
rect 2742 21494 2746 21564
rect 2766 21494 2770 21564
rect 2790 21494 2794 21564
rect 2814 21494 2818 21564
rect 2838 21494 2842 21564
rect 2862 21542 2869 21563
rect 2886 21542 2890 21564
rect 2910 21542 2914 21564
rect 2934 21542 2938 21564
rect 2958 21542 2962 21564
rect 2982 21563 2986 21564
rect 2845 21540 2979 21542
rect 2845 21539 2859 21540
rect 2862 21539 2869 21540
rect 2862 21494 2866 21539
rect 2886 21494 2890 21540
rect 2910 21494 2914 21540
rect 2934 21494 2938 21540
rect 2958 21494 2962 21540
rect 2965 21539 2979 21540
rect 2982 21518 2989 21563
rect 3006 21518 3010 21564
rect 3030 21518 3034 21564
rect 3054 21518 3058 21564
rect 3078 21542 3085 21563
rect 3102 21542 3106 21564
rect 3126 21542 3130 21564
rect 3150 21542 3154 21564
rect 3174 21542 3178 21564
rect 3198 21542 3202 21564
rect 3222 21542 3226 21564
rect 3283 21557 3288 21564
rect 3301 21563 3315 21564
rect 3349 21563 3363 21564
rect 3293 21543 3298 21557
rect 3307 21553 3315 21557
rect 3355 21553 3363 21557
rect 3301 21543 3307 21553
rect 3349 21543 3355 21553
rect 3283 21542 3317 21543
rect 3061 21540 3317 21542
rect 3331 21542 3365 21543
rect 3366 21542 3373 21564
rect 3379 21557 3384 21564
rect 3397 21563 3411 21564
rect 3829 21563 3843 21564
rect 3389 21543 3394 21557
rect 3403 21553 3411 21557
rect 3835 21553 3843 21557
rect 3397 21543 3403 21553
rect 3829 21543 3835 21553
rect 3379 21542 3413 21543
rect 3331 21540 3413 21542
rect 3811 21542 3845 21543
rect 3846 21542 3853 21564
rect 3859 21557 3864 21564
rect 3877 21563 3891 21564
rect 4549 21563 4563 21564
rect 3869 21543 3874 21557
rect 3883 21553 3891 21557
rect 4555 21553 4563 21557
rect 3877 21543 3883 21553
rect 4549 21543 4555 21553
rect 3859 21542 3893 21543
rect 3811 21540 3893 21542
rect 4531 21542 4565 21543
rect 4566 21542 4573 21564
rect 4579 21557 4584 21564
rect 4597 21563 4611 21564
rect 4789 21563 4803 21564
rect 4589 21543 4594 21557
rect 4603 21553 4611 21557
rect 4795 21553 4803 21557
rect 4597 21543 4603 21553
rect 4789 21543 4795 21553
rect 4579 21542 4613 21543
rect 4531 21540 4613 21542
rect 4771 21542 4805 21543
rect 4806 21542 4813 21564
rect 4819 21557 4824 21564
rect 4837 21563 4851 21564
rect 6589 21563 6603 21564
rect 4829 21543 4834 21557
rect 4843 21553 4851 21557
rect 6595 21553 6603 21557
rect 4837 21543 4843 21553
rect 6589 21543 6595 21553
rect 4819 21542 4853 21543
rect 4771 21540 4853 21542
rect 6571 21542 6605 21543
rect 6606 21542 6613 21564
rect 6654 21542 6658 21564
rect 6702 21542 6706 21564
rect 6726 21542 6730 21564
rect 6750 21542 6754 21564
rect 6774 21542 6778 21564
rect 6798 21542 6802 21564
rect 6822 21542 6826 21564
rect 6846 21542 6850 21564
rect 6870 21542 6874 21564
rect 6894 21542 6898 21564
rect 6918 21542 6922 21564
rect 6942 21542 6946 21564
rect 6966 21542 6970 21564
rect 6990 21542 6994 21564
rect 7038 21542 7042 21564
rect 7099 21557 7104 21564
rect 7117 21563 7131 21564
rect 7501 21563 7515 21564
rect 7109 21543 7114 21557
rect 7123 21553 7131 21557
rect 7507 21553 7515 21557
rect 7117 21543 7123 21553
rect 7501 21543 7507 21553
rect 7099 21542 7133 21543
rect 6571 21540 7133 21542
rect 7483 21542 7517 21543
rect 7518 21542 7525 21564
rect 7531 21557 7536 21564
rect 7549 21563 7563 21564
rect 8245 21563 8259 21564
rect 7541 21543 7546 21557
rect 7555 21553 7563 21557
rect 8251 21553 8259 21557
rect 7549 21543 7555 21553
rect 8245 21543 8251 21553
rect 7531 21542 7565 21543
rect 7483 21540 7565 21542
rect 8227 21542 8261 21543
rect 8262 21542 8269 21564
rect 8275 21557 8280 21564
rect 8293 21563 8307 21564
rect 14533 21563 14547 21564
rect 14581 21563 14595 21564
rect 14749 21563 14763 21564
rect 8285 21543 8290 21557
rect 8299 21553 8307 21557
rect 8293 21543 8299 21553
rect 14549 21543 14554 21557
rect 14755 21553 14763 21557
rect 14749 21543 14755 21553
rect 8275 21542 8309 21543
rect 8227 21540 8309 21542
rect 14491 21540 14525 21543
rect 3061 21539 3075 21540
rect 3078 21539 3085 21540
rect 3078 21518 3082 21539
rect 3102 21518 3106 21540
rect 3126 21518 3130 21540
rect 3150 21518 3154 21540
rect 3174 21518 3178 21540
rect 3198 21518 3202 21540
rect 3222 21518 3226 21540
rect 3283 21533 3288 21540
rect 3301 21539 3315 21540
rect 3349 21539 3363 21540
rect 3293 21519 3298 21533
rect 3307 21529 3315 21533
rect 3355 21529 3363 21533
rect 3301 21519 3307 21529
rect 3349 21519 3355 21529
rect 3283 21518 3317 21519
rect 2965 21516 3317 21518
rect 3331 21518 3365 21519
rect 3366 21518 3373 21540
rect 3379 21533 3384 21540
rect 3397 21539 3411 21540
rect 3829 21539 3843 21540
rect 3389 21519 3394 21533
rect 3403 21529 3411 21533
rect 3835 21529 3843 21533
rect 3397 21519 3403 21529
rect 3829 21519 3835 21529
rect 3379 21518 3413 21519
rect 3331 21516 3413 21518
rect 3811 21518 3845 21519
rect 3846 21518 3853 21540
rect 3859 21533 3864 21540
rect 3877 21539 3891 21540
rect 4549 21539 4563 21540
rect 3869 21519 3874 21533
rect 3883 21529 3891 21533
rect 4555 21529 4563 21533
rect 3877 21519 3883 21529
rect 4549 21519 4555 21529
rect 3859 21518 3893 21519
rect 3811 21516 3893 21518
rect 4531 21518 4565 21519
rect 4566 21518 4573 21540
rect 4579 21533 4584 21540
rect 4597 21539 4611 21540
rect 4789 21539 4803 21540
rect 4589 21519 4594 21533
rect 4603 21529 4611 21533
rect 4795 21529 4803 21533
rect 4597 21519 4603 21529
rect 4789 21519 4795 21529
rect 4579 21518 4613 21519
rect 4531 21516 4613 21518
rect 4771 21518 4805 21519
rect 4806 21518 4813 21540
rect 4819 21533 4824 21540
rect 4837 21539 4851 21540
rect 6589 21539 6603 21540
rect 4829 21519 4834 21533
rect 4843 21529 4851 21533
rect 6595 21529 6603 21533
rect 4837 21519 4843 21529
rect 6589 21519 6595 21529
rect 4819 21518 4853 21519
rect 4771 21516 4853 21518
rect 6571 21518 6605 21519
rect 6606 21518 6613 21540
rect 6654 21518 6658 21540
rect 6571 21516 6675 21518
rect 6702 21516 6706 21540
rect 2965 21515 2979 21516
rect 2982 21515 2989 21516
rect 2982 21494 2986 21515
rect 3006 21494 3010 21516
rect 3030 21494 3034 21516
rect 3054 21494 3058 21516
rect 3078 21494 3082 21516
rect 3102 21494 3106 21516
rect 3126 21494 3130 21516
rect 3150 21494 3154 21516
rect 3174 21494 3178 21516
rect 3198 21494 3202 21516
rect 3222 21494 3226 21516
rect 3283 21509 3288 21516
rect 3301 21515 3315 21516
rect 3349 21515 3363 21516
rect 3293 21495 3298 21509
rect 3307 21505 3315 21509
rect 3355 21505 3363 21509
rect 3301 21495 3307 21505
rect 3349 21495 3355 21505
rect 3235 21494 3269 21495
rect 2659 21492 3269 21494
rect 2659 21485 2664 21492
rect 2670 21485 2674 21492
rect 2669 21471 2674 21485
rect 2659 21470 2693 21471
rect 2611 21468 2693 21470
rect 2611 21461 2616 21468
rect 2622 21461 2626 21468
rect 2621 21447 2626 21461
rect 2612 21434 2616 21444
rect 2622 21278 2626 21434
rect 2646 21395 2650 21468
rect 2659 21461 2664 21468
rect 2669 21447 2674 21461
rect 2646 21374 2653 21395
rect 2670 21374 2674 21447
rect 2694 21419 2698 21492
rect 2694 21398 2701 21419
rect 2718 21398 2722 21492
rect 2742 21398 2746 21492
rect 2766 21471 2770 21492
rect 2755 21470 2789 21471
rect 2790 21470 2794 21492
rect 2814 21484 2818 21492
rect 2803 21470 2837 21471
rect 2755 21468 2837 21470
rect 2755 21461 2760 21468
rect 2766 21461 2770 21468
rect 2765 21447 2770 21461
rect 2755 21446 2789 21447
rect 2790 21446 2794 21468
rect 2803 21461 2808 21468
rect 2813 21447 2818 21461
rect 2814 21446 2818 21447
rect 2838 21446 2842 21492
rect 2862 21446 2866 21492
rect 2886 21446 2890 21492
rect 2910 21446 2914 21492
rect 2934 21471 2938 21492
rect 2923 21470 2957 21471
rect 2958 21470 2962 21492
rect 2982 21484 2986 21492
rect 2971 21470 3005 21471
rect 2923 21468 3005 21470
rect 2923 21461 2928 21468
rect 2934 21461 2938 21468
rect 2933 21447 2938 21461
rect 2958 21446 2962 21468
rect 2971 21461 2976 21468
rect 2981 21447 2986 21461
rect 2982 21446 2986 21447
rect 3006 21446 3010 21492
rect 3030 21471 3034 21492
rect 3019 21470 3053 21471
rect 3054 21470 3058 21492
rect 3078 21484 3082 21492
rect 3102 21471 3106 21492
rect 3067 21470 3125 21471
rect 3126 21470 3130 21492
rect 3150 21484 3154 21492
rect 3139 21470 3173 21471
rect 3019 21468 3173 21470
rect 3019 21461 3024 21468
rect 3030 21461 3034 21468
rect 3029 21447 3034 21461
rect 3054 21446 3058 21468
rect 3067 21461 3072 21468
rect 3091 21461 3096 21468
rect 3102 21461 3106 21468
rect 3077 21447 3082 21461
rect 3101 21447 3106 21461
rect 3078 21446 3082 21447
rect 3126 21446 3130 21468
rect 3139 21461 3144 21468
rect 3149 21447 3154 21461
rect 3150 21446 3154 21447
rect 3174 21446 3178 21492
rect 3198 21446 3202 21492
rect 3222 21446 3226 21492
rect 3235 21485 3240 21492
rect 3245 21471 3250 21485
rect 3246 21447 3250 21471
rect 3301 21467 3314 21468
rect 3235 21446 3269 21447
rect 2755 21444 3269 21446
rect 2755 21437 2760 21444
rect 2765 21423 2770 21437
rect 2766 21398 2770 21423
rect 2790 21398 2794 21444
rect 2814 21398 2818 21444
rect 2838 21408 2842 21444
rect 2862 21398 2866 21444
rect 2886 21398 2890 21444
rect 2910 21398 2914 21444
rect 2924 21412 2928 21422
rect 2934 21398 2938 21412
rect 2958 21398 2962 21444
rect 2982 21398 2986 21444
rect 3006 21408 3010 21444
rect 3020 21412 3024 21422
rect 3030 21398 3034 21412
rect 3054 21398 3058 21444
rect 3078 21398 3082 21444
rect 3092 21412 3096 21422
rect 3102 21408 3106 21412
rect 3126 21398 3130 21444
rect 3150 21398 3154 21444
rect 3174 21408 3178 21444
rect 3198 21398 3202 21444
rect 3222 21398 3226 21444
rect 3235 21437 3240 21444
rect 3246 21437 3250 21444
rect 3245 21423 3250 21437
rect 3294 21424 3298 21448
rect 3304 21443 3315 21444
rect 3235 21422 3269 21423
rect 3366 21422 3373 21516
rect 3379 21509 3384 21516
rect 3397 21515 3411 21516
rect 3829 21515 3843 21516
rect 3389 21495 3394 21509
rect 3403 21505 3411 21509
rect 3835 21505 3843 21509
rect 3397 21495 3403 21505
rect 3829 21495 3835 21505
rect 3379 21422 3413 21423
rect 3235 21420 3315 21422
rect 3349 21420 3413 21422
rect 3811 21422 3845 21423
rect 3846 21422 3853 21516
rect 3859 21509 3864 21516
rect 3877 21515 3891 21516
rect 4549 21515 4563 21516
rect 3869 21495 3874 21509
rect 3883 21505 3891 21509
rect 4555 21505 4563 21509
rect 3877 21495 3883 21505
rect 4549 21495 4555 21505
rect 3859 21422 3893 21423
rect 3811 21420 3893 21422
rect 4531 21422 4565 21423
rect 4566 21422 4573 21516
rect 4579 21509 4584 21516
rect 4597 21515 4611 21516
rect 4789 21515 4803 21516
rect 4589 21495 4594 21509
rect 4603 21505 4611 21509
rect 4795 21505 4803 21509
rect 4597 21495 4603 21505
rect 4789 21495 4795 21505
rect 4579 21422 4613 21423
rect 4531 21420 4613 21422
rect 4771 21422 4805 21423
rect 4806 21422 4813 21516
rect 4819 21509 4824 21516
rect 4837 21515 4851 21516
rect 6589 21515 6603 21516
rect 4829 21495 4834 21509
rect 4843 21505 4851 21509
rect 6595 21505 6603 21509
rect 4837 21495 4843 21505
rect 6589 21495 6595 21505
rect 4819 21422 4853 21423
rect 4771 21420 4853 21422
rect 6571 21422 6605 21423
rect 6606 21422 6613 21516
rect 6654 21515 6658 21516
rect 6661 21515 6675 21516
rect 6654 21491 6661 21515
rect 6702 21491 6709 21515
rect 6726 21422 6730 21540
rect 6750 21422 6754 21540
rect 6774 21422 6778 21540
rect 6798 21422 6802 21540
rect 6822 21422 6826 21540
rect 6846 21422 6850 21540
rect 6870 21422 6874 21540
rect 6894 21422 6898 21540
rect 6918 21422 6922 21540
rect 6942 21422 6946 21540
rect 6966 21422 6970 21540
rect 6990 21422 6994 21540
rect 7014 21518 7021 21539
rect 7038 21518 7042 21540
rect 7099 21533 7104 21540
rect 7117 21539 7131 21540
rect 7501 21539 7515 21540
rect 7109 21519 7114 21533
rect 7123 21529 7131 21533
rect 7507 21529 7515 21533
rect 7117 21519 7123 21529
rect 7501 21519 7507 21529
rect 7099 21518 7133 21519
rect 6997 21516 7133 21518
rect 7483 21518 7517 21519
rect 7518 21518 7525 21540
rect 7531 21533 7536 21540
rect 7549 21539 7563 21540
rect 8245 21539 8259 21540
rect 7541 21519 7546 21533
rect 7555 21529 7563 21533
rect 8251 21529 8259 21533
rect 7549 21519 7555 21529
rect 8245 21519 8251 21529
rect 7531 21518 7565 21519
rect 7483 21516 7565 21518
rect 8227 21518 8261 21519
rect 8262 21518 8269 21540
rect 8275 21533 8280 21540
rect 8293 21539 8307 21540
rect 8285 21519 8290 21533
rect 8299 21529 8307 21533
rect 14515 21529 14523 21533
rect 8293 21519 8299 21529
rect 14509 21519 14515 21529
rect 8275 21518 8309 21519
rect 8227 21516 8309 21518
rect 14491 21518 14525 21519
rect 14526 21518 14533 21539
rect 14539 21533 14544 21543
rect 14558 21540 14573 21543
rect 14731 21542 14765 21543
rect 14766 21542 14773 21564
rect 14779 21557 14784 21564
rect 14797 21563 14811 21564
rect 14989 21563 15003 21564
rect 14789 21543 14794 21557
rect 14803 21553 14811 21557
rect 14995 21553 15003 21557
rect 14797 21543 14803 21553
rect 14989 21543 14995 21553
rect 14779 21542 14813 21543
rect 14731 21540 14813 21542
rect 14971 21542 15005 21543
rect 15006 21542 15013 21564
rect 15019 21557 15024 21564
rect 15037 21563 15051 21564
rect 15229 21563 15243 21564
rect 15029 21543 15034 21557
rect 15043 21553 15051 21557
rect 15235 21553 15243 21557
rect 15037 21543 15043 21553
rect 15229 21543 15235 21553
rect 15019 21542 15053 21543
rect 14971 21540 15053 21542
rect 15211 21542 15245 21543
rect 15246 21542 15253 21564
rect 15259 21557 15264 21564
rect 15277 21563 15291 21564
rect 15709 21563 15723 21564
rect 15269 21543 15274 21557
rect 15283 21553 15291 21557
rect 15715 21553 15723 21557
rect 15277 21543 15283 21553
rect 15709 21543 15715 21553
rect 15259 21542 15293 21543
rect 15211 21540 15293 21542
rect 15691 21542 15725 21543
rect 15726 21542 15733 21564
rect 15739 21557 15744 21564
rect 15757 21563 15771 21564
rect 15949 21563 15963 21564
rect 15749 21543 15754 21557
rect 15763 21553 15771 21557
rect 15955 21553 15963 21557
rect 15757 21543 15763 21553
rect 15949 21543 15955 21553
rect 15739 21542 15773 21543
rect 15691 21540 15773 21542
rect 15931 21542 15965 21543
rect 15966 21542 15973 21564
rect 15979 21557 15984 21564
rect 15997 21563 16011 21564
rect 16189 21563 16203 21564
rect 15989 21543 15994 21557
rect 16003 21553 16011 21557
rect 16195 21553 16203 21557
rect 15997 21543 16003 21553
rect 16189 21543 16195 21553
rect 15979 21542 16013 21543
rect 15931 21540 16013 21542
rect 16171 21542 16205 21543
rect 16206 21542 16213 21564
rect 16219 21557 16224 21564
rect 16237 21563 16251 21564
rect 16381 21563 16395 21564
rect 16229 21543 16234 21557
rect 16243 21553 16251 21557
rect 16387 21553 16395 21557
rect 16237 21543 16243 21553
rect 16381 21543 16387 21553
rect 16219 21542 16253 21543
rect 16171 21540 16253 21542
rect 16363 21542 16397 21543
rect 16398 21542 16405 21564
rect 16411 21557 16416 21564
rect 16429 21563 16443 21564
rect 16421 21543 16426 21557
rect 16435 21553 16443 21557
rect 25795 21553 25803 21557
rect 16429 21543 16435 21553
rect 25789 21543 25795 21553
rect 16411 21542 16445 21543
rect 16363 21540 16445 21542
rect 25771 21542 25805 21543
rect 25806 21542 25813 21563
rect 25819 21557 25824 21567
rect 25838 21564 25853 21567
rect 25939 21564 25973 21567
rect 25987 21564 26006 21567
rect 25829 21543 25834 21557
rect 25843 21553 25851 21557
rect 25837 21543 25843 21553
rect 25997 21543 26002 21557
rect 25819 21542 25853 21543
rect 25771 21540 25853 21542
rect 25939 21540 25973 21543
rect 14749 21539 14763 21540
rect 14549 21519 14554 21533
rect 14563 21529 14571 21533
rect 14755 21529 14763 21533
rect 14557 21519 14563 21529
rect 14749 21519 14755 21529
rect 14539 21518 14573 21519
rect 14491 21516 14573 21518
rect 14731 21518 14765 21519
rect 14766 21518 14773 21540
rect 14779 21533 14784 21540
rect 14797 21539 14811 21540
rect 14989 21539 15003 21540
rect 14789 21519 14794 21533
rect 14803 21529 14811 21533
rect 14995 21529 15003 21533
rect 14797 21519 14803 21529
rect 14989 21519 14995 21529
rect 14779 21518 14813 21519
rect 14731 21516 14813 21518
rect 14971 21518 15005 21519
rect 15006 21518 15013 21540
rect 15019 21533 15024 21540
rect 15037 21539 15051 21540
rect 15229 21539 15243 21540
rect 15029 21519 15034 21533
rect 15043 21529 15051 21533
rect 15235 21529 15243 21533
rect 15037 21519 15043 21529
rect 15229 21519 15235 21529
rect 15019 21518 15053 21519
rect 14971 21516 15053 21518
rect 15211 21518 15245 21519
rect 15246 21518 15253 21540
rect 15259 21533 15264 21540
rect 15277 21539 15291 21540
rect 15709 21539 15723 21540
rect 15269 21519 15274 21533
rect 15283 21529 15291 21533
rect 15715 21529 15723 21533
rect 15277 21519 15283 21529
rect 15709 21519 15715 21529
rect 15259 21518 15293 21519
rect 15211 21516 15293 21518
rect 15691 21518 15725 21519
rect 15726 21518 15733 21540
rect 15739 21533 15744 21540
rect 15757 21539 15771 21540
rect 15949 21539 15963 21540
rect 15749 21519 15754 21533
rect 15763 21529 15771 21533
rect 15955 21529 15963 21533
rect 15757 21519 15763 21529
rect 15949 21519 15955 21529
rect 15739 21518 15773 21519
rect 15691 21516 15773 21518
rect 15931 21518 15965 21519
rect 15966 21518 15973 21540
rect 15979 21533 15984 21540
rect 15997 21539 16011 21540
rect 16189 21539 16203 21540
rect 15989 21519 15994 21533
rect 16003 21529 16011 21533
rect 16195 21529 16203 21533
rect 15997 21519 16003 21529
rect 16189 21519 16195 21529
rect 15979 21518 16013 21519
rect 15931 21516 16013 21518
rect 16171 21518 16205 21519
rect 16206 21518 16213 21540
rect 16219 21533 16224 21540
rect 16237 21539 16251 21540
rect 16381 21539 16395 21540
rect 16229 21519 16234 21533
rect 16243 21529 16251 21533
rect 16387 21529 16395 21533
rect 16237 21519 16243 21529
rect 16381 21519 16387 21529
rect 16219 21518 16253 21519
rect 16171 21516 16253 21518
rect 16363 21518 16397 21519
rect 16398 21518 16405 21540
rect 16411 21533 16416 21540
rect 16429 21539 16443 21540
rect 25789 21539 25803 21540
rect 16421 21519 16426 21533
rect 16435 21529 16443 21533
rect 25795 21529 25803 21533
rect 16429 21519 16435 21529
rect 25789 21519 25795 21529
rect 16411 21518 16445 21519
rect 16363 21516 16445 21518
rect 25771 21518 25805 21519
rect 25806 21518 25813 21540
rect 25819 21533 25824 21540
rect 25837 21539 25851 21540
rect 25829 21519 25834 21533
rect 25843 21529 25851 21533
rect 25963 21529 25971 21533
rect 25837 21519 25843 21529
rect 25957 21519 25963 21529
rect 25819 21518 25853 21519
rect 25771 21516 25853 21518
rect 25939 21518 25973 21519
rect 25974 21518 25981 21539
rect 25987 21533 25992 21543
rect 26006 21540 26021 21543
rect 26683 21540 26717 21543
rect 26731 21540 26750 21543
rect 25997 21519 26002 21533
rect 26011 21529 26019 21533
rect 26005 21519 26011 21529
rect 26741 21519 26746 21533
rect 25987 21518 26021 21519
rect 25939 21516 26021 21518
rect 26683 21516 26717 21519
rect 6997 21515 7011 21516
rect 7014 21515 7021 21516
rect 7014 21422 7018 21515
rect 7038 21423 7042 21516
rect 7099 21509 7104 21516
rect 7117 21515 7131 21516
rect 7501 21515 7515 21516
rect 7109 21495 7114 21509
rect 7123 21505 7131 21509
rect 7507 21505 7515 21509
rect 7117 21495 7123 21505
rect 7501 21495 7507 21505
rect 7504 21491 7515 21492
rect 7518 21491 7525 21516
rect 7531 21509 7536 21516
rect 7549 21515 7563 21516
rect 8245 21515 8259 21516
rect 7541 21495 7546 21509
rect 7555 21505 7563 21509
rect 8251 21505 8259 21509
rect 7549 21495 7555 21505
rect 8245 21495 8251 21505
rect 8248 21491 8259 21492
rect 8262 21491 8269 21516
rect 8275 21509 8280 21516
rect 8293 21515 8307 21516
rect 14509 21515 14523 21516
rect 8285 21495 8290 21509
rect 8299 21505 8307 21509
rect 14515 21505 14523 21509
rect 8293 21495 8299 21505
rect 14509 21495 14515 21505
rect 7514 21461 7524 21467
rect 7526 21461 7534 21472
rect 8258 21461 8268 21467
rect 8270 21461 8278 21472
rect 14526 21461 14533 21516
rect 14539 21509 14544 21516
rect 14557 21515 14571 21516
rect 14749 21515 14763 21516
rect 14549 21495 14554 21509
rect 14563 21505 14571 21509
rect 14755 21505 14763 21509
rect 14557 21495 14563 21505
rect 14749 21495 14755 21505
rect 14766 21461 14773 21516
rect 14779 21509 14784 21516
rect 14797 21515 14811 21516
rect 14989 21515 15003 21516
rect 14789 21495 14794 21509
rect 14803 21505 14811 21509
rect 14995 21505 15003 21509
rect 14797 21495 14803 21505
rect 14989 21495 14995 21505
rect 15006 21461 15013 21516
rect 15019 21509 15024 21516
rect 15037 21515 15051 21516
rect 15229 21515 15243 21516
rect 15029 21495 15034 21509
rect 15043 21505 15051 21509
rect 15235 21505 15243 21509
rect 15037 21495 15043 21505
rect 15229 21495 15235 21505
rect 15246 21461 15253 21516
rect 15259 21509 15264 21516
rect 15277 21515 15291 21516
rect 15709 21515 15723 21516
rect 15269 21495 15274 21509
rect 15283 21505 15291 21509
rect 15715 21505 15723 21509
rect 15277 21495 15283 21505
rect 15709 21495 15715 21505
rect 15726 21461 15733 21516
rect 15739 21509 15744 21516
rect 15757 21515 15771 21516
rect 15949 21515 15963 21516
rect 15749 21495 15754 21509
rect 15763 21505 15771 21509
rect 15955 21505 15963 21509
rect 15757 21495 15763 21505
rect 15949 21495 15955 21505
rect 15952 21491 15963 21492
rect 15966 21491 15973 21516
rect 15979 21509 15984 21516
rect 15997 21515 16011 21516
rect 16189 21515 16203 21516
rect 15989 21495 15994 21509
rect 16003 21505 16011 21509
rect 16195 21505 16203 21509
rect 15997 21495 16003 21505
rect 16189 21495 16195 21505
rect 16192 21491 16203 21492
rect 16206 21491 16213 21516
rect 16219 21509 16224 21516
rect 16237 21515 16251 21516
rect 16381 21515 16395 21516
rect 16229 21495 16234 21509
rect 16243 21505 16251 21509
rect 16387 21505 16395 21509
rect 16237 21495 16243 21505
rect 16381 21495 16387 21505
rect 16384 21491 16395 21492
rect 16398 21491 16405 21516
rect 16411 21509 16416 21516
rect 16429 21515 16443 21516
rect 25789 21515 25803 21516
rect 16421 21495 16426 21509
rect 16435 21505 16443 21509
rect 25795 21505 25803 21509
rect 16429 21495 16435 21505
rect 25789 21495 25795 21505
rect 25792 21491 25803 21492
rect 25806 21491 25813 21516
rect 25819 21509 25824 21516
rect 25837 21515 25851 21516
rect 25957 21515 25971 21516
rect 25829 21495 25834 21509
rect 25843 21505 25851 21509
rect 25963 21505 25971 21509
rect 25837 21495 25843 21505
rect 25957 21495 25963 21505
rect 25960 21491 25971 21492
rect 25974 21491 25981 21516
rect 25987 21509 25992 21516
rect 26005 21515 26019 21516
rect 25997 21495 26002 21509
rect 26011 21505 26019 21509
rect 26707 21505 26715 21509
rect 26005 21495 26011 21505
rect 26701 21495 26707 21505
rect 26704 21491 26715 21492
rect 26718 21491 26725 21515
rect 26731 21509 26736 21519
rect 26750 21516 26765 21519
rect 27643 21516 27677 21519
rect 27691 21516 27710 21519
rect 26741 21495 26746 21509
rect 26755 21505 26763 21509
rect 26749 21495 26755 21505
rect 27701 21495 27706 21509
rect 15962 21461 15972 21467
rect 15974 21461 15982 21472
rect 16202 21461 16212 21467
rect 16214 21461 16222 21472
rect 16394 21461 16404 21467
rect 16406 21461 16414 21472
rect 25802 21461 25812 21467
rect 25814 21461 25822 21472
rect 25970 21461 25980 21467
rect 25982 21461 25990 21472
rect 26714 21461 26724 21467
rect 26726 21461 26734 21472
rect 27674 21461 27684 21467
rect 27686 21461 27694 21472
rect 28418 21461 28428 21467
rect 28430 21461 28438 21468
rect 29186 21461 29196 21464
rect 29978 21461 29988 21464
rect 7027 21422 7061 21423
rect 6571 21420 7061 21422
rect 3235 21413 3240 21420
rect 3301 21419 3315 21420
rect 3318 21419 3325 21420
rect 3349 21419 3363 21420
rect 3366 21419 3373 21420
rect 3245 21399 3250 21413
rect 3259 21409 3267 21413
rect 3253 21399 3259 21409
rect 3246 21398 3250 21399
rect 2677 21396 3267 21398
rect 2677 21395 2691 21396
rect 2629 21372 2691 21374
rect 2629 21371 2643 21372
rect 2646 21371 2653 21372
rect 2646 21278 2650 21368
rect 2670 21278 2674 21372
rect 2677 21371 2691 21372
rect 2694 21371 2701 21396
rect 2694 21278 2698 21371
rect 2718 21278 2722 21396
rect 2742 21278 2746 21396
rect 2766 21278 2770 21396
rect 2790 21395 2794 21396
rect 2790 21374 2797 21395
rect 2814 21374 2818 21396
rect 2773 21372 2835 21374
rect 2773 21371 2787 21372
rect 2790 21350 2797 21372
rect 2814 21350 2818 21372
rect 2821 21371 2835 21372
rect 2838 21371 2845 21395
rect 2838 21350 2842 21371
rect 2862 21350 2866 21396
rect 2886 21350 2890 21396
rect 2910 21350 2914 21396
rect 2934 21350 2938 21396
rect 2958 21395 2962 21396
rect 2958 21374 2965 21395
rect 2982 21374 2986 21396
rect 2941 21372 3003 21374
rect 2941 21371 2955 21372
rect 2958 21371 2965 21372
rect 2982 21350 2986 21372
rect 2989 21371 3003 21372
rect 3006 21371 3013 21395
rect 3006 21350 3010 21371
rect 3030 21350 3034 21396
rect 3054 21395 3058 21396
rect 3054 21374 3061 21395
rect 3078 21374 3082 21396
rect 3126 21395 3130 21396
rect 3102 21374 3109 21395
rect 3126 21374 3133 21395
rect 3150 21374 3154 21396
rect 3037 21372 3099 21374
rect 3037 21371 3051 21372
rect 3054 21371 3061 21372
rect 3078 21350 3082 21372
rect 3085 21371 3099 21372
rect 3102 21372 3171 21374
rect 3102 21371 3123 21372
rect 3126 21371 3133 21372
rect 3102 21351 3106 21371
rect 3091 21350 3125 21351
rect 2773 21348 3125 21350
rect 2773 21347 2787 21348
rect 2790 21347 2797 21348
rect 2790 21278 2794 21347
rect 2814 21278 2818 21348
rect 2838 21278 2842 21348
rect 2862 21278 2866 21348
rect 2886 21278 2890 21348
rect 2910 21278 2914 21348
rect 2934 21278 2938 21348
rect 2958 21278 2962 21346
rect 2982 21278 2986 21348
rect 3006 21278 3010 21348
rect 3030 21278 3034 21348
rect 3054 21278 3058 21346
rect 3078 21278 3082 21348
rect 3091 21341 3096 21348
rect 3102 21341 3106 21348
rect 3101 21327 3106 21341
rect 3115 21336 3120 21337
rect 3091 21317 3096 21327
rect 3101 21303 3106 21317
rect 3102 21278 3106 21303
rect 3126 21278 3130 21346
rect 3150 21278 3154 21372
rect 3157 21371 3171 21372
rect 3174 21371 3181 21395
rect 3174 21278 3178 21371
rect 3198 21278 3202 21396
rect 3222 21278 3226 21396
rect 3246 21278 3250 21396
rect 3253 21395 3267 21396
rect 3270 21395 3277 21419
rect 3379 21413 3384 21420
rect 3397 21419 3411 21420
rect 3829 21419 3843 21420
rect 3846 21419 3853 21420
rect 3859 21413 3864 21420
rect 3877 21419 3891 21420
rect 4549 21419 4563 21420
rect 4566 21419 4573 21420
rect 4579 21413 4584 21420
rect 4597 21419 4611 21420
rect 4789 21419 4803 21420
rect 4806 21419 4813 21420
rect 4819 21413 4824 21420
rect 4837 21419 4851 21420
rect 6589 21419 6603 21420
rect 6606 21419 6613 21420
rect 3389 21399 3394 21413
rect 3869 21399 3874 21413
rect 4589 21399 4594 21413
rect 4829 21399 4834 21413
rect 3270 21371 3274 21395
rect 3283 21372 3302 21375
rect 3270 21326 3277 21371
rect 3293 21351 3298 21365
rect 3318 21358 3322 21392
rect 3379 21389 3384 21399
rect 3859 21389 3864 21399
rect 4579 21389 4584 21399
rect 4819 21389 4824 21399
rect 3389 21375 3394 21389
rect 3869 21375 3874 21389
rect 4589 21375 4594 21389
rect 4829 21375 4834 21389
rect 3379 21365 3384 21375
rect 3859 21365 3864 21375
rect 4579 21365 4584 21375
rect 4819 21365 4824 21375
rect 3341 21351 3346 21365
rect 3389 21351 3394 21365
rect 3869 21351 3874 21365
rect 4589 21351 4594 21365
rect 4829 21351 4834 21365
rect 3294 21326 3298 21351
rect 3342 21326 3346 21351
rect 3380 21338 3384 21348
rect 3390 21326 3394 21338
rect 3835 21337 3843 21341
rect 3829 21327 3835 21337
rect 3403 21326 3437 21327
rect 3253 21324 3437 21326
rect 3811 21326 3845 21327
rect 3846 21326 3853 21347
rect 3859 21341 3864 21351
rect 3869 21327 3874 21341
rect 3883 21337 3891 21341
rect 4555 21337 4563 21341
rect 3877 21327 3883 21337
rect 4549 21327 4555 21337
rect 3859 21326 3893 21327
rect 3811 21324 3893 21326
rect 4531 21326 4565 21327
rect 4566 21326 4573 21347
rect 4579 21341 4584 21351
rect 4589 21327 4594 21341
rect 4603 21337 4611 21341
rect 4795 21337 4803 21341
rect 4597 21327 4603 21337
rect 4789 21327 4795 21337
rect 4579 21326 4613 21327
rect 4531 21324 4613 21326
rect 4771 21326 4805 21327
rect 4806 21326 4813 21347
rect 4819 21341 4824 21351
rect 4829 21327 4834 21341
rect 4843 21337 4851 21341
rect 6595 21337 6603 21341
rect 4837 21327 4843 21337
rect 6589 21327 6595 21337
rect 4819 21326 4853 21327
rect 4771 21324 4853 21326
rect 6571 21326 6605 21327
rect 6606 21326 6613 21347
rect 6726 21326 6730 21420
rect 6750 21326 6754 21420
rect 6774 21326 6778 21420
rect 6798 21326 6802 21420
rect 6822 21326 6826 21420
rect 6846 21326 6850 21420
rect 6870 21326 6874 21420
rect 6894 21326 6898 21420
rect 6918 21326 6922 21420
rect 6942 21327 6946 21420
rect 6955 21341 6960 21351
rect 6966 21341 6970 21420
rect 6979 21365 6984 21375
rect 6990 21365 6994 21420
rect 7003 21389 7008 21399
rect 7014 21389 7018 21420
rect 7027 21413 7032 21420
rect 7038 21413 7042 21420
rect 7037 21399 7042 21413
rect 7013 21375 7018 21389
rect 6989 21351 6994 21365
rect 6965 21327 6970 21341
rect 6931 21326 6965 21327
rect 6571 21324 6965 21326
rect 3253 21323 3267 21324
rect 3270 21323 3277 21324
rect 3270 21278 3274 21323
rect 3294 21278 3298 21324
rect -2393 21276 3315 21278
rect -2371 21254 -2366 21276
rect -2348 21254 -2343 21276
rect -2325 21254 -2320 21276
rect -2054 21275 -1906 21276
rect -2054 21274 -2036 21275
rect -2309 21260 -2301 21270
rect -2317 21254 -2309 21260
rect -2068 21259 -2038 21266
rect -2000 21258 -1992 21275
rect -1920 21274 -1906 21275
rect -1846 21268 -1794 21276
rect -1852 21261 -1804 21266
rect -1902 21259 -1804 21261
rect -1655 21260 -1647 21270
rect -2000 21256 -1975 21258
rect -1902 21257 -1852 21259
rect -2025 21254 -1975 21256
rect -1846 21254 -1804 21257
rect -1663 21254 -1655 21260
rect -1642 21254 -1637 21276
rect -1619 21254 -1614 21276
rect -1530 21254 -1526 21276
rect -1506 21254 -1502 21276
rect -1482 21254 -1478 21276
rect -1458 21254 -1454 21276
rect -1434 21254 -1430 21276
rect -1410 21254 -1406 21276
rect -1386 21254 -1382 21276
rect -1362 21254 -1358 21276
rect -1338 21254 -1334 21276
rect -1314 21254 -1310 21276
rect -1290 21254 -1286 21276
rect -1266 21254 -1262 21276
rect -1242 21254 -1238 21276
rect -1218 21254 -1214 21276
rect -1194 21254 -1190 21276
rect -1170 21254 -1166 21276
rect -1146 21254 -1142 21276
rect -1122 21254 -1118 21276
rect -1098 21254 -1094 21276
rect -1074 21254 -1070 21276
rect -1050 21254 -1046 21276
rect -1026 21254 -1022 21276
rect -1002 21254 -998 21276
rect -978 21254 -974 21276
rect -954 21254 -950 21276
rect -930 21254 -926 21276
rect -906 21254 -902 21276
rect -882 21254 -878 21276
rect -858 21254 -854 21276
rect -834 21254 -830 21276
rect -810 21254 -806 21276
rect -786 21254 -782 21276
rect -762 21254 -758 21276
rect -738 21254 -734 21276
rect -714 21254 -710 21276
rect -690 21254 -686 21276
rect -666 21254 -662 21276
rect -642 21254 -638 21276
rect -618 21254 -614 21276
rect -594 21254 -590 21276
rect -570 21254 -566 21276
rect -546 21254 -542 21276
rect -522 21254 -518 21276
rect -498 21254 -494 21276
rect -474 21254 -470 21276
rect -450 21254 -446 21276
rect -426 21254 -422 21276
rect -402 21254 -398 21276
rect -378 21254 -374 21276
rect -354 21254 -350 21276
rect -330 21254 -326 21276
rect -306 21254 -302 21276
rect -282 21254 -278 21276
rect -258 21254 -254 21276
rect -234 21254 -230 21276
rect -210 21254 -206 21276
rect -186 21254 -182 21276
rect -162 21254 -158 21276
rect -138 21254 -134 21276
rect -114 21254 -110 21276
rect -90 21254 -86 21276
rect -66 21254 -62 21276
rect -42 21254 -38 21276
rect -18 21254 -14 21276
rect 6 21254 10 21276
rect 30 21254 34 21276
rect 54 21254 58 21276
rect 78 21254 82 21276
rect 102 21254 106 21276
rect 126 21254 130 21276
rect 150 21254 154 21276
rect 174 21254 178 21276
rect 198 21254 202 21276
rect 222 21254 226 21276
rect 246 21254 250 21276
rect 270 21254 274 21276
rect 294 21254 298 21276
rect 318 21254 322 21276
rect 342 21254 346 21276
rect 366 21254 370 21276
rect 390 21254 394 21276
rect 414 21254 418 21276
rect 438 21254 442 21276
rect 462 21254 466 21276
rect 486 21254 490 21276
rect 510 21254 514 21276
rect 534 21254 538 21276
rect 558 21254 562 21276
rect 582 21254 586 21276
rect 606 21254 610 21276
rect 630 21254 634 21276
rect 654 21254 658 21276
rect 678 21254 682 21276
rect 702 21254 706 21276
rect 726 21254 730 21276
rect 750 21254 754 21276
rect 774 21254 778 21276
rect 798 21254 802 21276
rect 822 21254 826 21276
rect 846 21254 850 21276
rect 870 21254 874 21276
rect 894 21254 898 21276
rect 918 21254 922 21276
rect 942 21254 946 21276
rect 966 21254 970 21276
rect 990 21254 994 21276
rect 1014 21254 1018 21276
rect 1038 21254 1042 21276
rect 1062 21254 1066 21276
rect 1086 21254 1090 21276
rect 1110 21254 1114 21276
rect 1134 21254 1138 21276
rect 1158 21254 1162 21276
rect 1182 21254 1186 21276
rect 1206 21254 1210 21276
rect 1230 21254 1234 21276
rect 1254 21254 1258 21276
rect 1278 21254 1282 21276
rect 1302 21254 1306 21276
rect 1326 21254 1330 21276
rect 1350 21254 1354 21276
rect 1374 21254 1378 21276
rect 1398 21254 1402 21276
rect 1422 21254 1426 21276
rect 1446 21254 1450 21276
rect 1470 21255 1474 21276
rect 1459 21254 1493 21255
rect -2393 21252 1493 21254
rect -2371 21230 -2366 21252
rect -2348 21230 -2343 21252
rect -2325 21230 -2320 21252
rect -2054 21251 -2038 21252
rect -2000 21251 -1966 21252
rect -1846 21251 -1804 21252
rect -2000 21250 -1975 21251
rect -2076 21242 -2054 21249
rect -2309 21232 -2301 21242
rect -2044 21239 -2038 21244
rect -2028 21242 -2001 21249
rect -2054 21232 -2038 21239
rect -2015 21241 -2001 21242
rect -2015 21232 -2014 21241
rect -2317 21230 -2309 21232
rect -2044 21230 -2028 21232
rect -2000 21230 -1992 21250
rect -1982 21249 -1975 21250
rect -1862 21249 -1798 21250
rect -1985 21242 -1796 21249
rect -1862 21241 -1798 21242
rect -1852 21232 -1804 21239
rect -1655 21232 -1647 21242
rect -1976 21230 -1940 21231
rect -1663 21230 -1655 21232
rect -1642 21230 -1637 21252
rect -1619 21230 -1614 21252
rect -1530 21230 -1526 21252
rect -1506 21230 -1502 21252
rect -1482 21251 -1478 21252
rect -2393 21228 -1485 21230
rect -2371 21158 -2366 21228
rect -2348 21158 -2343 21228
rect -2325 21194 -2320 21228
rect -2317 21226 -2309 21228
rect -2076 21215 -2054 21222
rect -2325 21186 -2317 21194
rect -2060 21188 -2030 21191
rect -2325 21158 -2320 21186
rect -2317 21178 -2309 21186
rect -2060 21175 -2038 21186
rect -2033 21179 -2030 21188
rect -2028 21184 -2027 21188
rect -2068 21170 -2038 21173
rect -2000 21158 -1992 21228
rect -1846 21224 -1804 21228
rect -1663 21226 -1655 21228
rect -1846 21214 -1794 21223
rect -1912 21203 -1884 21205
rect -1852 21197 -1804 21201
rect -1844 21188 -1796 21191
rect -1671 21186 -1663 21194
rect -1844 21175 -1804 21186
rect -1663 21178 -1655 21186
rect -1852 21170 -1680 21174
rect -1642 21158 -1637 21228
rect -1619 21158 -1614 21228
rect -1530 21158 -1526 21228
rect -1506 21158 -1502 21228
rect -1499 21227 -1485 21228
rect -1482 21227 -1475 21251
rect -1482 21158 -1478 21227
rect -1458 21158 -1454 21252
rect -1434 21158 -1430 21252
rect -1410 21158 -1406 21252
rect -1386 21158 -1382 21252
rect -1362 21158 -1358 21252
rect -1338 21158 -1334 21252
rect -1314 21158 -1310 21252
rect -1290 21158 -1286 21252
rect -1266 21158 -1262 21252
rect -1242 21158 -1238 21252
rect -1218 21158 -1214 21252
rect -1194 21158 -1190 21252
rect -1170 21158 -1166 21252
rect -1146 21158 -1142 21252
rect -1122 21158 -1118 21252
rect -1098 21158 -1094 21252
rect -1074 21158 -1070 21252
rect -1050 21158 -1046 21252
rect -1026 21158 -1022 21252
rect -1002 21158 -998 21252
rect -978 21158 -974 21252
rect -954 21158 -950 21252
rect -930 21158 -926 21252
rect -906 21158 -902 21252
rect -882 21158 -878 21252
rect -858 21158 -854 21252
rect -834 21158 -830 21252
rect -810 21158 -806 21252
rect -786 21158 -782 21252
rect -762 21158 -758 21252
rect -738 21158 -734 21252
rect -714 21158 -710 21252
rect -690 21158 -686 21252
rect -666 21158 -662 21252
rect -642 21158 -638 21252
rect -618 21158 -614 21252
rect -594 21158 -590 21252
rect -570 21158 -566 21252
rect -546 21158 -542 21252
rect -522 21158 -518 21252
rect -498 21158 -494 21252
rect -474 21158 -470 21252
rect -450 21158 -446 21252
rect -426 21158 -422 21252
rect -402 21158 -398 21252
rect -378 21158 -374 21252
rect -354 21158 -350 21252
rect -330 21158 -326 21252
rect -306 21158 -302 21252
rect -282 21158 -278 21252
rect -258 21158 -254 21252
rect -234 21158 -230 21252
rect -210 21158 -206 21252
rect -186 21158 -182 21252
rect -162 21158 -158 21252
rect -138 21158 -134 21252
rect -114 21158 -110 21252
rect -90 21158 -86 21252
rect -66 21158 -62 21252
rect -42 21158 -38 21252
rect -18 21158 -14 21252
rect 6 21158 10 21252
rect 30 21158 34 21252
rect 54 21158 58 21252
rect 78 21158 82 21252
rect 102 21158 106 21252
rect 126 21158 130 21252
rect 150 21158 154 21252
rect 174 21158 178 21252
rect 198 21158 202 21252
rect 222 21158 226 21252
rect 246 21158 250 21252
rect 270 21158 274 21252
rect 294 21158 298 21252
rect 318 21158 322 21252
rect 342 21158 346 21252
rect 366 21158 370 21252
rect 390 21158 394 21252
rect 414 21158 418 21252
rect 438 21158 442 21252
rect 462 21158 466 21252
rect 486 21158 490 21252
rect 510 21158 514 21252
rect 534 21158 538 21252
rect 558 21158 562 21252
rect 582 21158 586 21252
rect 606 21158 610 21252
rect 630 21158 634 21252
rect 654 21158 658 21252
rect 678 21158 682 21252
rect 702 21158 706 21252
rect 726 21158 730 21252
rect 750 21158 754 21252
rect 774 21158 778 21252
rect 798 21158 802 21252
rect 822 21158 826 21252
rect 846 21158 850 21252
rect 870 21158 874 21252
rect 894 21158 898 21252
rect 918 21158 922 21252
rect 942 21158 946 21252
rect 966 21158 970 21252
rect 990 21158 994 21252
rect 1014 21158 1018 21252
rect 1038 21158 1042 21252
rect 1062 21158 1066 21252
rect 1086 21158 1090 21252
rect 1110 21158 1114 21252
rect 1134 21158 1138 21252
rect 1158 21158 1162 21252
rect 1182 21158 1186 21252
rect 1206 21158 1210 21252
rect 1230 21158 1234 21252
rect 1243 21197 1248 21207
rect 1254 21197 1258 21252
rect 1267 21221 1272 21231
rect 1278 21221 1282 21252
rect 1277 21207 1282 21221
rect 1267 21197 1272 21207
rect 1253 21183 1258 21197
rect 1277 21183 1282 21197
rect 1243 21182 1277 21183
rect 1278 21182 1282 21183
rect 1302 21182 1306 21252
rect 1326 21182 1330 21252
rect 1350 21182 1354 21252
rect 1374 21182 1378 21252
rect 1398 21182 1402 21252
rect 1422 21182 1426 21252
rect 1446 21182 1450 21252
rect 1459 21245 1464 21252
rect 1470 21245 1474 21252
rect 1469 21231 1474 21245
rect 1459 21221 1464 21231
rect 1469 21207 1474 21221
rect 1470 21182 1474 21207
rect 1494 21182 1498 21276
rect 1518 21182 1522 21276
rect 1542 21182 1546 21276
rect 1566 21182 1570 21276
rect 1590 21182 1594 21276
rect 1614 21182 1618 21276
rect 1638 21182 1642 21276
rect 1662 21182 1666 21276
rect 1686 21182 1690 21276
rect 1710 21182 1714 21276
rect 1734 21182 1738 21276
rect 1758 21182 1762 21276
rect 1782 21182 1786 21276
rect 1806 21182 1810 21276
rect 1830 21182 1834 21276
rect 1854 21182 1858 21276
rect 1878 21182 1882 21276
rect 1902 21182 1906 21276
rect 1926 21182 1930 21276
rect 1950 21182 1954 21276
rect 1974 21182 1978 21276
rect 1998 21182 2002 21276
rect 2022 21182 2026 21276
rect 2046 21182 2050 21276
rect 2070 21182 2074 21276
rect 2094 21182 2098 21276
rect 2118 21182 2122 21276
rect 2142 21182 2146 21276
rect 2166 21182 2170 21276
rect 2190 21182 2194 21276
rect 2214 21182 2218 21276
rect 2238 21182 2242 21276
rect 2262 21182 2266 21276
rect 2286 21182 2290 21276
rect 2310 21182 2314 21276
rect 2334 21182 2338 21276
rect 2358 21182 2362 21276
rect 2382 21182 2386 21276
rect 2406 21182 2410 21276
rect 2430 21182 2434 21276
rect 2454 21182 2458 21276
rect 2478 21182 2482 21276
rect 2502 21182 2506 21276
rect 2526 21182 2530 21276
rect 2550 21182 2554 21276
rect 2574 21182 2578 21276
rect 2598 21182 2602 21276
rect 2622 21182 2626 21276
rect 2646 21182 2650 21276
rect 2670 21182 2674 21276
rect 2694 21182 2698 21276
rect 2718 21182 2722 21276
rect 2742 21182 2746 21276
rect 2766 21182 2770 21276
rect 2790 21182 2794 21276
rect 2814 21182 2818 21276
rect 2838 21182 2842 21276
rect 2862 21182 2866 21276
rect 2886 21182 2890 21276
rect 2910 21182 2914 21276
rect 2934 21182 2938 21276
rect 2958 21182 2962 21276
rect 2982 21182 2986 21276
rect 3006 21182 3010 21276
rect 3030 21182 3034 21276
rect 3054 21182 3058 21276
rect 3078 21182 3082 21276
rect 3102 21182 3106 21276
rect 3126 21275 3130 21276
rect 3126 21230 3133 21275
rect 3150 21230 3154 21276
rect 3174 21230 3178 21276
rect 3198 21230 3202 21276
rect 3222 21230 3226 21276
rect 3246 21230 3250 21276
rect 3270 21230 3274 21276
rect 3294 21230 3298 21276
rect 3301 21275 3315 21276
rect 3318 21275 3325 21299
rect 3318 21230 3322 21275
rect 3342 21230 3346 21324
rect 3366 21278 3373 21299
rect 3390 21278 3394 21324
rect 3397 21323 3411 21324
rect 3829 21323 3843 21324
rect 3413 21310 3421 21317
rect 3835 21313 3843 21317
rect 3413 21304 3415 21310
rect 3413 21303 3421 21304
rect 3829 21303 3835 21313
rect 3811 21302 3845 21303
rect 3846 21302 3853 21324
rect 3859 21317 3864 21324
rect 3877 21323 3891 21324
rect 4549 21323 4563 21324
rect 3869 21303 3874 21317
rect 3883 21313 3891 21317
rect 4555 21313 4563 21317
rect 3877 21303 3883 21313
rect 4549 21303 4555 21313
rect 3859 21302 3893 21303
rect 3811 21300 3893 21302
rect 4531 21302 4565 21303
rect 4566 21302 4573 21324
rect 4579 21317 4584 21324
rect 4597 21323 4611 21324
rect 4789 21323 4803 21324
rect 4589 21303 4594 21317
rect 4603 21313 4611 21317
rect 4795 21313 4803 21317
rect 4597 21303 4603 21313
rect 4789 21303 4795 21313
rect 4579 21302 4613 21303
rect 4531 21300 4613 21302
rect 4771 21302 4805 21303
rect 4806 21302 4813 21324
rect 4819 21317 4824 21324
rect 4837 21323 4851 21324
rect 6589 21323 6603 21324
rect 4829 21303 4834 21317
rect 4843 21313 4851 21317
rect 6595 21313 6603 21317
rect 4837 21303 4843 21313
rect 6589 21303 6595 21313
rect 4819 21302 4853 21303
rect 4771 21300 4853 21302
rect 6571 21302 6605 21303
rect 6606 21302 6613 21324
rect 6726 21302 6730 21324
rect 6750 21302 6754 21324
rect 6774 21302 6778 21324
rect 6798 21302 6802 21324
rect 6822 21302 6826 21324
rect 6846 21302 6850 21324
rect 6870 21302 6874 21324
rect 6894 21302 6898 21324
rect 6918 21303 6922 21324
rect 6931 21317 6936 21324
rect 6942 21317 6946 21324
rect 6941 21303 6946 21317
rect 6907 21302 6941 21303
rect 6571 21300 6941 21302
rect 3404 21299 3411 21300
rect 3829 21299 3843 21300
rect 3414 21286 3421 21290
rect 3835 21289 3843 21293
rect 3829 21279 3835 21289
rect 3349 21276 3411 21278
rect 3427 21276 3461 21279
rect 3811 21278 3845 21279
rect 3846 21278 3853 21300
rect 3859 21293 3864 21300
rect 3877 21299 3891 21300
rect 4549 21299 4563 21300
rect 3869 21279 3874 21293
rect 3883 21289 3891 21293
rect 4555 21289 4563 21293
rect 3877 21279 3883 21289
rect 4549 21279 4555 21289
rect 3859 21278 3893 21279
rect 3811 21276 3893 21278
rect 4531 21278 4565 21279
rect 4566 21278 4573 21300
rect 4579 21293 4584 21300
rect 4597 21299 4611 21300
rect 4789 21299 4803 21300
rect 4589 21279 4594 21293
rect 4603 21289 4611 21293
rect 4795 21289 4803 21293
rect 4597 21279 4603 21289
rect 4789 21279 4795 21289
rect 4579 21278 4613 21279
rect 4531 21276 4613 21278
rect 4771 21278 4805 21279
rect 4806 21278 4813 21300
rect 4819 21293 4824 21300
rect 4837 21299 4851 21300
rect 6589 21299 6603 21300
rect 4829 21279 4834 21293
rect 4843 21289 4851 21293
rect 6595 21289 6603 21293
rect 4837 21279 4843 21289
rect 6589 21279 6595 21289
rect 4819 21278 4853 21279
rect 4771 21276 4853 21278
rect 6571 21278 6605 21279
rect 6606 21278 6613 21300
rect 6726 21278 6730 21300
rect 6750 21278 6754 21300
rect 6774 21278 6778 21300
rect 6798 21278 6802 21300
rect 6822 21278 6826 21300
rect 6846 21278 6850 21300
rect 6870 21278 6874 21300
rect 6894 21279 6898 21300
rect 6907 21293 6912 21300
rect 6918 21293 6922 21300
rect 6917 21279 6922 21293
rect 6883 21278 6917 21279
rect 6571 21276 6917 21278
rect 3349 21275 3363 21276
rect 3366 21275 3373 21276
rect 3366 21230 3370 21275
rect 3390 21230 3394 21276
rect 3397 21275 3411 21276
rect 3414 21275 3421 21276
rect 3829 21275 3843 21276
rect 3835 21265 3843 21269
rect 3829 21255 3835 21265
rect 3811 21254 3845 21255
rect 3846 21254 3853 21276
rect 3859 21269 3864 21276
rect 3877 21275 3891 21276
rect 4549 21275 4563 21276
rect 3869 21255 3874 21269
rect 3883 21265 3891 21269
rect 4555 21265 4563 21269
rect 3877 21255 3883 21265
rect 4549 21255 4555 21265
rect 3859 21254 3893 21255
rect 3811 21252 3893 21254
rect 4531 21254 4565 21255
rect 4566 21254 4573 21276
rect 4579 21269 4584 21276
rect 4597 21275 4611 21276
rect 4789 21275 4803 21276
rect 4589 21255 4594 21269
rect 4603 21265 4611 21269
rect 4795 21265 4803 21269
rect 4597 21255 4603 21265
rect 4789 21255 4795 21265
rect 4579 21254 4613 21255
rect 4531 21252 4613 21254
rect 4771 21254 4805 21255
rect 4806 21254 4813 21276
rect 4819 21269 4824 21276
rect 4837 21275 4851 21276
rect 6589 21275 6603 21276
rect 4829 21255 4834 21269
rect 4843 21265 4851 21269
rect 6595 21265 6603 21269
rect 4837 21255 4843 21265
rect 6589 21255 6595 21265
rect 4819 21254 4853 21255
rect 4771 21252 4853 21254
rect 6571 21254 6605 21255
rect 6606 21254 6613 21276
rect 6726 21254 6730 21276
rect 6750 21254 6754 21276
rect 6774 21254 6778 21276
rect 6798 21254 6802 21276
rect 6822 21254 6826 21276
rect 6846 21254 6850 21276
rect 6870 21255 6874 21276
rect 6883 21269 6888 21276
rect 6894 21269 6898 21276
rect 6893 21255 6898 21269
rect 6859 21254 6893 21255
rect 6571 21252 6893 21254
rect 3414 21230 3418 21252
rect 3829 21251 3843 21252
rect 3438 21238 3445 21251
rect 3835 21241 3843 21245
rect 3829 21231 3835 21241
rect 3109 21228 3435 21230
rect 3499 21228 3533 21231
rect 3811 21230 3845 21231
rect 3846 21230 3853 21252
rect 3859 21245 3864 21252
rect 3877 21251 3891 21252
rect 4549 21251 4563 21252
rect 3869 21231 3874 21245
rect 3883 21241 3891 21245
rect 4555 21241 4563 21245
rect 3877 21231 3883 21241
rect 4549 21231 4555 21241
rect 3859 21230 3893 21231
rect 3811 21228 3893 21230
rect 4531 21230 4565 21231
rect 4566 21230 4573 21252
rect 4579 21245 4584 21252
rect 4597 21251 4611 21252
rect 4789 21251 4803 21252
rect 4589 21231 4594 21245
rect 4603 21241 4611 21245
rect 4795 21241 4803 21245
rect 4597 21231 4603 21241
rect 4789 21231 4795 21241
rect 4579 21230 4613 21231
rect 4531 21228 4613 21230
rect 4771 21230 4805 21231
rect 4806 21230 4813 21252
rect 4819 21245 4824 21252
rect 4837 21251 4851 21252
rect 6589 21251 6603 21252
rect 4829 21231 4834 21245
rect 4843 21241 4851 21245
rect 6595 21241 6603 21245
rect 4837 21231 4843 21241
rect 6589 21231 6595 21241
rect 4819 21230 4853 21231
rect 4771 21228 4853 21230
rect 6571 21230 6605 21231
rect 6606 21230 6613 21252
rect 6726 21230 6730 21252
rect 6750 21230 6754 21252
rect 6774 21230 6778 21252
rect 6798 21230 6802 21252
rect 6822 21230 6826 21252
rect 6846 21231 6850 21252
rect 6859 21245 6864 21252
rect 6870 21245 6874 21252
rect 6869 21231 6874 21245
rect 6835 21230 6869 21231
rect 6571 21228 6869 21230
rect 3109 21227 3123 21228
rect 3126 21227 3133 21228
rect 3126 21182 3130 21227
rect 3150 21182 3154 21228
rect 3174 21182 3178 21228
rect 3198 21182 3202 21228
rect 3222 21182 3226 21228
rect 3246 21182 3250 21228
rect 3270 21182 3274 21228
rect 3294 21182 3298 21228
rect 3318 21182 3322 21228
rect 3342 21182 3346 21228
rect 3366 21182 3370 21228
rect 3390 21182 3394 21228
rect 3414 21182 3418 21228
rect 3421 21227 3435 21228
rect 3438 21227 3445 21228
rect 3829 21227 3843 21228
rect 3835 21217 3843 21221
rect 3829 21207 3835 21217
rect 3499 21204 3533 21207
rect 3811 21206 3845 21207
rect 3846 21206 3853 21228
rect 3859 21221 3864 21228
rect 3877 21227 3891 21228
rect 4549 21227 4563 21228
rect 3869 21207 3874 21221
rect 3883 21217 3891 21221
rect 4555 21217 4563 21221
rect 3877 21207 3883 21217
rect 4549 21207 4555 21217
rect 3859 21206 3893 21207
rect 3811 21204 3893 21206
rect 4531 21206 4565 21207
rect 4566 21206 4573 21228
rect 4579 21221 4584 21228
rect 4597 21227 4611 21228
rect 4789 21227 4803 21228
rect 4589 21207 4594 21221
rect 4603 21217 4611 21221
rect 4795 21217 4803 21221
rect 4597 21207 4603 21217
rect 4789 21207 4795 21217
rect 4579 21206 4613 21207
rect 4531 21204 4613 21206
rect 4771 21206 4805 21207
rect 4806 21206 4813 21228
rect 4819 21221 4824 21228
rect 4837 21227 4851 21228
rect 6589 21227 6603 21228
rect 4829 21207 4834 21221
rect 4843 21217 4851 21221
rect 6595 21217 6603 21221
rect 4837 21207 4843 21217
rect 6589 21207 6595 21217
rect 4819 21206 4853 21207
rect 4771 21204 4853 21206
rect 6571 21206 6605 21207
rect 6606 21206 6613 21228
rect 6726 21206 6730 21228
rect 6750 21206 6754 21228
rect 6774 21206 6778 21228
rect 6798 21206 6802 21228
rect 6822 21207 6826 21228
rect 6835 21221 6840 21228
rect 6846 21221 6850 21228
rect 6845 21207 6850 21221
rect 6811 21206 6845 21207
rect 6571 21204 6845 21206
rect 3438 21182 3442 21204
rect 3829 21203 3843 21204
rect 1243 21180 3459 21182
rect 1243 21173 1248 21180
rect 1253 21159 1258 21173
rect 1254 21158 1258 21159
rect 1278 21158 1282 21180
rect 1302 21158 1306 21180
rect 1326 21158 1330 21180
rect 1350 21158 1354 21180
rect 1374 21158 1378 21180
rect 1398 21158 1402 21180
rect 1422 21158 1426 21180
rect 1446 21158 1450 21180
rect 1470 21158 1474 21180
rect 1494 21179 1498 21180
rect -2393 21156 1491 21158
rect -2371 21134 -2366 21156
rect -2348 21134 -2343 21156
rect -2325 21134 -2320 21156
rect -2309 21138 -2301 21148
rect -2068 21139 -2062 21144
rect -2317 21134 -2309 21138
rect -2060 21134 -2050 21139
rect -2000 21134 -1992 21156
rect -1806 21148 -1680 21154
rect -1854 21139 -1806 21144
rect -1655 21138 -1647 21148
rect -1972 21134 -1964 21135
rect -1958 21134 -1942 21136
rect -1844 21134 -1806 21137
rect -1663 21134 -1655 21138
rect -1642 21134 -1637 21156
rect -1619 21134 -1614 21156
rect -1530 21134 -1526 21156
rect -1506 21134 -1502 21156
rect -1482 21134 -1478 21156
rect -1458 21134 -1454 21156
rect -1434 21134 -1430 21156
rect -1410 21134 -1406 21156
rect -1386 21134 -1382 21156
rect -1362 21134 -1358 21156
rect -1338 21134 -1334 21156
rect -1314 21134 -1310 21156
rect -1290 21134 -1286 21156
rect -1266 21134 -1262 21156
rect -1242 21134 -1238 21156
rect -1218 21134 -1214 21156
rect -1194 21134 -1190 21156
rect -1170 21134 -1166 21156
rect -1146 21134 -1142 21156
rect -1122 21134 -1118 21156
rect -1098 21134 -1094 21156
rect -1074 21134 -1070 21156
rect -1050 21134 -1046 21156
rect -1026 21134 -1022 21156
rect -1002 21134 -998 21156
rect -978 21134 -974 21156
rect -954 21134 -950 21156
rect -930 21134 -926 21156
rect -906 21134 -902 21156
rect -882 21134 -878 21156
rect -858 21134 -854 21156
rect -834 21134 -830 21156
rect -810 21134 -806 21156
rect -786 21134 -782 21156
rect -762 21134 -758 21156
rect -738 21134 -734 21156
rect -714 21134 -710 21156
rect -690 21134 -686 21156
rect -666 21134 -662 21156
rect -642 21134 -638 21156
rect -618 21134 -614 21156
rect -594 21134 -590 21156
rect -570 21134 -566 21156
rect -546 21134 -542 21156
rect -522 21134 -518 21156
rect -498 21134 -494 21156
rect -474 21134 -470 21156
rect -450 21134 -446 21156
rect -426 21134 -422 21156
rect -402 21134 -398 21156
rect -378 21134 -374 21156
rect -354 21134 -350 21156
rect -330 21134 -326 21156
rect -306 21134 -302 21156
rect -282 21134 -278 21156
rect -258 21134 -254 21156
rect -234 21134 -230 21156
rect -210 21134 -206 21156
rect -186 21134 -182 21156
rect -162 21134 -158 21156
rect -138 21134 -134 21156
rect -114 21134 -110 21156
rect -90 21134 -86 21156
rect -66 21134 -62 21156
rect -42 21134 -38 21156
rect -18 21134 -14 21156
rect 6 21134 10 21156
rect 30 21134 34 21156
rect 54 21134 58 21156
rect 78 21134 82 21156
rect 102 21134 106 21156
rect 126 21134 130 21156
rect 150 21134 154 21156
rect 174 21134 178 21156
rect 198 21134 202 21156
rect 222 21134 226 21156
rect 246 21134 250 21156
rect 270 21134 274 21156
rect 294 21134 298 21156
rect 318 21134 322 21156
rect 342 21134 346 21156
rect 366 21134 370 21156
rect 390 21134 394 21156
rect 414 21134 418 21156
rect 438 21134 442 21156
rect 462 21134 466 21156
rect 486 21134 490 21156
rect 510 21134 514 21156
rect 534 21134 538 21156
rect 558 21134 562 21156
rect 582 21134 586 21156
rect 606 21134 610 21156
rect 630 21134 634 21156
rect 654 21134 658 21156
rect 678 21134 682 21156
rect 702 21134 706 21156
rect 726 21134 730 21156
rect 750 21134 754 21156
rect 774 21134 778 21156
rect 798 21135 802 21156
rect 787 21134 821 21135
rect -2393 21132 821 21134
rect -2371 21110 -2366 21132
rect -2348 21110 -2343 21132
rect -2325 21110 -2320 21132
rect -2060 21126 -2050 21132
rect -2309 21110 -2301 21120
rect -2060 21119 -2030 21126
rect -2000 21122 -1992 21132
rect -1972 21130 -1942 21132
rect -1958 21129 -1942 21130
rect -1844 21128 -1806 21132
rect -2068 21112 -2062 21119
rect -2062 21110 -2036 21112
rect -2393 21108 -2036 21110
rect -2030 21110 -2012 21112
rect -2004 21110 -1990 21122
rect -1844 21121 -1798 21126
rect -1806 21119 -1798 21121
rect -1854 21117 -1844 21119
rect -1854 21112 -1806 21117
rect -1864 21110 -1796 21111
rect -1655 21110 -1647 21120
rect -1642 21110 -1637 21132
rect -1619 21110 -1614 21132
rect -1530 21110 -1526 21132
rect -1506 21110 -1502 21132
rect -1482 21110 -1478 21132
rect -1458 21110 -1454 21132
rect -1434 21110 -1430 21132
rect -1410 21110 -1406 21132
rect -1386 21110 -1382 21132
rect -1362 21110 -1358 21132
rect -1338 21110 -1334 21132
rect -1314 21110 -1310 21132
rect -1290 21110 -1286 21132
rect -1266 21110 -1262 21132
rect -1242 21110 -1238 21132
rect -1218 21110 -1214 21132
rect -1194 21110 -1190 21132
rect -1170 21110 -1166 21132
rect -1146 21110 -1142 21132
rect -1122 21110 -1118 21132
rect -1098 21110 -1094 21132
rect -1074 21110 -1070 21132
rect -1050 21110 -1046 21132
rect -1026 21110 -1022 21132
rect -1002 21110 -998 21132
rect -978 21110 -974 21132
rect -954 21110 -950 21132
rect -930 21110 -926 21132
rect -906 21110 -902 21132
rect -882 21110 -878 21132
rect -858 21110 -854 21132
rect -834 21110 -830 21132
rect -810 21110 -806 21132
rect -786 21110 -782 21132
rect -762 21110 -758 21132
rect -738 21110 -734 21132
rect -714 21110 -710 21132
rect -690 21110 -686 21132
rect -666 21110 -662 21132
rect -642 21110 -638 21132
rect -618 21110 -614 21132
rect -594 21110 -590 21132
rect -570 21110 -566 21132
rect -546 21110 -542 21132
rect -522 21110 -518 21132
rect -498 21110 -494 21132
rect -474 21110 -470 21132
rect -450 21110 -446 21132
rect -426 21110 -422 21132
rect -402 21110 -398 21132
rect -378 21110 -374 21132
rect -354 21110 -350 21132
rect -330 21110 -326 21132
rect -306 21110 -302 21132
rect -282 21110 -278 21132
rect -258 21110 -254 21132
rect -234 21110 -230 21132
rect -210 21110 -206 21132
rect -186 21110 -182 21132
rect -162 21110 -158 21132
rect -138 21110 -134 21132
rect -114 21110 -110 21132
rect -90 21110 -86 21132
rect -66 21110 -62 21132
rect -42 21110 -38 21132
rect -18 21110 -14 21132
rect 6 21110 10 21132
rect 30 21110 34 21132
rect 54 21110 58 21132
rect 78 21110 82 21132
rect 102 21110 106 21132
rect 126 21110 130 21132
rect 150 21110 154 21132
rect 174 21110 178 21132
rect 198 21110 202 21132
rect 222 21110 226 21132
rect 246 21110 250 21132
rect 270 21110 274 21132
rect 294 21110 298 21132
rect 318 21110 322 21132
rect 342 21110 346 21132
rect 366 21110 370 21132
rect 390 21110 394 21132
rect 414 21110 418 21132
rect 438 21110 442 21132
rect 462 21110 466 21132
rect 486 21110 490 21132
rect 510 21110 514 21132
rect 534 21110 538 21132
rect 558 21110 562 21132
rect 582 21110 586 21132
rect 606 21110 610 21132
rect 630 21110 634 21132
rect 654 21110 658 21132
rect 678 21110 682 21132
rect 702 21110 706 21132
rect 726 21110 730 21132
rect 750 21110 754 21132
rect 774 21110 778 21132
rect 787 21125 792 21132
rect 798 21125 802 21132
rect 797 21111 802 21125
rect 822 21110 826 21156
rect 846 21110 850 21156
rect 870 21110 874 21156
rect 894 21110 898 21156
rect 918 21110 922 21156
rect 942 21110 946 21156
rect 966 21110 970 21156
rect 990 21110 994 21156
rect 1014 21110 1018 21156
rect 1038 21110 1042 21156
rect 1062 21110 1066 21156
rect 1086 21110 1090 21156
rect 1110 21110 1114 21156
rect 1134 21110 1138 21156
rect 1158 21110 1162 21156
rect 1182 21110 1186 21156
rect 1206 21110 1210 21156
rect 1230 21110 1234 21156
rect 1254 21110 1258 21156
rect 1278 21131 1282 21156
rect 1302 21155 1306 21156
rect 1278 21110 1285 21131
rect 1302 21110 1309 21155
rect 1326 21110 1330 21156
rect 1350 21110 1354 21156
rect 1374 21110 1378 21156
rect 1398 21110 1402 21156
rect 1422 21110 1426 21156
rect 1446 21110 1450 21156
rect 1470 21110 1474 21156
rect 1477 21155 1491 21156
rect 1494 21131 1501 21179
rect 1494 21110 1498 21131
rect 1518 21110 1522 21180
rect 1542 21110 1546 21180
rect 1566 21110 1570 21180
rect 1590 21110 1594 21180
rect 1614 21110 1618 21180
rect 1638 21110 1642 21180
rect 1662 21110 1666 21180
rect 1686 21110 1690 21180
rect 1710 21110 1714 21180
rect 1734 21110 1738 21180
rect 1758 21110 1762 21180
rect 1782 21110 1786 21180
rect 1806 21110 1810 21180
rect 1830 21110 1834 21180
rect 1854 21111 1858 21180
rect 1843 21110 1877 21111
rect -2030 21108 1275 21110
rect -2371 21062 -2366 21108
rect -2348 21062 -2343 21108
rect -2325 21062 -2320 21108
rect -2317 21104 -2309 21108
rect -2060 21104 -2050 21108
rect -2060 21102 -2036 21104
rect -2060 21100 -2030 21102
rect -2292 21094 -2030 21100
rect -2092 21078 -2062 21080
rect -2094 21074 -2062 21078
rect -2000 21062 -1992 21108
rect -1844 21101 -1806 21108
rect -1663 21104 -1655 21108
rect -1844 21094 -1680 21100
rect -1854 21078 -1806 21080
rect -1854 21074 -1680 21078
rect -1642 21062 -1637 21108
rect -1619 21062 -1614 21108
rect -1530 21062 -1526 21108
rect -1506 21062 -1502 21108
rect -1482 21062 -1478 21108
rect -1458 21062 -1454 21108
rect -1434 21062 -1430 21108
rect -1410 21062 -1406 21108
rect -1386 21062 -1382 21108
rect -1362 21062 -1358 21108
rect -1338 21062 -1334 21108
rect -1314 21062 -1310 21108
rect -1290 21062 -1286 21108
rect -1266 21062 -1262 21108
rect -1242 21062 -1238 21108
rect -1218 21062 -1214 21108
rect -1194 21062 -1190 21108
rect -1170 21062 -1166 21108
rect -1146 21062 -1142 21108
rect -1122 21062 -1118 21108
rect -1098 21062 -1094 21108
rect -1074 21062 -1070 21108
rect -1050 21062 -1046 21108
rect -1026 21062 -1022 21108
rect -1002 21062 -998 21108
rect -978 21062 -974 21108
rect -954 21062 -950 21108
rect -930 21062 -926 21108
rect -906 21062 -902 21108
rect -882 21062 -878 21108
rect -858 21062 -854 21108
rect -834 21062 -830 21108
rect -810 21062 -806 21108
rect -786 21062 -782 21108
rect -762 21062 -758 21108
rect -738 21062 -734 21108
rect -714 21062 -710 21108
rect -690 21062 -686 21108
rect -666 21062 -662 21108
rect -642 21062 -638 21108
rect -618 21062 -614 21108
rect -594 21062 -590 21108
rect -570 21062 -566 21108
rect -546 21062 -542 21108
rect -522 21062 -518 21108
rect -498 21062 -494 21108
rect -474 21062 -470 21108
rect -450 21062 -446 21108
rect -426 21062 -422 21108
rect -402 21062 -398 21108
rect -378 21062 -374 21108
rect -354 21062 -350 21108
rect -330 21062 -326 21108
rect -306 21062 -302 21108
rect -282 21062 -278 21108
rect -258 21062 -254 21108
rect -234 21062 -230 21108
rect -210 21062 -206 21108
rect -186 21062 -182 21108
rect -162 21062 -158 21108
rect -138 21062 -134 21108
rect -114 21062 -110 21108
rect -90 21062 -86 21108
rect -66 21062 -62 21108
rect -42 21062 -38 21108
rect -18 21062 -14 21108
rect 6 21062 10 21108
rect 30 21062 34 21108
rect 54 21062 58 21108
rect 78 21062 82 21108
rect 102 21062 106 21108
rect 126 21062 130 21108
rect 150 21062 154 21108
rect 174 21062 178 21108
rect 198 21062 202 21108
rect 222 21062 226 21108
rect 246 21062 250 21108
rect 270 21062 274 21108
rect 294 21062 298 21108
rect 318 21062 322 21108
rect 342 21062 346 21108
rect 366 21062 370 21108
rect 390 21062 394 21108
rect 414 21062 418 21108
rect 438 21062 442 21108
rect 462 21062 466 21108
rect 486 21062 490 21108
rect 510 21062 514 21108
rect 534 21062 538 21108
rect 558 21062 562 21108
rect 582 21062 586 21108
rect 606 21062 610 21108
rect 630 21062 634 21108
rect 654 21062 658 21108
rect 678 21062 682 21108
rect 702 21062 706 21108
rect 726 21062 730 21108
rect 750 21062 754 21108
rect 774 21062 778 21108
rect 787 21077 792 21087
rect 797 21063 802 21077
rect 798 21062 802 21063
rect 822 21062 826 21108
rect 846 21062 850 21108
rect 870 21062 874 21108
rect 894 21062 898 21108
rect 918 21062 922 21108
rect 942 21062 946 21108
rect 966 21062 970 21108
rect 990 21062 994 21108
rect 1014 21062 1018 21108
rect 1038 21062 1042 21108
rect 1062 21062 1066 21108
rect 1086 21062 1090 21108
rect 1110 21062 1114 21108
rect 1134 21062 1138 21108
rect 1158 21062 1162 21108
rect 1182 21062 1186 21108
rect 1206 21062 1210 21108
rect 1230 21062 1234 21108
rect 1254 21062 1258 21108
rect 1261 21107 1275 21108
rect 1278 21108 1877 21110
rect 1278 21107 1299 21108
rect 1302 21107 1309 21108
rect 1278 21086 1285 21107
rect 1302 21086 1306 21107
rect 1326 21086 1330 21108
rect 1350 21086 1354 21108
rect 1374 21086 1378 21108
rect 1398 21086 1402 21108
rect 1422 21086 1426 21108
rect 1446 21086 1450 21108
rect 1470 21086 1474 21108
rect 1494 21086 1498 21108
rect 1518 21086 1522 21108
rect 1542 21086 1546 21108
rect 1566 21086 1570 21108
rect 1590 21086 1594 21108
rect 1614 21086 1618 21108
rect 1638 21086 1642 21108
rect 1662 21086 1666 21108
rect 1686 21086 1690 21108
rect 1710 21086 1714 21108
rect 1734 21086 1738 21108
rect 1758 21086 1762 21108
rect 1782 21086 1786 21108
rect 1806 21086 1810 21108
rect 1830 21086 1834 21108
rect 1843 21101 1848 21108
rect 1854 21101 1858 21108
rect 1853 21087 1858 21101
rect 1878 21086 1882 21180
rect 1902 21086 1906 21180
rect 1926 21086 1930 21180
rect 1950 21086 1954 21180
rect 1974 21086 1978 21180
rect 1998 21086 2002 21180
rect 2022 21086 2026 21180
rect 2046 21086 2050 21180
rect 2070 21086 2074 21180
rect 2094 21086 2098 21180
rect 2118 21086 2122 21180
rect 2142 21086 2146 21180
rect 2166 21086 2170 21180
rect 2190 21086 2194 21180
rect 2214 21086 2218 21180
rect 2238 21086 2242 21180
rect 2262 21086 2266 21180
rect 2286 21086 2290 21180
rect 2310 21086 2314 21180
rect 2334 21086 2338 21180
rect 2358 21086 2362 21180
rect 2382 21086 2386 21180
rect 2406 21086 2410 21180
rect 2430 21086 2434 21180
rect 2454 21086 2458 21180
rect 2478 21086 2482 21180
rect 2502 21086 2506 21180
rect 2526 21086 2530 21180
rect 2550 21086 2554 21180
rect 2574 21086 2578 21180
rect 2598 21086 2602 21180
rect 2622 21086 2626 21180
rect 2646 21086 2650 21180
rect 2670 21086 2674 21180
rect 2694 21086 2698 21180
rect 2718 21086 2722 21180
rect 2742 21086 2746 21180
rect 2766 21086 2770 21180
rect 2790 21086 2794 21180
rect 2814 21086 2818 21180
rect 2838 21086 2842 21180
rect 2862 21086 2866 21180
rect 2886 21086 2890 21180
rect 2910 21086 2914 21180
rect 2934 21086 2938 21180
rect 2958 21086 2962 21180
rect 2982 21086 2986 21180
rect 3006 21086 3010 21180
rect 3030 21086 3034 21180
rect 3054 21086 3058 21180
rect 3078 21086 3082 21180
rect 3102 21086 3106 21180
rect 3126 21086 3130 21180
rect 3150 21086 3154 21180
rect 3174 21086 3178 21180
rect 3198 21086 3202 21180
rect 3222 21086 3226 21180
rect 3246 21086 3250 21180
rect 3270 21086 3274 21180
rect 3294 21086 3298 21180
rect 3318 21086 3322 21180
rect 3342 21086 3346 21180
rect 3366 21086 3370 21180
rect 3390 21086 3394 21180
rect 3414 21086 3418 21180
rect 3438 21086 3442 21180
rect 3445 21179 3459 21180
rect 3462 21179 3469 21203
rect 3835 21193 3843 21197
rect 3829 21183 3835 21193
rect 3499 21180 3533 21183
rect 3811 21182 3845 21183
rect 3846 21182 3853 21204
rect 3859 21197 3864 21204
rect 3877 21203 3891 21204
rect 4549 21203 4563 21204
rect 3869 21183 3874 21197
rect 3883 21193 3891 21197
rect 4555 21193 4563 21197
rect 3877 21183 3883 21193
rect 4549 21183 4555 21193
rect 3859 21182 3893 21183
rect 3811 21180 3893 21182
rect 4531 21182 4565 21183
rect 4566 21182 4573 21204
rect 4579 21197 4584 21204
rect 4597 21203 4611 21204
rect 4789 21203 4803 21204
rect 4589 21183 4594 21197
rect 4603 21193 4611 21197
rect 4795 21193 4803 21197
rect 4597 21183 4603 21193
rect 4789 21183 4795 21193
rect 4579 21182 4613 21183
rect 4531 21180 4613 21182
rect 4771 21182 4805 21183
rect 4806 21182 4813 21204
rect 4819 21197 4824 21204
rect 4837 21203 4851 21204
rect 6589 21203 6603 21204
rect 4829 21183 4834 21197
rect 4843 21193 4851 21197
rect 6595 21193 6603 21197
rect 4837 21183 4843 21193
rect 6589 21183 6595 21193
rect 4819 21182 4853 21183
rect 4771 21180 4853 21182
rect 6571 21182 6605 21183
rect 6606 21182 6613 21204
rect 6726 21182 6730 21204
rect 6750 21182 6754 21204
rect 6774 21182 6778 21204
rect 6798 21183 6802 21204
rect 6811 21197 6816 21204
rect 6822 21197 6826 21204
rect 6821 21183 6826 21197
rect 6787 21182 6821 21183
rect 6571 21180 6821 21182
rect 3462 21086 3466 21179
rect 3486 21086 3490 21180
rect 3829 21179 3843 21180
rect 3835 21169 3843 21173
rect 3829 21159 3835 21169
rect 3499 21156 3533 21159
rect 3811 21158 3845 21159
rect 3846 21158 3853 21180
rect 3859 21173 3864 21180
rect 3877 21179 3891 21180
rect 4549 21179 4563 21180
rect 3869 21159 3874 21173
rect 3883 21169 3891 21173
rect 4555 21169 4563 21173
rect 3877 21159 3883 21169
rect 4549 21159 4555 21169
rect 3859 21158 3893 21159
rect 3811 21156 3893 21158
rect 4531 21158 4565 21159
rect 4566 21158 4573 21180
rect 4579 21173 4584 21180
rect 4597 21179 4611 21180
rect 4789 21179 4803 21180
rect 4589 21159 4594 21173
rect 4603 21169 4611 21173
rect 4795 21169 4803 21173
rect 4597 21159 4603 21169
rect 4789 21159 4795 21169
rect 4579 21158 4613 21159
rect 4531 21156 4613 21158
rect 4771 21158 4805 21159
rect 4806 21158 4813 21180
rect 4819 21173 4824 21180
rect 4837 21179 4851 21180
rect 6589 21179 6603 21180
rect 4829 21159 4834 21173
rect 4843 21169 4851 21173
rect 6595 21169 6603 21173
rect 4837 21159 4843 21169
rect 6589 21159 6595 21169
rect 4819 21158 4853 21159
rect 4771 21156 4853 21158
rect 6571 21158 6605 21159
rect 6606 21158 6613 21180
rect 6726 21158 6730 21180
rect 6750 21158 6754 21180
rect 6774 21159 6778 21180
rect 6787 21173 6792 21180
rect 6798 21173 6802 21180
rect 6797 21159 6802 21173
rect 6763 21158 6797 21159
rect 6571 21156 6797 21158
rect 3499 21149 3504 21156
rect 3829 21155 3843 21156
rect 3509 21135 3514 21149
rect 3523 21145 3531 21149
rect 3517 21135 3523 21145
rect 3534 21142 3541 21146
rect 3835 21145 3843 21149
rect 3829 21135 3835 21145
rect 3510 21086 3514 21135
rect 3811 21134 3845 21135
rect 3846 21134 3853 21156
rect 3859 21149 3864 21156
rect 3877 21155 3891 21156
rect 4549 21155 4563 21156
rect 3869 21135 3874 21149
rect 3883 21145 3891 21149
rect 4555 21145 4563 21149
rect 3877 21135 3883 21145
rect 4549 21135 4555 21145
rect 3859 21134 3893 21135
rect 3811 21132 3893 21134
rect 4531 21134 4565 21135
rect 4566 21134 4573 21156
rect 4579 21149 4584 21156
rect 4597 21155 4611 21156
rect 4789 21155 4803 21156
rect 4589 21135 4594 21149
rect 4603 21145 4611 21149
rect 4795 21145 4803 21149
rect 4597 21135 4603 21145
rect 4789 21135 4795 21145
rect 4579 21134 4613 21135
rect 4531 21132 4613 21134
rect 4771 21134 4805 21135
rect 4806 21134 4813 21156
rect 4819 21149 4824 21156
rect 4837 21155 4851 21156
rect 6589 21155 6603 21156
rect 4829 21135 4834 21149
rect 4843 21145 4851 21149
rect 6595 21145 6603 21149
rect 4837 21135 4843 21145
rect 6589 21135 6595 21145
rect 4819 21134 4853 21135
rect 4771 21132 4853 21134
rect 6571 21134 6605 21135
rect 6606 21134 6613 21156
rect 6726 21134 6730 21156
rect 6750 21135 6754 21156
rect 6763 21149 6768 21156
rect 6774 21149 6778 21156
rect 6773 21135 6778 21149
rect 6739 21134 6773 21135
rect 6571 21132 6773 21134
rect 3534 21118 3541 21132
rect 3829 21131 3843 21132
rect 3835 21121 3843 21125
rect 3829 21111 3835 21121
rect 3811 21110 3845 21111
rect 3846 21110 3853 21132
rect 3859 21125 3864 21132
rect 3877 21131 3891 21132
rect 4549 21131 4563 21132
rect 3869 21111 3874 21125
rect 3883 21121 3891 21125
rect 4555 21121 4563 21125
rect 3877 21111 3883 21121
rect 4549 21111 4555 21121
rect 3859 21110 3893 21111
rect 3811 21108 3893 21110
rect 4531 21110 4565 21111
rect 4566 21110 4573 21132
rect 4579 21125 4584 21132
rect 4597 21131 4611 21132
rect 4789 21131 4803 21132
rect 4589 21111 4594 21125
rect 4603 21121 4611 21125
rect 4795 21121 4803 21125
rect 4597 21111 4603 21121
rect 4789 21111 4795 21121
rect 4579 21110 4613 21111
rect 4531 21108 4613 21110
rect 4771 21110 4805 21111
rect 4806 21110 4813 21132
rect 4819 21125 4824 21132
rect 4837 21131 4851 21132
rect 6589 21131 6603 21132
rect 4829 21111 4834 21125
rect 4843 21121 4851 21125
rect 6595 21121 6603 21125
rect 4837 21111 4843 21121
rect 6589 21111 6595 21121
rect 4819 21110 4853 21111
rect 4771 21108 4853 21110
rect 6571 21110 6605 21111
rect 6606 21110 6613 21132
rect 6726 21111 6730 21132
rect 6739 21125 6744 21132
rect 6750 21125 6754 21132
rect 6749 21111 6754 21125
rect 6715 21110 6749 21111
rect 6571 21108 6749 21110
rect 3534 21094 3541 21108
rect 3829 21107 3843 21108
rect 3835 21097 3843 21101
rect 3829 21087 3835 21097
rect 1261 21084 3531 21086
rect 3595 21084 3629 21087
rect 3811 21086 3845 21087
rect 3846 21086 3853 21108
rect 3859 21101 3864 21108
rect 3877 21107 3891 21108
rect 4549 21107 4563 21108
rect 3869 21087 3874 21101
rect 3883 21097 3891 21101
rect 4555 21097 4563 21101
rect 3877 21087 3883 21097
rect 4549 21087 4555 21097
rect 3859 21086 3893 21087
rect 3811 21084 3893 21086
rect 4531 21086 4565 21087
rect 4566 21086 4573 21108
rect 4579 21101 4584 21108
rect 4597 21107 4611 21108
rect 4789 21107 4803 21108
rect 4589 21087 4594 21101
rect 4603 21097 4611 21101
rect 4795 21097 4803 21101
rect 4597 21087 4603 21097
rect 4789 21087 4795 21097
rect 4579 21086 4613 21087
rect 4531 21084 4613 21086
rect 4771 21086 4805 21087
rect 4806 21086 4813 21108
rect 4819 21101 4824 21108
rect 4837 21107 4851 21108
rect 6589 21107 6603 21108
rect 4829 21087 4834 21101
rect 4843 21097 4851 21101
rect 6595 21097 6603 21101
rect 4837 21087 4843 21097
rect 6589 21087 6595 21097
rect 4819 21086 4853 21087
rect 4771 21084 4853 21086
rect 6571 21086 6605 21087
rect 6606 21086 6613 21108
rect 6715 21101 6720 21108
rect 6726 21101 6730 21108
rect 6725 21087 6730 21101
rect 6667 21086 6701 21087
rect 6571 21084 6701 21086
rect 1261 21083 1275 21084
rect 1278 21083 1285 21084
rect 1278 21062 1282 21083
rect 1302 21062 1306 21084
rect 1326 21062 1330 21084
rect 1350 21062 1354 21084
rect 1374 21062 1378 21084
rect 1398 21062 1402 21084
rect 1422 21062 1426 21084
rect 1446 21062 1450 21084
rect 1470 21062 1474 21084
rect 1494 21062 1498 21084
rect 1518 21062 1522 21084
rect 1542 21062 1546 21084
rect 1566 21062 1570 21084
rect 1590 21062 1594 21084
rect 1614 21062 1618 21084
rect 1638 21062 1642 21084
rect 1662 21062 1666 21084
rect 1686 21062 1690 21084
rect 1710 21062 1714 21084
rect 1734 21062 1738 21084
rect 1758 21062 1762 21084
rect 1782 21062 1786 21084
rect 1806 21062 1810 21084
rect 1830 21062 1834 21084
rect 1843 21062 1877 21063
rect -2393 21060 1877 21062
rect -2371 21038 -2366 21060
rect -2348 21038 -2343 21060
rect -2325 21038 -2320 21060
rect -2072 21058 -2036 21059
rect -2072 21052 -2054 21058
rect -2309 21044 -2301 21052
rect -2317 21038 -2309 21044
rect -2092 21043 -2062 21048
rect -2000 21039 -1992 21060
rect -1938 21059 -1906 21060
rect -1920 21058 -1906 21059
rect -1806 21052 -1680 21058
rect -1854 21043 -1806 21048
rect -1655 21044 -1647 21052
rect -1982 21039 -1966 21040
rect -2000 21038 -1966 21039
rect -1846 21038 -1806 21041
rect -1663 21038 -1655 21044
rect -1642 21038 -1637 21060
rect -1619 21038 -1614 21060
rect -1530 21038 -1526 21060
rect -1506 21038 -1502 21060
rect -1482 21038 -1478 21060
rect -1458 21038 -1454 21060
rect -1434 21038 -1430 21060
rect -1410 21038 -1406 21060
rect -1386 21038 -1382 21060
rect -1362 21038 -1358 21060
rect -1338 21038 -1334 21060
rect -1314 21038 -1310 21060
rect -1290 21038 -1286 21060
rect -1266 21038 -1262 21060
rect -1242 21038 -1238 21060
rect -1218 21038 -1214 21060
rect -1194 21038 -1190 21060
rect -1170 21038 -1166 21060
rect -1146 21038 -1142 21060
rect -1122 21038 -1118 21060
rect -1098 21038 -1094 21060
rect -1074 21038 -1070 21060
rect -1050 21038 -1046 21060
rect -1026 21038 -1022 21060
rect -1002 21038 -998 21060
rect -978 21038 -974 21060
rect -954 21038 -950 21060
rect -930 21038 -926 21060
rect -906 21038 -902 21060
rect -882 21038 -878 21060
rect -858 21038 -854 21060
rect -834 21038 -830 21060
rect -810 21038 -806 21060
rect -786 21038 -782 21060
rect -762 21038 -758 21060
rect -738 21038 -734 21060
rect -714 21038 -710 21060
rect -690 21038 -686 21060
rect -666 21038 -662 21060
rect -642 21038 -638 21060
rect -618 21038 -614 21060
rect -594 21038 -590 21060
rect -570 21038 -566 21060
rect -546 21038 -542 21060
rect -522 21038 -518 21060
rect -498 21038 -494 21060
rect -474 21038 -470 21060
rect -450 21038 -446 21060
rect -426 21038 -422 21060
rect -402 21038 -398 21060
rect -378 21038 -374 21060
rect -354 21038 -350 21060
rect -330 21038 -326 21060
rect -306 21038 -302 21060
rect -282 21038 -278 21060
rect -258 21038 -254 21060
rect -234 21038 -230 21060
rect -210 21038 -206 21060
rect -186 21038 -182 21060
rect -162 21038 -158 21060
rect -138 21038 -134 21060
rect -114 21038 -110 21060
rect -90 21038 -86 21060
rect -66 21038 -62 21060
rect -42 21038 -38 21060
rect -18 21038 -14 21060
rect 6 21038 10 21060
rect 30 21038 34 21060
rect 54 21038 58 21060
rect 78 21038 82 21060
rect 102 21038 106 21060
rect 126 21038 130 21060
rect 150 21038 154 21060
rect 174 21038 178 21060
rect 198 21038 202 21060
rect 222 21038 226 21060
rect 246 21038 250 21060
rect 270 21038 274 21060
rect 294 21038 298 21060
rect 318 21038 322 21060
rect 342 21038 346 21060
rect 366 21038 370 21060
rect 390 21038 394 21060
rect 414 21038 418 21060
rect 438 21038 442 21060
rect 462 21038 466 21060
rect 486 21038 490 21060
rect 510 21038 514 21060
rect 534 21038 538 21060
rect 558 21038 562 21060
rect 582 21038 586 21060
rect 606 21038 610 21060
rect 630 21038 634 21060
rect 654 21038 658 21060
rect 678 21038 682 21060
rect 702 21038 706 21060
rect 726 21038 730 21060
rect 750 21038 754 21060
rect 774 21038 778 21060
rect 798 21038 802 21060
rect 822 21059 826 21060
rect -2393 21036 819 21038
rect -2371 21014 -2366 21036
rect -2348 21014 -2343 21036
rect -2325 21014 -2320 21036
rect -2000 21034 -1966 21036
rect -2309 21016 -2301 21024
rect -2062 21023 -2054 21030
rect -2092 21016 -2084 21023
rect -2062 21016 -2026 21018
rect -2317 21014 -2309 21016
rect -2062 21014 -2012 21016
rect -2000 21014 -1992 21034
rect -1982 21033 -1966 21034
rect -1846 21032 -1806 21036
rect -1846 21025 -1798 21030
rect -1806 21023 -1798 21025
rect -1854 21021 -1846 21023
rect -1854 21016 -1806 21021
rect -1655 21016 -1647 21024
rect -1864 21014 -1796 21015
rect -1663 21014 -1655 21016
rect -1642 21014 -1637 21036
rect -1619 21014 -1614 21036
rect -1530 21014 -1526 21036
rect -1506 21014 -1502 21036
rect -1482 21014 -1478 21036
rect -1458 21014 -1454 21036
rect -1434 21014 -1430 21036
rect -1410 21014 -1406 21036
rect -1386 21014 -1382 21036
rect -1362 21014 -1358 21036
rect -1338 21014 -1334 21036
rect -1314 21014 -1310 21036
rect -1290 21014 -1286 21036
rect -1266 21014 -1262 21036
rect -1242 21014 -1238 21036
rect -1218 21014 -1214 21036
rect -1194 21014 -1190 21036
rect -1170 21014 -1166 21036
rect -1146 21014 -1142 21036
rect -1122 21014 -1118 21036
rect -1098 21014 -1094 21036
rect -1074 21014 -1070 21036
rect -1050 21014 -1046 21036
rect -1026 21014 -1022 21036
rect -1002 21014 -998 21036
rect -978 21014 -974 21036
rect -954 21014 -950 21036
rect -930 21014 -926 21036
rect -906 21014 -902 21036
rect -882 21014 -878 21036
rect -858 21014 -854 21036
rect -834 21014 -830 21036
rect -810 21014 -806 21036
rect -786 21014 -782 21036
rect -762 21014 -758 21036
rect -738 21014 -734 21036
rect -714 21014 -710 21036
rect -690 21014 -686 21036
rect -666 21014 -662 21036
rect -642 21014 -638 21036
rect -618 21014 -614 21036
rect -594 21014 -590 21036
rect -570 21014 -566 21036
rect -546 21014 -542 21036
rect -522 21014 -518 21036
rect -498 21014 -494 21036
rect -474 21014 -470 21036
rect -450 21014 -446 21036
rect -426 21014 -422 21036
rect -402 21014 -398 21036
rect -378 21014 -374 21036
rect -354 21014 -350 21036
rect -330 21014 -326 21036
rect -306 21014 -302 21036
rect -282 21014 -278 21036
rect -258 21014 -254 21036
rect -234 21014 -230 21036
rect -210 21014 -206 21036
rect -186 21014 -182 21036
rect -162 21014 -158 21036
rect -138 21014 -134 21036
rect -114 21014 -110 21036
rect -90 21014 -86 21036
rect -66 21014 -62 21036
rect -42 21014 -38 21036
rect -18 21014 -14 21036
rect 6 21014 10 21036
rect 30 21014 34 21036
rect 54 21014 58 21036
rect 78 21014 82 21036
rect 102 21014 106 21036
rect 126 21014 130 21036
rect 150 21014 154 21036
rect 174 21014 178 21036
rect 198 21014 202 21036
rect 222 21014 226 21036
rect 246 21014 250 21036
rect 270 21014 274 21036
rect 294 21014 298 21036
rect 318 21014 322 21036
rect 342 21014 346 21036
rect 366 21014 370 21036
rect 390 21014 394 21036
rect 414 21014 418 21036
rect 438 21014 442 21036
rect 462 21014 466 21036
rect 486 21014 490 21036
rect 510 21014 514 21036
rect 534 21014 538 21036
rect 558 21014 562 21036
rect 582 21014 586 21036
rect 606 21014 610 21036
rect 630 21014 634 21036
rect 654 21014 658 21036
rect 678 21014 682 21036
rect 702 21015 706 21036
rect 691 21014 725 21015
rect -2393 21012 725 21014
rect -2371 20966 -2366 21012
rect -2348 20966 -2343 21012
rect -2325 20966 -2320 21012
rect -2317 21008 -2309 21012
rect -2062 21008 -2054 21012
rect -2154 21004 -2138 21006
rect -2057 21004 -2054 21008
rect -2292 20998 -2054 21004
rect -2052 20998 -2044 21008
rect -2092 20982 -2062 20984
rect -2094 20978 -2062 20982
rect -2000 20966 -1992 21012
rect -1846 21005 -1806 21012
rect -1663 21008 -1655 21012
rect -1846 20998 -1680 21004
rect -1854 20982 -1806 20984
rect -1854 20978 -1680 20982
rect -1926 20966 -1892 20969
rect -1642 20966 -1637 21012
rect -1619 20966 -1614 21012
rect -1530 20966 -1526 21012
rect -1506 20966 -1502 21012
rect -1482 20966 -1478 21012
rect -1458 20966 -1454 21012
rect -1434 20966 -1430 21012
rect -1410 20966 -1406 21012
rect -1386 20966 -1382 21012
rect -1362 20966 -1358 21012
rect -1338 20966 -1334 21012
rect -1314 20966 -1310 21012
rect -1290 20966 -1286 21012
rect -1266 20966 -1262 21012
rect -1242 20966 -1238 21012
rect -1218 20966 -1214 21012
rect -1194 20966 -1190 21012
rect -1170 20966 -1166 21012
rect -1146 20966 -1142 21012
rect -1122 20966 -1118 21012
rect -1098 20966 -1094 21012
rect -1074 20966 -1070 21012
rect -1050 20966 -1046 21012
rect -1026 20966 -1022 21012
rect -1002 20966 -998 21012
rect -978 20966 -974 21012
rect -954 20966 -950 21012
rect -930 20966 -926 21012
rect -906 20966 -902 21012
rect -882 20966 -878 21012
rect -858 20966 -854 21012
rect -834 20966 -830 21012
rect -810 20966 -806 21012
rect -786 20966 -782 21012
rect -762 20966 -758 21012
rect -738 20966 -734 21012
rect -714 20966 -710 21012
rect -690 20966 -686 21012
rect -666 20966 -662 21012
rect -642 20966 -638 21012
rect -618 20966 -614 21012
rect -594 20966 -590 21012
rect -570 20966 -566 21012
rect -546 20966 -542 21012
rect -522 20966 -518 21012
rect -498 20966 -494 21012
rect -474 20966 -470 21012
rect -450 20966 -446 21012
rect -426 20966 -422 21012
rect -402 20966 -398 21012
rect -378 20966 -374 21012
rect -354 20966 -350 21012
rect -330 20966 -326 21012
rect -306 20966 -302 21012
rect -282 20966 -278 21012
rect -258 20966 -254 21012
rect -234 20966 -230 21012
rect -210 20966 -206 21012
rect -186 20966 -182 21012
rect -162 20966 -158 21012
rect -138 20966 -134 21012
rect -114 20966 -110 21012
rect -90 20966 -86 21012
rect -66 20966 -62 21012
rect -42 20966 -38 21012
rect -18 20966 -14 21012
rect 6 20966 10 21012
rect 30 20966 34 21012
rect 54 20966 58 21012
rect 78 20966 82 21012
rect 102 20966 106 21012
rect 126 20966 130 21012
rect 150 20966 154 21012
rect 174 20966 178 21012
rect 198 20966 202 21012
rect 222 20966 226 21012
rect 246 20966 250 21012
rect 270 20966 274 21012
rect 294 20966 298 21012
rect 318 20966 322 21012
rect 342 20966 346 21012
rect 366 20966 370 21012
rect 390 20966 394 21012
rect 414 20966 418 21012
rect 438 20966 442 21012
rect 462 20966 466 21012
rect 486 20966 490 21012
rect 510 20966 514 21012
rect 534 20966 538 21012
rect 558 20966 562 21012
rect 582 20966 586 21012
rect 606 20966 610 21012
rect 630 20966 634 21012
rect 654 20966 658 21012
rect 678 20966 682 21012
rect 691 21005 696 21012
rect 702 21005 706 21012
rect 701 20991 706 21005
rect 691 20981 696 20991
rect 701 20967 706 20981
rect 702 20966 706 20967
rect 726 20966 730 21036
rect 750 20966 754 21036
rect 774 20966 778 21036
rect 798 20966 802 21036
rect 805 21035 819 21036
rect 822 21035 829 21059
rect 822 20990 829 21011
rect 846 20990 850 21060
rect 870 20990 874 21060
rect 894 20990 898 21060
rect 918 20990 922 21060
rect 942 20990 946 21060
rect 966 20990 970 21060
rect 990 20990 994 21060
rect 1014 20990 1018 21060
rect 1038 20990 1042 21060
rect 1062 20990 1066 21060
rect 1086 20990 1090 21060
rect 1099 21029 1104 21039
rect 1110 21029 1114 21060
rect 1109 21015 1114 21029
rect 1099 21014 1133 21015
rect 1134 21014 1138 21060
rect 1158 21014 1162 21060
rect 1182 21014 1186 21060
rect 1206 21014 1210 21060
rect 1230 21014 1234 21060
rect 1254 21014 1258 21060
rect 1278 21014 1282 21060
rect 1302 21014 1306 21060
rect 1326 21014 1330 21060
rect 1350 21014 1354 21060
rect 1374 21014 1378 21060
rect 1398 21014 1402 21060
rect 1422 21014 1426 21060
rect 1446 21014 1450 21060
rect 1470 21014 1474 21060
rect 1494 21014 1498 21060
rect 1518 21014 1522 21060
rect 1542 21014 1546 21060
rect 1566 21014 1570 21060
rect 1590 21014 1594 21060
rect 1614 21014 1618 21060
rect 1638 21014 1642 21060
rect 1662 21014 1666 21060
rect 1686 21014 1690 21060
rect 1710 21014 1714 21060
rect 1734 21014 1738 21060
rect 1758 21014 1762 21060
rect 1782 21014 1786 21060
rect 1806 21014 1810 21060
rect 1830 21014 1834 21060
rect 1843 21053 1848 21060
rect 1853 21039 1858 21053
rect 1854 21014 1858 21039
rect 1878 21035 1882 21084
rect 1099 21012 1875 21014
rect 1099 21005 1104 21012
rect 1109 20991 1114 21005
rect 1110 20990 1114 20991
rect 1134 20990 1138 21012
rect 1158 20990 1162 21012
rect 1182 20990 1186 21012
rect 1206 20990 1210 21012
rect 1230 20990 1234 21012
rect 1254 20990 1258 21012
rect 1278 20990 1282 21012
rect 1302 20990 1306 21012
rect 1326 20990 1330 21012
rect 1350 20990 1354 21012
rect 1374 20990 1378 21012
rect 1398 20990 1402 21012
rect 1422 20990 1426 21012
rect 1446 20990 1450 21012
rect 1470 20990 1474 21012
rect 1494 20990 1498 21012
rect 1518 20990 1522 21012
rect 1542 20990 1546 21012
rect 1566 20990 1570 21012
rect 1590 20990 1594 21012
rect 1614 20990 1618 21012
rect 1638 20990 1642 21012
rect 1662 20990 1666 21012
rect 1686 20990 1690 21012
rect 1710 20990 1714 21012
rect 1734 20990 1738 21012
rect 1758 20990 1762 21012
rect 1782 20990 1786 21012
rect 1806 20990 1810 21012
rect 1830 20990 1834 21012
rect 1854 20990 1858 21012
rect 1861 21011 1875 21012
rect 1878 21011 1885 21035
rect 1902 20990 1906 21084
rect 1926 20990 1930 21084
rect 1950 20990 1954 21084
rect 1974 20990 1978 21084
rect 1998 20990 2002 21084
rect 2022 20990 2026 21084
rect 2046 20990 2050 21084
rect 2070 20990 2074 21084
rect 2094 20990 2098 21084
rect 2118 20990 2122 21084
rect 2142 20990 2146 21084
rect 2166 20990 2170 21084
rect 2190 20990 2194 21084
rect 2214 20990 2218 21084
rect 2238 20990 2242 21084
rect 2262 20990 2266 21084
rect 2286 20990 2290 21084
rect 2310 20990 2314 21084
rect 2334 20990 2338 21084
rect 2358 20990 2362 21084
rect 2382 20990 2386 21084
rect 2406 20990 2410 21084
rect 2430 20990 2434 21084
rect 2454 20990 2458 21084
rect 2478 20990 2482 21084
rect 2502 20990 2506 21084
rect 2526 20990 2530 21084
rect 2550 20990 2554 21084
rect 2574 20990 2578 21084
rect 2598 20990 2602 21084
rect 2622 20990 2626 21084
rect 2646 20990 2650 21084
rect 2670 20990 2674 21084
rect 2694 20990 2698 21084
rect 2718 20990 2722 21084
rect 2742 20990 2746 21084
rect 2766 20990 2770 21084
rect 2790 20990 2794 21084
rect 2814 20990 2818 21084
rect 2838 20990 2842 21084
rect 2862 20990 2866 21084
rect 2886 20990 2890 21084
rect 2910 20990 2914 21084
rect 2934 20990 2938 21084
rect 2958 20990 2962 21084
rect 2982 20990 2986 21084
rect 3006 20990 3010 21084
rect 3030 20990 3034 21084
rect 3054 20990 3058 21084
rect 3078 20990 3082 21084
rect 3102 20990 3106 21084
rect 3126 20990 3130 21084
rect 3150 20990 3154 21084
rect 3174 20990 3178 21084
rect 3198 20990 3202 21084
rect 3222 20990 3226 21084
rect 3246 20990 3250 21084
rect 3270 20990 3274 21084
rect 3294 20990 3298 21084
rect 3318 20990 3322 21084
rect 3342 20990 3346 21084
rect 3366 20990 3370 21084
rect 3390 20990 3394 21084
rect 3414 20990 3418 21084
rect 3438 20990 3442 21084
rect 3462 20990 3466 21084
rect 3486 20990 3490 21084
rect 3510 20990 3514 21084
rect 3517 21083 3531 21084
rect 3534 21059 3541 21084
rect 3829 21083 3843 21084
rect 3835 21073 3843 21077
rect 3829 21063 3835 21073
rect 3811 21062 3845 21063
rect 3846 21062 3853 21084
rect 3859 21077 3864 21084
rect 3877 21083 3891 21084
rect 4549 21083 4563 21084
rect 3869 21063 3874 21077
rect 3883 21073 3891 21077
rect 4555 21073 4563 21077
rect 3877 21063 3883 21073
rect 4549 21063 4555 21073
rect 3859 21062 3893 21063
rect 3811 21060 3893 21062
rect 4531 21062 4565 21063
rect 4566 21062 4573 21084
rect 4579 21077 4584 21084
rect 4597 21083 4611 21084
rect 4789 21083 4803 21084
rect 4589 21063 4594 21077
rect 4603 21073 4611 21077
rect 4795 21073 4803 21077
rect 4597 21063 4603 21073
rect 4789 21063 4795 21073
rect 4579 21062 4613 21063
rect 4531 21060 4613 21062
rect 4771 21062 4805 21063
rect 4806 21062 4813 21084
rect 4819 21077 4824 21084
rect 4837 21083 4851 21084
rect 6589 21083 6603 21084
rect 4829 21063 4834 21077
rect 4843 21073 4851 21077
rect 6595 21073 6603 21077
rect 4837 21063 4843 21073
rect 6589 21063 6595 21073
rect 4819 21062 4853 21063
rect 4771 21060 4853 21062
rect 6571 21062 6605 21063
rect 6606 21062 6613 21084
rect 6667 21077 6672 21084
rect 6677 21063 6682 21077
rect 6619 21062 6653 21063
rect 6571 21060 6653 21062
rect 3534 20990 3538 21059
rect 3558 20990 3562 21060
rect 3829 21059 3843 21060
rect 3835 21049 3843 21053
rect 3829 21039 3835 21049
rect 3811 21038 3845 21039
rect 3846 21038 3853 21060
rect 3859 21053 3864 21060
rect 3877 21059 3891 21060
rect 4549 21059 4563 21060
rect 3869 21039 3874 21053
rect 3883 21049 3891 21053
rect 4555 21049 4563 21053
rect 3877 21039 3883 21049
rect 4549 21039 4555 21049
rect 3859 21038 3893 21039
rect 3811 21036 3893 21038
rect 4531 21038 4565 21039
rect 4566 21038 4573 21060
rect 4579 21053 4584 21060
rect 4597 21059 4611 21060
rect 4789 21059 4803 21060
rect 4589 21039 4594 21053
rect 4603 21049 4611 21053
rect 4795 21049 4803 21053
rect 4597 21039 4603 21049
rect 4789 21039 4795 21049
rect 4579 21038 4613 21039
rect 4531 21036 4613 21038
rect 4771 21038 4805 21039
rect 4806 21038 4813 21060
rect 4819 21053 4824 21060
rect 4837 21059 4851 21060
rect 6589 21059 6603 21060
rect 4829 21039 4834 21053
rect 4843 21049 4851 21053
rect 6595 21049 6603 21053
rect 4837 21039 4843 21049
rect 6589 21039 6595 21049
rect 4819 21038 4853 21039
rect 4771 21036 4853 21038
rect 3582 20990 3586 21036
rect 3829 21035 3843 21036
rect 3835 21025 3843 21029
rect 3829 21015 3835 21025
rect 3643 21012 3677 21015
rect 3811 21014 3845 21015
rect 3846 21014 3853 21036
rect 3859 21029 3864 21036
rect 3877 21035 3891 21036
rect 4549 21035 4563 21036
rect 3869 21015 3874 21029
rect 3883 21025 3891 21029
rect 4555 21025 4563 21029
rect 3877 21015 3883 21025
rect 4549 21015 4555 21025
rect 3859 21014 3893 21015
rect 3811 21012 3893 21014
rect 4531 21014 4565 21015
rect 4566 21014 4573 21036
rect 4579 21029 4584 21036
rect 4597 21035 4611 21036
rect 4789 21035 4803 21036
rect 4589 21015 4594 21029
rect 4603 21025 4611 21029
rect 4795 21025 4803 21029
rect 4597 21015 4603 21025
rect 4789 21015 4795 21025
rect 4579 21014 4613 21015
rect 4531 21012 4613 21014
rect 3606 20990 3610 21012
rect 3829 21011 3843 21012
rect 3630 20998 3637 21011
rect 3835 21001 3843 21005
rect 3829 20991 3835 21001
rect 805 20988 3627 20990
rect 3643 20988 3677 20991
rect 3811 20990 3845 20991
rect 3846 20990 3853 21012
rect 3859 21005 3864 21012
rect 3877 21011 3891 21012
rect 4549 21011 4563 21012
rect 3869 20991 3874 21005
rect 3883 21001 3891 21005
rect 4555 21001 4563 21005
rect 3877 20991 3883 21001
rect 4549 20991 4555 21001
rect 3859 20990 3893 20991
rect 3811 20988 3893 20990
rect 805 20987 819 20988
rect 822 20987 829 20988
rect 822 20966 826 20987
rect 846 20966 850 20988
rect 870 20966 874 20988
rect 894 20966 898 20988
rect 918 20966 922 20988
rect 942 20966 946 20988
rect 966 20966 970 20988
rect 990 20966 994 20988
rect 1014 20966 1018 20988
rect 1038 20966 1042 20988
rect 1062 20966 1066 20988
rect 1086 20966 1090 20988
rect 1110 20966 1114 20988
rect 1134 20966 1138 20988
rect 1158 20966 1162 20988
rect 1182 20966 1186 20988
rect 1206 20966 1210 20988
rect 1230 20966 1234 20988
rect 1254 20966 1258 20988
rect 1278 20966 1282 20988
rect 1302 20966 1306 20988
rect 1326 20966 1330 20988
rect 1350 20966 1354 20988
rect 1374 20966 1378 20988
rect 1398 20966 1402 20988
rect 1422 20966 1426 20988
rect 1446 20966 1450 20988
rect 1470 20966 1474 20988
rect 1494 20966 1498 20988
rect 1518 20966 1522 20988
rect 1542 20966 1546 20988
rect 1566 20966 1570 20988
rect 1590 20966 1594 20988
rect 1614 20966 1618 20988
rect 1638 20966 1642 20988
rect 1662 20966 1666 20988
rect 1686 20966 1690 20988
rect 1710 20966 1714 20988
rect 1734 20966 1738 20988
rect 1758 20966 1762 20988
rect 1782 20966 1786 20988
rect 1806 20966 1810 20988
rect 1830 20966 1834 20988
rect 1854 20966 1858 20988
rect -2393 20964 1875 20966
rect -2371 20942 -2366 20964
rect -2348 20942 -2343 20964
rect -2325 20942 -2320 20964
rect -2054 20963 -1906 20964
rect -2054 20962 -2036 20963
rect -2309 20948 -2301 20958
rect -2317 20942 -2309 20948
rect -2068 20947 -2038 20954
rect -2000 20946 -1992 20963
rect -1920 20962 -1906 20963
rect -1846 20956 -1794 20964
rect -1852 20949 -1804 20954
rect -1902 20947 -1804 20949
rect -1655 20948 -1647 20958
rect -2000 20944 -1975 20946
rect -1902 20945 -1852 20947
rect -2025 20942 -1975 20944
rect -1846 20942 -1804 20945
rect -1663 20942 -1655 20948
rect -1642 20942 -1637 20964
rect -1619 20942 -1614 20964
rect -1530 20942 -1526 20964
rect -1506 20942 -1502 20964
rect -1482 20942 -1478 20964
rect -1458 20942 -1454 20964
rect -1434 20942 -1430 20964
rect -1410 20942 -1406 20964
rect -1386 20942 -1382 20964
rect -1362 20942 -1358 20964
rect -1338 20942 -1334 20964
rect -1314 20942 -1310 20964
rect -1290 20942 -1286 20964
rect -1266 20942 -1262 20964
rect -1242 20942 -1238 20964
rect -1218 20942 -1214 20964
rect -1194 20942 -1190 20964
rect -1170 20942 -1166 20964
rect -1146 20942 -1142 20964
rect -1122 20942 -1118 20964
rect -1098 20942 -1094 20964
rect -1074 20942 -1070 20964
rect -1050 20942 -1046 20964
rect -1026 20942 -1022 20964
rect -1002 20942 -998 20964
rect -978 20942 -974 20964
rect -954 20942 -950 20964
rect -930 20942 -926 20964
rect -906 20942 -902 20964
rect -882 20942 -878 20964
rect -858 20942 -854 20964
rect -834 20942 -830 20964
rect -810 20942 -806 20964
rect -786 20942 -782 20964
rect -762 20942 -758 20964
rect -738 20942 -734 20964
rect -714 20942 -710 20964
rect -690 20942 -686 20964
rect -666 20942 -662 20964
rect -642 20942 -638 20964
rect -618 20942 -614 20964
rect -594 20942 -590 20964
rect -570 20942 -566 20964
rect -546 20942 -542 20964
rect -522 20942 -518 20964
rect -498 20942 -494 20964
rect -474 20942 -470 20964
rect -450 20942 -446 20964
rect -426 20942 -422 20964
rect -402 20942 -398 20964
rect -378 20942 -374 20964
rect -354 20942 -350 20964
rect -330 20942 -326 20964
rect -306 20942 -302 20964
rect -282 20942 -278 20964
rect -258 20942 -254 20964
rect -234 20942 -230 20964
rect -210 20942 -206 20964
rect -186 20942 -182 20964
rect -162 20942 -158 20964
rect -138 20942 -134 20964
rect -114 20942 -110 20964
rect -90 20942 -86 20964
rect -66 20942 -62 20964
rect -42 20942 -38 20964
rect -18 20942 -14 20964
rect 6 20942 10 20964
rect 30 20942 34 20964
rect 54 20942 58 20964
rect 78 20942 82 20964
rect 102 20942 106 20964
rect 126 20942 130 20964
rect 150 20942 154 20964
rect 174 20942 178 20964
rect 198 20942 202 20964
rect 222 20942 226 20964
rect 246 20942 250 20964
rect 270 20942 274 20964
rect 294 20942 298 20964
rect 318 20942 322 20964
rect 342 20942 346 20964
rect 366 20942 370 20964
rect 390 20942 394 20964
rect 414 20942 418 20964
rect 438 20942 442 20964
rect 462 20942 466 20964
rect 486 20942 490 20964
rect 510 20942 514 20964
rect 534 20942 538 20964
rect 558 20942 562 20964
rect 582 20942 586 20964
rect 606 20942 610 20964
rect 630 20942 634 20964
rect 654 20942 658 20964
rect 678 20942 682 20964
rect 702 20942 706 20964
rect 726 20942 730 20964
rect 750 20942 754 20964
rect 774 20942 778 20964
rect 798 20942 802 20964
rect 822 20942 826 20964
rect 846 20942 850 20964
rect 870 20942 874 20964
rect 894 20942 898 20964
rect 918 20942 922 20964
rect 942 20942 946 20964
rect 966 20942 970 20964
rect 990 20942 994 20964
rect 1014 20942 1018 20964
rect 1038 20942 1042 20964
rect 1062 20942 1066 20964
rect 1086 20942 1090 20964
rect 1110 20942 1114 20964
rect 1134 20963 1138 20964
rect -2393 20940 1131 20942
rect -2371 20918 -2366 20940
rect -2348 20918 -2343 20940
rect -2325 20918 -2320 20940
rect -2054 20939 -2038 20940
rect -2000 20939 -1966 20940
rect -1846 20939 -1804 20940
rect -2000 20938 -1975 20939
rect -2076 20930 -2054 20937
rect -2309 20920 -2301 20930
rect -2044 20927 -2038 20932
rect -2028 20930 -2001 20937
rect -2054 20920 -2038 20927
rect -2015 20929 -2001 20930
rect -2015 20920 -2014 20929
rect -2317 20918 -2309 20920
rect -2044 20918 -2028 20920
rect -2000 20918 -1992 20938
rect -1982 20937 -1975 20938
rect -1862 20937 -1798 20938
rect -1985 20930 -1796 20937
rect -1862 20929 -1798 20930
rect -1852 20920 -1804 20927
rect -1655 20920 -1647 20930
rect -1976 20918 -1940 20919
rect -1663 20918 -1655 20920
rect -1642 20918 -1637 20940
rect -1619 20918 -1614 20940
rect -1530 20918 -1526 20940
rect -1506 20918 -1502 20940
rect -1482 20918 -1478 20940
rect -1458 20918 -1454 20940
rect -1434 20918 -1430 20940
rect -1410 20918 -1406 20940
rect -1386 20918 -1382 20940
rect -1362 20918 -1358 20940
rect -1338 20918 -1334 20940
rect -1314 20918 -1310 20940
rect -1290 20918 -1286 20940
rect -1266 20918 -1262 20940
rect -1242 20918 -1238 20940
rect -1218 20918 -1214 20940
rect -1194 20918 -1190 20940
rect -1170 20918 -1166 20940
rect -1146 20918 -1142 20940
rect -1122 20918 -1118 20940
rect -1098 20918 -1094 20940
rect -1074 20918 -1070 20940
rect -1050 20918 -1046 20940
rect -1026 20918 -1022 20940
rect -1002 20918 -998 20940
rect -978 20918 -974 20940
rect -954 20918 -950 20940
rect -930 20918 -926 20940
rect -906 20918 -902 20940
rect -882 20918 -878 20940
rect -858 20918 -854 20940
rect -834 20918 -830 20940
rect -810 20918 -806 20940
rect -786 20918 -782 20940
rect -762 20918 -758 20940
rect -738 20918 -734 20940
rect -714 20918 -710 20940
rect -690 20918 -686 20940
rect -666 20918 -662 20940
rect -642 20918 -638 20940
rect -618 20918 -614 20940
rect -594 20918 -590 20940
rect -570 20918 -566 20940
rect -546 20918 -542 20940
rect -522 20918 -518 20940
rect -498 20918 -494 20940
rect -474 20918 -470 20940
rect -450 20918 -446 20940
rect -426 20918 -422 20940
rect -402 20918 -398 20940
rect -378 20918 -374 20940
rect -354 20918 -350 20940
rect -330 20918 -326 20940
rect -306 20918 -302 20940
rect -282 20918 -278 20940
rect -258 20918 -254 20940
rect -234 20918 -230 20940
rect -210 20918 -206 20940
rect -186 20918 -182 20940
rect -162 20918 -158 20940
rect -138 20918 -134 20940
rect -114 20918 -110 20940
rect -90 20918 -86 20940
rect -66 20918 -62 20940
rect -42 20918 -38 20940
rect -18 20918 -14 20940
rect 6 20918 10 20940
rect 30 20918 34 20940
rect 54 20918 58 20940
rect 78 20918 82 20940
rect 102 20918 106 20940
rect 126 20918 130 20940
rect 150 20918 154 20940
rect 174 20918 178 20940
rect 198 20918 202 20940
rect 222 20918 226 20940
rect 246 20918 250 20940
rect 270 20918 274 20940
rect 294 20918 298 20940
rect 318 20918 322 20940
rect 342 20918 346 20940
rect 366 20918 370 20940
rect 390 20918 394 20940
rect 414 20918 418 20940
rect 438 20918 442 20940
rect 462 20918 466 20940
rect 486 20918 490 20940
rect 510 20918 514 20940
rect 534 20918 538 20940
rect 558 20918 562 20940
rect 582 20918 586 20940
rect 606 20918 610 20940
rect 630 20918 634 20940
rect 654 20918 658 20940
rect 678 20918 682 20940
rect 702 20918 706 20940
rect 726 20939 730 20940
rect -2393 20916 723 20918
rect -2371 20846 -2366 20916
rect -2348 20846 -2343 20916
rect -2325 20882 -2320 20916
rect -2317 20914 -2309 20916
rect -2076 20903 -2054 20910
rect -2325 20874 -2317 20882
rect -2060 20876 -2030 20879
rect -2325 20846 -2320 20874
rect -2317 20866 -2309 20874
rect -2060 20863 -2038 20874
rect -2033 20867 -2030 20876
rect -2028 20872 -2027 20876
rect -2068 20858 -2038 20861
rect -2000 20846 -1992 20916
rect -1846 20912 -1804 20916
rect -1663 20914 -1655 20916
rect -1846 20902 -1794 20911
rect -1912 20891 -1884 20893
rect -1852 20885 -1804 20889
rect -1844 20876 -1796 20879
rect -1671 20874 -1663 20882
rect -1844 20863 -1804 20874
rect -1663 20866 -1655 20874
rect -1852 20858 -1680 20862
rect -1642 20846 -1637 20916
rect -1619 20846 -1614 20916
rect -1530 20846 -1526 20916
rect -1506 20846 -1502 20916
rect -1482 20846 -1478 20916
rect -1458 20846 -1454 20916
rect -1434 20846 -1430 20916
rect -1410 20846 -1406 20916
rect -1386 20846 -1382 20916
rect -1362 20846 -1358 20916
rect -1338 20846 -1334 20916
rect -1314 20846 -1310 20916
rect -1290 20846 -1286 20916
rect -1266 20846 -1262 20916
rect -1242 20846 -1238 20916
rect -1218 20846 -1214 20916
rect -1194 20846 -1190 20916
rect -1170 20846 -1166 20916
rect -1146 20846 -1142 20916
rect -1122 20846 -1118 20916
rect -1098 20846 -1094 20916
rect -1074 20846 -1070 20916
rect -1050 20846 -1046 20916
rect -1026 20846 -1022 20916
rect -1002 20846 -998 20916
rect -978 20846 -974 20916
rect -954 20846 -950 20916
rect -930 20846 -926 20916
rect -906 20846 -902 20916
rect -882 20846 -878 20916
rect -858 20846 -854 20916
rect -834 20846 -830 20916
rect -810 20846 -806 20916
rect -786 20846 -782 20916
rect -762 20846 -758 20916
rect -738 20846 -734 20916
rect -714 20846 -710 20916
rect -690 20846 -686 20916
rect -666 20846 -662 20916
rect -642 20846 -638 20916
rect -618 20846 -614 20916
rect -594 20846 -590 20916
rect -570 20846 -566 20916
rect -546 20846 -542 20916
rect -522 20846 -518 20916
rect -498 20846 -494 20916
rect -474 20846 -470 20916
rect -450 20846 -446 20916
rect -426 20846 -422 20916
rect -402 20846 -398 20916
rect -378 20846 -374 20916
rect -354 20846 -350 20916
rect -330 20846 -326 20916
rect -306 20846 -302 20916
rect -282 20846 -278 20916
rect -258 20846 -254 20916
rect -234 20846 -230 20916
rect -210 20846 -206 20916
rect -186 20846 -182 20916
rect -162 20846 -158 20916
rect -138 20846 -134 20916
rect -114 20846 -110 20916
rect -90 20846 -86 20916
rect -66 20846 -62 20916
rect -42 20846 -38 20916
rect -18 20846 -14 20916
rect 6 20846 10 20916
rect 30 20846 34 20916
rect 54 20846 58 20916
rect 78 20846 82 20916
rect 102 20846 106 20916
rect 126 20846 130 20916
rect 150 20846 154 20916
rect 174 20846 178 20916
rect 198 20846 202 20916
rect 222 20846 226 20916
rect 246 20846 250 20916
rect 270 20846 274 20916
rect 294 20846 298 20916
rect 318 20846 322 20916
rect 342 20846 346 20916
rect 366 20846 370 20916
rect 390 20846 394 20916
rect 414 20846 418 20916
rect 438 20846 442 20916
rect 462 20846 466 20916
rect 486 20846 490 20916
rect 510 20846 514 20916
rect 534 20846 538 20916
rect 558 20846 562 20916
rect 582 20846 586 20916
rect 606 20846 610 20916
rect 630 20846 634 20916
rect 654 20846 658 20916
rect 678 20846 682 20916
rect 702 20846 706 20916
rect 709 20915 723 20916
rect 726 20894 733 20939
rect 750 20894 754 20940
rect 774 20894 778 20940
rect 798 20894 802 20940
rect 822 20894 826 20940
rect 846 20894 850 20940
rect 870 20894 874 20940
rect 894 20894 898 20940
rect 918 20894 922 20940
rect 942 20894 946 20940
rect 966 20894 970 20940
rect 990 20894 994 20940
rect 1014 20894 1018 20940
rect 1038 20894 1042 20940
rect 1062 20894 1066 20940
rect 1086 20894 1090 20940
rect 1110 20894 1114 20940
rect 1117 20939 1131 20940
rect 1134 20918 1141 20963
rect 1158 20918 1162 20964
rect 1182 20918 1186 20964
rect 1206 20918 1210 20964
rect 1230 20918 1234 20964
rect 1254 20918 1258 20964
rect 1278 20918 1282 20964
rect 1302 20918 1306 20964
rect 1326 20918 1330 20964
rect 1350 20918 1354 20964
rect 1374 20918 1378 20964
rect 1398 20918 1402 20964
rect 1422 20918 1426 20964
rect 1446 20918 1450 20964
rect 1470 20918 1474 20964
rect 1494 20918 1498 20964
rect 1518 20918 1522 20964
rect 1542 20918 1546 20964
rect 1566 20918 1570 20964
rect 1590 20918 1594 20964
rect 1614 20918 1618 20964
rect 1638 20918 1642 20964
rect 1662 20918 1666 20964
rect 1686 20918 1690 20964
rect 1710 20918 1714 20964
rect 1734 20918 1738 20964
rect 1758 20918 1762 20964
rect 1782 20918 1786 20964
rect 1806 20918 1810 20964
rect 1830 20918 1834 20964
rect 1854 20918 1858 20964
rect 1861 20963 1875 20964
rect 1878 20963 1885 20987
rect 1878 20918 1882 20963
rect 1902 20918 1906 20988
rect 1926 20918 1930 20988
rect 1950 20918 1954 20988
rect 1974 20918 1978 20988
rect 1998 20918 2002 20988
rect 2022 20918 2026 20988
rect 2046 20918 2050 20988
rect 2070 20918 2074 20988
rect 2094 20918 2098 20988
rect 2118 20918 2122 20988
rect 2142 20918 2146 20988
rect 2166 20918 2170 20988
rect 2190 20918 2194 20988
rect 2214 20918 2218 20988
rect 2238 20918 2242 20988
rect 2262 20918 2266 20988
rect 2286 20918 2290 20988
rect 2310 20918 2314 20988
rect 2334 20918 2338 20988
rect 2358 20918 2362 20988
rect 2382 20918 2386 20988
rect 2406 20918 2410 20988
rect 2430 20918 2434 20988
rect 2454 20918 2458 20988
rect 2478 20918 2482 20988
rect 2502 20918 2506 20988
rect 2526 20918 2530 20988
rect 2550 20918 2554 20988
rect 2574 20918 2578 20988
rect 2598 20918 2602 20988
rect 2622 20918 2626 20988
rect 2646 20918 2650 20988
rect 2670 20918 2674 20988
rect 2694 20918 2698 20988
rect 2718 20918 2722 20988
rect 2742 20918 2746 20988
rect 2766 20918 2770 20988
rect 2790 20918 2794 20988
rect 2814 20919 2818 20988
rect 2803 20918 2837 20919
rect 1117 20916 2837 20918
rect 1117 20915 1131 20916
rect 1134 20915 1141 20916
rect 1134 20894 1138 20915
rect 1158 20894 1162 20916
rect 1182 20894 1186 20916
rect 1206 20894 1210 20916
rect 1230 20894 1234 20916
rect 1254 20894 1258 20916
rect 1278 20894 1282 20916
rect 1302 20894 1306 20916
rect 1326 20894 1330 20916
rect 1350 20894 1354 20916
rect 1374 20894 1378 20916
rect 1398 20894 1402 20916
rect 1422 20894 1426 20916
rect 1446 20894 1450 20916
rect 1470 20894 1474 20916
rect 1494 20894 1498 20916
rect 1518 20894 1522 20916
rect 1542 20894 1546 20916
rect 1566 20894 1570 20916
rect 1590 20894 1594 20916
rect 1614 20894 1618 20916
rect 1638 20894 1642 20916
rect 1662 20894 1666 20916
rect 1686 20894 1690 20916
rect 1710 20894 1714 20916
rect 1734 20895 1738 20916
rect 1723 20894 1757 20895
rect 709 20892 1757 20894
rect 709 20891 723 20892
rect 726 20891 733 20892
rect 726 20846 730 20891
rect 750 20846 754 20892
rect 774 20846 778 20892
rect 798 20846 802 20892
rect 822 20846 826 20892
rect 846 20846 850 20892
rect 870 20846 874 20892
rect 894 20846 898 20892
rect 918 20846 922 20892
rect 942 20846 946 20892
rect 966 20846 970 20892
rect 990 20846 994 20892
rect 1014 20846 1018 20892
rect 1038 20846 1042 20892
rect 1062 20846 1066 20892
rect 1086 20846 1090 20892
rect 1110 20846 1114 20892
rect 1134 20846 1138 20892
rect 1158 20846 1162 20892
rect 1182 20846 1186 20892
rect 1206 20846 1210 20892
rect 1230 20846 1234 20892
rect 1254 20846 1258 20892
rect 1278 20846 1282 20892
rect 1302 20846 1306 20892
rect 1326 20846 1330 20892
rect 1350 20846 1354 20892
rect 1374 20846 1378 20892
rect 1398 20846 1402 20892
rect 1422 20846 1426 20892
rect 1446 20846 1450 20892
rect 1470 20846 1474 20892
rect 1494 20846 1498 20892
rect 1518 20846 1522 20892
rect 1542 20846 1546 20892
rect 1566 20846 1570 20892
rect 1590 20846 1594 20892
rect 1614 20846 1618 20892
rect 1638 20846 1642 20892
rect 1662 20846 1666 20892
rect 1686 20846 1690 20892
rect 1710 20846 1714 20892
rect 1723 20885 1728 20892
rect 1734 20885 1738 20892
rect 1733 20871 1738 20885
rect 1734 20846 1738 20871
rect 1758 20846 1762 20916
rect 1782 20846 1786 20916
rect 1806 20846 1810 20916
rect 1830 20846 1834 20916
rect 1854 20846 1858 20916
rect 1878 20846 1882 20916
rect 1902 20846 1906 20916
rect 1926 20846 1930 20916
rect 1950 20846 1954 20916
rect 1974 20846 1978 20916
rect 1998 20846 2002 20916
rect 2022 20846 2026 20916
rect 2046 20846 2050 20916
rect 2070 20846 2074 20916
rect 2094 20846 2098 20916
rect 2118 20846 2122 20916
rect 2142 20846 2146 20916
rect 2166 20846 2170 20916
rect 2190 20846 2194 20916
rect 2214 20846 2218 20916
rect 2238 20846 2242 20916
rect 2262 20846 2266 20916
rect 2286 20846 2290 20916
rect 2310 20846 2314 20916
rect 2334 20846 2338 20916
rect 2358 20846 2362 20916
rect 2382 20846 2386 20916
rect 2406 20846 2410 20916
rect 2430 20846 2434 20916
rect 2454 20846 2458 20916
rect 2478 20846 2482 20916
rect 2502 20846 2506 20916
rect 2526 20846 2530 20916
rect 2550 20846 2554 20916
rect 2574 20846 2578 20916
rect 2598 20846 2602 20916
rect 2622 20846 2626 20916
rect 2646 20846 2650 20916
rect 2670 20846 2674 20916
rect 2694 20846 2698 20916
rect 2718 20846 2722 20916
rect 2742 20846 2746 20916
rect 2766 20846 2770 20916
rect 2790 20846 2794 20916
rect 2803 20909 2808 20916
rect 2814 20909 2818 20916
rect 2813 20895 2818 20909
rect 2814 20846 2818 20895
rect 2838 20846 2842 20988
rect 2862 20846 2866 20988
rect 2886 20846 2890 20988
rect 2910 20846 2914 20988
rect 2934 20846 2938 20988
rect 2958 20846 2962 20988
rect 2982 20846 2986 20988
rect 3006 20846 3010 20988
rect 3030 20846 3034 20988
rect 3054 20846 3058 20988
rect 3078 20846 3082 20988
rect 3102 20846 3106 20988
rect 3126 20846 3130 20988
rect 3150 20846 3154 20988
rect 3174 20846 3178 20988
rect 3198 20846 3202 20988
rect 3222 20846 3226 20988
rect 3246 20846 3250 20988
rect 3259 20933 3264 20943
rect 3270 20933 3274 20988
rect 3269 20919 3274 20933
rect 3270 20846 3274 20919
rect 3294 20867 3298 20988
rect -2393 20844 3291 20846
rect -2371 20822 -2366 20844
rect -2348 20822 -2343 20844
rect -2325 20822 -2320 20844
rect -2309 20826 -2301 20836
rect -2068 20827 -2062 20832
rect -2317 20822 -2309 20826
rect -2060 20822 -2050 20827
rect -2000 20822 -1992 20844
rect -1806 20836 -1680 20842
rect -1854 20827 -1806 20832
rect -1655 20826 -1647 20836
rect -1972 20822 -1964 20823
rect -1958 20822 -1942 20824
rect -1844 20822 -1806 20825
rect -1663 20822 -1655 20826
rect -1642 20822 -1637 20844
rect -1619 20822 -1614 20844
rect -1530 20822 -1526 20844
rect -1506 20822 -1502 20844
rect -1482 20822 -1478 20844
rect -1458 20822 -1454 20844
rect -1434 20822 -1430 20844
rect -1410 20822 -1406 20844
rect -1386 20822 -1382 20844
rect -1362 20822 -1358 20844
rect -1338 20822 -1334 20844
rect -1314 20822 -1310 20844
rect -1290 20822 -1286 20844
rect -1266 20822 -1262 20844
rect -1242 20822 -1238 20844
rect -1218 20822 -1214 20844
rect -1194 20822 -1190 20844
rect -1170 20822 -1166 20844
rect -1146 20822 -1142 20844
rect -1122 20822 -1118 20844
rect -1098 20822 -1094 20844
rect -1074 20822 -1070 20844
rect -1050 20822 -1046 20844
rect -1026 20822 -1022 20844
rect -1002 20822 -998 20844
rect -978 20822 -974 20844
rect -954 20822 -950 20844
rect -930 20822 -926 20844
rect -906 20822 -902 20844
rect -882 20822 -878 20844
rect -858 20822 -854 20844
rect -834 20822 -830 20844
rect -810 20822 -806 20844
rect -786 20822 -782 20844
rect -762 20822 -758 20844
rect -738 20822 -734 20844
rect -714 20822 -710 20844
rect -690 20822 -686 20844
rect -666 20822 -662 20844
rect -642 20822 -638 20844
rect -618 20822 -614 20844
rect -594 20822 -590 20844
rect -570 20822 -566 20844
rect -546 20822 -542 20844
rect -522 20822 -518 20844
rect -498 20822 -494 20844
rect -474 20822 -470 20844
rect -450 20822 -446 20844
rect -426 20822 -422 20844
rect -402 20822 -398 20844
rect -378 20822 -374 20844
rect -354 20822 -350 20844
rect -330 20822 -326 20844
rect -306 20822 -302 20844
rect -282 20822 -278 20844
rect -258 20822 -254 20844
rect -234 20822 -230 20844
rect -210 20822 -206 20844
rect -186 20822 -182 20844
rect -162 20822 -158 20844
rect -138 20822 -134 20844
rect -114 20822 -110 20844
rect -90 20822 -86 20844
rect -66 20822 -62 20844
rect -42 20822 -38 20844
rect -18 20822 -14 20844
rect 6 20822 10 20844
rect 30 20822 34 20844
rect 54 20822 58 20844
rect 78 20822 82 20844
rect 102 20822 106 20844
rect 126 20822 130 20844
rect 150 20822 154 20844
rect 174 20822 178 20844
rect 198 20822 202 20844
rect 222 20822 226 20844
rect 246 20822 250 20844
rect 270 20823 274 20844
rect 259 20822 293 20823
rect -2393 20820 293 20822
rect -2371 20798 -2366 20820
rect -2348 20798 -2343 20820
rect -2325 20798 -2320 20820
rect -2060 20814 -2050 20820
rect -2309 20798 -2301 20808
rect -2060 20807 -2030 20814
rect -2000 20810 -1992 20820
rect -1972 20818 -1942 20820
rect -1958 20817 -1942 20818
rect -1844 20816 -1806 20820
rect -2068 20800 -2062 20807
rect -2062 20798 -2036 20800
rect -2393 20796 -2036 20798
rect -2030 20798 -2012 20800
rect -2004 20798 -1990 20810
rect -1844 20809 -1798 20814
rect -1806 20807 -1798 20809
rect -1854 20805 -1844 20807
rect -1854 20800 -1806 20805
rect -1864 20798 -1796 20799
rect -1655 20798 -1647 20808
rect -1642 20798 -1637 20820
rect -1619 20798 -1614 20820
rect -1530 20798 -1526 20820
rect -1506 20798 -1502 20820
rect -1482 20798 -1478 20820
rect -1458 20798 -1454 20820
rect -1434 20798 -1430 20820
rect -1410 20798 -1406 20820
rect -1386 20798 -1382 20820
rect -1362 20798 -1358 20820
rect -1338 20798 -1334 20820
rect -1314 20798 -1310 20820
rect -1290 20798 -1286 20820
rect -1266 20798 -1262 20820
rect -1242 20798 -1238 20820
rect -1218 20798 -1214 20820
rect -1194 20798 -1190 20820
rect -1170 20798 -1166 20820
rect -1146 20798 -1142 20820
rect -1122 20798 -1118 20820
rect -1098 20798 -1094 20820
rect -1074 20798 -1070 20820
rect -1050 20798 -1046 20820
rect -1026 20798 -1022 20820
rect -1002 20798 -998 20820
rect -978 20798 -974 20820
rect -954 20798 -950 20820
rect -930 20798 -926 20820
rect -906 20798 -902 20820
rect -882 20798 -878 20820
rect -858 20798 -854 20820
rect -834 20798 -830 20820
rect -810 20798 -806 20820
rect -786 20798 -782 20820
rect -762 20798 -758 20820
rect -738 20798 -734 20820
rect -714 20798 -710 20820
rect -690 20798 -686 20820
rect -666 20798 -662 20820
rect -642 20798 -638 20820
rect -618 20798 -614 20820
rect -594 20798 -590 20820
rect -570 20798 -566 20820
rect -546 20798 -542 20820
rect -522 20798 -518 20820
rect -498 20798 -494 20820
rect -474 20798 -470 20820
rect -450 20798 -446 20820
rect -426 20798 -422 20820
rect -402 20798 -398 20820
rect -378 20798 -374 20820
rect -354 20798 -350 20820
rect -330 20798 -326 20820
rect -306 20798 -302 20820
rect -282 20798 -278 20820
rect -258 20798 -254 20820
rect -234 20798 -230 20820
rect -210 20798 -206 20820
rect -186 20798 -182 20820
rect -162 20798 -158 20820
rect -138 20798 -134 20820
rect -114 20798 -110 20820
rect -90 20798 -86 20820
rect -66 20798 -62 20820
rect -42 20798 -38 20820
rect -18 20798 -14 20820
rect 6 20798 10 20820
rect 30 20798 34 20820
rect 54 20798 58 20820
rect 78 20798 82 20820
rect 102 20798 106 20820
rect 126 20798 130 20820
rect 150 20798 154 20820
rect 174 20798 178 20820
rect 198 20798 202 20820
rect 222 20798 226 20820
rect 246 20798 250 20820
rect 259 20813 264 20820
rect 270 20813 274 20820
rect 269 20799 274 20813
rect 259 20798 293 20799
rect 294 20798 298 20844
rect 318 20798 322 20844
rect 342 20798 346 20844
rect 366 20798 370 20844
rect 390 20798 394 20844
rect 414 20798 418 20844
rect 438 20798 442 20844
rect 462 20798 466 20844
rect 486 20798 490 20844
rect 510 20798 514 20844
rect 534 20798 538 20844
rect 558 20798 562 20844
rect 582 20798 586 20844
rect 606 20798 610 20844
rect 630 20798 634 20844
rect 654 20798 658 20844
rect 678 20798 682 20844
rect 702 20798 706 20844
rect 726 20798 730 20844
rect 750 20798 754 20844
rect 774 20798 778 20844
rect 798 20798 802 20844
rect 822 20798 826 20844
rect 846 20798 850 20844
rect 870 20798 874 20844
rect 894 20798 898 20844
rect 918 20798 922 20844
rect 942 20798 946 20844
rect 966 20798 970 20844
rect 990 20798 994 20844
rect 1014 20798 1018 20844
rect 1038 20798 1042 20844
rect 1062 20798 1066 20844
rect 1086 20798 1090 20844
rect 1110 20798 1114 20844
rect 1134 20799 1138 20844
rect 1123 20798 1157 20799
rect -2030 20796 1157 20798
rect -2371 20750 -2366 20796
rect -2348 20750 -2343 20796
rect -2325 20750 -2320 20796
rect -2317 20792 -2309 20796
rect -2060 20792 -2050 20796
rect -2060 20790 -2036 20792
rect -2060 20788 -2030 20790
rect -2292 20782 -2030 20788
rect -2092 20766 -2062 20768
rect -2094 20762 -2062 20766
rect -2000 20750 -1992 20796
rect -1844 20789 -1806 20796
rect -1663 20792 -1655 20796
rect -1844 20782 -1680 20788
rect -1854 20766 -1806 20768
rect -1854 20762 -1680 20766
rect -1926 20750 -1892 20753
rect -1642 20750 -1637 20796
rect -1619 20750 -1614 20796
rect -1530 20750 -1526 20796
rect -1506 20750 -1502 20796
rect -1482 20750 -1478 20796
rect -1458 20750 -1454 20796
rect -1434 20750 -1430 20796
rect -1410 20750 -1406 20796
rect -1386 20750 -1382 20796
rect -1362 20750 -1358 20796
rect -1338 20750 -1334 20796
rect -1314 20750 -1310 20796
rect -1290 20750 -1286 20796
rect -1266 20750 -1262 20796
rect -1242 20750 -1238 20796
rect -1218 20750 -1214 20796
rect -1194 20750 -1190 20796
rect -1170 20750 -1166 20796
rect -1146 20750 -1142 20796
rect -1122 20750 -1118 20796
rect -1098 20750 -1094 20796
rect -1074 20750 -1070 20796
rect -1050 20750 -1046 20796
rect -1026 20750 -1022 20796
rect -1002 20750 -998 20796
rect -978 20750 -974 20796
rect -954 20750 -950 20796
rect -930 20750 -926 20796
rect -906 20750 -902 20796
rect -882 20750 -878 20796
rect -858 20750 -854 20796
rect -834 20750 -830 20796
rect -810 20750 -806 20796
rect -786 20750 -782 20796
rect -762 20750 -758 20796
rect -738 20750 -734 20796
rect -714 20750 -710 20796
rect -690 20750 -686 20796
rect -666 20750 -662 20796
rect -642 20750 -638 20796
rect -618 20750 -614 20796
rect -594 20750 -590 20796
rect -570 20750 -566 20796
rect -546 20750 -542 20796
rect -522 20750 -518 20796
rect -498 20750 -494 20796
rect -474 20750 -470 20796
rect -450 20750 -446 20796
rect -426 20750 -422 20796
rect -402 20750 -398 20796
rect -378 20750 -374 20796
rect -354 20750 -350 20796
rect -330 20750 -326 20796
rect -306 20750 -302 20796
rect -282 20750 -278 20796
rect -258 20750 -254 20796
rect -234 20750 -230 20796
rect -210 20750 -206 20796
rect -186 20750 -182 20796
rect -162 20750 -158 20796
rect -138 20750 -134 20796
rect -114 20750 -110 20796
rect -90 20750 -86 20796
rect -66 20750 -62 20796
rect -42 20750 -38 20796
rect -18 20750 -14 20796
rect 6 20750 10 20796
rect 30 20750 34 20796
rect 54 20750 58 20796
rect 78 20750 82 20796
rect 102 20750 106 20796
rect 126 20750 130 20796
rect 150 20750 154 20796
rect 174 20750 178 20796
rect 198 20750 202 20796
rect 222 20750 226 20796
rect 246 20750 250 20796
rect 259 20789 264 20796
rect 269 20775 274 20789
rect 270 20750 274 20775
rect 294 20750 298 20796
rect 318 20750 322 20796
rect 342 20750 346 20796
rect 366 20750 370 20796
rect 390 20750 394 20796
rect 414 20750 418 20796
rect 438 20750 442 20796
rect 462 20750 466 20796
rect 486 20750 490 20796
rect 510 20750 514 20796
rect 534 20750 538 20796
rect 558 20750 562 20796
rect 582 20750 586 20796
rect 606 20750 610 20796
rect 630 20750 634 20796
rect 654 20750 658 20796
rect 678 20750 682 20796
rect 702 20750 706 20796
rect 726 20750 730 20796
rect 750 20750 754 20796
rect 774 20750 778 20796
rect 798 20750 802 20796
rect 822 20750 826 20796
rect 846 20750 850 20796
rect 870 20750 874 20796
rect 894 20750 898 20796
rect 918 20750 922 20796
rect 942 20750 946 20796
rect 966 20750 970 20796
rect 990 20750 994 20796
rect 1014 20750 1018 20796
rect 1038 20750 1042 20796
rect 1062 20750 1066 20796
rect 1086 20750 1090 20796
rect 1110 20750 1114 20796
rect 1123 20789 1128 20796
rect 1134 20789 1138 20796
rect 1133 20775 1138 20789
rect 1123 20765 1128 20775
rect 1133 20751 1138 20765
rect 1134 20750 1138 20751
rect 1158 20750 1162 20844
rect 1182 20750 1186 20844
rect 1206 20750 1210 20844
rect 1230 20750 1234 20844
rect 1254 20750 1258 20844
rect 1278 20750 1282 20844
rect 1302 20750 1306 20844
rect 1326 20750 1330 20844
rect 1350 20750 1354 20844
rect 1374 20750 1378 20844
rect 1398 20750 1402 20844
rect 1422 20750 1426 20844
rect 1446 20750 1450 20844
rect 1470 20750 1474 20844
rect 1494 20750 1498 20844
rect 1518 20750 1522 20844
rect 1542 20750 1546 20844
rect 1566 20750 1570 20844
rect 1590 20750 1594 20844
rect 1614 20750 1618 20844
rect 1638 20750 1642 20844
rect 1662 20750 1666 20844
rect 1686 20750 1690 20844
rect 1710 20750 1714 20844
rect 1734 20750 1738 20844
rect 1758 20819 1762 20844
rect 1758 20795 1765 20819
rect 1758 20750 1762 20795
rect 1782 20750 1786 20844
rect 1806 20750 1810 20844
rect 1830 20750 1834 20844
rect 1854 20750 1858 20844
rect 1878 20750 1882 20844
rect 1902 20750 1906 20844
rect 1926 20750 1930 20844
rect 1950 20750 1954 20844
rect 1974 20750 1978 20844
rect 1998 20750 2002 20844
rect 2022 20750 2026 20844
rect 2046 20750 2050 20844
rect 2070 20750 2074 20844
rect 2094 20750 2098 20844
rect 2118 20750 2122 20844
rect 2142 20750 2146 20844
rect 2166 20750 2170 20844
rect 2190 20750 2194 20844
rect 2214 20750 2218 20844
rect 2238 20750 2242 20844
rect 2262 20750 2266 20844
rect 2286 20750 2290 20844
rect 2310 20750 2314 20844
rect 2334 20750 2338 20844
rect 2358 20750 2362 20844
rect 2382 20750 2386 20844
rect 2406 20750 2410 20844
rect 2430 20750 2434 20844
rect 2454 20750 2458 20844
rect 2478 20750 2482 20844
rect 2502 20750 2506 20844
rect 2526 20750 2530 20844
rect 2550 20750 2554 20844
rect 2574 20750 2578 20844
rect 2598 20750 2602 20844
rect 2622 20750 2626 20844
rect 2646 20750 2650 20844
rect 2670 20750 2674 20844
rect 2694 20750 2698 20844
rect 2718 20750 2722 20844
rect 2742 20750 2746 20844
rect 2766 20750 2770 20844
rect 2790 20750 2794 20844
rect 2814 20750 2818 20844
rect 2838 20843 2842 20844
rect 2838 20819 2845 20843
rect 2838 20750 2842 20819
rect 2862 20750 2866 20844
rect 2886 20750 2890 20844
rect 2910 20750 2914 20844
rect 2934 20750 2938 20844
rect 2958 20750 2962 20844
rect 2982 20750 2986 20844
rect 3006 20750 3010 20844
rect 3030 20750 3034 20844
rect 3054 20750 3058 20844
rect 3078 20750 3082 20844
rect 3102 20750 3106 20844
rect 3126 20750 3130 20844
rect 3150 20750 3154 20844
rect 3174 20750 3178 20844
rect 3198 20750 3202 20844
rect 3222 20750 3226 20844
rect 3246 20750 3250 20844
rect 3270 20750 3274 20844
rect 3277 20843 3291 20844
rect 3294 20843 3301 20867
rect 3294 20750 3298 20843
rect 3318 20750 3322 20988
rect 3342 20750 3346 20988
rect 3366 20750 3370 20988
rect 3390 20750 3394 20988
rect 3414 20750 3418 20988
rect 3438 20750 3442 20988
rect 3462 20750 3466 20988
rect 3486 20750 3490 20988
rect 3510 20750 3514 20988
rect 3534 20750 3538 20988
rect 3558 20750 3562 20988
rect 3582 20750 3586 20988
rect 3606 20750 3610 20988
rect 3613 20987 3627 20988
rect 3630 20987 3637 20988
rect 3829 20987 3843 20988
rect 3835 20977 3843 20981
rect 3829 20967 3835 20977
rect 3643 20964 3677 20967
rect 3630 20750 3634 20964
rect 3829 20963 3843 20964
rect 3846 20963 3853 20988
rect 3859 20981 3864 20988
rect 3877 20987 3891 20988
rect 4549 20987 4563 20988
rect 4566 20987 4573 21012
rect 4579 21005 4584 21012
rect 4597 21011 4611 21012
rect 4789 21011 4803 21012
rect 4806 21011 4813 21036
rect 4819 21029 4824 21036
rect 4837 21035 4851 21036
rect 6589 21035 6603 21036
rect 6606 21035 6613 21060
rect 6619 21053 6624 21060
rect 6629 21039 6634 21053
rect 4829 21015 4834 21029
rect 4843 21025 4851 21029
rect 4837 21015 4843 21025
rect 4589 20991 4594 21005
rect 4603 21001 4611 21005
rect 4597 20991 4603 21001
rect 3869 20967 3874 20981
rect 3883 20977 3891 20981
rect 3877 20967 3883 20977
rect 3654 20750 3658 20940
rect 3678 20926 3685 20939
rect 3678 20902 3685 20916
rect 3678 20867 3685 20892
rect 3678 20750 3682 20867
rect 3691 20837 3696 20847
rect 3701 20823 3706 20837
rect 3691 20765 3696 20775
rect 3702 20765 3706 20823
rect 3701 20751 3706 20765
rect 3715 20761 3723 20765
rect 3709 20751 3715 20761
rect 3691 20750 3723 20751
rect -2393 20748 3723 20750
rect -2371 20726 -2366 20748
rect -2348 20726 -2343 20748
rect -2325 20726 -2320 20748
rect -2054 20747 -1906 20748
rect -2054 20746 -2036 20747
rect -2309 20732 -2301 20742
rect -2317 20726 -2309 20732
rect -2068 20731 -2038 20738
rect -2000 20730 -1992 20747
rect -1920 20746 -1906 20747
rect -1846 20740 -1794 20748
rect -1852 20733 -1804 20738
rect -1902 20731 -1804 20733
rect -1655 20732 -1647 20742
rect -2000 20728 -1975 20730
rect -1902 20729 -1852 20731
rect -2025 20726 -1975 20728
rect -1846 20726 -1804 20729
rect -1663 20726 -1655 20732
rect -1642 20726 -1637 20748
rect -1619 20726 -1614 20748
rect -1530 20726 -1526 20748
rect -1506 20726 -1502 20748
rect -1482 20726 -1478 20748
rect -1458 20726 -1454 20748
rect -1434 20726 -1430 20748
rect -1410 20726 -1406 20748
rect -1386 20726 -1382 20748
rect -1362 20726 -1358 20748
rect -1338 20726 -1334 20748
rect -1314 20726 -1310 20748
rect -1290 20726 -1286 20748
rect -1266 20726 -1262 20748
rect -1242 20726 -1238 20748
rect -1218 20726 -1214 20748
rect -1194 20726 -1190 20748
rect -1170 20726 -1166 20748
rect -1146 20726 -1142 20748
rect -1122 20726 -1118 20748
rect -1098 20726 -1094 20748
rect -1074 20726 -1070 20748
rect -1050 20726 -1046 20748
rect -1026 20726 -1022 20748
rect -1002 20726 -998 20748
rect -978 20726 -974 20748
rect -954 20726 -950 20748
rect -930 20726 -926 20748
rect -906 20726 -902 20748
rect -882 20726 -878 20748
rect -858 20726 -854 20748
rect -834 20726 -830 20748
rect -810 20726 -806 20748
rect -786 20726 -782 20748
rect -762 20726 -758 20748
rect -738 20726 -734 20748
rect -714 20726 -710 20748
rect -690 20726 -686 20748
rect -666 20726 -662 20748
rect -642 20726 -638 20748
rect -618 20726 -614 20748
rect -594 20726 -590 20748
rect -570 20726 -566 20748
rect -546 20726 -542 20748
rect -522 20726 -518 20748
rect -498 20726 -494 20748
rect -474 20726 -470 20748
rect -450 20726 -446 20748
rect -426 20726 -422 20748
rect -402 20726 -398 20748
rect -378 20726 -374 20748
rect -354 20726 -350 20748
rect -330 20726 -326 20748
rect -306 20726 -302 20748
rect -282 20726 -278 20748
rect -258 20726 -254 20748
rect -234 20726 -230 20748
rect -210 20726 -206 20748
rect -186 20726 -182 20748
rect -162 20726 -158 20748
rect -138 20726 -134 20748
rect -114 20726 -110 20748
rect -90 20726 -86 20748
rect -66 20726 -62 20748
rect -42 20726 -38 20748
rect -18 20726 -14 20748
rect 6 20726 10 20748
rect 30 20726 34 20748
rect 54 20726 58 20748
rect 78 20726 82 20748
rect 102 20726 106 20748
rect 126 20726 130 20748
rect 150 20726 154 20748
rect 174 20726 178 20748
rect 198 20726 202 20748
rect 222 20726 226 20748
rect 246 20726 250 20748
rect 270 20726 274 20748
rect 294 20747 298 20748
rect -2393 20724 291 20726
rect -2371 20702 -2366 20724
rect -2348 20702 -2343 20724
rect -2325 20702 -2320 20724
rect -2054 20723 -2038 20724
rect -2000 20723 -1966 20724
rect -1846 20723 -1804 20724
rect -2000 20722 -1975 20723
rect -2076 20714 -2054 20721
rect -2309 20704 -2301 20714
rect -2044 20711 -2038 20716
rect -2028 20714 -2001 20721
rect -2054 20704 -2038 20711
rect -2015 20713 -2001 20714
rect -2015 20704 -2014 20713
rect -2317 20702 -2309 20704
rect -2044 20702 -2028 20704
rect -2000 20702 -1992 20722
rect -1982 20721 -1975 20722
rect -1862 20721 -1798 20722
rect -1985 20714 -1796 20721
rect -1862 20713 -1798 20714
rect -1852 20704 -1804 20711
rect -1655 20704 -1647 20714
rect -1976 20702 -1940 20703
rect -1663 20702 -1655 20704
rect -1642 20702 -1637 20724
rect -1619 20702 -1614 20724
rect -1530 20702 -1526 20724
rect -1506 20702 -1502 20724
rect -1482 20702 -1478 20724
rect -1458 20702 -1454 20724
rect -1434 20702 -1430 20724
rect -1410 20702 -1406 20724
rect -1386 20702 -1382 20724
rect -1362 20702 -1358 20724
rect -1338 20702 -1334 20724
rect -1314 20702 -1310 20724
rect -1290 20702 -1286 20724
rect -1266 20702 -1262 20724
rect -1242 20702 -1238 20724
rect -1218 20702 -1214 20724
rect -1194 20702 -1190 20724
rect -1170 20702 -1166 20724
rect -1146 20702 -1142 20724
rect -1122 20702 -1118 20724
rect -1098 20702 -1094 20724
rect -1074 20702 -1070 20724
rect -1050 20702 -1046 20724
rect -1026 20702 -1022 20724
rect -1002 20702 -998 20724
rect -978 20702 -974 20724
rect -954 20702 -950 20724
rect -930 20702 -926 20724
rect -906 20702 -902 20724
rect -882 20702 -878 20724
rect -858 20702 -854 20724
rect -834 20702 -830 20724
rect -810 20702 -806 20724
rect -786 20702 -782 20724
rect -762 20702 -758 20724
rect -738 20702 -734 20724
rect -714 20702 -710 20724
rect -690 20702 -686 20724
rect -666 20702 -662 20724
rect -642 20702 -638 20724
rect -618 20702 -614 20724
rect -594 20702 -590 20724
rect -570 20702 -566 20724
rect -546 20702 -542 20724
rect -522 20702 -518 20724
rect -498 20702 -494 20724
rect -474 20702 -470 20724
rect -450 20702 -446 20724
rect -426 20702 -422 20724
rect -402 20702 -398 20724
rect -378 20702 -374 20724
rect -354 20702 -350 20724
rect -330 20702 -326 20724
rect -306 20702 -302 20724
rect -282 20702 -278 20724
rect -258 20702 -254 20724
rect -234 20702 -230 20724
rect -210 20702 -206 20724
rect -186 20702 -182 20724
rect -162 20702 -158 20724
rect -138 20702 -134 20724
rect -114 20702 -110 20724
rect -90 20702 -86 20724
rect -66 20702 -62 20724
rect -42 20702 -38 20724
rect -18 20702 -14 20724
rect 6 20702 10 20724
rect 30 20702 34 20724
rect 54 20702 58 20724
rect 78 20702 82 20724
rect 102 20702 106 20724
rect 126 20702 130 20724
rect 150 20702 154 20724
rect 174 20702 178 20724
rect 198 20702 202 20724
rect 222 20702 226 20724
rect 246 20702 250 20724
rect 270 20702 274 20724
rect 277 20723 291 20724
rect 294 20702 301 20747
rect 318 20702 322 20748
rect 342 20702 346 20748
rect 366 20702 370 20748
rect 390 20702 394 20748
rect 414 20702 418 20748
rect 438 20702 442 20748
rect 462 20702 466 20748
rect 486 20702 490 20748
rect 510 20702 514 20748
rect 534 20702 538 20748
rect 558 20702 562 20748
rect 582 20702 586 20748
rect 606 20702 610 20748
rect 630 20702 634 20748
rect 654 20702 658 20748
rect 678 20702 682 20748
rect 702 20702 706 20748
rect 726 20702 730 20748
rect 750 20702 754 20748
rect 774 20702 778 20748
rect 798 20702 802 20748
rect 822 20702 826 20748
rect 846 20702 850 20748
rect 870 20702 874 20748
rect 894 20702 898 20748
rect 918 20702 922 20748
rect 942 20702 946 20748
rect 966 20702 970 20748
rect 990 20702 994 20748
rect 1014 20702 1018 20748
rect 1038 20702 1042 20748
rect 1062 20702 1066 20748
rect 1086 20703 1090 20748
rect 1075 20702 1109 20703
rect -2393 20700 1109 20702
rect -2371 20630 -2366 20700
rect -2348 20630 -2343 20700
rect -2325 20666 -2320 20700
rect -2317 20698 -2309 20700
rect -2076 20687 -2054 20694
rect -2325 20658 -2317 20666
rect -2060 20660 -2030 20663
rect -2325 20630 -2320 20658
rect -2317 20650 -2309 20658
rect -2060 20647 -2038 20658
rect -2033 20651 -2030 20660
rect -2028 20656 -2027 20660
rect -2068 20642 -2038 20645
rect -2000 20630 -1992 20700
rect -1846 20696 -1804 20700
rect -1663 20698 -1655 20700
rect -1846 20686 -1794 20695
rect -1912 20675 -1884 20677
rect -1852 20669 -1804 20673
rect -1844 20660 -1796 20663
rect -1671 20658 -1663 20666
rect -1844 20647 -1804 20658
rect -1663 20650 -1655 20658
rect -1852 20642 -1680 20646
rect -1979 20630 -1945 20632
rect -1642 20630 -1637 20700
rect -1619 20630 -1614 20700
rect -1530 20630 -1526 20700
rect -1506 20630 -1502 20700
rect -1482 20630 -1478 20700
rect -1458 20630 -1454 20700
rect -1434 20630 -1430 20700
rect -1410 20630 -1406 20700
rect -1386 20630 -1382 20700
rect -1362 20630 -1358 20700
rect -1338 20630 -1334 20700
rect -1314 20630 -1310 20700
rect -1290 20630 -1286 20700
rect -1266 20630 -1262 20700
rect -1242 20630 -1238 20700
rect -1218 20630 -1214 20700
rect -1194 20630 -1190 20700
rect -1170 20630 -1166 20700
rect -1146 20630 -1142 20700
rect -1122 20630 -1118 20700
rect -1098 20630 -1094 20700
rect -1074 20630 -1070 20700
rect -1050 20630 -1046 20700
rect -1026 20630 -1022 20700
rect -1002 20630 -998 20700
rect -978 20630 -974 20700
rect -954 20630 -950 20700
rect -930 20630 -926 20700
rect -906 20630 -902 20700
rect -882 20630 -878 20700
rect -858 20630 -854 20700
rect -834 20630 -830 20700
rect -810 20630 -806 20700
rect -786 20630 -782 20700
rect -762 20630 -758 20700
rect -738 20630 -734 20700
rect -714 20630 -710 20700
rect -690 20630 -686 20700
rect -666 20630 -662 20700
rect -642 20630 -638 20700
rect -618 20630 -614 20700
rect -594 20630 -590 20700
rect -570 20630 -566 20700
rect -546 20630 -542 20700
rect -522 20630 -518 20700
rect -498 20630 -494 20700
rect -474 20630 -470 20700
rect -450 20630 -446 20700
rect -426 20630 -422 20700
rect -402 20630 -398 20700
rect -378 20630 -374 20700
rect -354 20630 -350 20700
rect -330 20630 -326 20700
rect -306 20630 -302 20700
rect -282 20630 -278 20700
rect -258 20630 -254 20700
rect -234 20630 -230 20700
rect -210 20630 -206 20700
rect -186 20630 -182 20700
rect -162 20630 -158 20700
rect -138 20630 -134 20700
rect -114 20630 -110 20700
rect -90 20630 -86 20700
rect -66 20630 -62 20700
rect -42 20630 -38 20700
rect -18 20630 -14 20700
rect 6 20630 10 20700
rect 30 20630 34 20700
rect 54 20630 58 20700
rect 78 20630 82 20700
rect 102 20630 106 20700
rect 126 20630 130 20700
rect 150 20630 154 20700
rect 174 20630 178 20700
rect 198 20630 202 20700
rect 222 20630 226 20700
rect 246 20630 250 20700
rect 270 20630 274 20700
rect 277 20699 291 20700
rect 294 20699 301 20700
rect 294 20630 298 20699
rect 318 20630 322 20700
rect 342 20630 346 20700
rect 366 20630 370 20700
rect 390 20630 394 20700
rect 414 20630 418 20700
rect 438 20630 442 20700
rect 462 20630 466 20700
rect 486 20630 490 20700
rect 510 20630 514 20700
rect 534 20630 538 20700
rect 558 20630 562 20700
rect 582 20630 586 20700
rect 606 20630 610 20700
rect 630 20630 634 20700
rect 654 20630 658 20700
rect 678 20630 682 20700
rect 702 20630 706 20700
rect 726 20630 730 20700
rect 750 20630 754 20700
rect 774 20630 778 20700
rect 798 20630 802 20700
rect 822 20630 826 20700
rect 846 20630 850 20700
rect 870 20630 874 20700
rect 894 20630 898 20700
rect 918 20630 922 20700
rect 942 20630 946 20700
rect 966 20630 970 20700
rect 990 20630 994 20700
rect 1014 20630 1018 20700
rect 1038 20630 1042 20700
rect 1062 20630 1066 20700
rect 1075 20693 1080 20700
rect 1086 20693 1090 20700
rect 1085 20679 1090 20693
rect 1075 20654 1109 20655
rect 1110 20654 1114 20748
rect 1134 20654 1138 20748
rect 1158 20723 1162 20748
rect 1158 20678 1165 20723
rect 1182 20678 1186 20748
rect 1206 20678 1210 20748
rect 1230 20678 1234 20748
rect 1254 20678 1258 20748
rect 1278 20678 1282 20748
rect 1302 20678 1306 20748
rect 1326 20678 1330 20748
rect 1350 20678 1354 20748
rect 1374 20678 1378 20748
rect 1398 20678 1402 20748
rect 1422 20678 1426 20748
rect 1446 20678 1450 20748
rect 1470 20678 1474 20748
rect 1494 20678 1498 20748
rect 1518 20678 1522 20748
rect 1542 20678 1546 20748
rect 1566 20678 1570 20748
rect 1590 20678 1594 20748
rect 1614 20678 1618 20748
rect 1638 20678 1642 20748
rect 1662 20678 1666 20748
rect 1686 20678 1690 20748
rect 1710 20678 1714 20748
rect 1734 20678 1738 20748
rect 1758 20678 1762 20748
rect 1782 20678 1786 20748
rect 1806 20678 1810 20748
rect 1830 20678 1834 20748
rect 1854 20678 1858 20748
rect 1878 20678 1882 20748
rect 1902 20678 1906 20748
rect 1926 20678 1930 20748
rect 1950 20678 1954 20748
rect 1974 20678 1978 20748
rect 1998 20678 2002 20748
rect 2011 20717 2016 20727
rect 2022 20717 2026 20748
rect 2021 20703 2026 20717
rect 2011 20693 2016 20703
rect 2021 20679 2026 20693
rect 2046 20679 2050 20748
rect 2022 20678 2026 20679
rect 2035 20678 2069 20679
rect 1141 20676 2069 20678
rect 1141 20675 1155 20676
rect 1158 20675 1165 20676
rect 1158 20654 1162 20675
rect 1182 20654 1186 20676
rect 1206 20654 1210 20676
rect 1230 20654 1234 20676
rect 1254 20654 1258 20676
rect 1278 20654 1282 20676
rect 1302 20654 1306 20676
rect 1326 20654 1330 20676
rect 1350 20654 1354 20676
rect 1374 20654 1378 20676
rect 1398 20654 1402 20676
rect 1422 20654 1426 20676
rect 1446 20654 1450 20676
rect 1470 20654 1474 20676
rect 1494 20654 1498 20676
rect 1518 20654 1522 20676
rect 1542 20654 1546 20676
rect 1566 20654 1570 20676
rect 1590 20654 1594 20676
rect 1614 20654 1618 20676
rect 1638 20654 1642 20676
rect 1662 20654 1666 20676
rect 1686 20654 1690 20676
rect 1710 20654 1714 20676
rect 1734 20654 1738 20676
rect 1758 20654 1762 20676
rect 1782 20654 1786 20676
rect 1806 20654 1810 20676
rect 1830 20654 1834 20676
rect 1854 20654 1858 20676
rect 1878 20654 1882 20676
rect 1902 20654 1906 20676
rect 1926 20654 1930 20676
rect 1950 20654 1954 20676
rect 1974 20654 1978 20676
rect 1998 20654 2002 20676
rect 2022 20654 2026 20676
rect 2035 20669 2040 20676
rect 2046 20669 2050 20676
rect 2045 20655 2050 20669
rect 2070 20654 2074 20748
rect 2094 20654 2098 20748
rect 2118 20654 2122 20748
rect 2142 20654 2146 20748
rect 2166 20654 2170 20748
rect 2190 20654 2194 20748
rect 2214 20654 2218 20748
rect 2238 20654 2242 20748
rect 2262 20654 2266 20748
rect 2286 20654 2290 20748
rect 2310 20654 2314 20748
rect 2334 20654 2338 20748
rect 2358 20654 2362 20748
rect 2382 20654 2386 20748
rect 2406 20654 2410 20748
rect 2430 20654 2434 20748
rect 2454 20654 2458 20748
rect 2478 20654 2482 20748
rect 2502 20654 2506 20748
rect 2526 20654 2530 20748
rect 2550 20654 2554 20748
rect 2574 20654 2578 20748
rect 2598 20654 2602 20748
rect 2622 20654 2626 20748
rect 2646 20654 2650 20748
rect 2670 20654 2674 20748
rect 2694 20654 2698 20748
rect 2718 20654 2722 20748
rect 2742 20654 2746 20748
rect 2766 20654 2770 20748
rect 2790 20654 2794 20748
rect 2814 20654 2818 20748
rect 2838 20654 2842 20748
rect 2862 20654 2866 20748
rect 2886 20654 2890 20748
rect 2910 20654 2914 20748
rect 2934 20654 2938 20748
rect 2958 20654 2962 20748
rect 2982 20654 2986 20748
rect 3006 20654 3010 20748
rect 3030 20654 3034 20748
rect 3054 20654 3058 20748
rect 3078 20654 3082 20748
rect 3102 20654 3106 20748
rect 3126 20654 3130 20748
rect 3150 20654 3154 20748
rect 3174 20654 3178 20748
rect 3198 20654 3202 20748
rect 3222 20654 3226 20748
rect 3246 20654 3250 20748
rect 3270 20654 3274 20748
rect 3294 20654 3298 20748
rect 3318 20654 3322 20748
rect 3342 20654 3346 20748
rect 3366 20654 3370 20748
rect 3390 20654 3394 20748
rect 3414 20654 3418 20748
rect 3438 20654 3442 20748
rect 3462 20654 3466 20748
rect 3486 20654 3490 20748
rect 3510 20654 3514 20748
rect 3534 20654 3538 20748
rect 3558 20654 3562 20748
rect 3582 20654 3586 20748
rect 3606 20654 3610 20748
rect 3630 20654 3634 20748
rect 3654 20654 3658 20748
rect 3678 20655 3682 20748
rect 3691 20741 3696 20748
rect 3709 20747 3723 20748
rect 3701 20727 3706 20741
rect 3691 20693 3696 20703
rect 3702 20693 3706 20727
rect 3701 20679 3706 20693
rect 3715 20689 3723 20693
rect 3709 20679 3715 20689
rect 3667 20654 3701 20655
rect 1075 20652 3701 20654
rect 1075 20645 1080 20652
rect 1085 20631 1090 20645
rect 1086 20630 1090 20631
rect 1110 20630 1114 20652
rect 1134 20630 1138 20652
rect 1158 20630 1162 20652
rect 1182 20630 1186 20652
rect 1206 20630 1210 20652
rect 1230 20630 1234 20652
rect 1254 20630 1258 20652
rect 1278 20630 1282 20652
rect 1302 20630 1306 20652
rect 1326 20630 1330 20652
rect 1350 20630 1354 20652
rect 1374 20630 1378 20652
rect 1398 20630 1402 20652
rect 1422 20630 1426 20652
rect 1446 20630 1450 20652
rect 1470 20630 1474 20652
rect 1494 20630 1498 20652
rect 1518 20630 1522 20652
rect 1542 20630 1546 20652
rect 1566 20630 1570 20652
rect 1590 20630 1594 20652
rect 1614 20630 1618 20652
rect 1638 20630 1642 20652
rect 1662 20630 1666 20652
rect 1686 20630 1690 20652
rect 1710 20630 1714 20652
rect 1734 20630 1738 20652
rect 1758 20630 1762 20652
rect 1782 20630 1786 20652
rect 1806 20630 1810 20652
rect 1830 20630 1834 20652
rect 1854 20630 1858 20652
rect 1878 20630 1882 20652
rect 1902 20630 1906 20652
rect 1926 20630 1930 20652
rect 1950 20630 1954 20652
rect 1974 20630 1978 20652
rect 1998 20630 2002 20652
rect 2022 20630 2026 20652
rect 2035 20630 2043 20631
rect -2393 20628 2043 20630
rect -2371 20582 -2366 20628
rect -2348 20582 -2343 20628
rect -2325 20582 -2320 20628
rect -2309 20610 -2301 20618
rect -2068 20611 -2040 20618
rect -2317 20602 -2309 20610
rect -2000 20601 -1992 20628
rect -1850 20620 -1844 20628
rect -1840 20620 -1792 20628
rect -1894 20618 -1850 20619
rect -1958 20616 -1955 20617
rect -1969 20610 -1955 20616
rect -1894 20611 -1802 20618
rect -1894 20610 -1850 20611
rect -1655 20610 -1647 20618
rect -1969 20608 -1942 20610
rect -1955 20601 -1942 20608
rect -1844 20603 -1802 20609
rect -1663 20602 -1655 20610
rect -1860 20601 -1796 20602
rect -2040 20594 -2020 20601
rect -2004 20594 -1945 20601
rect -1929 20599 -1794 20601
rect -1929 20594 -1850 20599
rect -1844 20594 -1794 20599
rect -2309 20582 -2301 20590
rect -2136 20582 -2129 20592
rect -2068 20584 -2040 20591
rect -2020 20582 -2004 20584
rect -2000 20582 -1992 20594
rect -1844 20593 -1796 20594
rect -1850 20584 -1802 20591
rect -1978 20582 -1942 20583
rect -1655 20582 -1647 20590
rect -1642 20582 -1637 20628
rect -1619 20582 -1614 20628
rect -1530 20582 -1526 20628
rect -1506 20582 -1502 20628
rect -1482 20582 -1478 20628
rect -1458 20582 -1454 20628
rect -1434 20582 -1430 20628
rect -1410 20582 -1406 20628
rect -1386 20582 -1382 20628
rect -1362 20582 -1358 20628
rect -1338 20582 -1334 20628
rect -1314 20582 -1310 20628
rect -1290 20582 -1286 20628
rect -1266 20582 -1262 20628
rect -1242 20582 -1238 20628
rect -1218 20582 -1214 20628
rect -1194 20582 -1190 20628
rect -1170 20582 -1166 20628
rect -1146 20582 -1142 20628
rect -1122 20582 -1118 20628
rect -1098 20582 -1094 20628
rect -1074 20582 -1070 20628
rect -1050 20582 -1046 20628
rect -1026 20582 -1022 20628
rect -1002 20582 -998 20628
rect -978 20582 -974 20628
rect -954 20582 -950 20628
rect -930 20582 -926 20628
rect -906 20582 -902 20628
rect -882 20582 -878 20628
rect -858 20582 -854 20628
rect -834 20582 -830 20628
rect -810 20582 -806 20628
rect -786 20582 -782 20628
rect -762 20582 -758 20628
rect -738 20582 -734 20628
rect -714 20582 -710 20628
rect -690 20582 -686 20628
rect -666 20582 -662 20628
rect -642 20582 -638 20628
rect -618 20582 -614 20628
rect -594 20582 -590 20628
rect -570 20582 -566 20628
rect -546 20582 -542 20628
rect -522 20582 -518 20628
rect -498 20582 -494 20628
rect -474 20582 -470 20628
rect -450 20582 -446 20628
rect -426 20582 -422 20628
rect -402 20582 -398 20628
rect -378 20582 -374 20628
rect -354 20582 -350 20628
rect -330 20582 -326 20628
rect -306 20582 -302 20628
rect -282 20582 -278 20628
rect -258 20582 -254 20628
rect -234 20582 -230 20628
rect -210 20582 -206 20628
rect -186 20582 -182 20628
rect -162 20582 -158 20628
rect -138 20582 -134 20628
rect -114 20582 -110 20628
rect -90 20582 -86 20628
rect -66 20582 -62 20628
rect -42 20582 -38 20628
rect -18 20582 -14 20628
rect 6 20582 10 20628
rect 30 20582 34 20628
rect 54 20582 58 20628
rect 78 20582 82 20628
rect 102 20582 106 20628
rect 126 20582 130 20628
rect 150 20582 154 20628
rect 174 20582 178 20628
rect 198 20582 202 20628
rect 222 20582 226 20628
rect 246 20582 250 20628
rect 270 20583 274 20628
rect 259 20582 293 20583
rect -2393 20580 293 20582
rect -2371 20486 -2366 20580
rect -2348 20486 -2343 20580
rect -2325 20542 -2320 20580
rect -2317 20574 -2309 20580
rect -2124 20576 -2117 20580
rect -2060 20576 -2040 20580
rect -2060 20567 -2030 20574
rect -2062 20542 -2032 20543
rect -2000 20542 -1992 20580
rect -1844 20576 -1802 20580
rect -1844 20566 -1792 20575
rect -1663 20574 -1655 20580
rect -1942 20544 -1937 20556
rect -1850 20553 -1822 20554
rect -1850 20549 -1802 20553
rect -2325 20534 -2317 20542
rect -2062 20540 -1961 20542
rect -2325 20514 -2320 20534
rect -2317 20526 -2309 20534
rect -2062 20527 -2040 20538
rect -2032 20533 -1961 20540
rect -1947 20534 -1942 20542
rect -1842 20540 -1794 20543
rect -2070 20522 -2022 20526
rect -2325 20502 -2317 20514
rect -2325 20486 -2320 20502
rect -2317 20498 -2309 20502
rect -2309 20486 -2301 20498
rect -2068 20491 -2038 20498
rect -2000 20488 -1992 20533
rect -1942 20532 -1937 20534
rect -1932 20524 -1927 20532
rect -1912 20529 -1896 20535
rect -1842 20527 -1802 20538
rect -1671 20534 -1663 20542
rect -1663 20526 -1655 20534
rect -1850 20522 -1680 20526
rect -1937 20508 -1934 20510
rect -1926 20508 -1921 20513
rect -1926 20503 -1924 20508
rect -1916 20500 -1914 20503
rect -1842 20500 -1794 20509
rect -1671 20502 -1663 20514
rect -1924 20490 -1916 20499
rect -1663 20498 -1655 20502
rect -1852 20491 -1804 20498
rect -1916 20489 -1914 20490
rect -2025 20487 -1991 20488
rect -2025 20486 -1975 20487
rect -1842 20486 -1804 20489
rect -1655 20486 -1647 20498
rect -1642 20486 -1637 20580
rect -1619 20486 -1614 20580
rect -1530 20486 -1526 20580
rect -1506 20486 -1502 20580
rect -1482 20486 -1478 20580
rect -1458 20486 -1454 20580
rect -1434 20486 -1430 20580
rect -1410 20486 -1406 20580
rect -1397 20549 -1392 20559
rect -1386 20549 -1382 20580
rect -1387 20535 -1382 20549
rect -1386 20486 -1382 20535
rect -1362 20486 -1358 20580
rect -1338 20486 -1334 20580
rect -1314 20486 -1310 20580
rect -1290 20486 -1286 20580
rect -1266 20486 -1262 20580
rect -1242 20486 -1238 20580
rect -1218 20486 -1214 20580
rect -1194 20486 -1190 20580
rect -1170 20486 -1166 20580
rect -1146 20486 -1142 20580
rect -1122 20486 -1118 20580
rect -1098 20486 -1094 20580
rect -1074 20486 -1070 20580
rect -1050 20486 -1046 20580
rect -1026 20486 -1022 20580
rect -1002 20486 -998 20580
rect -978 20486 -974 20580
rect -954 20486 -950 20580
rect -930 20486 -926 20580
rect -906 20486 -902 20580
rect -882 20486 -878 20580
rect -858 20486 -854 20580
rect -834 20486 -830 20580
rect -810 20486 -806 20580
rect -786 20486 -782 20580
rect -762 20486 -758 20580
rect -738 20486 -734 20580
rect -714 20486 -710 20580
rect -690 20486 -686 20580
rect -666 20486 -662 20580
rect -642 20486 -638 20580
rect -618 20486 -614 20580
rect -594 20486 -590 20580
rect -570 20486 -566 20580
rect -546 20486 -542 20580
rect -522 20486 -518 20580
rect -498 20486 -494 20580
rect -474 20486 -470 20580
rect -450 20486 -446 20580
rect -426 20486 -422 20580
rect -402 20486 -398 20580
rect -378 20486 -374 20580
rect -354 20486 -350 20580
rect -330 20486 -326 20580
rect -306 20486 -302 20580
rect -282 20486 -278 20580
rect -258 20486 -254 20580
rect -234 20486 -230 20580
rect -210 20486 -206 20580
rect -186 20486 -182 20580
rect -162 20486 -158 20580
rect -138 20486 -134 20580
rect -114 20486 -110 20580
rect -90 20486 -86 20580
rect -66 20486 -62 20580
rect -42 20486 -38 20580
rect -18 20486 -14 20580
rect 6 20486 10 20580
rect 30 20486 34 20580
rect 54 20486 58 20580
rect 78 20486 82 20580
rect 102 20486 106 20580
rect 126 20486 130 20580
rect 150 20486 154 20580
rect 174 20486 178 20580
rect 198 20486 202 20580
rect 222 20486 226 20580
rect 246 20486 250 20580
rect 259 20573 264 20580
rect 270 20573 274 20580
rect 269 20559 274 20573
rect 270 20486 274 20559
rect 294 20507 298 20628
rect -2393 20484 291 20486
rect -2371 20462 -2366 20484
rect -2348 20462 -2343 20484
rect -2325 20474 -2317 20484
rect -2076 20474 -2068 20481
rect -2062 20474 -2001 20481
rect -2325 20462 -2320 20474
rect -2317 20470 -2309 20474
rect -2015 20473 -2001 20474
rect -2309 20462 -2301 20470
rect -2068 20464 -2062 20471
rect -2000 20466 -1992 20484
rect -1974 20482 -1960 20484
rect -1842 20483 -1804 20484
rect -1862 20481 -1794 20482
rect -1985 20479 -1794 20481
rect -1985 20474 -1852 20479
rect -1842 20473 -1794 20479
rect -1671 20474 -1663 20484
rect -2015 20464 -1985 20466
rect -1852 20464 -1804 20471
rect -1663 20470 -1655 20474
rect -2000 20462 -1992 20464
rect -1976 20462 -1940 20463
rect -1655 20462 -1647 20470
rect -1642 20462 -1637 20484
rect -1619 20462 -1614 20484
rect -1530 20462 -1526 20484
rect -1506 20462 -1502 20484
rect -1482 20462 -1478 20484
rect -1458 20462 -1454 20484
rect -1434 20462 -1430 20484
rect -1410 20462 -1406 20484
rect -1386 20462 -1382 20484
rect -1362 20483 -1358 20484
rect -2393 20460 -1365 20462
rect -2371 20390 -2366 20460
rect -2348 20390 -2343 20460
rect -2325 20458 -2320 20460
rect -2309 20458 -2301 20460
rect -2325 20446 -2317 20458
rect -2062 20447 -2032 20454
rect -2325 20426 -2320 20446
rect -2317 20442 -2309 20446
rect -2325 20418 -2317 20426
rect -2060 20420 -2030 20423
rect -2325 20390 -2320 20418
rect -2317 20410 -2309 20418
rect -2060 20407 -2038 20418
rect -2033 20411 -2030 20420
rect -2028 20416 -2027 20420
rect -2068 20402 -2038 20405
rect -2000 20390 -1992 20460
rect -1888 20455 -1874 20460
rect -1842 20456 -1804 20460
rect -1655 20458 -1647 20460
rect -1902 20453 -1874 20455
rect -1842 20446 -1794 20455
rect -1671 20446 -1663 20458
rect -1663 20442 -1655 20446
rect -1912 20435 -1884 20437
rect -1852 20429 -1804 20433
rect -1844 20420 -1796 20423
rect -1671 20418 -1663 20426
rect -1844 20407 -1804 20418
rect -1663 20410 -1655 20418
rect -1852 20402 -1680 20406
rect -1979 20390 -1945 20392
rect -1642 20390 -1637 20460
rect -1619 20390 -1614 20460
rect -1530 20390 -1526 20460
rect -1506 20390 -1502 20460
rect -1482 20390 -1478 20460
rect -1458 20390 -1454 20460
rect -1434 20390 -1430 20460
rect -1410 20390 -1406 20460
rect -1386 20390 -1382 20460
rect -1379 20459 -1365 20460
rect -1362 20459 -1355 20483
rect -1362 20390 -1358 20459
rect -1338 20390 -1334 20484
rect -1314 20390 -1310 20484
rect -1290 20390 -1286 20484
rect -1266 20390 -1262 20484
rect -1242 20390 -1238 20484
rect -1218 20390 -1214 20484
rect -1194 20390 -1190 20484
rect -1170 20390 -1166 20484
rect -1146 20390 -1142 20484
rect -1122 20390 -1118 20484
rect -1098 20390 -1094 20484
rect -1074 20390 -1070 20484
rect -1050 20390 -1046 20484
rect -1026 20390 -1022 20484
rect -1002 20390 -998 20484
rect -978 20390 -974 20484
rect -954 20390 -950 20484
rect -930 20390 -926 20484
rect -906 20390 -902 20484
rect -882 20390 -878 20484
rect -858 20390 -854 20484
rect -834 20390 -830 20484
rect -810 20390 -806 20484
rect -786 20390 -782 20484
rect -762 20390 -758 20484
rect -738 20390 -734 20484
rect -714 20390 -710 20484
rect -690 20390 -686 20484
rect -666 20390 -662 20484
rect -642 20390 -638 20484
rect -618 20390 -614 20484
rect -594 20390 -590 20484
rect -570 20390 -566 20484
rect -546 20390 -542 20484
rect -522 20390 -518 20484
rect -498 20390 -494 20484
rect -474 20390 -470 20484
rect -450 20390 -446 20484
rect -426 20390 -422 20484
rect -402 20390 -398 20484
rect -378 20390 -374 20484
rect -354 20390 -350 20484
rect -330 20390 -326 20484
rect -306 20390 -302 20484
rect -282 20390 -278 20484
rect -258 20390 -254 20484
rect -234 20390 -230 20484
rect -210 20390 -206 20484
rect -186 20390 -182 20484
rect -162 20390 -158 20484
rect -138 20390 -134 20484
rect -114 20390 -110 20484
rect -90 20390 -86 20484
rect -66 20390 -62 20484
rect -42 20390 -38 20484
rect -18 20390 -14 20484
rect 6 20390 10 20484
rect 30 20390 34 20484
rect 54 20390 58 20484
rect 78 20390 82 20484
rect 102 20390 106 20484
rect 126 20390 130 20484
rect 150 20390 154 20484
rect 174 20390 178 20484
rect 198 20390 202 20484
rect 222 20390 226 20484
rect 246 20390 250 20484
rect 270 20390 274 20484
rect 277 20483 291 20484
rect 294 20483 301 20507
rect 294 20390 298 20483
rect 318 20390 322 20628
rect 342 20390 346 20628
rect 366 20390 370 20628
rect 390 20390 394 20628
rect 414 20390 418 20628
rect 438 20390 442 20628
rect 462 20390 466 20628
rect 486 20390 490 20628
rect 510 20390 514 20628
rect 534 20390 538 20628
rect 558 20390 562 20628
rect 582 20390 586 20628
rect 606 20390 610 20628
rect 630 20390 634 20628
rect 654 20390 658 20628
rect 678 20390 682 20628
rect 702 20390 706 20628
rect 726 20390 730 20628
rect 750 20390 754 20628
rect 774 20390 778 20628
rect 798 20390 802 20628
rect 822 20390 826 20628
rect 846 20390 850 20628
rect 870 20390 874 20628
rect 894 20390 898 20628
rect 918 20390 922 20628
rect 942 20390 946 20628
rect 966 20390 970 20628
rect 990 20390 994 20628
rect 1014 20390 1018 20628
rect 1038 20390 1042 20628
rect 1062 20390 1066 20628
rect 1086 20390 1090 20628
rect 1110 20627 1114 20628
rect 1110 20603 1117 20627
rect 1110 20555 1117 20579
rect 1110 20390 1114 20555
rect 1134 20390 1138 20628
rect 1158 20390 1162 20628
rect 1182 20390 1186 20628
rect 1206 20390 1210 20628
rect 1230 20390 1234 20628
rect 1254 20390 1258 20628
rect 1278 20390 1282 20628
rect 1302 20390 1306 20628
rect 1326 20390 1330 20628
rect 1350 20390 1354 20628
rect 1374 20390 1378 20628
rect 1398 20390 1402 20628
rect 1422 20390 1426 20628
rect 1446 20390 1450 20628
rect 1470 20390 1474 20628
rect 1494 20390 1498 20628
rect 1518 20390 1522 20628
rect 1542 20390 1546 20628
rect 1566 20390 1570 20628
rect 1590 20390 1594 20628
rect 1614 20390 1618 20628
rect 1638 20390 1642 20628
rect 1662 20390 1666 20628
rect 1686 20390 1690 20628
rect 1710 20390 1714 20628
rect 1734 20390 1738 20628
rect 1758 20390 1762 20628
rect 1782 20390 1786 20628
rect 1806 20390 1810 20628
rect 1830 20390 1834 20628
rect 1854 20390 1858 20628
rect 1878 20390 1882 20628
rect 1902 20390 1906 20628
rect 1926 20390 1930 20628
rect 1950 20390 1954 20628
rect 1974 20390 1978 20628
rect 1998 20390 2002 20628
rect 2022 20390 2026 20628
rect 2029 20627 2043 20628
rect 2045 20607 2053 20621
rect 2046 20603 2053 20607
rect 2070 20603 2074 20652
rect 2046 20390 2050 20603
rect 2070 20579 2077 20603
rect 2070 20531 2077 20555
rect 2070 20390 2074 20531
rect 2094 20390 2098 20652
rect 2118 20390 2122 20652
rect 2142 20390 2146 20652
rect 2166 20390 2170 20652
rect 2190 20390 2194 20652
rect 2214 20390 2218 20652
rect 2238 20390 2242 20652
rect 2262 20390 2266 20652
rect 2286 20390 2290 20652
rect 2310 20390 2314 20652
rect 2334 20390 2338 20652
rect 2358 20390 2362 20652
rect 2382 20390 2386 20652
rect 2406 20390 2410 20652
rect 2430 20390 2434 20652
rect 2454 20390 2458 20652
rect 2478 20390 2482 20652
rect 2502 20390 2506 20652
rect 2526 20390 2530 20652
rect 2550 20390 2554 20652
rect 2574 20390 2578 20652
rect 2598 20390 2602 20652
rect 2622 20390 2626 20652
rect 2646 20390 2650 20652
rect 2670 20390 2674 20652
rect 2694 20390 2698 20652
rect 2718 20390 2722 20652
rect 2742 20390 2746 20652
rect 2766 20390 2770 20652
rect 2790 20390 2794 20652
rect 2803 20453 2808 20463
rect 2814 20453 2818 20652
rect 2813 20439 2818 20453
rect 2803 20429 2808 20439
rect 2813 20415 2818 20429
rect 2814 20390 2818 20415
rect 2838 20390 2842 20652
rect 2862 20390 2866 20652
rect 2886 20390 2890 20652
rect 2910 20390 2914 20652
rect 2934 20390 2938 20652
rect 2958 20390 2962 20652
rect 2982 20390 2986 20652
rect 3006 20390 3010 20652
rect 3019 20429 3024 20439
rect 3030 20429 3034 20652
rect 3029 20415 3034 20429
rect 3019 20414 3053 20415
rect 3054 20414 3058 20652
rect 3078 20414 3082 20652
rect 3102 20414 3106 20652
rect 3126 20414 3130 20652
rect 3150 20414 3154 20652
rect 3174 20414 3178 20652
rect 3198 20414 3202 20652
rect 3222 20414 3226 20652
rect 3246 20414 3250 20652
rect 3259 20477 3264 20487
rect 3270 20477 3274 20652
rect 3269 20463 3274 20477
rect 3270 20414 3274 20463
rect 3294 20414 3298 20652
rect 3318 20414 3322 20652
rect 3342 20414 3346 20652
rect 3366 20414 3370 20652
rect 3390 20414 3394 20652
rect 3414 20414 3418 20652
rect 3438 20414 3442 20652
rect 3462 20414 3466 20652
rect 3486 20414 3490 20652
rect 3510 20414 3514 20652
rect 3534 20414 3538 20652
rect 3558 20414 3562 20652
rect 3582 20414 3586 20652
rect 3606 20414 3610 20652
rect 3630 20414 3634 20652
rect 3654 20414 3658 20652
rect 3667 20645 3672 20652
rect 3678 20645 3682 20652
rect 3677 20631 3682 20645
rect 3667 20501 3672 20511
rect 3677 20487 3682 20501
rect 3678 20415 3682 20487
rect 3667 20414 3699 20415
rect 3019 20412 3699 20414
rect 3019 20405 3024 20412
rect 3029 20391 3034 20405
rect 3030 20390 3034 20391
rect 3054 20390 3058 20412
rect 3078 20390 3082 20412
rect 3102 20390 3106 20412
rect 3126 20390 3130 20412
rect 3150 20390 3154 20412
rect 3174 20390 3178 20412
rect 3198 20390 3202 20412
rect 3222 20390 3226 20412
rect 3246 20390 3250 20412
rect 3270 20390 3274 20412
rect 3294 20411 3298 20412
rect -2393 20388 3291 20390
rect -2371 20342 -2366 20388
rect -2348 20342 -2343 20388
rect -2325 20342 -2320 20388
rect -2309 20370 -2301 20378
rect -2068 20371 -2040 20378
rect -2317 20362 -2309 20370
rect -2000 20361 -1992 20388
rect -1850 20380 -1844 20388
rect -1840 20380 -1792 20388
rect -1894 20378 -1850 20379
rect -1958 20376 -1955 20377
rect -1969 20370 -1955 20376
rect -1894 20371 -1802 20378
rect -1894 20370 -1850 20371
rect -1655 20370 -1647 20378
rect -1969 20368 -1942 20370
rect -1955 20361 -1942 20368
rect -1844 20363 -1802 20369
rect -1663 20362 -1655 20370
rect -1860 20361 -1796 20362
rect -2040 20354 -2020 20361
rect -2004 20354 -1945 20361
rect -1929 20359 -1794 20361
rect -1929 20354 -1850 20359
rect -1844 20354 -1794 20359
rect -2309 20342 -2301 20350
rect -2136 20342 -2129 20352
rect -2068 20344 -2040 20351
rect -2020 20342 -2004 20344
rect -2000 20342 -1992 20354
rect -1844 20353 -1796 20354
rect -1850 20344 -1802 20351
rect -1978 20342 -1942 20343
rect -1655 20342 -1647 20350
rect -1642 20342 -1637 20388
rect -1619 20342 -1614 20388
rect -1530 20342 -1526 20388
rect -1506 20342 -1502 20388
rect -1482 20342 -1478 20388
rect -1458 20342 -1454 20388
rect -1434 20342 -1430 20388
rect -1410 20342 -1406 20388
rect -1386 20342 -1382 20388
rect -1362 20342 -1358 20388
rect -1338 20342 -1334 20388
rect -1314 20342 -1310 20388
rect -1290 20342 -1286 20388
rect -1266 20342 -1262 20388
rect -1242 20342 -1238 20388
rect -1218 20342 -1214 20388
rect -1194 20342 -1190 20388
rect -1170 20342 -1166 20388
rect -1146 20342 -1142 20388
rect -1122 20342 -1118 20388
rect -1098 20342 -1094 20388
rect -1074 20342 -1070 20388
rect -1050 20342 -1046 20388
rect -1026 20342 -1022 20388
rect -1002 20342 -998 20388
rect -978 20342 -974 20388
rect -954 20342 -950 20388
rect -930 20342 -926 20388
rect -906 20342 -902 20388
rect -882 20342 -878 20388
rect -858 20342 -854 20388
rect -834 20342 -830 20388
rect -810 20342 -806 20388
rect -786 20342 -782 20388
rect -762 20342 -758 20388
rect -738 20342 -734 20388
rect -714 20342 -710 20388
rect -690 20342 -686 20388
rect -666 20342 -662 20388
rect -642 20342 -638 20388
rect -618 20342 -614 20388
rect -594 20342 -590 20388
rect -570 20342 -566 20388
rect -546 20342 -542 20388
rect -522 20342 -518 20388
rect -498 20342 -494 20388
rect -474 20342 -470 20388
rect -450 20342 -446 20388
rect -426 20342 -422 20388
rect -402 20342 -398 20388
rect -378 20342 -374 20388
rect -354 20342 -350 20388
rect -330 20342 -326 20388
rect -306 20342 -302 20388
rect -282 20342 -278 20388
rect -258 20342 -254 20388
rect -234 20342 -230 20388
rect -210 20342 -206 20388
rect -186 20342 -182 20388
rect -162 20342 -158 20388
rect -138 20342 -134 20388
rect -114 20342 -110 20388
rect -90 20342 -86 20388
rect -66 20342 -62 20388
rect -42 20342 -38 20388
rect -18 20342 -14 20388
rect 6 20342 10 20388
rect 30 20342 34 20388
rect 54 20342 58 20388
rect 78 20342 82 20388
rect 102 20342 106 20388
rect 126 20342 130 20388
rect 150 20342 154 20388
rect 174 20342 178 20388
rect 198 20342 202 20388
rect 222 20342 226 20388
rect 246 20342 250 20388
rect 270 20343 274 20388
rect 259 20342 293 20343
rect -2393 20340 293 20342
rect -2371 20222 -2366 20340
rect -2348 20222 -2343 20340
rect -2325 20302 -2320 20340
rect -2317 20334 -2309 20340
rect -2124 20336 -2117 20340
rect -2060 20336 -2040 20340
rect -2060 20327 -2030 20334
rect -2062 20302 -2032 20303
rect -2000 20302 -1992 20340
rect -1844 20336 -1802 20340
rect -1844 20326 -1792 20335
rect -1663 20334 -1655 20340
rect -1942 20304 -1937 20316
rect -1850 20313 -1822 20314
rect -1850 20309 -1802 20313
rect -2325 20294 -2317 20302
rect -2062 20300 -1961 20302
rect -2325 20274 -2320 20294
rect -2317 20286 -2309 20294
rect -2062 20287 -2040 20298
rect -2032 20293 -1961 20300
rect -1947 20294 -1942 20302
rect -1842 20300 -1794 20303
rect -2070 20282 -2022 20286
rect -2325 20258 -2317 20274
rect -2080 20260 -2032 20269
rect -2325 20242 -2320 20258
rect -2309 20246 -2301 20258
rect -2070 20251 -2040 20258
rect -2317 20242 -2309 20246
rect -2325 20230 -2317 20242
rect -2000 20241 -1992 20293
rect -1942 20292 -1937 20294
rect -1932 20284 -1927 20292
rect -1912 20289 -1896 20295
rect -1842 20287 -1802 20298
rect -1671 20294 -1663 20302
rect -1663 20286 -1655 20294
rect -1850 20282 -1680 20286
rect -1937 20268 -1934 20270
rect -1924 20268 -1921 20270
rect -1850 20260 -1842 20270
rect -1840 20260 -1792 20269
rect -1924 20258 -1850 20259
rect -1671 20258 -1663 20274
rect -1960 20256 -1955 20257
rect -1969 20250 -1955 20256
rect -1924 20251 -1802 20258
rect -1924 20250 -1850 20251
rect -1969 20248 -1944 20250
rect -1955 20241 -1944 20248
rect -1842 20243 -1802 20249
rect -1655 20246 -1647 20258
rect -1663 20242 -1655 20246
rect -1860 20241 -1794 20242
rect -2040 20234 -1945 20241
rect -1929 20239 -1794 20241
rect -1929 20234 -1850 20239
rect -2325 20222 -2320 20230
rect -2309 20222 -2301 20230
rect -2070 20224 -2040 20231
rect -2000 20222 -1992 20234
rect -1842 20233 -1794 20239
rect -1945 20224 -1942 20226
rect -1850 20224 -1802 20231
rect -1671 20230 -1663 20242
rect -1978 20222 -1942 20223
rect -1655 20222 -1647 20230
rect -1642 20222 -1637 20340
rect -1619 20222 -1614 20340
rect -1530 20222 -1526 20340
rect -1506 20222 -1502 20340
rect -1482 20222 -1478 20340
rect -1458 20222 -1454 20340
rect -1434 20222 -1430 20340
rect -1410 20222 -1406 20340
rect -1386 20222 -1382 20340
rect -1362 20222 -1358 20340
rect -1338 20222 -1334 20340
rect -1314 20222 -1310 20340
rect -1290 20222 -1286 20340
rect -1266 20222 -1262 20340
rect -1242 20222 -1238 20340
rect -1218 20222 -1214 20340
rect -1194 20222 -1190 20340
rect -1170 20222 -1166 20340
rect -1146 20222 -1142 20340
rect -1122 20222 -1118 20340
rect -1098 20222 -1094 20340
rect -1074 20222 -1070 20340
rect -1050 20222 -1046 20340
rect -1026 20222 -1022 20340
rect -1002 20222 -998 20340
rect -978 20222 -974 20340
rect -954 20222 -950 20340
rect -930 20222 -926 20340
rect -906 20222 -902 20340
rect -882 20222 -878 20340
rect -858 20222 -854 20340
rect -834 20222 -830 20340
rect -810 20222 -806 20340
rect -786 20222 -782 20340
rect -762 20222 -758 20340
rect -738 20222 -734 20340
rect -714 20222 -710 20340
rect -690 20222 -686 20340
rect -666 20222 -662 20340
rect -642 20222 -638 20340
rect -629 20309 -624 20319
rect -618 20309 -614 20340
rect -619 20295 -614 20309
rect -618 20222 -614 20295
rect -594 20243 -590 20340
rect -2393 20220 -597 20222
rect -2371 20126 -2366 20220
rect -2348 20126 -2343 20220
rect -2325 20214 -2320 20220
rect -2309 20218 -2301 20220
rect -2317 20214 -2309 20218
rect -2062 20216 -2040 20220
rect -2325 20202 -2317 20214
rect -2062 20207 -2032 20214
rect -2325 20182 -2320 20202
rect -2062 20182 -2032 20183
rect -2000 20182 -1992 20220
rect -1888 20215 -1874 20220
rect -1842 20216 -1802 20220
rect -1655 20218 -1647 20220
rect -1932 20206 -1924 20215
rect -1904 20213 -1874 20215
rect -1842 20206 -1792 20215
rect -1663 20214 -1655 20218
rect -1671 20202 -1663 20214
rect -1942 20184 -1937 20196
rect -1850 20193 -1822 20194
rect -1850 20189 -1802 20193
rect -2325 20174 -2317 20182
rect -2062 20180 -1961 20182
rect -2325 20154 -2320 20174
rect -2317 20166 -2309 20174
rect -2062 20167 -2040 20178
rect -2032 20173 -1961 20180
rect -1947 20174 -1942 20182
rect -1842 20180 -1794 20183
rect -2070 20162 -2022 20166
rect -2325 20142 -2317 20154
rect -2325 20126 -2320 20142
rect -2317 20138 -2309 20142
rect -2309 20126 -2301 20138
rect -2068 20131 -2038 20138
rect -2000 20128 -1992 20173
rect -1942 20172 -1937 20174
rect -1932 20164 -1927 20172
rect -1912 20169 -1896 20175
rect -1842 20167 -1802 20178
rect -1671 20174 -1663 20182
rect -1663 20166 -1655 20174
rect -1850 20162 -1680 20166
rect -1937 20148 -1934 20150
rect -1926 20148 -1921 20153
rect -1926 20143 -1924 20148
rect -1916 20140 -1914 20143
rect -1842 20140 -1794 20149
rect -1671 20142 -1663 20154
rect -1924 20130 -1916 20139
rect -1663 20138 -1655 20142
rect -1852 20131 -1804 20138
rect -1916 20129 -1914 20130
rect -2025 20127 -1991 20128
rect -2025 20126 -1975 20127
rect -1842 20126 -1804 20129
rect -1655 20126 -1647 20138
rect -1642 20126 -1637 20220
rect -1619 20126 -1614 20220
rect -1530 20126 -1526 20220
rect -1506 20126 -1502 20220
rect -1482 20126 -1478 20220
rect -1458 20126 -1454 20220
rect -1434 20126 -1430 20220
rect -1410 20126 -1406 20220
rect -1386 20126 -1382 20220
rect -1362 20126 -1358 20220
rect -1338 20126 -1334 20220
rect -1314 20126 -1310 20220
rect -1290 20126 -1286 20220
rect -1266 20126 -1262 20220
rect -1242 20126 -1238 20220
rect -1218 20126 -1214 20220
rect -1194 20126 -1190 20220
rect -1170 20126 -1166 20220
rect -1146 20126 -1142 20220
rect -1122 20126 -1118 20220
rect -1098 20126 -1094 20220
rect -1074 20126 -1070 20220
rect -1050 20126 -1046 20220
rect -1026 20126 -1022 20220
rect -1002 20126 -998 20220
rect -978 20126 -974 20220
rect -954 20126 -950 20220
rect -930 20126 -926 20220
rect -906 20126 -902 20220
rect -882 20126 -878 20220
rect -858 20126 -854 20220
rect -834 20126 -830 20220
rect -810 20126 -806 20220
rect -786 20126 -782 20220
rect -762 20126 -758 20220
rect -738 20126 -734 20220
rect -714 20126 -710 20220
rect -690 20126 -686 20220
rect -666 20126 -662 20220
rect -642 20126 -638 20220
rect -618 20126 -614 20220
rect -611 20219 -597 20220
rect -594 20219 -587 20243
rect -594 20126 -590 20219
rect -570 20126 -566 20340
rect -546 20126 -542 20340
rect -522 20126 -518 20340
rect -498 20126 -494 20340
rect -474 20126 -470 20340
rect -450 20126 -446 20340
rect -426 20126 -422 20340
rect -402 20126 -398 20340
rect -378 20126 -374 20340
rect -354 20126 -350 20340
rect -330 20126 -326 20340
rect -306 20126 -302 20340
rect -282 20126 -278 20340
rect -258 20126 -254 20340
rect -234 20126 -230 20340
rect -210 20126 -206 20340
rect -186 20126 -182 20340
rect -162 20126 -158 20340
rect -138 20126 -134 20340
rect -114 20126 -110 20340
rect -90 20126 -86 20340
rect -66 20126 -62 20340
rect -42 20126 -38 20340
rect -18 20126 -14 20340
rect 6 20126 10 20340
rect 30 20126 34 20340
rect 54 20126 58 20340
rect 78 20126 82 20340
rect 102 20126 106 20340
rect 126 20126 130 20340
rect 150 20126 154 20340
rect 174 20126 178 20340
rect 198 20126 202 20340
rect 222 20126 226 20340
rect 246 20126 250 20340
rect 259 20333 264 20340
rect 270 20333 274 20340
rect 269 20319 274 20333
rect 259 20189 264 20199
rect 270 20189 274 20319
rect 269 20175 274 20189
rect 270 20126 274 20175
rect 294 20267 298 20388
rect 294 20243 301 20267
rect 294 20126 298 20243
rect 318 20126 322 20388
rect 342 20126 346 20388
rect 366 20126 370 20388
rect 390 20126 394 20388
rect 414 20126 418 20388
rect 438 20126 442 20388
rect 462 20126 466 20388
rect 486 20127 490 20388
rect 475 20126 509 20127
rect -2393 20124 509 20126
rect -2371 20102 -2366 20124
rect -2348 20102 -2343 20124
rect -2325 20114 -2317 20124
rect -2076 20114 -2068 20121
rect -2062 20114 -2001 20121
rect -2325 20102 -2320 20114
rect -2317 20110 -2309 20114
rect -2015 20113 -2001 20114
rect -2309 20102 -2301 20110
rect -2068 20104 -2062 20111
rect -2000 20106 -1992 20124
rect -1974 20122 -1960 20124
rect -1842 20123 -1804 20124
rect -1862 20121 -1794 20122
rect -1985 20119 -1794 20121
rect -1985 20114 -1852 20119
rect -1842 20113 -1794 20119
rect -1671 20114 -1663 20124
rect -2015 20104 -1985 20106
rect -1852 20104 -1804 20111
rect -1663 20110 -1655 20114
rect -2000 20102 -1992 20104
rect -1976 20102 -1940 20103
rect -1655 20102 -1647 20110
rect -1642 20102 -1637 20124
rect -1619 20102 -1614 20124
rect -1530 20102 -1526 20124
rect -1506 20103 -1502 20124
rect -1517 20102 -1483 20103
rect -2393 20100 -1483 20102
rect -2371 20030 -2366 20100
rect -2348 20030 -2343 20100
rect -2325 20098 -2320 20100
rect -2309 20098 -2301 20100
rect -2325 20086 -2317 20098
rect -2062 20087 -2032 20094
rect -2325 20066 -2320 20086
rect -2317 20082 -2309 20086
rect -2325 20058 -2317 20066
rect -2060 20060 -2030 20063
rect -2325 20038 -2320 20058
rect -2317 20050 -2309 20058
rect -2060 20047 -2038 20058
rect -2033 20051 -2030 20060
rect -2028 20056 -2027 20060
rect -2068 20042 -2038 20045
rect -2325 20030 -2317 20038
rect -2000 20030 -1992 20100
rect -1888 20095 -1874 20100
rect -1842 20096 -1804 20100
rect -1655 20098 -1647 20100
rect -1902 20093 -1874 20095
rect -1842 20086 -1794 20095
rect -1671 20086 -1663 20098
rect -1663 20082 -1655 20086
rect -1912 20075 -1884 20077
rect -1852 20069 -1804 20073
rect -1844 20060 -1796 20063
rect -1671 20058 -1663 20066
rect -1844 20047 -1804 20058
rect -1663 20050 -1655 20058
rect -1852 20042 -1680 20046
rect -1926 20030 -1892 20033
rect -1671 20030 -1663 20038
rect -1642 20030 -1637 20100
rect -1619 20030 -1614 20100
rect -1530 20030 -1526 20100
rect -1517 20093 -1512 20100
rect -1506 20093 -1502 20100
rect -1507 20079 -1502 20093
rect -1506 20030 -1502 20079
rect -1482 20030 -1478 20124
rect -1458 20030 -1454 20124
rect -1434 20030 -1430 20124
rect -1410 20030 -1406 20124
rect -1386 20030 -1382 20124
rect -1362 20030 -1358 20124
rect -1338 20030 -1334 20124
rect -1314 20030 -1310 20124
rect -1290 20030 -1286 20124
rect -1266 20030 -1262 20124
rect -1242 20030 -1238 20124
rect -1218 20030 -1214 20124
rect -1194 20030 -1190 20124
rect -1170 20030 -1166 20124
rect -1146 20030 -1142 20124
rect -1122 20030 -1118 20124
rect -1098 20030 -1094 20124
rect -1074 20030 -1070 20124
rect -1050 20030 -1046 20124
rect -1026 20030 -1022 20124
rect -1002 20030 -998 20124
rect -978 20030 -974 20124
rect -954 20030 -950 20124
rect -930 20030 -926 20124
rect -906 20030 -902 20124
rect -882 20030 -878 20124
rect -858 20030 -854 20124
rect -834 20030 -830 20124
rect -810 20030 -806 20124
rect -786 20030 -782 20124
rect -762 20030 -758 20124
rect -738 20030 -734 20124
rect -714 20030 -710 20124
rect -690 20030 -686 20124
rect -666 20030 -662 20124
rect -642 20030 -638 20124
rect -618 20030 -614 20124
rect -594 20030 -590 20124
rect -570 20030 -566 20124
rect -546 20030 -542 20124
rect -522 20030 -518 20124
rect -498 20030 -494 20124
rect -474 20030 -470 20124
rect -450 20030 -446 20124
rect -426 20030 -422 20124
rect -402 20030 -398 20124
rect -378 20030 -374 20124
rect -354 20030 -350 20124
rect -330 20030 -326 20124
rect -306 20030 -302 20124
rect -282 20030 -278 20124
rect -258 20030 -254 20124
rect -234 20030 -230 20124
rect -210 20030 -206 20124
rect -186 20030 -182 20124
rect -162 20030 -158 20124
rect -138 20030 -134 20124
rect -114 20030 -110 20124
rect -90 20030 -86 20124
rect -66 20030 -62 20124
rect -42 20030 -38 20124
rect -18 20030 -14 20124
rect 6 20030 10 20124
rect 30 20030 34 20124
rect 54 20030 58 20124
rect 78 20030 82 20124
rect 102 20030 106 20124
rect 126 20030 130 20124
rect 150 20030 154 20124
rect 174 20030 178 20124
rect 198 20030 202 20124
rect 222 20030 226 20124
rect 246 20030 250 20124
rect 259 20069 264 20079
rect 270 20069 274 20124
rect 269 20055 274 20069
rect 270 20030 274 20055
rect 294 20123 298 20124
rect 294 20099 301 20123
rect 294 20030 298 20099
rect 318 20030 322 20124
rect 342 20030 346 20124
rect 366 20030 370 20124
rect 390 20030 394 20124
rect 414 20030 418 20124
rect 438 20030 442 20124
rect 462 20030 466 20124
rect 475 20117 480 20124
rect 486 20117 490 20124
rect 485 20103 490 20117
rect 486 20030 490 20103
rect 510 20051 514 20388
rect -2393 20028 507 20030
rect -2371 20006 -2366 20028
rect -2348 20006 -2343 20028
rect -2325 20022 -2317 20028
rect -2325 20006 -2320 20022
rect -2309 20010 -2301 20022
rect -2068 20011 -2038 20018
rect -2317 20006 -2309 20010
rect -2000 20008 -1992 20028
rect -1844 20020 -1794 20028
rect -1671 20022 -1663 20028
rect -1852 20011 -1804 20018
rect -1655 20010 -1647 20022
rect -2025 20007 -1991 20008
rect -2025 20006 -1975 20007
rect -1844 20006 -1804 20009
rect -1663 20006 -1655 20010
rect -1642 20006 -1637 20028
rect -1619 20006 -1614 20028
rect -1530 20006 -1526 20028
rect -1506 20006 -1502 20028
rect -1482 20027 -1478 20028
rect -2393 20004 -1485 20006
rect -2371 19982 -2366 20004
rect -2348 19982 -2343 20004
rect -2325 19994 -2317 20004
rect -2060 19994 -2020 20001
rect -2004 19996 -2001 20001
rect -2015 19994 -2001 19996
rect -2000 19994 -1992 20004
rect -1972 20002 -1958 20004
rect -1844 20003 -1804 20004
rect -1862 20001 -1796 20002
rect -1985 19999 -1796 20001
rect -1985 19994 -1852 19999
rect -2325 19982 -2320 19994
rect -2309 19982 -2301 19994
rect -2068 19984 -2060 19991
rect -2015 19984 -1990 19994
rect -1844 19993 -1796 19999
rect -1671 19994 -1663 20004
rect -1852 19984 -1804 19991
rect -2020 19982 -2004 19984
rect -2000 19982 -1992 19984
rect -1976 19982 -1940 19983
rect -1655 19982 -1647 19994
rect -1642 19982 -1637 20004
rect -1619 19982 -1614 20004
rect -1530 19982 -1526 20004
rect -1506 19982 -1502 20004
rect -1499 20003 -1485 20004
rect -1482 20003 -1475 20027
rect -1482 19982 -1478 20003
rect -1458 19982 -1454 20028
rect -1434 19982 -1430 20028
rect -1410 19982 -1406 20028
rect -1386 19982 -1382 20028
rect -1362 19982 -1358 20028
rect -1338 19982 -1334 20028
rect -1314 19982 -1310 20028
rect -1290 19982 -1286 20028
rect -1266 19982 -1262 20028
rect -1242 19982 -1238 20028
rect -1218 19982 -1214 20028
rect -1194 19982 -1190 20028
rect -1170 19982 -1166 20028
rect -1146 19982 -1142 20028
rect -1122 19982 -1118 20028
rect -1098 19982 -1094 20028
rect -1074 19982 -1070 20028
rect -1050 19982 -1046 20028
rect -1026 19982 -1022 20028
rect -1002 19982 -998 20028
rect -978 19982 -974 20028
rect -954 19982 -950 20028
rect -930 19982 -926 20028
rect -906 19982 -902 20028
rect -882 19982 -878 20028
rect -858 19982 -854 20028
rect -834 19982 -830 20028
rect -810 19982 -806 20028
rect -786 19982 -782 20028
rect -762 19982 -758 20028
rect -738 19982 -734 20028
rect -714 19982 -710 20028
rect -690 19982 -686 20028
rect -666 19982 -662 20028
rect -642 19982 -638 20028
rect -618 19982 -614 20028
rect -594 19982 -590 20028
rect -570 19982 -566 20028
rect -546 19982 -542 20028
rect -522 19982 -518 20028
rect -498 19982 -494 20028
rect -474 19982 -470 20028
rect -450 19983 -446 20028
rect -461 19982 -427 19983
rect -2393 19980 -427 19982
rect -2371 19910 -2366 19980
rect -2348 19910 -2343 19980
rect -2325 19978 -2320 19980
rect -2317 19978 -2309 19980
rect -2325 19966 -2317 19978
rect -2060 19967 -2030 19974
rect -2325 19946 -2320 19966
rect -2325 19938 -2317 19946
rect -2060 19940 -2030 19943
rect -2325 19918 -2320 19938
rect -2317 19930 -2309 19938
rect -2060 19927 -2038 19938
rect -2033 19931 -2030 19940
rect -2028 19936 -2027 19940
rect -2068 19922 -2038 19925
rect -2325 19910 -2317 19918
rect -2000 19910 -1992 19980
rect -1844 19976 -1804 19980
rect -1663 19978 -1655 19980
rect -1844 19966 -1794 19975
rect -1671 19966 -1663 19978
rect -1912 19955 -1884 19957
rect -1852 19949 -1804 19953
rect -1844 19940 -1796 19943
rect -1671 19938 -1663 19946
rect -1844 19927 -1804 19938
rect -1663 19930 -1655 19938
rect -1852 19922 -1680 19926
rect -1671 19910 -1663 19918
rect -1642 19910 -1637 19980
rect -1619 19910 -1614 19980
rect -1530 19910 -1526 19980
rect -1506 19910 -1502 19980
rect -1482 19910 -1478 19980
rect -1458 19910 -1454 19980
rect -1434 19910 -1430 19980
rect -1410 19910 -1406 19980
rect -1386 19910 -1382 19980
rect -1362 19910 -1358 19980
rect -1338 19910 -1334 19980
rect -1314 19910 -1310 19980
rect -1290 19910 -1286 19980
rect -1266 19910 -1262 19980
rect -1242 19910 -1238 19980
rect -1218 19910 -1214 19980
rect -1194 19910 -1190 19980
rect -1170 19910 -1166 19980
rect -1146 19910 -1142 19980
rect -1122 19910 -1118 19980
rect -1098 19910 -1094 19980
rect -1074 19910 -1070 19980
rect -1050 19910 -1046 19980
rect -1026 19910 -1022 19980
rect -1002 19910 -998 19980
rect -978 19910 -974 19980
rect -954 19910 -950 19980
rect -930 19910 -926 19980
rect -906 19910 -902 19980
rect -882 19910 -878 19980
rect -858 19910 -854 19980
rect -834 19910 -830 19980
rect -810 19910 -806 19980
rect -786 19910 -782 19980
rect -762 19910 -758 19980
rect -738 19910 -734 19980
rect -714 19910 -710 19980
rect -690 19910 -686 19980
rect -666 19910 -662 19980
rect -642 19910 -638 19980
rect -618 19910 -614 19980
rect -594 19910 -590 19980
rect -570 19910 -566 19980
rect -546 19910 -542 19980
rect -522 19910 -518 19980
rect -498 19910 -494 19980
rect -474 19910 -470 19980
rect -461 19973 -456 19980
rect -450 19973 -446 19980
rect -451 19959 -446 19973
rect -450 19910 -446 19959
rect -426 19910 -422 20028
rect -402 19910 -398 20028
rect -378 19910 -374 20028
rect -354 19910 -350 20028
rect -330 19910 -326 20028
rect -306 19910 -302 20028
rect -282 19910 -278 20028
rect -258 19910 -254 20028
rect -234 19910 -230 20028
rect -210 19910 -206 20028
rect -186 19910 -182 20028
rect -162 19910 -158 20028
rect -138 19910 -134 20028
rect -114 19910 -110 20028
rect -90 19910 -86 20028
rect -66 19910 -62 20028
rect -42 19910 -38 20028
rect -18 19910 -14 20028
rect 6 19910 10 20028
rect 30 19910 34 20028
rect 54 19910 58 20028
rect 78 19910 82 20028
rect 102 19910 106 20028
rect 126 19910 130 20028
rect 150 19910 154 20028
rect 174 19910 178 20028
rect 198 19910 202 20028
rect 222 19910 226 20028
rect 246 19910 250 20028
rect 270 19910 274 20028
rect 294 20003 298 20028
rect 294 19979 301 20003
rect 294 19910 298 19979
rect 318 19910 322 20028
rect 342 19910 346 20028
rect 366 19910 370 20028
rect 390 19910 394 20028
rect 414 19910 418 20028
rect 438 19910 442 20028
rect 462 19910 466 20028
rect 486 19910 490 20028
rect 493 20027 507 20028
rect 510 20027 517 20051
rect 510 19910 514 20027
rect 534 19910 538 20388
rect 558 19910 562 20388
rect 582 19910 586 20388
rect 606 19910 610 20388
rect 630 19910 634 20388
rect 654 19910 658 20388
rect 678 19910 682 20388
rect 702 19910 706 20388
rect 726 19910 730 20388
rect 750 19910 754 20388
rect 774 19910 778 20388
rect 798 19910 802 20388
rect 822 19910 826 20388
rect 846 19910 850 20388
rect 870 19910 874 20388
rect 894 19910 898 20388
rect 918 19910 922 20388
rect 942 19910 946 20388
rect 966 19910 970 20388
rect 990 19910 994 20388
rect 1014 19910 1018 20388
rect 1038 19910 1042 20388
rect 1062 19910 1066 20388
rect 1086 19910 1090 20388
rect 1110 19910 1114 20388
rect 1134 19910 1138 20388
rect 1158 19910 1162 20388
rect 1182 19910 1186 20388
rect 1206 19910 1210 20388
rect 1230 19910 1234 20388
rect 1254 19910 1258 20388
rect 1278 19910 1282 20388
rect 1302 19910 1306 20388
rect 1326 19910 1330 20388
rect 1350 19910 1354 20388
rect 1374 19910 1378 20388
rect 1398 19910 1402 20388
rect 1422 19910 1426 20388
rect 1446 19910 1450 20388
rect 1470 19910 1474 20388
rect 1494 19910 1498 20388
rect 1518 19910 1522 20388
rect 1542 19910 1546 20388
rect 1566 19910 1570 20388
rect 1590 19910 1594 20388
rect 1614 19910 1618 20388
rect 1638 19910 1642 20388
rect 1662 19910 1666 20388
rect 1686 19910 1690 20388
rect 1710 19910 1714 20388
rect 1734 19910 1738 20388
rect 1758 19910 1762 20388
rect 1782 19910 1786 20388
rect 1806 19910 1810 20388
rect 1830 19910 1834 20388
rect 1854 19910 1858 20388
rect 1867 19997 1872 20007
rect 1878 19997 1882 20388
rect 1877 19983 1882 19997
rect 1878 19910 1882 19983
rect 1902 19931 1906 20388
rect -2393 19908 1899 19910
rect -2371 19862 -2366 19908
rect -2348 19862 -2343 19908
rect -2325 19902 -2317 19908
rect -2325 19886 -2320 19902
rect -2309 19890 -2301 19902
rect -2317 19886 -2309 19890
rect -2000 19886 -1992 19908
rect -1671 19902 -1663 19908
rect -1977 19891 -1929 19897
rect -2325 19874 -2317 19886
rect -2030 19884 -1992 19886
rect -2030 19882 -1980 19884
rect -1972 19882 -1942 19891
rect -1655 19890 -1647 19902
rect -1663 19886 -1655 19890
rect -2059 19878 -2045 19882
rect -2325 19862 -2320 19874
rect -2309 19862 -2301 19874
rect -2025 19872 -2020 19876
rect -2292 19871 -2095 19872
rect -2025 19866 -2009 19872
rect -2000 19866 -1992 19882
rect -1958 19881 -1942 19882
rect -1671 19874 -1663 19886
rect -1977 19869 -1929 19871
rect -2033 19864 -1992 19866
rect -2060 19862 -1992 19864
rect -1655 19862 -1647 19874
rect -1642 19862 -1637 19908
rect -1619 19862 -1614 19908
rect -1530 19862 -1526 19908
rect -1506 19862 -1502 19908
rect -1482 19862 -1478 19908
rect -1458 19862 -1454 19908
rect -1434 19862 -1430 19908
rect -1410 19862 -1406 19908
rect -1386 19862 -1382 19908
rect -1362 19862 -1358 19908
rect -1338 19862 -1334 19908
rect -1314 19862 -1310 19908
rect -1290 19862 -1286 19908
rect -1266 19862 -1262 19908
rect -1242 19862 -1238 19908
rect -1218 19862 -1214 19908
rect -1194 19862 -1190 19908
rect -1170 19862 -1166 19908
rect -1146 19862 -1142 19908
rect -1122 19862 -1118 19908
rect -1098 19862 -1094 19908
rect -1074 19862 -1070 19908
rect -1050 19862 -1046 19908
rect -1026 19862 -1022 19908
rect -1002 19862 -998 19908
rect -978 19862 -974 19908
rect -954 19862 -950 19908
rect -930 19862 -926 19908
rect -906 19862 -902 19908
rect -882 19862 -878 19908
rect -858 19862 -854 19908
rect -834 19862 -830 19908
rect -810 19862 -806 19908
rect -786 19862 -782 19908
rect -762 19862 -758 19908
rect -738 19862 -734 19908
rect -714 19862 -710 19908
rect -690 19862 -686 19908
rect -666 19862 -662 19908
rect -642 19862 -638 19908
rect -618 19862 -614 19908
rect -594 19862 -590 19908
rect -570 19862 -566 19908
rect -546 19862 -542 19908
rect -522 19863 -518 19908
rect -533 19862 -499 19863
rect -2393 19860 -499 19862
rect -2371 19742 -2366 19860
rect -2348 19742 -2343 19860
rect -2325 19858 -2320 19860
rect -2317 19858 -2309 19860
rect -2325 19846 -2317 19858
rect -2124 19846 -2108 19860
rect -2025 19856 -2020 19860
rect -2060 19846 -2030 19847
rect -2023 19846 -2020 19856
rect -2325 19826 -2320 19846
rect -2325 19818 -2317 19826
rect -2325 19798 -2320 19818
rect -2317 19810 -2309 19818
rect -2117 19809 -2095 19819
rect -2045 19816 -2037 19830
rect -2325 19782 -2317 19798
rect -2325 19766 -2320 19782
rect -2309 19770 -2301 19782
rect -2317 19766 -2309 19770
rect -2117 19768 -2095 19775
rect -2069 19774 -2041 19782
rect -2017 19780 -2015 19782
rect -2325 19754 -2317 19766
rect -2125 19759 -2095 19766
rect -2047 19764 -2011 19766
rect -2059 19762 -2011 19764
rect -2000 19762 -1992 19860
rect -1663 19858 -1655 19860
rect -1671 19846 -1663 19858
rect -1969 19809 -1929 19821
rect -1671 19818 -1663 19826
rect -1663 19810 -1655 19818
rect -1671 19782 -1663 19798
rect -1655 19770 -1647 19782
rect -1663 19766 -1655 19770
rect -2125 19757 -2117 19759
rect -2059 19758 -2045 19762
rect -2021 19759 -1992 19762
rect -1977 19759 -1929 19766
rect -2325 19742 -2320 19754
rect -2309 19742 -2301 19754
rect -2131 19749 -2129 19754
rect -2125 19751 -2095 19757
rect -2021 19752 -2009 19756
rect -2125 19749 -2117 19751
rect -2133 19742 -2129 19749
rect -2117 19742 -2087 19749
rect -2025 19746 -2021 19752
rect -2000 19746 -1992 19759
rect -1969 19751 -1929 19757
rect -1671 19754 -1663 19766
rect -2033 19742 -1992 19746
rect -1969 19742 -1921 19749
rect -1655 19742 -1647 19754
rect -1642 19742 -1637 19860
rect -1619 19742 -1614 19860
rect -1530 19742 -1526 19860
rect -1506 19742 -1502 19860
rect -1482 19742 -1478 19860
rect -1458 19742 -1454 19860
rect -1434 19742 -1430 19860
rect -1410 19742 -1406 19860
rect -1386 19742 -1382 19860
rect -1362 19742 -1358 19860
rect -1338 19742 -1334 19860
rect -1314 19742 -1310 19860
rect -1290 19742 -1286 19860
rect -1266 19742 -1262 19860
rect -1242 19742 -1238 19860
rect -1218 19742 -1214 19860
rect -1194 19742 -1190 19860
rect -1170 19742 -1166 19860
rect -1146 19742 -1142 19860
rect -1122 19742 -1118 19860
rect -1098 19742 -1094 19860
rect -1074 19742 -1070 19860
rect -1050 19742 -1046 19860
rect -1026 19742 -1022 19860
rect -1002 19742 -998 19860
rect -978 19742 -974 19860
rect -954 19742 -950 19860
rect -930 19742 -926 19860
rect -906 19742 -902 19860
rect -882 19742 -878 19860
rect -858 19742 -854 19860
rect -834 19742 -830 19860
rect -810 19742 -806 19860
rect -786 19742 -782 19860
rect -762 19742 -758 19860
rect -738 19742 -734 19860
rect -714 19742 -710 19860
rect -690 19742 -686 19860
rect -666 19742 -662 19860
rect -642 19742 -638 19860
rect -618 19742 -614 19860
rect -594 19742 -590 19860
rect -570 19742 -566 19860
rect -546 19742 -542 19860
rect -533 19853 -528 19860
rect -522 19853 -518 19860
rect -523 19839 -518 19853
rect -522 19742 -518 19839
rect -498 19787 -494 19908
rect -498 19763 -491 19787
rect -498 19742 -494 19763
rect -474 19742 -470 19908
rect -450 19742 -446 19908
rect -426 19907 -422 19908
rect -426 19883 -419 19907
rect -426 19742 -422 19883
rect -402 19742 -398 19908
rect -378 19742 -374 19908
rect -354 19742 -350 19908
rect -330 19742 -326 19908
rect -306 19742 -302 19908
rect -282 19742 -278 19908
rect -258 19742 -254 19908
rect -234 19742 -230 19908
rect -210 19742 -206 19908
rect -186 19742 -182 19908
rect -162 19742 -158 19908
rect -138 19742 -134 19908
rect -114 19742 -110 19908
rect -90 19742 -86 19908
rect -66 19742 -62 19908
rect -42 19742 -38 19908
rect -18 19742 -14 19908
rect 6 19742 10 19908
rect 30 19742 34 19908
rect 54 19742 58 19908
rect 78 19742 82 19908
rect 102 19742 106 19908
rect 126 19742 130 19908
rect 150 19742 154 19908
rect 174 19742 178 19908
rect 198 19742 202 19908
rect 222 19742 226 19908
rect 246 19742 250 19908
rect 270 19742 274 19908
rect 294 19742 298 19908
rect 318 19742 322 19908
rect 342 19742 346 19908
rect 366 19742 370 19908
rect 390 19742 394 19908
rect 414 19742 418 19908
rect 438 19742 442 19908
rect 462 19742 466 19908
rect 486 19742 490 19908
rect 510 19742 514 19908
rect 534 19742 538 19908
rect 558 19742 562 19908
rect 582 19742 586 19908
rect 606 19742 610 19908
rect 630 19742 634 19908
rect 654 19742 658 19908
rect 678 19742 682 19908
rect 702 19742 706 19908
rect 726 19742 730 19908
rect 750 19742 754 19908
rect 774 19742 778 19908
rect 798 19742 802 19908
rect 822 19742 826 19908
rect 846 19742 850 19908
rect 870 19742 874 19908
rect 894 19742 898 19908
rect 918 19742 922 19908
rect 942 19742 946 19908
rect 966 19742 970 19908
rect 990 19742 994 19908
rect 1014 19742 1018 19908
rect 1038 19742 1042 19908
rect 1062 19742 1066 19908
rect 1086 19742 1090 19908
rect 1110 19742 1114 19908
rect 1134 19742 1138 19908
rect 1158 19742 1162 19908
rect 1182 19742 1186 19908
rect 1206 19742 1210 19908
rect 1230 19742 1234 19908
rect 1254 19742 1258 19908
rect 1278 19742 1282 19908
rect 1302 19742 1306 19908
rect 1326 19742 1330 19908
rect 1350 19742 1354 19908
rect 1374 19742 1378 19908
rect 1398 19742 1402 19908
rect 1411 19829 1416 19839
rect 1422 19829 1426 19908
rect 1421 19815 1426 19829
rect 1422 19742 1426 19815
rect 1446 19763 1450 19908
rect -2393 19740 1443 19742
rect -2371 19646 -2366 19740
rect -2348 19646 -2343 19740
rect -2325 19738 -2320 19740
rect -2317 19738 -2309 19740
rect -2131 19738 -2129 19740
rect -2125 19738 -2095 19740
rect -2325 19726 -2317 19738
rect -2117 19733 -2095 19738
rect -2325 19706 -2320 19726
rect -2325 19698 -2317 19706
rect -2325 19646 -2320 19698
rect -2317 19690 -2309 19698
rect -2117 19689 -2095 19699
rect -2045 19696 -2037 19710
rect -2309 19650 -2301 19658
rect -2317 19646 -2309 19650
rect -2000 19646 -1992 19740
rect -1663 19738 -1655 19740
rect -1671 19726 -1663 19738
rect -1969 19689 -1929 19701
rect -1671 19698 -1663 19706
rect -1663 19690 -1655 19698
rect -1655 19650 -1647 19658
rect -1663 19646 -1655 19650
rect -1642 19646 -1637 19740
rect -1619 19646 -1614 19740
rect -1530 19646 -1526 19740
rect -1506 19646 -1502 19740
rect -1482 19646 -1478 19740
rect -1458 19646 -1454 19740
rect -1434 19646 -1430 19740
rect -1410 19646 -1406 19740
rect -1386 19646 -1382 19740
rect -1362 19646 -1358 19740
rect -1338 19646 -1334 19740
rect -1314 19646 -1310 19740
rect -1290 19646 -1286 19740
rect -1266 19646 -1262 19740
rect -1242 19646 -1238 19740
rect -1218 19646 -1214 19740
rect -1194 19646 -1190 19740
rect -1170 19646 -1166 19740
rect -1146 19646 -1142 19740
rect -1122 19646 -1118 19740
rect -1098 19646 -1094 19740
rect -1074 19646 -1070 19740
rect -1050 19646 -1046 19740
rect -1026 19646 -1022 19740
rect -1002 19646 -998 19740
rect -978 19646 -974 19740
rect -954 19646 -950 19740
rect -930 19646 -926 19740
rect -906 19646 -902 19740
rect -882 19646 -878 19740
rect -858 19646 -854 19740
rect -834 19646 -830 19740
rect -810 19646 -806 19740
rect -786 19646 -782 19740
rect -762 19646 -758 19740
rect -738 19646 -734 19740
rect -714 19646 -710 19740
rect -690 19646 -686 19740
rect -666 19646 -662 19740
rect -642 19646 -638 19740
rect -618 19646 -614 19740
rect -594 19646 -590 19740
rect -570 19646 -566 19740
rect -546 19646 -542 19740
rect -522 19646 -518 19740
rect -498 19646 -494 19740
rect -474 19646 -470 19740
rect -450 19646 -446 19740
rect -426 19646 -422 19740
rect -402 19646 -398 19740
rect -378 19646 -374 19740
rect -354 19646 -350 19740
rect -330 19646 -326 19740
rect -306 19646 -302 19740
rect -282 19646 -278 19740
rect -258 19646 -254 19740
rect -234 19646 -230 19740
rect -210 19646 -206 19740
rect -186 19646 -182 19740
rect -162 19646 -158 19740
rect -138 19646 -134 19740
rect -114 19646 -110 19740
rect -90 19646 -86 19740
rect -66 19646 -62 19740
rect -42 19646 -38 19740
rect -18 19646 -14 19740
rect 6 19646 10 19740
rect 30 19646 34 19740
rect 54 19646 58 19740
rect 78 19646 82 19740
rect 102 19646 106 19740
rect 126 19646 130 19740
rect 150 19646 154 19740
rect 174 19646 178 19740
rect 198 19646 202 19740
rect 222 19646 226 19740
rect 246 19646 250 19740
rect 270 19646 274 19740
rect 294 19646 298 19740
rect 318 19646 322 19740
rect 342 19646 346 19740
rect 366 19646 370 19740
rect 390 19646 394 19740
rect 414 19646 418 19740
rect 438 19646 442 19740
rect 462 19646 466 19740
rect 486 19646 490 19740
rect 510 19646 514 19740
rect 534 19646 538 19740
rect 558 19646 562 19740
rect 582 19646 586 19740
rect 606 19646 610 19740
rect 630 19646 634 19740
rect 654 19646 658 19740
rect 678 19646 682 19740
rect 702 19646 706 19740
rect 726 19646 730 19740
rect 750 19646 754 19740
rect 774 19646 778 19740
rect 798 19646 802 19740
rect 822 19646 826 19740
rect 846 19646 850 19740
rect 870 19646 874 19740
rect 894 19646 898 19740
rect 918 19646 922 19740
rect 942 19646 946 19740
rect 966 19646 970 19740
rect 990 19646 994 19740
rect 1014 19646 1018 19740
rect 1038 19646 1042 19740
rect 1062 19646 1066 19740
rect 1086 19646 1090 19740
rect 1110 19646 1114 19740
rect 1134 19646 1138 19740
rect 1158 19646 1162 19740
rect 1182 19646 1186 19740
rect 1206 19646 1210 19740
rect 1230 19646 1234 19740
rect 1254 19646 1258 19740
rect 1278 19646 1282 19740
rect 1302 19646 1306 19740
rect 1326 19646 1330 19740
rect 1350 19646 1354 19740
rect 1374 19646 1378 19740
rect 1398 19646 1402 19740
rect 1422 19646 1426 19740
rect 1429 19739 1443 19740
rect 1446 19739 1453 19763
rect 1446 19646 1450 19739
rect 1470 19646 1474 19908
rect 1494 19646 1498 19908
rect 1518 19646 1522 19908
rect 1542 19646 1546 19908
rect 1566 19646 1570 19908
rect 1590 19646 1594 19908
rect 1614 19646 1618 19908
rect 1638 19646 1642 19908
rect 1662 19646 1666 19908
rect 1686 19646 1690 19908
rect 1710 19646 1714 19908
rect 1734 19646 1738 19908
rect 1758 19646 1762 19908
rect 1782 19646 1786 19908
rect 1806 19646 1810 19908
rect 1830 19646 1834 19908
rect 1854 19646 1858 19908
rect 1878 19646 1882 19908
rect 1885 19907 1899 19908
rect 1902 19907 1909 19931
rect 1902 19646 1906 19907
rect 1926 19646 1930 20388
rect 1950 19646 1954 20388
rect 1963 19709 1968 19719
rect 1974 19709 1978 20388
rect 1987 19949 1992 19959
rect 1998 19949 2002 20388
rect 1997 19935 2002 19949
rect 1987 19934 2021 19935
rect 2022 19934 2026 20388
rect 2046 19934 2050 20388
rect 2070 19934 2074 20388
rect 2094 19934 2098 20388
rect 2118 19934 2122 20388
rect 2142 19934 2146 20388
rect 2166 19934 2170 20388
rect 2190 19934 2194 20388
rect 2214 19934 2218 20388
rect 2238 19934 2242 20388
rect 2262 19934 2266 20388
rect 2286 19934 2290 20388
rect 2310 19934 2314 20388
rect 2334 19934 2338 20388
rect 2358 19934 2362 20388
rect 2382 19934 2386 20388
rect 2406 19934 2410 20388
rect 2430 19934 2434 20388
rect 2454 19934 2458 20388
rect 2478 19934 2482 20388
rect 2502 19934 2506 20388
rect 2526 19934 2530 20388
rect 2550 19934 2554 20388
rect 2574 19934 2578 20388
rect 2598 19934 2602 20388
rect 2622 19934 2626 20388
rect 2646 19934 2650 20388
rect 2670 19934 2674 20388
rect 2694 19934 2698 20388
rect 2718 19934 2722 20388
rect 2742 19934 2746 20388
rect 2766 19934 2770 20388
rect 2790 19934 2794 20388
rect 2814 19934 2818 20388
rect 2838 20387 2842 20388
rect 2838 20339 2845 20387
rect 2838 19934 2842 20339
rect 2862 19934 2866 20388
rect 2886 19934 2890 20388
rect 2910 19934 2914 20388
rect 2934 19934 2938 20388
rect 2958 19934 2962 20388
rect 2982 19934 2986 20388
rect 3006 19934 3010 20388
rect 3030 19934 3034 20388
rect 3054 20363 3058 20388
rect 3054 20315 3061 20363
rect 3054 19934 3058 20315
rect 3078 19934 3082 20388
rect 3102 19934 3106 20388
rect 3126 19934 3130 20388
rect 3150 19934 3154 20388
rect 3174 19934 3178 20388
rect 3198 19934 3202 20388
rect 3222 19934 3226 20388
rect 3246 19934 3250 20388
rect 3259 20213 3264 20223
rect 3270 20213 3274 20388
rect 3277 20387 3291 20388
rect 3294 20387 3301 20411
rect 3269 20199 3274 20213
rect 3259 20189 3264 20199
rect 3269 20175 3274 20189
rect 3270 19934 3274 20175
rect 3294 20147 3298 20387
rect 3294 20099 3301 20147
rect 3294 19934 3298 20099
rect 3318 19934 3322 20412
rect 3342 19934 3346 20412
rect 3366 19934 3370 20412
rect 3390 19934 3394 20412
rect 3414 19934 3418 20412
rect 3438 19934 3442 20412
rect 3462 19934 3466 20412
rect 3486 19934 3490 20412
rect 3510 19934 3514 20412
rect 3534 19934 3538 20412
rect 3558 19934 3562 20412
rect 3582 19934 3586 20412
rect 3606 19934 3610 20412
rect 3630 19934 3634 20412
rect 3654 19934 3658 20412
rect 3667 20405 3672 20412
rect 3678 20405 3682 20412
rect 3685 20411 3699 20412
rect 3677 20391 3682 20405
rect 3667 20381 3672 20391
rect 3677 20367 3682 20381
rect 3678 19934 3682 20367
rect 3691 20261 3696 20271
rect 3701 20247 3706 20261
rect 3691 20189 3696 20199
rect 3702 20189 3706 20247
rect 3701 20175 3706 20189
rect 3715 20185 3723 20189
rect 3709 20175 3715 20185
rect 3691 20141 3696 20151
rect 3701 20127 3706 20141
rect 3702 19934 3706 20127
rect 3715 20021 3720 20031
rect 3725 20007 3730 20021
rect 3726 19935 3730 20007
rect 3715 19934 3747 19935
rect 1987 19932 3747 19934
rect 1987 19925 1992 19932
rect 1997 19911 2002 19925
rect 1973 19695 1978 19709
rect 1963 19694 1997 19695
rect 1998 19694 2002 19911
rect 2022 19883 2026 19932
rect 2022 19835 2029 19883
rect 2022 19694 2026 19835
rect 2046 19694 2050 19932
rect 2070 19694 2074 19932
rect 2094 19694 2098 19932
rect 2107 19733 2112 19743
rect 2118 19733 2122 19932
rect 2117 19719 2122 19733
rect 2107 19709 2112 19719
rect 2117 19695 2122 19709
rect 2118 19694 2122 19695
rect 2142 19694 2146 19932
rect 2166 19694 2170 19932
rect 2190 19694 2194 19932
rect 2214 19694 2218 19932
rect 2238 19694 2242 19932
rect 2262 19694 2266 19932
rect 2286 19694 2290 19932
rect 2310 19694 2314 19932
rect 2334 19694 2338 19932
rect 2358 19694 2362 19932
rect 2382 19694 2386 19932
rect 2406 19694 2410 19932
rect 2430 19694 2434 19932
rect 2454 19694 2458 19932
rect 2478 19694 2482 19932
rect 2502 19694 2506 19932
rect 2526 19694 2530 19932
rect 2550 19694 2554 19932
rect 2574 19694 2578 19932
rect 2598 19694 2602 19932
rect 2622 19694 2626 19932
rect 2646 19694 2650 19932
rect 2670 19694 2674 19932
rect 2694 19694 2698 19932
rect 2718 19694 2722 19932
rect 2742 19694 2746 19932
rect 2766 19694 2770 19932
rect 2790 19694 2794 19932
rect 2814 19694 2818 19932
rect 2838 19694 2842 19932
rect 2862 19694 2866 19932
rect 2886 19694 2890 19932
rect 2910 19694 2914 19932
rect 2934 19694 2938 19932
rect 2958 19694 2962 19932
rect 2982 19694 2986 19932
rect 3006 19694 3010 19932
rect 3030 19694 3034 19932
rect 3054 19694 3058 19932
rect 3078 19694 3082 19932
rect 3102 19694 3106 19932
rect 3126 19694 3130 19932
rect 3150 19694 3154 19932
rect 3174 19694 3178 19932
rect 3198 19694 3202 19932
rect 3222 19694 3226 19932
rect 3246 19694 3250 19932
rect 3270 19694 3274 19932
rect 3294 19694 3298 19932
rect 3318 19694 3322 19932
rect 3342 19694 3346 19932
rect 3366 19694 3370 19932
rect 3390 19694 3394 19932
rect 3414 19694 3418 19932
rect 3438 19694 3442 19932
rect 3462 19694 3466 19932
rect 3486 19694 3490 19932
rect 3510 19694 3514 19932
rect 3534 19694 3538 19932
rect 3558 19694 3562 19932
rect 3582 19694 3586 19932
rect 3606 19694 3610 19932
rect 3630 19694 3634 19932
rect 3654 19694 3658 19932
rect 3678 19694 3682 19932
rect 3702 19694 3706 19932
rect 3715 19925 3720 19932
rect 3726 19925 3730 19932
rect 3733 19931 3747 19932
rect 3725 19911 3730 19925
rect 3715 19901 3720 19911
rect 3725 19887 3730 19901
rect 3726 19695 3730 19887
rect 3739 19781 3744 19791
rect 3749 19767 3754 19781
rect 3739 19709 3744 19719
rect 3750 19709 3754 19767
rect 3749 19695 3754 19709
rect 3763 19705 3771 19709
rect 3757 19695 3763 19705
rect 3715 19694 3749 19695
rect 1963 19692 3749 19694
rect 1963 19685 1968 19692
rect 1973 19671 1978 19685
rect 1974 19646 1978 19671
rect 1998 19646 2002 19692
rect 2022 19646 2026 19692
rect 2046 19646 2050 19692
rect 2070 19646 2074 19692
rect 2094 19646 2098 19692
rect 2118 19646 2122 19692
rect 2142 19667 2146 19692
rect -2393 19644 -2026 19646
rect -2021 19644 2139 19646
rect -2371 19550 -2366 19644
rect -2348 19550 -2343 19644
rect -2325 19582 -2320 19644
rect -2317 19642 -2309 19644
rect -2309 19622 -2301 19630
rect -2317 19614 -2309 19622
rect -2123 19617 -2116 19622
rect -2123 19615 -2092 19617
rect -2091 19616 -2087 19632
rect -2026 19624 -2021 19636
rect -2037 19620 -2021 19624
rect -2292 19613 -2087 19615
rect -2123 19611 -2116 19613
rect -2325 19574 -2317 19582
rect -2325 19554 -2320 19574
rect -2317 19566 -2309 19574
rect -2325 19550 -2317 19554
rect -2000 19550 -1992 19644
rect -1663 19642 -1655 19644
rect -1969 19616 -1932 19632
rect -1655 19622 -1647 19630
rect -1969 19613 -1680 19615
rect -1663 19614 -1655 19622
rect -1671 19574 -1663 19582
rect -1663 19566 -1655 19574
rect -1926 19550 -1892 19553
rect -1671 19550 -1663 19554
rect -1642 19550 -1637 19644
rect -1619 19550 -1614 19644
rect -1530 19550 -1526 19644
rect -1506 19550 -1502 19644
rect -1482 19550 -1478 19644
rect -1458 19550 -1454 19644
rect -1434 19550 -1430 19644
rect -1410 19550 -1406 19644
rect -1386 19550 -1382 19644
rect -1362 19550 -1358 19644
rect -1338 19550 -1334 19644
rect -1314 19550 -1310 19644
rect -1290 19550 -1286 19644
rect -1266 19550 -1262 19644
rect -1242 19550 -1238 19644
rect -1218 19550 -1214 19644
rect -1194 19550 -1190 19644
rect -1170 19550 -1166 19644
rect -1146 19550 -1142 19644
rect -1122 19550 -1118 19644
rect -1098 19550 -1094 19644
rect -1074 19550 -1070 19644
rect -1050 19550 -1046 19644
rect -1026 19550 -1022 19644
rect -1002 19550 -998 19644
rect -978 19550 -974 19644
rect -954 19550 -950 19644
rect -930 19550 -926 19644
rect -906 19550 -902 19644
rect -882 19550 -878 19644
rect -858 19550 -854 19644
rect -834 19550 -830 19644
rect -810 19550 -806 19644
rect -786 19550 -782 19644
rect -762 19550 -758 19644
rect -738 19550 -734 19644
rect -714 19550 -710 19644
rect -690 19550 -686 19644
rect -666 19550 -662 19644
rect -642 19550 -638 19644
rect -618 19550 -614 19644
rect -594 19550 -590 19644
rect -570 19550 -566 19644
rect -546 19550 -542 19644
rect -522 19550 -518 19644
rect -498 19550 -494 19644
rect -474 19550 -470 19644
rect -450 19550 -446 19644
rect -426 19550 -422 19644
rect -402 19550 -398 19644
rect -378 19550 -374 19644
rect -354 19550 -350 19644
rect -330 19550 -326 19644
rect -306 19550 -302 19644
rect -282 19550 -278 19644
rect -258 19550 -254 19644
rect -234 19550 -230 19644
rect -210 19550 -206 19644
rect -186 19550 -182 19644
rect -162 19550 -158 19644
rect -138 19550 -134 19644
rect -114 19550 -110 19644
rect -90 19550 -86 19644
rect -66 19550 -62 19644
rect -42 19550 -38 19644
rect -18 19550 -14 19644
rect 6 19550 10 19644
rect 30 19550 34 19644
rect 54 19550 58 19644
rect 78 19550 82 19644
rect 102 19550 106 19644
rect 126 19550 130 19644
rect 150 19550 154 19644
rect 174 19550 178 19644
rect 198 19550 202 19644
rect 222 19550 226 19644
rect 246 19550 250 19644
rect 270 19550 274 19644
rect 294 19550 298 19644
rect 318 19550 322 19644
rect 342 19550 346 19644
rect 366 19550 370 19644
rect 390 19550 394 19644
rect 414 19550 418 19644
rect 438 19550 442 19644
rect 462 19550 466 19644
rect 486 19550 490 19644
rect 510 19550 514 19644
rect 534 19550 538 19644
rect 558 19550 562 19644
rect 582 19550 586 19644
rect 606 19550 610 19644
rect 630 19550 634 19644
rect 654 19550 658 19644
rect 678 19550 682 19644
rect 702 19550 706 19644
rect 726 19550 730 19644
rect 750 19550 754 19644
rect 774 19550 778 19644
rect 798 19550 802 19644
rect 822 19550 826 19644
rect 846 19550 850 19644
rect 870 19550 874 19644
rect 894 19550 898 19644
rect 918 19550 922 19644
rect 942 19550 946 19644
rect 966 19550 970 19644
rect 990 19550 994 19644
rect 1014 19550 1018 19644
rect 1038 19550 1042 19644
rect 1062 19550 1066 19644
rect 1086 19550 1090 19644
rect 1110 19550 1114 19644
rect 1134 19550 1138 19644
rect 1158 19550 1162 19644
rect 1182 19550 1186 19644
rect 1206 19550 1210 19644
rect 1230 19550 1234 19644
rect 1254 19550 1258 19644
rect 1278 19550 1282 19644
rect 1302 19550 1306 19644
rect 1326 19550 1330 19644
rect 1350 19550 1354 19644
rect 1374 19550 1378 19644
rect 1387 19589 1392 19599
rect 1398 19589 1402 19644
rect 1397 19575 1402 19589
rect 1387 19565 1392 19575
rect 1397 19551 1402 19565
rect 1398 19550 1402 19551
rect 1422 19550 1426 19644
rect 1446 19550 1450 19644
rect 1470 19550 1474 19644
rect 1494 19550 1498 19644
rect 1518 19550 1522 19644
rect 1542 19550 1546 19644
rect 1566 19550 1570 19644
rect 1590 19550 1594 19644
rect 1614 19550 1618 19644
rect 1638 19550 1642 19644
rect 1662 19550 1666 19644
rect 1686 19550 1690 19644
rect 1710 19550 1714 19644
rect 1734 19550 1738 19644
rect 1758 19550 1762 19644
rect 1782 19550 1786 19644
rect 1806 19550 1810 19644
rect 1830 19550 1834 19644
rect 1854 19550 1858 19644
rect 1878 19550 1882 19644
rect 1902 19550 1906 19644
rect 1926 19550 1930 19644
rect 1950 19550 1954 19644
rect 1974 19550 1978 19644
rect 1998 19643 2002 19644
rect 1998 19595 2005 19643
rect 1998 19550 2002 19595
rect 2022 19550 2026 19644
rect 2046 19550 2050 19644
rect 2070 19550 2074 19644
rect 2094 19550 2098 19644
rect 2118 19550 2122 19644
rect 2125 19643 2139 19644
rect 2142 19619 2149 19667
rect 2142 19550 2146 19619
rect 2166 19550 2170 19692
rect 2190 19550 2194 19692
rect 2214 19550 2218 19692
rect 2238 19550 2242 19692
rect 2262 19550 2266 19692
rect 2286 19550 2290 19692
rect 2310 19550 2314 19692
rect 2334 19550 2338 19692
rect 2358 19550 2362 19692
rect 2382 19550 2386 19692
rect 2406 19550 2410 19692
rect 2430 19550 2434 19692
rect 2454 19550 2458 19692
rect 2478 19550 2482 19692
rect 2502 19550 2506 19692
rect 2526 19550 2530 19692
rect 2550 19550 2554 19692
rect 2574 19550 2578 19692
rect 2598 19550 2602 19692
rect 2622 19550 2626 19692
rect 2646 19550 2650 19692
rect 2670 19550 2674 19692
rect 2694 19550 2698 19692
rect 2718 19550 2722 19692
rect 2742 19550 2746 19692
rect 2766 19550 2770 19692
rect 2790 19550 2794 19692
rect 2814 19550 2818 19692
rect 2838 19550 2842 19692
rect 2862 19550 2866 19692
rect 2886 19550 2890 19692
rect 2910 19550 2914 19692
rect 2934 19550 2938 19692
rect 2958 19550 2962 19692
rect 2982 19550 2986 19692
rect 3006 19550 3010 19692
rect 3030 19550 3034 19692
rect 3054 19550 3058 19692
rect 3078 19550 3082 19692
rect 3102 19550 3106 19692
rect 3126 19550 3130 19692
rect 3150 19550 3154 19692
rect 3174 19550 3178 19692
rect 3198 19550 3202 19692
rect 3222 19550 3226 19692
rect 3246 19550 3250 19692
rect 3270 19550 3274 19692
rect 3294 19550 3298 19692
rect 3318 19550 3322 19692
rect 3342 19550 3346 19692
rect 3366 19550 3370 19692
rect 3390 19550 3394 19692
rect 3414 19550 3418 19692
rect 3438 19550 3442 19692
rect 3462 19550 3466 19692
rect 3486 19550 3490 19692
rect 3510 19550 3514 19692
rect 3534 19550 3538 19692
rect 3558 19550 3562 19692
rect 3582 19550 3586 19692
rect 3606 19550 3610 19692
rect 3630 19550 3634 19692
rect 3654 19550 3658 19692
rect 3678 19550 3682 19692
rect 3702 19550 3706 19692
rect 3715 19685 3720 19692
rect 3726 19685 3730 19692
rect 3725 19671 3730 19685
rect 3715 19637 3720 19647
rect 3725 19623 3730 19637
rect 3715 19565 3720 19575
rect 3726 19565 3730 19623
rect 3725 19551 3730 19565
rect 3739 19561 3747 19565
rect 3733 19551 3739 19561
rect 3715 19550 3747 19551
rect -2393 19548 3747 19550
rect -2371 19502 -2366 19548
rect -2348 19502 -2343 19548
rect -2325 19542 -2317 19548
rect -2053 19546 -1972 19548
rect -2325 19526 -2320 19542
rect -2317 19538 -2309 19542
rect -2069 19538 -2068 19539
rect -2309 19526 -2301 19538
rect -2069 19531 -2038 19538
rect -2069 19529 -2068 19531
rect -2000 19530 -1992 19546
rect -1926 19543 -1924 19548
rect -1916 19540 -1914 19543
rect -1671 19542 -1663 19548
rect -1982 19530 -1916 19539
rect -1663 19538 -1655 19542
rect -2325 19514 -2317 19526
rect -2068 19523 -2053 19529
rect -2027 19528 -1992 19530
rect -2076 19514 -2053 19521
rect -2011 19520 -2002 19528
rect -2000 19520 -1992 19528
rect -1655 19526 -1647 19538
rect -2003 19518 -1992 19520
rect -2325 19502 -2320 19514
rect -2317 19510 -2309 19514
rect -2309 19502 -2301 19510
rect -2015 19506 -2003 19518
rect -2000 19502 -1992 19518
rect -1972 19514 -1924 19521
rect -1862 19513 -1680 19522
rect -1671 19514 -1663 19526
rect -1663 19510 -1655 19514
rect -1976 19502 -1940 19503
rect -1655 19502 -1647 19510
rect -1642 19502 -1637 19548
rect -1619 19502 -1614 19548
rect -1530 19502 -1526 19548
rect -1506 19502 -1502 19548
rect -1482 19502 -1478 19548
rect -1458 19502 -1454 19548
rect -1434 19502 -1430 19548
rect -1410 19502 -1406 19548
rect -1386 19502 -1382 19548
rect -1362 19502 -1358 19548
rect -1338 19502 -1334 19548
rect -1314 19502 -1310 19548
rect -1290 19502 -1286 19548
rect -1266 19502 -1262 19548
rect -1242 19502 -1238 19548
rect -1218 19502 -1214 19548
rect -1194 19502 -1190 19548
rect -1170 19502 -1166 19548
rect -1146 19502 -1142 19548
rect -1122 19502 -1118 19548
rect -1098 19502 -1094 19548
rect -1074 19502 -1070 19548
rect -1050 19502 -1046 19548
rect -1026 19502 -1022 19548
rect -1002 19502 -998 19548
rect -978 19502 -974 19548
rect -954 19502 -950 19548
rect -930 19502 -926 19548
rect -906 19502 -902 19548
rect -882 19502 -878 19548
rect -858 19502 -854 19548
rect -834 19502 -830 19548
rect -810 19502 -806 19548
rect -786 19502 -782 19548
rect -762 19502 -758 19548
rect -738 19502 -734 19548
rect -714 19502 -710 19548
rect -690 19502 -686 19548
rect -666 19502 -662 19548
rect -642 19502 -638 19548
rect -618 19502 -614 19548
rect -594 19502 -590 19548
rect -570 19502 -566 19548
rect -546 19502 -542 19548
rect -522 19502 -518 19548
rect -498 19502 -494 19548
rect -474 19502 -470 19548
rect -450 19502 -446 19548
rect -426 19502 -422 19548
rect -402 19502 -398 19548
rect -378 19502 -374 19548
rect -354 19503 -350 19548
rect -365 19502 -331 19503
rect -2393 19500 -331 19502
rect -2371 19430 -2366 19500
rect -2348 19430 -2343 19500
rect -2325 19498 -2320 19500
rect -2309 19498 -2301 19500
rect -2325 19486 -2317 19498
rect -2325 19466 -2320 19486
rect -2317 19482 -2309 19486
rect -2325 19458 -2317 19466
rect -2060 19460 -2030 19463
rect -2325 19430 -2320 19458
rect -2317 19450 -2309 19458
rect -2060 19447 -2038 19458
rect -2033 19451 -2030 19460
rect -2028 19456 -2027 19460
rect -2068 19442 -2038 19445
rect -2000 19430 -1992 19500
rect -1655 19498 -1647 19500
rect -1671 19486 -1663 19498
rect -1663 19482 -1655 19486
rect -1912 19475 -1884 19477
rect -1852 19469 -1804 19473
rect -1844 19460 -1796 19463
rect -1671 19458 -1663 19466
rect -1844 19447 -1804 19458
rect -1663 19450 -1655 19458
rect -1852 19442 -1680 19446
rect -1642 19430 -1637 19500
rect -1619 19430 -1614 19500
rect -1530 19430 -1526 19500
rect -1506 19430 -1502 19500
rect -1482 19430 -1478 19500
rect -1458 19430 -1454 19500
rect -1434 19430 -1430 19500
rect -1410 19430 -1406 19500
rect -1386 19430 -1382 19500
rect -1362 19430 -1358 19500
rect -1338 19430 -1334 19500
rect -1314 19430 -1310 19500
rect -1290 19430 -1286 19500
rect -1266 19430 -1262 19500
rect -1242 19430 -1238 19500
rect -1218 19430 -1214 19500
rect -1194 19430 -1190 19500
rect -1170 19430 -1166 19500
rect -1146 19430 -1142 19500
rect -1122 19430 -1118 19500
rect -1098 19430 -1094 19500
rect -1074 19430 -1070 19500
rect -1050 19430 -1046 19500
rect -1026 19430 -1022 19500
rect -1002 19430 -998 19500
rect -978 19430 -974 19500
rect -954 19430 -950 19500
rect -930 19430 -926 19500
rect -906 19430 -902 19500
rect -893 19469 -888 19479
rect -882 19469 -878 19500
rect -883 19455 -878 19469
rect -882 19430 -878 19455
rect -858 19430 -854 19500
rect -834 19430 -830 19500
rect -810 19430 -806 19500
rect -786 19430 -782 19500
rect -762 19430 -758 19500
rect -738 19430 -734 19500
rect -714 19430 -710 19500
rect -690 19430 -686 19500
rect -666 19430 -662 19500
rect -642 19430 -638 19500
rect -618 19430 -614 19500
rect -594 19430 -590 19500
rect -570 19430 -566 19500
rect -546 19430 -542 19500
rect -522 19430 -518 19500
rect -498 19430 -494 19500
rect -474 19430 -470 19500
rect -450 19430 -446 19500
rect -426 19430 -422 19500
rect -402 19430 -398 19500
rect -378 19430 -374 19500
rect -365 19493 -360 19500
rect -354 19493 -350 19500
rect -355 19479 -350 19493
rect -365 19469 -360 19479
rect -355 19455 -350 19469
rect -354 19430 -350 19455
rect -330 19430 -326 19548
rect -306 19430 -302 19548
rect -282 19430 -278 19548
rect -258 19430 -254 19548
rect -234 19430 -230 19548
rect -210 19430 -206 19548
rect -197 19517 -192 19527
rect -186 19517 -182 19548
rect -187 19503 -182 19517
rect -197 19502 -163 19503
rect -162 19502 -158 19548
rect -138 19502 -134 19548
rect -114 19502 -110 19548
rect -90 19502 -86 19548
rect -66 19502 -62 19548
rect -42 19502 -38 19548
rect -18 19502 -14 19548
rect 6 19502 10 19548
rect 30 19502 34 19548
rect 54 19502 58 19548
rect 78 19502 82 19548
rect 102 19502 106 19548
rect 126 19502 130 19548
rect 150 19502 154 19548
rect 174 19502 178 19548
rect 198 19502 202 19548
rect 222 19502 226 19548
rect 246 19502 250 19548
rect 270 19502 274 19548
rect 294 19502 298 19548
rect 318 19502 322 19548
rect 342 19502 346 19548
rect 366 19502 370 19548
rect 390 19502 394 19548
rect 414 19502 418 19548
rect 438 19502 442 19548
rect 462 19502 466 19548
rect 486 19502 490 19548
rect 510 19502 514 19548
rect 534 19502 538 19548
rect 558 19502 562 19548
rect 582 19502 586 19548
rect 606 19502 610 19548
rect 630 19502 634 19548
rect 654 19502 658 19548
rect 678 19502 682 19548
rect 702 19502 706 19548
rect 726 19502 730 19548
rect 750 19502 754 19548
rect 774 19502 778 19548
rect 798 19502 802 19548
rect 822 19502 826 19548
rect 846 19502 850 19548
rect 870 19502 874 19548
rect 894 19502 898 19548
rect 918 19502 922 19548
rect 942 19502 946 19548
rect 966 19502 970 19548
rect 990 19502 994 19548
rect 1014 19502 1018 19548
rect 1038 19502 1042 19548
rect 1062 19502 1066 19548
rect 1086 19502 1090 19548
rect 1110 19502 1114 19548
rect 1134 19502 1138 19548
rect 1158 19502 1162 19548
rect 1182 19502 1186 19548
rect 1206 19502 1210 19548
rect 1230 19502 1234 19548
rect 1254 19502 1258 19548
rect 1278 19502 1282 19548
rect 1302 19502 1306 19548
rect 1326 19502 1330 19548
rect 1350 19502 1354 19548
rect 1374 19502 1378 19548
rect 1398 19502 1402 19548
rect 1422 19523 1426 19548
rect -197 19500 1419 19502
rect -197 19493 -192 19500
rect -187 19479 -182 19493
rect -186 19430 -182 19479
rect -162 19451 -158 19500
rect -2393 19428 -165 19430
rect -2371 19406 -2366 19428
rect -2348 19406 -2343 19428
rect -2325 19406 -2320 19428
rect -2309 19410 -2301 19420
rect -2068 19411 -2062 19416
rect -2317 19406 -2309 19410
rect -2060 19406 -2050 19411
rect -2000 19406 -1992 19428
rect -1806 19420 -1680 19426
rect -1854 19411 -1806 19416
rect -1655 19410 -1647 19420
rect -1972 19406 -1964 19407
rect -1958 19406 -1942 19408
rect -1844 19406 -1806 19409
rect -1663 19406 -1655 19410
rect -1642 19406 -1637 19428
rect -1619 19406 -1614 19428
rect -1530 19406 -1526 19428
rect -1506 19406 -1502 19428
rect -1482 19406 -1478 19428
rect -1458 19406 -1454 19428
rect -1434 19406 -1430 19428
rect -1410 19406 -1406 19428
rect -1386 19406 -1382 19428
rect -1362 19406 -1358 19428
rect -1338 19406 -1334 19428
rect -1314 19406 -1310 19428
rect -1290 19406 -1286 19428
rect -1266 19406 -1262 19428
rect -1242 19406 -1238 19428
rect -1218 19406 -1214 19428
rect -1194 19406 -1190 19428
rect -1170 19406 -1166 19428
rect -1146 19406 -1142 19428
rect -1122 19406 -1118 19428
rect -1098 19406 -1094 19428
rect -1074 19406 -1070 19428
rect -1050 19406 -1046 19428
rect -1026 19406 -1022 19428
rect -1002 19406 -998 19428
rect -978 19406 -974 19428
rect -954 19406 -950 19428
rect -930 19406 -926 19428
rect -906 19406 -902 19428
rect -882 19406 -878 19428
rect -858 19406 -854 19428
rect -834 19406 -830 19428
rect -810 19406 -806 19428
rect -786 19406 -782 19428
rect -762 19406 -758 19428
rect -738 19406 -734 19428
rect -714 19406 -710 19428
rect -690 19406 -686 19428
rect -666 19406 -662 19428
rect -642 19406 -638 19428
rect -618 19406 -614 19428
rect -594 19406 -590 19428
rect -570 19406 -566 19428
rect -546 19406 -542 19428
rect -522 19406 -518 19428
rect -498 19406 -494 19428
rect -474 19406 -470 19428
rect -450 19406 -446 19428
rect -426 19406 -422 19428
rect -402 19406 -398 19428
rect -378 19406 -374 19428
rect -354 19406 -350 19428
rect -330 19427 -326 19428
rect -2393 19404 -333 19406
rect -2371 19382 -2366 19404
rect -2348 19382 -2343 19404
rect -2325 19382 -2320 19404
rect -2060 19398 -2050 19404
rect -2309 19382 -2301 19392
rect -2060 19391 -2030 19398
rect -2000 19394 -1992 19404
rect -1972 19402 -1942 19404
rect -1958 19401 -1942 19402
rect -1844 19400 -1806 19404
rect -2068 19384 -2062 19391
rect -2062 19382 -2036 19384
rect -2393 19380 -2036 19382
rect -2030 19382 -2012 19384
rect -2004 19382 -1990 19394
rect -1844 19393 -1798 19398
rect -1806 19391 -1798 19393
rect -1854 19389 -1844 19391
rect -1854 19384 -1806 19389
rect -1864 19382 -1796 19383
rect -1655 19382 -1647 19392
rect -1642 19382 -1637 19404
rect -1619 19382 -1614 19404
rect -1530 19382 -1526 19404
rect -1506 19382 -1502 19404
rect -1482 19382 -1478 19404
rect -1458 19382 -1454 19404
rect -1434 19382 -1430 19404
rect -1410 19382 -1406 19404
rect -1386 19382 -1382 19404
rect -1362 19382 -1358 19404
rect -1338 19382 -1334 19404
rect -1314 19382 -1310 19404
rect -1290 19382 -1286 19404
rect -1266 19382 -1262 19404
rect -1242 19382 -1238 19404
rect -1218 19382 -1214 19404
rect -1194 19382 -1190 19404
rect -1170 19382 -1166 19404
rect -1146 19382 -1142 19404
rect -1122 19382 -1118 19404
rect -1098 19382 -1094 19404
rect -1074 19382 -1070 19404
rect -1050 19382 -1046 19404
rect -1026 19382 -1022 19404
rect -1002 19382 -998 19404
rect -978 19382 -974 19404
rect -954 19382 -950 19404
rect -930 19382 -926 19404
rect -906 19382 -902 19404
rect -882 19382 -878 19404
rect -858 19403 -854 19404
rect -2030 19380 -861 19382
rect -2371 19334 -2366 19380
rect -2348 19334 -2343 19380
rect -2325 19334 -2320 19380
rect -2317 19376 -2309 19380
rect -2060 19376 -2050 19380
rect -2060 19374 -2036 19376
rect -2060 19372 -2030 19374
rect -2292 19366 -2030 19372
rect -2092 19350 -2062 19352
rect -2094 19346 -2062 19350
rect -2000 19334 -1992 19380
rect -1844 19373 -1806 19380
rect -1663 19376 -1655 19380
rect -1844 19366 -1680 19372
rect -1854 19350 -1806 19352
rect -1854 19346 -1680 19350
rect -1979 19334 -1945 19336
rect -1642 19334 -1637 19380
rect -1619 19334 -1614 19380
rect -1530 19334 -1526 19380
rect -1506 19334 -1502 19380
rect -1482 19334 -1478 19380
rect -1458 19334 -1454 19380
rect -1434 19334 -1430 19380
rect -1410 19334 -1406 19380
rect -1386 19334 -1382 19380
rect -1362 19334 -1358 19380
rect -1338 19334 -1334 19380
rect -1314 19334 -1310 19380
rect -1290 19334 -1286 19380
rect -1266 19334 -1262 19380
rect -1242 19334 -1238 19380
rect -1218 19334 -1214 19380
rect -1194 19334 -1190 19380
rect -1170 19334 -1166 19380
rect -1146 19334 -1142 19380
rect -1122 19334 -1118 19380
rect -1098 19334 -1094 19380
rect -1074 19334 -1070 19380
rect -1050 19334 -1046 19380
rect -1026 19334 -1022 19380
rect -1002 19334 -998 19380
rect -978 19334 -974 19380
rect -954 19334 -950 19380
rect -930 19334 -926 19380
rect -906 19334 -902 19380
rect -882 19334 -878 19380
rect -875 19379 -861 19380
rect -858 19379 -851 19403
rect -858 19334 -854 19379
rect -834 19334 -830 19404
rect -810 19334 -806 19404
rect -786 19334 -782 19404
rect -762 19334 -758 19404
rect -738 19334 -734 19404
rect -714 19334 -710 19404
rect -690 19334 -686 19404
rect -666 19334 -662 19404
rect -642 19334 -638 19404
rect -618 19334 -614 19404
rect -594 19334 -590 19404
rect -570 19334 -566 19404
rect -546 19334 -542 19404
rect -522 19334 -518 19404
rect -498 19334 -494 19404
rect -474 19334 -470 19404
rect -450 19334 -446 19404
rect -426 19334 -422 19404
rect -402 19334 -398 19404
rect -378 19334 -374 19404
rect -354 19334 -350 19404
rect -347 19403 -333 19404
rect -330 19382 -323 19427
rect -306 19382 -302 19428
rect -282 19382 -278 19428
rect -258 19382 -254 19428
rect -234 19382 -230 19428
rect -210 19382 -206 19428
rect -186 19382 -182 19428
rect -179 19427 -165 19428
rect -162 19407 -155 19451
rect -173 19406 -139 19407
rect -179 19404 -139 19406
rect -179 19403 -165 19404
rect -162 19403 -155 19404
rect -173 19397 -168 19403
rect -162 19397 -158 19403
rect -163 19383 -158 19397
rect -173 19382 -139 19383
rect -138 19382 -134 19500
rect -114 19382 -110 19500
rect -90 19382 -86 19500
rect -66 19382 -62 19500
rect -42 19382 -38 19500
rect -18 19382 -14 19500
rect 6 19382 10 19500
rect 30 19382 34 19500
rect 54 19382 58 19500
rect 78 19382 82 19500
rect 102 19382 106 19500
rect 126 19382 130 19500
rect 150 19382 154 19500
rect 174 19382 178 19500
rect 198 19382 202 19500
rect 222 19382 226 19500
rect 246 19382 250 19500
rect 270 19382 274 19500
rect 294 19382 298 19500
rect 318 19382 322 19500
rect 342 19382 346 19500
rect 366 19382 370 19500
rect 390 19382 394 19500
rect 414 19382 418 19500
rect 438 19382 442 19500
rect 462 19382 466 19500
rect 486 19382 490 19500
rect 510 19382 514 19500
rect 534 19382 538 19500
rect 558 19382 562 19500
rect 582 19382 586 19500
rect 606 19382 610 19500
rect 630 19382 634 19500
rect 654 19382 658 19500
rect 678 19382 682 19500
rect 702 19382 706 19500
rect 726 19382 730 19500
rect 750 19382 754 19500
rect 774 19382 778 19500
rect 798 19382 802 19500
rect 822 19382 826 19500
rect 846 19382 850 19500
rect 870 19382 874 19500
rect 894 19382 898 19500
rect 918 19382 922 19500
rect 942 19382 946 19500
rect 966 19382 970 19500
rect 990 19382 994 19500
rect 1014 19382 1018 19500
rect 1038 19382 1042 19500
rect 1062 19382 1066 19500
rect 1086 19382 1090 19500
rect 1110 19382 1114 19500
rect 1134 19382 1138 19500
rect 1158 19382 1162 19500
rect 1182 19382 1186 19500
rect 1206 19382 1210 19500
rect 1230 19382 1234 19500
rect 1254 19382 1258 19500
rect 1278 19382 1282 19500
rect 1302 19382 1306 19500
rect 1326 19382 1330 19500
rect 1350 19382 1354 19500
rect 1374 19382 1378 19500
rect 1398 19382 1402 19500
rect 1405 19499 1419 19500
rect 1422 19478 1429 19523
rect 1446 19478 1450 19548
rect 1470 19478 1474 19548
rect 1494 19478 1498 19548
rect 1518 19478 1522 19548
rect 1542 19478 1546 19548
rect 1566 19478 1570 19548
rect 1590 19478 1594 19548
rect 1614 19478 1618 19548
rect 1638 19478 1642 19548
rect 1662 19478 1666 19548
rect 1686 19478 1690 19548
rect 1710 19478 1714 19548
rect 1734 19478 1738 19548
rect 1758 19478 1762 19548
rect 1782 19478 1786 19548
rect 1806 19478 1810 19548
rect 1830 19478 1834 19548
rect 1854 19478 1858 19548
rect 1878 19478 1882 19548
rect 1902 19478 1906 19548
rect 1926 19478 1930 19548
rect 1950 19478 1954 19548
rect 1974 19478 1978 19548
rect 1998 19478 2002 19548
rect 2022 19478 2026 19548
rect 2046 19478 2050 19548
rect 2070 19478 2074 19548
rect 2094 19478 2098 19548
rect 2118 19478 2122 19548
rect 2142 19478 2146 19548
rect 2166 19478 2170 19548
rect 2190 19478 2194 19548
rect 2214 19478 2218 19548
rect 2238 19478 2242 19548
rect 2262 19478 2266 19548
rect 2286 19478 2290 19548
rect 2310 19478 2314 19548
rect 2334 19478 2338 19548
rect 2358 19478 2362 19548
rect 2382 19478 2386 19548
rect 2406 19478 2410 19548
rect 2430 19478 2434 19548
rect 2454 19478 2458 19548
rect 2478 19478 2482 19548
rect 2502 19478 2506 19548
rect 2526 19478 2530 19548
rect 2550 19478 2554 19548
rect 2574 19478 2578 19548
rect 2598 19478 2602 19548
rect 2622 19478 2626 19548
rect 2646 19478 2650 19548
rect 2670 19478 2674 19548
rect 2694 19478 2698 19548
rect 2718 19478 2722 19548
rect 2742 19478 2746 19548
rect 2766 19478 2770 19548
rect 2790 19478 2794 19548
rect 2814 19478 2818 19548
rect 2838 19478 2842 19548
rect 2862 19478 2866 19548
rect 2886 19478 2890 19548
rect 2910 19478 2914 19548
rect 2934 19478 2938 19548
rect 2958 19478 2962 19548
rect 2982 19478 2986 19548
rect 3006 19478 3010 19548
rect 3030 19478 3034 19548
rect 3054 19478 3058 19548
rect 3078 19478 3082 19548
rect 3102 19478 3106 19548
rect 3126 19478 3130 19548
rect 3150 19478 3154 19548
rect 3174 19478 3178 19548
rect 3198 19478 3202 19548
rect 3222 19478 3226 19548
rect 3246 19478 3250 19548
rect 3270 19478 3274 19548
rect 3294 19478 3298 19548
rect 3318 19478 3322 19548
rect 3342 19478 3346 19548
rect 3366 19478 3370 19548
rect 3390 19478 3394 19548
rect 3414 19478 3418 19548
rect 3438 19478 3442 19548
rect 3462 19478 3466 19548
rect 3486 19478 3490 19548
rect 3510 19478 3514 19548
rect 3534 19478 3538 19548
rect 3558 19478 3562 19548
rect 3582 19478 3586 19548
rect 3606 19478 3610 19548
rect 3630 19478 3634 19548
rect 3654 19478 3658 19548
rect 3678 19478 3682 19548
rect 3702 19479 3706 19548
rect 3715 19541 3720 19548
rect 3733 19547 3747 19548
rect 3725 19527 3730 19541
rect 3715 19493 3720 19503
rect 3726 19493 3730 19527
rect 3725 19479 3730 19493
rect 3739 19489 3747 19493
rect 3733 19479 3739 19489
rect 3691 19478 3725 19479
rect 1405 19476 3725 19478
rect 1405 19475 1419 19476
rect 1422 19475 1429 19476
rect 1422 19382 1426 19475
rect 1446 19382 1450 19476
rect 1470 19382 1474 19476
rect 1494 19383 1498 19476
rect 1483 19382 1517 19383
rect -347 19380 1517 19382
rect -347 19379 -333 19380
rect -330 19379 -323 19380
rect -330 19334 -326 19379
rect -306 19334 -302 19380
rect -282 19334 -278 19380
rect -258 19334 -254 19380
rect -234 19334 -230 19380
rect -210 19334 -206 19380
rect -186 19334 -182 19380
rect -173 19373 -168 19380
rect -163 19359 -158 19373
rect -162 19334 -158 19359
rect -138 19334 -134 19380
rect -114 19334 -110 19380
rect -90 19334 -86 19380
rect -66 19334 -62 19380
rect -42 19334 -38 19380
rect -18 19334 -14 19380
rect 6 19334 10 19380
rect 30 19334 34 19380
rect 54 19334 58 19380
rect 78 19334 82 19380
rect 102 19334 106 19380
rect 126 19334 130 19380
rect 150 19334 154 19380
rect 174 19334 178 19380
rect 198 19334 202 19380
rect 222 19334 226 19380
rect 246 19334 250 19380
rect 270 19334 274 19380
rect 294 19334 298 19380
rect 318 19334 322 19380
rect 342 19334 346 19380
rect 366 19334 370 19380
rect 390 19334 394 19380
rect 414 19334 418 19380
rect 438 19334 442 19380
rect 462 19334 466 19380
rect 486 19334 490 19380
rect 510 19334 514 19380
rect 534 19334 538 19380
rect 558 19334 562 19380
rect 582 19334 586 19380
rect 606 19334 610 19380
rect 630 19334 634 19380
rect 654 19334 658 19380
rect 678 19334 682 19380
rect 702 19334 706 19380
rect 726 19334 730 19380
rect 750 19334 754 19380
rect 774 19334 778 19380
rect 798 19334 802 19380
rect 822 19334 826 19380
rect 846 19334 850 19380
rect 870 19334 874 19380
rect 894 19334 898 19380
rect 918 19334 922 19380
rect 942 19334 946 19380
rect 966 19334 970 19380
rect 990 19334 994 19380
rect 1014 19334 1018 19380
rect 1038 19334 1042 19380
rect 1062 19334 1066 19380
rect 1086 19334 1090 19380
rect 1110 19334 1114 19380
rect 1134 19334 1138 19380
rect 1158 19334 1162 19380
rect 1182 19334 1186 19380
rect 1206 19334 1210 19380
rect 1230 19334 1234 19380
rect 1254 19334 1258 19380
rect 1278 19334 1282 19380
rect 1302 19334 1306 19380
rect 1326 19334 1330 19380
rect 1350 19334 1354 19380
rect 1374 19334 1378 19380
rect 1398 19334 1402 19380
rect 1422 19334 1426 19380
rect 1446 19334 1450 19380
rect 1470 19334 1474 19380
rect 1483 19373 1488 19380
rect 1494 19373 1498 19380
rect 1493 19359 1498 19373
rect 1483 19349 1488 19359
rect 1493 19335 1498 19349
rect 1494 19334 1498 19335
rect 1518 19334 1522 19476
rect 1542 19334 1546 19476
rect 1566 19334 1570 19476
rect 1590 19334 1594 19476
rect 1614 19334 1618 19476
rect 1638 19334 1642 19476
rect 1662 19334 1666 19476
rect 1686 19334 1690 19476
rect 1710 19334 1714 19476
rect 1734 19334 1738 19476
rect 1758 19334 1762 19476
rect 1782 19334 1786 19476
rect 1806 19334 1810 19476
rect 1830 19334 1834 19476
rect 1854 19334 1858 19476
rect 1878 19334 1882 19476
rect 1902 19334 1906 19476
rect 1926 19334 1930 19476
rect 1950 19334 1954 19476
rect 1974 19334 1978 19476
rect 1998 19334 2002 19476
rect 2022 19334 2026 19476
rect 2046 19334 2050 19476
rect 2070 19334 2074 19476
rect 2094 19334 2098 19476
rect 2118 19334 2122 19476
rect 2142 19334 2146 19476
rect 2166 19334 2170 19476
rect 2190 19334 2194 19476
rect 2214 19334 2218 19476
rect 2238 19334 2242 19476
rect 2262 19334 2266 19476
rect 2286 19334 2290 19476
rect 2310 19334 2314 19476
rect 2334 19334 2338 19476
rect 2358 19334 2362 19476
rect 2382 19334 2386 19476
rect 2406 19334 2410 19476
rect 2430 19334 2434 19476
rect 2454 19334 2458 19476
rect 2478 19334 2482 19476
rect 2502 19334 2506 19476
rect 2526 19334 2530 19476
rect 2550 19334 2554 19476
rect 2574 19334 2578 19476
rect 2598 19334 2602 19476
rect 2622 19334 2626 19476
rect 2646 19334 2650 19476
rect 2670 19334 2674 19476
rect 2694 19334 2698 19476
rect 2718 19334 2722 19476
rect 2742 19334 2746 19476
rect 2766 19334 2770 19476
rect 2790 19334 2794 19476
rect 2814 19334 2818 19476
rect 2838 19334 2842 19476
rect 2862 19334 2866 19476
rect 2886 19334 2890 19476
rect 2910 19334 2914 19476
rect 2934 19334 2938 19476
rect 2958 19334 2962 19476
rect 2982 19334 2986 19476
rect 3006 19334 3010 19476
rect 3030 19334 3034 19476
rect 3054 19334 3058 19476
rect 3078 19334 3082 19476
rect 3102 19334 3106 19476
rect 3126 19334 3130 19476
rect 3150 19334 3154 19476
rect 3174 19334 3178 19476
rect 3198 19334 3202 19476
rect 3222 19334 3226 19476
rect 3246 19334 3250 19476
rect 3270 19334 3274 19476
rect 3294 19334 3298 19476
rect 3318 19334 3322 19476
rect 3342 19334 3346 19476
rect 3366 19334 3370 19476
rect 3390 19334 3394 19476
rect 3414 19334 3418 19476
rect 3438 19334 3442 19476
rect 3462 19334 3466 19476
rect 3486 19334 3490 19476
rect 3510 19334 3514 19476
rect 3534 19334 3538 19476
rect 3558 19334 3562 19476
rect 3582 19334 3586 19476
rect 3606 19334 3610 19476
rect 3630 19334 3634 19476
rect 3654 19334 3658 19476
rect 3678 19334 3682 19476
rect 3691 19469 3696 19476
rect 3702 19469 3706 19476
rect 3701 19455 3706 19469
rect 3691 19421 3696 19431
rect 3701 19407 3706 19421
rect 3691 19349 3696 19359
rect 3702 19349 3706 19407
rect 3701 19335 3706 19349
rect 3715 19345 3723 19349
rect 3709 19335 3715 19345
rect 3691 19334 3723 19335
rect -2393 19332 3723 19334
rect -2371 19286 -2366 19332
rect -2348 19286 -2343 19332
rect -2325 19286 -2320 19332
rect -2080 19331 -1906 19332
rect -2080 19330 -2036 19331
rect -2080 19324 -2054 19330
rect -2309 19316 -2301 19322
rect -2317 19306 -2309 19316
rect -2070 19315 -2040 19322
rect -2054 19307 -2040 19310
rect -2000 19305 -1992 19331
rect -1920 19330 -1906 19331
rect -1850 19324 -1846 19332
rect -1840 19324 -1792 19332
rect -1969 19312 -1966 19321
rect -1850 19317 -1802 19322
rect -1906 19315 -1802 19317
rect -1655 19316 -1647 19322
rect -1906 19314 -1850 19315
rect -1846 19307 -1802 19313
rect -1663 19306 -1655 19316
rect -1860 19305 -1798 19306
rect -2078 19298 -2070 19305
rect -2309 19288 -2301 19294
rect -2317 19286 -2309 19288
rect -2154 19286 -2145 19296
rect -2044 19295 -2040 19300
rect -2028 19298 -1945 19305
rect -1929 19298 -1794 19305
rect -2070 19288 -2040 19295
rect -2044 19286 -2028 19288
rect -2000 19286 -1992 19298
rect -1860 19297 -1798 19298
rect -1850 19288 -1802 19295
rect -1655 19288 -1647 19294
rect -1978 19286 -1942 19287
rect -1663 19286 -1655 19288
rect -1642 19286 -1637 19332
rect -1619 19286 -1614 19332
rect -1530 19286 -1526 19332
rect -1506 19286 -1502 19332
rect -1482 19286 -1478 19332
rect -1458 19286 -1454 19332
rect -1434 19286 -1430 19332
rect -1410 19286 -1406 19332
rect -1386 19286 -1382 19332
rect -1362 19286 -1358 19332
rect -1338 19286 -1334 19332
rect -1314 19286 -1310 19332
rect -1290 19286 -1286 19332
rect -1266 19286 -1262 19332
rect -1242 19286 -1238 19332
rect -1218 19286 -1214 19332
rect -1194 19286 -1190 19332
rect -1170 19286 -1166 19332
rect -1146 19286 -1142 19332
rect -1122 19286 -1118 19332
rect -1098 19286 -1094 19332
rect -1074 19286 -1070 19332
rect -1050 19286 -1046 19332
rect -1026 19286 -1022 19332
rect -1002 19286 -998 19332
rect -978 19286 -974 19332
rect -954 19286 -950 19332
rect -930 19286 -926 19332
rect -906 19286 -902 19332
rect -882 19286 -878 19332
rect -858 19286 -854 19332
rect -834 19286 -830 19332
rect -810 19286 -806 19332
rect -786 19286 -782 19332
rect -762 19286 -758 19332
rect -738 19286 -734 19332
rect -714 19286 -710 19332
rect -690 19286 -686 19332
rect -666 19286 -662 19332
rect -642 19286 -638 19332
rect -618 19286 -614 19332
rect -594 19286 -590 19332
rect -570 19286 -566 19332
rect -546 19286 -542 19332
rect -522 19286 -518 19332
rect -498 19286 -494 19332
rect -474 19286 -470 19332
rect -450 19286 -446 19332
rect -426 19286 -422 19332
rect -402 19286 -398 19332
rect -378 19286 -374 19332
rect -354 19286 -350 19332
rect -330 19286 -326 19332
rect -306 19286 -302 19332
rect -282 19286 -278 19332
rect -258 19286 -254 19332
rect -234 19286 -230 19332
rect -210 19286 -206 19332
rect -186 19286 -182 19332
rect -162 19286 -158 19332
rect -138 19331 -134 19332
rect -138 19286 -131 19331
rect -114 19286 -110 19332
rect -90 19286 -86 19332
rect -66 19286 -62 19332
rect -42 19286 -38 19332
rect -18 19286 -14 19332
rect 6 19286 10 19332
rect 30 19286 34 19332
rect 54 19286 58 19332
rect 78 19286 82 19332
rect 102 19286 106 19332
rect 126 19286 130 19332
rect 150 19286 154 19332
rect 174 19286 178 19332
rect 198 19286 202 19332
rect 222 19286 226 19332
rect 246 19286 250 19332
rect 270 19286 274 19332
rect 294 19286 298 19332
rect 318 19286 322 19332
rect 342 19286 346 19332
rect 366 19286 370 19332
rect 390 19286 394 19332
rect 414 19286 418 19332
rect 438 19286 442 19332
rect 462 19286 466 19332
rect 486 19286 490 19332
rect 510 19286 514 19332
rect 534 19286 538 19332
rect 558 19286 562 19332
rect 582 19286 586 19332
rect 606 19286 610 19332
rect 630 19286 634 19332
rect 654 19286 658 19332
rect 678 19286 682 19332
rect 702 19286 706 19332
rect 726 19286 730 19332
rect 750 19286 754 19332
rect 774 19286 778 19332
rect 798 19286 802 19332
rect 822 19286 826 19332
rect 846 19286 850 19332
rect 870 19286 874 19332
rect 894 19286 898 19332
rect 918 19286 922 19332
rect 942 19286 946 19332
rect 966 19286 970 19332
rect 990 19286 994 19332
rect 1014 19286 1018 19332
rect 1038 19286 1042 19332
rect 1062 19286 1066 19332
rect 1086 19286 1090 19332
rect 1110 19286 1114 19332
rect 1134 19286 1138 19332
rect 1158 19286 1162 19332
rect 1182 19286 1186 19332
rect 1206 19287 1210 19332
rect 1195 19286 1229 19287
rect -2393 19284 1229 19286
rect -2371 18843 -2366 19284
rect -2361 18863 -2353 18873
rect -2348 18863 -2343 19284
rect -2351 18847 -2343 18863
rect -2371 18817 -2363 18843
rect -2383 18645 -2376 18655
rect -2371 18645 -2366 18817
rect -2373 18634 -2366 18645
rect -2348 18634 -2343 18847
rect -2325 19246 -2320 19284
rect -2317 19278 -2309 19284
rect -2145 19280 -2138 19284
rect -2070 19280 -2054 19284
rect -2078 19271 -2054 19278
rect -2062 19246 -2032 19247
rect -2000 19246 -1992 19284
rect -1846 19280 -1802 19284
rect -1846 19270 -1792 19279
rect -1663 19278 -1655 19284
rect -1942 19248 -1937 19260
rect -1850 19257 -1822 19258
rect -1850 19253 -1802 19257
rect -2325 19238 -2317 19246
rect -2062 19244 -1961 19246
rect -2325 19218 -2320 19238
rect -2317 19230 -2309 19238
rect -2062 19231 -2040 19242
rect -2032 19237 -1961 19244
rect -1947 19238 -1942 19246
rect -1842 19244 -1794 19247
rect -2070 19226 -2022 19230
rect -2325 19206 -2317 19218
rect -2325 19189 -2320 19206
rect -2317 19202 -2309 19206
rect -2309 19190 -2301 19202
rect -2317 19189 -2309 19190
rect -2325 19177 -2317 19189
rect -2325 19160 -2320 19177
rect -2317 19174 -2309 19177
rect -2309 19162 -2301 19174
rect -2062 19163 -2032 19168
rect -2317 19160 -2309 19162
rect -2325 19148 -2317 19160
rect -2325 19129 -2320 19148
rect -2317 19146 -2309 19148
rect -2325 19119 -2317 19129
rect -2325 19100 -2320 19119
rect -2317 19113 -2309 19119
rect -2243 19102 -2221 19110
rect -2211 19102 -2201 19122
rect -2073 19102 -2065 19120
rect -2000 19102 -1992 19237
rect -1942 19236 -1937 19238
rect -1932 19228 -1927 19236
rect -1912 19233 -1896 19239
rect -1842 19231 -1802 19242
rect -1671 19238 -1663 19246
rect -1663 19230 -1655 19238
rect -1850 19226 -1680 19230
rect -1842 19204 -1837 19206
rect -1789 19204 -1680 19206
rect -1671 19202 -1663 19218
rect -1837 19195 -1789 19196
rect -1895 19181 -1878 19183
rect -1895 19180 -1864 19181
rect -1837 19180 -1794 19193
rect -1655 19190 -1647 19202
rect -1663 19186 -1655 19190
rect -1794 19170 -1789 19175
rect -1671 19174 -1663 19186
rect -1837 19168 -1794 19170
rect -1842 19166 -1837 19168
rect -1842 19163 -1794 19166
rect -1655 19162 -1647 19174
rect -1837 19150 -1794 19160
rect -1663 19158 -1655 19162
rect -1671 19146 -1663 19158
rect -1671 19118 -1663 19126
rect -1655 19118 -1647 19120
rect -1663 19110 -1647 19118
rect -1642 19110 -1637 19284
rect -1885 19102 -1877 19104
rect -1708 19102 -1672 19104
rect -2243 19101 -2213 19102
rect -2325 19091 -2317 19100
rect -2259 19095 -2211 19101
rect -2183 19095 -1877 19102
rect -1869 19095 -1758 19102
rect -1710 19096 -1672 19102
rect -1710 19095 -1692 19096
rect -2211 19091 -2201 19095
rect -2325 19071 -2320 19091
rect -2317 19084 -2309 19091
rect -2211 19084 -2198 19091
rect -2325 19063 -2317 19071
rect -2300 19064 -2292 19074
rect -2243 19065 -2228 19076
rect -2211 19068 -2181 19084
rect -2211 19065 -2201 19068
rect -2325 19043 -2320 19063
rect -2317 19055 -2309 19063
rect -2325 19035 -2317 19043
rect -2325 19015 -2320 19035
rect -2317 19027 -2309 19035
rect -2325 19006 -2317 19015
rect -2325 18987 -2320 19006
rect -2317 18999 -2309 19006
rect -2325 18978 -2317 18987
rect -2325 18958 -2320 18978
rect -2317 18971 -2309 18978
rect -2325 18950 -2317 18958
rect -2290 18951 -2282 19064
rect -2251 19054 -2240 19058
rect -2211 19054 -2181 19058
rect -2251 19051 -2181 19054
rect -2176 19044 -2173 19046
rect -2240 19037 -2173 19044
rect -2169 19039 -2163 19094
rect -2073 19058 -2065 19095
rect -2073 19054 -2043 19058
rect -2000 19054 -1992 19095
rect -1915 19064 -1907 19073
rect -1963 19058 -1955 19064
rect -1963 19054 -1915 19058
rect -1885 19054 -1877 19095
rect -1875 19090 -1869 19094
rect -1829 19072 -1781 19074
rect -1847 19068 -1781 19072
rect -1778 19068 -1771 19094
rect -1758 19087 -1710 19094
rect -1718 19080 -1710 19087
rect -1768 19070 -1760 19080
rect -1718 19078 -1700 19080
rect -2146 19051 -2135 19054
rect -2105 19051 -2043 19054
rect -2035 19051 -1989 19054
rect -1973 19051 -1915 19054
rect -1907 19051 -1854 19054
rect -2073 19049 -2043 19051
rect -2135 19037 -2105 19044
rect -2065 19042 -2043 19049
rect -2243 19026 -2240 19035
rect -2221 19029 -2213 19037
rect -2211 19029 -2208 19037
rect -2203 19030 -2173 19037
rect -2251 19019 -2240 19026
rect -2211 19026 -2203 19029
rect -2211 19019 -2181 19026
rect -2073 19019 -2043 19026
rect -2203 18996 -2173 19003
rect -2262 18978 -2240 18988
rect -2203 18987 -2176 18996
rect -2083 18985 -2075 18995
rect -2040 18985 -2035 18989
rect -2073 18973 -2043 18985
rect -2028 18973 -2023 18985
rect -2000 18978 -1992 19051
rect -1963 19048 -1955 19051
rect -1963 19047 -1915 19048
rect -1955 19037 -1907 19044
rect -1885 19040 -1877 19051
rect -1837 19046 -1828 19062
rect -1758 19055 -1750 19070
rect -1758 19054 -1692 19055
rect -1837 19044 -1833 19046
rect -1837 19042 -1835 19044
rect -1887 19037 -1851 19040
rect -1750 19037 -1702 19044
rect -1885 19032 -1877 19037
rect -1963 19019 -1915 19026
rect -1905 18987 -1897 19032
rect -1857 19014 -1851 19037
rect -1760 19029 -1758 19030
rect -1837 19019 -1789 19026
rect -1758 19020 -1750 19026
rect -1758 19019 -1710 19020
rect -1955 18984 -1915 18987
rect -1963 18978 -1962 18980
rect -2000 18975 -1981 18978
rect -1965 18975 -1962 18978
rect -1955 18978 -1907 18982
rect -1885 18978 -1877 18997
rect -1857 18984 -1851 18996
rect -1750 18992 -1702 18999
rect -1829 18984 -1789 18986
rect -1766 18982 -1760 18992
rect -1829 18978 -1781 18982
rect -1756 18978 -1740 18982
rect -1680 18978 -1672 19096
rect -1671 19090 -1663 19098
rect -1645 19094 -1637 19110
rect -1663 19082 -1655 19090
rect -1671 19062 -1663 19070
rect -1663 19054 -1655 19062
rect -1671 19034 -1663 19042
rect -1671 19018 -1669 19031
rect -1663 19026 -1655 19034
rect -1671 19006 -1663 19014
rect -1663 18998 -1655 19006
rect -1671 18978 -1663 18986
rect -1955 18975 -1837 18978
rect -1829 18975 -1740 18978
rect -2206 18965 -2176 18968
rect -2206 18962 -2203 18965
rect -2161 18963 -2145 18972
rect -2073 18970 -2065 18973
rect -2073 18969 -2043 18970
rect -2028 18969 -2012 18973
rect -2073 18962 -2065 18968
rect -2203 18961 -2176 18962
rect -2065 18961 -2043 18962
rect -2262 18955 -2232 18961
rect -2176 18955 -2173 18961
rect -2043 18955 -2035 18961
rect -2325 18930 -2320 18950
rect -2317 18942 -2309 18950
rect -2153 18949 -2146 18953
rect -2325 18922 -2317 18930
rect -2300 18926 -2292 18936
rect -2325 18902 -2320 18922
rect -2317 18914 -2309 18922
rect -2325 18894 -2317 18902
rect -2325 18874 -2320 18894
rect -2317 18886 -2309 18894
rect -2290 18893 -2282 18926
rect -2273 18922 -2264 18927
rect -2206 18922 -2176 18927
rect -2262 18915 -2232 18920
rect -2198 18911 -2176 18922
rect -2198 18897 -2176 18905
rect -2166 18889 -2158 18937
rect -2143 18933 -2136 18949
rect -2143 18922 -2113 18927
rect -2073 18922 -2065 18927
rect -2065 18920 -2043 18922
rect -2043 18915 -2035 18920
rect -2065 18894 -2043 18909
rect -2006 18893 -2004 18909
rect -2265 18879 -2260 18885
rect -2143 18879 -2113 18886
rect -2270 18878 -2240 18879
rect -2270 18875 -2265 18878
rect -2325 18866 -2317 18874
rect -2325 18846 -2320 18866
rect -2317 18858 -2309 18866
rect -2113 18863 -2105 18873
rect -2291 18851 -2270 18858
rect -2198 18856 -2168 18858
rect -2135 18857 -2105 18858
rect -2103 18857 -2095 18863
rect -2113 18856 -2105 18857
rect -2065 18856 -2035 18858
rect -2000 18856 -1992 18975
rect -1963 18968 -1960 18975
rect -1915 18971 -1905 18975
rect -1963 18967 -1955 18968
rect -1963 18961 -1915 18967
rect -1989 18934 -1973 18937
rect -1915 18934 -1907 18941
rect -1990 18899 -1989 18920
rect -1983 18856 -1981 18919
rect -1885 18910 -1877 18975
rect -1789 18970 -1778 18975
rect -1837 18967 -1829 18968
rect -1837 18961 -1789 18967
rect -1756 18966 -1740 18975
rect -1837 18951 -1829 18961
rect -1872 18932 -1867 18942
rect -1789 18934 -1781 18941
rect -1776 18934 -1769 18951
rect -1756 18944 -1750 18966
rect -1671 18962 -1669 18973
rect -1663 18970 -1655 18978
rect -1671 18950 -1663 18958
rect -1663 18942 -1655 18950
rect -1702 18932 -1696 18938
rect -1955 18908 -1915 18910
rect -1963 18906 -1955 18908
rect -1963 18899 -1915 18906
rect -1963 18891 -1955 18899
rect -1963 18890 -1915 18891
rect -1973 18884 -1965 18887
rect -1955 18884 -1907 18888
rect -1974 18881 -1907 18884
rect -1973 18877 -1965 18881
rect -1963 18877 -1960 18879
rect -1963 18873 -1915 18877
rect -1963 18865 -1955 18873
rect -1963 18861 -1915 18865
rect -1963 18858 -1955 18861
rect -2240 18851 -2206 18856
rect -2198 18851 -2143 18856
rect -2113 18851 -1981 18856
rect -1915 18851 -1907 18858
rect -2270 18846 -2266 18850
rect -2086 18847 -2070 18851
rect -2325 18838 -2317 18846
rect -2270 18839 -2240 18846
rect -2206 18839 -2176 18846
rect -2325 18818 -2320 18838
rect -2317 18830 -2309 18838
rect -2270 18834 -2266 18839
rect -2270 18830 -2266 18833
rect -2198 18830 -2176 18837
rect -2166 18830 -2158 18847
rect -2143 18839 -2113 18846
rect -2198 18821 -2168 18825
rect -2325 18810 -2317 18818
rect -2143 18816 -2136 18830
rect -2085 18825 -2060 18826
rect -2039 18825 -2035 18834
rect -2135 18818 -2105 18825
rect -2085 18818 -2035 18825
rect -2029 18818 -2025 18825
rect -2325 18797 -2320 18810
rect -2317 18802 -2309 18810
rect -2235 18800 -2232 18803
rect -2325 18771 -2317 18797
rect -2325 18762 -2320 18771
rect -2325 18754 -2317 18762
rect -2135 18754 -2119 18767
rect -2000 18759 -1992 18851
rect -1983 18833 -1981 18851
rect -1955 18833 -1915 18834
rect -1862 18830 -1857 18932
rect -1706 18928 -1702 18932
rect -1829 18916 -1789 18924
rect -1671 18922 -1663 18930
rect -1849 18908 -1842 18916
rect -1790 18908 -1781 18916
rect -1663 18914 -1655 18922
rect -1837 18899 -1829 18906
rect -1758 18899 -1732 18906
rect -1748 18890 -1732 18899
rect -1671 18894 -1663 18902
rect -1829 18881 -1781 18888
rect -1663 18886 -1655 18894
rect -1829 18875 -1789 18879
rect -1768 18876 -1760 18886
rect -1758 18875 -1750 18876
rect -1671 18866 -1663 18874
rect -1837 18863 -1780 18866
rect -1758 18860 -1748 18866
rect -1708 18860 -1690 18866
rect -1829 18851 -1781 18858
rect -1680 18849 -1672 18866
rect -1663 18858 -1655 18866
rect -1829 18840 -1791 18846
rect -1758 18840 -1710 18842
rect -1758 18833 -1692 18840
rect -1671 18838 -1663 18846
rect -1955 18822 -1907 18825
rect -1791 18822 -1781 18825
rect -1991 18818 -1839 18822
rect -1791 18818 -1780 18822
rect -1680 18815 -1672 18833
rect -1663 18830 -1655 18838
rect -1839 18805 -1791 18812
rect -1671 18810 -1663 18818
rect -1829 18799 -1791 18803
rect -1671 18800 -1669 18810
rect -1663 18802 -1655 18810
rect -1680 18784 -1672 18799
rect -1642 18784 -1637 19094
rect -1619 19044 -1614 19284
rect -1619 19018 -1611 19044
rect -1768 18768 -1760 18778
rect -1758 18761 -1710 18768
rect -2325 18734 -2320 18754
rect -2317 18746 -2306 18754
rect -2031 18751 -1992 18759
rect -1750 18757 -1710 18761
rect -1674 18756 -1663 18762
rect -2307 18738 -2306 18746
rect -2149 18749 -2135 18750
rect -2149 18745 -2119 18749
rect -2024 18740 -2021 18749
rect -2325 18726 -2317 18734
rect -2325 18678 -2320 18726
rect -2317 18718 -2306 18726
rect -2185 18724 -2169 18736
rect -2056 18733 -2040 18737
rect -2021 18733 -2008 18740
rect -2056 18722 -2054 18732
rect -2056 18721 -2048 18722
rect -2307 18682 -2306 18690
rect -2111 18689 -2054 18695
rect -2325 18670 -2314 18678
rect -2104 18671 -2101 18675
rect -2325 18650 -2320 18670
rect -2314 18662 -2306 18670
rect -2104 18668 -2101 18670
rect -2084 18668 -2054 18669
rect -2000 18668 -1992 18751
rect -1758 18750 -1750 18751
rect -1758 18749 -1749 18750
rect -1758 18748 -1710 18749
rect -1663 18746 -1658 18756
rect -1831 18738 -1783 18742
rect -1784 18725 -1783 18738
rect -1674 18728 -1663 18734
rect -1826 18723 -1796 18724
rect -1663 18718 -1658 18728
rect -1654 18724 -1647 18734
rect -1644 18710 -1637 18724
rect -1758 18692 -1750 18695
rect -1758 18689 -1710 18692
rect -1844 18677 -1828 18679
rect -1844 18676 -1792 18677
rect -1828 18675 -1792 18676
rect -1772 18675 -1758 18683
rect -1750 18680 -1702 18687
rect -1750 18672 -1710 18676
rect -1700 18672 -1692 18692
rect -1674 18684 -1665 18692
rect -1674 18672 -1666 18680
rect -1758 18668 -1710 18669
rect -2307 18654 -2306 18662
rect -2139 18658 -2123 18667
rect -2111 18662 -2016 18668
rect -2139 18651 -2111 18658
rect -2325 18642 -2314 18650
rect -2177 18644 -2161 18645
rect -2141 18644 -2119 18646
rect -2104 18644 -2101 18662
rect -2076 18651 -2046 18656
rect -2325 18634 -2320 18642
rect -2314 18634 -2306 18642
rect -2076 18640 -2054 18646
rect -2021 18643 -2016 18662
rect -2000 18662 -1818 18668
rect -1802 18662 -1776 18668
rect -1760 18662 -1710 18668
rect -1666 18664 -1658 18672
rect -2189 18634 -2175 18639
rect -2373 18632 -2175 18634
rect -2373 18631 -2359 18632
rect -2371 18494 -2366 18631
rect -2348 18579 -2343 18632
rect -2325 18622 -2320 18632
rect -2307 18626 -2306 18632
rect -2189 18631 -2175 18632
rect -2149 18630 -2119 18639
rect -2084 18638 -2036 18639
rect -2000 18638 -1992 18662
rect -1758 18660 -1710 18662
rect -1758 18658 -1755 18660
rect -1828 18651 -1792 18658
rect -1768 18649 -1760 18656
rect -1758 18651 -1757 18658
rect -1710 18657 -1702 18658
rect -1750 18651 -1702 18657
rect -1674 18656 -1665 18664
rect -1768 18646 -1764 18649
rect -1758 18646 -1755 18651
rect -1818 18638 -1789 18646
rect -1758 18639 -1754 18646
rect -1750 18641 -1710 18646
rect -1674 18644 -1666 18652
rect -1758 18638 -1692 18639
rect -2084 18636 -1692 18638
rect -1666 18636 -1658 18644
rect -2084 18633 -1690 18636
rect -2084 18630 -2054 18633
rect -2046 18631 -1710 18633
rect -2325 18614 -2314 18622
rect -2076 18621 -2046 18628
rect -2325 18594 -2320 18614
rect -2314 18606 -2306 18614
rect -2076 18613 -2054 18619
rect -2084 18609 -2054 18611
rect -2104 18606 -2054 18609
rect -2307 18598 -2306 18606
rect -2084 18603 -2054 18606
rect -2325 18580 -2314 18594
rect -2348 18555 -2341 18579
rect -2325 18564 -2320 18580
rect -2314 18578 -2309 18580
rect -2309 18566 -2298 18578
rect -2092 18575 -2060 18576
rect -2062 18570 -2060 18575
rect -2314 18564 -2309 18566
rect -2348 18494 -2343 18555
rect -2325 18552 -2314 18564
rect -2076 18560 -2062 18570
rect -2076 18554 -2046 18558
rect -2014 18557 -2003 18566
rect -2062 18552 -2046 18554
rect -2325 18536 -2320 18552
rect -2314 18550 -2309 18552
rect -2076 18551 -2062 18552
rect -2309 18538 -2298 18550
rect -2092 18545 -2076 18551
rect -2046 18545 -2026 18546
rect -2314 18536 -2309 18538
rect -2046 18536 -2042 18537
rect -2325 18524 -2314 18536
rect -2141 18532 -2134 18534
rect -2052 18532 -2046 18536
rect -2292 18527 -2111 18532
rect -2096 18530 -2046 18532
rect -2076 18527 -2046 18530
rect -2325 18494 -2320 18524
rect -2314 18522 -2309 18524
rect -2092 18510 -2062 18512
rect -2094 18506 -2062 18510
rect -2000 18494 -1992 18631
rect -1758 18630 -1710 18631
rect -1680 18628 -1665 18636
rect -1750 18621 -1702 18628
rect -1680 18624 -1672 18628
rect -1680 18619 -1666 18624
rect -1836 18615 -1820 18616
rect -1837 18611 -1820 18615
rect -1750 18613 -1710 18619
rect -1674 18616 -1666 18619
rect -1837 18604 -1789 18611
rect -1758 18610 -1710 18611
rect -1760 18607 -1692 18610
rect -1666 18608 -1658 18616
rect -1837 18603 -1820 18604
rect -1764 18603 -1692 18607
rect -1674 18603 -1665 18608
rect -1680 18600 -1665 18603
rect -1750 18584 -1702 18586
rect -1680 18576 -1672 18600
rect -1671 18580 -1666 18596
rect -1854 18575 -1806 18576
rect -1829 18560 -1806 18570
rect -1655 18568 -1650 18580
rect -1666 18564 -1655 18568
rect -1829 18554 -1798 18558
rect -1680 18557 -1672 18560
rect -1806 18552 -1798 18554
rect -1671 18552 -1666 18564
rect -1829 18551 -1806 18552
rect -1854 18549 -1829 18551
rect -1854 18545 -1806 18549
rect -1829 18533 -1806 18543
rect -1655 18540 -1650 18552
rect -1666 18536 -1655 18540
rect -1829 18527 -1680 18532
rect -1671 18524 -1666 18536
rect -1854 18510 -1806 18512
rect -1854 18506 -1680 18510
rect -1926 18494 -1892 18497
rect -1642 18494 -1637 18710
rect -1619 18708 -1614 19018
rect -1619 18634 -1612 18658
rect -1619 18494 -1614 18634
rect -1530 18494 -1526 19284
rect -1506 18494 -1502 19284
rect -1482 18494 -1478 19284
rect -1458 18494 -1454 19284
rect -1434 18494 -1430 19284
rect -1410 18494 -1406 19284
rect -1386 18494 -1382 19284
rect -1362 18494 -1358 19284
rect -1338 18494 -1334 19284
rect -1314 18494 -1310 19284
rect -1290 18494 -1286 19284
rect -1266 18494 -1262 19284
rect -1242 18494 -1238 19284
rect -1218 18494 -1214 19284
rect -1194 18494 -1190 19284
rect -1170 18494 -1166 19284
rect -1146 18494 -1142 19284
rect -1122 18494 -1118 19284
rect -1098 18494 -1094 19284
rect -1074 18494 -1070 19284
rect -1061 18557 -1056 18567
rect -1050 18557 -1046 19284
rect -1051 18543 -1046 18557
rect -1061 18533 -1056 18543
rect -1051 18519 -1046 18533
rect -1050 18494 -1046 18519
rect -1026 18494 -1022 19284
rect -1002 18494 -998 19284
rect -978 18494 -974 19284
rect -954 18494 -950 19284
rect -930 18494 -926 19284
rect -906 18494 -902 19284
rect -882 18494 -878 19284
rect -858 18494 -854 19284
rect -834 18494 -830 19284
rect -821 19109 -816 19119
rect -810 19109 -806 19284
rect -811 19095 -806 19109
rect -810 18494 -806 19095
rect -786 19043 -782 19284
rect -786 19019 -779 19043
rect -786 18494 -782 19019
rect -762 18494 -758 19284
rect -738 18494 -734 19284
rect -714 18494 -710 19284
rect -690 18494 -686 19284
rect -666 18494 -662 19284
rect -642 18494 -638 19284
rect -618 18494 -614 19284
rect -594 18494 -590 19284
rect -570 18494 -566 19284
rect -546 18494 -542 19284
rect -522 18494 -518 19284
rect -498 18494 -494 19284
rect -474 18494 -470 19284
rect -450 18494 -446 19284
rect -426 18494 -422 19284
rect -402 18494 -398 19284
rect -378 18494 -374 19284
rect -354 18494 -350 19284
rect -330 18494 -326 19284
rect -306 18494 -302 19284
rect -282 18494 -278 19284
rect -258 18494 -254 19284
rect -234 18494 -230 19284
rect -210 18494 -206 19284
rect -186 18494 -182 19284
rect -162 18494 -158 19284
rect -155 19283 -141 19284
rect -138 19283 -131 19284
rect -138 18494 -134 19283
rect -114 18494 -110 19284
rect -90 18494 -86 19284
rect -66 18494 -62 19284
rect -42 18494 -38 19284
rect -18 18494 -14 19284
rect 6 18494 10 19284
rect 30 18494 34 19284
rect 54 18494 58 19284
rect 78 18494 82 19284
rect 102 18494 106 19284
rect 126 18494 130 19284
rect 150 18494 154 19284
rect 174 18494 178 19284
rect 198 18494 202 19284
rect 222 18494 226 19284
rect 246 18494 250 19284
rect 270 18494 274 19284
rect 294 18494 298 19284
rect 318 18494 322 19284
rect 342 18494 346 19284
rect 366 18494 370 19284
rect 390 18494 394 19284
rect 414 18494 418 19284
rect 438 18494 442 19284
rect 462 18494 466 19284
rect 486 18494 490 19284
rect 510 18494 514 19284
rect 534 18494 538 19284
rect 558 18494 562 19284
rect 582 18494 586 19284
rect 606 18494 610 19284
rect 630 18494 634 19284
rect 654 18494 658 19284
rect 678 18494 682 19284
rect 702 18494 706 19284
rect 726 18494 730 19284
rect 750 18494 754 19284
rect 774 18494 778 19284
rect 798 18494 802 19284
rect 822 18494 826 19284
rect 846 18494 850 19284
rect 870 18494 874 19284
rect 894 18494 898 19284
rect 918 18494 922 19284
rect 942 18494 946 19284
rect 955 19253 960 19263
rect 966 19253 970 19284
rect 965 19239 970 19253
rect 955 19238 989 19239
rect 990 19238 994 19284
rect 1014 19238 1018 19284
rect 1038 19238 1042 19284
rect 1062 19238 1066 19284
rect 1086 19238 1090 19284
rect 1110 19238 1114 19284
rect 1134 19238 1138 19284
rect 1158 19238 1162 19284
rect 1182 19238 1186 19284
rect 1195 19277 1200 19284
rect 1206 19277 1210 19284
rect 1205 19263 1210 19277
rect 1195 19253 1200 19263
rect 1205 19239 1210 19253
rect 1206 19238 1210 19239
rect 1230 19238 1234 19332
rect 1254 19238 1258 19332
rect 1278 19238 1282 19332
rect 1302 19238 1306 19332
rect 1326 19238 1330 19332
rect 1350 19238 1354 19332
rect 1374 19238 1378 19332
rect 1398 19238 1402 19332
rect 1422 19238 1426 19332
rect 1446 19238 1450 19332
rect 1470 19238 1474 19332
rect 1494 19238 1498 19332
rect 1518 19307 1522 19332
rect 1518 19262 1525 19307
rect 1542 19262 1546 19332
rect 1566 19262 1570 19332
rect 1590 19262 1594 19332
rect 1614 19262 1618 19332
rect 1638 19262 1642 19332
rect 1662 19262 1666 19332
rect 1686 19262 1690 19332
rect 1710 19262 1714 19332
rect 1734 19262 1738 19332
rect 1758 19262 1762 19332
rect 1782 19262 1786 19332
rect 1806 19262 1810 19332
rect 1830 19262 1834 19332
rect 1854 19262 1858 19332
rect 1878 19262 1882 19332
rect 1902 19262 1906 19332
rect 1926 19262 1930 19332
rect 1950 19262 1954 19332
rect 1974 19262 1978 19332
rect 1998 19262 2002 19332
rect 2022 19262 2026 19332
rect 2046 19262 2050 19332
rect 2070 19262 2074 19332
rect 2094 19262 2098 19332
rect 2118 19262 2122 19332
rect 2142 19262 2146 19332
rect 2166 19262 2170 19332
rect 2190 19262 2194 19332
rect 2214 19262 2218 19332
rect 2238 19262 2242 19332
rect 2262 19262 2266 19332
rect 2286 19262 2290 19332
rect 2310 19262 2314 19332
rect 2334 19262 2338 19332
rect 2358 19262 2362 19332
rect 2382 19262 2386 19332
rect 2406 19262 2410 19332
rect 2430 19262 2434 19332
rect 2454 19262 2458 19332
rect 2478 19262 2482 19332
rect 2502 19262 2506 19332
rect 2526 19262 2530 19332
rect 2550 19262 2554 19332
rect 2574 19262 2578 19332
rect 2598 19262 2602 19332
rect 2622 19262 2626 19332
rect 2646 19262 2650 19332
rect 2670 19262 2674 19332
rect 2694 19262 2698 19332
rect 2718 19262 2722 19332
rect 2742 19262 2746 19332
rect 2766 19262 2770 19332
rect 2790 19262 2794 19332
rect 2814 19262 2818 19332
rect 2838 19262 2842 19332
rect 2862 19262 2866 19332
rect 2886 19262 2890 19332
rect 2910 19262 2914 19332
rect 2934 19262 2938 19332
rect 2958 19262 2962 19332
rect 2982 19262 2986 19332
rect 3006 19262 3010 19332
rect 3030 19262 3034 19332
rect 3054 19262 3058 19332
rect 3078 19262 3082 19332
rect 3102 19262 3106 19332
rect 3126 19262 3130 19332
rect 3150 19262 3154 19332
rect 3174 19262 3178 19332
rect 3198 19262 3202 19332
rect 3222 19262 3226 19332
rect 3246 19262 3250 19332
rect 3270 19262 3274 19332
rect 3294 19262 3298 19332
rect 3318 19262 3322 19332
rect 3342 19262 3346 19332
rect 3366 19262 3370 19332
rect 3390 19262 3394 19332
rect 3414 19262 3418 19332
rect 3438 19262 3442 19332
rect 3462 19262 3466 19332
rect 3486 19262 3490 19332
rect 3510 19262 3514 19332
rect 3534 19262 3538 19332
rect 3558 19262 3562 19332
rect 3582 19262 3586 19332
rect 3606 19262 3610 19332
rect 3630 19262 3634 19332
rect 3654 19262 3658 19332
rect 3678 19262 3682 19332
rect 3691 19325 3696 19332
rect 3709 19331 3723 19332
rect 3701 19311 3706 19325
rect 3702 19263 3706 19311
rect 3691 19262 3723 19263
rect 1501 19260 3723 19262
rect 1501 19259 1515 19260
rect 1518 19259 1525 19260
rect 1518 19238 1522 19259
rect 1542 19238 1546 19260
rect 1566 19238 1570 19260
rect 1590 19238 1594 19260
rect 1614 19238 1618 19260
rect 1638 19238 1642 19260
rect 1662 19238 1666 19260
rect 1686 19238 1690 19260
rect 1710 19238 1714 19260
rect 1734 19238 1738 19260
rect 1758 19238 1762 19260
rect 1782 19238 1786 19260
rect 1806 19238 1810 19260
rect 1830 19238 1834 19260
rect 1854 19238 1858 19260
rect 1878 19238 1882 19260
rect 1902 19238 1906 19260
rect 1926 19238 1930 19260
rect 1950 19238 1954 19260
rect 1974 19238 1978 19260
rect 1998 19238 2002 19260
rect 2022 19238 2026 19260
rect 2046 19238 2050 19260
rect 2070 19238 2074 19260
rect 2094 19238 2098 19260
rect 2118 19238 2122 19260
rect 2142 19238 2146 19260
rect 2166 19238 2170 19260
rect 2190 19238 2194 19260
rect 2214 19238 2218 19260
rect 2238 19238 2242 19260
rect 2262 19238 2266 19260
rect 2286 19238 2290 19260
rect 2310 19238 2314 19260
rect 2334 19238 2338 19260
rect 2358 19238 2362 19260
rect 2382 19238 2386 19260
rect 2406 19238 2410 19260
rect 2430 19238 2434 19260
rect 2454 19238 2458 19260
rect 2478 19238 2482 19260
rect 2502 19238 2506 19260
rect 2526 19238 2530 19260
rect 2550 19238 2554 19260
rect 2574 19238 2578 19260
rect 2598 19238 2602 19260
rect 2622 19238 2626 19260
rect 2646 19238 2650 19260
rect 2670 19238 2674 19260
rect 2694 19238 2698 19260
rect 2718 19238 2722 19260
rect 2742 19238 2746 19260
rect 2766 19238 2770 19260
rect 2790 19238 2794 19260
rect 2814 19238 2818 19260
rect 2838 19238 2842 19260
rect 2862 19238 2866 19260
rect 2886 19238 2890 19260
rect 2910 19238 2914 19260
rect 2934 19238 2938 19260
rect 2958 19238 2962 19260
rect 2982 19238 2986 19260
rect 3006 19238 3010 19260
rect 3030 19238 3034 19260
rect 3054 19238 3058 19260
rect 3078 19238 3082 19260
rect 3102 19238 3106 19260
rect 3126 19238 3130 19260
rect 3150 19238 3154 19260
rect 3174 19238 3178 19260
rect 3198 19238 3202 19260
rect 3222 19238 3226 19260
rect 3246 19238 3250 19260
rect 3270 19238 3274 19260
rect 3294 19238 3298 19260
rect 3318 19238 3322 19260
rect 3342 19238 3346 19260
rect 3366 19238 3370 19260
rect 3390 19238 3394 19260
rect 3414 19238 3418 19260
rect 3438 19238 3442 19260
rect 3462 19238 3466 19260
rect 3486 19238 3490 19260
rect 3510 19238 3514 19260
rect 3534 19238 3538 19260
rect 3558 19238 3562 19260
rect 3582 19238 3586 19260
rect 3606 19238 3610 19260
rect 3630 19238 3634 19260
rect 3654 19238 3658 19260
rect 3678 19239 3682 19260
rect 3691 19253 3696 19260
rect 3702 19253 3706 19260
rect 3709 19259 3723 19260
rect 3701 19239 3706 19253
rect 3715 19249 3723 19253
rect 3709 19239 3715 19249
rect 3667 19238 3701 19239
rect 955 19236 3701 19238
rect 955 19229 960 19236
rect 965 19215 970 19229
rect 966 18494 970 19215
rect 990 19187 994 19236
rect 990 19139 997 19187
rect 990 18494 994 19139
rect 1014 18494 1018 19236
rect 1038 18494 1042 19236
rect 1062 18494 1066 19236
rect 1086 18494 1090 19236
rect 1110 18494 1114 19236
rect 1134 18494 1138 19236
rect 1158 18494 1162 19236
rect 1182 18494 1186 19236
rect 1206 18494 1210 19236
rect 1230 19211 1234 19236
rect 1230 19163 1237 19211
rect 1230 18494 1234 19163
rect 1254 18494 1258 19236
rect 1278 18494 1282 19236
rect 1302 18494 1306 19236
rect 1326 18494 1330 19236
rect 1350 18494 1354 19236
rect 1374 18494 1378 19236
rect 1398 18494 1402 19236
rect 1422 18494 1426 19236
rect 1446 18494 1450 19236
rect 1470 18494 1474 19236
rect 1494 18494 1498 19236
rect 1518 18494 1522 19236
rect 1542 18494 1546 19236
rect 1566 18494 1570 19236
rect 1590 18494 1594 19236
rect 1614 18494 1618 19236
rect 1638 18494 1642 19236
rect 1662 18494 1666 19236
rect 1686 18494 1690 19236
rect 1710 18494 1714 19236
rect 1734 18494 1738 19236
rect 1758 18494 1762 19236
rect 1782 18494 1786 19236
rect 1806 18494 1810 19236
rect 1830 18494 1834 19236
rect 1854 18494 1858 19236
rect 1878 18494 1882 19236
rect 1902 18494 1906 19236
rect 1926 18494 1930 19236
rect 1950 18494 1954 19236
rect 1974 18494 1978 19236
rect 1998 18494 2002 19236
rect 2022 18494 2026 19236
rect 2046 18494 2050 19236
rect 2070 18494 2074 19236
rect 2094 18494 2098 19236
rect 2118 18494 2122 19236
rect 2142 18494 2146 19236
rect 2166 18494 2170 19236
rect 2190 18494 2194 19236
rect 2214 18494 2218 19236
rect 2238 18494 2242 19236
rect 2262 18494 2266 19236
rect 2286 18494 2290 19236
rect 2310 18494 2314 19236
rect 2334 18494 2338 19236
rect 2358 18494 2362 19236
rect 2382 18494 2386 19236
rect 2406 18494 2410 19236
rect 2430 18494 2434 19236
rect 2454 18494 2458 19236
rect 2478 18494 2482 19236
rect 2502 18494 2506 19236
rect 2526 18494 2530 19236
rect 2550 18494 2554 19236
rect 2574 18494 2578 19236
rect 2598 18494 2602 19236
rect 2622 18494 2626 19236
rect 2646 18494 2650 19236
rect 2670 18494 2674 19236
rect 2694 18494 2698 19236
rect 2718 18494 2722 19236
rect 2742 18494 2746 19236
rect 2766 18494 2770 19236
rect 2790 18494 2794 19236
rect 2814 18494 2818 19236
rect 2838 18494 2842 19236
rect 2862 18494 2866 19236
rect 2886 18494 2890 19236
rect 2910 18494 2914 19236
rect 2934 18494 2938 19236
rect 2958 18494 2962 19236
rect 2982 18494 2986 19236
rect 3006 18494 3010 19236
rect 3030 18494 3034 19236
rect 3054 18494 3058 19236
rect 3078 18494 3082 19236
rect 3102 18494 3106 19236
rect 3126 18494 3130 19236
rect 3150 18494 3154 19236
rect 3174 18494 3178 19236
rect 3198 18494 3202 19236
rect 3211 18533 3216 18543
rect 3222 18533 3226 19236
rect 3221 18519 3226 18533
rect 3211 18509 3216 18519
rect 3221 18495 3226 18509
rect 3222 18494 3226 18495
rect 3246 18494 3250 19236
rect 3270 18494 3274 19236
rect 3294 18494 3298 19236
rect 3318 18494 3322 19236
rect 3342 18494 3346 19236
rect 3366 18494 3370 19236
rect 3390 18494 3394 19236
rect 3414 18494 3418 19236
rect 3427 18701 3432 18711
rect 3438 18701 3442 19236
rect 3437 18687 3442 18701
rect 3427 18677 3432 18687
rect 3437 18663 3442 18677
rect 3438 18494 3442 18663
rect 3462 18635 3466 19236
rect 3462 18590 3469 18635
rect 3486 18590 3490 19236
rect 3510 18590 3514 19236
rect 3534 18590 3538 19236
rect 3558 18590 3562 19236
rect 3582 18590 3586 19236
rect 3606 18590 3610 19236
rect 3630 18590 3634 19236
rect 3643 18677 3648 18687
rect 3654 18677 3658 19236
rect 3667 19229 3672 19236
rect 3678 19229 3682 19236
rect 3677 19215 3682 19229
rect 3653 18663 3658 18677
rect 3643 18590 3675 18591
rect 3445 18588 3675 18590
rect 3445 18587 3459 18588
rect 3462 18587 3469 18588
rect 3462 18494 3466 18587
rect 3486 18494 3490 18588
rect 3510 18494 3514 18588
rect 3534 18494 3538 18588
rect 3558 18494 3562 18588
rect 3582 18494 3586 18588
rect 3606 18494 3610 18588
rect 3630 18494 3634 18588
rect 3643 18581 3648 18588
rect 3661 18587 3675 18588
rect 3653 18567 3658 18581
rect 3643 18509 3648 18519
rect 3654 18509 3658 18567
rect 3653 18495 3658 18509
rect 3667 18505 3675 18509
rect 3661 18495 3667 18505
rect 3643 18494 3675 18495
rect -2393 18492 3675 18494
rect -2371 18470 -2366 18492
rect -2348 18470 -2343 18492
rect -2325 18470 -2320 18492
rect -2054 18491 -1906 18492
rect -2054 18490 -2036 18491
rect -2309 18476 -2301 18486
rect -2317 18470 -2309 18476
rect -2068 18475 -2038 18482
rect -2000 18474 -1992 18491
rect -1920 18490 -1906 18491
rect -1846 18484 -1794 18492
rect -1852 18477 -1804 18482
rect -1902 18475 -1804 18477
rect -1655 18476 -1647 18486
rect -2000 18472 -1975 18474
rect -1902 18473 -1852 18475
rect -2025 18470 -1975 18472
rect -1846 18470 -1804 18473
rect -1663 18470 -1655 18476
rect -1642 18470 -1637 18492
rect -1619 18470 -1614 18492
rect -1530 18470 -1526 18492
rect -1506 18470 -1502 18492
rect -1482 18470 -1478 18492
rect -1458 18470 -1454 18492
rect -1434 18470 -1430 18492
rect -1410 18470 -1406 18492
rect -1386 18470 -1382 18492
rect -1362 18470 -1358 18492
rect -1338 18470 -1334 18492
rect -1314 18470 -1310 18492
rect -1290 18470 -1286 18492
rect -1266 18470 -1262 18492
rect -1242 18470 -1238 18492
rect -1218 18470 -1214 18492
rect -1194 18470 -1190 18492
rect -1170 18470 -1166 18492
rect -1146 18470 -1142 18492
rect -1122 18470 -1118 18492
rect -1098 18470 -1094 18492
rect -1074 18470 -1070 18492
rect -1050 18470 -1046 18492
rect -1026 18491 -1022 18492
rect -2393 18468 -1029 18470
rect -2371 18446 -2366 18468
rect -2348 18446 -2343 18468
rect -2325 18446 -2320 18468
rect -2054 18467 -2038 18468
rect -2000 18467 -1966 18468
rect -1846 18467 -1804 18468
rect -2000 18466 -1975 18467
rect -2076 18458 -2054 18465
rect -2309 18448 -2301 18458
rect -2044 18455 -2038 18460
rect -2028 18458 -2001 18465
rect -2054 18448 -2038 18455
rect -2015 18457 -2001 18458
rect -2015 18448 -2014 18457
rect -2317 18446 -2309 18448
rect -2044 18446 -2028 18448
rect -2000 18446 -1992 18466
rect -1982 18465 -1975 18466
rect -1862 18465 -1798 18466
rect -1985 18458 -1796 18465
rect -1862 18457 -1798 18458
rect -1852 18448 -1804 18455
rect -1655 18448 -1647 18458
rect -1976 18446 -1940 18447
rect -1663 18446 -1655 18448
rect -1642 18446 -1637 18468
rect -1619 18446 -1614 18468
rect -1530 18446 -1526 18468
rect -1506 18446 -1502 18468
rect -1482 18446 -1478 18468
rect -1458 18446 -1454 18468
rect -1434 18446 -1430 18468
rect -1410 18446 -1406 18468
rect -1386 18446 -1382 18468
rect -1362 18446 -1358 18468
rect -1338 18446 -1334 18468
rect -1314 18446 -1310 18468
rect -1290 18446 -1286 18468
rect -1266 18446 -1262 18468
rect -1242 18446 -1238 18468
rect -1218 18446 -1214 18468
rect -1194 18446 -1190 18468
rect -1170 18446 -1166 18468
rect -1146 18446 -1142 18468
rect -1122 18446 -1118 18468
rect -1098 18446 -1094 18468
rect -1074 18446 -1070 18468
rect -1050 18446 -1046 18468
rect -1043 18467 -1029 18468
rect -1026 18446 -1019 18491
rect -1002 18446 -998 18492
rect -978 18446 -974 18492
rect -954 18446 -950 18492
rect -930 18446 -926 18492
rect -906 18446 -902 18492
rect -882 18446 -878 18492
rect -858 18446 -854 18492
rect -834 18446 -830 18492
rect -810 18446 -806 18492
rect -786 18446 -782 18492
rect -762 18446 -758 18492
rect -738 18446 -734 18492
rect -714 18446 -710 18492
rect -690 18446 -686 18492
rect -666 18446 -662 18492
rect -642 18446 -638 18492
rect -618 18446 -614 18492
rect -594 18446 -590 18492
rect -570 18446 -566 18492
rect -546 18446 -542 18492
rect -522 18446 -518 18492
rect -498 18446 -494 18492
rect -474 18446 -470 18492
rect -450 18446 -446 18492
rect -426 18446 -422 18492
rect -402 18446 -398 18492
rect -378 18446 -374 18492
rect -354 18446 -350 18492
rect -330 18446 -326 18492
rect -306 18446 -302 18492
rect -282 18447 -278 18492
rect -293 18446 -259 18447
rect -2393 18444 -259 18446
rect -2371 18374 -2366 18444
rect -2348 18374 -2343 18444
rect -2325 18410 -2320 18444
rect -2317 18442 -2309 18444
rect -2076 18431 -2054 18438
rect -2325 18402 -2317 18410
rect -2060 18404 -2030 18407
rect -2325 18374 -2320 18402
rect -2317 18394 -2309 18402
rect -2060 18391 -2038 18402
rect -2033 18395 -2030 18404
rect -2028 18400 -2027 18404
rect -2068 18386 -2038 18389
rect -2000 18374 -1992 18444
rect -1846 18440 -1804 18444
rect -1663 18442 -1655 18444
rect -1846 18430 -1794 18439
rect -1912 18419 -1884 18421
rect -1852 18413 -1804 18417
rect -1844 18404 -1796 18407
rect -1671 18402 -1663 18410
rect -1844 18391 -1804 18402
rect -1663 18394 -1655 18402
rect -1852 18386 -1680 18390
rect -1642 18374 -1637 18444
rect -1619 18374 -1614 18444
rect -1530 18374 -1526 18444
rect -1506 18374 -1502 18444
rect -1482 18374 -1478 18444
rect -1458 18374 -1454 18444
rect -1434 18374 -1430 18444
rect -1410 18374 -1406 18444
rect -1386 18374 -1382 18444
rect -1362 18374 -1358 18444
rect -1338 18374 -1334 18444
rect -1314 18374 -1310 18444
rect -1290 18374 -1286 18444
rect -1266 18374 -1262 18444
rect -1242 18374 -1238 18444
rect -1218 18374 -1214 18444
rect -1194 18374 -1190 18444
rect -1170 18374 -1166 18444
rect -1146 18374 -1142 18444
rect -1122 18374 -1118 18444
rect -1098 18374 -1094 18444
rect -1074 18374 -1070 18444
rect -1050 18374 -1046 18444
rect -1043 18443 -1029 18444
rect -1026 18443 -1019 18444
rect -1026 18374 -1022 18443
rect -1002 18374 -998 18444
rect -978 18374 -974 18444
rect -954 18374 -950 18444
rect -930 18374 -926 18444
rect -906 18374 -902 18444
rect -882 18374 -878 18444
rect -858 18374 -854 18444
rect -834 18374 -830 18444
rect -810 18374 -806 18444
rect -786 18374 -782 18444
rect -773 18413 -768 18423
rect -762 18413 -758 18444
rect -763 18399 -758 18413
rect -762 18374 -758 18399
rect -738 18374 -734 18444
rect -714 18374 -710 18444
rect -690 18374 -686 18444
rect -666 18374 -662 18444
rect -642 18374 -638 18444
rect -618 18374 -614 18444
rect -594 18374 -590 18444
rect -570 18374 -566 18444
rect -546 18374 -542 18444
rect -522 18374 -518 18444
rect -498 18374 -494 18444
rect -474 18374 -470 18444
rect -450 18374 -446 18444
rect -426 18374 -422 18444
rect -402 18374 -398 18444
rect -378 18374 -374 18444
rect -354 18374 -350 18444
rect -330 18374 -326 18444
rect -306 18374 -302 18444
rect -293 18437 -288 18444
rect -282 18437 -278 18444
rect -283 18423 -278 18437
rect -282 18374 -278 18423
rect -258 18374 -254 18492
rect -234 18374 -230 18492
rect -210 18374 -206 18492
rect -186 18374 -182 18492
rect -162 18374 -158 18492
rect -138 18374 -134 18492
rect -114 18374 -110 18492
rect -90 18374 -86 18492
rect -66 18374 -62 18492
rect -42 18374 -38 18492
rect -18 18374 -14 18492
rect 6 18374 10 18492
rect 30 18374 34 18492
rect 54 18374 58 18492
rect 78 18374 82 18492
rect 102 18374 106 18492
rect 126 18374 130 18492
rect 150 18374 154 18492
rect 174 18374 178 18492
rect 198 18374 202 18492
rect 222 18374 226 18492
rect 246 18374 250 18492
rect 270 18374 274 18492
rect 294 18374 298 18492
rect 318 18374 322 18492
rect 342 18374 346 18492
rect 366 18374 370 18492
rect 390 18374 394 18492
rect 414 18374 418 18492
rect 438 18374 442 18492
rect 462 18374 466 18492
rect 486 18374 490 18492
rect 510 18374 514 18492
rect 534 18374 538 18492
rect 558 18374 562 18492
rect 582 18374 586 18492
rect 606 18374 610 18492
rect 630 18374 634 18492
rect 654 18374 658 18492
rect 678 18374 682 18492
rect 702 18374 706 18492
rect 726 18374 730 18492
rect 750 18374 754 18492
rect 774 18374 778 18492
rect 798 18374 802 18492
rect 822 18374 826 18492
rect 846 18374 850 18492
rect 870 18374 874 18492
rect 894 18374 898 18492
rect 918 18374 922 18492
rect 931 18461 936 18471
rect 942 18461 946 18492
rect 941 18447 946 18461
rect 942 18374 946 18447
rect 966 18395 970 18492
rect -2393 18372 963 18374
rect -2371 18350 -2366 18372
rect -2348 18350 -2343 18372
rect -2325 18350 -2320 18372
rect -2309 18354 -2301 18364
rect -2068 18355 -2062 18360
rect -2317 18350 -2309 18354
rect -2060 18350 -2050 18355
rect -2000 18350 -1992 18372
rect -1806 18364 -1680 18370
rect -1854 18355 -1806 18360
rect -1655 18354 -1647 18364
rect -1972 18350 -1964 18351
rect -1958 18350 -1942 18352
rect -1844 18350 -1806 18353
rect -1663 18350 -1655 18354
rect -1642 18350 -1637 18372
rect -1619 18350 -1614 18372
rect -1530 18350 -1526 18372
rect -1506 18350 -1502 18372
rect -1482 18350 -1478 18372
rect -1458 18351 -1454 18372
rect -1469 18350 -1435 18351
rect -2393 18348 -1435 18350
rect -2371 18326 -2366 18348
rect -2348 18326 -2343 18348
rect -2325 18326 -2320 18348
rect -2060 18342 -2050 18348
rect -2309 18326 -2301 18336
rect -2060 18335 -2030 18342
rect -2000 18338 -1992 18348
rect -1972 18346 -1942 18348
rect -1958 18345 -1942 18346
rect -1844 18344 -1806 18348
rect -2068 18328 -2062 18335
rect -2062 18326 -2036 18328
rect -2393 18324 -2036 18326
rect -2030 18326 -2012 18328
rect -2004 18326 -1990 18338
rect -1844 18337 -1798 18342
rect -1806 18335 -1798 18337
rect -1854 18333 -1844 18335
rect -1854 18328 -1806 18333
rect -1864 18326 -1796 18327
rect -1655 18326 -1647 18336
rect -1642 18326 -1637 18348
rect -1619 18326 -1614 18348
rect -1530 18326 -1526 18348
rect -1506 18326 -1502 18348
rect -1482 18326 -1478 18348
rect -1469 18341 -1464 18348
rect -1458 18341 -1454 18348
rect -1459 18327 -1454 18341
rect -1458 18326 -1454 18327
rect -1434 18326 -1430 18372
rect -1410 18326 -1406 18372
rect -1386 18326 -1382 18372
rect -1362 18326 -1358 18372
rect -1338 18326 -1334 18372
rect -1314 18326 -1310 18372
rect -1290 18326 -1286 18372
rect -1266 18326 -1262 18372
rect -1242 18326 -1238 18372
rect -1218 18326 -1214 18372
rect -1194 18326 -1190 18372
rect -1170 18326 -1166 18372
rect -1146 18326 -1142 18372
rect -1122 18327 -1118 18372
rect -1133 18326 -1099 18327
rect -2030 18324 -1099 18326
rect -2371 18278 -2366 18324
rect -2348 18278 -2343 18324
rect -2325 18278 -2320 18324
rect -2317 18320 -2309 18324
rect -2060 18320 -2050 18324
rect -2060 18318 -2036 18320
rect -2060 18316 -2030 18318
rect -2292 18310 -2030 18316
rect -2092 18294 -2062 18296
rect -2094 18290 -2062 18294
rect -2000 18278 -1992 18324
rect -1844 18317 -1806 18324
rect -1663 18320 -1655 18324
rect -1844 18310 -1680 18316
rect -1854 18294 -1806 18296
rect -1854 18290 -1680 18294
rect -1642 18278 -1637 18324
rect -1619 18278 -1614 18324
rect -1530 18278 -1526 18324
rect -1506 18278 -1502 18324
rect -1482 18278 -1478 18324
rect -1458 18278 -1454 18324
rect -1434 18278 -1430 18324
rect -1410 18278 -1406 18324
rect -1386 18278 -1382 18324
rect -1362 18278 -1358 18324
rect -1338 18278 -1334 18324
rect -1314 18278 -1310 18324
rect -1290 18278 -1286 18324
rect -1266 18278 -1262 18324
rect -1242 18278 -1238 18324
rect -1218 18278 -1214 18324
rect -1194 18278 -1190 18324
rect -1170 18278 -1166 18324
rect -1146 18278 -1142 18324
rect -1133 18317 -1128 18324
rect -1122 18317 -1118 18324
rect -1123 18303 -1118 18317
rect -1122 18278 -1118 18303
rect -1098 18278 -1094 18372
rect -1074 18278 -1070 18372
rect -1050 18278 -1046 18372
rect -1026 18278 -1022 18372
rect -1002 18278 -998 18372
rect -978 18278 -974 18372
rect -954 18278 -950 18372
rect -930 18278 -926 18372
rect -906 18278 -902 18372
rect -882 18278 -878 18372
rect -858 18278 -854 18372
rect -834 18278 -830 18372
rect -810 18278 -806 18372
rect -786 18278 -782 18372
rect -762 18278 -758 18372
rect -738 18347 -734 18372
rect -738 18323 -731 18347
rect -738 18278 -734 18323
rect -714 18278 -710 18372
rect -690 18278 -686 18372
rect -666 18278 -662 18372
rect -642 18278 -638 18372
rect -618 18278 -614 18372
rect -594 18278 -590 18372
rect -570 18278 -566 18372
rect -546 18278 -542 18372
rect -522 18278 -518 18372
rect -498 18278 -494 18372
rect -474 18278 -470 18372
rect -450 18278 -446 18372
rect -426 18278 -422 18372
rect -402 18278 -398 18372
rect -378 18278 -374 18372
rect -354 18278 -350 18372
rect -330 18278 -326 18372
rect -306 18278 -302 18372
rect -282 18278 -278 18372
rect -258 18371 -254 18372
rect -258 18347 -251 18371
rect -258 18278 -254 18347
rect -234 18278 -230 18372
rect -210 18278 -206 18372
rect -186 18278 -182 18372
rect -162 18278 -158 18372
rect -138 18278 -134 18372
rect -114 18278 -110 18372
rect -90 18278 -86 18372
rect -66 18278 -62 18372
rect -42 18278 -38 18372
rect -18 18278 -14 18372
rect 6 18278 10 18372
rect 30 18278 34 18372
rect 54 18278 58 18372
rect 78 18278 82 18372
rect 102 18278 106 18372
rect 126 18278 130 18372
rect 150 18278 154 18372
rect 174 18278 178 18372
rect 198 18278 202 18372
rect 222 18278 226 18372
rect 246 18278 250 18372
rect 270 18278 274 18372
rect 294 18278 298 18372
rect 318 18278 322 18372
rect 342 18278 346 18372
rect 366 18278 370 18372
rect 390 18278 394 18372
rect 414 18278 418 18372
rect 438 18278 442 18372
rect 462 18278 466 18372
rect 486 18278 490 18372
rect 510 18278 514 18372
rect 534 18278 538 18372
rect 558 18278 562 18372
rect 582 18278 586 18372
rect 606 18278 610 18372
rect 630 18278 634 18372
rect 654 18278 658 18372
rect 678 18278 682 18372
rect 702 18278 706 18372
rect 726 18278 730 18372
rect 750 18278 754 18372
rect 774 18278 778 18372
rect 798 18278 802 18372
rect 822 18278 826 18372
rect 846 18278 850 18372
rect 870 18278 874 18372
rect 894 18278 898 18372
rect 918 18278 922 18372
rect 942 18278 946 18372
rect 949 18371 963 18372
rect 966 18371 973 18395
rect 966 18278 970 18371
rect 990 18278 994 18492
rect 1014 18278 1018 18492
rect 1038 18278 1042 18492
rect 1062 18278 1066 18492
rect 1086 18278 1090 18492
rect 1110 18278 1114 18492
rect 1134 18278 1138 18492
rect 1158 18278 1162 18492
rect 1182 18278 1186 18492
rect 1206 18278 1210 18492
rect 1230 18278 1234 18492
rect 1254 18278 1258 18492
rect 1278 18278 1282 18492
rect 1302 18278 1306 18492
rect 1326 18278 1330 18492
rect 1350 18278 1354 18492
rect 1374 18278 1378 18492
rect 1398 18278 1402 18492
rect 1422 18278 1426 18492
rect 1446 18278 1450 18492
rect 1470 18278 1474 18492
rect 1494 18278 1498 18492
rect 1518 18278 1522 18492
rect 1542 18278 1546 18492
rect 1566 18278 1570 18492
rect 1590 18278 1594 18492
rect 1614 18278 1618 18492
rect 1638 18278 1642 18492
rect 1662 18278 1666 18492
rect 1686 18278 1690 18492
rect 1710 18278 1714 18492
rect 1734 18278 1738 18492
rect 1758 18278 1762 18492
rect 1782 18278 1786 18492
rect 1806 18278 1810 18492
rect 1830 18278 1834 18492
rect 1854 18278 1858 18492
rect 1878 18278 1882 18492
rect 1902 18278 1906 18492
rect 1926 18278 1930 18492
rect 1950 18278 1954 18492
rect 1974 18278 1978 18492
rect 1998 18278 2002 18492
rect 2022 18278 2026 18492
rect 2046 18278 2050 18492
rect 2070 18278 2074 18492
rect 2094 18278 2098 18492
rect 2118 18278 2122 18492
rect 2142 18278 2146 18492
rect 2166 18278 2170 18492
rect 2190 18278 2194 18492
rect 2214 18278 2218 18492
rect 2238 18278 2242 18492
rect 2262 18278 2266 18492
rect 2286 18278 2290 18492
rect 2310 18278 2314 18492
rect 2334 18278 2338 18492
rect 2358 18278 2362 18492
rect 2382 18278 2386 18492
rect 2406 18278 2410 18492
rect 2430 18278 2434 18492
rect 2454 18278 2458 18492
rect 2478 18278 2482 18492
rect 2502 18278 2506 18492
rect 2526 18278 2530 18492
rect 2550 18278 2554 18492
rect 2574 18278 2578 18492
rect 2598 18278 2602 18492
rect 2622 18278 2626 18492
rect 2646 18278 2650 18492
rect 2670 18278 2674 18492
rect 2694 18278 2698 18492
rect 2718 18278 2722 18492
rect 2742 18278 2746 18492
rect 2766 18278 2770 18492
rect 2790 18278 2794 18492
rect 2814 18278 2818 18492
rect 2838 18278 2842 18492
rect 2862 18278 2866 18492
rect 2886 18278 2890 18492
rect 2910 18278 2914 18492
rect 2934 18278 2938 18492
rect 2958 18278 2962 18492
rect 2982 18278 2986 18492
rect 3006 18278 3010 18492
rect 3030 18278 3034 18492
rect 3054 18278 3058 18492
rect 3078 18278 3082 18492
rect 3102 18278 3106 18492
rect 3126 18278 3130 18492
rect 3150 18278 3154 18492
rect 3174 18278 3178 18492
rect 3198 18278 3202 18492
rect 3222 18278 3226 18492
rect 3246 18467 3250 18492
rect 3246 18419 3253 18467
rect 3246 18278 3250 18419
rect 3270 18278 3274 18492
rect 3294 18278 3298 18492
rect 3318 18278 3322 18492
rect 3342 18278 3346 18492
rect 3366 18278 3370 18492
rect 3390 18278 3394 18492
rect 3414 18278 3418 18492
rect 3438 18278 3442 18492
rect 3462 18278 3466 18492
rect 3486 18278 3490 18492
rect 3510 18278 3514 18492
rect 3534 18278 3538 18492
rect 3558 18278 3562 18492
rect 3582 18278 3586 18492
rect 3606 18278 3610 18492
rect 3630 18278 3634 18492
rect 3643 18485 3648 18492
rect 3661 18491 3675 18492
rect 3653 18471 3658 18485
rect 3654 18278 3658 18471
rect 3667 18365 3672 18375
rect 3677 18351 3682 18365
rect 3678 18278 3682 18351
rect 3691 18278 3699 18279
rect -2393 18276 3699 18278
rect -2371 18254 -2366 18276
rect -2348 18254 -2343 18276
rect -2325 18254 -2320 18276
rect -2072 18274 -2036 18275
rect -2072 18268 -2054 18274
rect -2309 18260 -2301 18268
rect -2317 18254 -2309 18260
rect -2092 18259 -2062 18264
rect -2000 18255 -1992 18276
rect -1938 18275 -1906 18276
rect -1920 18274 -1906 18275
rect -1806 18268 -1680 18274
rect -1854 18259 -1806 18264
rect -1655 18260 -1647 18268
rect -1982 18255 -1966 18256
rect -2000 18254 -1966 18255
rect -1846 18254 -1806 18257
rect -1663 18254 -1655 18260
rect -1642 18254 -1637 18276
rect -1619 18254 -1614 18276
rect -1589 18254 -1555 18255
rect -2393 18252 -1555 18254
rect -2371 18230 -2366 18252
rect -2348 18230 -2343 18252
rect -2325 18230 -2320 18252
rect -2000 18250 -1966 18252
rect -2309 18232 -2301 18240
rect -2062 18239 -2054 18246
rect -2092 18232 -2084 18239
rect -2062 18232 -2026 18234
rect -2317 18230 -2309 18232
rect -2062 18230 -2012 18232
rect -2000 18230 -1992 18250
rect -1982 18249 -1966 18250
rect -1846 18248 -1806 18252
rect -1846 18241 -1798 18246
rect -1806 18239 -1798 18241
rect -1854 18237 -1846 18239
rect -1854 18232 -1806 18237
rect -1655 18232 -1647 18240
rect -1864 18230 -1796 18231
rect -1663 18230 -1655 18232
rect -1642 18230 -1637 18252
rect -1619 18230 -1614 18252
rect -1530 18230 -1526 18276
rect -1506 18230 -1502 18276
rect -1482 18230 -1478 18276
rect -1458 18230 -1454 18276
rect -1434 18275 -1430 18276
rect -1434 18251 -1427 18275
rect -1434 18230 -1430 18251
rect -1410 18230 -1406 18276
rect -1386 18230 -1382 18276
rect -1362 18230 -1358 18276
rect -1338 18230 -1334 18276
rect -1314 18230 -1310 18276
rect -1290 18230 -1286 18276
rect -1266 18230 -1262 18276
rect -1242 18230 -1238 18276
rect -1218 18230 -1214 18276
rect -1194 18230 -1190 18276
rect -1170 18230 -1166 18276
rect -1146 18230 -1142 18276
rect -1122 18230 -1118 18276
rect -1098 18251 -1094 18276
rect -2393 18228 -1101 18230
rect -2371 18182 -2366 18228
rect -2348 18182 -2343 18228
rect -2325 18182 -2320 18228
rect -2317 18224 -2309 18228
rect -2062 18224 -2054 18228
rect -2154 18220 -2138 18222
rect -2057 18220 -2054 18224
rect -2292 18214 -2054 18220
rect -2052 18214 -2044 18224
rect -2092 18198 -2062 18200
rect -2094 18194 -2062 18198
rect -2000 18182 -1992 18228
rect -1846 18221 -1806 18228
rect -1663 18224 -1655 18228
rect -1846 18214 -1680 18220
rect -1854 18198 -1806 18200
rect -1854 18194 -1680 18198
rect -1642 18182 -1637 18228
rect -1619 18182 -1614 18228
rect -1530 18182 -1526 18228
rect -1506 18182 -1502 18228
rect -1482 18182 -1478 18228
rect -1458 18182 -1454 18228
rect -1434 18182 -1430 18228
rect -1410 18182 -1406 18228
rect -1386 18182 -1382 18228
rect -1362 18182 -1358 18228
rect -1338 18182 -1334 18228
rect -1314 18182 -1310 18228
rect -1290 18182 -1286 18228
rect -1266 18182 -1262 18228
rect -1242 18182 -1238 18228
rect -1218 18182 -1214 18228
rect -1194 18182 -1190 18228
rect -1170 18182 -1166 18228
rect -1146 18182 -1142 18228
rect -1122 18182 -1118 18228
rect -1115 18227 -1101 18228
rect -1098 18227 -1091 18251
rect -1098 18182 -1094 18227
rect -1074 18182 -1070 18276
rect -1061 18221 -1056 18231
rect -1050 18221 -1046 18276
rect -1051 18207 -1046 18221
rect -1050 18182 -1046 18207
rect -1026 18182 -1022 18276
rect -1002 18182 -998 18276
rect -978 18182 -974 18276
rect -954 18182 -950 18276
rect -930 18182 -926 18276
rect -906 18182 -902 18276
rect -882 18182 -878 18276
rect -858 18182 -854 18276
rect -834 18182 -830 18276
rect -810 18182 -806 18276
rect -786 18182 -782 18276
rect -762 18182 -758 18276
rect -738 18182 -734 18276
rect -714 18182 -710 18276
rect -690 18182 -686 18276
rect -666 18182 -662 18276
rect -642 18182 -638 18276
rect -618 18182 -614 18276
rect -594 18182 -590 18276
rect -570 18182 -566 18276
rect -546 18182 -542 18276
rect -522 18182 -518 18276
rect -498 18182 -494 18276
rect -474 18182 -470 18276
rect -450 18182 -446 18276
rect -426 18182 -422 18276
rect -402 18182 -398 18276
rect -378 18182 -374 18276
rect -354 18182 -350 18276
rect -330 18182 -326 18276
rect -306 18182 -302 18276
rect -282 18182 -278 18276
rect -258 18182 -254 18276
rect -234 18182 -230 18276
rect -210 18182 -206 18276
rect -186 18182 -182 18276
rect -162 18182 -158 18276
rect -138 18182 -134 18276
rect -114 18182 -110 18276
rect -90 18182 -86 18276
rect -66 18182 -62 18276
rect -42 18182 -38 18276
rect -18 18182 -14 18276
rect 6 18182 10 18276
rect 30 18182 34 18276
rect 54 18182 58 18276
rect 78 18182 82 18276
rect 102 18182 106 18276
rect 126 18182 130 18276
rect 150 18182 154 18276
rect 174 18182 178 18276
rect 198 18182 202 18276
rect 222 18182 226 18276
rect 246 18182 250 18276
rect 270 18182 274 18276
rect 294 18182 298 18276
rect 318 18182 322 18276
rect 342 18182 346 18276
rect 366 18182 370 18276
rect 390 18182 394 18276
rect 414 18182 418 18276
rect 438 18182 442 18276
rect 462 18182 466 18276
rect 486 18182 490 18276
rect 510 18182 514 18276
rect 534 18182 538 18276
rect 558 18182 562 18276
rect 582 18182 586 18276
rect 606 18182 610 18276
rect 630 18182 634 18276
rect 654 18182 658 18276
rect 678 18182 682 18276
rect 702 18182 706 18276
rect 726 18182 730 18276
rect 750 18182 754 18276
rect 774 18182 778 18276
rect 798 18182 802 18276
rect 822 18182 826 18276
rect 846 18182 850 18276
rect 870 18182 874 18276
rect 894 18182 898 18276
rect 918 18182 922 18276
rect 942 18182 946 18276
rect 966 18182 970 18276
rect 990 18182 994 18276
rect 1014 18182 1018 18276
rect 1038 18182 1042 18276
rect 1062 18182 1066 18276
rect 1086 18182 1090 18276
rect 1110 18182 1114 18276
rect 1134 18182 1138 18276
rect 1158 18182 1162 18276
rect 1182 18182 1186 18276
rect 1206 18182 1210 18276
rect 1230 18182 1234 18276
rect 1254 18182 1258 18276
rect 1278 18182 1282 18276
rect 1302 18182 1306 18276
rect 1326 18182 1330 18276
rect 1350 18182 1354 18276
rect 1374 18182 1378 18276
rect 1398 18182 1402 18276
rect 1422 18182 1426 18276
rect 1446 18182 1450 18276
rect 1470 18182 1474 18276
rect 1494 18182 1498 18276
rect 1518 18182 1522 18276
rect 1542 18182 1546 18276
rect 1566 18182 1570 18276
rect 1590 18182 1594 18276
rect 1614 18182 1618 18276
rect 1638 18182 1642 18276
rect 1662 18182 1666 18276
rect 1686 18182 1690 18276
rect 1710 18182 1714 18276
rect 1734 18182 1738 18276
rect 1758 18182 1762 18276
rect 1782 18182 1786 18276
rect 1806 18182 1810 18276
rect 1830 18182 1834 18276
rect 1854 18182 1858 18276
rect 1878 18182 1882 18276
rect 1902 18182 1906 18276
rect 1926 18182 1930 18276
rect 1950 18182 1954 18276
rect 1974 18182 1978 18276
rect 1998 18182 2002 18276
rect 2022 18182 2026 18276
rect 2046 18182 2050 18276
rect 2070 18182 2074 18276
rect 2094 18182 2098 18276
rect 2118 18182 2122 18276
rect 2142 18182 2146 18276
rect 2166 18182 2170 18276
rect 2190 18182 2194 18276
rect 2214 18182 2218 18276
rect 2238 18182 2242 18276
rect 2262 18182 2266 18276
rect 2286 18182 2290 18276
rect 2310 18182 2314 18276
rect 2334 18182 2338 18276
rect 2358 18182 2362 18276
rect 2382 18182 2386 18276
rect 2406 18182 2410 18276
rect 2430 18182 2434 18276
rect 2454 18182 2458 18276
rect 2478 18182 2482 18276
rect 2502 18182 2506 18276
rect 2526 18182 2530 18276
rect 2550 18182 2554 18276
rect 2574 18182 2578 18276
rect 2598 18182 2602 18276
rect 2622 18182 2626 18276
rect 2646 18182 2650 18276
rect 2670 18182 2674 18276
rect 2694 18182 2698 18276
rect 2718 18182 2722 18276
rect 2742 18182 2746 18276
rect 2766 18182 2770 18276
rect 2790 18182 2794 18276
rect 2814 18182 2818 18276
rect 2838 18182 2842 18276
rect 2862 18182 2866 18276
rect 2886 18182 2890 18276
rect 2910 18182 2914 18276
rect 2934 18182 2938 18276
rect 2958 18182 2962 18276
rect 2982 18182 2986 18276
rect 3006 18182 3010 18276
rect 3030 18182 3034 18276
rect 3054 18182 3058 18276
rect 3078 18182 3082 18276
rect 3102 18182 3106 18276
rect 3126 18182 3130 18276
rect 3150 18182 3154 18276
rect 3174 18182 3178 18276
rect 3198 18182 3202 18276
rect 3222 18182 3226 18276
rect 3246 18182 3250 18276
rect 3270 18182 3274 18276
rect 3294 18182 3298 18276
rect 3318 18182 3322 18276
rect 3342 18182 3346 18276
rect 3366 18182 3370 18276
rect 3390 18182 3394 18276
rect 3414 18182 3418 18276
rect 3438 18182 3442 18276
rect 3462 18182 3466 18276
rect 3486 18182 3490 18276
rect 3510 18182 3514 18276
rect 3534 18182 3538 18276
rect 3558 18182 3562 18276
rect 3582 18182 3586 18276
rect 3606 18182 3610 18276
rect 3630 18182 3634 18276
rect 3654 18182 3658 18276
rect 3678 18182 3682 18276
rect 3685 18275 3699 18276
rect 3691 18269 3696 18275
rect 3701 18255 3706 18269
rect 3702 18182 3706 18255
rect 3715 18182 3723 18183
rect -2393 18180 3723 18182
rect -2371 18158 -2366 18180
rect -2348 18158 -2343 18180
rect -2325 18158 -2320 18180
rect -2072 18178 -2036 18179
rect -2072 18172 -2054 18178
rect -2309 18164 -2301 18172
rect -2317 18158 -2309 18164
rect -2092 18163 -2062 18168
rect -2000 18159 -1992 18180
rect -1938 18179 -1906 18180
rect -1920 18178 -1906 18179
rect -1806 18172 -1680 18178
rect -1854 18163 -1806 18168
rect -1655 18164 -1647 18172
rect -1982 18159 -1966 18160
rect -2000 18158 -1966 18159
rect -1846 18158 -1806 18161
rect -1663 18158 -1655 18164
rect -1642 18158 -1637 18180
rect -1619 18158 -1614 18180
rect -1554 18166 -1547 18179
rect -2393 18156 -1557 18158
rect -2371 18134 -2366 18156
rect -2348 18134 -2343 18156
rect -2325 18134 -2320 18156
rect -2000 18154 -1966 18156
rect -2309 18136 -2301 18144
rect -2062 18143 -2054 18150
rect -2092 18136 -2084 18143
rect -2062 18136 -2026 18138
rect -2317 18134 -2309 18136
rect -2062 18134 -2012 18136
rect -2000 18134 -1992 18154
rect -1982 18153 -1966 18154
rect -1846 18152 -1806 18156
rect -1846 18145 -1798 18150
rect -1806 18143 -1798 18145
rect -1854 18141 -1846 18143
rect -1854 18136 -1806 18141
rect -1655 18136 -1647 18144
rect -1864 18134 -1796 18135
rect -1663 18134 -1655 18136
rect -1642 18134 -1637 18156
rect -1619 18134 -1614 18156
rect -1571 18155 -1557 18156
rect -1554 18155 -1547 18156
rect -1530 18134 -1526 18180
rect -1506 18134 -1502 18180
rect -1482 18134 -1478 18180
rect -1469 18149 -1464 18159
rect -1458 18149 -1454 18180
rect -1459 18135 -1454 18149
rect -1458 18134 -1454 18135
rect -1434 18134 -1430 18180
rect -1410 18134 -1406 18180
rect -1386 18134 -1382 18180
rect -1362 18134 -1358 18180
rect -1338 18134 -1334 18180
rect -1314 18134 -1310 18180
rect -1290 18134 -1286 18180
rect -1266 18134 -1262 18180
rect -1242 18134 -1238 18180
rect -1218 18134 -1214 18180
rect -1194 18134 -1190 18180
rect -1170 18134 -1166 18180
rect -1146 18134 -1142 18180
rect -1122 18134 -1118 18180
rect -1098 18134 -1094 18180
rect -1074 18134 -1070 18180
rect -1050 18134 -1046 18180
rect -1026 18155 -1022 18180
rect -2393 18132 -1029 18134
rect -2371 18086 -2366 18132
rect -2348 18086 -2343 18132
rect -2325 18086 -2320 18132
rect -2317 18128 -2309 18132
rect -2062 18128 -2054 18132
rect -2154 18124 -2138 18126
rect -2057 18124 -2054 18128
rect -2292 18118 -2054 18124
rect -2052 18118 -2044 18128
rect -2092 18102 -2062 18104
rect -2094 18098 -2062 18102
rect -2000 18086 -1992 18132
rect -1846 18125 -1806 18132
rect -1663 18128 -1655 18132
rect -1846 18118 -1680 18124
rect -1854 18102 -1806 18104
rect -1854 18098 -1680 18102
rect -1642 18086 -1637 18132
rect -1619 18086 -1614 18132
rect -1530 18086 -1526 18132
rect -1506 18086 -1502 18132
rect -1482 18086 -1478 18132
rect -1458 18086 -1454 18132
rect -1434 18086 -1430 18132
rect -1410 18086 -1406 18132
rect -1386 18086 -1382 18132
rect -1362 18086 -1358 18132
rect -1338 18086 -1334 18132
rect -1314 18086 -1310 18132
rect -1290 18086 -1286 18132
rect -1266 18086 -1262 18132
rect -1242 18086 -1238 18132
rect -1218 18086 -1214 18132
rect -1194 18086 -1190 18132
rect -1170 18086 -1166 18132
rect -1146 18086 -1142 18132
rect -1122 18086 -1118 18132
rect -1098 18086 -1094 18132
rect -1074 18086 -1070 18132
rect -1050 18086 -1046 18132
rect -1043 18131 -1029 18132
rect -1026 18131 -1019 18155
rect -1026 18086 -1022 18131
rect -1002 18086 -998 18180
rect -978 18086 -974 18180
rect -954 18086 -950 18180
rect -930 18086 -926 18180
rect -906 18086 -902 18180
rect -882 18086 -878 18180
rect -858 18086 -854 18180
rect -834 18086 -830 18180
rect -810 18086 -806 18180
rect -786 18086 -782 18180
rect -762 18086 -758 18180
rect -738 18086 -734 18180
rect -725 18125 -720 18135
rect -714 18125 -710 18180
rect -715 18111 -710 18125
rect -714 18086 -710 18111
rect -690 18086 -686 18180
rect -666 18086 -662 18180
rect -642 18086 -638 18180
rect -618 18086 -614 18180
rect -594 18086 -590 18180
rect -570 18086 -566 18180
rect -546 18086 -542 18180
rect -522 18086 -518 18180
rect -498 18086 -494 18180
rect -474 18086 -470 18180
rect -450 18086 -446 18180
rect -426 18086 -422 18180
rect -402 18086 -398 18180
rect -378 18086 -374 18180
rect -354 18086 -350 18180
rect -330 18086 -326 18180
rect -306 18086 -302 18180
rect -282 18086 -278 18180
rect -258 18086 -254 18180
rect -234 18086 -230 18180
rect -210 18086 -206 18180
rect -186 18086 -182 18180
rect -162 18086 -158 18180
rect -138 18086 -134 18180
rect -114 18086 -110 18180
rect -90 18086 -86 18180
rect -66 18086 -62 18180
rect -42 18086 -38 18180
rect -18 18086 -14 18180
rect 6 18086 10 18180
rect 30 18086 34 18180
rect 54 18086 58 18180
rect 78 18086 82 18180
rect 102 18086 106 18180
rect 126 18086 130 18180
rect 150 18086 154 18180
rect 174 18086 178 18180
rect 198 18086 202 18180
rect 222 18086 226 18180
rect 246 18086 250 18180
rect 270 18086 274 18180
rect 294 18086 298 18180
rect 318 18086 322 18180
rect 342 18086 346 18180
rect 366 18086 370 18180
rect 390 18086 394 18180
rect 414 18086 418 18180
rect 438 18086 442 18180
rect 462 18086 466 18180
rect 486 18086 490 18180
rect 510 18086 514 18180
rect 534 18086 538 18180
rect 558 18086 562 18180
rect 582 18086 586 18180
rect 606 18086 610 18180
rect 630 18086 634 18180
rect 654 18086 658 18180
rect 678 18086 682 18180
rect 702 18086 706 18180
rect 726 18086 730 18180
rect 750 18086 754 18180
rect 774 18086 778 18180
rect 798 18086 802 18180
rect 822 18086 826 18180
rect 846 18086 850 18180
rect 870 18086 874 18180
rect 894 18086 898 18180
rect 918 18086 922 18180
rect 942 18086 946 18180
rect 966 18086 970 18180
rect 990 18086 994 18180
rect 1014 18086 1018 18180
rect 1038 18086 1042 18180
rect 1062 18086 1066 18180
rect 1086 18086 1090 18180
rect 1110 18086 1114 18180
rect 1134 18086 1138 18180
rect 1158 18086 1162 18180
rect 1182 18086 1186 18180
rect 1206 18086 1210 18180
rect 1230 18086 1234 18180
rect 1254 18086 1258 18180
rect 1278 18086 1282 18180
rect 1302 18086 1306 18180
rect 1326 18086 1330 18180
rect 1350 18086 1354 18180
rect 1374 18086 1378 18180
rect 1398 18086 1402 18180
rect 1422 18086 1426 18180
rect 1446 18086 1450 18180
rect 1470 18086 1474 18180
rect 1494 18086 1498 18180
rect 1518 18086 1522 18180
rect 1542 18086 1546 18180
rect 1566 18086 1570 18180
rect 1590 18086 1594 18180
rect 1614 18086 1618 18180
rect 1638 18086 1642 18180
rect 1662 18086 1666 18180
rect 1686 18086 1690 18180
rect 1710 18086 1714 18180
rect 1734 18086 1738 18180
rect 1758 18086 1762 18180
rect 1782 18086 1786 18180
rect 1806 18086 1810 18180
rect 1830 18086 1834 18180
rect 1854 18086 1858 18180
rect 1878 18086 1882 18180
rect 1902 18086 1906 18180
rect 1926 18086 1930 18180
rect 1950 18086 1954 18180
rect 1974 18086 1978 18180
rect 1998 18086 2002 18180
rect 2022 18086 2026 18180
rect 2046 18086 2050 18180
rect 2070 18086 2074 18180
rect 2094 18086 2098 18180
rect 2118 18086 2122 18180
rect 2142 18086 2146 18180
rect 2166 18086 2170 18180
rect 2190 18086 2194 18180
rect 2214 18086 2218 18180
rect 2238 18086 2242 18180
rect 2262 18086 2266 18180
rect 2286 18086 2290 18180
rect 2310 18086 2314 18180
rect 2334 18086 2338 18180
rect 2358 18086 2362 18180
rect 2382 18086 2386 18180
rect 2406 18086 2410 18180
rect 2430 18086 2434 18180
rect 2454 18086 2458 18180
rect 2478 18086 2482 18180
rect 2502 18086 2506 18180
rect 2526 18086 2530 18180
rect 2550 18086 2554 18180
rect 2574 18086 2578 18180
rect 2598 18086 2602 18180
rect 2622 18086 2626 18180
rect 2646 18086 2650 18180
rect 2670 18086 2674 18180
rect 2694 18086 2698 18180
rect 2718 18086 2722 18180
rect 2742 18086 2746 18180
rect 2766 18086 2770 18180
rect 2790 18086 2794 18180
rect 2814 18086 2818 18180
rect 2838 18086 2842 18180
rect 2862 18086 2866 18180
rect 2886 18086 2890 18180
rect 2910 18086 2914 18180
rect 2934 18086 2938 18180
rect 2958 18086 2962 18180
rect 2982 18086 2986 18180
rect 3006 18086 3010 18180
rect 3030 18086 3034 18180
rect 3054 18086 3058 18180
rect 3078 18086 3082 18180
rect 3102 18086 3106 18180
rect 3126 18086 3130 18180
rect 3150 18086 3154 18180
rect 3174 18086 3178 18180
rect 3198 18086 3202 18180
rect 3222 18086 3226 18180
rect 3246 18086 3250 18180
rect 3270 18086 3274 18180
rect 3294 18086 3298 18180
rect 3318 18086 3322 18180
rect 3342 18086 3346 18180
rect 3366 18086 3370 18180
rect 3390 18086 3394 18180
rect 3414 18086 3418 18180
rect 3438 18086 3442 18180
rect 3462 18086 3466 18180
rect 3486 18086 3490 18180
rect 3510 18086 3514 18180
rect 3534 18086 3538 18180
rect 3558 18086 3562 18180
rect 3582 18086 3586 18180
rect 3606 18086 3610 18180
rect 3630 18086 3634 18180
rect 3654 18086 3658 18180
rect 3678 18086 3682 18180
rect 3702 18086 3706 18180
rect 3709 18179 3723 18180
rect 3715 18173 3720 18179
rect 3725 18159 3730 18173
rect 3726 18086 3730 18159
rect 3739 18086 3747 18087
rect -2393 18084 3747 18086
rect -2371 18062 -2366 18084
rect -2348 18062 -2343 18084
rect -2325 18062 -2320 18084
rect -2072 18082 -2036 18083
rect -2072 18076 -2054 18082
rect -2309 18068 -2301 18076
rect -2317 18062 -2309 18068
rect -2092 18067 -2062 18072
rect -2000 18063 -1992 18084
rect -1938 18083 -1906 18084
rect -1920 18082 -1906 18083
rect -1806 18076 -1680 18082
rect -1854 18067 -1806 18072
rect -1655 18068 -1647 18076
rect -1982 18063 -1966 18064
rect -2000 18062 -1966 18063
rect -1846 18062 -1806 18065
rect -1663 18062 -1655 18068
rect -1642 18062 -1637 18084
rect -1619 18062 -1614 18084
rect -1530 18062 -1526 18084
rect -1506 18062 -1502 18084
rect -1482 18062 -1478 18084
rect -1458 18062 -1454 18084
rect -1434 18083 -1430 18084
rect -2393 18060 -1437 18062
rect -2371 18038 -2366 18060
rect -2348 18038 -2343 18060
rect -2325 18038 -2320 18060
rect -2000 18058 -1966 18060
rect -2309 18040 -2301 18048
rect -2062 18047 -2054 18054
rect -2092 18040 -2084 18047
rect -2062 18040 -2026 18042
rect -2317 18038 -2309 18040
rect -2062 18038 -2012 18040
rect -2000 18038 -1992 18058
rect -1982 18057 -1966 18058
rect -1846 18056 -1806 18060
rect -1846 18049 -1798 18054
rect -1806 18047 -1798 18049
rect -1854 18045 -1846 18047
rect -1854 18040 -1806 18045
rect -1655 18040 -1647 18048
rect -1864 18038 -1796 18039
rect -1663 18038 -1655 18040
rect -1642 18038 -1637 18060
rect -1619 18038 -1614 18060
rect -1530 18038 -1526 18060
rect -1506 18038 -1502 18060
rect -1482 18038 -1478 18060
rect -1458 18038 -1454 18060
rect -1451 18059 -1437 18060
rect -1434 18059 -1427 18083
rect -1434 18038 -1430 18059
rect -1410 18038 -1406 18084
rect -1386 18038 -1382 18084
rect -1362 18038 -1358 18084
rect -1338 18038 -1334 18084
rect -1314 18038 -1310 18084
rect -1290 18038 -1286 18084
rect -1266 18038 -1262 18084
rect -1242 18038 -1238 18084
rect -1218 18038 -1214 18084
rect -1194 18038 -1190 18084
rect -1170 18038 -1166 18084
rect -1146 18038 -1142 18084
rect -1122 18038 -1118 18084
rect -1098 18038 -1094 18084
rect -1074 18038 -1070 18084
rect -1050 18038 -1046 18084
rect -1026 18038 -1022 18084
rect -1002 18038 -998 18084
rect -978 18038 -974 18084
rect -954 18038 -950 18084
rect -930 18038 -926 18084
rect -906 18038 -902 18084
rect -882 18038 -878 18084
rect -858 18038 -854 18084
rect -834 18038 -830 18084
rect -810 18038 -806 18084
rect -786 18038 -782 18084
rect -762 18038 -758 18084
rect -738 18038 -734 18084
rect -714 18038 -710 18084
rect -690 18059 -686 18084
rect -2393 18036 -693 18038
rect -2371 17990 -2366 18036
rect -2348 17990 -2343 18036
rect -2325 17990 -2320 18036
rect -2317 18032 -2309 18036
rect -2062 18032 -2054 18036
rect -2154 18028 -2138 18030
rect -2057 18028 -2054 18032
rect -2292 18022 -2054 18028
rect -2052 18022 -2044 18032
rect -2092 18006 -2062 18008
rect -2094 18002 -2062 18006
rect -2000 17990 -1992 18036
rect -1846 18029 -1806 18036
rect -1663 18032 -1655 18036
rect -1846 18022 -1680 18028
rect -1854 18006 -1806 18008
rect -1854 18002 -1680 18006
rect -1642 17990 -1637 18036
rect -1619 17990 -1614 18036
rect -1530 17990 -1526 18036
rect -1506 17990 -1502 18036
rect -1482 17990 -1478 18036
rect -1458 17990 -1454 18036
rect -1434 17990 -1430 18036
rect -1410 17990 -1406 18036
rect -1386 17990 -1382 18036
rect -1362 17990 -1358 18036
rect -1338 17990 -1334 18036
rect -1314 17990 -1310 18036
rect -1290 17990 -1286 18036
rect -1266 17990 -1262 18036
rect -1242 17990 -1238 18036
rect -1218 17990 -1214 18036
rect -1194 17990 -1190 18036
rect -1170 17990 -1166 18036
rect -1146 17990 -1142 18036
rect -1122 17990 -1118 18036
rect -1098 17990 -1094 18036
rect -1074 17990 -1070 18036
rect -1050 17990 -1046 18036
rect -1026 17990 -1022 18036
rect -1002 17990 -998 18036
rect -978 17990 -974 18036
rect -954 17990 -950 18036
rect -930 17990 -926 18036
rect -906 17990 -902 18036
rect -882 17990 -878 18036
rect -858 17990 -854 18036
rect -834 17990 -830 18036
rect -810 17990 -806 18036
rect -786 17990 -782 18036
rect -762 17990 -758 18036
rect -738 17990 -734 18036
rect -714 17990 -710 18036
rect -707 18035 -693 18036
rect -690 18035 -683 18059
rect -690 17990 -686 18035
rect -666 17990 -662 18084
rect -642 17990 -638 18084
rect -618 17990 -614 18084
rect -594 17990 -590 18084
rect -570 17990 -566 18084
rect -546 17990 -542 18084
rect -533 18053 -528 18063
rect -522 18053 -518 18084
rect -523 18039 -518 18053
rect -522 17990 -518 18039
rect -498 17990 -494 18084
rect -474 17990 -470 18084
rect -450 17990 -446 18084
rect -426 17990 -422 18084
rect -402 17990 -398 18084
rect -378 17990 -374 18084
rect -354 17990 -350 18084
rect -330 17990 -326 18084
rect -306 17990 -302 18084
rect -282 17990 -278 18084
rect -258 17990 -254 18084
rect -234 17990 -230 18084
rect -210 17990 -206 18084
rect -186 17990 -182 18084
rect -173 18029 -168 18039
rect -162 18029 -158 18084
rect -163 18015 -158 18029
rect -173 18005 -168 18015
rect -163 17991 -158 18005
rect -162 17990 -158 17991
rect -138 17990 -134 18084
rect -114 17990 -110 18084
rect -90 17990 -86 18084
rect -66 17990 -62 18084
rect -42 17990 -38 18084
rect -18 17990 -14 18084
rect 6 17990 10 18084
rect 30 17990 34 18084
rect 54 17990 58 18084
rect 78 17990 82 18084
rect 102 17990 106 18084
rect 126 17990 130 18084
rect 150 17990 154 18084
rect 174 17990 178 18084
rect 198 17990 202 18084
rect 222 17990 226 18084
rect 246 17990 250 18084
rect 270 17990 274 18084
rect 294 17990 298 18084
rect 318 17990 322 18084
rect 342 17990 346 18084
rect 366 17990 370 18084
rect 390 17990 394 18084
rect 414 17990 418 18084
rect 438 17990 442 18084
rect 462 17990 466 18084
rect 486 17990 490 18084
rect 510 17990 514 18084
rect 534 17990 538 18084
rect 558 17990 562 18084
rect 582 17990 586 18084
rect 606 17990 610 18084
rect 630 17990 634 18084
rect 654 17990 658 18084
rect 678 17990 682 18084
rect 702 17990 706 18084
rect 726 17990 730 18084
rect 750 17990 754 18084
rect 774 17990 778 18084
rect 798 17990 802 18084
rect 822 17990 826 18084
rect 846 17990 850 18084
rect 870 17990 874 18084
rect 894 17990 898 18084
rect 918 17990 922 18084
rect 942 17990 946 18084
rect 966 17990 970 18084
rect 990 17990 994 18084
rect 1014 17990 1018 18084
rect 1038 17990 1042 18084
rect 1062 17990 1066 18084
rect 1086 17990 1090 18084
rect 1110 17990 1114 18084
rect 1134 17990 1138 18084
rect 1158 17990 1162 18084
rect 1182 17990 1186 18084
rect 1206 17990 1210 18084
rect 1230 17990 1234 18084
rect 1254 17990 1258 18084
rect 1278 17990 1282 18084
rect 1302 17990 1306 18084
rect 1326 17990 1330 18084
rect 1350 17990 1354 18084
rect 1374 17990 1378 18084
rect 1398 17990 1402 18084
rect 1422 17990 1426 18084
rect 1446 17990 1450 18084
rect 1470 17990 1474 18084
rect 1494 17990 1498 18084
rect 1518 17990 1522 18084
rect 1542 17990 1546 18084
rect 1566 17990 1570 18084
rect 1590 17990 1594 18084
rect 1614 17990 1618 18084
rect 1638 17990 1642 18084
rect 1662 17990 1666 18084
rect 1686 17990 1690 18084
rect 1710 17990 1714 18084
rect 1734 17990 1738 18084
rect 1758 17990 1762 18084
rect 1782 17990 1786 18084
rect 1806 17990 1810 18084
rect 1830 17990 1834 18084
rect 1854 17990 1858 18084
rect 1878 17990 1882 18084
rect 1902 17990 1906 18084
rect 1926 17990 1930 18084
rect 1950 17990 1954 18084
rect 1974 17990 1978 18084
rect 1998 17990 2002 18084
rect 2022 17990 2026 18084
rect 2046 17990 2050 18084
rect 2070 17990 2074 18084
rect 2094 17990 2098 18084
rect 2118 17990 2122 18084
rect 2142 17990 2146 18084
rect 2166 17990 2170 18084
rect 2190 17990 2194 18084
rect 2214 17990 2218 18084
rect 2238 17990 2242 18084
rect 2262 17990 2266 18084
rect 2286 17990 2290 18084
rect 2310 17990 2314 18084
rect 2334 17990 2338 18084
rect 2358 17990 2362 18084
rect 2382 17990 2386 18084
rect 2406 17990 2410 18084
rect 2430 17990 2434 18084
rect 2454 17990 2458 18084
rect 2478 17990 2482 18084
rect 2502 17990 2506 18084
rect 2526 17990 2530 18084
rect 2550 17990 2554 18084
rect 2574 17990 2578 18084
rect 2598 17990 2602 18084
rect 2622 17990 2626 18084
rect 2646 17990 2650 18084
rect 2670 17990 2674 18084
rect 2694 17990 2698 18084
rect 2718 17990 2722 18084
rect 2742 17990 2746 18084
rect 2766 17990 2770 18084
rect 2790 17990 2794 18084
rect 2814 17990 2818 18084
rect 2838 17990 2842 18084
rect 2862 17990 2866 18084
rect 2886 17990 2890 18084
rect 2910 17990 2914 18084
rect 2934 17990 2938 18084
rect 2958 17990 2962 18084
rect 2982 17990 2986 18084
rect 3006 17990 3010 18084
rect 3030 17990 3034 18084
rect 3054 17990 3058 18084
rect 3078 17990 3082 18084
rect 3102 17990 3106 18084
rect 3126 17990 3130 18084
rect 3150 17990 3154 18084
rect 3174 17990 3178 18084
rect 3198 17990 3202 18084
rect 3222 17990 3226 18084
rect 3246 17990 3250 18084
rect 3270 17990 3274 18084
rect 3294 17990 3298 18084
rect 3318 17990 3322 18084
rect 3342 17990 3346 18084
rect 3366 17990 3370 18084
rect 3390 17990 3394 18084
rect 3414 17990 3418 18084
rect 3438 17990 3442 18084
rect 3462 17990 3466 18084
rect 3486 17990 3490 18084
rect 3510 17990 3514 18084
rect 3534 17990 3538 18084
rect 3558 17990 3562 18084
rect 3582 17990 3586 18084
rect 3606 17990 3610 18084
rect 3630 17990 3634 18084
rect 3654 17990 3658 18084
rect 3678 17990 3682 18084
rect 3702 17990 3706 18084
rect 3726 17990 3730 18084
rect 3733 18083 3747 18084
rect 3739 18077 3744 18083
rect 3749 18063 3754 18077
rect 3739 18005 3744 18015
rect 3750 18005 3754 18063
rect 3749 17991 3754 18005
rect 3763 18001 3771 18005
rect 3757 17991 3763 18001
rect 3739 17990 3771 17991
rect -2393 17988 3771 17990
rect -2371 17966 -2366 17988
rect -2348 17966 -2343 17988
rect -2325 17966 -2320 17988
rect -2072 17986 -2036 17987
rect -2072 17980 -2054 17986
rect -2309 17972 -2301 17980
rect -2317 17966 -2309 17972
rect -2092 17971 -2062 17976
rect -2000 17967 -1992 17988
rect -1938 17987 -1906 17988
rect -1920 17986 -1906 17987
rect -1806 17980 -1680 17986
rect -1854 17971 -1806 17976
rect -1655 17972 -1647 17980
rect -1982 17967 -1966 17968
rect -2000 17966 -1966 17967
rect -1846 17966 -1806 17969
rect -1663 17966 -1655 17972
rect -1642 17966 -1637 17988
rect -1619 17966 -1614 17988
rect -1530 17966 -1526 17988
rect -1506 17966 -1502 17988
rect -1482 17966 -1478 17988
rect -1458 17966 -1454 17988
rect -1434 17966 -1430 17988
rect -1410 17966 -1406 17988
rect -1386 17966 -1382 17988
rect -1362 17966 -1358 17988
rect -1338 17966 -1334 17988
rect -1314 17966 -1310 17988
rect -1290 17966 -1286 17988
rect -1266 17966 -1262 17988
rect -1242 17966 -1238 17988
rect -1218 17966 -1214 17988
rect -1194 17966 -1190 17988
rect -1170 17966 -1166 17988
rect -1146 17966 -1142 17988
rect -1122 17966 -1118 17988
rect -1098 17966 -1094 17988
rect -1074 17966 -1070 17988
rect -1050 17966 -1046 17988
rect -1026 17966 -1022 17988
rect -1002 17966 -998 17988
rect -978 17966 -974 17988
rect -954 17966 -950 17988
rect -930 17966 -926 17988
rect -906 17966 -902 17988
rect -882 17966 -878 17988
rect -858 17966 -854 17988
rect -834 17966 -830 17988
rect -810 17966 -806 17988
rect -786 17966 -782 17988
rect -762 17966 -758 17988
rect -738 17966 -734 17988
rect -714 17966 -710 17988
rect -690 17966 -686 17988
rect -666 17966 -662 17988
rect -642 17966 -638 17988
rect -618 17966 -614 17988
rect -594 17966 -590 17988
rect -570 17966 -566 17988
rect -546 17966 -542 17988
rect -522 17966 -518 17988
rect -498 17987 -494 17988
rect -2393 17964 -501 17966
rect -2371 17942 -2366 17964
rect -2348 17942 -2343 17964
rect -2325 17942 -2320 17964
rect -2000 17962 -1966 17964
rect -2309 17944 -2301 17952
rect -2062 17951 -2054 17958
rect -2092 17944 -2084 17951
rect -2062 17944 -2026 17946
rect -2317 17942 -2309 17944
rect -2062 17942 -2012 17944
rect -2000 17942 -1992 17962
rect -1982 17961 -1966 17962
rect -1846 17960 -1806 17964
rect -1846 17953 -1798 17958
rect -1806 17951 -1798 17953
rect -1854 17949 -1846 17951
rect -1854 17944 -1806 17949
rect -1655 17944 -1647 17952
rect -1864 17942 -1796 17943
rect -1663 17942 -1655 17944
rect -1642 17942 -1637 17964
rect -1619 17942 -1614 17964
rect -1530 17942 -1526 17964
rect -1506 17942 -1502 17964
rect -1482 17942 -1478 17964
rect -1458 17942 -1454 17964
rect -1434 17942 -1430 17964
rect -1410 17942 -1406 17964
rect -1386 17942 -1382 17964
rect -1362 17942 -1358 17964
rect -1338 17942 -1334 17964
rect -1314 17942 -1310 17964
rect -1290 17942 -1286 17964
rect -1266 17942 -1262 17964
rect -1242 17942 -1238 17964
rect -1218 17942 -1214 17964
rect -1194 17942 -1190 17964
rect -1170 17942 -1166 17964
rect -1146 17942 -1142 17964
rect -1122 17942 -1118 17964
rect -1098 17942 -1094 17964
rect -1074 17942 -1070 17964
rect -1050 17943 -1046 17964
rect -1061 17942 -1027 17943
rect -2393 17940 -1027 17942
rect -2371 17894 -2366 17940
rect -2348 17894 -2343 17940
rect -2325 17894 -2320 17940
rect -2317 17936 -2309 17940
rect -2062 17936 -2054 17940
rect -2154 17932 -2138 17934
rect -2057 17932 -2054 17936
rect -2292 17926 -2054 17932
rect -2052 17926 -2044 17936
rect -2092 17910 -2062 17912
rect -2094 17906 -2062 17910
rect -2000 17894 -1992 17940
rect -1846 17933 -1806 17940
rect -1663 17936 -1655 17940
rect -1846 17926 -1680 17932
rect -1854 17910 -1806 17912
rect -1854 17906 -1680 17910
rect -1642 17894 -1637 17940
rect -1619 17894 -1614 17940
rect -1530 17894 -1526 17940
rect -1506 17894 -1502 17940
rect -1482 17894 -1478 17940
rect -1458 17894 -1454 17940
rect -1434 17894 -1430 17940
rect -1410 17894 -1406 17940
rect -1386 17894 -1382 17940
rect -1362 17894 -1358 17940
rect -1338 17894 -1334 17940
rect -1314 17894 -1310 17940
rect -1290 17894 -1286 17940
rect -1266 17894 -1262 17940
rect -1242 17894 -1238 17940
rect -1218 17894 -1214 17940
rect -1194 17894 -1190 17940
rect -1170 17894 -1166 17940
rect -1146 17894 -1142 17940
rect -1122 17894 -1118 17940
rect -1098 17894 -1094 17940
rect -1074 17894 -1070 17940
rect -1061 17933 -1056 17940
rect -1050 17933 -1046 17940
rect -1051 17919 -1046 17933
rect -1050 17894 -1046 17919
rect -1026 17894 -1022 17964
rect -1002 17894 -998 17964
rect -978 17894 -974 17964
rect -954 17894 -950 17964
rect -930 17894 -926 17964
rect -906 17894 -902 17964
rect -882 17894 -878 17964
rect -858 17894 -854 17964
rect -834 17894 -830 17964
rect -810 17894 -806 17964
rect -786 17894 -782 17964
rect -762 17894 -758 17964
rect -738 17894 -734 17964
rect -714 17894 -710 17964
rect -690 17894 -686 17964
rect -666 17894 -662 17964
rect -642 17894 -638 17964
rect -618 17894 -614 17964
rect -594 17894 -590 17964
rect -570 17894 -566 17964
rect -546 17894 -542 17964
rect -522 17894 -518 17964
rect -515 17963 -501 17964
rect -498 17963 -491 17987
rect -498 17894 -494 17963
rect -474 17894 -470 17988
rect -450 17894 -446 17988
rect -426 17894 -422 17988
rect -402 17894 -398 17988
rect -378 17894 -374 17988
rect -354 17894 -350 17988
rect -330 17894 -326 17988
rect -306 17894 -302 17988
rect -282 17894 -278 17988
rect -258 17894 -254 17988
rect -234 17894 -230 17988
rect -210 17894 -206 17988
rect -186 17894 -182 17988
rect -162 17894 -158 17988
rect -138 17963 -134 17988
rect -138 17915 -131 17963
rect -138 17894 -134 17915
rect -114 17894 -110 17988
rect -90 17894 -86 17988
rect -66 17894 -62 17988
rect -42 17894 -38 17988
rect -18 17894 -14 17988
rect 6 17894 10 17988
rect 30 17894 34 17988
rect 54 17894 58 17988
rect 78 17894 82 17988
rect 102 17894 106 17988
rect 126 17894 130 17988
rect 150 17894 154 17988
rect 174 17894 178 17988
rect 198 17894 202 17988
rect 222 17894 226 17988
rect 246 17894 250 17988
rect 270 17894 274 17988
rect 294 17894 298 17988
rect 318 17894 322 17988
rect 342 17894 346 17988
rect 366 17894 370 17988
rect 390 17894 394 17988
rect 414 17894 418 17988
rect 438 17894 442 17988
rect 462 17894 466 17988
rect 486 17894 490 17988
rect 510 17894 514 17988
rect 534 17894 538 17988
rect 558 17894 562 17988
rect 582 17894 586 17988
rect 606 17894 610 17988
rect 630 17894 634 17988
rect 654 17894 658 17988
rect 678 17894 682 17988
rect 702 17894 706 17988
rect 726 17894 730 17988
rect 750 17894 754 17988
rect 774 17894 778 17988
rect 798 17894 802 17988
rect 822 17894 826 17988
rect 846 17894 850 17988
rect 870 17894 874 17988
rect 894 17894 898 17988
rect 918 17894 922 17988
rect 942 17894 946 17988
rect 966 17894 970 17988
rect 990 17894 994 17988
rect 1014 17894 1018 17988
rect 1038 17894 1042 17988
rect 1062 17894 1066 17988
rect 1086 17894 1090 17988
rect 1110 17894 1114 17988
rect 1134 17894 1138 17988
rect 1158 17894 1162 17988
rect 1182 17894 1186 17988
rect 1206 17894 1210 17988
rect 1230 17894 1234 17988
rect 1254 17894 1258 17988
rect 1278 17894 1282 17988
rect 1302 17894 1306 17988
rect 1326 17894 1330 17988
rect 1350 17894 1354 17988
rect 1374 17894 1378 17988
rect 1398 17894 1402 17988
rect 1422 17894 1426 17988
rect 1446 17894 1450 17988
rect 1470 17894 1474 17988
rect 1494 17894 1498 17988
rect 1518 17894 1522 17988
rect 1542 17894 1546 17988
rect 1566 17894 1570 17988
rect 1590 17894 1594 17988
rect 1614 17894 1618 17988
rect 1638 17894 1642 17988
rect 1662 17894 1666 17988
rect 1686 17894 1690 17988
rect 1710 17894 1714 17988
rect 1734 17894 1738 17988
rect 1758 17894 1762 17988
rect 1782 17894 1786 17988
rect 1806 17894 1810 17988
rect 1830 17894 1834 17988
rect 1854 17894 1858 17988
rect 1878 17894 1882 17988
rect 1902 17894 1906 17988
rect 1926 17894 1930 17988
rect 1950 17894 1954 17988
rect 1974 17894 1978 17988
rect 1998 17894 2002 17988
rect 2022 17894 2026 17988
rect 2046 17894 2050 17988
rect 2070 17894 2074 17988
rect 2094 17894 2098 17988
rect 2118 17894 2122 17988
rect 2142 17894 2146 17988
rect 2155 17957 2160 17967
rect 2166 17957 2170 17988
rect 2165 17943 2170 17957
rect 2155 17933 2160 17943
rect 2165 17919 2170 17933
rect 2166 17894 2170 17919
rect 2190 17894 2194 17988
rect 2214 17894 2218 17988
rect 2238 17894 2242 17988
rect 2262 17894 2266 17988
rect 2286 17894 2290 17988
rect 2310 17894 2314 17988
rect 2334 17894 2338 17988
rect 2358 17894 2362 17988
rect 2382 17894 2386 17988
rect 2406 17894 2410 17988
rect 2430 17894 2434 17988
rect 2454 17894 2458 17988
rect 2478 17894 2482 17988
rect 2502 17894 2506 17988
rect 2526 17894 2530 17988
rect 2550 17894 2554 17988
rect 2574 17894 2578 17988
rect 2598 17894 2602 17988
rect 2622 17894 2626 17988
rect 2646 17894 2650 17988
rect 2670 17894 2674 17988
rect 2694 17894 2698 17988
rect 2718 17894 2722 17988
rect 2742 17894 2746 17988
rect 2766 17894 2770 17988
rect 2790 17894 2794 17988
rect 2814 17894 2818 17988
rect 2838 17894 2842 17988
rect 2862 17894 2866 17988
rect 2886 17894 2890 17988
rect 2910 17894 2914 17988
rect 2934 17894 2938 17988
rect 2958 17894 2962 17988
rect 2982 17894 2986 17988
rect 3006 17894 3010 17988
rect 3030 17894 3034 17988
rect 3054 17894 3058 17988
rect 3078 17894 3082 17988
rect 3102 17894 3106 17988
rect 3126 17894 3130 17988
rect 3150 17894 3154 17988
rect 3174 17894 3178 17988
rect 3198 17894 3202 17988
rect 3222 17894 3226 17988
rect 3246 17894 3250 17988
rect 3270 17894 3274 17988
rect 3294 17894 3298 17988
rect 3318 17894 3322 17988
rect 3342 17894 3346 17988
rect 3366 17894 3370 17988
rect 3390 17894 3394 17988
rect 3414 17894 3418 17988
rect 3438 17894 3442 17988
rect 3462 17894 3466 17988
rect 3486 17894 3490 17988
rect 3510 17894 3514 17988
rect 3534 17894 3538 17988
rect 3558 17894 3562 17988
rect 3582 17894 3586 17988
rect 3606 17894 3610 17988
rect 3630 17894 3634 17988
rect 3654 17894 3658 17988
rect 3678 17894 3682 17988
rect 3702 17894 3706 17988
rect 3726 17894 3730 17988
rect 3739 17981 3744 17988
rect 3757 17987 3771 17988
rect 3749 17967 3754 17981
rect 3739 17933 3744 17943
rect 3750 17933 3754 17967
rect 3749 17919 3754 17933
rect 3763 17929 3771 17933
rect 3757 17919 3763 17929
rect 3739 17894 3771 17895
rect -2393 17892 3771 17894
rect -2371 17870 -2366 17892
rect -2348 17870 -2343 17892
rect -2325 17870 -2320 17892
rect -2072 17890 -2036 17891
rect -2072 17884 -2054 17890
rect -2309 17876 -2301 17884
rect -2317 17870 -2309 17876
rect -2092 17875 -2062 17880
rect -2000 17871 -1992 17892
rect -1938 17891 -1906 17892
rect -1920 17890 -1906 17891
rect -1806 17884 -1680 17890
rect -1854 17875 -1806 17880
rect -1655 17876 -1647 17884
rect -1982 17871 -1966 17872
rect -2000 17870 -1966 17871
rect -1846 17870 -1806 17873
rect -1663 17870 -1655 17876
rect -1642 17870 -1637 17892
rect -1619 17870 -1614 17892
rect -1530 17870 -1526 17892
rect -1506 17870 -1502 17892
rect -1482 17870 -1478 17892
rect -1458 17870 -1454 17892
rect -1434 17870 -1430 17892
rect -1410 17870 -1406 17892
rect -1386 17870 -1382 17892
rect -1362 17870 -1358 17892
rect -1338 17870 -1334 17892
rect -1314 17870 -1310 17892
rect -1290 17870 -1286 17892
rect -1266 17870 -1262 17892
rect -1242 17870 -1238 17892
rect -1218 17870 -1214 17892
rect -1194 17870 -1190 17892
rect -1170 17870 -1166 17892
rect -1146 17870 -1142 17892
rect -1122 17870 -1118 17892
rect -1098 17870 -1094 17892
rect -1074 17870 -1070 17892
rect -1050 17870 -1046 17892
rect -1026 17870 -1022 17892
rect -1002 17870 -998 17892
rect -978 17870 -974 17892
rect -954 17870 -950 17892
rect -930 17870 -926 17892
rect -906 17870 -902 17892
rect -882 17870 -878 17892
rect -858 17870 -854 17892
rect -834 17870 -830 17892
rect -810 17870 -806 17892
rect -786 17870 -782 17892
rect -762 17870 -758 17892
rect -738 17870 -734 17892
rect -714 17870 -710 17892
rect -690 17870 -686 17892
rect -666 17870 -662 17892
rect -642 17870 -638 17892
rect -618 17870 -614 17892
rect -594 17870 -590 17892
rect -570 17870 -566 17892
rect -546 17870 -542 17892
rect -522 17870 -518 17892
rect -498 17870 -494 17892
rect -474 17870 -470 17892
rect -450 17870 -446 17892
rect -426 17870 -422 17892
rect -402 17870 -398 17892
rect -378 17870 -374 17892
rect -354 17870 -350 17892
rect -330 17870 -326 17892
rect -306 17870 -302 17892
rect -282 17870 -278 17892
rect -258 17870 -254 17892
rect -234 17870 -230 17892
rect -210 17870 -206 17892
rect -186 17870 -182 17892
rect -162 17870 -158 17892
rect -138 17870 -134 17892
rect -114 17870 -110 17892
rect -90 17870 -86 17892
rect -66 17870 -62 17892
rect -42 17870 -38 17892
rect -18 17870 -14 17892
rect 6 17870 10 17892
rect 30 17870 34 17892
rect 54 17870 58 17892
rect 78 17870 82 17892
rect 102 17870 106 17892
rect 126 17870 130 17892
rect 150 17870 154 17892
rect 174 17870 178 17892
rect 198 17870 202 17892
rect 222 17870 226 17892
rect 246 17870 250 17892
rect 270 17871 274 17892
rect 259 17870 293 17871
rect -2393 17868 293 17870
rect -2371 17846 -2366 17868
rect -2348 17846 -2343 17868
rect -2325 17846 -2320 17868
rect -2000 17866 -1966 17868
rect -2309 17848 -2301 17856
rect -2062 17855 -2054 17862
rect -2092 17848 -2084 17855
rect -2062 17848 -2026 17850
rect -2317 17846 -2309 17848
rect -2062 17846 -2012 17848
rect -2000 17846 -1992 17866
rect -1982 17865 -1966 17866
rect -1846 17864 -1806 17868
rect -1846 17857 -1798 17862
rect -1806 17855 -1798 17857
rect -1854 17853 -1846 17855
rect -1854 17848 -1806 17853
rect -1655 17848 -1647 17856
rect -1864 17846 -1796 17847
rect -1663 17846 -1655 17848
rect -1642 17846 -1637 17868
rect -1619 17846 -1614 17868
rect -1530 17846 -1526 17868
rect -1506 17846 -1502 17868
rect -1482 17846 -1478 17868
rect -1458 17846 -1454 17868
rect -1434 17846 -1430 17868
rect -1410 17846 -1406 17868
rect -1386 17846 -1382 17868
rect -1362 17846 -1358 17868
rect -1338 17846 -1334 17868
rect -1314 17846 -1310 17868
rect -1290 17846 -1286 17868
rect -1266 17846 -1262 17868
rect -1242 17846 -1238 17868
rect -1218 17846 -1214 17868
rect -1194 17846 -1190 17868
rect -1170 17846 -1166 17868
rect -1146 17846 -1142 17868
rect -1122 17846 -1118 17868
rect -1098 17846 -1094 17868
rect -1074 17846 -1070 17868
rect -1050 17847 -1046 17868
rect -1026 17867 -1022 17868
rect -1061 17846 -1029 17847
rect -2393 17844 -1029 17846
rect -2371 17798 -2366 17844
rect -2348 17798 -2343 17844
rect -2325 17798 -2320 17844
rect -2317 17840 -2309 17844
rect -2062 17840 -2054 17844
rect -2154 17836 -2138 17838
rect -2057 17836 -2054 17840
rect -2292 17830 -2054 17836
rect -2052 17830 -2044 17840
rect -2092 17814 -2062 17816
rect -2094 17810 -2062 17814
rect -2000 17798 -1992 17844
rect -1846 17837 -1806 17844
rect -1663 17840 -1655 17844
rect -1846 17830 -1680 17836
rect -1854 17814 -1806 17816
rect -1854 17810 -1680 17814
rect -1642 17798 -1637 17844
rect -1619 17798 -1614 17844
rect -1530 17798 -1526 17844
rect -1506 17798 -1502 17844
rect -1482 17798 -1478 17844
rect -1458 17798 -1454 17844
rect -1434 17798 -1430 17844
rect -1410 17798 -1406 17844
rect -1386 17798 -1382 17844
rect -1362 17798 -1358 17844
rect -1338 17798 -1334 17844
rect -1314 17798 -1310 17844
rect -1290 17798 -1286 17844
rect -1266 17798 -1262 17844
rect -1242 17798 -1238 17844
rect -1218 17798 -1214 17844
rect -1194 17798 -1190 17844
rect -1170 17798 -1166 17844
rect -1146 17798 -1142 17844
rect -1122 17798 -1118 17844
rect -1098 17798 -1094 17844
rect -1074 17798 -1070 17844
rect -1061 17837 -1056 17844
rect -1050 17837 -1046 17844
rect -1043 17843 -1029 17844
rect -1026 17843 -1019 17867
rect -1051 17823 -1046 17837
rect -1050 17798 -1046 17823
rect -1026 17798 -1022 17843
rect -1002 17798 -998 17868
rect -978 17798 -974 17868
rect -954 17798 -950 17868
rect -930 17798 -926 17868
rect -906 17798 -902 17868
rect -882 17798 -878 17868
rect -858 17798 -854 17868
rect -834 17798 -830 17868
rect -810 17798 -806 17868
rect -786 17798 -782 17868
rect -762 17798 -758 17868
rect -738 17798 -734 17868
rect -714 17798 -710 17868
rect -690 17798 -686 17868
rect -666 17798 -662 17868
rect -642 17798 -638 17868
rect -618 17798 -614 17868
rect -594 17798 -590 17868
rect -570 17798 -566 17868
rect -546 17798 -542 17868
rect -522 17798 -518 17868
rect -498 17798 -494 17868
rect -474 17798 -470 17868
rect -450 17798 -446 17868
rect -426 17798 -422 17868
rect -402 17798 -398 17868
rect -378 17798 -374 17868
rect -354 17798 -350 17868
rect -330 17798 -326 17868
rect -306 17798 -302 17868
rect -282 17798 -278 17868
rect -258 17798 -254 17868
rect -234 17798 -230 17868
rect -210 17798 -206 17868
rect -186 17798 -182 17868
rect -162 17798 -158 17868
rect -138 17798 -134 17868
rect -114 17798 -110 17868
rect -90 17798 -86 17868
rect -66 17798 -62 17868
rect -42 17798 -38 17868
rect -18 17798 -14 17868
rect 6 17798 10 17868
rect 30 17798 34 17868
rect 54 17798 58 17868
rect 78 17798 82 17868
rect 102 17798 106 17868
rect 126 17798 130 17868
rect 150 17798 154 17868
rect 174 17798 178 17868
rect 198 17798 202 17868
rect 222 17798 226 17868
rect 246 17798 250 17868
rect 259 17861 264 17868
rect 270 17861 274 17868
rect 269 17847 274 17861
rect 259 17837 264 17847
rect 269 17823 274 17837
rect 270 17798 274 17823
rect 294 17798 298 17892
rect 318 17798 322 17892
rect 342 17798 346 17892
rect 366 17798 370 17892
rect 390 17798 394 17892
rect 414 17798 418 17892
rect 438 17798 442 17892
rect 462 17798 466 17892
rect 486 17798 490 17892
rect 510 17798 514 17892
rect 534 17798 538 17892
rect 558 17798 562 17892
rect 582 17798 586 17892
rect 606 17798 610 17892
rect 630 17798 634 17892
rect 654 17798 658 17892
rect 678 17798 682 17892
rect 702 17798 706 17892
rect 726 17798 730 17892
rect 750 17798 754 17892
rect 774 17798 778 17892
rect 798 17798 802 17892
rect 822 17798 826 17892
rect 846 17798 850 17892
rect 870 17798 874 17892
rect 894 17798 898 17892
rect 918 17798 922 17892
rect 942 17798 946 17892
rect 966 17798 970 17892
rect 990 17798 994 17892
rect 1014 17798 1018 17892
rect 1038 17798 1042 17892
rect 1062 17798 1066 17892
rect 1086 17798 1090 17892
rect 1110 17798 1114 17892
rect 1134 17798 1138 17892
rect 1158 17798 1162 17892
rect 1182 17798 1186 17892
rect 1206 17798 1210 17892
rect 1230 17798 1234 17892
rect 1254 17798 1258 17892
rect 1278 17798 1282 17892
rect 1302 17798 1306 17892
rect 1326 17798 1330 17892
rect 1350 17798 1354 17892
rect 1374 17798 1378 17892
rect 1398 17798 1402 17892
rect 1422 17798 1426 17892
rect 1446 17798 1450 17892
rect 1470 17798 1474 17892
rect 1494 17798 1498 17892
rect 1518 17798 1522 17892
rect 1542 17798 1546 17892
rect 1566 17798 1570 17892
rect 1590 17798 1594 17892
rect 1614 17798 1618 17892
rect 1638 17798 1642 17892
rect 1662 17798 1666 17892
rect 1686 17798 1690 17892
rect 1710 17798 1714 17892
rect 1734 17798 1738 17892
rect 1758 17798 1762 17892
rect 1782 17798 1786 17892
rect 1806 17798 1810 17892
rect 1830 17798 1834 17892
rect 1854 17798 1858 17892
rect 1878 17798 1882 17892
rect 1902 17798 1906 17892
rect 1926 17798 1930 17892
rect 1950 17798 1954 17892
rect 1974 17798 1978 17892
rect 1998 17798 2002 17892
rect 2022 17798 2026 17892
rect 2046 17798 2050 17892
rect 2070 17798 2074 17892
rect 2094 17798 2098 17892
rect 2118 17798 2122 17892
rect 2142 17798 2146 17892
rect 2166 17798 2170 17892
rect 2190 17891 2194 17892
rect 2190 17846 2197 17891
rect 2214 17846 2218 17892
rect 2238 17846 2242 17892
rect 2262 17846 2266 17892
rect 2286 17846 2290 17892
rect 2310 17846 2314 17892
rect 2334 17846 2338 17892
rect 2358 17846 2362 17892
rect 2382 17846 2386 17892
rect 2406 17846 2410 17892
rect 2430 17846 2434 17892
rect 2454 17846 2458 17892
rect 2478 17846 2482 17892
rect 2502 17846 2506 17892
rect 2526 17846 2530 17892
rect 2550 17846 2554 17892
rect 2574 17846 2578 17892
rect 2598 17846 2602 17892
rect 2622 17846 2626 17892
rect 2646 17846 2650 17892
rect 2670 17846 2674 17892
rect 2694 17846 2698 17892
rect 2718 17846 2722 17892
rect 2742 17846 2746 17892
rect 2766 17846 2770 17892
rect 2790 17846 2794 17892
rect 2814 17846 2818 17892
rect 2838 17846 2842 17892
rect 2862 17846 2866 17892
rect 2886 17846 2890 17892
rect 2910 17846 2914 17892
rect 2934 17846 2938 17892
rect 2958 17846 2962 17892
rect 2982 17846 2986 17892
rect 3006 17846 3010 17892
rect 3030 17846 3034 17892
rect 3054 17846 3058 17892
rect 3078 17846 3082 17892
rect 3102 17846 3106 17892
rect 3126 17846 3130 17892
rect 3150 17846 3154 17892
rect 3174 17846 3178 17892
rect 3198 17846 3202 17892
rect 3222 17846 3226 17892
rect 3246 17846 3250 17892
rect 3270 17846 3274 17892
rect 3294 17846 3298 17892
rect 3318 17846 3322 17892
rect 3342 17846 3346 17892
rect 3366 17846 3370 17892
rect 3390 17846 3394 17892
rect 3414 17846 3418 17892
rect 3438 17846 3442 17892
rect 3462 17846 3466 17892
rect 3486 17846 3490 17892
rect 3510 17846 3514 17892
rect 3534 17846 3538 17892
rect 3558 17846 3562 17892
rect 3582 17846 3586 17892
rect 3606 17846 3610 17892
rect 3630 17846 3634 17892
rect 3654 17846 3658 17892
rect 3678 17846 3682 17892
rect 3702 17846 3706 17892
rect 3726 17846 3730 17892
rect 3739 17885 3744 17892
rect 3757 17891 3771 17892
rect 3749 17871 3754 17885
rect 3750 17847 3754 17871
rect 3739 17846 3771 17847
rect 2173 17844 3771 17846
rect 2173 17843 2187 17844
rect 2190 17843 2197 17844
rect 2190 17798 2194 17843
rect 2214 17798 2218 17844
rect 2238 17798 2242 17844
rect 2262 17798 2266 17844
rect 2286 17798 2290 17844
rect 2310 17798 2314 17844
rect 2334 17798 2338 17844
rect 2358 17798 2362 17844
rect 2382 17798 2386 17844
rect 2406 17798 2410 17844
rect 2430 17798 2434 17844
rect 2454 17798 2458 17844
rect 2478 17798 2482 17844
rect 2502 17798 2506 17844
rect 2526 17798 2530 17844
rect 2550 17798 2554 17844
rect 2574 17798 2578 17844
rect 2598 17798 2602 17844
rect 2622 17798 2626 17844
rect 2646 17798 2650 17844
rect 2670 17798 2674 17844
rect 2694 17798 2698 17844
rect 2718 17798 2722 17844
rect 2742 17798 2746 17844
rect 2766 17798 2770 17844
rect 2790 17798 2794 17844
rect 2814 17798 2818 17844
rect 2838 17798 2842 17844
rect 2862 17798 2866 17844
rect 2886 17798 2890 17844
rect 2910 17798 2914 17844
rect 2934 17798 2938 17844
rect 2958 17798 2962 17844
rect 2982 17798 2986 17844
rect 3006 17798 3010 17844
rect 3030 17798 3034 17844
rect 3054 17798 3058 17844
rect 3078 17798 3082 17844
rect 3102 17798 3106 17844
rect 3126 17798 3130 17844
rect 3150 17798 3154 17844
rect 3174 17798 3178 17844
rect 3198 17798 3202 17844
rect 3222 17798 3226 17844
rect 3246 17798 3250 17844
rect 3270 17798 3274 17844
rect 3294 17798 3298 17844
rect 3318 17798 3322 17844
rect 3342 17798 3346 17844
rect 3366 17798 3370 17844
rect 3390 17798 3394 17844
rect 3414 17798 3418 17844
rect 3438 17798 3442 17844
rect 3462 17798 3466 17844
rect 3486 17798 3490 17844
rect 3510 17798 3514 17844
rect 3534 17798 3538 17844
rect 3558 17798 3562 17844
rect 3582 17798 3586 17844
rect 3606 17798 3610 17844
rect 3630 17798 3634 17844
rect 3654 17798 3658 17844
rect 3678 17798 3682 17844
rect 3702 17798 3706 17844
rect 3726 17798 3730 17844
rect 3739 17837 3744 17844
rect 3750 17837 3754 17844
rect 3757 17843 3771 17844
rect 3749 17823 3754 17837
rect 3739 17798 3771 17799
rect -2393 17796 3771 17798
rect -2371 17774 -2366 17796
rect -2348 17774 -2343 17796
rect -2325 17774 -2320 17796
rect -2072 17794 -2036 17795
rect -2072 17788 -2054 17794
rect -2309 17780 -2301 17788
rect -2317 17774 -2309 17780
rect -2092 17779 -2062 17784
rect -2000 17775 -1992 17796
rect -1938 17795 -1906 17796
rect -1920 17794 -1906 17795
rect -1806 17788 -1680 17794
rect -1854 17779 -1806 17784
rect -1655 17780 -1647 17788
rect -1982 17775 -1966 17776
rect -2000 17774 -1966 17775
rect -1846 17774 -1806 17777
rect -1663 17774 -1655 17780
rect -1642 17774 -1637 17796
rect -1619 17774 -1614 17796
rect -1530 17774 -1526 17796
rect -1506 17774 -1502 17796
rect -1482 17774 -1478 17796
rect -1458 17774 -1454 17796
rect -1434 17774 -1430 17796
rect -1410 17775 -1406 17796
rect -1421 17774 -1387 17775
rect -2393 17772 -1387 17774
rect -2371 17750 -2366 17772
rect -2348 17750 -2343 17772
rect -2325 17750 -2320 17772
rect -2000 17770 -1966 17772
rect -2309 17752 -2301 17760
rect -2062 17759 -2054 17766
rect -2092 17752 -2084 17759
rect -2062 17752 -2026 17754
rect -2317 17750 -2309 17752
rect -2062 17750 -2012 17752
rect -2000 17750 -1992 17770
rect -1982 17769 -1966 17770
rect -1846 17768 -1806 17772
rect -1846 17761 -1798 17766
rect -1806 17759 -1798 17761
rect -1854 17757 -1846 17759
rect -1854 17752 -1806 17757
rect -1655 17752 -1647 17760
rect -1864 17750 -1796 17751
rect -1663 17750 -1655 17752
rect -1642 17750 -1637 17772
rect -1619 17750 -1614 17772
rect -1530 17750 -1526 17772
rect -1506 17750 -1502 17772
rect -1482 17750 -1478 17772
rect -1458 17750 -1454 17772
rect -1434 17750 -1430 17772
rect -1421 17765 -1416 17772
rect -1410 17765 -1406 17772
rect -1411 17751 -1406 17765
rect -1410 17750 -1406 17751
rect -1386 17750 -1382 17796
rect -1362 17750 -1358 17796
rect -1338 17750 -1334 17796
rect -1314 17750 -1310 17796
rect -1290 17750 -1286 17796
rect -1266 17750 -1262 17796
rect -1242 17750 -1238 17796
rect -1218 17750 -1214 17796
rect -1194 17750 -1190 17796
rect -1170 17750 -1166 17796
rect -1146 17750 -1142 17796
rect -1122 17750 -1118 17796
rect -1098 17750 -1094 17796
rect -1074 17750 -1070 17796
rect -1050 17751 -1046 17796
rect -1026 17771 -1022 17796
rect -1061 17750 -1029 17751
rect -2393 17748 -1029 17750
rect -2371 17702 -2366 17748
rect -2348 17702 -2343 17748
rect -2325 17702 -2320 17748
rect -2317 17744 -2309 17748
rect -2062 17744 -2054 17748
rect -2154 17740 -2138 17742
rect -2057 17740 -2054 17744
rect -2292 17734 -2054 17740
rect -2052 17734 -2044 17744
rect -2092 17718 -2062 17720
rect -2094 17714 -2062 17718
rect -2000 17702 -1992 17748
rect -1846 17741 -1806 17748
rect -1663 17744 -1655 17748
rect -1846 17734 -1680 17740
rect -1854 17718 -1806 17720
rect -1854 17714 -1680 17718
rect -1642 17702 -1637 17748
rect -1619 17702 -1614 17748
rect -1530 17702 -1526 17748
rect -1506 17702 -1502 17748
rect -1482 17702 -1478 17748
rect -1458 17702 -1454 17748
rect -1434 17702 -1430 17748
rect -1410 17702 -1406 17748
rect -1386 17702 -1382 17748
rect -1362 17702 -1358 17748
rect -1338 17702 -1334 17748
rect -1314 17702 -1310 17748
rect -1290 17702 -1286 17748
rect -1266 17702 -1262 17748
rect -1242 17702 -1238 17748
rect -1218 17702 -1214 17748
rect -1194 17702 -1190 17748
rect -1170 17702 -1166 17748
rect -1146 17702 -1142 17748
rect -1122 17702 -1118 17748
rect -1098 17702 -1094 17748
rect -1074 17702 -1070 17748
rect -1061 17741 -1056 17748
rect -1050 17741 -1046 17748
rect -1043 17747 -1029 17748
rect -1026 17747 -1019 17771
rect -1051 17727 -1046 17741
rect -1050 17702 -1046 17727
rect -1026 17702 -1022 17747
rect -1002 17702 -998 17796
rect -978 17702 -974 17796
rect -954 17702 -950 17796
rect -930 17702 -926 17796
rect -906 17702 -902 17796
rect -882 17702 -878 17796
rect -858 17702 -854 17796
rect -834 17702 -830 17796
rect -810 17702 -806 17796
rect -786 17702 -782 17796
rect -762 17702 -758 17796
rect -738 17702 -734 17796
rect -714 17702 -710 17796
rect -690 17702 -686 17796
rect -666 17702 -662 17796
rect -642 17702 -638 17796
rect -618 17702 -614 17796
rect -594 17702 -590 17796
rect -570 17702 -566 17796
rect -546 17702 -542 17796
rect -522 17702 -518 17796
rect -498 17702 -494 17796
rect -474 17702 -470 17796
rect -450 17702 -446 17796
rect -426 17702 -422 17796
rect -402 17702 -398 17796
rect -378 17702 -374 17796
rect -354 17702 -350 17796
rect -330 17702 -326 17796
rect -306 17702 -302 17796
rect -282 17702 -278 17796
rect -258 17702 -254 17796
rect -234 17702 -230 17796
rect -210 17702 -206 17796
rect -186 17702 -182 17796
rect -162 17702 -158 17796
rect -138 17702 -134 17796
rect -114 17702 -110 17796
rect -90 17702 -86 17796
rect -66 17702 -62 17796
rect -42 17702 -38 17796
rect -18 17702 -14 17796
rect 6 17702 10 17796
rect 30 17702 34 17796
rect 54 17702 58 17796
rect 78 17702 82 17796
rect 102 17702 106 17796
rect 126 17702 130 17796
rect 150 17702 154 17796
rect 174 17702 178 17796
rect 198 17702 202 17796
rect 222 17702 226 17796
rect 246 17702 250 17796
rect 270 17702 274 17796
rect 294 17795 298 17796
rect 294 17747 301 17795
rect 294 17702 298 17747
rect 318 17702 322 17796
rect 342 17702 346 17796
rect 366 17702 370 17796
rect 390 17702 394 17796
rect 414 17702 418 17796
rect 438 17702 442 17796
rect 462 17702 466 17796
rect 486 17702 490 17796
rect 510 17702 514 17796
rect 534 17702 538 17796
rect 558 17702 562 17796
rect 582 17702 586 17796
rect 606 17702 610 17796
rect 630 17702 634 17796
rect 654 17702 658 17796
rect 678 17702 682 17796
rect 702 17702 706 17796
rect 726 17702 730 17796
rect 750 17702 754 17796
rect 774 17702 778 17796
rect 798 17702 802 17796
rect 822 17702 826 17796
rect 846 17702 850 17796
rect 870 17702 874 17796
rect 894 17702 898 17796
rect 918 17702 922 17796
rect 942 17702 946 17796
rect 966 17702 970 17796
rect 990 17702 994 17796
rect 1014 17702 1018 17796
rect 1038 17702 1042 17796
rect 1062 17702 1066 17796
rect 1086 17702 1090 17796
rect 1110 17702 1114 17796
rect 1134 17702 1138 17796
rect 1158 17702 1162 17796
rect 1182 17702 1186 17796
rect 1206 17702 1210 17796
rect 1230 17702 1234 17796
rect 1254 17702 1258 17796
rect 1278 17702 1282 17796
rect 1302 17702 1306 17796
rect 1326 17702 1330 17796
rect 1350 17702 1354 17796
rect 1374 17702 1378 17796
rect 1398 17702 1402 17796
rect 1422 17702 1426 17796
rect 1446 17702 1450 17796
rect 1470 17702 1474 17796
rect 1494 17702 1498 17796
rect 1518 17702 1522 17796
rect 1542 17702 1546 17796
rect 1566 17702 1570 17796
rect 1590 17702 1594 17796
rect 1614 17702 1618 17796
rect 1638 17702 1642 17796
rect 1662 17702 1666 17796
rect 1686 17702 1690 17796
rect 1710 17702 1714 17796
rect 1734 17702 1738 17796
rect 1758 17702 1762 17796
rect 1782 17702 1786 17796
rect 1806 17702 1810 17796
rect 1830 17702 1834 17796
rect 1854 17702 1858 17796
rect 1878 17702 1882 17796
rect 1902 17702 1906 17796
rect 1926 17702 1930 17796
rect 1950 17702 1954 17796
rect 1974 17702 1978 17796
rect 1998 17702 2002 17796
rect 2022 17702 2026 17796
rect 2046 17702 2050 17796
rect 2070 17702 2074 17796
rect 2094 17702 2098 17796
rect 2118 17702 2122 17796
rect 2142 17702 2146 17796
rect 2166 17702 2170 17796
rect 2190 17702 2194 17796
rect 2214 17702 2218 17796
rect 2238 17702 2242 17796
rect 2262 17702 2266 17796
rect 2286 17702 2290 17796
rect 2310 17702 2314 17796
rect 2334 17702 2338 17796
rect 2358 17702 2362 17796
rect 2382 17702 2386 17796
rect 2406 17702 2410 17796
rect 2430 17702 2434 17796
rect 2454 17702 2458 17796
rect 2478 17702 2482 17796
rect 2502 17702 2506 17796
rect 2526 17702 2530 17796
rect 2550 17702 2554 17796
rect 2574 17702 2578 17796
rect 2598 17702 2602 17796
rect 2622 17702 2626 17796
rect 2646 17702 2650 17796
rect 2670 17702 2674 17796
rect 2694 17702 2698 17796
rect 2718 17702 2722 17796
rect 2742 17702 2746 17796
rect 2766 17702 2770 17796
rect 2790 17702 2794 17796
rect 2814 17702 2818 17796
rect 2838 17702 2842 17796
rect 2862 17702 2866 17796
rect 2886 17702 2890 17796
rect 2910 17702 2914 17796
rect 2934 17702 2938 17796
rect 2958 17702 2962 17796
rect 2982 17702 2986 17796
rect 3006 17702 3010 17796
rect 3030 17702 3034 17796
rect 3054 17702 3058 17796
rect 3078 17702 3082 17796
rect 3102 17702 3106 17796
rect 3126 17702 3130 17796
rect 3150 17702 3154 17796
rect 3174 17702 3178 17796
rect 3198 17702 3202 17796
rect 3222 17702 3226 17796
rect 3246 17702 3250 17796
rect 3270 17702 3274 17796
rect 3294 17702 3298 17796
rect 3318 17702 3322 17796
rect 3342 17702 3346 17796
rect 3366 17702 3370 17796
rect 3390 17702 3394 17796
rect 3414 17702 3418 17796
rect 3438 17702 3442 17796
rect 3462 17702 3466 17796
rect 3486 17702 3490 17796
rect 3510 17702 3514 17796
rect 3534 17702 3538 17796
rect 3558 17702 3562 17796
rect 3582 17702 3586 17796
rect 3606 17702 3610 17796
rect 3630 17702 3634 17796
rect 3654 17702 3658 17796
rect 3678 17702 3682 17796
rect 3702 17702 3706 17796
rect 3726 17702 3730 17796
rect 3739 17789 3744 17796
rect 3757 17795 3771 17796
rect 3749 17775 3754 17789
rect 3750 17702 3754 17775
rect 3763 17702 3771 17703
rect -2393 17700 3771 17702
rect -2371 17678 -2366 17700
rect -2348 17678 -2343 17700
rect -2325 17678 -2320 17700
rect -2072 17698 -2036 17699
rect -2072 17692 -2054 17698
rect -2309 17684 -2301 17692
rect -2317 17678 -2309 17684
rect -2092 17683 -2062 17688
rect -2000 17679 -1992 17700
rect -1938 17699 -1906 17700
rect -1920 17698 -1906 17699
rect -1806 17692 -1680 17698
rect -1854 17683 -1806 17688
rect -1655 17684 -1647 17692
rect -1982 17679 -1966 17680
rect -2000 17678 -1966 17679
rect -1846 17678 -1806 17681
rect -1663 17678 -1655 17684
rect -1642 17678 -1637 17700
rect -1619 17678 -1614 17700
rect -1530 17678 -1526 17700
rect -1506 17678 -1502 17700
rect -1482 17678 -1478 17700
rect -1458 17678 -1454 17700
rect -1434 17678 -1430 17700
rect -1410 17678 -1406 17700
rect -1386 17699 -1382 17700
rect -2393 17676 -1389 17678
rect -2371 17654 -2366 17676
rect -2348 17654 -2343 17676
rect -2325 17654 -2320 17676
rect -2000 17674 -1966 17676
rect -2309 17656 -2301 17664
rect -2062 17663 -2054 17670
rect -2092 17656 -2084 17663
rect -2062 17656 -2026 17658
rect -2317 17654 -2309 17656
rect -2062 17654 -2012 17656
rect -2000 17654 -1992 17674
rect -1982 17673 -1966 17674
rect -1846 17672 -1806 17676
rect -1846 17665 -1798 17670
rect -1806 17663 -1798 17665
rect -1854 17661 -1846 17663
rect -1854 17656 -1806 17661
rect -1655 17656 -1647 17664
rect -1864 17654 -1796 17655
rect -1663 17654 -1655 17656
rect -1642 17654 -1637 17676
rect -1619 17654 -1614 17676
rect -1530 17654 -1526 17676
rect -1506 17654 -1502 17676
rect -1482 17654 -1478 17676
rect -1458 17654 -1454 17676
rect -1434 17654 -1430 17676
rect -1410 17654 -1406 17676
rect -1403 17675 -1389 17676
rect -1386 17675 -1379 17699
rect -1386 17654 -1382 17675
rect -1362 17654 -1358 17700
rect -1338 17654 -1334 17700
rect -1314 17654 -1310 17700
rect -1290 17654 -1286 17700
rect -1266 17654 -1262 17700
rect -1242 17654 -1238 17700
rect -1218 17654 -1214 17700
rect -1194 17654 -1190 17700
rect -1170 17654 -1166 17700
rect -1146 17654 -1142 17700
rect -1122 17654 -1118 17700
rect -1098 17654 -1094 17700
rect -1074 17654 -1070 17700
rect -1050 17654 -1046 17700
rect -1026 17675 -1022 17700
rect -2393 17652 -1029 17654
rect -2371 17606 -2366 17652
rect -2348 17606 -2343 17652
rect -2325 17606 -2320 17652
rect -2317 17648 -2309 17652
rect -2062 17648 -2054 17652
rect -2154 17644 -2138 17646
rect -2057 17644 -2054 17648
rect -2292 17638 -2054 17644
rect -2052 17638 -2044 17648
rect -2092 17622 -2062 17624
rect -2094 17618 -2062 17622
rect -2000 17606 -1992 17652
rect -1846 17645 -1806 17652
rect -1663 17648 -1655 17652
rect -1846 17638 -1680 17644
rect -1854 17622 -1806 17624
rect -1854 17618 -1680 17622
rect -1642 17606 -1637 17652
rect -1619 17606 -1614 17652
rect -1530 17606 -1526 17652
rect -1506 17606 -1502 17652
rect -1482 17606 -1478 17652
rect -1458 17606 -1454 17652
rect -1434 17606 -1430 17652
rect -1410 17606 -1406 17652
rect -1386 17606 -1382 17652
rect -1362 17606 -1358 17652
rect -1338 17606 -1334 17652
rect -1314 17606 -1310 17652
rect -1290 17606 -1286 17652
rect -1266 17606 -1262 17652
rect -1242 17606 -1238 17652
rect -1218 17606 -1214 17652
rect -1194 17606 -1190 17652
rect -1170 17606 -1166 17652
rect -1146 17606 -1142 17652
rect -1122 17606 -1118 17652
rect -1098 17606 -1094 17652
rect -1074 17606 -1070 17652
rect -1050 17606 -1046 17652
rect -1043 17651 -1029 17652
rect -1026 17651 -1019 17675
rect -1026 17606 -1022 17651
rect -1002 17606 -998 17700
rect -978 17606 -974 17700
rect -954 17606 -950 17700
rect -930 17606 -926 17700
rect -906 17606 -902 17700
rect -882 17606 -878 17700
rect -858 17606 -854 17700
rect -845 17645 -840 17655
rect -834 17645 -830 17700
rect -835 17631 -830 17645
rect -834 17606 -830 17631
rect -810 17606 -806 17700
rect -786 17606 -782 17700
rect -762 17606 -758 17700
rect -738 17606 -734 17700
rect -714 17606 -710 17700
rect -690 17606 -686 17700
rect -666 17606 -662 17700
rect -642 17606 -638 17700
rect -618 17606 -614 17700
rect -594 17606 -590 17700
rect -570 17606 -566 17700
rect -546 17606 -542 17700
rect -522 17606 -518 17700
rect -498 17606 -494 17700
rect -474 17606 -470 17700
rect -450 17606 -446 17700
rect -426 17606 -422 17700
rect -402 17606 -398 17700
rect -378 17606 -374 17700
rect -354 17606 -350 17700
rect -330 17606 -326 17700
rect -306 17606 -302 17700
rect -282 17606 -278 17700
rect -258 17606 -254 17700
rect -234 17606 -230 17700
rect -210 17606 -206 17700
rect -186 17606 -182 17700
rect -162 17606 -158 17700
rect -138 17606 -134 17700
rect -114 17606 -110 17700
rect -90 17606 -86 17700
rect -66 17606 -62 17700
rect -42 17606 -38 17700
rect -18 17606 -14 17700
rect 6 17606 10 17700
rect 30 17606 34 17700
rect 54 17606 58 17700
rect 78 17606 82 17700
rect 102 17606 106 17700
rect 126 17606 130 17700
rect 150 17606 154 17700
rect 174 17606 178 17700
rect 198 17606 202 17700
rect 222 17606 226 17700
rect 246 17606 250 17700
rect 270 17606 274 17700
rect 294 17606 298 17700
rect 318 17606 322 17700
rect 342 17606 346 17700
rect 366 17606 370 17700
rect 390 17606 394 17700
rect 414 17606 418 17700
rect 438 17606 442 17700
rect 462 17606 466 17700
rect 486 17606 490 17700
rect 510 17606 514 17700
rect 534 17606 538 17700
rect 558 17606 562 17700
rect 582 17606 586 17700
rect 606 17606 610 17700
rect 630 17606 634 17700
rect 654 17606 658 17700
rect 678 17606 682 17700
rect 702 17606 706 17700
rect 726 17606 730 17700
rect 750 17606 754 17700
rect 774 17606 778 17700
rect 798 17606 802 17700
rect 822 17606 826 17700
rect 846 17606 850 17700
rect 870 17606 874 17700
rect 894 17606 898 17700
rect 918 17606 922 17700
rect 942 17606 946 17700
rect 966 17606 970 17700
rect 990 17606 994 17700
rect 1014 17606 1018 17700
rect 1038 17606 1042 17700
rect 1062 17606 1066 17700
rect 1086 17606 1090 17700
rect 1110 17606 1114 17700
rect 1134 17606 1138 17700
rect 1158 17606 1162 17700
rect 1182 17606 1186 17700
rect 1206 17606 1210 17700
rect 1230 17606 1234 17700
rect 1254 17606 1258 17700
rect 1278 17606 1282 17700
rect 1302 17606 1306 17700
rect 1326 17606 1330 17700
rect 1350 17606 1354 17700
rect 1374 17606 1378 17700
rect 1398 17606 1402 17700
rect 1422 17606 1426 17700
rect 1446 17606 1450 17700
rect 1470 17606 1474 17700
rect 1494 17606 1498 17700
rect 1518 17606 1522 17700
rect 1542 17606 1546 17700
rect 1566 17606 1570 17700
rect 1590 17606 1594 17700
rect 1614 17606 1618 17700
rect 1638 17606 1642 17700
rect 1662 17606 1666 17700
rect 1686 17606 1690 17700
rect 1710 17606 1714 17700
rect 1734 17606 1738 17700
rect 1758 17606 1762 17700
rect 1782 17606 1786 17700
rect 1806 17606 1810 17700
rect 1830 17606 1834 17700
rect 1854 17606 1858 17700
rect 1878 17606 1882 17700
rect 1902 17606 1906 17700
rect 1926 17606 1930 17700
rect 1950 17606 1954 17700
rect 1974 17606 1978 17700
rect 1998 17606 2002 17700
rect 2022 17606 2026 17700
rect 2046 17606 2050 17700
rect 2070 17606 2074 17700
rect 2094 17606 2098 17700
rect 2118 17606 2122 17700
rect 2142 17606 2146 17700
rect 2166 17606 2170 17700
rect 2190 17606 2194 17700
rect 2214 17606 2218 17700
rect 2238 17606 2242 17700
rect 2262 17606 2266 17700
rect 2286 17606 2290 17700
rect 2310 17606 2314 17700
rect 2334 17606 2338 17700
rect 2358 17606 2362 17700
rect 2382 17606 2386 17700
rect 2406 17606 2410 17700
rect 2430 17606 2434 17700
rect 2454 17606 2458 17700
rect 2478 17606 2482 17700
rect 2502 17606 2506 17700
rect 2526 17606 2530 17700
rect 2550 17606 2554 17700
rect 2574 17606 2578 17700
rect 2598 17606 2602 17700
rect 2622 17606 2626 17700
rect 2646 17606 2650 17700
rect 2670 17606 2674 17700
rect 2694 17606 2698 17700
rect 2718 17606 2722 17700
rect 2742 17606 2746 17700
rect 2766 17606 2770 17700
rect 2790 17606 2794 17700
rect 2814 17606 2818 17700
rect 2838 17606 2842 17700
rect 2862 17606 2866 17700
rect 2886 17606 2890 17700
rect 2910 17606 2914 17700
rect 2934 17606 2938 17700
rect 2958 17606 2962 17700
rect 2982 17606 2986 17700
rect 3006 17606 3010 17700
rect 3030 17606 3034 17700
rect 3054 17606 3058 17700
rect 3078 17606 3082 17700
rect 3102 17606 3106 17700
rect 3126 17606 3130 17700
rect 3150 17606 3154 17700
rect 3174 17606 3178 17700
rect 3198 17606 3202 17700
rect 3222 17606 3226 17700
rect 3246 17606 3250 17700
rect 3270 17606 3274 17700
rect 3294 17606 3298 17700
rect 3318 17606 3322 17700
rect 3342 17606 3346 17700
rect 3355 17669 3360 17679
rect 3366 17669 3370 17700
rect 3365 17655 3370 17669
rect 3355 17645 3360 17655
rect 3365 17631 3370 17645
rect 3366 17606 3370 17631
rect 3390 17606 3394 17700
rect 3414 17606 3418 17700
rect 3438 17606 3442 17700
rect 3462 17606 3466 17700
rect 3486 17606 3490 17700
rect 3510 17606 3514 17700
rect 3534 17606 3538 17700
rect 3558 17606 3562 17700
rect 3582 17606 3586 17700
rect 3606 17606 3610 17700
rect 3630 17606 3634 17700
rect 3654 17606 3658 17700
rect 3678 17606 3682 17700
rect 3702 17606 3706 17700
rect 3726 17606 3730 17700
rect 3750 17606 3754 17700
rect 3757 17699 3771 17700
rect 3763 17693 3768 17699
rect 3773 17679 3778 17693
rect 3763 17645 3768 17655
rect 3774 17645 3778 17679
rect 3773 17631 3778 17645
rect 3763 17606 3795 17607
rect -2393 17604 3795 17606
rect -2371 17582 -2366 17604
rect -2348 17582 -2343 17604
rect -2325 17582 -2320 17604
rect -2072 17602 -2036 17603
rect -2072 17596 -2054 17602
rect -2309 17588 -2301 17596
rect -2317 17582 -2309 17588
rect -2092 17587 -2062 17592
rect -2000 17583 -1992 17604
rect -1938 17603 -1906 17604
rect -1920 17602 -1906 17603
rect -1806 17596 -1680 17602
rect -1854 17587 -1806 17592
rect -1655 17588 -1647 17596
rect -1982 17583 -1966 17584
rect -2000 17582 -1966 17583
rect -1846 17582 -1806 17585
rect -1663 17582 -1655 17588
rect -1642 17582 -1637 17604
rect -1619 17582 -1614 17604
rect -1530 17582 -1526 17604
rect -1506 17582 -1502 17604
rect -1482 17582 -1478 17604
rect -1458 17582 -1454 17604
rect -1434 17582 -1430 17604
rect -1410 17582 -1406 17604
rect -1386 17582 -1382 17604
rect -1362 17582 -1358 17604
rect -1338 17582 -1334 17604
rect -1314 17582 -1310 17604
rect -1290 17582 -1286 17604
rect -1266 17582 -1262 17604
rect -1242 17582 -1238 17604
rect -1218 17582 -1214 17604
rect -1194 17582 -1190 17604
rect -1170 17582 -1166 17604
rect -1146 17582 -1142 17604
rect -1122 17582 -1118 17604
rect -1098 17582 -1094 17604
rect -1074 17582 -1070 17604
rect -1050 17582 -1046 17604
rect -1026 17582 -1022 17604
rect -1002 17582 -998 17604
rect -978 17582 -974 17604
rect -954 17582 -950 17604
rect -930 17582 -926 17604
rect -906 17582 -902 17604
rect -882 17582 -878 17604
rect -858 17582 -854 17604
rect -834 17582 -830 17604
rect -810 17582 -806 17604
rect -786 17582 -782 17604
rect -762 17582 -758 17604
rect -738 17582 -734 17604
rect -714 17582 -710 17604
rect -690 17582 -686 17604
rect -666 17582 -662 17604
rect -642 17582 -638 17604
rect -618 17582 -614 17604
rect -594 17582 -590 17604
rect -570 17582 -566 17604
rect -546 17582 -542 17604
rect -522 17582 -518 17604
rect -498 17582 -494 17604
rect -474 17582 -470 17604
rect -450 17582 -446 17604
rect -426 17582 -422 17604
rect -402 17582 -398 17604
rect -378 17582 -374 17604
rect -354 17582 -350 17604
rect -330 17582 -326 17604
rect -306 17582 -302 17604
rect -282 17582 -278 17604
rect -258 17582 -254 17604
rect -234 17582 -230 17604
rect -210 17582 -206 17604
rect -186 17582 -182 17604
rect -162 17582 -158 17604
rect -138 17582 -134 17604
rect -114 17582 -110 17604
rect -90 17582 -86 17604
rect -66 17582 -62 17604
rect -42 17582 -38 17604
rect -18 17582 -14 17604
rect 6 17582 10 17604
rect 30 17582 34 17604
rect 54 17582 58 17604
rect 78 17582 82 17604
rect 102 17582 106 17604
rect 126 17582 130 17604
rect 150 17582 154 17604
rect 174 17582 178 17604
rect 198 17582 202 17604
rect 222 17582 226 17604
rect 246 17582 250 17604
rect 270 17582 274 17604
rect 294 17582 298 17604
rect 318 17582 322 17604
rect 342 17582 346 17604
rect 366 17582 370 17604
rect 390 17582 394 17604
rect 414 17582 418 17604
rect 438 17582 442 17604
rect 462 17582 466 17604
rect 486 17582 490 17604
rect 510 17582 514 17604
rect 534 17582 538 17604
rect 558 17582 562 17604
rect 582 17582 586 17604
rect 606 17582 610 17604
rect 630 17582 634 17604
rect 654 17582 658 17604
rect 678 17582 682 17604
rect 702 17582 706 17604
rect 726 17582 730 17604
rect 750 17582 754 17604
rect 774 17582 778 17604
rect 798 17582 802 17604
rect 822 17582 826 17604
rect 846 17582 850 17604
rect 870 17582 874 17604
rect 894 17582 898 17604
rect 918 17582 922 17604
rect 942 17582 946 17604
rect 966 17582 970 17604
rect 990 17582 994 17604
rect 1014 17582 1018 17604
rect 1038 17582 1042 17604
rect 1062 17582 1066 17604
rect 1086 17582 1090 17604
rect 1110 17582 1114 17604
rect 1134 17582 1138 17604
rect 1158 17582 1162 17604
rect 1182 17582 1186 17604
rect 1206 17582 1210 17604
rect 1230 17582 1234 17604
rect 1254 17582 1258 17604
rect 1278 17582 1282 17604
rect 1302 17582 1306 17604
rect 1326 17582 1330 17604
rect 1350 17582 1354 17604
rect 1374 17582 1378 17604
rect 1398 17582 1402 17604
rect 1422 17582 1426 17604
rect 1446 17582 1450 17604
rect 1470 17582 1474 17604
rect 1494 17582 1498 17604
rect 1518 17582 1522 17604
rect 1542 17582 1546 17604
rect 1566 17582 1570 17604
rect 1590 17582 1594 17604
rect 1614 17583 1618 17604
rect 1603 17582 1637 17583
rect -2393 17580 1637 17582
rect -2371 17558 -2366 17580
rect -2348 17558 -2343 17580
rect -2325 17558 -2320 17580
rect -2000 17578 -1966 17580
rect -2309 17560 -2301 17568
rect -2062 17567 -2054 17574
rect -2092 17560 -2084 17567
rect -2062 17560 -2026 17562
rect -2317 17558 -2309 17560
rect -2062 17558 -2012 17560
rect -2000 17558 -1992 17578
rect -1982 17577 -1966 17578
rect -1846 17576 -1806 17580
rect -1846 17569 -1798 17574
rect -1806 17567 -1798 17569
rect -1854 17565 -1846 17567
rect -1854 17560 -1806 17565
rect -1655 17560 -1647 17568
rect -1864 17558 -1796 17559
rect -1663 17558 -1655 17560
rect -1642 17558 -1637 17580
rect -1619 17558 -1614 17580
rect -1530 17558 -1526 17580
rect -1506 17558 -1502 17580
rect -1482 17558 -1478 17580
rect -1458 17558 -1454 17580
rect -1434 17558 -1430 17580
rect -1410 17558 -1406 17580
rect -1386 17558 -1382 17580
rect -1362 17558 -1358 17580
rect -1338 17558 -1334 17580
rect -1314 17558 -1310 17580
rect -1290 17558 -1286 17580
rect -1266 17558 -1262 17580
rect -1242 17558 -1238 17580
rect -1218 17558 -1214 17580
rect -1194 17558 -1190 17580
rect -1170 17558 -1166 17580
rect -1146 17558 -1142 17580
rect -1122 17558 -1118 17580
rect -1098 17558 -1094 17580
rect -1074 17558 -1070 17580
rect -1050 17558 -1046 17580
rect -1026 17558 -1022 17580
rect -1002 17558 -998 17580
rect -978 17558 -974 17580
rect -954 17558 -950 17580
rect -930 17558 -926 17580
rect -906 17558 -902 17580
rect -882 17558 -878 17580
rect -858 17558 -854 17580
rect -834 17559 -830 17580
rect -810 17579 -806 17580
rect -845 17558 -813 17559
rect -2393 17556 -813 17558
rect -2371 17510 -2366 17556
rect -2348 17510 -2343 17556
rect -2325 17510 -2320 17556
rect -2317 17552 -2309 17556
rect -2062 17552 -2054 17556
rect -2154 17548 -2138 17550
rect -2057 17548 -2054 17552
rect -2292 17542 -2054 17548
rect -2052 17542 -2044 17552
rect -2092 17526 -2062 17528
rect -2094 17522 -2062 17526
rect -2000 17510 -1992 17556
rect -1846 17549 -1806 17556
rect -1663 17552 -1655 17556
rect -1846 17542 -1680 17548
rect -1854 17526 -1806 17528
rect -1854 17522 -1680 17526
rect -1979 17510 -1945 17512
rect -1642 17510 -1637 17556
rect -1619 17510 -1614 17556
rect -1530 17510 -1526 17556
rect -1506 17510 -1502 17556
rect -1482 17510 -1478 17556
rect -1458 17510 -1454 17556
rect -1434 17510 -1430 17556
rect -1410 17510 -1406 17556
rect -1386 17510 -1382 17556
rect -1362 17510 -1358 17556
rect -1338 17510 -1334 17556
rect -1314 17510 -1310 17556
rect -1290 17510 -1286 17556
rect -1266 17510 -1262 17556
rect -1242 17510 -1238 17556
rect -1218 17510 -1214 17556
rect -1194 17510 -1190 17556
rect -1170 17510 -1166 17556
rect -1146 17510 -1142 17556
rect -1122 17510 -1118 17556
rect -1098 17510 -1094 17556
rect -1074 17510 -1070 17556
rect -1050 17510 -1046 17556
rect -1026 17510 -1022 17556
rect -1002 17510 -998 17556
rect -978 17510 -974 17556
rect -954 17510 -950 17556
rect -930 17510 -926 17556
rect -906 17510 -902 17556
rect -882 17510 -878 17556
rect -858 17510 -854 17556
rect -845 17549 -840 17556
rect -834 17549 -830 17556
rect -827 17555 -813 17556
rect -810 17555 -803 17579
rect -835 17535 -830 17549
rect -834 17510 -830 17535
rect -810 17510 -806 17555
rect -786 17510 -782 17580
rect -762 17510 -758 17580
rect -738 17510 -734 17580
rect -714 17510 -710 17580
rect -690 17510 -686 17580
rect -666 17510 -662 17580
rect -642 17510 -638 17580
rect -618 17510 -614 17580
rect -594 17510 -590 17580
rect -570 17510 -566 17580
rect -546 17510 -542 17580
rect -522 17510 -518 17580
rect -498 17510 -494 17580
rect -474 17510 -470 17580
rect -450 17510 -446 17580
rect -426 17510 -422 17580
rect -402 17510 -398 17580
rect -378 17510 -374 17580
rect -354 17510 -350 17580
rect -330 17510 -326 17580
rect -306 17510 -302 17580
rect -282 17510 -278 17580
rect -258 17510 -254 17580
rect -234 17510 -230 17580
rect -210 17510 -206 17580
rect -186 17510 -182 17580
rect -162 17510 -158 17580
rect -138 17510 -134 17580
rect -114 17510 -110 17580
rect -90 17510 -86 17580
rect -66 17510 -62 17580
rect -42 17510 -38 17580
rect -18 17510 -14 17580
rect 6 17510 10 17580
rect 30 17510 34 17580
rect 54 17510 58 17580
rect 78 17510 82 17580
rect 102 17510 106 17580
rect 126 17510 130 17580
rect 150 17510 154 17580
rect 174 17510 178 17580
rect 198 17510 202 17580
rect 222 17510 226 17580
rect 246 17510 250 17580
rect 270 17510 274 17580
rect 294 17510 298 17580
rect 318 17510 322 17580
rect 342 17510 346 17580
rect 366 17510 370 17580
rect 390 17510 394 17580
rect 414 17510 418 17580
rect 438 17510 442 17580
rect 462 17510 466 17580
rect 486 17510 490 17580
rect 510 17510 514 17580
rect 534 17510 538 17580
rect 558 17510 562 17580
rect 582 17510 586 17580
rect 606 17510 610 17580
rect 630 17510 634 17580
rect 654 17510 658 17580
rect 678 17510 682 17580
rect 702 17510 706 17580
rect 726 17510 730 17580
rect 750 17510 754 17580
rect 774 17510 778 17580
rect 798 17510 802 17580
rect 822 17510 826 17580
rect 846 17510 850 17580
rect 870 17510 874 17580
rect 894 17510 898 17580
rect 918 17510 922 17580
rect 942 17510 946 17580
rect 966 17510 970 17580
rect 990 17510 994 17580
rect 1014 17510 1018 17580
rect 1038 17510 1042 17580
rect 1062 17510 1066 17580
rect 1086 17510 1090 17580
rect 1110 17510 1114 17580
rect 1134 17510 1138 17580
rect 1158 17510 1162 17580
rect 1182 17510 1186 17580
rect 1206 17510 1210 17580
rect 1230 17510 1234 17580
rect 1254 17510 1258 17580
rect 1278 17510 1282 17580
rect 1302 17510 1306 17580
rect 1326 17510 1330 17580
rect 1350 17510 1354 17580
rect 1374 17510 1378 17580
rect 1398 17510 1402 17580
rect 1422 17510 1426 17580
rect 1446 17510 1450 17580
rect 1470 17510 1474 17580
rect 1494 17510 1498 17580
rect 1518 17510 1522 17580
rect 1542 17510 1546 17580
rect 1566 17510 1570 17580
rect 1590 17510 1594 17580
rect 1603 17573 1608 17580
rect 1614 17573 1618 17580
rect 1613 17559 1618 17573
rect 1614 17510 1618 17559
rect 1638 17510 1642 17604
rect 1662 17510 1666 17604
rect 1686 17510 1690 17604
rect 1710 17510 1714 17604
rect 1734 17510 1738 17604
rect 1758 17510 1762 17604
rect 1782 17510 1786 17604
rect 1806 17510 1810 17604
rect 1830 17510 1834 17604
rect 1854 17510 1858 17604
rect 1878 17510 1882 17604
rect 1902 17510 1906 17604
rect 1926 17510 1930 17604
rect 1950 17510 1954 17604
rect 1974 17510 1978 17604
rect 1998 17510 2002 17604
rect 2022 17510 2026 17604
rect 2046 17510 2050 17604
rect 2070 17510 2074 17604
rect 2094 17510 2098 17604
rect 2118 17510 2122 17604
rect 2142 17510 2146 17604
rect 2166 17510 2170 17604
rect 2190 17510 2194 17604
rect 2214 17510 2218 17604
rect 2238 17510 2242 17604
rect 2262 17510 2266 17604
rect 2286 17510 2290 17604
rect 2310 17510 2314 17604
rect 2334 17510 2338 17604
rect 2358 17510 2362 17604
rect 2382 17510 2386 17604
rect 2406 17510 2410 17604
rect 2430 17510 2434 17604
rect 2454 17510 2458 17604
rect 2478 17510 2482 17604
rect 2502 17510 2506 17604
rect 2526 17510 2530 17604
rect 2550 17510 2554 17604
rect 2574 17510 2578 17604
rect 2598 17510 2602 17604
rect 2622 17510 2626 17604
rect 2646 17510 2650 17604
rect 2670 17510 2674 17604
rect 2694 17510 2698 17604
rect 2718 17510 2722 17604
rect 2742 17510 2746 17604
rect 2766 17510 2770 17604
rect 2790 17510 2794 17604
rect 2814 17510 2818 17604
rect 2838 17510 2842 17604
rect 2862 17510 2866 17604
rect 2886 17510 2890 17604
rect 2910 17510 2914 17604
rect 2934 17510 2938 17604
rect 2958 17510 2962 17604
rect 2982 17510 2986 17604
rect 3006 17510 3010 17604
rect 3030 17510 3034 17604
rect 3054 17510 3058 17604
rect 3078 17510 3082 17604
rect 3102 17510 3106 17604
rect 3126 17510 3130 17604
rect 3150 17510 3154 17604
rect 3174 17510 3178 17604
rect 3198 17510 3202 17604
rect 3222 17510 3226 17604
rect 3246 17510 3250 17604
rect 3270 17510 3274 17604
rect 3294 17510 3298 17604
rect 3318 17510 3322 17604
rect 3342 17510 3346 17604
rect 3366 17510 3370 17604
rect 3390 17603 3394 17604
rect 3390 17555 3397 17603
rect 3390 17510 3394 17555
rect 3414 17510 3418 17604
rect 3438 17510 3442 17604
rect 3462 17510 3466 17604
rect 3486 17510 3490 17604
rect 3510 17510 3514 17604
rect 3534 17510 3538 17604
rect 3558 17510 3562 17604
rect 3582 17510 3586 17604
rect 3606 17510 3610 17604
rect 3630 17510 3634 17604
rect 3654 17510 3658 17604
rect 3678 17510 3682 17604
rect 3702 17510 3706 17604
rect 3726 17510 3730 17604
rect 3750 17510 3754 17604
rect 3763 17597 3768 17604
rect 3781 17603 3795 17604
rect 3773 17583 3778 17597
rect 3774 17510 3778 17583
rect 3787 17510 3795 17511
rect -2393 17508 3795 17510
rect -2371 17462 -2366 17508
rect -2348 17462 -2343 17508
rect -2325 17462 -2320 17508
rect -2080 17507 -1906 17508
rect -2080 17506 -2036 17507
rect -2080 17500 -2054 17506
rect -2309 17492 -2301 17498
rect -2317 17482 -2309 17492
rect -2070 17491 -2040 17498
rect -2054 17483 -2040 17486
rect -2000 17481 -1992 17507
rect -1920 17506 -1906 17507
rect -1850 17500 -1846 17508
rect -1840 17500 -1792 17508
rect -1969 17488 -1966 17497
rect -1850 17493 -1802 17498
rect -1906 17491 -1802 17493
rect -1655 17492 -1647 17498
rect -1906 17490 -1850 17491
rect -1846 17483 -1802 17489
rect -1663 17482 -1655 17492
rect -1860 17481 -1798 17482
rect -2078 17474 -2070 17481
rect -2309 17464 -2301 17470
rect -2317 17462 -2309 17464
rect -2154 17462 -2145 17472
rect -2044 17471 -2040 17476
rect -2028 17474 -1945 17481
rect -1929 17474 -1794 17481
rect -2070 17464 -2040 17471
rect -2044 17462 -2028 17464
rect -2000 17462 -1992 17474
rect -1860 17473 -1798 17474
rect -1850 17464 -1802 17471
rect -1655 17464 -1647 17470
rect -1978 17462 -1942 17463
rect -1663 17462 -1655 17464
rect -1642 17462 -1637 17508
rect -1619 17462 -1614 17508
rect -1530 17462 -1526 17508
rect -1506 17462 -1502 17508
rect -1482 17462 -1478 17508
rect -1458 17462 -1454 17508
rect -1434 17462 -1430 17508
rect -1410 17462 -1406 17508
rect -1386 17462 -1382 17508
rect -1362 17462 -1358 17508
rect -1338 17462 -1334 17508
rect -1314 17462 -1310 17508
rect -1290 17462 -1286 17508
rect -1266 17462 -1262 17508
rect -1242 17463 -1238 17508
rect -1253 17462 -1219 17463
rect -2393 17460 -1219 17462
rect -2371 17366 -2366 17460
rect -2348 17366 -2343 17460
rect -2325 17422 -2320 17460
rect -2317 17454 -2309 17460
rect -2145 17456 -2138 17460
rect -2070 17456 -2054 17460
rect -2078 17447 -2054 17454
rect -2062 17422 -2032 17423
rect -2000 17422 -1992 17460
rect -1846 17456 -1802 17460
rect -1846 17446 -1792 17455
rect -1663 17454 -1655 17460
rect -1942 17424 -1937 17436
rect -1850 17433 -1822 17434
rect -1850 17429 -1802 17433
rect -2325 17414 -2317 17422
rect -2062 17420 -1961 17422
rect -2325 17394 -2320 17414
rect -2317 17406 -2309 17414
rect -2062 17407 -2040 17418
rect -2032 17413 -1961 17420
rect -1947 17414 -1942 17422
rect -1842 17420 -1794 17423
rect -2070 17402 -2022 17406
rect -2325 17380 -2317 17394
rect -2072 17386 -2032 17387
rect -2102 17380 -2032 17386
rect -2325 17366 -2320 17380
rect -2317 17378 -2309 17380
rect -2309 17366 -2301 17378
rect -2070 17371 -2062 17376
rect -2000 17366 -1992 17413
rect -1942 17412 -1937 17414
rect -1932 17404 -1927 17412
rect -1912 17409 -1896 17415
rect -1842 17407 -1802 17418
rect -1671 17414 -1663 17422
rect -1663 17406 -1655 17414
rect -1850 17402 -1680 17406
rect -1924 17388 -1921 17390
rect -1806 17380 -1680 17386
rect -1671 17380 -1663 17394
rect -1663 17378 -1655 17380
rect -1854 17371 -1806 17376
rect -1974 17366 -1964 17367
rect -1960 17366 -1944 17368
rect -1842 17366 -1806 17369
rect -1655 17366 -1647 17378
rect -1642 17366 -1637 17460
rect -1619 17366 -1614 17460
rect -1530 17366 -1526 17460
rect -1506 17366 -1502 17460
rect -1482 17366 -1478 17460
rect -1458 17366 -1454 17460
rect -1434 17366 -1430 17460
rect -1410 17366 -1406 17460
rect -1386 17366 -1382 17460
rect -1362 17366 -1358 17460
rect -1338 17366 -1334 17460
rect -1314 17366 -1310 17460
rect -1290 17366 -1286 17460
rect -1266 17366 -1262 17460
rect -1253 17453 -1248 17460
rect -1242 17453 -1238 17460
rect -1243 17439 -1238 17453
rect -1242 17366 -1238 17439
rect -1218 17387 -1214 17508
rect -2393 17364 -1221 17366
rect -2371 17342 -2366 17364
rect -2348 17342 -2343 17364
rect -2325 17352 -2317 17364
rect -2325 17342 -2320 17352
rect -2317 17350 -2309 17352
rect -2062 17351 -2032 17358
rect -2309 17342 -2301 17350
rect -2070 17344 -2062 17351
rect -2000 17346 -1992 17364
rect -1974 17362 -1944 17364
rect -1960 17361 -1944 17362
rect -1842 17360 -1806 17364
rect -1842 17353 -1798 17358
rect -1806 17351 -1798 17353
rect -1671 17352 -1663 17364
rect -1854 17349 -1842 17351
rect -1663 17350 -1655 17352
rect -2062 17342 -2036 17344
rect -2393 17340 -2036 17342
rect -2032 17342 -2012 17344
rect -2004 17342 -1974 17346
rect -1854 17344 -1806 17349
rect -1864 17342 -1796 17343
rect -1655 17342 -1647 17350
rect -1642 17342 -1637 17364
rect -1619 17342 -1614 17364
rect -1530 17342 -1526 17364
rect -1506 17342 -1502 17364
rect -1482 17342 -1478 17364
rect -1458 17342 -1454 17364
rect -1434 17342 -1430 17364
rect -1410 17342 -1406 17364
rect -1386 17342 -1382 17364
rect -1362 17342 -1358 17364
rect -1338 17342 -1334 17364
rect -1314 17342 -1310 17364
rect -1290 17342 -1286 17364
rect -1266 17342 -1262 17364
rect -1242 17342 -1238 17364
rect -1235 17363 -1221 17364
rect -1218 17363 -1211 17387
rect -1218 17342 -1214 17363
rect -1194 17342 -1190 17508
rect -1170 17342 -1166 17508
rect -1146 17342 -1142 17508
rect -1122 17342 -1118 17508
rect -1098 17342 -1094 17508
rect -1074 17342 -1070 17508
rect -1050 17342 -1046 17508
rect -1026 17342 -1022 17508
rect -1002 17342 -998 17508
rect -978 17342 -974 17508
rect -954 17342 -950 17508
rect -930 17342 -926 17508
rect -906 17342 -902 17508
rect -882 17342 -878 17508
rect -858 17342 -854 17508
rect -845 17429 -840 17439
rect -834 17429 -830 17508
rect -835 17415 -830 17429
rect -834 17342 -830 17415
rect -810 17483 -806 17508
rect -810 17459 -803 17483
rect -810 17363 -806 17459
rect -2032 17340 -813 17342
rect -2371 17294 -2366 17340
rect -2348 17294 -2343 17340
rect -2325 17336 -2320 17340
rect -2309 17338 -2301 17340
rect -2317 17336 -2309 17338
rect -2325 17324 -2317 17336
rect -2052 17334 -2036 17336
rect -2052 17332 -2032 17334
rect -2062 17326 -2032 17332
rect -2325 17294 -2320 17324
rect -2317 17322 -2309 17324
rect -2092 17310 -2062 17312
rect -2094 17306 -2062 17310
rect -2000 17294 -1992 17340
rect -1904 17333 -1874 17340
rect -1842 17333 -1806 17340
rect -1655 17338 -1647 17340
rect -1663 17336 -1655 17338
rect -1842 17326 -1680 17332
rect -1671 17324 -1663 17336
rect -1663 17322 -1655 17324
rect -1854 17310 -1806 17312
rect -1854 17306 -1680 17310
rect -1642 17294 -1637 17340
rect -1619 17294 -1614 17340
rect -1530 17294 -1526 17340
rect -1506 17294 -1502 17340
rect -1482 17294 -1478 17340
rect -1458 17294 -1454 17340
rect -1434 17294 -1430 17340
rect -1410 17294 -1406 17340
rect -1386 17294 -1382 17340
rect -1362 17294 -1358 17340
rect -1338 17294 -1334 17340
rect -1314 17294 -1310 17340
rect -1290 17294 -1286 17340
rect -1266 17294 -1262 17340
rect -1242 17294 -1238 17340
rect -1218 17294 -1214 17340
rect -1194 17294 -1190 17340
rect -1170 17294 -1166 17340
rect -1146 17294 -1142 17340
rect -1122 17294 -1118 17340
rect -1098 17294 -1094 17340
rect -1074 17294 -1070 17340
rect -1050 17294 -1046 17340
rect -1026 17294 -1022 17340
rect -1002 17294 -998 17340
rect -978 17294 -974 17340
rect -954 17294 -950 17340
rect -930 17294 -926 17340
rect -906 17294 -902 17340
rect -882 17294 -878 17340
rect -858 17294 -854 17340
rect -834 17294 -830 17340
rect -827 17339 -813 17340
rect -810 17339 -803 17363
rect -810 17294 -806 17339
rect -786 17294 -782 17508
rect -762 17294 -758 17508
rect -738 17294 -734 17508
rect -714 17294 -710 17508
rect -690 17294 -686 17508
rect -666 17294 -662 17508
rect -642 17294 -638 17508
rect -618 17294 -614 17508
rect -594 17294 -590 17508
rect -570 17294 -566 17508
rect -546 17294 -542 17508
rect -522 17294 -518 17508
rect -498 17294 -494 17508
rect -474 17294 -470 17508
rect -450 17294 -446 17508
rect -426 17294 -422 17508
rect -402 17294 -398 17508
rect -378 17294 -374 17508
rect -354 17294 -350 17508
rect -330 17294 -326 17508
rect -306 17294 -302 17508
rect -282 17294 -278 17508
rect -258 17294 -254 17508
rect -245 17333 -240 17343
rect -234 17333 -230 17508
rect -235 17319 -230 17333
rect -234 17294 -230 17319
rect -210 17294 -206 17508
rect -186 17294 -182 17508
rect -162 17294 -158 17508
rect -138 17294 -134 17508
rect -114 17294 -110 17508
rect -90 17294 -86 17508
rect -66 17294 -62 17508
rect -42 17294 -38 17508
rect -18 17294 -14 17508
rect 6 17294 10 17508
rect 30 17294 34 17508
rect 54 17294 58 17508
rect 78 17294 82 17508
rect 102 17294 106 17508
rect 126 17294 130 17508
rect 150 17294 154 17508
rect 174 17294 178 17508
rect 198 17294 202 17508
rect 222 17294 226 17508
rect 246 17294 250 17508
rect 270 17294 274 17508
rect 294 17294 298 17508
rect 318 17294 322 17508
rect 342 17294 346 17508
rect 366 17294 370 17508
rect 390 17294 394 17508
rect 414 17294 418 17508
rect 438 17294 442 17508
rect 462 17294 466 17508
rect 486 17294 490 17508
rect 510 17294 514 17508
rect 534 17294 538 17508
rect 558 17294 562 17508
rect 582 17294 586 17508
rect 606 17294 610 17508
rect 630 17294 634 17508
rect 654 17294 658 17508
rect 678 17294 682 17508
rect 702 17294 706 17508
rect 726 17294 730 17508
rect 750 17294 754 17508
rect 774 17294 778 17508
rect 798 17294 802 17508
rect 822 17294 826 17508
rect 846 17294 850 17508
rect 870 17294 874 17508
rect 894 17294 898 17508
rect 918 17294 922 17508
rect 942 17294 946 17508
rect 966 17294 970 17508
rect 990 17294 994 17508
rect 1014 17294 1018 17508
rect 1038 17294 1042 17508
rect 1062 17294 1066 17508
rect 1086 17294 1090 17508
rect 1110 17294 1114 17508
rect 1134 17294 1138 17508
rect 1158 17294 1162 17508
rect 1182 17294 1186 17508
rect 1206 17294 1210 17508
rect 1230 17294 1234 17508
rect 1254 17294 1258 17508
rect 1278 17294 1282 17508
rect 1302 17294 1306 17508
rect 1326 17294 1330 17508
rect 1350 17294 1354 17508
rect 1374 17294 1378 17508
rect 1398 17294 1402 17508
rect 1422 17294 1426 17508
rect 1446 17294 1450 17508
rect 1470 17294 1474 17508
rect 1494 17294 1498 17508
rect 1518 17294 1522 17508
rect 1542 17294 1546 17508
rect 1566 17294 1570 17508
rect 1590 17294 1594 17508
rect 1603 17357 1608 17367
rect 1614 17357 1618 17508
rect 1613 17343 1618 17357
rect 1638 17507 1642 17508
rect 1638 17483 1645 17507
rect 1603 17333 1608 17343
rect 1613 17319 1618 17333
rect 1614 17294 1618 17319
rect 1638 17294 1642 17483
rect 1662 17294 1666 17508
rect 1686 17294 1690 17508
rect 1710 17294 1714 17508
rect 1734 17294 1738 17508
rect 1758 17294 1762 17508
rect 1782 17294 1786 17508
rect 1806 17294 1810 17508
rect 1830 17294 1834 17508
rect 1854 17294 1858 17508
rect 1878 17294 1882 17508
rect 1902 17294 1906 17508
rect 1926 17294 1930 17508
rect 1950 17294 1954 17508
rect 1974 17294 1978 17508
rect 1998 17294 2002 17508
rect 2022 17294 2026 17508
rect 2046 17294 2050 17508
rect 2070 17294 2074 17508
rect 2094 17294 2098 17508
rect 2118 17294 2122 17508
rect 2142 17294 2146 17508
rect 2166 17294 2170 17508
rect 2190 17294 2194 17508
rect 2214 17294 2218 17508
rect 2238 17294 2242 17508
rect 2262 17294 2266 17508
rect 2286 17294 2290 17508
rect 2310 17294 2314 17508
rect 2334 17294 2338 17508
rect 2358 17294 2362 17508
rect 2382 17294 2386 17508
rect 2406 17294 2410 17508
rect 2430 17294 2434 17508
rect 2454 17294 2458 17508
rect 2478 17294 2482 17508
rect 2502 17294 2506 17508
rect 2526 17294 2530 17508
rect 2550 17294 2554 17508
rect 2574 17294 2578 17508
rect 2598 17294 2602 17508
rect 2622 17294 2626 17508
rect 2646 17294 2650 17508
rect 2670 17294 2674 17508
rect 2694 17294 2698 17508
rect 2718 17294 2722 17508
rect 2742 17294 2746 17508
rect 2766 17294 2770 17508
rect 2790 17294 2794 17508
rect 2814 17294 2818 17508
rect 2838 17294 2842 17508
rect 2862 17294 2866 17508
rect 2886 17294 2890 17508
rect 2910 17294 2914 17508
rect 2934 17294 2938 17508
rect 2958 17294 2962 17508
rect 2982 17294 2986 17508
rect 3006 17294 3010 17508
rect 3030 17294 3034 17508
rect 3054 17294 3058 17508
rect 3078 17294 3082 17508
rect 3102 17294 3106 17508
rect 3126 17294 3130 17508
rect 3150 17294 3154 17508
rect 3174 17294 3178 17508
rect 3198 17294 3202 17508
rect 3222 17294 3226 17508
rect 3246 17294 3250 17508
rect 3270 17294 3274 17508
rect 3294 17294 3298 17508
rect 3318 17294 3322 17508
rect 3342 17294 3346 17508
rect 3366 17294 3370 17508
rect 3390 17294 3394 17508
rect 3414 17294 3418 17508
rect 3438 17294 3442 17508
rect 3462 17294 3466 17508
rect 3486 17294 3490 17508
rect 3510 17294 3514 17508
rect 3534 17294 3538 17508
rect 3558 17294 3562 17508
rect 3582 17294 3586 17508
rect 3606 17294 3610 17508
rect 3630 17294 3634 17508
rect 3654 17294 3658 17508
rect 3678 17294 3682 17508
rect 3702 17294 3706 17508
rect 3726 17294 3730 17508
rect 3750 17294 3754 17508
rect 3774 17294 3778 17508
rect 3781 17507 3795 17508
rect 3787 17501 3792 17507
rect 3797 17487 3802 17501
rect 3798 17294 3802 17487
rect 3811 17381 3816 17391
rect 3821 17367 3826 17381
rect 3811 17333 3816 17343
rect 3822 17333 3826 17367
rect 3821 17319 3826 17333
rect 3811 17294 3843 17295
rect -2393 17292 3843 17294
rect -2371 17270 -2366 17292
rect -2348 17270 -2343 17292
rect -2325 17270 -2320 17292
rect -2072 17290 -2036 17291
rect -2072 17284 -2054 17290
rect -2309 17276 -2301 17284
rect -2317 17270 -2309 17276
rect -2092 17275 -2062 17280
rect -2000 17271 -1992 17292
rect -1938 17291 -1906 17292
rect -1920 17290 -1906 17291
rect -1806 17284 -1680 17290
rect -1854 17275 -1806 17280
rect -1655 17276 -1647 17284
rect -1982 17271 -1966 17272
rect -2000 17270 -1966 17271
rect -1846 17270 -1806 17273
rect -1663 17270 -1655 17276
rect -1642 17270 -1637 17292
rect -1619 17270 -1614 17292
rect -1530 17271 -1526 17292
rect -1541 17270 -1507 17271
rect -2393 17268 -1507 17270
rect -2371 17246 -2366 17268
rect -2348 17246 -2343 17268
rect -2325 17246 -2320 17268
rect -2000 17266 -1966 17268
rect -2309 17248 -2301 17256
rect -2062 17255 -2054 17262
rect -2092 17248 -2084 17255
rect -2062 17248 -2026 17250
rect -2317 17246 -2309 17248
rect -2062 17246 -2012 17248
rect -2000 17246 -1992 17266
rect -1982 17265 -1966 17266
rect -1846 17264 -1806 17268
rect -1846 17257 -1798 17262
rect -1806 17255 -1798 17257
rect -1854 17253 -1846 17255
rect -1854 17248 -1806 17253
rect -1655 17248 -1647 17256
rect -1864 17246 -1796 17247
rect -1663 17246 -1655 17248
rect -1642 17246 -1637 17268
rect -1619 17246 -1614 17268
rect -1541 17261 -1536 17268
rect -1530 17261 -1526 17268
rect -1531 17247 -1526 17261
rect -1541 17246 -1507 17247
rect -1506 17246 -1502 17292
rect -1482 17246 -1478 17292
rect -1458 17246 -1454 17292
rect -1434 17246 -1430 17292
rect -1410 17246 -1406 17292
rect -1386 17246 -1382 17292
rect -1362 17246 -1358 17292
rect -1338 17246 -1334 17292
rect -1314 17246 -1310 17292
rect -1290 17246 -1286 17292
rect -1266 17246 -1262 17292
rect -1242 17246 -1238 17292
rect -1218 17246 -1214 17292
rect -1194 17246 -1190 17292
rect -1170 17246 -1166 17292
rect -1146 17246 -1142 17292
rect -1122 17246 -1118 17292
rect -1098 17246 -1094 17292
rect -1074 17246 -1070 17292
rect -1050 17246 -1046 17292
rect -1026 17246 -1022 17292
rect -1002 17246 -998 17292
rect -978 17246 -974 17292
rect -954 17246 -950 17292
rect -930 17246 -926 17292
rect -906 17246 -902 17292
rect -882 17246 -878 17292
rect -858 17246 -854 17292
rect -834 17246 -830 17292
rect -810 17246 -806 17292
rect -786 17246 -782 17292
rect -762 17246 -758 17292
rect -738 17246 -734 17292
rect -714 17246 -710 17292
rect -690 17246 -686 17292
rect -666 17246 -662 17292
rect -642 17246 -638 17292
rect -618 17246 -614 17292
rect -594 17246 -590 17292
rect -570 17246 -566 17292
rect -546 17246 -542 17292
rect -522 17246 -518 17292
rect -498 17246 -494 17292
rect -474 17246 -470 17292
rect -450 17246 -446 17292
rect -426 17246 -422 17292
rect -402 17246 -398 17292
rect -378 17246 -374 17292
rect -354 17246 -350 17292
rect -330 17246 -326 17292
rect -306 17246 -302 17292
rect -282 17246 -278 17292
rect -258 17246 -254 17292
rect -234 17247 -230 17292
rect -210 17267 -206 17292
rect -245 17246 -213 17247
rect -2393 17244 -213 17246
rect -2371 17198 -2366 17244
rect -2348 17198 -2343 17244
rect -2325 17198 -2320 17244
rect -2317 17240 -2309 17244
rect -2062 17240 -2054 17244
rect -2154 17236 -2138 17238
rect -2057 17236 -2054 17240
rect -2292 17230 -2054 17236
rect -2052 17230 -2044 17240
rect -2092 17214 -2062 17216
rect -2094 17210 -2062 17214
rect -2000 17198 -1992 17244
rect -1846 17237 -1806 17244
rect -1663 17240 -1655 17244
rect -1846 17230 -1680 17236
rect -1854 17214 -1806 17216
rect -1854 17210 -1680 17214
rect -1642 17198 -1637 17244
rect -1619 17198 -1614 17244
rect -1541 17237 -1536 17244
rect -1531 17223 -1526 17237
rect -1530 17198 -1526 17223
rect -1506 17198 -1502 17244
rect -1482 17198 -1478 17244
rect -1458 17198 -1454 17244
rect -1434 17198 -1430 17244
rect -1410 17198 -1406 17244
rect -1386 17198 -1382 17244
rect -1362 17198 -1358 17244
rect -1338 17198 -1334 17244
rect -1314 17198 -1310 17244
rect -1290 17198 -1286 17244
rect -1266 17198 -1262 17244
rect -1242 17198 -1238 17244
rect -1218 17198 -1214 17244
rect -1194 17198 -1190 17244
rect -1170 17198 -1166 17244
rect -1146 17198 -1142 17244
rect -1122 17198 -1118 17244
rect -1098 17198 -1094 17244
rect -1074 17198 -1070 17244
rect -1050 17198 -1046 17244
rect -1026 17198 -1022 17244
rect -1002 17198 -998 17244
rect -978 17198 -974 17244
rect -954 17198 -950 17244
rect -930 17198 -926 17244
rect -906 17198 -902 17244
rect -882 17198 -878 17244
rect -858 17198 -854 17244
rect -834 17198 -830 17244
rect -810 17198 -806 17244
rect -786 17198 -782 17244
rect -762 17198 -758 17244
rect -738 17198 -734 17244
rect -714 17198 -710 17244
rect -690 17198 -686 17244
rect -666 17198 -662 17244
rect -642 17198 -638 17244
rect -618 17198 -614 17244
rect -594 17198 -590 17244
rect -570 17198 -566 17244
rect -546 17198 -542 17244
rect -522 17198 -518 17244
rect -498 17198 -494 17244
rect -474 17198 -470 17244
rect -450 17198 -446 17244
rect -426 17198 -422 17244
rect -402 17198 -398 17244
rect -378 17198 -374 17244
rect -354 17198 -350 17244
rect -330 17198 -326 17244
rect -306 17198 -302 17244
rect -282 17198 -278 17244
rect -258 17198 -254 17244
rect -245 17237 -240 17244
rect -234 17237 -230 17244
rect -227 17243 -213 17244
rect -210 17243 -203 17267
rect -235 17223 -230 17237
rect -245 17213 -240 17223
rect -235 17199 -230 17213
rect -234 17198 -230 17199
rect -210 17198 -206 17243
rect -186 17198 -182 17292
rect -162 17198 -158 17292
rect -138 17198 -134 17292
rect -114 17198 -110 17292
rect -90 17198 -86 17292
rect -66 17198 -62 17292
rect -42 17198 -38 17292
rect -18 17198 -14 17292
rect 6 17198 10 17292
rect 30 17198 34 17292
rect 54 17198 58 17292
rect 78 17198 82 17292
rect 102 17198 106 17292
rect 126 17198 130 17292
rect 150 17198 154 17292
rect 174 17198 178 17292
rect 198 17198 202 17292
rect 222 17198 226 17292
rect 246 17198 250 17292
rect 270 17198 274 17292
rect 294 17198 298 17292
rect 318 17198 322 17292
rect 342 17198 346 17292
rect 366 17198 370 17292
rect 390 17198 394 17292
rect 414 17198 418 17292
rect 438 17198 442 17292
rect 462 17198 466 17292
rect 486 17198 490 17292
rect 510 17198 514 17292
rect 534 17198 538 17292
rect 558 17198 562 17292
rect 582 17198 586 17292
rect 606 17198 610 17292
rect 630 17198 634 17292
rect 654 17198 658 17292
rect 678 17198 682 17292
rect 702 17198 706 17292
rect 726 17198 730 17292
rect 750 17198 754 17292
rect 774 17198 778 17292
rect 798 17198 802 17292
rect 822 17198 826 17292
rect 846 17198 850 17292
rect 870 17198 874 17292
rect 894 17198 898 17292
rect 918 17198 922 17292
rect 942 17198 946 17292
rect 966 17198 970 17292
rect 990 17198 994 17292
rect 1014 17198 1018 17292
rect 1038 17198 1042 17292
rect 1062 17198 1066 17292
rect 1086 17198 1090 17292
rect 1110 17198 1114 17292
rect 1134 17198 1138 17292
rect 1158 17198 1162 17292
rect 1182 17198 1186 17292
rect 1206 17198 1210 17292
rect 1230 17198 1234 17292
rect 1254 17198 1258 17292
rect 1278 17198 1282 17292
rect 1302 17198 1306 17292
rect 1326 17198 1330 17292
rect 1350 17198 1354 17292
rect 1374 17198 1378 17292
rect 1398 17198 1402 17292
rect 1422 17198 1426 17292
rect 1446 17198 1450 17292
rect 1470 17198 1474 17292
rect 1494 17198 1498 17292
rect 1518 17198 1522 17292
rect 1542 17198 1546 17292
rect 1566 17198 1570 17292
rect 1590 17198 1594 17292
rect 1614 17198 1618 17292
rect 1638 17291 1642 17292
rect 1638 17243 1645 17291
rect 1638 17198 1642 17243
rect 1662 17198 1666 17292
rect 1686 17198 1690 17292
rect 1710 17198 1714 17292
rect 1734 17198 1738 17292
rect 1758 17198 1762 17292
rect 1782 17198 1786 17292
rect 1806 17198 1810 17292
rect 1830 17198 1834 17292
rect 1854 17198 1858 17292
rect 1878 17198 1882 17292
rect 1902 17198 1906 17292
rect 1926 17198 1930 17292
rect 1950 17198 1954 17292
rect 1974 17198 1978 17292
rect 1998 17198 2002 17292
rect 2022 17198 2026 17292
rect 2046 17198 2050 17292
rect 2070 17198 2074 17292
rect 2094 17198 2098 17292
rect 2118 17198 2122 17292
rect 2142 17198 2146 17292
rect 2166 17198 2170 17292
rect 2190 17198 2194 17292
rect 2214 17198 2218 17292
rect 2238 17198 2242 17292
rect 2262 17198 2266 17292
rect 2286 17198 2290 17292
rect 2310 17198 2314 17292
rect 2334 17198 2338 17292
rect 2358 17198 2362 17292
rect 2382 17198 2386 17292
rect 2406 17198 2410 17292
rect 2430 17198 2434 17292
rect 2454 17198 2458 17292
rect 2478 17198 2482 17292
rect 2502 17198 2506 17292
rect 2526 17198 2530 17292
rect 2550 17198 2554 17292
rect 2574 17198 2578 17292
rect 2598 17198 2602 17292
rect 2622 17198 2626 17292
rect 2646 17198 2650 17292
rect 2670 17198 2674 17292
rect 2694 17198 2698 17292
rect 2718 17198 2722 17292
rect 2742 17198 2746 17292
rect 2766 17198 2770 17292
rect 2790 17198 2794 17292
rect 2814 17198 2818 17292
rect 2838 17198 2842 17292
rect 2862 17198 2866 17292
rect 2886 17198 2890 17292
rect 2910 17198 2914 17292
rect 2934 17198 2938 17292
rect 2958 17198 2962 17292
rect 2982 17198 2986 17292
rect 3006 17198 3010 17292
rect 3030 17198 3034 17292
rect 3054 17198 3058 17292
rect 3078 17198 3082 17292
rect 3102 17198 3106 17292
rect 3126 17198 3130 17292
rect 3150 17198 3154 17292
rect 3174 17198 3178 17292
rect 3198 17198 3202 17292
rect 3222 17198 3226 17292
rect 3246 17198 3250 17292
rect 3270 17198 3274 17292
rect 3294 17198 3298 17292
rect 3318 17198 3322 17292
rect 3342 17198 3346 17292
rect 3366 17198 3370 17292
rect 3390 17198 3394 17292
rect 3414 17198 3418 17292
rect 3438 17198 3442 17292
rect 3462 17198 3466 17292
rect 3486 17198 3490 17292
rect 3510 17198 3514 17292
rect 3534 17198 3538 17292
rect 3558 17198 3562 17292
rect 3582 17198 3586 17292
rect 3606 17198 3610 17292
rect 3630 17198 3634 17292
rect 3654 17198 3658 17292
rect 3678 17198 3682 17292
rect 3702 17198 3706 17292
rect 3726 17198 3730 17292
rect 3750 17198 3754 17292
rect 3774 17198 3778 17292
rect 3798 17198 3802 17292
rect 3811 17285 3816 17292
rect 3829 17291 3843 17292
rect 3821 17271 3826 17285
rect 3811 17213 3816 17223
rect 3822 17213 3826 17271
rect 3821 17199 3826 17213
rect 3835 17209 3843 17213
rect 3829 17199 3835 17209
rect 3811 17198 3843 17199
rect -2393 17196 3843 17198
rect -2371 17174 -2366 17196
rect -2348 17174 -2343 17196
rect -2325 17174 -2320 17196
rect -2072 17194 -2036 17195
rect -2072 17188 -2054 17194
rect -2309 17180 -2301 17188
rect -2317 17174 -2309 17180
rect -2092 17179 -2062 17184
rect -2000 17175 -1992 17196
rect -1938 17195 -1906 17196
rect -1920 17194 -1906 17195
rect -1806 17188 -1680 17194
rect -1854 17179 -1806 17184
rect -1655 17180 -1647 17188
rect -1982 17175 -1966 17176
rect -2000 17174 -1966 17175
rect -1846 17174 -1806 17177
rect -1663 17174 -1655 17180
rect -1642 17174 -1637 17196
rect -1619 17174 -1614 17196
rect -1530 17174 -1526 17196
rect -1506 17195 -1502 17196
rect -2393 17172 -1509 17174
rect -2371 17150 -2366 17172
rect -2348 17150 -2343 17172
rect -2325 17150 -2320 17172
rect -2000 17170 -1966 17172
rect -2309 17152 -2301 17160
rect -2062 17159 -2054 17166
rect -2092 17152 -2084 17159
rect -2062 17152 -2026 17154
rect -2317 17150 -2309 17152
rect -2062 17150 -2012 17152
rect -2000 17150 -1992 17170
rect -1982 17169 -1966 17170
rect -1846 17168 -1806 17172
rect -1846 17161 -1798 17166
rect -1806 17159 -1798 17161
rect -1854 17157 -1846 17159
rect -1854 17152 -1806 17157
rect -1655 17152 -1647 17160
rect -1864 17150 -1796 17151
rect -1663 17150 -1655 17152
rect -1642 17150 -1637 17172
rect -1619 17150 -1614 17172
rect -1530 17150 -1526 17172
rect -1523 17171 -1509 17172
rect -1506 17150 -1499 17195
rect -1482 17150 -1478 17196
rect -1458 17150 -1454 17196
rect -1434 17150 -1430 17196
rect -1410 17150 -1406 17196
rect -1386 17150 -1382 17196
rect -1362 17150 -1358 17196
rect -1338 17150 -1334 17196
rect -1314 17150 -1310 17196
rect -1290 17150 -1286 17196
rect -1266 17150 -1262 17196
rect -1242 17150 -1238 17196
rect -1218 17150 -1214 17196
rect -1194 17150 -1190 17196
rect -1170 17150 -1166 17196
rect -1146 17150 -1142 17196
rect -1122 17150 -1118 17196
rect -1098 17150 -1094 17196
rect -1074 17150 -1070 17196
rect -1050 17150 -1046 17196
rect -1026 17150 -1022 17196
rect -1002 17150 -998 17196
rect -978 17150 -974 17196
rect -954 17150 -950 17196
rect -930 17150 -926 17196
rect -906 17150 -902 17196
rect -882 17150 -878 17196
rect -858 17150 -854 17196
rect -834 17150 -830 17196
rect -810 17150 -806 17196
rect -786 17150 -782 17196
rect -762 17150 -758 17196
rect -738 17150 -734 17196
rect -714 17150 -710 17196
rect -690 17150 -686 17196
rect -666 17150 -662 17196
rect -642 17150 -638 17196
rect -618 17150 -614 17196
rect -594 17150 -590 17196
rect -570 17150 -566 17196
rect -546 17150 -542 17196
rect -522 17150 -518 17196
rect -498 17150 -494 17196
rect -474 17150 -470 17196
rect -450 17150 -446 17196
rect -426 17150 -422 17196
rect -402 17150 -398 17196
rect -378 17150 -374 17196
rect -354 17150 -350 17196
rect -330 17150 -326 17196
rect -306 17150 -302 17196
rect -282 17150 -278 17196
rect -258 17150 -254 17196
rect -234 17150 -230 17196
rect -210 17171 -206 17196
rect -2393 17148 -213 17150
rect -2371 17102 -2366 17148
rect -2348 17102 -2343 17148
rect -2325 17102 -2320 17148
rect -2317 17144 -2309 17148
rect -2062 17144 -2054 17148
rect -2154 17140 -2138 17142
rect -2057 17140 -2054 17144
rect -2292 17134 -2054 17140
rect -2052 17134 -2044 17144
rect -2092 17118 -2062 17120
rect -2094 17114 -2062 17118
rect -2000 17102 -1992 17148
rect -1846 17141 -1806 17148
rect -1663 17144 -1655 17148
rect -1846 17134 -1680 17140
rect -1854 17118 -1806 17120
rect -1854 17114 -1680 17118
rect -1642 17102 -1637 17148
rect -1619 17102 -1614 17148
rect -1530 17102 -1526 17148
rect -1523 17147 -1509 17148
rect -1506 17147 -1499 17148
rect -1506 17102 -1502 17147
rect -1482 17102 -1478 17148
rect -1458 17102 -1454 17148
rect -1434 17102 -1430 17148
rect -1410 17102 -1406 17148
rect -1386 17102 -1382 17148
rect -1362 17102 -1358 17148
rect -1338 17102 -1334 17148
rect -1314 17102 -1310 17148
rect -1290 17102 -1286 17148
rect -1266 17102 -1262 17148
rect -1242 17102 -1238 17148
rect -1218 17102 -1214 17148
rect -1194 17102 -1190 17148
rect -1170 17102 -1166 17148
rect -1146 17102 -1142 17148
rect -1122 17102 -1118 17148
rect -1098 17102 -1094 17148
rect -1074 17102 -1070 17148
rect -1050 17102 -1046 17148
rect -1026 17102 -1022 17148
rect -1002 17102 -998 17148
rect -978 17102 -974 17148
rect -954 17102 -950 17148
rect -930 17102 -926 17148
rect -906 17102 -902 17148
rect -882 17102 -878 17148
rect -858 17102 -854 17148
rect -834 17102 -830 17148
rect -810 17102 -806 17148
rect -786 17102 -782 17148
rect -762 17102 -758 17148
rect -738 17102 -734 17148
rect -714 17102 -710 17148
rect -690 17102 -686 17148
rect -666 17102 -662 17148
rect -642 17102 -638 17148
rect -618 17102 -614 17148
rect -594 17102 -590 17148
rect -570 17102 -566 17148
rect -546 17102 -542 17148
rect -522 17102 -518 17148
rect -498 17102 -494 17148
rect -474 17102 -470 17148
rect -450 17102 -446 17148
rect -426 17102 -422 17148
rect -402 17102 -398 17148
rect -378 17102 -374 17148
rect -354 17102 -350 17148
rect -330 17102 -326 17148
rect -306 17102 -302 17148
rect -282 17102 -278 17148
rect -258 17102 -254 17148
rect -234 17102 -230 17148
rect -227 17147 -213 17148
rect -210 17123 -203 17171
rect -210 17102 -206 17123
rect -186 17102 -182 17196
rect -162 17102 -158 17196
rect -138 17102 -134 17196
rect -114 17102 -110 17196
rect -90 17102 -86 17196
rect -66 17102 -62 17196
rect -42 17102 -38 17196
rect -18 17102 -14 17196
rect 6 17102 10 17196
rect 30 17102 34 17196
rect 54 17102 58 17196
rect 78 17102 82 17196
rect 102 17102 106 17196
rect 126 17102 130 17196
rect 150 17102 154 17196
rect 174 17102 178 17196
rect 198 17102 202 17196
rect 222 17102 226 17196
rect 246 17102 250 17196
rect 270 17102 274 17196
rect 294 17102 298 17196
rect 318 17102 322 17196
rect 342 17102 346 17196
rect 366 17102 370 17196
rect 390 17102 394 17196
rect 414 17102 418 17196
rect 438 17102 442 17196
rect 462 17102 466 17196
rect 486 17102 490 17196
rect 510 17102 514 17196
rect 534 17102 538 17196
rect 558 17102 562 17196
rect 582 17102 586 17196
rect 606 17102 610 17196
rect 630 17102 634 17196
rect 654 17102 658 17196
rect 678 17102 682 17196
rect 702 17102 706 17196
rect 726 17102 730 17196
rect 750 17102 754 17196
rect 774 17102 778 17196
rect 798 17102 802 17196
rect 822 17102 826 17196
rect 846 17102 850 17196
rect 870 17102 874 17196
rect 894 17102 898 17196
rect 918 17102 922 17196
rect 942 17102 946 17196
rect 966 17102 970 17196
rect 990 17102 994 17196
rect 1014 17102 1018 17196
rect 1038 17102 1042 17196
rect 1062 17102 1066 17196
rect 1086 17102 1090 17196
rect 1110 17102 1114 17196
rect 1134 17102 1138 17196
rect 1158 17102 1162 17196
rect 1182 17102 1186 17196
rect 1206 17102 1210 17196
rect 1230 17102 1234 17196
rect 1254 17102 1258 17196
rect 1278 17102 1282 17196
rect 1302 17102 1306 17196
rect 1326 17102 1330 17196
rect 1350 17102 1354 17196
rect 1374 17102 1378 17196
rect 1398 17102 1402 17196
rect 1422 17102 1426 17196
rect 1435 17165 1440 17175
rect 1446 17165 1450 17196
rect 1445 17151 1450 17165
rect 1435 17126 1469 17127
rect 1470 17126 1474 17196
rect 1494 17126 1498 17196
rect 1518 17126 1522 17196
rect 1542 17126 1546 17196
rect 1566 17126 1570 17196
rect 1590 17126 1594 17196
rect 1614 17126 1618 17196
rect 1638 17126 1642 17196
rect 1662 17126 1666 17196
rect 1686 17126 1690 17196
rect 1710 17126 1714 17196
rect 1734 17126 1738 17196
rect 1758 17126 1762 17196
rect 1771 17141 1776 17151
rect 1782 17141 1786 17196
rect 1781 17127 1786 17141
rect 1806 17126 1810 17196
rect 1830 17126 1834 17196
rect 1854 17126 1858 17196
rect 1878 17126 1882 17196
rect 1902 17126 1906 17196
rect 1926 17126 1930 17196
rect 1950 17126 1954 17196
rect 1974 17126 1978 17196
rect 1998 17126 2002 17196
rect 2022 17126 2026 17196
rect 2046 17126 2050 17196
rect 2070 17126 2074 17196
rect 2094 17126 2098 17196
rect 2118 17126 2122 17196
rect 2142 17126 2146 17196
rect 2166 17126 2170 17196
rect 2190 17126 2194 17196
rect 2214 17126 2218 17196
rect 2238 17126 2242 17196
rect 2262 17126 2266 17196
rect 2286 17126 2290 17196
rect 2310 17126 2314 17196
rect 2334 17126 2338 17196
rect 2358 17126 2362 17196
rect 2382 17126 2386 17196
rect 2406 17126 2410 17196
rect 2430 17126 2434 17196
rect 2454 17126 2458 17196
rect 2478 17126 2482 17196
rect 2502 17126 2506 17196
rect 2526 17126 2530 17196
rect 2550 17126 2554 17196
rect 2574 17126 2578 17196
rect 2598 17126 2602 17196
rect 2622 17126 2626 17196
rect 2646 17126 2650 17196
rect 2670 17126 2674 17196
rect 2694 17126 2698 17196
rect 2718 17126 2722 17196
rect 2742 17126 2746 17196
rect 2766 17126 2770 17196
rect 2790 17126 2794 17196
rect 2814 17126 2818 17196
rect 2838 17126 2842 17196
rect 2862 17126 2866 17196
rect 2886 17126 2890 17196
rect 2910 17126 2914 17196
rect 2934 17126 2938 17196
rect 2958 17126 2962 17196
rect 2982 17126 2986 17196
rect 3006 17126 3010 17196
rect 3030 17126 3034 17196
rect 3054 17126 3058 17196
rect 3078 17126 3082 17196
rect 3102 17126 3106 17196
rect 3126 17126 3130 17196
rect 3150 17126 3154 17196
rect 3174 17126 3178 17196
rect 3198 17126 3202 17196
rect 3222 17126 3226 17196
rect 3246 17126 3250 17196
rect 3270 17126 3274 17196
rect 3294 17126 3298 17196
rect 3318 17126 3322 17196
rect 3342 17126 3346 17196
rect 3366 17126 3370 17196
rect 3390 17126 3394 17196
rect 3414 17126 3418 17196
rect 3438 17126 3442 17196
rect 3462 17126 3466 17196
rect 3486 17126 3490 17196
rect 3510 17126 3514 17196
rect 3534 17126 3538 17196
rect 3558 17126 3562 17196
rect 3582 17126 3586 17196
rect 3606 17126 3610 17196
rect 3630 17126 3634 17196
rect 3654 17126 3658 17196
rect 3678 17126 3682 17196
rect 3702 17126 3706 17196
rect 3726 17126 3730 17196
rect 3750 17126 3754 17196
rect 3774 17126 3778 17196
rect 3798 17126 3802 17196
rect 3811 17189 3816 17196
rect 3829 17195 3843 17196
rect 3821 17175 3826 17189
rect 3822 17127 3826 17175
rect 3811 17126 3843 17127
rect 1435 17124 3843 17126
rect 1435 17117 1440 17124
rect 1445 17103 1450 17117
rect 1446 17102 1450 17103
rect 1470 17102 1474 17124
rect 1494 17102 1498 17124
rect 1518 17102 1522 17124
rect 1542 17102 1546 17124
rect 1566 17102 1570 17124
rect 1590 17102 1594 17124
rect 1614 17102 1618 17124
rect 1638 17102 1642 17124
rect 1662 17102 1666 17124
rect 1686 17102 1690 17124
rect 1710 17102 1714 17124
rect 1734 17102 1738 17124
rect 1758 17102 1762 17124
rect 1771 17102 1805 17103
rect -2393 17100 1805 17102
rect -2371 17078 -2366 17100
rect -2348 17078 -2343 17100
rect -2325 17078 -2320 17100
rect -2072 17098 -2036 17099
rect -2072 17092 -2054 17098
rect -2309 17084 -2301 17092
rect -2317 17078 -2309 17084
rect -2092 17083 -2062 17088
rect -2000 17079 -1992 17100
rect -1938 17099 -1906 17100
rect -1920 17098 -1906 17099
rect -1806 17092 -1680 17098
rect -1854 17083 -1806 17088
rect -1655 17084 -1647 17092
rect -1982 17079 -1966 17080
rect -2000 17078 -1966 17079
rect -1846 17078 -1806 17081
rect -1663 17078 -1655 17084
rect -1642 17078 -1637 17100
rect -1619 17078 -1614 17100
rect -1530 17078 -1526 17100
rect -1506 17078 -1502 17100
rect -1482 17078 -1478 17100
rect -1458 17078 -1454 17100
rect -1434 17078 -1430 17100
rect -1410 17078 -1406 17100
rect -1386 17078 -1382 17100
rect -1362 17078 -1358 17100
rect -1338 17078 -1334 17100
rect -1314 17078 -1310 17100
rect -1290 17078 -1286 17100
rect -1266 17078 -1262 17100
rect -1242 17078 -1238 17100
rect -1218 17078 -1214 17100
rect -1194 17078 -1190 17100
rect -1170 17078 -1166 17100
rect -1146 17078 -1142 17100
rect -1122 17078 -1118 17100
rect -1098 17078 -1094 17100
rect -1074 17078 -1070 17100
rect -1050 17078 -1046 17100
rect -1026 17078 -1022 17100
rect -1002 17078 -998 17100
rect -978 17078 -974 17100
rect -954 17078 -950 17100
rect -930 17078 -926 17100
rect -906 17078 -902 17100
rect -882 17078 -878 17100
rect -858 17078 -854 17100
rect -834 17078 -830 17100
rect -810 17078 -806 17100
rect -786 17078 -782 17100
rect -762 17078 -758 17100
rect -738 17078 -734 17100
rect -714 17078 -710 17100
rect -690 17078 -686 17100
rect -666 17078 -662 17100
rect -642 17078 -638 17100
rect -618 17078 -614 17100
rect -594 17078 -590 17100
rect -570 17078 -566 17100
rect -546 17078 -542 17100
rect -522 17078 -518 17100
rect -498 17078 -494 17100
rect -474 17078 -470 17100
rect -450 17078 -446 17100
rect -426 17078 -422 17100
rect -402 17078 -398 17100
rect -378 17078 -374 17100
rect -354 17078 -350 17100
rect -330 17078 -326 17100
rect -306 17078 -302 17100
rect -282 17078 -278 17100
rect -258 17078 -254 17100
rect -234 17078 -230 17100
rect -210 17078 -206 17100
rect -186 17078 -182 17100
rect -162 17078 -158 17100
rect -138 17078 -134 17100
rect -114 17078 -110 17100
rect -90 17078 -86 17100
rect -66 17078 -62 17100
rect -42 17078 -38 17100
rect -18 17078 -14 17100
rect 6 17078 10 17100
rect 30 17078 34 17100
rect 54 17078 58 17100
rect 78 17078 82 17100
rect 102 17078 106 17100
rect 126 17078 130 17100
rect 150 17078 154 17100
rect 174 17078 178 17100
rect 198 17078 202 17100
rect 222 17078 226 17100
rect 246 17078 250 17100
rect 270 17078 274 17100
rect 294 17078 298 17100
rect 318 17078 322 17100
rect 342 17078 346 17100
rect 366 17078 370 17100
rect 390 17078 394 17100
rect 414 17078 418 17100
rect 438 17078 442 17100
rect 462 17078 466 17100
rect 486 17078 490 17100
rect 510 17078 514 17100
rect 534 17078 538 17100
rect 558 17078 562 17100
rect 582 17078 586 17100
rect 606 17078 610 17100
rect 630 17078 634 17100
rect 654 17078 658 17100
rect 678 17078 682 17100
rect 702 17078 706 17100
rect 726 17078 730 17100
rect 750 17078 754 17100
rect 774 17078 778 17100
rect 798 17078 802 17100
rect 822 17078 826 17100
rect 846 17078 850 17100
rect 870 17078 874 17100
rect 894 17078 898 17100
rect 918 17078 922 17100
rect 942 17078 946 17100
rect 966 17078 970 17100
rect 990 17078 994 17100
rect 1014 17078 1018 17100
rect 1038 17078 1042 17100
rect 1062 17078 1066 17100
rect 1086 17078 1090 17100
rect 1110 17078 1114 17100
rect 1134 17078 1138 17100
rect 1158 17078 1162 17100
rect 1182 17078 1186 17100
rect 1206 17078 1210 17100
rect 1230 17078 1234 17100
rect 1254 17078 1258 17100
rect 1278 17078 1282 17100
rect 1302 17078 1306 17100
rect 1326 17078 1330 17100
rect 1350 17078 1354 17100
rect 1374 17078 1378 17100
rect 1398 17078 1402 17100
rect 1422 17078 1426 17100
rect 1446 17078 1450 17100
rect 1470 17099 1474 17100
rect -2393 17076 1467 17078
rect -2371 17054 -2366 17076
rect -2348 17054 -2343 17076
rect -2325 17054 -2320 17076
rect -2000 17074 -1966 17076
rect -2309 17056 -2301 17064
rect -2062 17063 -2054 17070
rect -2092 17056 -2084 17063
rect -2062 17056 -2026 17058
rect -2317 17054 -2309 17056
rect -2062 17054 -2012 17056
rect -2000 17054 -1992 17074
rect -1982 17073 -1966 17074
rect -1846 17072 -1806 17076
rect -1846 17065 -1798 17070
rect -1806 17063 -1798 17065
rect -1854 17061 -1846 17063
rect -1854 17056 -1806 17061
rect -1655 17056 -1647 17064
rect -1864 17054 -1796 17055
rect -1663 17054 -1655 17056
rect -1642 17054 -1637 17076
rect -1619 17054 -1614 17076
rect -1530 17054 -1526 17076
rect -1506 17054 -1502 17076
rect -1482 17054 -1478 17076
rect -1458 17054 -1454 17076
rect -1434 17054 -1430 17076
rect -1410 17054 -1406 17076
rect -1386 17054 -1382 17076
rect -1362 17054 -1358 17076
rect -1338 17054 -1334 17076
rect -1314 17054 -1310 17076
rect -1290 17054 -1286 17076
rect -1266 17054 -1262 17076
rect -1242 17054 -1238 17076
rect -1218 17054 -1214 17076
rect -1194 17054 -1190 17076
rect -1170 17054 -1166 17076
rect -1146 17054 -1142 17076
rect -1122 17054 -1118 17076
rect -1098 17054 -1094 17076
rect -1074 17054 -1070 17076
rect -1050 17054 -1046 17076
rect -1026 17054 -1022 17076
rect -1002 17054 -998 17076
rect -978 17054 -974 17076
rect -954 17054 -950 17076
rect -930 17054 -926 17076
rect -906 17054 -902 17076
rect -882 17054 -878 17076
rect -858 17054 -854 17076
rect -834 17055 -830 17076
rect -845 17054 -811 17055
rect -2393 17052 -811 17054
rect -2371 17006 -2366 17052
rect -2348 17006 -2343 17052
rect -2325 17006 -2320 17052
rect -2317 17048 -2309 17052
rect -2062 17048 -2054 17052
rect -2154 17044 -2138 17046
rect -2057 17044 -2054 17048
rect -2292 17038 -2054 17044
rect -2052 17038 -2044 17048
rect -2092 17022 -2062 17024
rect -2094 17018 -2062 17022
rect -2000 17006 -1992 17052
rect -1846 17045 -1806 17052
rect -1663 17048 -1655 17052
rect -1846 17038 -1680 17044
rect -1854 17022 -1806 17024
rect -1854 17018 -1680 17022
rect -1642 17006 -1637 17052
rect -1619 17006 -1614 17052
rect -1530 17006 -1526 17052
rect -1506 17006 -1502 17052
rect -1482 17006 -1478 17052
rect -1458 17006 -1454 17052
rect -1434 17006 -1430 17052
rect -1410 17006 -1406 17052
rect -1386 17006 -1382 17052
rect -1362 17006 -1358 17052
rect -1338 17006 -1334 17052
rect -1314 17006 -1310 17052
rect -1290 17006 -1286 17052
rect -1266 17006 -1262 17052
rect -1242 17006 -1238 17052
rect -1218 17006 -1214 17052
rect -1194 17006 -1190 17052
rect -1170 17006 -1166 17052
rect -1146 17006 -1142 17052
rect -1122 17006 -1118 17052
rect -1098 17006 -1094 17052
rect -1074 17006 -1070 17052
rect -1050 17006 -1046 17052
rect -1026 17006 -1022 17052
rect -1002 17006 -998 17052
rect -978 17006 -974 17052
rect -954 17006 -950 17052
rect -930 17006 -926 17052
rect -906 17006 -902 17052
rect -882 17006 -878 17052
rect -858 17006 -854 17052
rect -845 17045 -840 17052
rect -834 17045 -830 17052
rect -835 17031 -830 17045
rect -834 17006 -830 17031
rect -810 17006 -806 17076
rect -786 17006 -782 17076
rect -762 17006 -758 17076
rect -738 17006 -734 17076
rect -714 17006 -710 17076
rect -690 17006 -686 17076
rect -666 17006 -662 17076
rect -642 17006 -638 17076
rect -618 17006 -614 17076
rect -594 17006 -590 17076
rect -570 17006 -566 17076
rect -546 17006 -542 17076
rect -522 17006 -518 17076
rect -498 17006 -494 17076
rect -474 17006 -470 17076
rect -450 17006 -446 17076
rect -426 17006 -422 17076
rect -402 17006 -398 17076
rect -378 17006 -374 17076
rect -354 17006 -350 17076
rect -330 17006 -326 17076
rect -306 17006 -302 17076
rect -282 17006 -278 17076
rect -258 17006 -254 17076
rect -234 17006 -230 17076
rect -210 17006 -206 17076
rect -186 17006 -182 17076
rect -162 17006 -158 17076
rect -138 17006 -134 17076
rect -114 17006 -110 17076
rect -90 17006 -86 17076
rect -66 17006 -62 17076
rect -42 17006 -38 17076
rect -18 17006 -14 17076
rect 6 17006 10 17076
rect 30 17006 34 17076
rect 54 17006 58 17076
rect 78 17006 82 17076
rect 102 17006 106 17076
rect 126 17006 130 17076
rect 150 17006 154 17076
rect 174 17006 178 17076
rect 198 17006 202 17076
rect 222 17006 226 17076
rect 246 17006 250 17076
rect 270 17006 274 17076
rect 294 17006 298 17076
rect 318 17006 322 17076
rect 342 17006 346 17076
rect 366 17006 370 17076
rect 390 17006 394 17076
rect 414 17006 418 17076
rect 438 17006 442 17076
rect 462 17006 466 17076
rect 486 17006 490 17076
rect 510 17006 514 17076
rect 534 17006 538 17076
rect 558 17006 562 17076
rect 582 17006 586 17076
rect 606 17006 610 17076
rect 630 17006 634 17076
rect 654 17006 658 17076
rect 678 17006 682 17076
rect 702 17006 706 17076
rect 726 17006 730 17076
rect 750 17006 754 17076
rect 774 17006 778 17076
rect 798 17006 802 17076
rect 822 17006 826 17076
rect 846 17006 850 17076
rect 870 17006 874 17076
rect 894 17006 898 17076
rect 918 17006 922 17076
rect 942 17006 946 17076
rect 966 17006 970 17076
rect 990 17006 994 17076
rect 1014 17006 1018 17076
rect 1038 17006 1042 17076
rect 1062 17006 1066 17076
rect 1086 17006 1090 17076
rect 1110 17006 1114 17076
rect 1134 17006 1138 17076
rect 1158 17006 1162 17076
rect 1182 17006 1186 17076
rect 1206 17006 1210 17076
rect 1230 17006 1234 17076
rect 1254 17006 1258 17076
rect 1278 17006 1282 17076
rect 1302 17006 1306 17076
rect 1326 17006 1330 17076
rect 1350 17006 1354 17076
rect 1374 17006 1378 17076
rect 1398 17006 1402 17076
rect 1422 17006 1426 17076
rect 1446 17006 1450 17076
rect 1453 17075 1467 17076
rect 1470 17075 1477 17099
rect 1470 17027 1477 17051
rect 1470 17006 1474 17027
rect 1494 17006 1498 17100
rect 1518 17006 1522 17100
rect 1542 17006 1546 17100
rect 1566 17006 1570 17100
rect 1590 17006 1594 17100
rect 1614 17006 1618 17100
rect 1638 17006 1642 17100
rect 1662 17006 1666 17100
rect 1686 17006 1690 17100
rect 1710 17006 1714 17100
rect 1734 17006 1738 17100
rect 1758 17006 1762 17100
rect 1771 17093 1776 17100
rect 1781 17079 1786 17093
rect 1782 17006 1786 17079
rect 1806 17075 1810 17124
rect 1806 17051 1813 17075
rect -2393 17004 1803 17006
rect -2371 16982 -2366 17004
rect -2348 16982 -2343 17004
rect -2325 16982 -2320 17004
rect -2072 17002 -2036 17003
rect -2072 16996 -2054 17002
rect -2309 16988 -2301 16996
rect -2317 16982 -2309 16988
rect -2092 16987 -2062 16992
rect -2000 16983 -1992 17004
rect -1938 17003 -1906 17004
rect -1920 17002 -1906 17003
rect -1806 16996 -1680 17002
rect -1854 16987 -1806 16992
rect -1655 16988 -1647 16996
rect -1982 16983 -1966 16984
rect -2000 16982 -1966 16983
rect -1846 16982 -1806 16985
rect -1663 16982 -1655 16988
rect -1642 16982 -1637 17004
rect -1619 16982 -1614 17004
rect -1530 16982 -1526 17004
rect -1506 16982 -1502 17004
rect -1482 16982 -1478 17004
rect -1458 16982 -1454 17004
rect -1434 16982 -1430 17004
rect -1410 16982 -1406 17004
rect -1386 16982 -1382 17004
rect -1362 16982 -1358 17004
rect -1338 16982 -1334 17004
rect -1314 16982 -1310 17004
rect -1290 16982 -1286 17004
rect -1266 16982 -1262 17004
rect -1242 16982 -1238 17004
rect -1218 16982 -1214 17004
rect -1194 16982 -1190 17004
rect -1170 16982 -1166 17004
rect -1146 16982 -1142 17004
rect -1122 16982 -1118 17004
rect -1098 16982 -1094 17004
rect -1074 16982 -1070 17004
rect -1050 16982 -1046 17004
rect -1026 16982 -1022 17004
rect -1002 16982 -998 17004
rect -978 16982 -974 17004
rect -954 16982 -950 17004
rect -930 16982 -926 17004
rect -906 16982 -902 17004
rect -882 16982 -878 17004
rect -858 16982 -854 17004
rect -834 16982 -830 17004
rect -810 16982 -806 17004
rect -786 16982 -782 17004
rect -762 16982 -758 17004
rect -738 16982 -734 17004
rect -714 16982 -710 17004
rect -690 16982 -686 17004
rect -666 16982 -662 17004
rect -642 16982 -638 17004
rect -618 16982 -614 17004
rect -594 16982 -590 17004
rect -570 16982 -566 17004
rect -546 16982 -542 17004
rect -522 16982 -518 17004
rect -498 16982 -494 17004
rect -474 16982 -470 17004
rect -450 16982 -446 17004
rect -426 16982 -422 17004
rect -402 16982 -398 17004
rect -378 16982 -374 17004
rect -354 16982 -350 17004
rect -330 16982 -326 17004
rect -306 16982 -302 17004
rect -282 16982 -278 17004
rect -258 16982 -254 17004
rect -234 16982 -230 17004
rect -210 16982 -206 17004
rect -186 16982 -182 17004
rect -162 16982 -158 17004
rect -138 16982 -134 17004
rect -114 16982 -110 17004
rect -90 16982 -86 17004
rect -66 16982 -62 17004
rect -42 16982 -38 17004
rect -18 16982 -14 17004
rect 6 16982 10 17004
rect 30 16982 34 17004
rect 54 16982 58 17004
rect 78 16982 82 17004
rect 102 16982 106 17004
rect 126 16982 130 17004
rect 150 16982 154 17004
rect 174 16982 178 17004
rect 198 16982 202 17004
rect 222 16982 226 17004
rect 246 16982 250 17004
rect 270 16982 274 17004
rect 294 16982 298 17004
rect 318 16982 322 17004
rect 342 16982 346 17004
rect 366 16982 370 17004
rect 390 16982 394 17004
rect 414 16982 418 17004
rect 438 16982 442 17004
rect 462 16982 466 17004
rect 486 16982 490 17004
rect 510 16982 514 17004
rect 534 16982 538 17004
rect 558 16982 562 17004
rect 582 16982 586 17004
rect 606 16982 610 17004
rect 630 16982 634 17004
rect 654 16982 658 17004
rect 678 16982 682 17004
rect 702 16982 706 17004
rect 726 16982 730 17004
rect 750 16982 754 17004
rect 774 16982 778 17004
rect 798 16982 802 17004
rect 822 16982 826 17004
rect 846 16982 850 17004
rect 870 16982 874 17004
rect 894 16982 898 17004
rect 918 16982 922 17004
rect 942 16982 946 17004
rect 966 16982 970 17004
rect 990 16982 994 17004
rect 1014 16982 1018 17004
rect 1038 16982 1042 17004
rect 1062 16982 1066 17004
rect 1086 16982 1090 17004
rect 1110 16982 1114 17004
rect 1134 16982 1138 17004
rect 1158 16982 1162 17004
rect 1182 16982 1186 17004
rect 1206 16982 1210 17004
rect 1230 16982 1234 17004
rect 1254 16982 1258 17004
rect 1278 16982 1282 17004
rect 1302 16982 1306 17004
rect 1326 16982 1330 17004
rect 1350 16982 1354 17004
rect 1374 16982 1378 17004
rect 1398 16982 1402 17004
rect 1422 16982 1426 17004
rect 1446 16982 1450 17004
rect 1470 16982 1474 17004
rect 1494 16982 1498 17004
rect 1518 16982 1522 17004
rect 1542 16982 1546 17004
rect 1566 16982 1570 17004
rect 1590 16982 1594 17004
rect 1614 16982 1618 17004
rect 1638 16982 1642 17004
rect 1662 16982 1666 17004
rect 1686 16982 1690 17004
rect 1710 16982 1714 17004
rect 1734 16982 1738 17004
rect 1758 16982 1762 17004
rect 1782 16982 1786 17004
rect 1789 17003 1803 17004
rect 1806 17003 1813 17027
rect 1806 16982 1810 17003
rect 1830 16982 1834 17124
rect 1854 16982 1858 17124
rect 1878 16982 1882 17124
rect 1902 16982 1906 17124
rect 1926 16982 1930 17124
rect 1950 16982 1954 17124
rect 1974 16982 1978 17124
rect 1998 16982 2002 17124
rect 2022 16982 2026 17124
rect 2046 16982 2050 17124
rect 2070 16982 2074 17124
rect 2094 16982 2098 17124
rect 2118 16982 2122 17124
rect 2142 16982 2146 17124
rect 2166 16982 2170 17124
rect 2190 16982 2194 17124
rect 2214 16982 2218 17124
rect 2238 16982 2242 17124
rect 2262 16982 2266 17124
rect 2286 16982 2290 17124
rect 2310 16982 2314 17124
rect 2334 16982 2338 17124
rect 2358 16982 2362 17124
rect 2382 16982 2386 17124
rect 2406 16982 2410 17124
rect 2430 16982 2434 17124
rect 2454 16982 2458 17124
rect 2478 16982 2482 17124
rect 2502 16982 2506 17124
rect 2526 16982 2530 17124
rect 2550 16982 2554 17124
rect 2574 16982 2578 17124
rect 2598 16982 2602 17124
rect 2622 16982 2626 17124
rect 2646 16982 2650 17124
rect 2670 16982 2674 17124
rect 2694 16982 2698 17124
rect 2718 16982 2722 17124
rect 2742 16982 2746 17124
rect 2766 16982 2770 17124
rect 2790 16982 2794 17124
rect 2814 16982 2818 17124
rect 2838 16982 2842 17124
rect 2862 16982 2866 17124
rect 2886 16982 2890 17124
rect 2910 16982 2914 17124
rect 2934 16983 2938 17124
rect 2923 16982 2957 16983
rect -2393 16980 2957 16982
rect -2371 16958 -2366 16980
rect -2348 16958 -2343 16980
rect -2325 16958 -2320 16980
rect -2000 16978 -1966 16980
rect -2309 16960 -2301 16968
rect -2062 16967 -2054 16974
rect -2092 16960 -2084 16967
rect -2062 16960 -2026 16962
rect -2317 16958 -2309 16960
rect -2062 16958 -2012 16960
rect -2000 16958 -1992 16978
rect -1982 16977 -1966 16978
rect -1846 16976 -1806 16980
rect -1846 16969 -1798 16974
rect -1806 16967 -1798 16969
rect -1854 16965 -1846 16967
rect -1854 16960 -1806 16965
rect -1655 16960 -1647 16968
rect -1864 16958 -1796 16959
rect -1663 16958 -1655 16960
rect -1642 16958 -1637 16980
rect -1619 16958 -1614 16980
rect -1530 16958 -1526 16980
rect -1506 16958 -1502 16980
rect -1482 16958 -1478 16980
rect -1458 16958 -1454 16980
rect -1434 16958 -1430 16980
rect -1410 16958 -1406 16980
rect -1386 16958 -1382 16980
rect -1362 16958 -1358 16980
rect -1338 16958 -1334 16980
rect -1314 16958 -1310 16980
rect -1290 16958 -1286 16980
rect -1266 16958 -1262 16980
rect -1242 16958 -1238 16980
rect -1218 16958 -1214 16980
rect -1194 16958 -1190 16980
rect -1170 16958 -1166 16980
rect -1146 16958 -1142 16980
rect -1122 16958 -1118 16980
rect -1098 16958 -1094 16980
rect -1074 16958 -1070 16980
rect -1050 16958 -1046 16980
rect -1026 16958 -1022 16980
rect -1002 16958 -998 16980
rect -978 16958 -974 16980
rect -954 16958 -950 16980
rect -930 16958 -926 16980
rect -906 16958 -902 16980
rect -882 16958 -878 16980
rect -858 16958 -854 16980
rect -834 16958 -830 16980
rect -810 16979 -806 16980
rect -2393 16956 -813 16958
rect -2371 16910 -2366 16956
rect -2348 16910 -2343 16956
rect -2325 16920 -2320 16956
rect -2317 16952 -2309 16956
rect -2062 16952 -2054 16956
rect -2154 16948 -2138 16950
rect -2057 16948 -2054 16952
rect -2292 16942 -2054 16948
rect -2052 16942 -2044 16952
rect -2092 16926 -2062 16928
rect -2094 16922 -2062 16926
rect -2325 16910 -2317 16920
rect -2095 16912 -2084 16916
rect -2000 16913 -1992 16956
rect -1846 16949 -1806 16956
rect -1663 16952 -1655 16956
rect -1846 16942 -1680 16948
rect -1854 16926 -1806 16928
rect -1854 16922 -1680 16926
rect -2119 16910 -2069 16912
rect -2054 16910 -1892 16913
rect -1671 16910 -1663 16920
rect -1642 16910 -1637 16956
rect -1619 16910 -1614 16956
rect -1530 16910 -1526 16956
rect -1506 16910 -1502 16956
rect -1482 16910 -1478 16956
rect -1458 16910 -1454 16956
rect -1434 16910 -1430 16956
rect -1410 16910 -1406 16956
rect -1386 16910 -1382 16956
rect -1362 16910 -1358 16956
rect -1338 16910 -1334 16956
rect -1314 16910 -1310 16956
rect -1290 16910 -1286 16956
rect -1266 16910 -1262 16956
rect -1242 16910 -1238 16956
rect -1218 16910 -1214 16956
rect -1194 16910 -1190 16956
rect -1170 16910 -1166 16956
rect -1146 16910 -1142 16956
rect -1122 16910 -1118 16956
rect -1098 16910 -1094 16956
rect -1074 16910 -1070 16956
rect -1050 16910 -1046 16956
rect -1026 16910 -1022 16956
rect -1002 16910 -998 16956
rect -978 16910 -974 16956
rect -954 16910 -950 16956
rect -930 16910 -926 16956
rect -906 16910 -902 16956
rect -882 16910 -878 16956
rect -858 16910 -854 16956
rect -834 16910 -830 16956
rect -827 16955 -813 16956
rect -810 16955 -803 16979
rect -810 16910 -806 16955
rect -786 16910 -782 16980
rect -762 16910 -758 16980
rect -738 16910 -734 16980
rect -714 16910 -710 16980
rect -690 16910 -686 16980
rect -666 16910 -662 16980
rect -642 16910 -638 16980
rect -618 16910 -614 16980
rect -594 16910 -590 16980
rect -570 16910 -566 16980
rect -546 16910 -542 16980
rect -522 16910 -518 16980
rect -498 16910 -494 16980
rect -474 16910 -470 16980
rect -450 16910 -446 16980
rect -426 16910 -422 16980
rect -402 16910 -398 16980
rect -378 16910 -374 16980
rect -354 16910 -350 16980
rect -330 16910 -326 16980
rect -306 16910 -302 16980
rect -282 16910 -278 16980
rect -258 16910 -254 16980
rect -234 16910 -230 16980
rect -210 16910 -206 16980
rect -186 16910 -182 16980
rect -162 16910 -158 16980
rect -138 16910 -134 16980
rect -114 16910 -110 16980
rect -90 16910 -86 16980
rect -66 16910 -62 16980
rect -42 16910 -38 16980
rect -18 16910 -14 16980
rect 6 16910 10 16980
rect 30 16910 34 16980
rect 54 16910 58 16980
rect 78 16910 82 16980
rect 102 16910 106 16980
rect 126 16910 130 16980
rect 150 16910 154 16980
rect 174 16910 178 16980
rect 198 16910 202 16980
rect 222 16910 226 16980
rect 246 16910 250 16980
rect 270 16910 274 16980
rect 294 16910 298 16980
rect 318 16910 322 16980
rect 342 16910 346 16980
rect 366 16910 370 16980
rect 390 16910 394 16980
rect 414 16910 418 16980
rect 438 16910 442 16980
rect 462 16910 466 16980
rect 486 16910 490 16980
rect 510 16910 514 16980
rect 534 16910 538 16980
rect 558 16910 562 16980
rect 582 16910 586 16980
rect 606 16910 610 16980
rect 630 16910 634 16980
rect 654 16910 658 16980
rect 678 16910 682 16980
rect 702 16910 706 16980
rect 726 16910 730 16980
rect 750 16910 754 16980
rect 774 16910 778 16980
rect 798 16910 802 16980
rect 822 16910 826 16980
rect 846 16910 850 16980
rect 870 16910 874 16980
rect 894 16910 898 16980
rect 918 16910 922 16980
rect 942 16910 946 16980
rect 966 16910 970 16980
rect 990 16910 994 16980
rect 1014 16910 1018 16980
rect 1038 16910 1042 16980
rect 1062 16910 1066 16980
rect 1086 16910 1090 16980
rect 1110 16910 1114 16980
rect 1134 16910 1138 16980
rect 1158 16910 1162 16980
rect 1182 16910 1186 16980
rect 1206 16910 1210 16980
rect 1230 16910 1234 16980
rect 1254 16910 1258 16980
rect 1278 16910 1282 16980
rect 1302 16910 1306 16980
rect 1326 16910 1330 16980
rect 1350 16910 1354 16980
rect 1374 16910 1378 16980
rect 1398 16910 1402 16980
rect 1422 16910 1426 16980
rect 1446 16910 1450 16980
rect 1470 16910 1474 16980
rect 1494 16910 1498 16980
rect 1518 16910 1522 16980
rect 1542 16910 1546 16980
rect 1566 16910 1570 16980
rect 1590 16910 1594 16980
rect 1614 16910 1618 16980
rect 1638 16910 1642 16980
rect 1662 16910 1666 16980
rect 1686 16910 1690 16980
rect 1710 16910 1714 16980
rect 1734 16910 1738 16980
rect 1758 16910 1762 16980
rect 1782 16910 1786 16980
rect 1806 16910 1810 16980
rect 1830 16910 1834 16980
rect 1854 16910 1858 16980
rect 1878 16910 1882 16980
rect 1902 16910 1906 16980
rect 1915 16949 1920 16959
rect 1926 16949 1930 16980
rect 1925 16935 1930 16949
rect 1926 16910 1930 16935
rect 1950 16910 1954 16980
rect 1974 16910 1978 16980
rect 1998 16910 2002 16980
rect 2022 16910 2026 16980
rect 2046 16910 2050 16980
rect 2070 16910 2074 16980
rect 2094 16910 2098 16980
rect 2118 16910 2122 16980
rect 2142 16910 2146 16980
rect 2166 16910 2170 16980
rect 2190 16910 2194 16980
rect 2214 16910 2218 16980
rect 2238 16910 2242 16980
rect 2262 16910 2266 16980
rect 2286 16910 2290 16980
rect 2310 16910 2314 16980
rect 2334 16910 2338 16980
rect 2358 16910 2362 16980
rect 2382 16910 2386 16980
rect 2406 16910 2410 16980
rect 2430 16910 2434 16980
rect 2454 16910 2458 16980
rect 2478 16910 2482 16980
rect 2502 16910 2506 16980
rect 2526 16910 2530 16980
rect 2550 16910 2554 16980
rect 2574 16910 2578 16980
rect 2598 16910 2602 16980
rect 2622 16910 2626 16980
rect 2646 16910 2650 16980
rect 2670 16910 2674 16980
rect 2694 16910 2698 16980
rect 2718 16910 2722 16980
rect 2742 16910 2746 16980
rect 2766 16910 2770 16980
rect 2790 16910 2794 16980
rect 2814 16910 2818 16980
rect 2838 16910 2842 16980
rect 2862 16910 2866 16980
rect 2886 16910 2890 16980
rect 2910 16910 2914 16980
rect 2923 16973 2928 16980
rect 2934 16973 2938 16980
rect 2933 16959 2938 16973
rect 2934 16910 2938 16959
rect 2958 16910 2962 17124
rect 2982 16910 2986 17124
rect 3006 16910 3010 17124
rect 3030 16910 3034 17124
rect 3054 16910 3058 17124
rect 3078 16910 3082 17124
rect 3102 16910 3106 17124
rect 3126 16910 3130 17124
rect 3150 16910 3154 17124
rect 3174 16910 3178 17124
rect 3198 16910 3202 17124
rect 3222 16910 3226 17124
rect 3246 16910 3250 17124
rect 3270 16910 3274 17124
rect 3294 16910 3298 17124
rect 3307 17069 3312 17079
rect 3318 17069 3322 17124
rect 3317 17055 3322 17069
rect 3307 17045 3312 17055
rect 3317 17031 3322 17045
rect 3318 16910 3322 17031
rect 3342 17003 3346 17124
rect 3342 16955 3349 17003
rect 3342 16910 3346 16955
rect 3366 16910 3370 17124
rect 3390 16910 3394 17124
rect 3414 16910 3418 17124
rect 3438 16910 3442 17124
rect 3462 16910 3466 17124
rect 3486 16910 3490 17124
rect 3510 16910 3514 17124
rect 3534 16910 3538 17124
rect 3558 16910 3562 17124
rect 3582 16910 3586 17124
rect 3606 16910 3610 17124
rect 3630 16910 3634 17124
rect 3654 16910 3658 17124
rect 3678 16910 3682 17124
rect 3702 16910 3706 17124
rect 3726 16910 3730 17124
rect 3750 16910 3754 17124
rect 3774 16910 3778 17124
rect 3787 17045 3792 17055
rect 3798 17045 3802 17124
rect 3811 17117 3816 17124
rect 3822 17117 3826 17124
rect 3829 17123 3843 17124
rect 3821 17103 3826 17117
rect 3835 17113 3843 17117
rect 3829 17103 3835 17113
rect 3797 17031 3802 17045
rect 3787 16997 3792 17007
rect 3797 16983 3802 16997
rect 3798 16910 3802 16983
rect 3811 16910 3819 16911
rect -2393 16908 3819 16910
rect -2371 16886 -2366 16908
rect -2348 16886 -2343 16908
rect -2325 16904 -2317 16908
rect -2325 16888 -2320 16904
rect -2309 16892 -2301 16904
rect -2095 16902 -2084 16908
rect -2054 16907 -1906 16908
rect -2054 16906 -2036 16907
rect -2084 16900 -2079 16902
rect -2317 16888 -2309 16892
rect -2092 16891 -2079 16898
rect -2000 16894 -1992 16907
rect -1920 16906 -1906 16907
rect -1671 16904 -1663 16908
rect -1846 16900 -1806 16902
rect -1854 16894 -1806 16898
rect -2054 16891 -1982 16894
rect -1966 16891 -1806 16894
rect -1655 16892 -1647 16904
rect -2003 16888 -1992 16891
rect -1904 16889 -1902 16891
rect -1854 16889 -1846 16891
rect -2325 16886 -2317 16888
rect -2033 16886 -1992 16888
rect -1854 16887 -1806 16889
rect -1663 16888 -1655 16892
rect -1864 16886 -1796 16887
rect -1671 16886 -1663 16888
rect -1642 16886 -1637 16908
rect -1619 16886 -1614 16908
rect -1530 16886 -1526 16908
rect -1506 16886 -1502 16908
rect -1482 16886 -1478 16908
rect -1458 16886 -1454 16908
rect -1434 16886 -1430 16908
rect -1410 16886 -1406 16908
rect -1386 16886 -1382 16908
rect -1362 16886 -1358 16908
rect -1338 16886 -1334 16908
rect -1314 16886 -1310 16908
rect -1290 16886 -1286 16908
rect -1266 16886 -1262 16908
rect -1242 16886 -1238 16908
rect -1218 16886 -1214 16908
rect -1194 16886 -1190 16908
rect -1170 16886 -1166 16908
rect -1146 16886 -1142 16908
rect -1122 16886 -1118 16908
rect -1098 16886 -1094 16908
rect -1074 16886 -1070 16908
rect -1050 16886 -1046 16908
rect -1026 16886 -1022 16908
rect -1002 16886 -998 16908
rect -978 16886 -974 16908
rect -954 16886 -950 16908
rect -930 16886 -926 16908
rect -906 16886 -902 16908
rect -882 16886 -878 16908
rect -858 16886 -854 16908
rect -834 16886 -830 16908
rect -810 16886 -806 16908
rect -786 16886 -782 16908
rect -762 16886 -758 16908
rect -738 16886 -734 16908
rect -714 16886 -710 16908
rect -690 16886 -686 16908
rect -666 16886 -662 16908
rect -642 16886 -638 16908
rect -618 16886 -614 16908
rect -594 16886 -590 16908
rect -570 16886 -566 16908
rect -546 16886 -542 16908
rect -522 16886 -518 16908
rect -498 16886 -494 16908
rect -474 16886 -470 16908
rect -450 16886 -446 16908
rect -426 16886 -422 16908
rect -402 16886 -398 16908
rect -378 16886 -374 16908
rect -354 16886 -350 16908
rect -330 16886 -326 16908
rect -306 16886 -302 16908
rect -282 16886 -278 16908
rect -258 16886 -254 16908
rect -234 16886 -230 16908
rect -210 16886 -206 16908
rect -186 16886 -182 16908
rect -162 16886 -158 16908
rect -138 16886 -134 16908
rect -114 16886 -110 16908
rect -90 16886 -86 16908
rect -66 16886 -62 16908
rect -42 16886 -38 16908
rect -18 16886 -14 16908
rect 6 16886 10 16908
rect 30 16886 34 16908
rect 54 16886 58 16908
rect 78 16886 82 16908
rect 102 16886 106 16908
rect 126 16886 130 16908
rect 150 16886 154 16908
rect 174 16886 178 16908
rect 198 16886 202 16908
rect 222 16886 226 16908
rect 246 16886 250 16908
rect 270 16886 274 16908
rect 294 16886 298 16908
rect 318 16886 322 16908
rect 342 16886 346 16908
rect 366 16886 370 16908
rect 390 16886 394 16908
rect 414 16886 418 16908
rect 438 16886 442 16908
rect 462 16886 466 16908
rect 486 16886 490 16908
rect 510 16886 514 16908
rect 534 16886 538 16908
rect 558 16886 562 16908
rect 582 16886 586 16908
rect 606 16886 610 16908
rect 630 16886 634 16908
rect 654 16886 658 16908
rect 678 16886 682 16908
rect 702 16886 706 16908
rect 726 16886 730 16908
rect 750 16886 754 16908
rect 774 16886 778 16908
rect 798 16886 802 16908
rect 822 16886 826 16908
rect 846 16886 850 16908
rect 870 16886 874 16908
rect 894 16886 898 16908
rect 918 16886 922 16908
rect 942 16886 946 16908
rect 966 16886 970 16908
rect 990 16886 994 16908
rect 1014 16886 1018 16908
rect 1038 16886 1042 16908
rect 1062 16886 1066 16908
rect 1086 16886 1090 16908
rect 1110 16886 1114 16908
rect 1134 16886 1138 16908
rect 1158 16886 1162 16908
rect 1182 16886 1186 16908
rect 1206 16886 1210 16908
rect 1230 16886 1234 16908
rect 1254 16886 1258 16908
rect 1278 16886 1282 16908
rect 1302 16886 1306 16908
rect 1326 16886 1330 16908
rect 1350 16886 1354 16908
rect 1374 16886 1378 16908
rect 1398 16886 1402 16908
rect 1422 16886 1426 16908
rect 1446 16886 1450 16908
rect 1470 16886 1474 16908
rect 1494 16886 1498 16908
rect 1518 16886 1522 16908
rect 1542 16886 1546 16908
rect 1566 16886 1570 16908
rect 1590 16886 1594 16908
rect 1614 16886 1618 16908
rect 1638 16886 1642 16908
rect 1662 16886 1666 16908
rect 1686 16886 1690 16908
rect 1710 16886 1714 16908
rect 1734 16886 1738 16908
rect 1758 16886 1762 16908
rect 1782 16886 1786 16908
rect 1806 16886 1810 16908
rect 1830 16886 1834 16908
rect 1854 16886 1858 16908
rect 1878 16886 1882 16908
rect 1902 16886 1906 16908
rect 1926 16886 1930 16908
rect 1950 16886 1954 16908
rect 1974 16886 1978 16908
rect 1998 16886 2002 16908
rect 2022 16886 2026 16908
rect 2046 16886 2050 16908
rect 2070 16886 2074 16908
rect 2094 16886 2098 16908
rect 2118 16886 2122 16908
rect 2142 16886 2146 16908
rect 2166 16886 2170 16908
rect 2190 16886 2194 16908
rect 2214 16886 2218 16908
rect 2238 16886 2242 16908
rect 2262 16886 2266 16908
rect 2286 16886 2290 16908
rect 2310 16886 2314 16908
rect 2334 16886 2338 16908
rect 2358 16886 2362 16908
rect 2382 16886 2386 16908
rect 2406 16886 2410 16908
rect 2430 16886 2434 16908
rect 2454 16886 2458 16908
rect 2478 16886 2482 16908
rect 2502 16886 2506 16908
rect 2526 16886 2530 16908
rect 2550 16886 2554 16908
rect 2574 16886 2578 16908
rect 2598 16886 2602 16908
rect 2622 16887 2626 16908
rect 2611 16886 2645 16887
rect -2393 16884 2645 16886
rect -2371 16862 -2366 16884
rect -2348 16862 -2343 16884
rect -2325 16876 -2317 16884
rect -2079 16881 -2018 16884
rect -2003 16883 -1966 16884
rect -2000 16882 -1982 16883
rect -2000 16881 -1992 16882
rect -2084 16877 -2009 16881
rect -2028 16876 -2009 16877
rect -2000 16877 -1854 16881
rect -1846 16877 -1798 16884
rect -2325 16862 -2320 16876
rect -2309 16864 -2301 16876
rect -2028 16874 -2018 16876
rect -2092 16864 -2084 16871
rect -2023 16867 -2014 16874
rect -2000 16867 -1992 16877
rect -1671 16876 -1663 16884
rect -1846 16873 -1806 16875
rect -1854 16867 -1806 16871
rect -2054 16864 -1806 16867
rect -1655 16864 -1647 16876
rect -2317 16862 -2309 16864
rect -2054 16862 -2024 16864
rect -2000 16862 -1992 16864
rect -1663 16862 -1655 16864
rect -1642 16862 -1637 16884
rect -1619 16862 -1614 16884
rect -1530 16862 -1526 16884
rect -1506 16862 -1502 16884
rect -1482 16862 -1478 16884
rect -1458 16862 -1454 16884
rect -1434 16862 -1430 16884
rect -1410 16862 -1406 16884
rect -1386 16862 -1382 16884
rect -1362 16862 -1358 16884
rect -1338 16862 -1334 16884
rect -1314 16862 -1310 16884
rect -1290 16862 -1286 16884
rect -1266 16862 -1262 16884
rect -1242 16862 -1238 16884
rect -1218 16862 -1214 16884
rect -1194 16862 -1190 16884
rect -1170 16862 -1166 16884
rect -1146 16862 -1142 16884
rect -1122 16862 -1118 16884
rect -1098 16862 -1094 16884
rect -1074 16862 -1070 16884
rect -1050 16862 -1046 16884
rect -1026 16862 -1022 16884
rect -1002 16862 -998 16884
rect -978 16862 -974 16884
rect -954 16862 -950 16884
rect -930 16862 -926 16884
rect -906 16862 -902 16884
rect -882 16862 -878 16884
rect -858 16862 -854 16884
rect -834 16862 -830 16884
rect -810 16862 -806 16884
rect -786 16862 -782 16884
rect -762 16862 -758 16884
rect -738 16862 -734 16884
rect -714 16862 -710 16884
rect -690 16862 -686 16884
rect -666 16862 -662 16884
rect -642 16862 -638 16884
rect -618 16862 -614 16884
rect -594 16862 -590 16884
rect -570 16862 -566 16884
rect -546 16862 -542 16884
rect -522 16862 -518 16884
rect -498 16862 -494 16884
rect -474 16862 -470 16884
rect -450 16862 -446 16884
rect -426 16862 -422 16884
rect -402 16862 -398 16884
rect -378 16862 -374 16884
rect -354 16862 -350 16884
rect -330 16862 -326 16884
rect -306 16862 -302 16884
rect -282 16862 -278 16884
rect -258 16862 -254 16884
rect -234 16862 -230 16884
rect -210 16862 -206 16884
rect -186 16862 -182 16884
rect -162 16862 -158 16884
rect -138 16862 -134 16884
rect -114 16862 -110 16884
rect -90 16862 -86 16884
rect -66 16862 -62 16884
rect -42 16862 -38 16884
rect -18 16862 -14 16884
rect 6 16862 10 16884
rect 30 16862 34 16884
rect 54 16862 58 16884
rect 78 16862 82 16884
rect 102 16862 106 16884
rect 126 16862 130 16884
rect 150 16862 154 16884
rect 174 16862 178 16884
rect 198 16862 202 16884
rect 222 16862 226 16884
rect 246 16862 250 16884
rect 270 16862 274 16884
rect 294 16862 298 16884
rect 318 16862 322 16884
rect 342 16862 346 16884
rect 366 16862 370 16884
rect 390 16862 394 16884
rect 414 16862 418 16884
rect 438 16862 442 16884
rect 462 16862 466 16884
rect 486 16862 490 16884
rect 510 16862 514 16884
rect 534 16862 538 16884
rect 558 16862 562 16884
rect 582 16862 586 16884
rect 606 16862 610 16884
rect 630 16862 634 16884
rect 654 16862 658 16884
rect 678 16862 682 16884
rect 702 16862 706 16884
rect 726 16862 730 16884
rect 750 16862 754 16884
rect 774 16862 778 16884
rect 798 16862 802 16884
rect 822 16862 826 16884
rect 846 16862 850 16884
rect 870 16862 874 16884
rect 894 16862 898 16884
rect 918 16862 922 16884
rect 942 16862 946 16884
rect 966 16862 970 16884
rect 990 16862 994 16884
rect 1014 16862 1018 16884
rect 1038 16862 1042 16884
rect 1062 16862 1066 16884
rect 1086 16862 1090 16884
rect 1110 16862 1114 16884
rect 1134 16862 1138 16884
rect 1158 16862 1162 16884
rect 1182 16862 1186 16884
rect 1206 16862 1210 16884
rect 1230 16862 1234 16884
rect 1254 16862 1258 16884
rect 1278 16862 1282 16884
rect 1302 16862 1306 16884
rect 1326 16862 1330 16884
rect 1350 16862 1354 16884
rect 1374 16862 1378 16884
rect 1398 16862 1402 16884
rect 1422 16862 1426 16884
rect 1446 16862 1450 16884
rect 1470 16862 1474 16884
rect 1494 16862 1498 16884
rect 1518 16862 1522 16884
rect 1542 16862 1546 16884
rect 1566 16862 1570 16884
rect 1590 16862 1594 16884
rect 1614 16862 1618 16884
rect 1638 16862 1642 16884
rect 1662 16862 1666 16884
rect 1686 16862 1690 16884
rect 1710 16862 1714 16884
rect 1734 16862 1738 16884
rect 1758 16863 1762 16884
rect 1747 16862 1781 16863
rect -2393 16860 -2064 16862
rect -2060 16860 1781 16862
rect -2371 16814 -2366 16860
rect -2348 16814 -2343 16860
rect -2325 16848 -2317 16860
rect -2060 16857 -2054 16860
rect -2084 16850 -2054 16857
rect -2050 16854 -2044 16856
rect -2325 16828 -2320 16848
rect -2064 16846 -2054 16850
rect -2325 16820 -2317 16828
rect -2101 16823 -2071 16826
rect -2325 16814 -2320 16820
rect -2317 16814 -2309 16820
rect -2000 16818 -1992 16860
rect -1846 16859 -1806 16860
rect -1846 16850 -1798 16857
rect -1671 16848 -1663 16860
rect -1846 16846 -1806 16848
rect -1854 16832 -1680 16836
rect -1846 16823 -1798 16826
rect -2079 16817 -2043 16818
rect -2007 16817 -1991 16818
rect -2079 16816 -2071 16817
rect -2079 16814 -2029 16816
rect -2011 16814 -1991 16817
rect -1846 16815 -1806 16821
rect -1671 16820 -1663 16828
rect -1864 16814 -1796 16815
rect -1663 16814 -1655 16820
rect -1642 16814 -1637 16860
rect -1619 16814 -1614 16860
rect -1530 16814 -1526 16860
rect -1506 16814 -1502 16860
rect -1482 16814 -1478 16860
rect -1458 16814 -1454 16860
rect -1434 16814 -1430 16860
rect -1410 16814 -1406 16860
rect -1386 16814 -1382 16860
rect -1362 16814 -1358 16860
rect -1338 16814 -1334 16860
rect -1314 16814 -1310 16860
rect -1290 16814 -1286 16860
rect -1266 16814 -1262 16860
rect -1242 16814 -1238 16860
rect -1218 16814 -1214 16860
rect -1194 16814 -1190 16860
rect -1170 16814 -1166 16860
rect -1146 16814 -1142 16860
rect -1122 16814 -1118 16860
rect -1098 16814 -1094 16860
rect -1074 16814 -1070 16860
rect -1050 16814 -1046 16860
rect -1026 16814 -1022 16860
rect -1002 16814 -998 16860
rect -978 16814 -974 16860
rect -954 16814 -950 16860
rect -930 16814 -926 16860
rect -906 16814 -902 16860
rect -882 16814 -878 16860
rect -858 16814 -854 16860
rect -834 16814 -830 16860
rect -810 16814 -806 16860
rect -786 16814 -782 16860
rect -762 16814 -758 16860
rect -738 16814 -734 16860
rect -714 16814 -710 16860
rect -690 16814 -686 16860
rect -666 16814 -662 16860
rect -642 16814 -638 16860
rect -618 16814 -614 16860
rect -594 16814 -590 16860
rect -570 16814 -566 16860
rect -546 16814 -542 16860
rect -522 16814 -518 16860
rect -498 16814 -494 16860
rect -474 16814 -470 16860
rect -450 16814 -446 16860
rect -426 16814 -422 16860
rect -402 16814 -398 16860
rect -378 16814 -374 16860
rect -354 16814 -350 16860
rect -330 16814 -326 16860
rect -306 16814 -302 16860
rect -282 16814 -278 16860
rect -258 16814 -254 16860
rect -234 16814 -230 16860
rect -210 16814 -206 16860
rect -186 16814 -182 16860
rect -162 16814 -158 16860
rect -138 16814 -134 16860
rect -114 16814 -110 16860
rect -90 16814 -86 16860
rect -66 16814 -62 16860
rect -42 16814 -38 16860
rect -18 16814 -14 16860
rect 6 16814 10 16860
rect 30 16814 34 16860
rect 54 16814 58 16860
rect 78 16814 82 16860
rect 102 16814 106 16860
rect 126 16814 130 16860
rect 150 16814 154 16860
rect 174 16814 178 16860
rect 198 16814 202 16860
rect 222 16814 226 16860
rect 246 16814 250 16860
rect 270 16814 274 16860
rect 294 16814 298 16860
rect 318 16814 322 16860
rect 342 16814 346 16860
rect 366 16814 370 16860
rect 390 16814 394 16860
rect 414 16814 418 16860
rect 438 16814 442 16860
rect 462 16814 466 16860
rect 486 16814 490 16860
rect 510 16814 514 16860
rect 534 16814 538 16860
rect 558 16814 562 16860
rect 582 16814 586 16860
rect 606 16814 610 16860
rect 630 16814 634 16860
rect 654 16814 658 16860
rect 678 16814 682 16860
rect 702 16814 706 16860
rect 726 16814 730 16860
rect 750 16814 754 16860
rect 774 16814 778 16860
rect 798 16814 802 16860
rect 822 16814 826 16860
rect 846 16814 850 16860
rect 870 16814 874 16860
rect 894 16814 898 16860
rect 918 16814 922 16860
rect 942 16814 946 16860
rect 966 16814 970 16860
rect 990 16814 994 16860
rect 1014 16814 1018 16860
rect 1038 16814 1042 16860
rect 1062 16814 1066 16860
rect 1086 16814 1090 16860
rect 1110 16814 1114 16860
rect 1134 16814 1138 16860
rect 1158 16814 1162 16860
rect 1182 16815 1186 16860
rect 1171 16814 1205 16815
rect -2393 16812 1205 16814
rect -2371 16766 -2366 16812
rect -2348 16766 -2343 16812
rect -2325 16800 -2320 16812
rect -2079 16810 -2071 16812
rect -2072 16808 -2071 16810
rect -2109 16803 -2101 16808
rect -2101 16801 -2079 16803
rect -2069 16801 -2068 16808
rect -2325 16792 -2317 16800
rect -2079 16796 -2071 16801
rect -2325 16772 -2320 16792
rect -2317 16784 -2309 16792
rect -2074 16787 -2071 16796
rect -2069 16792 -2068 16796
rect -2109 16778 -2079 16781
rect -2325 16766 -2317 16772
rect -2000 16766 -1992 16812
rect -1846 16810 -1806 16812
rect -1854 16805 -1806 16809
rect -1854 16803 -1846 16805
rect -1846 16801 -1806 16803
rect -1806 16799 -1798 16801
rect -1846 16796 -1798 16799
rect -1846 16783 -1806 16794
rect -1671 16792 -1663 16800
rect -1663 16784 -1655 16792
rect -1854 16778 -1680 16782
rect -1671 16766 -1663 16772
rect -1642 16766 -1637 16812
rect -1619 16766 -1614 16812
rect -1530 16766 -1526 16812
rect -1506 16766 -1502 16812
rect -1482 16766 -1478 16812
rect -1458 16766 -1454 16812
rect -1434 16766 -1430 16812
rect -1410 16766 -1406 16812
rect -1386 16766 -1382 16812
rect -1362 16766 -1358 16812
rect -1338 16766 -1334 16812
rect -1314 16766 -1310 16812
rect -1290 16766 -1286 16812
rect -1266 16766 -1262 16812
rect -1242 16766 -1238 16812
rect -1218 16766 -1214 16812
rect -1194 16766 -1190 16812
rect -1170 16766 -1166 16812
rect -1146 16766 -1142 16812
rect -1122 16766 -1118 16812
rect -1098 16766 -1094 16812
rect -1074 16766 -1070 16812
rect -1050 16766 -1046 16812
rect -1026 16766 -1022 16812
rect -1002 16766 -998 16812
rect -978 16766 -974 16812
rect -954 16766 -950 16812
rect -930 16766 -926 16812
rect -906 16766 -902 16812
rect -882 16766 -878 16812
rect -858 16766 -854 16812
rect -834 16766 -830 16812
rect -810 16766 -806 16812
rect -786 16766 -782 16812
rect -762 16766 -758 16812
rect -738 16766 -734 16812
rect -714 16766 -710 16812
rect -690 16766 -686 16812
rect -666 16766 -662 16812
rect -642 16766 -638 16812
rect -618 16766 -614 16812
rect -594 16766 -590 16812
rect -570 16766 -566 16812
rect -546 16766 -542 16812
rect -522 16766 -518 16812
rect -498 16766 -494 16812
rect -474 16766 -470 16812
rect -450 16766 -446 16812
rect -426 16766 -422 16812
rect -402 16766 -398 16812
rect -378 16766 -374 16812
rect -354 16766 -350 16812
rect -330 16766 -326 16812
rect -306 16766 -302 16812
rect -282 16766 -278 16812
rect -258 16766 -254 16812
rect -234 16766 -230 16812
rect -210 16766 -206 16812
rect -186 16766 -182 16812
rect -162 16766 -158 16812
rect -138 16766 -134 16812
rect -114 16766 -110 16812
rect -90 16766 -86 16812
rect -66 16766 -62 16812
rect -42 16766 -38 16812
rect -18 16766 -14 16812
rect 6 16766 10 16812
rect 30 16766 34 16812
rect 54 16766 58 16812
rect 78 16766 82 16812
rect 102 16766 106 16812
rect 126 16766 130 16812
rect 150 16766 154 16812
rect 174 16766 178 16812
rect 198 16766 202 16812
rect 222 16766 226 16812
rect 246 16766 250 16812
rect 270 16766 274 16812
rect 294 16766 298 16812
rect 318 16766 322 16812
rect 342 16766 346 16812
rect 366 16766 370 16812
rect 390 16766 394 16812
rect 414 16766 418 16812
rect 438 16766 442 16812
rect 462 16766 466 16812
rect 486 16766 490 16812
rect 510 16766 514 16812
rect 534 16766 538 16812
rect 558 16766 562 16812
rect 582 16766 586 16812
rect 606 16766 610 16812
rect 630 16766 634 16812
rect 654 16766 658 16812
rect 678 16766 682 16812
rect 702 16766 706 16812
rect 726 16766 730 16812
rect 750 16766 754 16812
rect 774 16766 778 16812
rect 798 16766 802 16812
rect 822 16766 826 16812
rect 846 16766 850 16812
rect 870 16766 874 16812
rect 894 16766 898 16812
rect 918 16766 922 16812
rect 942 16766 946 16812
rect 966 16766 970 16812
rect 990 16766 994 16812
rect 1014 16766 1018 16812
rect 1038 16766 1042 16812
rect 1062 16766 1066 16812
rect 1086 16766 1090 16812
rect 1110 16766 1114 16812
rect 1134 16766 1138 16812
rect 1158 16766 1162 16812
rect 1171 16805 1176 16812
rect 1182 16805 1186 16812
rect 1181 16791 1186 16805
rect 1171 16790 1205 16791
rect 1206 16790 1210 16860
rect 1230 16790 1234 16860
rect 1254 16790 1258 16860
rect 1278 16790 1282 16860
rect 1302 16790 1306 16860
rect 1326 16790 1330 16860
rect 1350 16790 1354 16860
rect 1374 16790 1378 16860
rect 1398 16790 1402 16860
rect 1422 16790 1426 16860
rect 1446 16790 1450 16860
rect 1470 16790 1474 16860
rect 1494 16790 1498 16860
rect 1518 16790 1522 16860
rect 1542 16790 1546 16860
rect 1566 16790 1570 16860
rect 1590 16790 1594 16860
rect 1614 16790 1618 16860
rect 1638 16790 1642 16860
rect 1662 16790 1666 16860
rect 1686 16790 1690 16860
rect 1710 16790 1714 16860
rect 1734 16790 1738 16860
rect 1747 16853 1752 16860
rect 1758 16853 1762 16860
rect 1757 16839 1762 16853
rect 1747 16814 1781 16815
rect 1782 16814 1786 16884
rect 1806 16814 1810 16884
rect 1830 16814 1834 16884
rect 1854 16814 1858 16884
rect 1878 16814 1882 16884
rect 1902 16814 1906 16884
rect 1926 16814 1930 16884
rect 1950 16883 1954 16884
rect 1950 16859 1957 16883
rect 1950 16814 1954 16859
rect 1974 16814 1978 16884
rect 1998 16814 2002 16884
rect 2022 16814 2026 16884
rect 2046 16814 2050 16884
rect 2070 16814 2074 16884
rect 2094 16814 2098 16884
rect 2118 16814 2122 16884
rect 2142 16814 2146 16884
rect 2166 16814 2170 16884
rect 2190 16814 2194 16884
rect 2214 16814 2218 16884
rect 2238 16814 2242 16884
rect 2262 16814 2266 16884
rect 2286 16814 2290 16884
rect 2310 16814 2314 16884
rect 2334 16814 2338 16884
rect 2358 16814 2362 16884
rect 2382 16814 2386 16884
rect 2406 16814 2410 16884
rect 2430 16814 2434 16884
rect 2454 16814 2458 16884
rect 2478 16814 2482 16884
rect 2502 16814 2506 16884
rect 2526 16814 2530 16884
rect 2550 16814 2554 16884
rect 2574 16814 2578 16884
rect 2598 16814 2602 16884
rect 2611 16877 2616 16884
rect 2622 16877 2626 16884
rect 2621 16863 2626 16877
rect 2611 16853 2616 16863
rect 2621 16839 2626 16853
rect 2622 16814 2626 16839
rect 2646 16814 2650 16908
rect 2670 16814 2674 16908
rect 2694 16814 2698 16908
rect 2718 16814 2722 16908
rect 2742 16814 2746 16908
rect 2766 16814 2770 16908
rect 2790 16814 2794 16908
rect 2814 16814 2818 16908
rect 2838 16814 2842 16908
rect 2862 16814 2866 16908
rect 2886 16814 2890 16908
rect 2910 16814 2914 16908
rect 2934 16814 2938 16908
rect 2958 16907 2962 16908
rect 2958 16883 2965 16907
rect 2958 16814 2962 16883
rect 2971 16829 2976 16839
rect 2982 16829 2986 16908
rect 2981 16815 2986 16829
rect 3006 16814 3010 16908
rect 3030 16814 3034 16908
rect 3054 16814 3058 16908
rect 3078 16814 3082 16908
rect 3102 16814 3106 16908
rect 3126 16814 3130 16908
rect 3150 16814 3154 16908
rect 3174 16814 3178 16908
rect 3198 16814 3202 16908
rect 3222 16814 3226 16908
rect 3246 16814 3250 16908
rect 3270 16814 3274 16908
rect 3294 16814 3298 16908
rect 3318 16814 3322 16908
rect 3342 16814 3346 16908
rect 3366 16814 3370 16908
rect 3390 16814 3394 16908
rect 3414 16814 3418 16908
rect 3438 16814 3442 16908
rect 3462 16814 3466 16908
rect 3486 16814 3490 16908
rect 3510 16814 3514 16908
rect 3534 16814 3538 16908
rect 3558 16814 3562 16908
rect 3582 16814 3586 16908
rect 3606 16814 3610 16908
rect 3630 16814 3634 16908
rect 3654 16814 3658 16908
rect 3678 16814 3682 16908
rect 3702 16814 3706 16908
rect 3726 16814 3730 16908
rect 3750 16814 3754 16908
rect 3774 16814 3778 16908
rect 3798 16815 3802 16908
rect 3805 16907 3819 16908
rect 3811 16901 3816 16907
rect 3821 16887 3826 16901
rect 3811 16853 3816 16863
rect 3822 16853 3826 16887
rect 3821 16839 3826 16853
rect 3787 16814 3821 16815
rect 1747 16812 3821 16814
rect 1747 16805 1752 16812
rect 1757 16791 1762 16805
rect 1758 16790 1762 16791
rect 1782 16790 1786 16812
rect 1806 16790 1810 16812
rect 1830 16790 1834 16812
rect 1854 16790 1858 16812
rect 1878 16790 1882 16812
rect 1902 16790 1906 16812
rect 1926 16790 1930 16812
rect 1950 16790 1954 16812
rect 1974 16790 1978 16812
rect 1998 16790 2002 16812
rect 2022 16790 2026 16812
rect 2046 16790 2050 16812
rect 2070 16790 2074 16812
rect 2094 16790 2098 16812
rect 2118 16790 2122 16812
rect 2142 16790 2146 16812
rect 2166 16790 2170 16812
rect 2190 16790 2194 16812
rect 2214 16790 2218 16812
rect 2238 16790 2242 16812
rect 2262 16790 2266 16812
rect 2286 16790 2290 16812
rect 2310 16790 2314 16812
rect 2334 16790 2338 16812
rect 2358 16790 2362 16812
rect 2382 16790 2386 16812
rect 2406 16790 2410 16812
rect 2430 16790 2434 16812
rect 2454 16790 2458 16812
rect 2478 16790 2482 16812
rect 2502 16790 2506 16812
rect 2526 16790 2530 16812
rect 2550 16790 2554 16812
rect 2574 16790 2578 16812
rect 2598 16790 2602 16812
rect 2622 16790 2626 16812
rect 2646 16811 2650 16812
rect 1171 16788 2643 16790
rect 1171 16781 1176 16788
rect 1181 16767 1186 16781
rect 1182 16766 1186 16767
rect 1206 16766 1210 16788
rect 1230 16766 1234 16788
rect 1254 16766 1258 16788
rect 1278 16766 1282 16788
rect 1302 16766 1306 16788
rect 1326 16766 1330 16788
rect 1350 16766 1354 16788
rect 1374 16766 1378 16788
rect 1398 16766 1402 16788
rect 1422 16766 1426 16788
rect 1446 16766 1450 16788
rect 1470 16766 1474 16788
rect 1494 16766 1498 16788
rect 1518 16766 1522 16788
rect 1542 16766 1546 16788
rect 1566 16766 1570 16788
rect 1590 16766 1594 16788
rect 1614 16766 1618 16788
rect 1638 16766 1642 16788
rect 1662 16766 1666 16788
rect 1686 16766 1690 16788
rect 1710 16766 1714 16788
rect 1734 16766 1738 16788
rect 1758 16766 1762 16788
rect 1782 16787 1786 16788
rect -2393 16764 1779 16766
rect -2371 16742 -2366 16764
rect -2348 16742 -2343 16764
rect -2325 16756 -2317 16764
rect -2325 16742 -2320 16756
rect -2309 16744 -2301 16756
rect -2092 16747 -2062 16752
rect -2000 16744 -1992 16764
rect -2317 16742 -2309 16744
rect -2000 16742 -1983 16744
rect -1906 16742 -1904 16764
rect -1806 16756 -1680 16762
rect -1671 16756 -1663 16764
rect -1854 16747 -1806 16752
rect -1846 16742 -1806 16745
rect -1655 16744 -1647 16756
rect -1663 16742 -1655 16744
rect -1642 16742 -1637 16764
rect -1619 16742 -1614 16764
rect -1530 16742 -1526 16764
rect -1506 16742 -1502 16764
rect -1482 16742 -1478 16764
rect -1458 16742 -1454 16764
rect -1434 16742 -1430 16764
rect -1410 16742 -1406 16764
rect -1386 16742 -1382 16764
rect -1362 16742 -1358 16764
rect -1338 16742 -1334 16764
rect -1314 16742 -1310 16764
rect -1290 16742 -1286 16764
rect -1266 16742 -1262 16764
rect -1242 16742 -1238 16764
rect -1218 16742 -1214 16764
rect -1194 16742 -1190 16764
rect -1170 16742 -1166 16764
rect -1146 16742 -1142 16764
rect -1122 16742 -1118 16764
rect -1098 16742 -1094 16764
rect -1074 16742 -1070 16764
rect -1050 16742 -1046 16764
rect -1026 16742 -1022 16764
rect -1002 16742 -998 16764
rect -978 16742 -974 16764
rect -954 16742 -950 16764
rect -930 16742 -926 16764
rect -906 16742 -902 16764
rect -882 16742 -878 16764
rect -858 16742 -854 16764
rect -834 16742 -830 16764
rect -810 16742 -806 16764
rect -786 16742 -782 16764
rect -762 16742 -758 16764
rect -738 16742 -734 16764
rect -714 16742 -710 16764
rect -690 16742 -686 16764
rect -666 16742 -662 16764
rect -642 16742 -638 16764
rect -618 16742 -614 16764
rect -594 16742 -590 16764
rect -570 16742 -566 16764
rect -546 16742 -542 16764
rect -522 16742 -518 16764
rect -498 16742 -494 16764
rect -474 16742 -470 16764
rect -450 16742 -446 16764
rect -426 16742 -422 16764
rect -402 16742 -398 16764
rect -378 16742 -374 16764
rect -354 16742 -350 16764
rect -330 16742 -326 16764
rect -306 16742 -302 16764
rect -282 16742 -278 16764
rect -258 16742 -254 16764
rect -234 16742 -230 16764
rect -210 16742 -206 16764
rect -186 16742 -182 16764
rect -162 16742 -158 16764
rect -138 16742 -134 16764
rect -114 16742 -110 16764
rect -90 16742 -86 16764
rect -66 16742 -62 16764
rect -42 16742 -38 16764
rect -18 16742 -14 16764
rect 6 16743 10 16764
rect -5 16742 29 16743
rect -2393 16740 29 16742
rect -2371 16718 -2366 16740
rect -2348 16718 -2343 16740
rect -2325 16728 -2317 16740
rect -2071 16736 -2062 16740
rect -2013 16738 -1983 16740
rect -2000 16737 -1983 16738
rect -2325 16718 -2320 16728
rect -2309 16718 -2301 16728
rect -2100 16727 -2092 16734
rect -2064 16732 -2062 16735
rect -2061 16727 -2059 16732
rect -2071 16722 -2062 16727
rect -2071 16720 -2026 16722
rect -2066 16718 -2012 16720
rect -2000 16718 -1992 16737
rect -1906 16735 -1904 16740
rect -1846 16736 -1806 16740
rect -1846 16729 -1798 16734
rect -1806 16727 -1798 16729
rect -1671 16728 -1663 16740
rect -1854 16725 -1846 16727
rect -1854 16720 -1806 16725
rect -1864 16718 -1796 16719
rect -1655 16718 -1647 16728
rect -1642 16718 -1637 16740
rect -1619 16718 -1614 16740
rect -1530 16718 -1526 16740
rect -1506 16719 -1502 16740
rect -1517 16718 -1483 16719
rect -2393 16716 -1483 16718
rect -2371 16670 -2366 16716
rect -2348 16670 -2343 16716
rect -2325 16712 -2320 16716
rect -2317 16712 -2309 16716
rect -2325 16700 -2317 16712
rect -2066 16711 -2062 16716
rect -2147 16708 -2134 16710
rect -2292 16702 -2071 16708
rect -2325 16670 -2320 16700
rect -2092 16686 -2062 16688
rect -2094 16682 -2062 16686
rect -2000 16670 -1992 16716
rect -1846 16709 -1806 16716
rect -1663 16712 -1655 16716
rect -1846 16702 -1680 16708
rect -1671 16700 -1663 16712
rect -1854 16686 -1806 16688
rect -1854 16682 -1680 16686
rect -1926 16670 -1892 16673
rect -1642 16670 -1637 16716
rect -1619 16670 -1614 16716
rect -1530 16670 -1526 16716
rect -1517 16709 -1512 16716
rect -1506 16709 -1502 16716
rect -1507 16695 -1502 16709
rect -1506 16670 -1502 16695
rect -1482 16670 -1478 16740
rect -1458 16670 -1454 16740
rect -1434 16670 -1430 16740
rect -1410 16670 -1406 16740
rect -1386 16670 -1382 16740
rect -1362 16670 -1358 16740
rect -1338 16670 -1334 16740
rect -1314 16670 -1310 16740
rect -1290 16670 -1286 16740
rect -1266 16670 -1262 16740
rect -1242 16670 -1238 16740
rect -1218 16670 -1214 16740
rect -1194 16670 -1190 16740
rect -1170 16670 -1166 16740
rect -1146 16670 -1142 16740
rect -1122 16670 -1118 16740
rect -1098 16670 -1094 16740
rect -1074 16670 -1070 16740
rect -1050 16670 -1046 16740
rect -1026 16670 -1022 16740
rect -1002 16670 -998 16740
rect -978 16670 -974 16740
rect -954 16670 -950 16740
rect -930 16670 -926 16740
rect -906 16670 -902 16740
rect -882 16670 -878 16740
rect -858 16670 -854 16740
rect -834 16670 -830 16740
rect -810 16670 -806 16740
rect -786 16670 -782 16740
rect -762 16670 -758 16740
rect -738 16670 -734 16740
rect -714 16670 -710 16740
rect -690 16670 -686 16740
rect -666 16670 -662 16740
rect -642 16670 -638 16740
rect -618 16670 -614 16740
rect -594 16670 -590 16740
rect -570 16670 -566 16740
rect -546 16670 -542 16740
rect -522 16670 -518 16740
rect -498 16670 -494 16740
rect -474 16670 -470 16740
rect -450 16670 -446 16740
rect -426 16670 -422 16740
rect -402 16670 -398 16740
rect -378 16670 -374 16740
rect -354 16670 -350 16740
rect -330 16670 -326 16740
rect -306 16670 -302 16740
rect -282 16670 -278 16740
rect -258 16670 -254 16740
rect -234 16670 -230 16740
rect -210 16670 -206 16740
rect -186 16670 -182 16740
rect -162 16670 -158 16740
rect -138 16670 -134 16740
rect -114 16670 -110 16740
rect -90 16670 -86 16740
rect -66 16670 -62 16740
rect -42 16670 -38 16740
rect -18 16670 -14 16740
rect -5 16733 0 16740
rect 6 16733 10 16740
rect 5 16719 10 16733
rect -5 16718 29 16719
rect 30 16718 34 16764
rect 54 16718 58 16764
rect 78 16718 82 16764
rect 102 16718 106 16764
rect 126 16718 130 16764
rect 150 16718 154 16764
rect 174 16718 178 16764
rect 198 16718 202 16764
rect 222 16718 226 16764
rect 246 16718 250 16764
rect 270 16718 274 16764
rect 294 16718 298 16764
rect 318 16718 322 16764
rect 342 16718 346 16764
rect 366 16718 370 16764
rect 390 16718 394 16764
rect 414 16718 418 16764
rect 438 16718 442 16764
rect 462 16718 466 16764
rect 486 16718 490 16764
rect 510 16718 514 16764
rect 534 16718 538 16764
rect 558 16718 562 16764
rect 582 16718 586 16764
rect 606 16718 610 16764
rect 630 16718 634 16764
rect 654 16718 658 16764
rect 678 16718 682 16764
rect 702 16718 706 16764
rect 726 16718 730 16764
rect 750 16718 754 16764
rect 774 16718 778 16764
rect 798 16718 802 16764
rect 822 16718 826 16764
rect 846 16718 850 16764
rect 870 16718 874 16764
rect 894 16718 898 16764
rect 918 16718 922 16764
rect 942 16718 946 16764
rect 966 16718 970 16764
rect 990 16718 994 16764
rect 1014 16718 1018 16764
rect 1038 16718 1042 16764
rect 1062 16718 1066 16764
rect 1086 16718 1090 16764
rect 1110 16718 1114 16764
rect 1134 16718 1138 16764
rect 1158 16718 1162 16764
rect 1182 16718 1186 16764
rect 1206 16739 1210 16764
rect -5 16716 1203 16718
rect -5 16709 0 16716
rect 5 16695 10 16709
rect 6 16670 10 16695
rect 30 16670 34 16716
rect 54 16670 58 16716
rect 78 16670 82 16716
rect 102 16670 106 16716
rect 126 16670 130 16716
rect 150 16670 154 16716
rect 174 16670 178 16716
rect 198 16670 202 16716
rect 222 16670 226 16716
rect 246 16670 250 16716
rect 270 16670 274 16716
rect 294 16670 298 16716
rect 318 16670 322 16716
rect 342 16670 346 16716
rect 366 16670 370 16716
rect 390 16670 394 16716
rect 414 16670 418 16716
rect 438 16670 442 16716
rect 462 16670 466 16716
rect 486 16670 490 16716
rect 510 16670 514 16716
rect 534 16670 538 16716
rect 558 16670 562 16716
rect 582 16670 586 16716
rect 606 16670 610 16716
rect 630 16670 634 16716
rect 654 16670 658 16716
rect 678 16670 682 16716
rect 702 16670 706 16716
rect 726 16670 730 16716
rect 750 16670 754 16716
rect 774 16670 778 16716
rect 798 16670 802 16716
rect 822 16670 826 16716
rect 846 16670 850 16716
rect 870 16670 874 16716
rect 894 16670 898 16716
rect 918 16670 922 16716
rect 942 16670 946 16716
rect 966 16670 970 16716
rect 990 16670 994 16716
rect 1014 16670 1018 16716
rect 1038 16670 1042 16716
rect 1062 16670 1066 16716
rect 1086 16670 1090 16716
rect 1110 16670 1114 16716
rect 1134 16670 1138 16716
rect 1158 16670 1162 16716
rect 1182 16670 1186 16716
rect 1189 16715 1203 16716
rect 1206 16691 1213 16739
rect 1206 16670 1210 16691
rect 1230 16670 1234 16764
rect 1254 16670 1258 16764
rect 1278 16670 1282 16764
rect 1302 16670 1306 16764
rect 1326 16670 1330 16764
rect 1350 16670 1354 16764
rect 1374 16670 1378 16764
rect 1398 16670 1402 16764
rect 1422 16670 1426 16764
rect 1446 16670 1450 16764
rect 1470 16670 1474 16764
rect 1494 16670 1498 16764
rect 1518 16670 1522 16764
rect 1542 16670 1546 16764
rect 1566 16670 1570 16764
rect 1590 16670 1594 16764
rect 1614 16670 1618 16764
rect 1638 16670 1642 16764
rect 1662 16670 1666 16764
rect 1686 16670 1690 16764
rect 1710 16670 1714 16764
rect 1734 16670 1738 16764
rect 1758 16670 1762 16764
rect 1765 16763 1779 16764
rect 1782 16763 1789 16787
rect 1782 16718 1789 16739
rect 1806 16718 1810 16788
rect 1830 16718 1834 16788
rect 1854 16718 1858 16788
rect 1878 16718 1882 16788
rect 1902 16718 1906 16788
rect 1926 16718 1930 16788
rect 1950 16718 1954 16788
rect 1974 16718 1978 16788
rect 1998 16718 2002 16788
rect 2022 16718 2026 16788
rect 2046 16718 2050 16788
rect 2070 16718 2074 16788
rect 2094 16718 2098 16788
rect 2118 16718 2122 16788
rect 2142 16718 2146 16788
rect 2166 16718 2170 16788
rect 2190 16718 2194 16788
rect 2214 16718 2218 16788
rect 2238 16718 2242 16788
rect 2262 16718 2266 16788
rect 2286 16718 2290 16788
rect 2310 16718 2314 16788
rect 2334 16718 2338 16788
rect 2358 16718 2362 16788
rect 2382 16718 2386 16788
rect 2406 16718 2410 16788
rect 2430 16718 2434 16788
rect 2454 16718 2458 16788
rect 2478 16718 2482 16788
rect 2502 16718 2506 16788
rect 2526 16718 2530 16788
rect 2550 16718 2554 16788
rect 2574 16718 2578 16788
rect 2598 16718 2602 16788
rect 2622 16718 2626 16788
rect 2629 16787 2643 16788
rect 2646 16766 2653 16811
rect 2670 16766 2674 16812
rect 2694 16766 2698 16812
rect 2718 16766 2722 16812
rect 2742 16766 2746 16812
rect 2766 16766 2770 16812
rect 2790 16766 2794 16812
rect 2814 16766 2818 16812
rect 2838 16766 2842 16812
rect 2862 16766 2866 16812
rect 2886 16766 2890 16812
rect 2910 16766 2914 16812
rect 2934 16766 2938 16812
rect 2958 16766 2962 16812
rect 2971 16766 3005 16767
rect 2629 16764 3005 16766
rect 2629 16763 2643 16764
rect 2646 16763 2653 16764
rect 2646 16718 2650 16763
rect 2670 16718 2674 16764
rect 2694 16718 2698 16764
rect 2718 16718 2722 16764
rect 2742 16718 2746 16764
rect 2766 16718 2770 16764
rect 2790 16718 2794 16764
rect 2814 16718 2818 16764
rect 2838 16718 2842 16764
rect 2862 16718 2866 16764
rect 2886 16718 2890 16764
rect 2910 16718 2914 16764
rect 2934 16718 2938 16764
rect 2958 16718 2962 16764
rect 2971 16757 2976 16764
rect 3006 16763 3010 16812
rect 2981 16743 2986 16757
rect 2995 16753 3003 16757
rect 2989 16743 2995 16753
rect 2982 16718 2986 16743
rect 3006 16739 3013 16763
rect 3030 16718 3034 16812
rect 3054 16718 3058 16812
rect 3078 16718 3082 16812
rect 3102 16718 3106 16812
rect 3126 16718 3130 16812
rect 3150 16718 3154 16812
rect 3174 16718 3178 16812
rect 3198 16718 3202 16812
rect 3222 16718 3226 16812
rect 3246 16718 3250 16812
rect 3270 16718 3274 16812
rect 3294 16718 3298 16812
rect 3318 16718 3322 16812
rect 3342 16718 3346 16812
rect 3366 16718 3370 16812
rect 3390 16718 3394 16812
rect 3414 16718 3418 16812
rect 3438 16718 3442 16812
rect 3462 16718 3466 16812
rect 3486 16718 3490 16812
rect 3510 16718 3514 16812
rect 3534 16718 3538 16812
rect 3558 16718 3562 16812
rect 3582 16718 3586 16812
rect 3606 16718 3610 16812
rect 3630 16718 3634 16812
rect 3654 16718 3658 16812
rect 3678 16718 3682 16812
rect 3702 16718 3706 16812
rect 3726 16718 3730 16812
rect 3750 16719 3754 16812
rect 3763 16781 3768 16791
rect 3774 16781 3778 16812
rect 3787 16805 3792 16812
rect 3798 16805 3802 16812
rect 3797 16791 3802 16805
rect 3773 16767 3778 16781
rect 3739 16718 3773 16719
rect 1765 16716 3773 16718
rect 1765 16715 1779 16716
rect 1782 16715 1789 16716
rect 1782 16670 1786 16715
rect 1806 16670 1810 16716
rect 1830 16670 1834 16716
rect 1854 16670 1858 16716
rect 1878 16670 1882 16716
rect 1902 16670 1906 16716
rect 1926 16670 1930 16716
rect 1950 16670 1954 16716
rect 1974 16670 1978 16716
rect 1998 16670 2002 16716
rect 2022 16670 2026 16716
rect 2046 16670 2050 16716
rect 2070 16670 2074 16716
rect 2094 16670 2098 16716
rect 2118 16670 2122 16716
rect 2142 16670 2146 16716
rect 2166 16670 2170 16716
rect 2190 16670 2194 16716
rect 2214 16670 2218 16716
rect 2238 16670 2242 16716
rect 2262 16670 2266 16716
rect 2286 16670 2290 16716
rect 2310 16670 2314 16716
rect 2334 16670 2338 16716
rect 2358 16670 2362 16716
rect 2382 16670 2386 16716
rect 2406 16670 2410 16716
rect 2430 16670 2434 16716
rect 2454 16670 2458 16716
rect 2478 16670 2482 16716
rect 2502 16670 2506 16716
rect 2526 16670 2530 16716
rect 2550 16670 2554 16716
rect 2574 16670 2578 16716
rect 2598 16670 2602 16716
rect 2622 16670 2626 16716
rect 2646 16670 2650 16716
rect 2670 16670 2674 16716
rect 2694 16670 2698 16716
rect 2718 16670 2722 16716
rect 2742 16670 2746 16716
rect 2766 16670 2770 16716
rect 2790 16670 2794 16716
rect 2814 16670 2818 16716
rect 2838 16670 2842 16716
rect 2862 16670 2866 16716
rect 2886 16670 2890 16716
rect 2910 16670 2914 16716
rect 2934 16670 2938 16716
rect 2958 16670 2962 16716
rect 2982 16670 2986 16716
rect -2393 16668 3003 16670
rect -2371 16646 -2366 16668
rect -2348 16646 -2343 16668
rect -2325 16646 -2320 16668
rect -2054 16667 -1906 16668
rect -2054 16666 -2036 16667
rect -2309 16652 -2301 16662
rect -2317 16646 -2309 16652
rect -2068 16651 -2038 16658
rect -2000 16650 -1992 16667
rect -1920 16666 -1906 16667
rect -1846 16660 -1794 16668
rect -1852 16653 -1804 16658
rect -1902 16651 -1804 16653
rect -1655 16652 -1647 16662
rect -2000 16648 -1975 16650
rect -1902 16649 -1852 16651
rect -2025 16646 -1975 16648
rect -1846 16646 -1804 16649
rect -1663 16646 -1655 16652
rect -1642 16646 -1637 16668
rect -1619 16646 -1614 16668
rect -1530 16646 -1526 16668
rect -1506 16646 -1502 16668
rect -1482 16646 -1478 16668
rect -1458 16646 -1454 16668
rect -1434 16646 -1430 16668
rect -1410 16646 -1406 16668
rect -1386 16646 -1382 16668
rect -1362 16646 -1358 16668
rect -1338 16646 -1334 16668
rect -1314 16646 -1310 16668
rect -1290 16646 -1286 16668
rect -1266 16646 -1262 16668
rect -1242 16646 -1238 16668
rect -1218 16646 -1214 16668
rect -1194 16646 -1190 16668
rect -1170 16646 -1166 16668
rect -1146 16646 -1142 16668
rect -1122 16646 -1118 16668
rect -1098 16646 -1094 16668
rect -1074 16646 -1070 16668
rect -1050 16646 -1046 16668
rect -1026 16646 -1022 16668
rect -1002 16646 -998 16668
rect -978 16646 -974 16668
rect -954 16646 -950 16668
rect -930 16646 -926 16668
rect -906 16646 -902 16668
rect -882 16646 -878 16668
rect -858 16646 -854 16668
rect -834 16646 -830 16668
rect -810 16646 -806 16668
rect -786 16646 -782 16668
rect -762 16646 -758 16668
rect -738 16646 -734 16668
rect -714 16646 -710 16668
rect -690 16646 -686 16668
rect -666 16646 -662 16668
rect -642 16646 -638 16668
rect -618 16646 -614 16668
rect -594 16646 -590 16668
rect -570 16646 -566 16668
rect -546 16646 -542 16668
rect -522 16646 -518 16668
rect -498 16646 -494 16668
rect -474 16646 -470 16668
rect -450 16646 -446 16668
rect -426 16646 -422 16668
rect -402 16646 -398 16668
rect -378 16646 -374 16668
rect -354 16646 -350 16668
rect -330 16646 -326 16668
rect -306 16646 -302 16668
rect -282 16646 -278 16668
rect -258 16646 -254 16668
rect -234 16646 -230 16668
rect -210 16646 -206 16668
rect -186 16646 -182 16668
rect -162 16646 -158 16668
rect -138 16646 -134 16668
rect -114 16646 -110 16668
rect -90 16646 -86 16668
rect -66 16646 -62 16668
rect -42 16646 -38 16668
rect -18 16646 -14 16668
rect 6 16646 10 16668
rect 30 16667 34 16668
rect -2393 16644 27 16646
rect -2371 16622 -2366 16644
rect -2348 16622 -2343 16644
rect -2325 16622 -2320 16644
rect -2054 16643 -2038 16644
rect -2000 16643 -1966 16644
rect -1846 16643 -1804 16644
rect -2000 16642 -1975 16643
rect -2076 16634 -2054 16641
rect -2309 16624 -2301 16634
rect -2044 16631 -2038 16636
rect -2028 16634 -2001 16641
rect -2054 16624 -2038 16631
rect -2015 16633 -2001 16634
rect -2015 16624 -2014 16633
rect -2317 16622 -2309 16624
rect -2044 16622 -2028 16624
rect -2000 16622 -1992 16642
rect -1982 16641 -1975 16642
rect -1862 16641 -1798 16642
rect -1985 16634 -1796 16641
rect -1862 16633 -1798 16634
rect -1852 16624 -1804 16631
rect -1655 16624 -1647 16634
rect -1976 16622 -1940 16623
rect -1663 16622 -1655 16624
rect -1642 16622 -1637 16644
rect -1619 16622 -1614 16644
rect -1530 16622 -1526 16644
rect -1506 16622 -1502 16644
rect -1482 16643 -1478 16644
rect -2393 16620 -1485 16622
rect -2371 16550 -2366 16620
rect -2348 16550 -2343 16620
rect -2325 16586 -2320 16620
rect -2317 16618 -2309 16620
rect -2076 16607 -2054 16614
rect -2325 16578 -2317 16586
rect -2060 16580 -2030 16583
rect -2325 16550 -2320 16578
rect -2317 16570 -2309 16578
rect -2060 16567 -2038 16578
rect -2033 16571 -2030 16580
rect -2028 16576 -2027 16580
rect -2068 16562 -2038 16565
rect -2000 16550 -1992 16620
rect -1846 16616 -1804 16620
rect -1663 16618 -1655 16620
rect -1846 16606 -1794 16615
rect -1912 16595 -1884 16597
rect -1852 16589 -1804 16593
rect -1844 16580 -1796 16583
rect -1671 16578 -1663 16586
rect -1844 16567 -1804 16578
rect -1663 16570 -1655 16578
rect -1852 16562 -1680 16566
rect -1642 16550 -1637 16620
rect -1619 16550 -1614 16620
rect -1530 16550 -1526 16620
rect -1506 16550 -1502 16620
rect -1499 16619 -1485 16620
rect -1482 16619 -1475 16643
rect -1482 16550 -1478 16619
rect -1458 16550 -1454 16644
rect -1434 16550 -1430 16644
rect -1410 16550 -1406 16644
rect -1386 16550 -1382 16644
rect -1362 16550 -1358 16644
rect -1338 16550 -1334 16644
rect -1314 16550 -1310 16644
rect -1290 16550 -1286 16644
rect -1266 16550 -1262 16644
rect -1242 16550 -1238 16644
rect -1218 16550 -1214 16644
rect -1194 16550 -1190 16644
rect -1170 16550 -1166 16644
rect -1146 16550 -1142 16644
rect -1122 16550 -1118 16644
rect -1098 16550 -1094 16644
rect -1074 16550 -1070 16644
rect -1050 16550 -1046 16644
rect -1026 16550 -1022 16644
rect -1002 16550 -998 16644
rect -978 16550 -974 16644
rect -954 16550 -950 16644
rect -930 16550 -926 16644
rect -906 16550 -902 16644
rect -882 16550 -878 16644
rect -858 16550 -854 16644
rect -834 16550 -830 16644
rect -810 16550 -806 16644
rect -786 16550 -782 16644
rect -773 16589 -768 16599
rect -762 16589 -758 16644
rect -763 16575 -758 16589
rect -773 16574 -739 16575
rect -738 16574 -734 16644
rect -714 16574 -710 16644
rect -690 16574 -686 16644
rect -666 16574 -662 16644
rect -642 16574 -638 16644
rect -618 16574 -614 16644
rect -594 16574 -590 16644
rect -570 16574 -566 16644
rect -546 16574 -542 16644
rect -522 16574 -518 16644
rect -498 16574 -494 16644
rect -474 16574 -470 16644
rect -450 16574 -446 16644
rect -426 16574 -422 16644
rect -402 16574 -398 16644
rect -378 16574 -374 16644
rect -354 16574 -350 16644
rect -330 16574 -326 16644
rect -306 16574 -302 16644
rect -293 16613 -288 16623
rect -282 16613 -278 16644
rect -283 16599 -278 16613
rect -282 16574 -278 16599
rect -258 16574 -254 16644
rect -234 16574 -230 16644
rect -210 16574 -206 16644
rect -186 16574 -182 16644
rect -162 16574 -158 16644
rect -138 16574 -134 16644
rect -114 16574 -110 16644
rect -90 16574 -86 16644
rect -66 16574 -62 16644
rect -42 16574 -38 16644
rect -18 16574 -14 16644
rect 6 16574 10 16644
rect 13 16643 27 16644
rect 30 16619 37 16667
rect 30 16574 34 16619
rect 54 16574 58 16668
rect 78 16574 82 16668
rect 102 16574 106 16668
rect 126 16574 130 16668
rect 150 16574 154 16668
rect 174 16574 178 16668
rect 198 16574 202 16668
rect 222 16574 226 16668
rect 246 16574 250 16668
rect 270 16574 274 16668
rect 294 16574 298 16668
rect 318 16574 322 16668
rect 342 16574 346 16668
rect 366 16574 370 16668
rect 390 16574 394 16668
rect 414 16574 418 16668
rect 438 16574 442 16668
rect 462 16574 466 16668
rect 486 16574 490 16668
rect 510 16574 514 16668
rect 534 16574 538 16668
rect 558 16574 562 16668
rect 582 16574 586 16668
rect 606 16574 610 16668
rect 630 16574 634 16668
rect 654 16574 658 16668
rect 678 16574 682 16668
rect 702 16574 706 16668
rect 726 16574 730 16668
rect 750 16574 754 16668
rect 774 16574 778 16668
rect 798 16574 802 16668
rect 822 16574 826 16668
rect 846 16574 850 16668
rect 870 16574 874 16668
rect 894 16574 898 16668
rect 918 16574 922 16668
rect 942 16574 946 16668
rect 966 16574 970 16668
rect 990 16574 994 16668
rect 1014 16574 1018 16668
rect 1038 16574 1042 16668
rect 1062 16574 1066 16668
rect 1086 16574 1090 16668
rect 1110 16574 1114 16668
rect 1134 16574 1138 16668
rect 1158 16574 1162 16668
rect 1182 16574 1186 16668
rect 1206 16574 1210 16668
rect 1230 16574 1234 16668
rect 1254 16574 1258 16668
rect 1278 16574 1282 16668
rect 1302 16574 1306 16668
rect 1326 16574 1330 16668
rect 1350 16574 1354 16668
rect 1374 16574 1378 16668
rect 1398 16574 1402 16668
rect 1422 16574 1426 16668
rect 1446 16574 1450 16668
rect 1470 16574 1474 16668
rect 1494 16574 1498 16668
rect 1518 16574 1522 16668
rect 1542 16574 1546 16668
rect 1566 16574 1570 16668
rect 1590 16574 1594 16668
rect 1614 16574 1618 16668
rect 1638 16574 1642 16668
rect 1662 16574 1666 16668
rect 1686 16574 1690 16668
rect 1710 16574 1714 16668
rect 1734 16574 1738 16668
rect 1758 16574 1762 16668
rect 1782 16574 1786 16668
rect 1806 16574 1810 16668
rect 1830 16574 1834 16668
rect 1854 16574 1858 16668
rect 1878 16574 1882 16668
rect 1902 16574 1906 16668
rect 1926 16574 1930 16668
rect 1950 16574 1954 16668
rect 1974 16574 1978 16668
rect 1998 16574 2002 16668
rect 2022 16574 2026 16668
rect 2046 16574 2050 16668
rect 2070 16574 2074 16668
rect 2094 16574 2098 16668
rect 2118 16574 2122 16668
rect 2142 16574 2146 16668
rect 2166 16574 2170 16668
rect 2190 16574 2194 16668
rect 2214 16574 2218 16668
rect 2238 16574 2242 16668
rect 2262 16574 2266 16668
rect 2286 16574 2290 16668
rect 2310 16574 2314 16668
rect 2334 16574 2338 16668
rect 2358 16574 2362 16668
rect 2382 16574 2386 16668
rect 2406 16574 2410 16668
rect 2430 16574 2434 16668
rect 2454 16574 2458 16668
rect 2478 16574 2482 16668
rect 2502 16574 2506 16668
rect 2526 16574 2530 16668
rect 2539 16637 2544 16647
rect 2550 16637 2554 16668
rect 2549 16623 2554 16637
rect 2550 16574 2554 16623
rect 2574 16574 2578 16668
rect 2598 16574 2602 16668
rect 2622 16574 2626 16668
rect 2646 16574 2650 16668
rect 2670 16574 2674 16668
rect 2694 16574 2698 16668
rect 2718 16574 2722 16668
rect 2742 16574 2746 16668
rect 2766 16574 2770 16668
rect 2790 16574 2794 16668
rect 2814 16574 2818 16668
rect 2838 16574 2842 16668
rect 2862 16574 2866 16668
rect 2886 16574 2890 16668
rect 2910 16574 2914 16668
rect 2934 16574 2938 16668
rect 2958 16574 2962 16668
rect 2982 16574 2986 16668
rect 2989 16667 3003 16668
rect 3006 16667 3013 16691
rect 3006 16574 3010 16667
rect 3030 16574 3034 16716
rect 3054 16574 3058 16716
rect 3078 16574 3082 16716
rect 3102 16574 3106 16716
rect 3126 16574 3130 16716
rect 3150 16574 3154 16716
rect 3174 16574 3178 16716
rect 3198 16574 3202 16716
rect 3222 16574 3226 16716
rect 3246 16574 3250 16716
rect 3270 16574 3274 16716
rect 3294 16574 3298 16716
rect 3318 16574 3322 16716
rect 3342 16574 3346 16716
rect 3366 16574 3370 16716
rect 3390 16574 3394 16716
rect 3414 16574 3418 16716
rect 3438 16574 3442 16716
rect 3462 16574 3466 16716
rect 3486 16574 3490 16716
rect 3510 16574 3514 16716
rect 3534 16574 3538 16716
rect 3558 16574 3562 16716
rect 3582 16574 3586 16716
rect 3606 16574 3610 16716
rect 3630 16574 3634 16716
rect 3654 16574 3658 16716
rect 3678 16574 3682 16716
rect 3702 16574 3706 16716
rect 3726 16574 3730 16716
rect 3739 16709 3744 16716
rect 3750 16709 3754 16716
rect 3749 16695 3754 16709
rect 3739 16661 3744 16671
rect 3749 16647 3754 16661
rect 3750 16575 3754 16647
rect 3739 16574 3771 16575
rect -773 16572 3771 16574
rect -773 16565 -768 16572
rect -763 16551 -758 16565
rect -762 16550 -758 16551
rect -738 16550 -734 16572
rect -714 16550 -710 16572
rect -690 16550 -686 16572
rect -666 16550 -662 16572
rect -642 16550 -638 16572
rect -618 16550 -614 16572
rect -594 16550 -590 16572
rect -570 16550 -566 16572
rect -546 16550 -542 16572
rect -522 16550 -518 16572
rect -498 16550 -494 16572
rect -474 16550 -470 16572
rect -450 16550 -446 16572
rect -426 16550 -422 16572
rect -402 16550 -398 16572
rect -378 16550 -374 16572
rect -354 16550 -350 16572
rect -330 16550 -326 16572
rect -306 16550 -302 16572
rect -282 16550 -278 16572
rect -258 16550 -254 16572
rect -234 16550 -230 16572
rect -210 16550 -206 16572
rect -186 16550 -182 16572
rect -162 16550 -158 16572
rect -138 16550 -134 16572
rect -114 16550 -110 16572
rect -90 16550 -86 16572
rect -66 16550 -62 16572
rect -42 16550 -38 16572
rect -18 16550 -14 16572
rect 6 16550 10 16572
rect 30 16550 34 16572
rect 54 16550 58 16572
rect 78 16550 82 16572
rect 102 16550 106 16572
rect 126 16550 130 16572
rect 150 16550 154 16572
rect 174 16550 178 16572
rect 198 16550 202 16572
rect 222 16550 226 16572
rect 246 16550 250 16572
rect 270 16550 274 16572
rect 294 16550 298 16572
rect 318 16550 322 16572
rect 342 16550 346 16572
rect 366 16550 370 16572
rect 390 16550 394 16572
rect 414 16550 418 16572
rect 438 16550 442 16572
rect 462 16550 466 16572
rect 486 16550 490 16572
rect 510 16550 514 16572
rect 534 16550 538 16572
rect 558 16550 562 16572
rect 582 16550 586 16572
rect 606 16550 610 16572
rect 630 16550 634 16572
rect 654 16550 658 16572
rect 678 16550 682 16572
rect 702 16550 706 16572
rect 726 16550 730 16572
rect 750 16550 754 16572
rect 774 16550 778 16572
rect 798 16550 802 16572
rect 822 16550 826 16572
rect 846 16550 850 16572
rect 870 16550 874 16572
rect 894 16550 898 16572
rect 918 16550 922 16572
rect 942 16550 946 16572
rect 966 16550 970 16572
rect 990 16550 994 16572
rect 1014 16550 1018 16572
rect 1038 16550 1042 16572
rect 1062 16550 1066 16572
rect 1086 16550 1090 16572
rect 1110 16550 1114 16572
rect 1134 16550 1138 16572
rect 1158 16550 1162 16572
rect 1182 16550 1186 16572
rect 1206 16550 1210 16572
rect 1230 16550 1234 16572
rect 1254 16550 1258 16572
rect 1278 16550 1282 16572
rect 1302 16550 1306 16572
rect 1326 16550 1330 16572
rect 1350 16550 1354 16572
rect 1374 16550 1378 16572
rect 1398 16550 1402 16572
rect 1422 16550 1426 16572
rect 1446 16550 1450 16572
rect 1470 16550 1474 16572
rect 1494 16550 1498 16572
rect 1518 16550 1522 16572
rect 1542 16550 1546 16572
rect 1566 16550 1570 16572
rect 1590 16550 1594 16572
rect 1614 16550 1618 16572
rect 1638 16550 1642 16572
rect 1662 16550 1666 16572
rect 1686 16550 1690 16572
rect 1710 16550 1714 16572
rect 1734 16550 1738 16572
rect 1758 16550 1762 16572
rect 1782 16550 1786 16572
rect 1806 16550 1810 16572
rect 1830 16550 1834 16572
rect 1854 16550 1858 16572
rect 1878 16550 1882 16572
rect 1902 16550 1906 16572
rect 1926 16550 1930 16572
rect 1950 16550 1954 16572
rect 1974 16550 1978 16572
rect 1998 16550 2002 16572
rect 2022 16550 2026 16572
rect 2046 16550 2050 16572
rect 2070 16550 2074 16572
rect 2094 16550 2098 16572
rect 2118 16550 2122 16572
rect 2142 16550 2146 16572
rect 2166 16550 2170 16572
rect 2190 16550 2194 16572
rect 2214 16550 2218 16572
rect 2238 16550 2242 16572
rect 2262 16550 2266 16572
rect 2286 16550 2290 16572
rect 2310 16550 2314 16572
rect 2334 16550 2338 16572
rect 2358 16550 2362 16572
rect 2382 16550 2386 16572
rect 2406 16550 2410 16572
rect 2430 16550 2434 16572
rect 2454 16550 2458 16572
rect 2478 16550 2482 16572
rect 2502 16550 2506 16572
rect 2526 16550 2530 16572
rect 2550 16550 2554 16572
rect 2574 16571 2578 16572
rect -2393 16548 2571 16550
rect -2371 16526 -2366 16548
rect -2348 16526 -2343 16548
rect -2325 16526 -2320 16548
rect -2309 16530 -2301 16540
rect -2068 16531 -2062 16536
rect -2317 16526 -2309 16530
rect -2060 16526 -2050 16531
rect -2000 16526 -1992 16548
rect -1806 16540 -1680 16546
rect -1854 16531 -1806 16536
rect -1655 16530 -1647 16540
rect -1972 16526 -1964 16527
rect -1958 16526 -1942 16528
rect -1844 16526 -1806 16529
rect -1663 16526 -1655 16530
rect -1642 16526 -1637 16548
rect -1619 16526 -1614 16548
rect -1530 16526 -1526 16548
rect -1506 16526 -1502 16548
rect -1482 16526 -1478 16548
rect -1458 16526 -1454 16548
rect -1434 16526 -1430 16548
rect -1410 16526 -1406 16548
rect -1386 16526 -1382 16548
rect -1362 16526 -1358 16548
rect -1338 16526 -1334 16548
rect -1314 16526 -1310 16548
rect -1290 16526 -1286 16548
rect -1266 16526 -1262 16548
rect -1242 16526 -1238 16548
rect -1218 16526 -1214 16548
rect -1194 16526 -1190 16548
rect -1170 16526 -1166 16548
rect -1146 16526 -1142 16548
rect -1122 16526 -1118 16548
rect -1098 16526 -1094 16548
rect -1074 16526 -1070 16548
rect -1050 16526 -1046 16548
rect -1026 16526 -1022 16548
rect -1002 16526 -998 16548
rect -978 16526 -974 16548
rect -954 16526 -950 16548
rect -930 16526 -926 16548
rect -906 16526 -902 16548
rect -882 16526 -878 16548
rect -858 16526 -854 16548
rect -834 16526 -830 16548
rect -810 16526 -806 16548
rect -786 16526 -782 16548
rect -762 16526 -758 16548
rect -738 16526 -734 16548
rect -714 16526 -710 16548
rect -690 16526 -686 16548
rect -666 16526 -662 16548
rect -642 16526 -638 16548
rect -618 16526 -614 16548
rect -594 16526 -590 16548
rect -570 16526 -566 16548
rect -546 16526 -542 16548
rect -522 16526 -518 16548
rect -498 16526 -494 16548
rect -474 16526 -470 16548
rect -450 16527 -446 16548
rect -461 16526 -427 16527
rect -2393 16524 -427 16526
rect -2371 16502 -2366 16524
rect -2348 16502 -2343 16524
rect -2325 16502 -2320 16524
rect -2060 16518 -2050 16524
rect -2309 16502 -2301 16512
rect -2060 16511 -2030 16518
rect -2000 16514 -1992 16524
rect -1972 16522 -1942 16524
rect -1958 16521 -1942 16522
rect -1844 16520 -1806 16524
rect -2068 16504 -2062 16511
rect -2062 16502 -2036 16504
rect -2393 16500 -2036 16502
rect -2030 16502 -2012 16504
rect -2004 16502 -1990 16514
rect -1844 16513 -1798 16518
rect -1806 16511 -1798 16513
rect -1854 16509 -1844 16511
rect -1854 16504 -1806 16509
rect -1864 16502 -1796 16503
rect -1655 16502 -1647 16512
rect -1642 16502 -1637 16524
rect -1619 16502 -1614 16524
rect -1530 16502 -1526 16524
rect -1506 16502 -1502 16524
rect -1482 16502 -1478 16524
rect -1458 16502 -1454 16524
rect -1434 16502 -1430 16524
rect -1410 16502 -1406 16524
rect -1386 16502 -1382 16524
rect -1362 16502 -1358 16524
rect -1338 16502 -1334 16524
rect -1314 16502 -1310 16524
rect -1290 16502 -1286 16524
rect -1266 16502 -1262 16524
rect -1242 16502 -1238 16524
rect -1218 16502 -1214 16524
rect -1194 16502 -1190 16524
rect -1170 16502 -1166 16524
rect -1146 16502 -1142 16524
rect -1122 16502 -1118 16524
rect -1098 16502 -1094 16524
rect -1074 16502 -1070 16524
rect -1050 16502 -1046 16524
rect -1026 16502 -1022 16524
rect -1002 16503 -998 16524
rect -1013 16502 -979 16503
rect -2030 16500 -979 16502
rect -2371 16454 -2366 16500
rect -2348 16454 -2343 16500
rect -2325 16454 -2320 16500
rect -2317 16496 -2309 16500
rect -2060 16496 -2050 16500
rect -2060 16494 -2036 16496
rect -2060 16492 -2030 16494
rect -2292 16486 -2030 16492
rect -2092 16470 -2062 16472
rect -2094 16466 -2062 16470
rect -2000 16454 -1992 16500
rect -1844 16493 -1806 16500
rect -1663 16496 -1655 16500
rect -1844 16486 -1680 16492
rect -1854 16470 -1806 16472
rect -1854 16466 -1680 16470
rect -1926 16454 -1892 16457
rect -1642 16454 -1637 16500
rect -1619 16454 -1614 16500
rect -1530 16454 -1526 16500
rect -1506 16454 -1502 16500
rect -1482 16454 -1478 16500
rect -1458 16454 -1454 16500
rect -1434 16454 -1430 16500
rect -1410 16454 -1406 16500
rect -1386 16454 -1382 16500
rect -1362 16454 -1358 16500
rect -1338 16454 -1334 16500
rect -1314 16454 -1310 16500
rect -1290 16454 -1286 16500
rect -1266 16454 -1262 16500
rect -1242 16454 -1238 16500
rect -1218 16454 -1214 16500
rect -1194 16454 -1190 16500
rect -1170 16454 -1166 16500
rect -1146 16454 -1142 16500
rect -1122 16454 -1118 16500
rect -1098 16454 -1094 16500
rect -1074 16454 -1070 16500
rect -1050 16454 -1046 16500
rect -1026 16454 -1022 16500
rect -1013 16493 -1008 16500
rect -1002 16493 -998 16500
rect -1003 16479 -998 16493
rect -1013 16469 -1008 16479
rect -1003 16455 -998 16469
rect -1002 16454 -998 16455
rect -978 16454 -974 16524
rect -954 16454 -950 16524
rect -930 16454 -926 16524
rect -906 16454 -902 16524
rect -882 16454 -878 16524
rect -858 16454 -854 16524
rect -834 16454 -830 16524
rect -810 16454 -806 16524
rect -786 16454 -782 16524
rect -762 16454 -758 16524
rect -738 16523 -734 16524
rect -738 16478 -731 16523
rect -714 16478 -710 16524
rect -690 16478 -686 16524
rect -666 16478 -662 16524
rect -642 16478 -638 16524
rect -618 16478 -614 16524
rect -594 16478 -590 16524
rect -570 16478 -566 16524
rect -546 16478 -542 16524
rect -522 16478 -518 16524
rect -498 16478 -494 16524
rect -474 16478 -470 16524
rect -461 16517 -456 16524
rect -450 16517 -446 16524
rect -451 16503 -446 16517
rect -461 16493 -456 16503
rect -451 16479 -446 16493
rect -450 16478 -446 16479
rect -426 16478 -422 16548
rect -402 16478 -398 16548
rect -378 16478 -374 16548
rect -354 16478 -350 16548
rect -330 16478 -326 16548
rect -306 16478 -302 16548
rect -282 16478 -278 16548
rect -258 16547 -254 16548
rect -258 16523 -251 16547
rect -258 16478 -254 16523
rect -234 16478 -230 16548
rect -210 16478 -206 16548
rect -186 16478 -182 16548
rect -162 16478 -158 16548
rect -138 16478 -134 16548
rect -114 16478 -110 16548
rect -90 16478 -86 16548
rect -66 16478 -62 16548
rect -42 16478 -38 16548
rect -18 16478 -14 16548
rect 6 16478 10 16548
rect 30 16478 34 16548
rect 54 16478 58 16548
rect 78 16478 82 16548
rect 102 16478 106 16548
rect 126 16478 130 16548
rect 150 16478 154 16548
rect 174 16478 178 16548
rect 198 16478 202 16548
rect 222 16478 226 16548
rect 246 16478 250 16548
rect 270 16478 274 16548
rect 294 16478 298 16548
rect 318 16478 322 16548
rect 342 16478 346 16548
rect 366 16478 370 16548
rect 390 16478 394 16548
rect 414 16478 418 16548
rect 438 16478 442 16548
rect 462 16478 466 16548
rect 486 16478 490 16548
rect 510 16478 514 16548
rect 534 16478 538 16548
rect 558 16478 562 16548
rect 582 16478 586 16548
rect 606 16478 610 16548
rect 630 16478 634 16548
rect 654 16478 658 16548
rect 678 16478 682 16548
rect 702 16478 706 16548
rect 726 16478 730 16548
rect 750 16478 754 16548
rect 774 16478 778 16548
rect 798 16478 802 16548
rect 822 16478 826 16548
rect 846 16478 850 16548
rect 870 16478 874 16548
rect 894 16478 898 16548
rect 918 16478 922 16548
rect 942 16478 946 16548
rect 966 16478 970 16548
rect 990 16478 994 16548
rect 1014 16478 1018 16548
rect 1038 16478 1042 16548
rect 1062 16478 1066 16548
rect 1086 16478 1090 16548
rect 1110 16478 1114 16548
rect 1134 16478 1138 16548
rect 1158 16478 1162 16548
rect 1182 16478 1186 16548
rect 1206 16478 1210 16548
rect 1230 16478 1234 16548
rect 1254 16478 1258 16548
rect 1278 16478 1282 16548
rect 1302 16478 1306 16548
rect 1326 16478 1330 16548
rect 1350 16478 1354 16548
rect 1374 16478 1378 16548
rect 1398 16478 1402 16548
rect 1422 16478 1426 16548
rect 1446 16478 1450 16548
rect 1470 16478 1474 16548
rect 1494 16478 1498 16548
rect 1518 16478 1522 16548
rect 1542 16478 1546 16548
rect 1566 16478 1570 16548
rect 1590 16478 1594 16548
rect 1614 16478 1618 16548
rect 1638 16478 1642 16548
rect 1662 16478 1666 16548
rect 1686 16478 1690 16548
rect 1710 16478 1714 16548
rect 1734 16478 1738 16548
rect 1758 16478 1762 16548
rect 1782 16478 1786 16548
rect 1806 16478 1810 16548
rect 1830 16478 1834 16548
rect 1854 16478 1858 16548
rect 1878 16478 1882 16548
rect 1902 16478 1906 16548
rect 1926 16478 1930 16548
rect 1950 16478 1954 16548
rect 1974 16478 1978 16548
rect 1998 16478 2002 16548
rect 2022 16478 2026 16548
rect 2046 16478 2050 16548
rect 2070 16478 2074 16548
rect 2094 16478 2098 16548
rect 2118 16478 2122 16548
rect 2142 16478 2146 16548
rect 2166 16478 2170 16548
rect 2190 16478 2194 16548
rect 2214 16478 2218 16548
rect 2238 16478 2242 16548
rect 2262 16478 2266 16548
rect 2286 16478 2290 16548
rect 2310 16478 2314 16548
rect 2334 16478 2338 16548
rect 2358 16478 2362 16548
rect 2382 16478 2386 16548
rect 2406 16478 2410 16548
rect 2430 16478 2434 16548
rect 2454 16478 2458 16548
rect 2478 16478 2482 16548
rect 2502 16478 2506 16548
rect 2526 16478 2530 16548
rect 2550 16478 2554 16548
rect 2557 16547 2571 16548
rect 2574 16547 2581 16571
rect 2574 16478 2578 16547
rect 2598 16478 2602 16572
rect 2622 16478 2626 16572
rect 2646 16478 2650 16572
rect 2670 16478 2674 16572
rect 2694 16478 2698 16572
rect 2718 16478 2722 16572
rect 2742 16478 2746 16572
rect 2766 16478 2770 16572
rect 2790 16478 2794 16572
rect 2814 16478 2818 16572
rect 2838 16478 2842 16572
rect 2862 16478 2866 16572
rect 2886 16478 2890 16572
rect 2910 16478 2914 16572
rect 2934 16478 2938 16572
rect 2958 16478 2962 16572
rect 2982 16478 2986 16572
rect 3006 16478 3010 16572
rect 3030 16478 3034 16572
rect 3054 16478 3058 16572
rect 3078 16478 3082 16572
rect 3102 16478 3106 16572
rect 3126 16478 3130 16572
rect 3150 16478 3154 16572
rect 3174 16478 3178 16572
rect 3198 16478 3202 16572
rect 3222 16478 3226 16572
rect 3246 16478 3250 16572
rect 3270 16478 3274 16572
rect 3294 16478 3298 16572
rect 3318 16478 3322 16572
rect 3342 16478 3346 16572
rect 3366 16478 3370 16572
rect 3390 16478 3394 16572
rect 3414 16478 3418 16572
rect 3438 16478 3442 16572
rect 3462 16478 3466 16572
rect 3486 16478 3490 16572
rect 3510 16478 3514 16572
rect 3534 16478 3538 16572
rect 3558 16478 3562 16572
rect 3582 16478 3586 16572
rect 3606 16478 3610 16572
rect 3630 16478 3634 16572
rect 3654 16478 3658 16572
rect 3678 16478 3682 16572
rect 3702 16478 3706 16572
rect 3726 16479 3730 16572
rect 3739 16565 3744 16572
rect 3750 16565 3754 16572
rect 3757 16571 3771 16572
rect 3749 16551 3754 16565
rect 3739 16541 3744 16551
rect 3749 16527 3754 16541
rect 3739 16493 3744 16503
rect 3750 16493 3754 16527
rect 3749 16479 3754 16493
rect 3763 16489 3771 16493
rect 3757 16479 3763 16489
rect 3715 16478 3749 16479
rect -755 16476 3749 16478
rect -755 16475 -741 16476
rect -738 16475 -731 16476
rect -738 16454 -734 16475
rect -714 16454 -710 16476
rect -690 16454 -686 16476
rect -666 16454 -662 16476
rect -642 16454 -638 16476
rect -618 16454 -614 16476
rect -594 16454 -590 16476
rect -570 16454 -566 16476
rect -546 16454 -542 16476
rect -522 16454 -518 16476
rect -498 16454 -494 16476
rect -474 16454 -470 16476
rect -450 16454 -446 16476
rect -426 16454 -422 16476
rect -402 16454 -398 16476
rect -378 16454 -374 16476
rect -354 16454 -350 16476
rect -330 16454 -326 16476
rect -306 16454 -302 16476
rect -282 16454 -278 16476
rect -258 16454 -254 16476
rect -234 16454 -230 16476
rect -210 16454 -206 16476
rect -186 16454 -182 16476
rect -162 16454 -158 16476
rect -138 16454 -134 16476
rect -114 16454 -110 16476
rect -90 16454 -86 16476
rect -66 16454 -62 16476
rect -42 16454 -38 16476
rect -18 16454 -14 16476
rect 6 16454 10 16476
rect 30 16454 34 16476
rect 54 16454 58 16476
rect 78 16454 82 16476
rect 102 16454 106 16476
rect 126 16454 130 16476
rect 150 16454 154 16476
rect 174 16454 178 16476
rect 198 16454 202 16476
rect 222 16454 226 16476
rect 246 16454 250 16476
rect 270 16454 274 16476
rect 294 16454 298 16476
rect 318 16454 322 16476
rect 342 16454 346 16476
rect 366 16454 370 16476
rect 390 16454 394 16476
rect 414 16454 418 16476
rect 438 16454 442 16476
rect 462 16454 466 16476
rect 486 16454 490 16476
rect 510 16454 514 16476
rect 534 16454 538 16476
rect 558 16454 562 16476
rect 582 16454 586 16476
rect 606 16454 610 16476
rect 630 16454 634 16476
rect 654 16454 658 16476
rect 678 16454 682 16476
rect 702 16454 706 16476
rect 726 16454 730 16476
rect 750 16454 754 16476
rect 774 16454 778 16476
rect 798 16454 802 16476
rect 822 16454 826 16476
rect 846 16454 850 16476
rect 870 16454 874 16476
rect 894 16454 898 16476
rect 918 16454 922 16476
rect 942 16454 946 16476
rect 966 16454 970 16476
rect 990 16454 994 16476
rect 1014 16454 1018 16476
rect 1038 16454 1042 16476
rect 1062 16454 1066 16476
rect 1086 16454 1090 16476
rect 1110 16454 1114 16476
rect 1134 16454 1138 16476
rect 1158 16454 1162 16476
rect 1182 16454 1186 16476
rect 1206 16454 1210 16476
rect 1230 16454 1234 16476
rect 1254 16454 1258 16476
rect 1278 16454 1282 16476
rect 1302 16454 1306 16476
rect 1326 16454 1330 16476
rect 1350 16454 1354 16476
rect 1374 16454 1378 16476
rect 1398 16454 1402 16476
rect 1422 16454 1426 16476
rect 1446 16454 1450 16476
rect 1470 16454 1474 16476
rect 1494 16454 1498 16476
rect 1518 16454 1522 16476
rect 1542 16454 1546 16476
rect 1566 16454 1570 16476
rect 1590 16454 1594 16476
rect 1614 16454 1618 16476
rect 1638 16454 1642 16476
rect 1662 16454 1666 16476
rect 1686 16454 1690 16476
rect 1710 16454 1714 16476
rect 1734 16454 1738 16476
rect 1758 16454 1762 16476
rect 1782 16454 1786 16476
rect 1806 16454 1810 16476
rect 1830 16454 1834 16476
rect 1854 16454 1858 16476
rect 1878 16454 1882 16476
rect 1902 16454 1906 16476
rect 1926 16454 1930 16476
rect 1950 16454 1954 16476
rect 1974 16454 1978 16476
rect 1998 16454 2002 16476
rect 2022 16454 2026 16476
rect 2046 16454 2050 16476
rect 2070 16454 2074 16476
rect 2094 16454 2098 16476
rect 2118 16454 2122 16476
rect 2142 16454 2146 16476
rect 2166 16454 2170 16476
rect 2190 16454 2194 16476
rect 2214 16454 2218 16476
rect 2238 16454 2242 16476
rect 2262 16454 2266 16476
rect 2286 16454 2290 16476
rect 2310 16454 2314 16476
rect 2334 16454 2338 16476
rect 2358 16454 2362 16476
rect 2382 16454 2386 16476
rect 2406 16454 2410 16476
rect 2430 16454 2434 16476
rect 2454 16454 2458 16476
rect 2478 16454 2482 16476
rect 2502 16454 2506 16476
rect 2526 16454 2530 16476
rect 2550 16454 2554 16476
rect 2574 16454 2578 16476
rect 2598 16454 2602 16476
rect 2622 16454 2626 16476
rect 2646 16454 2650 16476
rect 2670 16454 2674 16476
rect 2694 16454 2698 16476
rect 2718 16454 2722 16476
rect 2742 16454 2746 16476
rect 2766 16454 2770 16476
rect 2790 16454 2794 16476
rect 2814 16454 2818 16476
rect 2838 16454 2842 16476
rect 2862 16454 2866 16476
rect 2886 16454 2890 16476
rect 2910 16454 2914 16476
rect 2934 16454 2938 16476
rect 2958 16454 2962 16476
rect 2982 16454 2986 16476
rect 3006 16454 3010 16476
rect 3030 16454 3034 16476
rect 3054 16454 3058 16476
rect 3078 16454 3082 16476
rect 3102 16454 3106 16476
rect 3126 16454 3130 16476
rect 3150 16454 3154 16476
rect 3174 16454 3178 16476
rect 3198 16454 3202 16476
rect 3222 16454 3226 16476
rect 3246 16454 3250 16476
rect 3270 16454 3274 16476
rect 3294 16454 3298 16476
rect 3318 16454 3322 16476
rect 3342 16454 3346 16476
rect 3366 16454 3370 16476
rect 3390 16454 3394 16476
rect 3414 16454 3418 16476
rect 3438 16454 3442 16476
rect 3462 16454 3466 16476
rect 3486 16454 3490 16476
rect 3510 16454 3514 16476
rect 3534 16454 3538 16476
rect 3558 16454 3562 16476
rect 3582 16454 3586 16476
rect 3606 16454 3610 16476
rect 3630 16454 3634 16476
rect 3654 16454 3658 16476
rect 3678 16454 3682 16476
rect 3702 16454 3706 16476
rect 3715 16469 3720 16476
rect 3726 16469 3730 16476
rect 3725 16455 3730 16469
rect 3715 16454 3749 16455
rect -2393 16452 3749 16454
rect -2371 16430 -2366 16452
rect -2348 16430 -2343 16452
rect -2325 16430 -2320 16452
rect -2054 16451 -1906 16452
rect -2054 16450 -2036 16451
rect -2309 16436 -2301 16446
rect -2317 16430 -2309 16436
rect -2068 16435 -2038 16442
rect -2000 16434 -1992 16451
rect -1920 16450 -1906 16451
rect -1846 16444 -1794 16452
rect -1852 16437 -1804 16442
rect -1902 16435 -1804 16437
rect -1655 16436 -1647 16446
rect -2000 16432 -1975 16434
rect -1902 16433 -1852 16435
rect -2025 16430 -1975 16432
rect -1846 16430 -1804 16433
rect -1663 16430 -1655 16436
rect -1642 16430 -1637 16452
rect -1619 16430 -1614 16452
rect -1530 16430 -1526 16452
rect -1506 16430 -1502 16452
rect -1482 16430 -1478 16452
rect -1458 16430 -1454 16452
rect -1434 16430 -1430 16452
rect -1410 16430 -1406 16452
rect -1386 16430 -1382 16452
rect -1362 16430 -1358 16452
rect -1338 16430 -1334 16452
rect -1314 16430 -1310 16452
rect -1290 16430 -1286 16452
rect -1266 16430 -1262 16452
rect -1242 16430 -1238 16452
rect -1218 16430 -1214 16452
rect -1194 16430 -1190 16452
rect -1170 16430 -1166 16452
rect -1146 16430 -1142 16452
rect -1122 16430 -1118 16452
rect -1098 16430 -1094 16452
rect -1074 16430 -1070 16452
rect -1050 16430 -1046 16452
rect -1026 16430 -1022 16452
rect -1002 16430 -998 16452
rect -978 16430 -974 16452
rect -954 16430 -950 16452
rect -930 16430 -926 16452
rect -906 16430 -902 16452
rect -882 16430 -878 16452
rect -858 16430 -854 16452
rect -834 16430 -830 16452
rect -810 16430 -806 16452
rect -786 16430 -782 16452
rect -762 16430 -758 16452
rect -738 16430 -734 16452
rect -714 16430 -710 16452
rect -690 16430 -686 16452
rect -666 16430 -662 16452
rect -642 16430 -638 16452
rect -618 16430 -614 16452
rect -594 16430 -590 16452
rect -570 16430 -566 16452
rect -546 16430 -542 16452
rect -522 16430 -518 16452
rect -498 16430 -494 16452
rect -474 16430 -470 16452
rect -450 16430 -446 16452
rect -426 16451 -422 16452
rect -2393 16428 -429 16430
rect -2371 16406 -2366 16428
rect -2348 16406 -2343 16428
rect -2325 16406 -2320 16428
rect -2054 16427 -2038 16428
rect -2000 16427 -1966 16428
rect -1846 16427 -1804 16428
rect -2000 16426 -1975 16427
rect -2076 16418 -2054 16425
rect -2309 16408 -2301 16418
rect -2044 16415 -2038 16420
rect -2028 16418 -2001 16425
rect -2054 16408 -2038 16415
rect -2015 16417 -2001 16418
rect -2015 16408 -2014 16417
rect -2317 16406 -2309 16408
rect -2044 16406 -2028 16408
rect -2000 16406 -1992 16426
rect -1982 16425 -1975 16426
rect -1862 16425 -1798 16426
rect -1985 16418 -1796 16425
rect -1862 16417 -1798 16418
rect -1852 16408 -1804 16415
rect -1655 16408 -1647 16418
rect -1976 16406 -1940 16407
rect -1663 16406 -1655 16408
rect -1642 16406 -1637 16428
rect -1619 16406 -1614 16428
rect -1530 16406 -1526 16428
rect -1506 16406 -1502 16428
rect -1482 16406 -1478 16428
rect -1458 16406 -1454 16428
rect -1434 16406 -1430 16428
rect -1410 16406 -1406 16428
rect -1386 16406 -1382 16428
rect -1362 16406 -1358 16428
rect -1338 16406 -1334 16428
rect -1314 16406 -1310 16428
rect -1290 16406 -1286 16428
rect -1266 16406 -1262 16428
rect -1242 16406 -1238 16428
rect -1218 16406 -1214 16428
rect -1194 16406 -1190 16428
rect -1170 16406 -1166 16428
rect -1146 16406 -1142 16428
rect -1122 16406 -1118 16428
rect -1098 16406 -1094 16428
rect -1074 16406 -1070 16428
rect -1050 16406 -1046 16428
rect -1026 16406 -1022 16428
rect -1002 16406 -998 16428
rect -978 16427 -974 16428
rect -2393 16404 -981 16406
rect -2371 16334 -2366 16404
rect -2348 16334 -2343 16404
rect -2325 16370 -2320 16404
rect -2317 16402 -2309 16404
rect -2076 16391 -2054 16398
rect -2325 16362 -2317 16370
rect -2060 16364 -2030 16367
rect -2325 16342 -2320 16362
rect -2317 16354 -2309 16362
rect -2060 16351 -2038 16362
rect -2033 16355 -2030 16364
rect -2028 16360 -2027 16364
rect -2068 16346 -2038 16349
rect -2325 16334 -2317 16342
rect -2000 16334 -1992 16404
rect -1846 16400 -1804 16404
rect -1663 16402 -1655 16404
rect -1846 16390 -1794 16399
rect -1912 16379 -1884 16381
rect -1852 16373 -1804 16377
rect -1844 16364 -1796 16367
rect -1671 16362 -1663 16370
rect -1844 16351 -1804 16362
rect -1663 16354 -1655 16362
rect -1852 16346 -1680 16350
rect -1926 16334 -1892 16337
rect -1671 16334 -1663 16342
rect -1642 16334 -1637 16404
rect -1619 16334 -1614 16404
rect -1530 16334 -1526 16404
rect -1506 16334 -1502 16404
rect -1482 16334 -1478 16404
rect -1458 16334 -1454 16404
rect -1434 16334 -1430 16404
rect -1410 16334 -1406 16404
rect -1386 16334 -1382 16404
rect -1362 16334 -1358 16404
rect -1338 16334 -1334 16404
rect -1314 16334 -1310 16404
rect -1290 16334 -1286 16404
rect -1266 16334 -1262 16404
rect -1242 16334 -1238 16404
rect -1218 16334 -1214 16404
rect -1194 16334 -1190 16404
rect -1170 16334 -1166 16404
rect -1146 16334 -1142 16404
rect -1122 16334 -1118 16404
rect -1098 16334 -1094 16404
rect -1074 16334 -1070 16404
rect -1050 16334 -1046 16404
rect -1026 16334 -1022 16404
rect -1002 16334 -998 16404
rect -995 16403 -981 16404
rect -978 16382 -971 16427
rect -954 16382 -950 16428
rect -930 16382 -926 16428
rect -906 16382 -902 16428
rect -882 16382 -878 16428
rect -869 16397 -864 16407
rect -858 16397 -854 16428
rect -859 16383 -854 16397
rect -858 16382 -854 16383
rect -834 16382 -830 16428
rect -810 16382 -806 16428
rect -786 16382 -782 16428
rect -762 16382 -758 16428
rect -738 16382 -734 16428
rect -714 16382 -710 16428
rect -690 16382 -686 16428
rect -666 16382 -662 16428
rect -642 16382 -638 16428
rect -618 16382 -614 16428
rect -594 16382 -590 16428
rect -570 16382 -566 16428
rect -546 16382 -542 16428
rect -522 16382 -518 16428
rect -498 16382 -494 16428
rect -474 16382 -470 16428
rect -450 16382 -446 16428
rect -443 16427 -429 16428
rect -426 16403 -419 16451
rect -426 16382 -422 16403
rect -402 16382 -398 16452
rect -378 16382 -374 16452
rect -354 16382 -350 16452
rect -330 16382 -326 16452
rect -306 16382 -302 16452
rect -282 16382 -278 16452
rect -258 16382 -254 16452
rect -234 16382 -230 16452
rect -210 16382 -206 16452
rect -186 16382 -182 16452
rect -162 16382 -158 16452
rect -138 16382 -134 16452
rect -114 16382 -110 16452
rect -90 16382 -86 16452
rect -66 16382 -62 16452
rect -42 16382 -38 16452
rect -18 16382 -14 16452
rect 6 16382 10 16452
rect 30 16382 34 16452
rect 54 16382 58 16452
rect 78 16382 82 16452
rect 102 16382 106 16452
rect 126 16382 130 16452
rect 150 16382 154 16452
rect 174 16382 178 16452
rect 198 16382 202 16452
rect 222 16382 226 16452
rect 246 16382 250 16452
rect 270 16382 274 16452
rect 294 16382 298 16452
rect 318 16382 322 16452
rect 342 16382 346 16452
rect 366 16382 370 16452
rect 390 16382 394 16452
rect 414 16382 418 16452
rect 438 16382 442 16452
rect 462 16382 466 16452
rect 475 16421 480 16431
rect 486 16421 490 16452
rect 485 16407 490 16421
rect 486 16382 490 16407
rect 510 16382 514 16452
rect 534 16382 538 16452
rect 558 16382 562 16452
rect 582 16382 586 16452
rect 606 16382 610 16452
rect 630 16382 634 16452
rect 654 16382 658 16452
rect 678 16382 682 16452
rect 702 16382 706 16452
rect 726 16382 730 16452
rect 750 16382 754 16452
rect 774 16382 778 16452
rect 798 16382 802 16452
rect 822 16382 826 16452
rect 846 16382 850 16452
rect 870 16382 874 16452
rect 894 16382 898 16452
rect 918 16382 922 16452
rect 942 16382 946 16452
rect 966 16382 970 16452
rect 990 16382 994 16452
rect 1014 16382 1018 16452
rect 1038 16382 1042 16452
rect 1062 16382 1066 16452
rect 1086 16382 1090 16452
rect 1110 16382 1114 16452
rect 1134 16382 1138 16452
rect 1158 16382 1162 16452
rect 1182 16382 1186 16452
rect 1206 16382 1210 16452
rect 1230 16382 1234 16452
rect 1254 16382 1258 16452
rect 1278 16382 1282 16452
rect 1302 16382 1306 16452
rect 1326 16382 1330 16452
rect 1350 16382 1354 16452
rect 1374 16382 1378 16452
rect 1398 16382 1402 16452
rect 1422 16382 1426 16452
rect 1446 16382 1450 16452
rect 1470 16382 1474 16452
rect 1494 16382 1498 16452
rect 1518 16382 1522 16452
rect 1542 16382 1546 16452
rect 1566 16382 1570 16452
rect 1590 16382 1594 16452
rect 1614 16382 1618 16452
rect 1638 16382 1642 16452
rect 1662 16382 1666 16452
rect 1686 16382 1690 16452
rect 1710 16382 1714 16452
rect 1734 16382 1738 16452
rect 1758 16382 1762 16452
rect 1782 16382 1786 16452
rect 1806 16382 1810 16452
rect 1830 16382 1834 16452
rect 1854 16382 1858 16452
rect 1878 16382 1882 16452
rect 1902 16382 1906 16452
rect 1926 16382 1930 16452
rect 1950 16382 1954 16452
rect 1974 16382 1978 16452
rect 1998 16382 2002 16452
rect 2022 16382 2026 16452
rect 2046 16382 2050 16452
rect 2070 16382 2074 16452
rect 2094 16382 2098 16452
rect 2118 16382 2122 16452
rect 2142 16382 2146 16452
rect 2166 16382 2170 16452
rect 2190 16382 2194 16452
rect 2214 16382 2218 16452
rect 2238 16382 2242 16452
rect 2262 16382 2266 16452
rect 2286 16382 2290 16452
rect 2310 16382 2314 16452
rect 2334 16382 2338 16452
rect 2358 16382 2362 16452
rect 2382 16382 2386 16452
rect 2406 16382 2410 16452
rect 2430 16382 2434 16452
rect 2454 16382 2458 16452
rect 2478 16382 2482 16452
rect 2502 16382 2506 16452
rect 2526 16382 2530 16452
rect 2550 16382 2554 16452
rect 2574 16382 2578 16452
rect 2598 16382 2602 16452
rect 2622 16382 2626 16452
rect 2646 16382 2650 16452
rect 2670 16382 2674 16452
rect 2694 16382 2698 16452
rect 2718 16382 2722 16452
rect 2742 16382 2746 16452
rect 2766 16382 2770 16452
rect 2790 16382 2794 16452
rect 2814 16382 2818 16452
rect 2838 16382 2842 16452
rect 2862 16382 2866 16452
rect 2886 16382 2890 16452
rect 2910 16382 2914 16452
rect 2934 16382 2938 16452
rect 2958 16382 2962 16452
rect 2982 16382 2986 16452
rect 3006 16382 3010 16452
rect 3030 16382 3034 16452
rect 3054 16382 3058 16452
rect 3078 16382 3082 16452
rect 3102 16382 3106 16452
rect 3126 16382 3130 16452
rect 3150 16382 3154 16452
rect 3174 16382 3178 16452
rect 3198 16382 3202 16452
rect 3222 16382 3226 16452
rect 3246 16382 3250 16452
rect 3270 16383 3274 16452
rect 3259 16382 3293 16383
rect -995 16380 3293 16382
rect -995 16379 -981 16380
rect -978 16379 -971 16380
rect -978 16334 -974 16379
rect -954 16334 -950 16380
rect -930 16334 -926 16380
rect -906 16334 -902 16380
rect -882 16334 -878 16380
rect -858 16334 -854 16380
rect -834 16334 -830 16380
rect -810 16334 -806 16380
rect -786 16334 -782 16380
rect -762 16334 -758 16380
rect -738 16334 -734 16380
rect -714 16334 -710 16380
rect -690 16334 -686 16380
rect -666 16334 -662 16380
rect -642 16334 -638 16380
rect -618 16334 -614 16380
rect -594 16334 -590 16380
rect -570 16334 -566 16380
rect -546 16334 -542 16380
rect -522 16334 -518 16380
rect -498 16334 -494 16380
rect -474 16334 -470 16380
rect -450 16334 -446 16380
rect -426 16334 -422 16380
rect -402 16334 -398 16380
rect -378 16334 -374 16380
rect -354 16334 -350 16380
rect -330 16334 -326 16380
rect -306 16334 -302 16380
rect -282 16334 -278 16380
rect -258 16334 -254 16380
rect -234 16334 -230 16380
rect -210 16334 -206 16380
rect -186 16334 -182 16380
rect -162 16334 -158 16380
rect -138 16334 -134 16380
rect -114 16334 -110 16380
rect -90 16334 -86 16380
rect -66 16334 -62 16380
rect -42 16334 -38 16380
rect -18 16334 -14 16380
rect 6 16334 10 16380
rect 30 16334 34 16380
rect 54 16334 58 16380
rect 78 16334 82 16380
rect 102 16334 106 16380
rect 126 16334 130 16380
rect 150 16334 154 16380
rect 174 16334 178 16380
rect 198 16334 202 16380
rect 222 16334 226 16380
rect 246 16334 250 16380
rect 270 16334 274 16380
rect 294 16334 298 16380
rect 318 16334 322 16380
rect 342 16334 346 16380
rect 366 16334 370 16380
rect 390 16334 394 16380
rect 414 16334 418 16380
rect 438 16334 442 16380
rect 462 16334 466 16380
rect 486 16334 490 16380
rect 510 16355 514 16380
rect -2393 16332 507 16334
rect -2371 16310 -2366 16332
rect -2348 16310 -2343 16332
rect -2325 16326 -2317 16332
rect -2325 16310 -2320 16326
rect -2309 16314 -2301 16326
rect -2068 16315 -2038 16322
rect -2317 16310 -2309 16314
rect -2000 16312 -1992 16332
rect -1844 16324 -1794 16332
rect -1671 16326 -1663 16332
rect -1852 16315 -1804 16322
rect -1655 16314 -1647 16326
rect -2025 16311 -1991 16312
rect -2025 16310 -1975 16311
rect -1844 16310 -1804 16313
rect -1663 16310 -1655 16314
rect -1642 16310 -1637 16332
rect -1619 16310 -1614 16332
rect -1530 16310 -1526 16332
rect -1506 16310 -1502 16332
rect -1482 16310 -1478 16332
rect -1458 16310 -1454 16332
rect -1434 16310 -1430 16332
rect -1410 16310 -1406 16332
rect -1386 16310 -1382 16332
rect -1362 16310 -1358 16332
rect -1338 16310 -1334 16332
rect -1314 16310 -1310 16332
rect -1290 16310 -1286 16332
rect -1266 16310 -1262 16332
rect -1242 16310 -1238 16332
rect -1218 16310 -1214 16332
rect -1194 16310 -1190 16332
rect -1170 16310 -1166 16332
rect -1146 16310 -1142 16332
rect -1122 16310 -1118 16332
rect -1098 16310 -1094 16332
rect -1074 16310 -1070 16332
rect -1050 16310 -1046 16332
rect -1026 16310 -1022 16332
rect -1002 16310 -998 16332
rect -978 16310 -974 16332
rect -954 16310 -950 16332
rect -930 16310 -926 16332
rect -906 16310 -902 16332
rect -882 16310 -878 16332
rect -858 16310 -854 16332
rect -834 16331 -830 16332
rect -2393 16308 -837 16310
rect -2371 16286 -2366 16308
rect -2348 16286 -2343 16308
rect -2325 16298 -2317 16308
rect -2060 16298 -2020 16305
rect -2004 16300 -2001 16305
rect -2015 16298 -2001 16300
rect -2000 16298 -1992 16308
rect -1972 16306 -1958 16308
rect -1844 16307 -1804 16308
rect -1862 16305 -1796 16306
rect -1985 16303 -1796 16305
rect -1985 16298 -1852 16303
rect -2325 16286 -2320 16298
rect -2309 16286 -2301 16298
rect -2068 16288 -2060 16295
rect -2015 16288 -1990 16298
rect -1844 16297 -1796 16303
rect -1671 16298 -1663 16308
rect -1852 16288 -1804 16295
rect -2020 16286 -2004 16288
rect -2000 16286 -1992 16288
rect -1976 16286 -1940 16287
rect -1655 16286 -1647 16298
rect -1642 16286 -1637 16308
rect -1619 16286 -1614 16308
rect -1530 16286 -1526 16308
rect -1506 16286 -1502 16308
rect -1482 16286 -1478 16308
rect -1458 16286 -1454 16308
rect -1434 16286 -1430 16308
rect -1410 16286 -1406 16308
rect -1386 16286 -1382 16308
rect -1362 16286 -1358 16308
rect -1338 16286 -1334 16308
rect -1314 16286 -1310 16308
rect -1290 16286 -1286 16308
rect -1266 16286 -1262 16308
rect -1242 16286 -1238 16308
rect -1218 16286 -1214 16308
rect -1194 16286 -1190 16308
rect -1170 16286 -1166 16308
rect -1146 16286 -1142 16308
rect -1122 16286 -1118 16308
rect -1098 16286 -1094 16308
rect -1074 16286 -1070 16308
rect -1050 16286 -1046 16308
rect -1026 16286 -1022 16308
rect -1002 16286 -998 16308
rect -978 16286 -974 16308
rect -954 16286 -950 16308
rect -930 16286 -926 16308
rect -906 16286 -902 16308
rect -882 16286 -878 16308
rect -858 16286 -854 16308
rect -851 16307 -837 16308
rect -834 16307 -827 16331
rect -834 16286 -830 16307
rect -810 16286 -806 16332
rect -786 16286 -782 16332
rect -762 16286 -758 16332
rect -738 16286 -734 16332
rect -714 16286 -710 16332
rect -690 16286 -686 16332
rect -666 16286 -662 16332
rect -642 16286 -638 16332
rect -618 16286 -614 16332
rect -594 16286 -590 16332
rect -570 16286 -566 16332
rect -546 16286 -542 16332
rect -522 16286 -518 16332
rect -498 16286 -494 16332
rect -474 16286 -470 16332
rect -450 16286 -446 16332
rect -426 16286 -422 16332
rect -402 16286 -398 16332
rect -378 16286 -374 16332
rect -354 16286 -350 16332
rect -330 16286 -326 16332
rect -306 16286 -302 16332
rect -282 16286 -278 16332
rect -258 16286 -254 16332
rect -234 16286 -230 16332
rect -210 16286 -206 16332
rect -186 16286 -182 16332
rect -162 16286 -158 16332
rect -138 16286 -134 16332
rect -114 16286 -110 16332
rect -90 16286 -86 16332
rect -66 16286 -62 16332
rect -42 16286 -38 16332
rect -18 16286 -14 16332
rect 6 16286 10 16332
rect 30 16286 34 16332
rect 54 16286 58 16332
rect 78 16286 82 16332
rect 102 16286 106 16332
rect 126 16286 130 16332
rect 150 16286 154 16332
rect 174 16286 178 16332
rect 198 16286 202 16332
rect 222 16286 226 16332
rect 246 16286 250 16332
rect 270 16286 274 16332
rect 294 16286 298 16332
rect 318 16286 322 16332
rect 342 16286 346 16332
rect 366 16286 370 16332
rect 390 16286 394 16332
rect 414 16286 418 16332
rect 438 16286 442 16332
rect 462 16286 466 16332
rect 486 16286 490 16332
rect 493 16331 507 16332
rect 510 16331 517 16355
rect 510 16286 514 16331
rect 534 16286 538 16380
rect 558 16286 562 16380
rect 582 16286 586 16380
rect 606 16286 610 16380
rect 630 16286 634 16380
rect 654 16286 658 16380
rect 678 16286 682 16380
rect 702 16286 706 16380
rect 726 16286 730 16380
rect 750 16286 754 16380
rect 774 16286 778 16380
rect 798 16286 802 16380
rect 822 16286 826 16380
rect 846 16286 850 16380
rect 870 16286 874 16380
rect 894 16286 898 16380
rect 918 16286 922 16380
rect 931 16301 936 16311
rect 942 16301 946 16380
rect 941 16287 946 16301
rect 966 16286 970 16380
rect 990 16286 994 16380
rect 1014 16286 1018 16380
rect 1038 16286 1042 16380
rect 1062 16286 1066 16380
rect 1086 16286 1090 16380
rect 1110 16286 1114 16380
rect 1134 16286 1138 16380
rect 1158 16286 1162 16380
rect 1182 16286 1186 16380
rect 1206 16286 1210 16380
rect 1230 16286 1234 16380
rect 1254 16286 1258 16380
rect 1278 16286 1282 16380
rect 1302 16286 1306 16380
rect 1326 16286 1330 16380
rect 1350 16286 1354 16380
rect 1374 16286 1378 16380
rect 1398 16286 1402 16380
rect 1422 16286 1426 16380
rect 1446 16286 1450 16380
rect 1470 16286 1474 16380
rect 1494 16286 1498 16380
rect 1518 16286 1522 16380
rect 1542 16286 1546 16380
rect 1566 16286 1570 16380
rect 1590 16286 1594 16380
rect 1614 16286 1618 16380
rect 1638 16286 1642 16380
rect 1662 16286 1666 16380
rect 1686 16286 1690 16380
rect 1710 16286 1714 16380
rect 1734 16286 1738 16380
rect 1758 16286 1762 16380
rect 1782 16286 1786 16380
rect 1806 16286 1810 16380
rect 1830 16286 1834 16380
rect 1854 16286 1858 16380
rect 1878 16286 1882 16380
rect 1902 16286 1906 16380
rect 1926 16287 1930 16380
rect 1915 16286 1949 16287
rect -2393 16284 1949 16286
rect -2371 16214 -2366 16284
rect -2348 16214 -2343 16284
rect -2325 16282 -2320 16284
rect -2317 16282 -2309 16284
rect -2325 16270 -2317 16282
rect -2060 16271 -2030 16278
rect -2325 16250 -2320 16270
rect -2325 16242 -2317 16250
rect -2060 16244 -2030 16247
rect -2325 16214 -2320 16242
rect -2317 16234 -2309 16242
rect -2060 16231 -2038 16242
rect -2033 16235 -2030 16244
rect -2028 16240 -2027 16244
rect -2068 16226 -2038 16229
rect -2000 16214 -1992 16284
rect -1844 16280 -1804 16284
rect -1663 16282 -1655 16284
rect -1844 16270 -1794 16279
rect -1671 16270 -1663 16282
rect -1912 16259 -1884 16261
rect -1852 16253 -1804 16257
rect -1844 16244 -1796 16247
rect -1671 16242 -1663 16250
rect -1844 16231 -1804 16242
rect -1663 16234 -1655 16242
rect -1852 16226 -1680 16230
rect -1979 16214 -1945 16216
rect -1642 16214 -1637 16284
rect -1619 16214 -1614 16284
rect -1530 16214 -1526 16284
rect -1506 16214 -1502 16284
rect -1482 16214 -1478 16284
rect -1458 16214 -1454 16284
rect -1434 16214 -1430 16284
rect -1410 16214 -1406 16284
rect -1386 16214 -1382 16284
rect -1362 16214 -1358 16284
rect -1338 16214 -1334 16284
rect -1314 16214 -1310 16284
rect -1290 16214 -1286 16284
rect -1266 16214 -1262 16284
rect -1242 16214 -1238 16284
rect -1218 16214 -1214 16284
rect -1194 16214 -1190 16284
rect -1170 16214 -1166 16284
rect -1146 16214 -1142 16284
rect -1122 16214 -1118 16284
rect -1098 16214 -1094 16284
rect -1074 16214 -1070 16284
rect -1050 16214 -1046 16284
rect -1026 16214 -1022 16284
rect -1002 16214 -998 16284
rect -978 16214 -974 16284
rect -954 16214 -950 16284
rect -930 16214 -926 16284
rect -906 16214 -902 16284
rect -882 16214 -878 16284
rect -858 16214 -854 16284
rect -834 16214 -830 16284
rect -810 16214 -806 16284
rect -786 16214 -782 16284
rect -762 16214 -758 16284
rect -738 16214 -734 16284
rect -714 16214 -710 16284
rect -690 16214 -686 16284
rect -666 16214 -662 16284
rect -642 16214 -638 16284
rect -618 16214 -614 16284
rect -594 16214 -590 16284
rect -570 16214 -566 16284
rect -546 16214 -542 16284
rect -522 16214 -518 16284
rect -498 16214 -494 16284
rect -474 16214 -470 16284
rect -450 16214 -446 16284
rect -426 16214 -422 16284
rect -402 16214 -398 16284
rect -378 16214 -374 16284
rect -354 16214 -350 16284
rect -330 16214 -326 16284
rect -306 16214 -302 16284
rect -282 16214 -278 16284
rect -258 16214 -254 16284
rect -234 16214 -230 16284
rect -210 16214 -206 16284
rect -186 16214 -182 16284
rect -162 16214 -158 16284
rect -138 16214 -134 16284
rect -114 16214 -110 16284
rect -90 16214 -86 16284
rect -66 16214 -62 16284
rect -42 16214 -38 16284
rect -18 16214 -14 16284
rect 6 16214 10 16284
rect 30 16214 34 16284
rect 54 16214 58 16284
rect 78 16214 82 16284
rect 102 16214 106 16284
rect 126 16214 130 16284
rect 150 16214 154 16284
rect 174 16214 178 16284
rect 198 16214 202 16284
rect 222 16214 226 16284
rect 246 16214 250 16284
rect 270 16214 274 16284
rect 294 16214 298 16284
rect 318 16214 322 16284
rect 342 16214 346 16284
rect 366 16214 370 16284
rect 390 16214 394 16284
rect 414 16214 418 16284
rect 438 16214 442 16284
rect 462 16214 466 16284
rect 486 16214 490 16284
rect 510 16214 514 16284
rect 534 16214 538 16284
rect 558 16214 562 16284
rect 582 16214 586 16284
rect 606 16214 610 16284
rect 630 16214 634 16284
rect 654 16214 658 16284
rect 678 16214 682 16284
rect 702 16214 706 16284
rect 726 16214 730 16284
rect 750 16214 754 16284
rect 774 16214 778 16284
rect 798 16214 802 16284
rect 822 16214 826 16284
rect 846 16214 850 16284
rect 870 16214 874 16284
rect 894 16214 898 16284
rect 918 16214 922 16284
rect 931 16253 936 16263
rect 941 16239 946 16253
rect 942 16214 946 16239
rect 966 16235 970 16284
rect -2393 16212 963 16214
rect -2371 16166 -2366 16212
rect -2348 16166 -2343 16212
rect -2325 16166 -2320 16212
rect -2309 16194 -2301 16202
rect -2068 16195 -2040 16202
rect -2317 16186 -2309 16194
rect -2000 16185 -1992 16212
rect -1850 16204 -1844 16212
rect -1840 16204 -1792 16212
rect -1894 16202 -1850 16203
rect -1958 16200 -1955 16201
rect -1969 16194 -1955 16200
rect -1894 16195 -1802 16202
rect -1894 16194 -1850 16195
rect -1655 16194 -1647 16202
rect -1969 16192 -1942 16194
rect -1955 16185 -1942 16192
rect -1844 16187 -1802 16193
rect -1663 16186 -1655 16194
rect -1860 16185 -1796 16186
rect -2040 16178 -2020 16185
rect -2004 16178 -1945 16185
rect -1929 16183 -1794 16185
rect -1929 16178 -1850 16183
rect -1844 16178 -1794 16183
rect -2309 16166 -2301 16174
rect -2136 16166 -2129 16176
rect -2068 16168 -2040 16175
rect -2020 16166 -2004 16168
rect -2000 16166 -1992 16178
rect -1844 16177 -1796 16178
rect -1850 16168 -1802 16175
rect -1978 16166 -1942 16167
rect -1655 16166 -1647 16174
rect -1642 16166 -1637 16212
rect -1619 16166 -1614 16212
rect -1530 16166 -1526 16212
rect -1506 16166 -1502 16212
rect -1482 16166 -1478 16212
rect -1458 16166 -1454 16212
rect -1434 16166 -1430 16212
rect -1410 16166 -1406 16212
rect -1386 16166 -1382 16212
rect -1362 16166 -1358 16212
rect -1338 16166 -1334 16212
rect -1314 16166 -1310 16212
rect -1290 16166 -1286 16212
rect -1266 16166 -1262 16212
rect -1242 16166 -1238 16212
rect -1218 16166 -1214 16212
rect -1194 16166 -1190 16212
rect -1170 16166 -1166 16212
rect -1146 16166 -1142 16212
rect -1122 16166 -1118 16212
rect -1098 16166 -1094 16212
rect -1074 16166 -1070 16212
rect -1050 16166 -1046 16212
rect -1026 16166 -1022 16212
rect -1002 16166 -998 16212
rect -978 16166 -974 16212
rect -954 16166 -950 16212
rect -930 16166 -926 16212
rect -906 16166 -902 16212
rect -882 16166 -878 16212
rect -858 16166 -854 16212
rect -834 16166 -830 16212
rect -810 16166 -806 16212
rect -786 16166 -782 16212
rect -762 16166 -758 16212
rect -738 16166 -734 16212
rect -714 16166 -710 16212
rect -690 16166 -686 16212
rect -666 16166 -662 16212
rect -642 16166 -638 16212
rect -618 16166 -614 16212
rect -594 16166 -590 16212
rect -570 16166 -566 16212
rect -546 16166 -542 16212
rect -522 16166 -518 16212
rect -498 16166 -494 16212
rect -474 16166 -470 16212
rect -450 16166 -446 16212
rect -426 16166 -422 16212
rect -402 16166 -398 16212
rect -378 16166 -374 16212
rect -354 16166 -350 16212
rect -330 16166 -326 16212
rect -306 16166 -302 16212
rect -282 16166 -278 16212
rect -258 16166 -254 16212
rect -234 16166 -230 16212
rect -210 16166 -206 16212
rect -186 16166 -182 16212
rect -162 16166 -158 16212
rect -138 16166 -134 16212
rect -114 16166 -110 16212
rect -90 16166 -86 16212
rect -66 16166 -62 16212
rect -42 16166 -38 16212
rect -18 16166 -14 16212
rect 6 16166 10 16212
rect 30 16167 34 16212
rect 19 16166 53 16167
rect -2393 16164 53 16166
rect -2371 16070 -2366 16164
rect -2348 16070 -2343 16164
rect -2325 16126 -2320 16164
rect -2317 16158 -2309 16164
rect -2124 16160 -2117 16164
rect -2060 16160 -2040 16164
rect -2060 16151 -2030 16158
rect -2062 16126 -2032 16127
rect -2000 16126 -1992 16164
rect -1844 16160 -1802 16164
rect -1844 16150 -1792 16159
rect -1663 16158 -1655 16164
rect -1942 16128 -1937 16140
rect -1850 16137 -1822 16138
rect -1850 16133 -1802 16137
rect -2325 16118 -2317 16126
rect -2062 16124 -1961 16126
rect -2325 16098 -2320 16118
rect -2317 16110 -2309 16118
rect -2062 16111 -2040 16122
rect -2032 16117 -1961 16124
rect -1947 16118 -1942 16126
rect -1842 16124 -1794 16127
rect -2070 16106 -2022 16110
rect -2325 16086 -2317 16098
rect -2325 16070 -2320 16086
rect -2317 16082 -2309 16086
rect -2309 16070 -2301 16082
rect -2068 16075 -2038 16082
rect -2000 16072 -1992 16117
rect -1942 16116 -1937 16118
rect -1932 16108 -1927 16116
rect -1912 16113 -1896 16119
rect -1842 16111 -1802 16122
rect -1671 16118 -1663 16126
rect -1663 16110 -1655 16118
rect -1850 16106 -1680 16110
rect -1937 16092 -1934 16094
rect -1926 16092 -1921 16097
rect -1926 16087 -1924 16092
rect -1916 16084 -1914 16087
rect -1842 16084 -1794 16093
rect -1671 16086 -1663 16098
rect -1924 16074 -1916 16083
rect -1663 16082 -1655 16086
rect -1852 16075 -1804 16082
rect -1916 16073 -1914 16074
rect -2025 16071 -1991 16072
rect -2025 16070 -1975 16071
rect -1842 16070 -1804 16073
rect -1655 16070 -1647 16082
rect -1642 16070 -1637 16164
rect -1619 16070 -1614 16164
rect -1530 16070 -1526 16164
rect -1506 16070 -1502 16164
rect -1482 16070 -1478 16164
rect -1458 16070 -1454 16164
rect -1434 16070 -1430 16164
rect -1410 16070 -1406 16164
rect -1386 16070 -1382 16164
rect -1362 16070 -1358 16164
rect -1338 16070 -1334 16164
rect -1314 16070 -1310 16164
rect -1290 16070 -1286 16164
rect -1266 16070 -1262 16164
rect -1242 16071 -1238 16164
rect -1253 16070 -1219 16071
rect -2393 16068 -1219 16070
rect -2371 16046 -2366 16068
rect -2348 16046 -2343 16068
rect -2325 16058 -2317 16068
rect -2076 16058 -2068 16065
rect -2062 16058 -2001 16065
rect -2325 16046 -2320 16058
rect -2317 16054 -2309 16058
rect -2015 16057 -2001 16058
rect -2309 16046 -2301 16054
rect -2068 16048 -2062 16055
rect -2000 16050 -1992 16068
rect -1974 16066 -1960 16068
rect -1842 16067 -1804 16068
rect -1862 16065 -1794 16066
rect -1985 16063 -1794 16065
rect -1985 16058 -1852 16063
rect -1842 16057 -1794 16063
rect -1671 16058 -1663 16068
rect -2015 16048 -1985 16050
rect -1852 16048 -1804 16055
rect -1663 16054 -1655 16058
rect -2000 16046 -1992 16048
rect -1976 16046 -1940 16047
rect -1655 16046 -1647 16054
rect -1642 16046 -1637 16068
rect -1619 16046 -1614 16068
rect -1530 16047 -1526 16068
rect -1541 16046 -1507 16047
rect -2393 16044 -1507 16046
rect -2371 15974 -2366 16044
rect -2348 15974 -2343 16044
rect -2325 16042 -2320 16044
rect -2309 16042 -2301 16044
rect -2325 16030 -2317 16042
rect -2062 16031 -2032 16038
rect -2325 16010 -2320 16030
rect -2317 16026 -2309 16030
rect -2325 16002 -2317 16010
rect -2060 16004 -2030 16007
rect -2325 15974 -2320 16002
rect -2317 15994 -2309 16002
rect -2060 15991 -2038 16002
rect -2033 15995 -2030 16004
rect -2028 16000 -2027 16004
rect -2068 15986 -2038 15989
rect -2000 15974 -1992 16044
rect -1888 16039 -1874 16044
rect -1842 16040 -1804 16044
rect -1655 16042 -1647 16044
rect -1902 16037 -1874 16039
rect -1842 16030 -1794 16039
rect -1671 16030 -1663 16042
rect -1663 16026 -1655 16030
rect -1912 16019 -1884 16021
rect -1852 16013 -1804 16017
rect -1844 16004 -1796 16007
rect -1671 16002 -1663 16010
rect -1844 15991 -1804 16002
rect -1663 15994 -1655 16002
rect -1852 15986 -1680 15990
rect -1979 15974 -1945 15976
rect -1642 15974 -1637 16044
rect -1619 15974 -1614 16044
rect -1541 16037 -1536 16044
rect -1530 16037 -1526 16044
rect -1531 16023 -1526 16037
rect -1530 15974 -1526 16023
rect -1506 15974 -1502 16068
rect -1482 15974 -1478 16068
rect -1458 15974 -1454 16068
rect -1434 15974 -1430 16068
rect -1410 15974 -1406 16068
rect -1386 15974 -1382 16068
rect -1362 15974 -1358 16068
rect -1338 15974 -1334 16068
rect -1314 15974 -1310 16068
rect -1290 15974 -1286 16068
rect -1266 15974 -1262 16068
rect -1253 16061 -1248 16068
rect -1242 16061 -1238 16068
rect -1243 16047 -1238 16061
rect -1253 16046 -1219 16047
rect -1218 16046 -1214 16164
rect -1194 16046 -1190 16164
rect -1170 16046 -1166 16164
rect -1146 16046 -1142 16164
rect -1122 16046 -1118 16164
rect -1098 16046 -1094 16164
rect -1074 16046 -1070 16164
rect -1050 16046 -1046 16164
rect -1026 16046 -1022 16164
rect -1002 16046 -998 16164
rect -978 16046 -974 16164
rect -954 16046 -950 16164
rect -930 16046 -926 16164
rect -906 16046 -902 16164
rect -882 16046 -878 16164
rect -858 16046 -854 16164
rect -834 16046 -830 16164
rect -810 16046 -806 16164
rect -786 16046 -782 16164
rect -762 16046 -758 16164
rect -738 16046 -734 16164
rect -714 16046 -710 16164
rect -690 16046 -686 16164
rect -666 16046 -662 16164
rect -642 16046 -638 16164
rect -618 16046 -614 16164
rect -594 16046 -590 16164
rect -570 16046 -566 16164
rect -546 16046 -542 16164
rect -522 16046 -518 16164
rect -498 16046 -494 16164
rect -474 16046 -470 16164
rect -450 16046 -446 16164
rect -426 16046 -422 16164
rect -402 16046 -398 16164
rect -378 16046 -374 16164
rect -354 16046 -350 16164
rect -330 16046 -326 16164
rect -306 16046 -302 16164
rect -282 16046 -278 16164
rect -258 16046 -254 16164
rect -234 16046 -230 16164
rect -210 16046 -206 16164
rect -186 16046 -182 16164
rect -162 16046 -158 16164
rect -138 16046 -134 16164
rect -114 16046 -110 16164
rect -90 16046 -86 16164
rect -66 16046 -62 16164
rect -42 16046 -38 16164
rect -18 16046 -14 16164
rect 6 16046 10 16164
rect 19 16157 24 16164
rect 30 16157 34 16164
rect 29 16143 34 16157
rect 19 16118 53 16119
rect 54 16118 58 16212
rect 78 16118 82 16212
rect 102 16118 106 16212
rect 126 16118 130 16212
rect 150 16118 154 16212
rect 174 16118 178 16212
rect 198 16118 202 16212
rect 222 16118 226 16212
rect 246 16118 250 16212
rect 270 16118 274 16212
rect 294 16118 298 16212
rect 318 16118 322 16212
rect 342 16118 346 16212
rect 366 16118 370 16212
rect 390 16118 394 16212
rect 414 16118 418 16212
rect 438 16118 442 16212
rect 462 16118 466 16212
rect 486 16118 490 16212
rect 510 16118 514 16212
rect 534 16118 538 16212
rect 558 16118 562 16212
rect 582 16118 586 16212
rect 606 16118 610 16212
rect 630 16118 634 16212
rect 654 16118 658 16212
rect 678 16118 682 16212
rect 702 16118 706 16212
rect 726 16118 730 16212
rect 750 16118 754 16212
rect 774 16118 778 16212
rect 798 16118 802 16212
rect 822 16118 826 16212
rect 846 16118 850 16212
rect 870 16118 874 16212
rect 894 16118 898 16212
rect 918 16118 922 16212
rect 942 16118 946 16212
rect 949 16211 963 16212
rect 966 16211 973 16235
rect 966 16163 973 16187
rect 966 16118 970 16163
rect 990 16118 994 16284
rect 1014 16118 1018 16284
rect 1038 16118 1042 16284
rect 1062 16118 1066 16284
rect 1086 16118 1090 16284
rect 1110 16118 1114 16284
rect 1134 16118 1138 16284
rect 1158 16118 1162 16284
rect 1182 16118 1186 16284
rect 1206 16118 1210 16284
rect 1230 16118 1234 16284
rect 1254 16118 1258 16284
rect 1278 16118 1282 16284
rect 1302 16118 1306 16284
rect 1326 16118 1330 16284
rect 1350 16118 1354 16284
rect 1374 16118 1378 16284
rect 1398 16118 1402 16284
rect 1422 16118 1426 16284
rect 1446 16118 1450 16284
rect 1470 16118 1474 16284
rect 1494 16118 1498 16284
rect 1518 16118 1522 16284
rect 1542 16118 1546 16284
rect 1566 16118 1570 16284
rect 1590 16118 1594 16284
rect 1614 16118 1618 16284
rect 1638 16118 1642 16284
rect 1662 16118 1666 16284
rect 1686 16118 1690 16284
rect 1710 16118 1714 16284
rect 1734 16118 1738 16284
rect 1758 16118 1762 16284
rect 1782 16118 1786 16284
rect 1806 16118 1810 16284
rect 1830 16118 1834 16284
rect 1854 16118 1858 16284
rect 1878 16118 1882 16284
rect 1902 16118 1906 16284
rect 1915 16277 1920 16284
rect 1926 16277 1930 16284
rect 1925 16263 1930 16277
rect 1915 16238 1949 16239
rect 1950 16238 1954 16380
rect 1974 16238 1978 16380
rect 1998 16238 2002 16380
rect 2022 16238 2026 16380
rect 2046 16238 2050 16380
rect 2070 16238 2074 16380
rect 2094 16238 2098 16380
rect 2118 16238 2122 16380
rect 2142 16238 2146 16380
rect 2166 16238 2170 16380
rect 2190 16238 2194 16380
rect 2214 16238 2218 16380
rect 2238 16238 2242 16380
rect 2262 16238 2266 16380
rect 2286 16238 2290 16380
rect 2310 16238 2314 16380
rect 2334 16238 2338 16380
rect 2358 16238 2362 16380
rect 2382 16238 2386 16380
rect 2406 16238 2410 16380
rect 2430 16238 2434 16380
rect 2454 16238 2458 16380
rect 2478 16238 2482 16380
rect 2502 16238 2506 16380
rect 2526 16238 2530 16380
rect 2550 16238 2554 16380
rect 2574 16238 2578 16380
rect 2598 16238 2602 16380
rect 2622 16238 2626 16380
rect 2646 16238 2650 16380
rect 2670 16238 2674 16380
rect 2694 16238 2698 16380
rect 2718 16238 2722 16380
rect 2742 16238 2746 16380
rect 2766 16238 2770 16380
rect 2790 16238 2794 16380
rect 2814 16238 2818 16380
rect 2838 16238 2842 16380
rect 2862 16238 2866 16380
rect 2886 16238 2890 16380
rect 2910 16238 2914 16380
rect 2923 16253 2928 16263
rect 2934 16253 2938 16380
rect 2933 16239 2938 16253
rect 2958 16238 2962 16380
rect 2982 16238 2986 16380
rect 3006 16238 3010 16380
rect 3030 16238 3034 16380
rect 3054 16238 3058 16380
rect 3078 16238 3082 16380
rect 3102 16238 3106 16380
rect 3126 16238 3130 16380
rect 3150 16238 3154 16380
rect 3174 16238 3178 16380
rect 3198 16238 3202 16380
rect 3222 16238 3226 16380
rect 3246 16238 3250 16380
rect 3259 16373 3264 16380
rect 3270 16373 3274 16380
rect 3269 16359 3274 16373
rect 3270 16238 3274 16359
rect 3294 16307 3298 16452
rect 3294 16283 3301 16307
rect 3294 16238 3298 16283
rect 3318 16238 3322 16452
rect 3342 16238 3346 16452
rect 3366 16238 3370 16452
rect 3390 16238 3394 16452
rect 3414 16238 3418 16452
rect 3438 16238 3442 16452
rect 3462 16238 3466 16452
rect 3486 16238 3490 16452
rect 3510 16238 3514 16452
rect 3534 16238 3538 16452
rect 3558 16238 3562 16452
rect 3582 16238 3586 16452
rect 3606 16238 3610 16452
rect 3630 16238 3634 16452
rect 3654 16238 3658 16452
rect 3678 16238 3682 16452
rect 3702 16238 3706 16452
rect 3715 16445 3720 16452
rect 3725 16431 3730 16445
rect 3726 16238 3730 16431
rect 3739 16325 3744 16335
rect 3749 16311 3754 16325
rect 3750 16239 3754 16311
rect 3739 16238 3771 16239
rect 1915 16236 3771 16238
rect 1915 16229 1920 16236
rect 1925 16215 1930 16229
rect 1926 16118 1930 16215
rect 1950 16211 1954 16236
rect 1950 16187 1957 16211
rect 1950 16142 1957 16163
rect 1974 16142 1978 16236
rect 1998 16143 2002 16236
rect 1987 16142 2021 16143
rect 1933 16140 2021 16142
rect 1933 16139 1947 16140
rect 1950 16139 1957 16140
rect 1950 16118 1954 16139
rect 1974 16118 1978 16140
rect 1987 16133 1992 16140
rect 1998 16133 2002 16140
rect 1997 16119 2002 16133
rect 2022 16118 2026 16236
rect 2046 16118 2050 16236
rect 2070 16118 2074 16236
rect 2094 16118 2098 16236
rect 2118 16118 2122 16236
rect 2142 16118 2146 16236
rect 2166 16118 2170 16236
rect 2190 16118 2194 16236
rect 2214 16118 2218 16236
rect 2238 16118 2242 16236
rect 2262 16118 2266 16236
rect 2286 16118 2290 16236
rect 2310 16118 2314 16236
rect 2334 16118 2338 16236
rect 2358 16118 2362 16236
rect 2382 16118 2386 16236
rect 2406 16118 2410 16236
rect 2430 16118 2434 16236
rect 2454 16118 2458 16236
rect 2478 16118 2482 16236
rect 2502 16118 2506 16236
rect 2526 16118 2530 16236
rect 2550 16118 2554 16236
rect 2574 16118 2578 16236
rect 2598 16118 2602 16236
rect 2622 16118 2626 16236
rect 2646 16118 2650 16236
rect 2670 16118 2674 16236
rect 2694 16118 2698 16236
rect 2718 16118 2722 16236
rect 2742 16118 2746 16236
rect 2766 16118 2770 16236
rect 2790 16118 2794 16236
rect 2814 16118 2818 16236
rect 2838 16118 2842 16236
rect 2862 16118 2866 16236
rect 2886 16118 2890 16236
rect 2910 16118 2914 16236
rect 2923 16205 2928 16215
rect 2933 16191 2938 16205
rect 2934 16118 2938 16191
rect 2958 16187 2962 16236
rect 2958 16163 2965 16187
rect 19 16116 2955 16118
rect 19 16109 24 16116
rect 29 16095 34 16109
rect 30 16046 34 16095
rect 54 16091 58 16116
rect 54 16067 61 16091
rect 78 16046 82 16116
rect 102 16046 106 16116
rect 126 16046 130 16116
rect 150 16046 154 16116
rect 174 16046 178 16116
rect 198 16046 202 16116
rect 222 16046 226 16116
rect 246 16046 250 16116
rect 270 16046 274 16116
rect 294 16046 298 16116
rect 318 16046 322 16116
rect 342 16046 346 16116
rect 366 16046 370 16116
rect 390 16046 394 16116
rect 414 16046 418 16116
rect 438 16046 442 16116
rect 462 16046 466 16116
rect 486 16046 490 16116
rect 510 16046 514 16116
rect 534 16046 538 16116
rect 558 16046 562 16116
rect 582 16046 586 16116
rect 606 16046 610 16116
rect 630 16046 634 16116
rect 654 16046 658 16116
rect 678 16046 682 16116
rect 702 16046 706 16116
rect 726 16046 730 16116
rect 750 16046 754 16116
rect 774 16046 778 16116
rect 798 16046 802 16116
rect 822 16046 826 16116
rect 846 16046 850 16116
rect 870 16046 874 16116
rect 894 16046 898 16116
rect 918 16046 922 16116
rect 942 16046 946 16116
rect 966 16046 970 16116
rect 990 16046 994 16116
rect 1014 16046 1018 16116
rect 1038 16046 1042 16116
rect 1062 16046 1066 16116
rect 1086 16046 1090 16116
rect 1110 16046 1114 16116
rect 1134 16046 1138 16116
rect 1158 16046 1162 16116
rect 1182 16046 1186 16116
rect 1206 16046 1210 16116
rect 1230 16046 1234 16116
rect 1254 16046 1258 16116
rect 1278 16046 1282 16116
rect 1302 16046 1306 16116
rect 1326 16046 1330 16116
rect 1350 16046 1354 16116
rect 1374 16046 1378 16116
rect 1398 16046 1402 16116
rect 1422 16046 1426 16116
rect 1446 16046 1450 16116
rect 1470 16046 1474 16116
rect 1494 16046 1498 16116
rect 1518 16046 1522 16116
rect 1542 16046 1546 16116
rect 1566 16046 1570 16116
rect 1590 16046 1594 16116
rect 1614 16046 1618 16116
rect 1638 16046 1642 16116
rect 1662 16046 1666 16116
rect 1686 16046 1690 16116
rect 1710 16046 1714 16116
rect 1734 16046 1738 16116
rect 1758 16046 1762 16116
rect 1782 16046 1786 16116
rect 1806 16046 1810 16116
rect 1830 16046 1834 16116
rect 1854 16046 1858 16116
rect 1878 16046 1882 16116
rect 1902 16046 1906 16116
rect 1926 16046 1930 16116
rect 1950 16046 1954 16116
rect 1974 16046 1978 16116
rect 1987 16085 1992 16095
rect 1997 16071 2002 16085
rect 1998 16046 2002 16071
rect 2022 16067 2026 16116
rect -1253 16044 2019 16046
rect -1253 16037 -1248 16044
rect -1243 16023 -1238 16037
rect -1242 15974 -1238 16023
rect -1218 15995 -1214 16044
rect -2393 15972 -1221 15974
rect -2371 15926 -2366 15972
rect -2348 15926 -2343 15972
rect -2325 15926 -2320 15972
rect -2309 15954 -2301 15962
rect -2068 15955 -2040 15962
rect -2317 15946 -2309 15954
rect -2000 15945 -1992 15972
rect -1850 15964 -1844 15972
rect -1840 15964 -1792 15972
rect -1894 15962 -1850 15963
rect -1958 15960 -1955 15961
rect -1969 15954 -1955 15960
rect -1894 15955 -1802 15962
rect -1894 15954 -1850 15955
rect -1655 15954 -1647 15962
rect -1969 15952 -1942 15954
rect -1955 15945 -1942 15952
rect -1844 15947 -1802 15953
rect -1663 15946 -1655 15954
rect -1860 15945 -1796 15946
rect -2040 15938 -2020 15945
rect -2004 15938 -1945 15945
rect -1929 15943 -1794 15945
rect -1929 15938 -1850 15943
rect -1844 15938 -1794 15943
rect -2309 15926 -2301 15934
rect -2136 15926 -2129 15936
rect -2068 15928 -2040 15935
rect -2020 15926 -2004 15928
rect -2000 15926 -1992 15938
rect -1844 15937 -1796 15938
rect -1850 15928 -1802 15935
rect -1978 15926 -1942 15927
rect -1655 15926 -1647 15934
rect -1642 15926 -1637 15972
rect -1619 15926 -1614 15972
rect -1530 15926 -1526 15972
rect -1506 15971 -1502 15972
rect -1506 15947 -1499 15971
rect -1506 15926 -1502 15947
rect -1482 15926 -1478 15972
rect -1458 15926 -1454 15972
rect -1434 15926 -1430 15972
rect -1410 15926 -1406 15972
rect -1386 15926 -1382 15972
rect -1362 15926 -1358 15972
rect -1338 15926 -1334 15972
rect -1314 15926 -1310 15972
rect -1290 15926 -1286 15972
rect -1266 15926 -1262 15972
rect -1242 15926 -1238 15972
rect -1235 15971 -1221 15972
rect -1218 15947 -1211 15995
rect -1218 15926 -1214 15947
rect -1194 15926 -1190 16044
rect -1170 15926 -1166 16044
rect -1146 15926 -1142 16044
rect -1122 15926 -1118 16044
rect -1098 15926 -1094 16044
rect -1074 15926 -1070 16044
rect -1050 15926 -1046 16044
rect -1026 15926 -1022 16044
rect -1002 15926 -998 16044
rect -978 15926 -974 16044
rect -954 15926 -950 16044
rect -930 15926 -926 16044
rect -906 15926 -902 16044
rect -882 15926 -878 16044
rect -858 15926 -854 16044
rect -834 15926 -830 16044
rect -810 15926 -806 16044
rect -786 15926 -782 16044
rect -762 15926 -758 16044
rect -738 15926 -734 16044
rect -714 15926 -710 16044
rect -690 15926 -686 16044
rect -666 15926 -662 16044
rect -642 15926 -638 16044
rect -618 15926 -614 16044
rect -594 15926 -590 16044
rect -570 15926 -566 16044
rect -546 15926 -542 16044
rect -522 15926 -518 16044
rect -498 15926 -494 16044
rect -474 15926 -470 16044
rect -450 15926 -446 16044
rect -426 15926 -422 16044
rect -402 15926 -398 16044
rect -378 15926 -374 16044
rect -354 15926 -350 16044
rect -330 15926 -326 16044
rect -306 15926 -302 16044
rect -282 15926 -278 16044
rect -258 15926 -254 16044
rect -234 15926 -230 16044
rect -210 15926 -206 16044
rect -186 15926 -182 16044
rect -162 15926 -158 16044
rect -138 15926 -134 16044
rect -114 15926 -110 16044
rect -90 15926 -86 16044
rect -66 15926 -62 16044
rect -42 15926 -38 16044
rect -18 15926 -14 16044
rect 6 15926 10 16044
rect 30 15926 34 16044
rect 54 16022 61 16043
rect 78 16022 82 16044
rect 102 16022 106 16044
rect 126 16022 130 16044
rect 150 16022 154 16044
rect 174 16022 178 16044
rect 198 16022 202 16044
rect 222 16022 226 16044
rect 246 16022 250 16044
rect 270 16022 274 16044
rect 294 16022 298 16044
rect 318 16022 322 16044
rect 342 16022 346 16044
rect 366 16022 370 16044
rect 390 16022 394 16044
rect 414 16022 418 16044
rect 438 16022 442 16044
rect 462 16022 466 16044
rect 486 16022 490 16044
rect 510 16022 514 16044
rect 534 16022 538 16044
rect 558 16022 562 16044
rect 582 16022 586 16044
rect 606 16022 610 16044
rect 630 16022 634 16044
rect 654 16022 658 16044
rect 678 16022 682 16044
rect 702 16022 706 16044
rect 726 16022 730 16044
rect 750 16022 754 16044
rect 774 16022 778 16044
rect 798 16022 802 16044
rect 822 16022 826 16044
rect 846 16022 850 16044
rect 870 16022 874 16044
rect 894 16022 898 16044
rect 918 16022 922 16044
rect 942 16022 946 16044
rect 966 16022 970 16044
rect 990 16022 994 16044
rect 1014 16022 1018 16044
rect 1038 16022 1042 16044
rect 1062 16022 1066 16044
rect 1086 16022 1090 16044
rect 1110 16022 1114 16044
rect 1134 16022 1138 16044
rect 1158 16022 1162 16044
rect 1182 16022 1186 16044
rect 1206 16022 1210 16044
rect 1230 16022 1234 16044
rect 1254 16022 1258 16044
rect 1278 16022 1282 16044
rect 1302 16022 1306 16044
rect 1326 16022 1330 16044
rect 1350 16022 1354 16044
rect 1374 16022 1378 16044
rect 1398 16022 1402 16044
rect 1422 16022 1426 16044
rect 1446 16022 1450 16044
rect 1470 16022 1474 16044
rect 1494 16022 1498 16044
rect 1518 16022 1522 16044
rect 1542 16022 1546 16044
rect 1566 16022 1570 16044
rect 1590 16022 1594 16044
rect 1614 16022 1618 16044
rect 1638 16022 1642 16044
rect 1662 16022 1666 16044
rect 1686 16022 1690 16044
rect 1710 16022 1714 16044
rect 1734 16022 1738 16044
rect 1758 16022 1762 16044
rect 1782 16022 1786 16044
rect 1806 16022 1810 16044
rect 1830 16022 1834 16044
rect 1854 16022 1858 16044
rect 1878 16022 1882 16044
rect 1902 16022 1906 16044
rect 1926 16022 1930 16044
rect 1950 16022 1954 16044
rect 1974 16022 1978 16044
rect 1998 16022 2002 16044
rect 2005 16043 2019 16044
rect 2022 16043 2029 16067
rect 2046 16022 2050 16116
rect 2070 16022 2074 16116
rect 2094 16022 2098 16116
rect 2118 16022 2122 16116
rect 2142 16022 2146 16116
rect 2166 16022 2170 16116
rect 2190 16022 2194 16116
rect 2214 16022 2218 16116
rect 2238 16022 2242 16116
rect 2262 16022 2266 16116
rect 2286 16022 2290 16116
rect 2310 16022 2314 16116
rect 2334 16022 2338 16116
rect 2358 16022 2362 16116
rect 2382 16022 2386 16116
rect 2406 16022 2410 16116
rect 2430 16022 2434 16116
rect 2454 16022 2458 16116
rect 2478 16022 2482 16116
rect 2502 16022 2506 16116
rect 2526 16022 2530 16116
rect 2550 16022 2554 16116
rect 2574 16022 2578 16116
rect 2598 16022 2602 16116
rect 2622 16022 2626 16116
rect 2646 16022 2650 16116
rect 2670 16022 2674 16116
rect 2694 16022 2698 16116
rect 2718 16022 2722 16116
rect 2742 16022 2746 16116
rect 2766 16022 2770 16116
rect 2790 16022 2794 16116
rect 2814 16022 2818 16116
rect 2838 16022 2842 16116
rect 2862 16022 2866 16116
rect 2886 16022 2890 16116
rect 2910 16022 2914 16116
rect 2934 16022 2938 16116
rect 2941 16115 2955 16116
rect 2958 16115 2965 16139
rect 2958 16022 2962 16115
rect 2982 16022 2986 16236
rect 3006 16022 3010 16236
rect 3030 16022 3034 16236
rect 3054 16022 3058 16236
rect 3078 16022 3082 16236
rect 3102 16022 3106 16236
rect 3126 16022 3130 16236
rect 3150 16022 3154 16236
rect 3174 16023 3178 16236
rect 3163 16022 3197 16023
rect 37 16020 3197 16022
rect 37 16019 51 16020
rect 54 16019 61 16020
rect 54 15926 58 16019
rect 78 15926 82 16020
rect 102 15926 106 16020
rect 126 15926 130 16020
rect 150 15926 154 16020
rect 174 15926 178 16020
rect 198 15926 202 16020
rect 222 15926 226 16020
rect 246 15926 250 16020
rect 270 15926 274 16020
rect 294 15926 298 16020
rect 318 15926 322 16020
rect 342 15926 346 16020
rect 366 15926 370 16020
rect 390 15926 394 16020
rect 414 15926 418 16020
rect 438 15926 442 16020
rect 462 15926 466 16020
rect 486 15926 490 16020
rect 510 15926 514 16020
rect 534 15926 538 16020
rect 558 15926 562 16020
rect 582 15926 586 16020
rect 606 15926 610 16020
rect 630 15926 634 16020
rect 654 15926 658 16020
rect 678 15926 682 16020
rect 702 15926 706 16020
rect 726 15926 730 16020
rect 750 15926 754 16020
rect 774 15926 778 16020
rect 798 15926 802 16020
rect 822 15926 826 16020
rect 846 15926 850 16020
rect 870 15926 874 16020
rect 894 15926 898 16020
rect 918 15926 922 16020
rect 942 15926 946 16020
rect 966 15926 970 16020
rect 990 15926 994 16020
rect 1014 15926 1018 16020
rect 1038 15926 1042 16020
rect 1062 15926 1066 16020
rect 1086 15926 1090 16020
rect 1110 15926 1114 16020
rect 1134 15926 1138 16020
rect 1158 15926 1162 16020
rect 1182 15926 1186 16020
rect 1206 15926 1210 16020
rect 1230 15926 1234 16020
rect 1254 15926 1258 16020
rect 1278 15926 1282 16020
rect 1302 15926 1306 16020
rect 1326 15926 1330 16020
rect 1350 15926 1354 16020
rect 1374 15926 1378 16020
rect 1398 15926 1402 16020
rect 1422 15926 1426 16020
rect 1446 15926 1450 16020
rect 1470 15926 1474 16020
rect 1494 15926 1498 16020
rect 1518 15926 1522 16020
rect 1542 15926 1546 16020
rect 1566 15926 1570 16020
rect 1590 15926 1594 16020
rect 1614 15926 1618 16020
rect 1638 15926 1642 16020
rect 1662 15926 1666 16020
rect 1686 15926 1690 16020
rect 1710 15926 1714 16020
rect 1734 15926 1738 16020
rect 1758 15926 1762 16020
rect 1782 15926 1786 16020
rect 1806 15926 1810 16020
rect 1830 15926 1834 16020
rect 1854 15926 1858 16020
rect 1878 15926 1882 16020
rect 1902 15926 1906 16020
rect 1926 15926 1930 16020
rect 1950 15926 1954 16020
rect 1974 15926 1978 16020
rect 1998 15926 2002 16020
rect 2022 15995 2029 16019
rect 2022 15926 2026 15995
rect 2046 15926 2050 16020
rect 2070 15927 2074 16020
rect 2059 15926 2093 15927
rect -2393 15924 2093 15926
rect -2371 15830 -2366 15924
rect -2348 15830 -2343 15924
rect -2325 15886 -2320 15924
rect -2317 15918 -2309 15924
rect -2124 15920 -2117 15924
rect -2060 15920 -2040 15924
rect -2060 15911 -2030 15918
rect -2062 15886 -2032 15887
rect -2000 15886 -1992 15924
rect -1844 15920 -1802 15924
rect -1844 15910 -1792 15919
rect -1663 15918 -1655 15924
rect -1942 15888 -1937 15900
rect -1850 15897 -1822 15898
rect -1850 15893 -1802 15897
rect -2325 15878 -2317 15886
rect -2062 15884 -1961 15886
rect -2325 15858 -2320 15878
rect -2317 15870 -2309 15878
rect -2062 15871 -2040 15882
rect -2032 15877 -1961 15884
rect -1947 15878 -1942 15886
rect -1842 15884 -1794 15887
rect -2070 15866 -2022 15870
rect -2325 15844 -2317 15858
rect -2072 15850 -2032 15851
rect -2102 15844 -2032 15850
rect -2325 15830 -2320 15844
rect -2317 15842 -2309 15844
rect -2309 15830 -2301 15842
rect -2070 15835 -2062 15840
rect -2000 15830 -1992 15877
rect -1942 15876 -1937 15878
rect -1932 15868 -1927 15876
rect -1912 15873 -1896 15879
rect -1842 15871 -1802 15882
rect -1671 15878 -1663 15886
rect -1663 15870 -1655 15878
rect -1850 15866 -1680 15870
rect -1924 15852 -1921 15854
rect -1806 15844 -1680 15850
rect -1671 15844 -1663 15858
rect -1663 15842 -1655 15844
rect -1854 15835 -1806 15840
rect -1974 15830 -1964 15831
rect -1960 15830 -1944 15832
rect -1842 15830 -1806 15833
rect -1655 15830 -1647 15842
rect -1642 15830 -1637 15924
rect -1619 15830 -1614 15924
rect -1530 15830 -1526 15924
rect -1506 15830 -1502 15924
rect -1482 15830 -1478 15924
rect -1458 15830 -1454 15924
rect -1434 15830 -1430 15924
rect -1410 15830 -1406 15924
rect -1386 15830 -1382 15924
rect -1362 15830 -1358 15924
rect -1338 15830 -1334 15924
rect -1314 15830 -1310 15924
rect -1290 15830 -1286 15924
rect -1266 15830 -1262 15924
rect -1242 15830 -1238 15924
rect -1218 15830 -1214 15924
rect -1194 15830 -1190 15924
rect -1170 15830 -1166 15924
rect -1146 15830 -1142 15924
rect -1122 15830 -1118 15924
rect -1098 15830 -1094 15924
rect -1074 15830 -1070 15924
rect -1050 15830 -1046 15924
rect -1026 15830 -1022 15924
rect -1002 15830 -998 15924
rect -978 15830 -974 15924
rect -954 15830 -950 15924
rect -930 15830 -926 15924
rect -906 15830 -902 15924
rect -882 15830 -878 15924
rect -858 15830 -854 15924
rect -834 15830 -830 15924
rect -810 15830 -806 15924
rect -786 15830 -782 15924
rect -762 15830 -758 15924
rect -738 15830 -734 15924
rect -714 15830 -710 15924
rect -690 15830 -686 15924
rect -666 15830 -662 15924
rect -642 15830 -638 15924
rect -618 15830 -614 15924
rect -594 15830 -590 15924
rect -570 15830 -566 15924
rect -546 15830 -542 15924
rect -522 15830 -518 15924
rect -498 15830 -494 15924
rect -474 15830 -470 15924
rect -450 15830 -446 15924
rect -426 15830 -422 15924
rect -402 15830 -398 15924
rect -378 15830 -374 15924
rect -354 15830 -350 15924
rect -330 15830 -326 15924
rect -306 15830 -302 15924
rect -282 15830 -278 15924
rect -258 15830 -254 15924
rect -234 15830 -230 15924
rect -210 15830 -206 15924
rect -186 15830 -182 15924
rect -162 15830 -158 15924
rect -138 15830 -134 15924
rect -114 15830 -110 15924
rect -90 15830 -86 15924
rect -66 15830 -62 15924
rect -42 15830 -38 15924
rect -18 15830 -14 15924
rect 6 15830 10 15924
rect 30 15830 34 15924
rect 54 15830 58 15924
rect 78 15830 82 15924
rect 102 15830 106 15924
rect 126 15830 130 15924
rect 150 15830 154 15924
rect 174 15830 178 15924
rect 198 15830 202 15924
rect 222 15830 226 15924
rect 246 15830 250 15924
rect 270 15830 274 15924
rect 294 15830 298 15924
rect 318 15830 322 15924
rect 342 15830 346 15924
rect 366 15830 370 15924
rect 390 15830 394 15924
rect 414 15830 418 15924
rect 438 15830 442 15924
rect 462 15830 466 15924
rect 486 15830 490 15924
rect 510 15830 514 15924
rect 534 15830 538 15924
rect 558 15830 562 15924
rect 582 15830 586 15924
rect 606 15830 610 15924
rect 630 15830 634 15924
rect 654 15830 658 15924
rect 678 15830 682 15924
rect 702 15830 706 15924
rect 726 15830 730 15924
rect 750 15830 754 15924
rect 774 15830 778 15924
rect 798 15830 802 15924
rect 822 15830 826 15924
rect 846 15830 850 15924
rect 870 15830 874 15924
rect 894 15830 898 15924
rect 918 15830 922 15924
rect 942 15830 946 15924
rect 955 15893 960 15903
rect 966 15893 970 15924
rect 965 15879 970 15893
rect 966 15830 970 15879
rect 990 15830 994 15924
rect 1014 15830 1018 15924
rect 1038 15830 1042 15924
rect 1062 15830 1066 15924
rect 1086 15830 1090 15924
rect 1110 15830 1114 15924
rect 1134 15830 1138 15924
rect 1158 15830 1162 15924
rect 1182 15830 1186 15924
rect 1206 15830 1210 15924
rect 1230 15830 1234 15924
rect 1254 15830 1258 15924
rect 1278 15830 1282 15924
rect 1302 15830 1306 15924
rect 1326 15830 1330 15924
rect 1350 15830 1354 15924
rect 1374 15830 1378 15924
rect 1398 15830 1402 15924
rect 1422 15830 1426 15924
rect 1446 15830 1450 15924
rect 1470 15830 1474 15924
rect 1494 15830 1498 15924
rect 1518 15830 1522 15924
rect 1542 15830 1546 15924
rect 1566 15830 1570 15924
rect 1590 15830 1594 15924
rect 1614 15830 1618 15924
rect 1638 15830 1642 15924
rect 1662 15830 1666 15924
rect 1686 15830 1690 15924
rect 1710 15830 1714 15924
rect 1734 15830 1738 15924
rect 1758 15830 1762 15924
rect 1782 15830 1786 15924
rect 1806 15830 1810 15924
rect 1830 15830 1834 15924
rect 1854 15830 1858 15924
rect 1878 15830 1882 15924
rect 1902 15830 1906 15924
rect 1926 15830 1930 15924
rect 1950 15830 1954 15924
rect 1974 15830 1978 15924
rect 1998 15830 2002 15924
rect 2022 15830 2026 15924
rect 2046 15830 2050 15924
rect 2059 15917 2064 15924
rect 2070 15917 2074 15924
rect 2069 15903 2074 15917
rect 2059 15893 2064 15903
rect 2069 15879 2074 15893
rect 2070 15830 2074 15879
rect 2094 15851 2098 16020
rect -2393 15828 2091 15830
rect -2371 15806 -2366 15828
rect -2348 15806 -2343 15828
rect -2325 15816 -2317 15828
rect -2325 15806 -2320 15816
rect -2317 15814 -2309 15816
rect -2062 15815 -2032 15822
rect -2309 15806 -2301 15814
rect -2070 15808 -2062 15815
rect -2000 15810 -1992 15828
rect -1974 15826 -1944 15828
rect -1960 15825 -1944 15826
rect -1842 15824 -1806 15828
rect -1842 15817 -1798 15822
rect -1806 15815 -1798 15817
rect -1671 15816 -1663 15828
rect -1854 15813 -1842 15815
rect -1663 15814 -1655 15816
rect -2062 15806 -2036 15808
rect -2393 15804 -2036 15806
rect -2032 15806 -2012 15808
rect -2004 15806 -1974 15810
rect -1854 15808 -1806 15813
rect -1864 15806 -1796 15807
rect -1655 15806 -1647 15814
rect -1642 15806 -1637 15828
rect -1619 15806 -1614 15828
rect -1530 15806 -1526 15828
rect -1506 15806 -1502 15828
rect -1482 15806 -1478 15828
rect -1458 15806 -1454 15828
rect -1434 15806 -1430 15828
rect -1410 15806 -1406 15828
rect -1386 15806 -1382 15828
rect -1362 15806 -1358 15828
rect -1338 15806 -1334 15828
rect -1314 15806 -1310 15828
rect -1290 15806 -1286 15828
rect -1266 15806 -1262 15828
rect -1242 15806 -1238 15828
rect -1218 15806 -1214 15828
rect -1194 15806 -1190 15828
rect -1170 15806 -1166 15828
rect -1146 15806 -1142 15828
rect -1122 15806 -1118 15828
rect -1098 15806 -1094 15828
rect -1074 15806 -1070 15828
rect -1050 15806 -1046 15828
rect -1026 15806 -1022 15828
rect -1002 15806 -998 15828
rect -978 15806 -974 15828
rect -954 15807 -950 15828
rect -965 15806 -931 15807
rect -2032 15804 -931 15806
rect -2371 15758 -2366 15804
rect -2348 15758 -2343 15804
rect -2325 15800 -2320 15804
rect -2309 15802 -2301 15804
rect -2317 15800 -2309 15802
rect -2325 15788 -2317 15800
rect -2052 15798 -2036 15800
rect -2052 15796 -2032 15798
rect -2062 15790 -2032 15796
rect -2325 15768 -2320 15788
rect -2317 15786 -2309 15788
rect -2092 15774 -2062 15776
rect -2094 15770 -2062 15774
rect -2325 15758 -2317 15768
rect -2095 15760 -2084 15764
rect -2000 15761 -1992 15804
rect -1904 15797 -1874 15804
rect -1842 15797 -1806 15804
rect -1655 15802 -1647 15804
rect -1663 15800 -1655 15802
rect -1842 15790 -1680 15796
rect -1671 15788 -1663 15800
rect -1663 15786 -1655 15788
rect -1854 15774 -1806 15776
rect -1854 15770 -1680 15774
rect -2119 15758 -2069 15760
rect -2054 15758 -1892 15761
rect -1671 15758 -1663 15768
rect -1642 15758 -1637 15804
rect -1619 15758 -1614 15804
rect -1530 15758 -1526 15804
rect -1506 15758 -1502 15804
rect -1482 15758 -1478 15804
rect -1458 15758 -1454 15804
rect -1434 15758 -1430 15804
rect -1410 15758 -1406 15804
rect -1386 15758 -1382 15804
rect -1362 15758 -1358 15804
rect -1338 15758 -1334 15804
rect -1314 15758 -1310 15804
rect -1290 15758 -1286 15804
rect -1266 15758 -1262 15804
rect -1242 15758 -1238 15804
rect -1218 15758 -1214 15804
rect -1194 15758 -1190 15804
rect -1170 15758 -1166 15804
rect -1146 15758 -1142 15804
rect -1122 15758 -1118 15804
rect -1098 15758 -1094 15804
rect -1074 15758 -1070 15804
rect -1050 15758 -1046 15804
rect -1026 15758 -1022 15804
rect -1002 15758 -998 15804
rect -978 15758 -974 15804
rect -965 15797 -960 15804
rect -954 15797 -950 15804
rect -955 15783 -950 15797
rect -954 15758 -950 15783
rect -930 15758 -926 15828
rect -906 15758 -902 15828
rect -882 15758 -878 15828
rect -858 15758 -854 15828
rect -834 15758 -830 15828
rect -810 15758 -806 15828
rect -786 15758 -782 15828
rect -762 15758 -758 15828
rect -738 15758 -734 15828
rect -714 15758 -710 15828
rect -690 15758 -686 15828
rect -666 15758 -662 15828
rect -642 15758 -638 15828
rect -618 15758 -614 15828
rect -594 15758 -590 15828
rect -570 15758 -566 15828
rect -546 15758 -542 15828
rect -522 15758 -518 15828
rect -498 15758 -494 15828
rect -474 15758 -470 15828
rect -450 15758 -446 15828
rect -426 15758 -422 15828
rect -402 15758 -398 15828
rect -378 15758 -374 15828
rect -354 15758 -350 15828
rect -330 15758 -326 15828
rect -306 15758 -302 15828
rect -282 15758 -278 15828
rect -258 15758 -254 15828
rect -234 15758 -230 15828
rect -210 15758 -206 15828
rect -186 15758 -182 15828
rect -162 15758 -158 15828
rect -138 15758 -134 15828
rect -114 15758 -110 15828
rect -90 15758 -86 15828
rect -66 15758 -62 15828
rect -42 15758 -38 15828
rect -18 15758 -14 15828
rect 6 15758 10 15828
rect 30 15758 34 15828
rect 54 15758 58 15828
rect 78 15758 82 15828
rect 102 15758 106 15828
rect 126 15758 130 15828
rect 150 15758 154 15828
rect 174 15758 178 15828
rect 198 15758 202 15828
rect 222 15758 226 15828
rect 246 15758 250 15828
rect 270 15758 274 15828
rect 294 15758 298 15828
rect 318 15758 322 15828
rect 342 15758 346 15828
rect 366 15758 370 15828
rect 390 15758 394 15828
rect 414 15758 418 15828
rect 438 15758 442 15828
rect 462 15758 466 15828
rect 486 15758 490 15828
rect 510 15758 514 15828
rect 534 15758 538 15828
rect 558 15758 562 15828
rect 582 15758 586 15828
rect 606 15758 610 15828
rect 630 15758 634 15828
rect 654 15758 658 15828
rect 678 15758 682 15828
rect 702 15758 706 15828
rect 726 15758 730 15828
rect 750 15758 754 15828
rect 774 15758 778 15828
rect 798 15758 802 15828
rect 822 15758 826 15828
rect 846 15758 850 15828
rect 870 15758 874 15828
rect 894 15758 898 15828
rect 918 15758 922 15828
rect 942 15758 946 15828
rect 966 15758 970 15828
rect 990 15827 994 15828
rect 990 15803 997 15827
rect 990 15758 994 15803
rect 1014 15758 1018 15828
rect 1038 15758 1042 15828
rect 1062 15758 1066 15828
rect 1086 15758 1090 15828
rect 1110 15758 1114 15828
rect 1134 15758 1138 15828
rect 1158 15758 1162 15828
rect 1182 15758 1186 15828
rect 1206 15758 1210 15828
rect 1230 15758 1234 15828
rect 1254 15758 1258 15828
rect 1278 15758 1282 15828
rect 1302 15758 1306 15828
rect 1326 15758 1330 15828
rect 1350 15758 1354 15828
rect 1374 15758 1378 15828
rect 1398 15758 1402 15828
rect 1422 15758 1426 15828
rect 1446 15758 1450 15828
rect 1470 15758 1474 15828
rect 1494 15758 1498 15828
rect 1518 15758 1522 15828
rect 1542 15758 1546 15828
rect 1566 15758 1570 15828
rect 1590 15758 1594 15828
rect 1614 15758 1618 15828
rect 1638 15758 1642 15828
rect 1662 15758 1666 15828
rect 1686 15758 1690 15828
rect 1710 15758 1714 15828
rect 1734 15758 1738 15828
rect 1758 15758 1762 15828
rect 1782 15758 1786 15828
rect 1806 15758 1810 15828
rect 1830 15758 1834 15828
rect 1854 15758 1858 15828
rect 1878 15758 1882 15828
rect 1902 15758 1906 15828
rect 1926 15758 1930 15828
rect 1950 15758 1954 15828
rect 1974 15758 1978 15828
rect 1998 15758 2002 15828
rect 2022 15758 2026 15828
rect 2046 15758 2050 15828
rect 2070 15758 2074 15828
rect 2077 15827 2091 15828
rect 2094 15803 2101 15851
rect 2094 15758 2098 15803
rect 2118 15758 2122 16020
rect 2142 15758 2146 16020
rect 2166 15758 2170 16020
rect 2190 15758 2194 16020
rect 2214 15758 2218 16020
rect 2238 15758 2242 16020
rect 2262 15758 2266 16020
rect 2286 15758 2290 16020
rect 2310 15758 2314 16020
rect 2334 15758 2338 16020
rect 2358 15758 2362 16020
rect 2382 15758 2386 16020
rect 2406 15758 2410 16020
rect 2430 15758 2434 16020
rect 2454 15758 2458 16020
rect 2478 15758 2482 16020
rect 2502 15758 2506 16020
rect 2526 15758 2530 16020
rect 2550 15758 2554 16020
rect 2574 15758 2578 16020
rect 2598 15758 2602 16020
rect 2622 15758 2626 16020
rect 2646 15758 2650 16020
rect 2670 15758 2674 16020
rect 2694 15758 2698 16020
rect 2718 15758 2722 16020
rect 2742 15758 2746 16020
rect 2766 15758 2770 16020
rect 2790 15758 2794 16020
rect 2814 15758 2818 16020
rect 2838 15758 2842 16020
rect 2862 15758 2866 16020
rect 2886 15758 2890 16020
rect 2910 15758 2914 16020
rect 2934 15758 2938 16020
rect 2958 15758 2962 16020
rect 2982 15758 2986 16020
rect 3006 15758 3010 16020
rect 3030 15758 3034 16020
rect 3054 15758 3058 16020
rect 3078 15758 3082 16020
rect 3102 15758 3106 16020
rect 3126 15758 3130 16020
rect 3150 15758 3154 16020
rect 3163 16013 3168 16020
rect 3174 16013 3178 16020
rect 3173 15999 3178 16013
rect 3163 15989 3168 15999
rect 3173 15975 3178 15989
rect 3174 15758 3178 15975
rect 3198 15947 3202 16236
rect 3198 15902 3205 15947
rect 3222 15902 3226 16236
rect 3246 15902 3250 16236
rect 3270 15902 3274 16236
rect 3294 15902 3298 16236
rect 3318 15902 3322 16236
rect 3342 15902 3346 16236
rect 3366 15902 3370 16236
rect 3390 15902 3394 16236
rect 3414 15902 3418 16236
rect 3438 15902 3442 16236
rect 3462 15902 3466 16236
rect 3486 15902 3490 16236
rect 3510 15902 3514 16236
rect 3534 15902 3538 16236
rect 3558 15902 3562 16236
rect 3582 15902 3586 16236
rect 3606 15902 3610 16236
rect 3630 15902 3634 16236
rect 3654 15902 3658 16236
rect 3667 15989 3672 15999
rect 3678 15989 3682 16236
rect 3691 16037 3696 16047
rect 3702 16037 3706 16236
rect 3715 16109 3720 16119
rect 3726 16109 3730 16236
rect 3739 16229 3744 16236
rect 3750 16229 3754 16236
rect 3757 16235 3771 16236
rect 3749 16215 3754 16229
rect 3725 16095 3730 16109
rect 3701 16023 3706 16037
rect 3677 15975 3682 15989
rect 3667 15965 3672 15975
rect 3677 15951 3682 15965
rect 3678 15903 3682 15951
rect 3667 15902 3699 15903
rect 3181 15900 3699 15902
rect 3181 15899 3195 15900
rect 3198 15899 3205 15900
rect 3198 15758 3202 15899
rect 3222 15758 3226 15900
rect 3246 15758 3250 15900
rect 3259 15821 3264 15831
rect 3270 15821 3274 15900
rect 3269 15807 3274 15821
rect 3270 15758 3274 15807
rect 3294 15758 3298 15900
rect 3318 15758 3322 15900
rect 3342 15758 3346 15900
rect 3366 15758 3370 15900
rect 3390 15758 3394 15900
rect 3414 15758 3418 15900
rect 3438 15758 3442 15900
rect 3462 15758 3466 15900
rect 3486 15758 3490 15900
rect 3510 15758 3514 15900
rect 3534 15758 3538 15900
rect 3558 15758 3562 15900
rect 3582 15758 3586 15900
rect 3606 15758 3610 15900
rect 3630 15758 3634 15900
rect 3654 15758 3658 15900
rect 3667 15893 3672 15900
rect 3678 15893 3682 15900
rect 3685 15899 3699 15900
rect 3677 15879 3682 15893
rect 3691 15889 3699 15893
rect 3685 15879 3691 15889
rect 3667 15845 3672 15855
rect 3677 15831 3682 15845
rect 3678 15758 3682 15831
rect 3691 15758 3699 15759
rect -2393 15756 3699 15758
rect -2371 15734 -2366 15756
rect -2348 15734 -2343 15756
rect -2325 15752 -2317 15756
rect -2325 15736 -2320 15752
rect -2309 15740 -2301 15752
rect -2095 15750 -2084 15756
rect -2054 15755 -1906 15756
rect -2054 15754 -2036 15755
rect -2084 15748 -2079 15750
rect -2317 15736 -2309 15740
rect -2092 15739 -2079 15746
rect -2000 15742 -1992 15755
rect -1920 15754 -1906 15755
rect -1671 15752 -1663 15756
rect -1846 15748 -1806 15750
rect -1854 15742 -1806 15746
rect -2054 15739 -1982 15742
rect -1966 15739 -1806 15742
rect -1655 15740 -1647 15752
rect -2003 15736 -1992 15739
rect -1904 15737 -1902 15739
rect -1854 15737 -1846 15739
rect -2325 15734 -2317 15736
rect -2033 15734 -1992 15736
rect -1854 15735 -1806 15737
rect -1663 15736 -1655 15740
rect -1864 15734 -1796 15735
rect -1671 15734 -1663 15736
rect -1642 15734 -1637 15756
rect -1619 15734 -1614 15756
rect -1530 15734 -1526 15756
rect -1506 15734 -1502 15756
rect -1482 15734 -1478 15756
rect -1458 15734 -1454 15756
rect -1434 15734 -1430 15756
rect -1410 15734 -1406 15756
rect -1386 15734 -1382 15756
rect -1362 15734 -1358 15756
rect -1338 15734 -1334 15756
rect -1314 15734 -1310 15756
rect -1290 15734 -1286 15756
rect -1266 15734 -1262 15756
rect -1242 15734 -1238 15756
rect -1218 15734 -1214 15756
rect -1194 15734 -1190 15756
rect -1170 15734 -1166 15756
rect -1146 15734 -1142 15756
rect -1122 15734 -1118 15756
rect -1098 15734 -1094 15756
rect -1074 15734 -1070 15756
rect -1050 15734 -1046 15756
rect -1026 15734 -1022 15756
rect -1002 15734 -998 15756
rect -978 15734 -974 15756
rect -954 15734 -950 15756
rect -930 15734 -926 15756
rect -906 15734 -902 15756
rect -882 15734 -878 15756
rect -858 15734 -854 15756
rect -834 15734 -830 15756
rect -810 15734 -806 15756
rect -786 15734 -782 15756
rect -762 15734 -758 15756
rect -738 15734 -734 15756
rect -714 15734 -710 15756
rect -690 15734 -686 15756
rect -666 15734 -662 15756
rect -642 15734 -638 15756
rect -618 15734 -614 15756
rect -594 15734 -590 15756
rect -570 15734 -566 15756
rect -546 15734 -542 15756
rect -522 15734 -518 15756
rect -498 15734 -494 15756
rect -474 15734 -470 15756
rect -450 15734 -446 15756
rect -426 15734 -422 15756
rect -402 15734 -398 15756
rect -378 15734 -374 15756
rect -354 15734 -350 15756
rect -330 15734 -326 15756
rect -306 15734 -302 15756
rect -282 15734 -278 15756
rect -258 15734 -254 15756
rect -234 15734 -230 15756
rect -210 15734 -206 15756
rect -186 15734 -182 15756
rect -162 15734 -158 15756
rect -138 15734 -134 15756
rect -114 15734 -110 15756
rect -90 15734 -86 15756
rect -66 15734 -62 15756
rect -42 15734 -38 15756
rect -18 15734 -14 15756
rect 6 15734 10 15756
rect 30 15734 34 15756
rect 54 15735 58 15756
rect 43 15734 77 15735
rect -2393 15732 77 15734
rect -2371 15710 -2366 15732
rect -2348 15710 -2343 15732
rect -2325 15724 -2317 15732
rect -2079 15729 -2018 15732
rect -2003 15731 -1966 15732
rect -2000 15730 -1982 15731
rect -2000 15729 -1992 15730
rect -2084 15725 -2009 15729
rect -2028 15724 -2009 15725
rect -2000 15725 -1854 15729
rect -1846 15725 -1798 15732
rect -2325 15710 -2320 15724
rect -2309 15712 -2301 15724
rect -2028 15722 -2018 15724
rect -2092 15712 -2084 15719
rect -2023 15715 -2014 15722
rect -2000 15715 -1992 15725
rect -1671 15724 -1663 15732
rect -1846 15721 -1806 15723
rect -1854 15715 -1806 15719
rect -2054 15712 -1806 15715
rect -1655 15712 -1647 15724
rect -2317 15710 -2309 15712
rect -2054 15710 -2024 15712
rect -2000 15710 -1992 15712
rect -1663 15710 -1655 15712
rect -1642 15710 -1637 15732
rect -1619 15710 -1614 15732
rect -1530 15710 -1526 15732
rect -1506 15710 -1502 15732
rect -1482 15710 -1478 15732
rect -1458 15710 -1454 15732
rect -1434 15710 -1430 15732
rect -1410 15710 -1406 15732
rect -1386 15710 -1382 15732
rect -1362 15710 -1358 15732
rect -1338 15710 -1334 15732
rect -1314 15710 -1310 15732
rect -1290 15710 -1286 15732
rect -1266 15710 -1262 15732
rect -1242 15710 -1238 15732
rect -1218 15710 -1214 15732
rect -1194 15710 -1190 15732
rect -1170 15710 -1166 15732
rect -1146 15710 -1142 15732
rect -1122 15710 -1118 15732
rect -1098 15710 -1094 15732
rect -1074 15710 -1070 15732
rect -1050 15710 -1046 15732
rect -1026 15710 -1022 15732
rect -1002 15710 -998 15732
rect -978 15710 -974 15732
rect -954 15710 -950 15732
rect -930 15731 -926 15732
rect -941 15710 -933 15711
rect -2393 15708 -2064 15710
rect -2060 15708 -933 15710
rect -2371 15662 -2366 15708
rect -2348 15662 -2343 15708
rect -2325 15696 -2317 15708
rect -2060 15705 -2054 15708
rect -2084 15698 -2054 15705
rect -2050 15702 -2044 15704
rect -2325 15676 -2320 15696
rect -2064 15694 -2054 15698
rect -2325 15668 -2317 15676
rect -2101 15671 -2071 15674
rect -2325 15662 -2320 15668
rect -2317 15662 -2309 15668
rect -2000 15666 -1992 15708
rect -1846 15707 -1806 15708
rect -1846 15698 -1798 15705
rect -1671 15696 -1663 15708
rect -1846 15694 -1806 15696
rect -1854 15680 -1680 15684
rect -1846 15671 -1798 15674
rect -2079 15665 -2043 15666
rect -2007 15665 -1991 15666
rect -2079 15664 -2071 15665
rect -2079 15662 -2029 15664
rect -2011 15662 -1991 15665
rect -1846 15663 -1806 15669
rect -1671 15668 -1663 15676
rect -1864 15662 -1796 15663
rect -1663 15662 -1655 15668
rect -1642 15662 -1637 15708
rect -1619 15662 -1614 15708
rect -1530 15662 -1526 15708
rect -1506 15662 -1502 15708
rect -1482 15662 -1478 15708
rect -1458 15662 -1454 15708
rect -1434 15662 -1430 15708
rect -1410 15662 -1406 15708
rect -1386 15662 -1382 15708
rect -1362 15662 -1358 15708
rect -1338 15662 -1334 15708
rect -1314 15662 -1310 15708
rect -1290 15662 -1286 15708
rect -1266 15662 -1262 15708
rect -1242 15662 -1238 15708
rect -1218 15662 -1214 15708
rect -1194 15662 -1190 15708
rect -1170 15662 -1166 15708
rect -1146 15662 -1142 15708
rect -1122 15662 -1118 15708
rect -1098 15662 -1094 15708
rect -1074 15662 -1070 15708
rect -1050 15662 -1046 15708
rect -1026 15662 -1022 15708
rect -1002 15662 -998 15708
rect -978 15663 -974 15708
rect -989 15662 -955 15663
rect -2393 15660 -955 15662
rect -2371 15614 -2366 15660
rect -2348 15614 -2343 15660
rect -2325 15648 -2320 15660
rect -2079 15658 -2071 15660
rect -2072 15656 -2071 15658
rect -2109 15651 -2101 15656
rect -2101 15649 -2079 15651
rect -2069 15649 -2068 15656
rect -2325 15640 -2317 15648
rect -2079 15644 -2071 15649
rect -2325 15620 -2320 15640
rect -2317 15632 -2309 15640
rect -2074 15635 -2071 15644
rect -2069 15640 -2068 15644
rect -2109 15626 -2079 15629
rect -2325 15614 -2317 15620
rect -2000 15614 -1992 15660
rect -1846 15658 -1806 15660
rect -1854 15653 -1806 15657
rect -1854 15651 -1846 15653
rect -1846 15649 -1806 15651
rect -1806 15647 -1798 15649
rect -1846 15644 -1798 15647
rect -1846 15631 -1806 15642
rect -1671 15640 -1663 15648
rect -1663 15632 -1655 15640
rect -1854 15626 -1680 15630
rect -1671 15614 -1663 15620
rect -1642 15614 -1637 15660
rect -1619 15614 -1614 15660
rect -1530 15614 -1526 15660
rect -1506 15614 -1502 15660
rect -1482 15614 -1478 15660
rect -1458 15614 -1454 15660
rect -1434 15614 -1430 15660
rect -1410 15614 -1406 15660
rect -1386 15614 -1382 15660
rect -1362 15614 -1358 15660
rect -1338 15614 -1334 15660
rect -1314 15614 -1310 15660
rect -1290 15614 -1286 15660
rect -1266 15614 -1262 15660
rect -1242 15614 -1238 15660
rect -1218 15614 -1214 15660
rect -1194 15614 -1190 15660
rect -1170 15614 -1166 15660
rect -1146 15614 -1142 15660
rect -1122 15614 -1118 15660
rect -1098 15614 -1094 15660
rect -1074 15614 -1070 15660
rect -1050 15614 -1046 15660
rect -1026 15614 -1022 15660
rect -1002 15614 -998 15660
rect -989 15653 -984 15660
rect -978 15653 -974 15660
rect -979 15639 -974 15653
rect -989 15638 -955 15639
rect -954 15638 -950 15708
rect -947 15707 -933 15708
rect -930 15707 -923 15731
rect -941 15701 -936 15707
rect -930 15701 -926 15707
rect -931 15687 -926 15701
rect -941 15662 -907 15663
rect -906 15662 -902 15732
rect -882 15662 -878 15732
rect -858 15662 -854 15732
rect -834 15662 -830 15732
rect -810 15662 -806 15732
rect -786 15662 -782 15732
rect -762 15662 -758 15732
rect -738 15662 -734 15732
rect -714 15662 -710 15732
rect -690 15662 -686 15732
rect -666 15662 -662 15732
rect -642 15662 -638 15732
rect -618 15662 -614 15732
rect -594 15662 -590 15732
rect -570 15662 -566 15732
rect -546 15662 -542 15732
rect -522 15662 -518 15732
rect -509 15677 -504 15687
rect -498 15677 -494 15732
rect -499 15663 -494 15677
rect -474 15662 -470 15732
rect -450 15662 -446 15732
rect -426 15662 -422 15732
rect -402 15662 -398 15732
rect -378 15662 -374 15732
rect -354 15662 -350 15732
rect -330 15662 -326 15732
rect -306 15662 -302 15732
rect -282 15662 -278 15732
rect -258 15662 -254 15732
rect -234 15662 -230 15732
rect -210 15662 -206 15732
rect -186 15662 -182 15732
rect -162 15662 -158 15732
rect -138 15662 -134 15732
rect -114 15662 -110 15732
rect -90 15662 -86 15732
rect -66 15662 -62 15732
rect -42 15662 -38 15732
rect -18 15662 -14 15732
rect 6 15662 10 15732
rect 30 15662 34 15732
rect 43 15725 48 15732
rect 54 15725 58 15732
rect 53 15711 58 15725
rect 43 15701 48 15711
rect 53 15687 58 15701
rect 54 15662 58 15687
rect 78 15662 82 15756
rect 102 15662 106 15756
rect 126 15662 130 15756
rect 150 15662 154 15756
rect 174 15662 178 15756
rect 198 15662 202 15756
rect 222 15662 226 15756
rect 246 15662 250 15756
rect 270 15662 274 15756
rect 294 15662 298 15756
rect 318 15662 322 15756
rect 342 15662 346 15756
rect 366 15662 370 15756
rect 390 15662 394 15756
rect 414 15662 418 15756
rect 438 15662 442 15756
rect 462 15662 466 15756
rect 486 15662 490 15756
rect 510 15662 514 15756
rect 534 15662 538 15756
rect 558 15662 562 15756
rect 582 15662 586 15756
rect 606 15662 610 15756
rect 630 15662 634 15756
rect 654 15662 658 15756
rect 678 15662 682 15756
rect 702 15662 706 15756
rect 726 15662 730 15756
rect 750 15662 754 15756
rect 774 15662 778 15756
rect 798 15662 802 15756
rect 822 15662 826 15756
rect 846 15662 850 15756
rect 870 15662 874 15756
rect 894 15662 898 15756
rect 918 15662 922 15756
rect 942 15662 946 15756
rect 966 15662 970 15756
rect 990 15662 994 15756
rect 1014 15662 1018 15756
rect 1038 15662 1042 15756
rect 1062 15662 1066 15756
rect 1086 15662 1090 15756
rect 1110 15662 1114 15756
rect 1134 15662 1138 15756
rect 1158 15662 1162 15756
rect 1182 15662 1186 15756
rect 1206 15662 1210 15756
rect 1230 15662 1234 15756
rect 1254 15662 1258 15756
rect 1278 15662 1282 15756
rect 1302 15662 1306 15756
rect 1326 15662 1330 15756
rect 1350 15662 1354 15756
rect 1374 15662 1378 15756
rect 1398 15662 1402 15756
rect 1422 15662 1426 15756
rect 1446 15662 1450 15756
rect 1470 15662 1474 15756
rect 1494 15662 1498 15756
rect 1518 15662 1522 15756
rect 1542 15662 1546 15756
rect 1566 15662 1570 15756
rect 1590 15662 1594 15756
rect 1614 15662 1618 15756
rect 1638 15662 1642 15756
rect 1662 15662 1666 15756
rect 1686 15662 1690 15756
rect 1710 15662 1714 15756
rect 1734 15662 1738 15756
rect 1758 15662 1762 15756
rect 1782 15662 1786 15756
rect 1806 15662 1810 15756
rect 1830 15662 1834 15756
rect 1854 15662 1858 15756
rect 1878 15662 1882 15756
rect 1902 15662 1906 15756
rect 1926 15662 1930 15756
rect 1950 15662 1954 15756
rect 1974 15662 1978 15756
rect 1998 15662 2002 15756
rect 2022 15662 2026 15756
rect 2046 15662 2050 15756
rect 2070 15662 2074 15756
rect 2094 15662 2098 15756
rect 2118 15662 2122 15756
rect 2142 15662 2146 15756
rect 2166 15662 2170 15756
rect 2190 15662 2194 15756
rect 2214 15662 2218 15756
rect 2238 15662 2242 15756
rect 2262 15662 2266 15756
rect 2286 15662 2290 15756
rect 2310 15662 2314 15756
rect 2334 15662 2338 15756
rect 2358 15662 2362 15756
rect 2382 15662 2386 15756
rect 2406 15662 2410 15756
rect 2430 15662 2434 15756
rect 2454 15662 2458 15756
rect 2478 15662 2482 15756
rect 2502 15662 2506 15756
rect 2526 15662 2530 15756
rect 2550 15662 2554 15756
rect 2574 15662 2578 15756
rect 2598 15662 2602 15756
rect 2622 15662 2626 15756
rect 2646 15662 2650 15756
rect 2670 15662 2674 15756
rect 2694 15662 2698 15756
rect 2718 15662 2722 15756
rect 2742 15662 2746 15756
rect 2766 15662 2770 15756
rect 2790 15662 2794 15756
rect 2814 15662 2818 15756
rect 2838 15662 2842 15756
rect 2862 15662 2866 15756
rect 2886 15662 2890 15756
rect 2910 15662 2914 15756
rect 2934 15662 2938 15756
rect 2958 15662 2962 15756
rect 2982 15662 2986 15756
rect 3006 15662 3010 15756
rect 3030 15662 3034 15756
rect 3054 15662 3058 15756
rect 3078 15662 3082 15756
rect 3102 15662 3106 15756
rect 3126 15662 3130 15756
rect 3150 15662 3154 15756
rect 3174 15662 3178 15756
rect 3198 15662 3202 15756
rect 3222 15662 3226 15756
rect 3246 15662 3250 15756
rect 3270 15662 3274 15756
rect 3294 15755 3298 15756
rect 3294 15731 3301 15755
rect 3294 15662 3298 15731
rect 3318 15662 3322 15756
rect 3342 15662 3346 15756
rect 3366 15662 3370 15756
rect 3390 15662 3394 15756
rect 3414 15662 3418 15756
rect 3438 15662 3442 15756
rect 3462 15662 3466 15756
rect 3486 15662 3490 15756
rect 3510 15662 3514 15756
rect 3534 15662 3538 15756
rect 3558 15662 3562 15756
rect 3582 15662 3586 15756
rect 3606 15662 3610 15756
rect 3630 15662 3634 15756
rect 3654 15662 3658 15756
rect 3678 15663 3682 15756
rect 3685 15755 3699 15756
rect 3691 15749 3696 15755
rect 3701 15735 3706 15749
rect 3691 15701 3696 15711
rect 3702 15701 3706 15735
rect 3701 15687 3706 15701
rect 3667 15662 3701 15663
rect -941 15660 3701 15662
rect -941 15653 -936 15660
rect -931 15639 -926 15653
rect -930 15638 -926 15639
rect -906 15638 -902 15660
rect -882 15638 -878 15660
rect -858 15638 -854 15660
rect -834 15638 -830 15660
rect -810 15638 -806 15660
rect -786 15638 -782 15660
rect -762 15638 -758 15660
rect -738 15638 -734 15660
rect -714 15638 -710 15660
rect -690 15638 -686 15660
rect -666 15638 -662 15660
rect -642 15638 -638 15660
rect -618 15638 -614 15660
rect -594 15638 -590 15660
rect -570 15638 -566 15660
rect -546 15638 -542 15660
rect -522 15638 -518 15660
rect -474 15638 -470 15660
rect -450 15638 -446 15660
rect -426 15638 -422 15660
rect -402 15638 -398 15660
rect -378 15638 -374 15660
rect -354 15638 -350 15660
rect -330 15638 -326 15660
rect -306 15638 -302 15660
rect -282 15638 -278 15660
rect -258 15638 -254 15660
rect -234 15638 -230 15660
rect -210 15638 -206 15660
rect -186 15638 -182 15660
rect -162 15638 -158 15660
rect -138 15638 -134 15660
rect -114 15638 -110 15660
rect -90 15638 -86 15660
rect -66 15638 -62 15660
rect -42 15638 -38 15660
rect -18 15638 -14 15660
rect 6 15638 10 15660
rect 30 15638 34 15660
rect 54 15638 58 15660
rect 78 15659 82 15660
rect -989 15636 75 15638
rect -989 15629 -984 15636
rect -979 15615 -974 15629
rect -978 15614 -974 15615
rect -954 15614 -950 15636
rect -930 15614 -926 15636
rect -906 15635 -902 15636
rect -2393 15612 -909 15614
rect -2371 15590 -2366 15612
rect -2348 15590 -2343 15612
rect -2325 15604 -2317 15612
rect -2325 15590 -2320 15604
rect -2309 15592 -2301 15604
rect -2092 15595 -2062 15600
rect -2000 15592 -1992 15612
rect -2317 15590 -2309 15592
rect -2000 15590 -1983 15592
rect -1906 15590 -1904 15612
rect -1806 15604 -1680 15610
rect -1671 15604 -1663 15612
rect -1854 15595 -1806 15600
rect -1846 15590 -1806 15593
rect -1655 15592 -1647 15604
rect -1663 15590 -1655 15592
rect -1642 15590 -1637 15612
rect -1619 15590 -1614 15612
rect -1530 15590 -1526 15612
rect -1506 15590 -1502 15612
rect -1482 15590 -1478 15612
rect -1458 15590 -1454 15612
rect -1434 15590 -1430 15612
rect -1410 15590 -1406 15612
rect -1386 15590 -1382 15612
rect -1362 15590 -1358 15612
rect -1338 15590 -1334 15612
rect -1314 15590 -1310 15612
rect -1290 15590 -1286 15612
rect -1266 15590 -1262 15612
rect -1242 15590 -1238 15612
rect -1218 15590 -1214 15612
rect -1194 15590 -1190 15612
rect -1170 15590 -1166 15612
rect -1146 15590 -1142 15612
rect -1122 15590 -1118 15612
rect -1098 15590 -1094 15612
rect -1074 15590 -1070 15612
rect -1050 15590 -1046 15612
rect -1026 15590 -1022 15612
rect -1002 15590 -998 15612
rect -978 15590 -974 15612
rect -954 15590 -950 15612
rect -930 15590 -926 15612
rect -923 15611 -909 15612
rect -906 15611 -899 15635
rect -882 15590 -878 15636
rect -858 15590 -854 15636
rect -834 15590 -830 15636
rect -810 15590 -806 15636
rect -786 15590 -782 15636
rect -762 15590 -758 15636
rect -738 15590 -734 15636
rect -714 15590 -710 15636
rect -690 15590 -686 15636
rect -666 15590 -662 15636
rect -642 15590 -638 15636
rect -618 15590 -614 15636
rect -594 15590 -590 15636
rect -570 15590 -566 15636
rect -546 15590 -542 15636
rect -522 15590 -518 15636
rect -509 15605 -504 15615
rect -474 15611 -470 15636
rect -499 15591 -494 15605
rect -485 15601 -477 15605
rect -491 15591 -485 15601
rect -498 15590 -494 15591
rect -2393 15588 -477 15590
rect -2371 15566 -2366 15588
rect -2348 15566 -2343 15588
rect -2325 15576 -2317 15588
rect -2071 15584 -2062 15588
rect -2013 15586 -1983 15588
rect -2000 15585 -1983 15586
rect -2325 15566 -2320 15576
rect -2309 15566 -2301 15576
rect -2100 15575 -2092 15582
rect -2064 15580 -2062 15583
rect -2061 15575 -2059 15580
rect -2071 15570 -2062 15575
rect -2071 15568 -2026 15570
rect -2066 15566 -2012 15568
rect -2000 15566 -1992 15585
rect -1906 15583 -1904 15588
rect -1846 15584 -1806 15588
rect -1846 15577 -1798 15582
rect -1806 15575 -1798 15577
rect -1671 15576 -1663 15588
rect -1854 15573 -1846 15575
rect -1854 15568 -1806 15573
rect -1864 15566 -1796 15567
rect -1655 15566 -1647 15576
rect -1642 15566 -1637 15588
rect -1619 15566 -1614 15588
rect -1530 15566 -1526 15588
rect -1506 15567 -1502 15588
rect -1517 15566 -1483 15567
rect -2393 15564 -1483 15566
rect -2371 15518 -2366 15564
rect -2348 15518 -2343 15564
rect -2325 15560 -2320 15564
rect -2317 15560 -2309 15564
rect -2325 15548 -2317 15560
rect -2066 15559 -2062 15564
rect -2147 15556 -2134 15558
rect -2292 15550 -2071 15556
rect -2325 15518 -2320 15548
rect -2092 15534 -2062 15536
rect -2094 15530 -2062 15534
rect -2000 15518 -1992 15564
rect -1846 15557 -1806 15564
rect -1663 15560 -1655 15564
rect -1846 15550 -1680 15556
rect -1671 15548 -1663 15560
rect -1854 15534 -1806 15536
rect -1854 15530 -1680 15534
rect -1642 15518 -1637 15564
rect -1619 15518 -1614 15564
rect -1530 15518 -1526 15564
rect -1517 15557 -1512 15564
rect -1506 15557 -1502 15564
rect -1507 15543 -1502 15557
rect -1506 15518 -1502 15543
rect -1482 15518 -1478 15588
rect -1458 15518 -1454 15588
rect -1434 15518 -1430 15588
rect -1410 15518 -1406 15588
rect -1386 15518 -1382 15588
rect -1362 15518 -1358 15588
rect -1338 15518 -1334 15588
rect -1314 15518 -1310 15588
rect -1290 15518 -1286 15588
rect -1266 15518 -1262 15588
rect -1242 15518 -1238 15588
rect -1218 15518 -1214 15588
rect -1194 15518 -1190 15588
rect -1170 15518 -1166 15588
rect -1146 15518 -1142 15588
rect -1122 15518 -1118 15588
rect -1098 15518 -1094 15588
rect -1074 15518 -1070 15588
rect -1050 15518 -1046 15588
rect -1026 15518 -1022 15588
rect -1002 15518 -998 15588
rect -978 15518 -974 15588
rect -954 15587 -950 15588
rect -954 15539 -947 15587
rect -954 15518 -950 15539
rect -930 15518 -926 15588
rect -906 15563 -899 15587
rect -906 15518 -902 15563
rect -882 15518 -878 15588
rect -858 15518 -854 15588
rect -834 15518 -830 15588
rect -810 15518 -806 15588
rect -786 15518 -782 15588
rect -762 15518 -758 15588
rect -738 15518 -734 15588
rect -714 15518 -710 15588
rect -690 15518 -686 15588
rect -666 15518 -662 15588
rect -642 15518 -638 15588
rect -618 15518 -614 15588
rect -594 15518 -590 15588
rect -570 15518 -566 15588
rect -546 15518 -542 15588
rect -522 15518 -518 15588
rect -498 15518 -494 15588
rect -491 15587 -477 15588
rect -474 15587 -467 15611
rect -2393 15516 -477 15518
rect -2371 15494 -2366 15516
rect -2348 15494 -2343 15516
rect -2325 15494 -2320 15516
rect -2072 15514 -2036 15515
rect -2072 15508 -2054 15514
rect -2309 15500 -2301 15508
rect -2317 15494 -2309 15500
rect -2092 15499 -2062 15504
rect -2000 15495 -1992 15516
rect -1938 15515 -1906 15516
rect -1920 15514 -1906 15515
rect -1806 15508 -1680 15514
rect -1854 15499 -1806 15504
rect -1655 15500 -1647 15508
rect -1982 15495 -1966 15496
rect -2000 15494 -1966 15495
rect -1846 15494 -1806 15497
rect -1663 15494 -1655 15500
rect -1642 15494 -1637 15516
rect -1619 15494 -1614 15516
rect -1530 15494 -1526 15516
rect -1506 15494 -1502 15516
rect -1482 15494 -1478 15516
rect -1458 15494 -1454 15516
rect -1434 15494 -1430 15516
rect -1410 15494 -1406 15516
rect -1386 15494 -1382 15516
rect -1362 15494 -1358 15516
rect -1338 15494 -1334 15516
rect -1314 15494 -1310 15516
rect -1290 15494 -1286 15516
rect -1266 15494 -1262 15516
rect -1242 15494 -1238 15516
rect -1218 15494 -1214 15516
rect -1194 15494 -1190 15516
rect -1170 15494 -1166 15516
rect -1146 15494 -1142 15516
rect -1122 15494 -1118 15516
rect -1098 15494 -1094 15516
rect -1074 15494 -1070 15516
rect -1050 15494 -1046 15516
rect -1026 15494 -1022 15516
rect -1002 15494 -998 15516
rect -978 15494 -974 15516
rect -954 15494 -950 15516
rect -930 15494 -926 15516
rect -906 15494 -902 15516
rect -882 15494 -878 15516
rect -858 15494 -854 15516
rect -834 15494 -830 15516
rect -810 15494 -806 15516
rect -786 15494 -782 15516
rect -762 15494 -758 15516
rect -738 15494 -734 15516
rect -714 15494 -710 15516
rect -690 15494 -686 15516
rect -666 15494 -662 15516
rect -642 15494 -638 15516
rect -618 15494 -614 15516
rect -594 15494 -590 15516
rect -570 15494 -566 15516
rect -546 15494 -542 15516
rect -522 15494 -518 15516
rect -498 15494 -494 15516
rect -491 15515 -477 15516
rect -474 15515 -467 15539
rect -474 15494 -470 15515
rect -450 15494 -446 15636
rect -426 15494 -422 15636
rect -402 15494 -398 15636
rect -378 15494 -374 15636
rect -354 15494 -350 15636
rect -330 15494 -326 15636
rect -306 15494 -302 15636
rect -282 15494 -278 15636
rect -258 15494 -254 15636
rect -234 15494 -230 15636
rect -210 15494 -206 15636
rect -197 15581 -192 15591
rect -186 15581 -182 15636
rect -187 15567 -182 15581
rect -197 15566 -163 15567
rect -162 15566 -158 15636
rect -138 15566 -134 15636
rect -114 15566 -110 15636
rect -90 15566 -86 15636
rect -66 15566 -62 15636
rect -42 15566 -38 15636
rect -18 15566 -14 15636
rect 6 15566 10 15636
rect 30 15566 34 15636
rect 54 15566 58 15636
rect 61 15635 75 15636
rect 78 15611 85 15659
rect 78 15566 82 15611
rect 102 15566 106 15660
rect 126 15566 130 15660
rect 150 15566 154 15660
rect 174 15566 178 15660
rect 198 15566 202 15660
rect 222 15566 226 15660
rect 246 15566 250 15660
rect 270 15566 274 15660
rect 294 15566 298 15660
rect 318 15566 322 15660
rect 342 15566 346 15660
rect 366 15566 370 15660
rect 390 15566 394 15660
rect 414 15566 418 15660
rect 438 15566 442 15660
rect 462 15566 466 15660
rect 486 15566 490 15660
rect 510 15566 514 15660
rect 534 15566 538 15660
rect 558 15566 562 15660
rect 582 15566 586 15660
rect 606 15566 610 15660
rect 630 15566 634 15660
rect 654 15566 658 15660
rect 678 15566 682 15660
rect 702 15566 706 15660
rect 726 15566 730 15660
rect 750 15566 754 15660
rect 774 15566 778 15660
rect 798 15566 802 15660
rect 822 15566 826 15660
rect 846 15566 850 15660
rect 870 15566 874 15660
rect 894 15566 898 15660
rect 918 15566 922 15660
rect 942 15566 946 15660
rect 966 15566 970 15660
rect 990 15566 994 15660
rect 1014 15566 1018 15660
rect 1038 15566 1042 15660
rect 1062 15566 1066 15660
rect 1086 15566 1090 15660
rect 1110 15566 1114 15660
rect 1134 15566 1138 15660
rect 1158 15566 1162 15660
rect 1182 15566 1186 15660
rect 1206 15566 1210 15660
rect 1230 15566 1234 15660
rect 1254 15566 1258 15660
rect 1278 15566 1282 15660
rect 1302 15566 1306 15660
rect 1326 15566 1330 15660
rect 1350 15566 1354 15660
rect 1374 15566 1378 15660
rect 1398 15566 1402 15660
rect 1422 15566 1426 15660
rect 1446 15566 1450 15660
rect 1470 15566 1474 15660
rect 1494 15566 1498 15660
rect 1518 15566 1522 15660
rect 1542 15566 1546 15660
rect 1566 15566 1570 15660
rect 1590 15566 1594 15660
rect 1614 15566 1618 15660
rect 1638 15566 1642 15660
rect 1662 15566 1666 15660
rect 1686 15566 1690 15660
rect 1710 15566 1714 15660
rect 1734 15566 1738 15660
rect 1758 15566 1762 15660
rect 1782 15566 1786 15660
rect 1806 15566 1810 15660
rect 1830 15566 1834 15660
rect 1854 15566 1858 15660
rect 1878 15566 1882 15660
rect 1902 15566 1906 15660
rect 1926 15566 1930 15660
rect 1950 15566 1954 15660
rect 1974 15566 1978 15660
rect 1998 15566 2002 15660
rect 2022 15566 2026 15660
rect 2046 15566 2050 15660
rect 2070 15566 2074 15660
rect 2094 15566 2098 15660
rect 2118 15566 2122 15660
rect 2142 15566 2146 15660
rect 2166 15566 2170 15660
rect 2190 15566 2194 15660
rect 2214 15566 2218 15660
rect 2238 15566 2242 15660
rect 2262 15566 2266 15660
rect 2286 15566 2290 15660
rect 2310 15566 2314 15660
rect 2334 15566 2338 15660
rect 2358 15566 2362 15660
rect 2382 15566 2386 15660
rect 2406 15566 2410 15660
rect 2430 15566 2434 15660
rect 2454 15566 2458 15660
rect 2478 15566 2482 15660
rect 2502 15566 2506 15660
rect 2526 15566 2530 15660
rect 2550 15566 2554 15660
rect 2574 15566 2578 15660
rect 2598 15566 2602 15660
rect 2622 15566 2626 15660
rect 2646 15566 2650 15660
rect 2670 15566 2674 15660
rect 2694 15566 2698 15660
rect 2718 15566 2722 15660
rect 2742 15566 2746 15660
rect 2766 15566 2770 15660
rect 2790 15566 2794 15660
rect 2814 15566 2818 15660
rect 2838 15566 2842 15660
rect 2862 15566 2866 15660
rect 2886 15566 2890 15660
rect 2910 15566 2914 15660
rect 2934 15566 2938 15660
rect 2958 15566 2962 15660
rect 2982 15566 2986 15660
rect 3006 15566 3010 15660
rect 3030 15566 3034 15660
rect 3054 15566 3058 15660
rect 3078 15566 3082 15660
rect 3102 15566 3106 15660
rect 3126 15566 3130 15660
rect 3150 15566 3154 15660
rect 3174 15566 3178 15660
rect 3198 15566 3202 15660
rect 3222 15566 3226 15660
rect 3246 15566 3250 15660
rect 3270 15566 3274 15660
rect 3294 15566 3298 15660
rect 3318 15566 3322 15660
rect 3342 15566 3346 15660
rect 3366 15566 3370 15660
rect 3390 15566 3394 15660
rect 3414 15566 3418 15660
rect 3438 15566 3442 15660
rect 3462 15566 3466 15660
rect 3486 15566 3490 15660
rect 3510 15566 3514 15660
rect 3534 15566 3538 15660
rect 3558 15566 3562 15660
rect 3582 15566 3586 15660
rect 3606 15566 3610 15660
rect 3630 15567 3634 15660
rect 3643 15629 3648 15639
rect 3654 15629 3658 15660
rect 3667 15653 3672 15660
rect 3678 15653 3682 15660
rect 3677 15639 3682 15653
rect 3653 15615 3658 15629
rect 3619 15566 3653 15567
rect -197 15564 3653 15566
rect -197 15557 -192 15564
rect -187 15543 -182 15557
rect -186 15494 -182 15543
rect -162 15515 -158 15564
rect -2393 15492 -165 15494
rect -2371 15470 -2366 15492
rect -2348 15470 -2343 15492
rect -2325 15470 -2320 15492
rect -2000 15490 -1966 15492
rect -2309 15472 -2301 15480
rect -2062 15479 -2054 15486
rect -2092 15472 -2084 15479
rect -2062 15472 -2026 15474
rect -2317 15470 -2309 15472
rect -2062 15470 -2012 15472
rect -2000 15470 -1992 15490
rect -1982 15489 -1966 15490
rect -1846 15488 -1806 15492
rect -1846 15481 -1798 15486
rect -1806 15479 -1798 15481
rect -1854 15477 -1846 15479
rect -1854 15472 -1806 15477
rect -1655 15472 -1647 15480
rect -1864 15470 -1796 15471
rect -1663 15470 -1655 15472
rect -1642 15470 -1637 15492
rect -1619 15470 -1614 15492
rect -1530 15470 -1526 15492
rect -1506 15470 -1502 15492
rect -1482 15491 -1478 15492
rect -2393 15468 -1485 15470
rect -2371 15051 -2366 15468
rect -2361 15071 -2353 15081
rect -2348 15071 -2343 15468
rect -2351 15055 -2343 15071
rect -2371 15025 -2363 15051
rect -2383 14853 -2376 14863
rect -2371 14853 -2366 15025
rect -2373 14842 -2366 14853
rect -2348 14842 -2343 15055
rect -2325 15337 -2320 15468
rect -2317 15464 -2309 15468
rect -2062 15464 -2054 15468
rect -2154 15460 -2138 15462
rect -2057 15460 -2054 15464
rect -2292 15454 -2054 15460
rect -2052 15454 -2044 15464
rect -2092 15438 -2062 15440
rect -2094 15434 -2062 15438
rect -2309 15404 -2301 15413
rect -2317 15397 -2309 15404
rect -2309 15376 -2301 15384
rect -2251 15378 -2093 15384
rect -2317 15368 -2309 15376
rect -2154 15371 -2138 15374
rect -2084 15371 -2054 15376
rect -2143 15358 -2138 15364
rect -2325 15327 -2317 15337
rect -2325 15308 -2320 15327
rect -2317 15321 -2309 15327
rect -2243 15310 -2221 15318
rect -2211 15310 -2201 15330
rect -2073 15310 -2065 15328
rect -2000 15310 -1992 15468
rect -1846 15461 -1806 15468
rect -1663 15464 -1655 15468
rect -1846 15454 -1680 15460
rect -1854 15438 -1806 15440
rect -1854 15434 -1680 15438
rect -1915 15404 -1906 15414
rect -1846 15412 -1837 15414
rect -1790 15412 -1680 15414
rect -1655 15404 -1647 15410
rect -1905 15395 -1896 15404
rect -1837 15403 -1790 15404
rect -1837 15388 -1798 15401
rect -1663 15394 -1655 15404
rect -1798 15378 -1790 15383
rect -1837 15376 -1798 15378
rect -1655 15376 -1647 15382
rect -1846 15374 -1837 15376
rect -1846 15371 -1798 15374
rect -1837 15358 -1798 15368
rect -1663 15366 -1655 15376
rect -1671 15326 -1663 15334
rect -1655 15326 -1647 15328
rect -1663 15318 -1647 15326
rect -1642 15318 -1637 15468
rect -1885 15310 -1877 15312
rect -1708 15310 -1672 15312
rect -2243 15309 -2213 15310
rect -2325 15299 -2317 15308
rect -2259 15303 -2211 15309
rect -2183 15303 -1877 15310
rect -1869 15303 -1758 15310
rect -1710 15304 -1672 15310
rect -1710 15303 -1692 15304
rect -2211 15299 -2201 15303
rect -2325 15279 -2320 15299
rect -2317 15292 -2309 15299
rect -2211 15292 -2198 15299
rect -2325 15271 -2317 15279
rect -2300 15272 -2292 15282
rect -2243 15273 -2228 15284
rect -2211 15276 -2181 15292
rect -2211 15273 -2201 15276
rect -2325 15251 -2320 15271
rect -2317 15263 -2309 15271
rect -2325 15243 -2317 15251
rect -2325 15223 -2320 15243
rect -2317 15235 -2309 15243
rect -2325 15214 -2317 15223
rect -2325 15195 -2320 15214
rect -2317 15207 -2309 15214
rect -2325 15186 -2317 15195
rect -2325 15166 -2320 15186
rect -2317 15179 -2309 15186
rect -2325 15158 -2317 15166
rect -2290 15159 -2282 15272
rect -2251 15262 -2240 15266
rect -2211 15262 -2181 15266
rect -2251 15259 -2181 15262
rect -2176 15252 -2173 15254
rect -2240 15245 -2173 15252
rect -2169 15247 -2163 15302
rect -2073 15266 -2065 15303
rect -2073 15262 -2043 15266
rect -2000 15262 -1992 15303
rect -1915 15272 -1907 15281
rect -1963 15266 -1955 15272
rect -1963 15262 -1915 15266
rect -1885 15262 -1877 15303
rect -1875 15298 -1869 15302
rect -1829 15280 -1781 15282
rect -1847 15276 -1781 15280
rect -1778 15276 -1771 15302
rect -1758 15295 -1710 15302
rect -1718 15288 -1710 15295
rect -1768 15278 -1760 15288
rect -1718 15286 -1700 15288
rect -2146 15259 -2135 15262
rect -2105 15259 -2043 15262
rect -2035 15259 -1989 15262
rect -1973 15259 -1915 15262
rect -1907 15259 -1854 15262
rect -2073 15257 -2043 15259
rect -2135 15245 -2105 15252
rect -2065 15250 -2043 15257
rect -2243 15234 -2240 15243
rect -2221 15237 -2213 15245
rect -2211 15237 -2208 15245
rect -2203 15238 -2173 15245
rect -2251 15227 -2240 15234
rect -2211 15234 -2203 15237
rect -2211 15227 -2181 15234
rect -2073 15227 -2043 15234
rect -2203 15204 -2173 15211
rect -2262 15186 -2240 15196
rect -2203 15195 -2176 15204
rect -2083 15193 -2075 15203
rect -2040 15193 -2035 15197
rect -2073 15181 -2043 15193
rect -2028 15181 -2023 15193
rect -2000 15186 -1992 15259
rect -1963 15256 -1955 15259
rect -1963 15255 -1915 15256
rect -1955 15245 -1907 15252
rect -1885 15248 -1877 15259
rect -1837 15254 -1828 15270
rect -1758 15263 -1750 15278
rect -1758 15262 -1692 15263
rect -1837 15252 -1833 15254
rect -1837 15250 -1835 15252
rect -1887 15245 -1851 15248
rect -1750 15245 -1702 15252
rect -1885 15240 -1877 15245
rect -1963 15227 -1915 15234
rect -1905 15195 -1897 15240
rect -1857 15222 -1851 15245
rect -1760 15237 -1758 15238
rect -1837 15227 -1789 15234
rect -1758 15228 -1750 15234
rect -1758 15227 -1710 15228
rect -1955 15192 -1915 15195
rect -1963 15186 -1962 15188
rect -2000 15183 -1981 15186
rect -1965 15183 -1962 15186
rect -1955 15186 -1907 15190
rect -1885 15186 -1877 15205
rect -1857 15192 -1851 15204
rect -1750 15200 -1702 15207
rect -1829 15192 -1789 15194
rect -1766 15190 -1760 15200
rect -1829 15186 -1781 15190
rect -1756 15186 -1740 15190
rect -1680 15186 -1672 15304
rect -1671 15298 -1663 15306
rect -1645 15302 -1637 15318
rect -1663 15290 -1655 15298
rect -1671 15270 -1663 15278
rect -1663 15262 -1655 15270
rect -1671 15242 -1663 15250
rect -1671 15226 -1669 15239
rect -1663 15234 -1655 15242
rect -1671 15214 -1663 15222
rect -1663 15206 -1655 15214
rect -1671 15186 -1663 15194
rect -1955 15183 -1837 15186
rect -1829 15183 -1740 15186
rect -2206 15173 -2176 15176
rect -2206 15170 -2203 15173
rect -2161 15171 -2145 15180
rect -2073 15178 -2065 15181
rect -2073 15177 -2043 15178
rect -2028 15177 -2012 15181
rect -2073 15170 -2065 15176
rect -2203 15169 -2176 15170
rect -2065 15169 -2043 15170
rect -2262 15163 -2232 15169
rect -2176 15163 -2173 15169
rect -2043 15163 -2035 15169
rect -2325 15138 -2320 15158
rect -2317 15150 -2309 15158
rect -2153 15157 -2146 15161
rect -2325 15130 -2317 15138
rect -2300 15134 -2292 15144
rect -2325 15110 -2320 15130
rect -2317 15122 -2309 15130
rect -2325 15102 -2317 15110
rect -2325 15082 -2320 15102
rect -2317 15094 -2309 15102
rect -2290 15101 -2282 15134
rect -2273 15130 -2264 15135
rect -2206 15130 -2176 15135
rect -2262 15123 -2232 15128
rect -2198 15119 -2176 15130
rect -2198 15105 -2176 15113
rect -2166 15097 -2158 15145
rect -2143 15141 -2136 15157
rect -2143 15130 -2113 15135
rect -2073 15130 -2065 15135
rect -2065 15128 -2043 15130
rect -2043 15123 -2035 15128
rect -2065 15102 -2043 15117
rect -2006 15101 -2004 15117
rect -2265 15087 -2260 15093
rect -2143 15087 -2113 15094
rect -2270 15086 -2240 15087
rect -2270 15083 -2265 15086
rect -2325 15074 -2317 15082
rect -2325 15054 -2320 15074
rect -2317 15066 -2309 15074
rect -2113 15071 -2105 15081
rect -2291 15059 -2270 15066
rect -2198 15064 -2168 15066
rect -2135 15065 -2105 15066
rect -2103 15065 -2095 15071
rect -2113 15064 -2105 15065
rect -2065 15064 -2035 15066
rect -2000 15064 -1992 15183
rect -1963 15176 -1960 15183
rect -1915 15179 -1905 15183
rect -1963 15175 -1955 15176
rect -1963 15169 -1915 15175
rect -1989 15142 -1973 15145
rect -1915 15142 -1907 15149
rect -1990 15107 -1989 15128
rect -1983 15064 -1981 15127
rect -1885 15118 -1877 15183
rect -1789 15178 -1778 15183
rect -1837 15175 -1829 15176
rect -1837 15169 -1789 15175
rect -1756 15174 -1740 15183
rect -1837 15159 -1829 15169
rect -1872 15140 -1867 15150
rect -1789 15142 -1781 15149
rect -1776 15142 -1769 15159
rect -1756 15152 -1750 15174
rect -1671 15170 -1669 15181
rect -1663 15178 -1655 15186
rect -1671 15158 -1663 15166
rect -1663 15150 -1655 15158
rect -1702 15140 -1696 15146
rect -1955 15116 -1915 15118
rect -1963 15114 -1955 15116
rect -1963 15107 -1915 15114
rect -1963 15099 -1955 15107
rect -1963 15098 -1915 15099
rect -1973 15092 -1965 15095
rect -1955 15092 -1907 15096
rect -1974 15089 -1907 15092
rect -1973 15085 -1965 15089
rect -1963 15085 -1960 15087
rect -1963 15081 -1915 15085
rect -1963 15073 -1955 15081
rect -1963 15069 -1915 15073
rect -1963 15066 -1955 15069
rect -2240 15059 -2206 15064
rect -2198 15059 -2143 15064
rect -2113 15059 -1981 15064
rect -1915 15059 -1907 15066
rect -2270 15054 -2266 15058
rect -2086 15055 -2070 15059
rect -2325 15046 -2317 15054
rect -2270 15047 -2240 15054
rect -2206 15047 -2176 15054
rect -2325 15026 -2320 15046
rect -2317 15038 -2309 15046
rect -2270 15042 -2266 15047
rect -2270 15038 -2266 15041
rect -2198 15038 -2176 15045
rect -2166 15038 -2158 15055
rect -2143 15047 -2113 15054
rect -2198 15029 -2168 15033
rect -2325 15018 -2317 15026
rect -2143 15024 -2136 15038
rect -2085 15033 -2060 15034
rect -2039 15033 -2035 15042
rect -2135 15026 -2105 15033
rect -2085 15026 -2035 15033
rect -2029 15026 -2025 15033
rect -2325 15005 -2320 15018
rect -2317 15010 -2309 15018
rect -2235 15008 -2232 15011
rect -2325 14979 -2317 15005
rect -2325 14970 -2320 14979
rect -2325 14962 -2317 14970
rect -2135 14962 -2119 14975
rect -2000 14967 -1992 15059
rect -1983 15041 -1981 15059
rect -1955 15041 -1915 15042
rect -1862 15038 -1857 15140
rect -1706 15136 -1702 15140
rect -1829 15124 -1789 15132
rect -1671 15130 -1663 15138
rect -1849 15116 -1842 15124
rect -1790 15116 -1781 15124
rect -1663 15122 -1655 15130
rect -1837 15107 -1829 15114
rect -1758 15107 -1732 15114
rect -1748 15098 -1732 15107
rect -1671 15102 -1663 15110
rect -1829 15089 -1781 15096
rect -1663 15094 -1655 15102
rect -1829 15083 -1789 15087
rect -1768 15084 -1760 15094
rect -1758 15083 -1750 15084
rect -1671 15074 -1663 15082
rect -1837 15071 -1780 15074
rect -1758 15068 -1748 15074
rect -1708 15068 -1690 15074
rect -1829 15059 -1781 15066
rect -1680 15057 -1672 15074
rect -1663 15066 -1655 15074
rect -1829 15048 -1791 15054
rect -1758 15048 -1710 15050
rect -1758 15041 -1692 15048
rect -1671 15046 -1663 15054
rect -1955 15030 -1907 15033
rect -1791 15030 -1781 15033
rect -1991 15026 -1839 15030
rect -1791 15026 -1780 15030
rect -1680 15023 -1672 15041
rect -1663 15038 -1655 15046
rect -1839 15013 -1791 15020
rect -1671 15018 -1663 15026
rect -1829 15007 -1791 15011
rect -1671 15008 -1669 15018
rect -1663 15010 -1655 15018
rect -1680 14992 -1672 15007
rect -1642 14992 -1637 15302
rect -1619 15252 -1614 15468
rect -1619 15226 -1611 15252
rect -1768 14976 -1760 14986
rect -1758 14969 -1710 14976
rect -2325 14942 -2320 14962
rect -2317 14954 -2306 14962
rect -2031 14959 -1992 14967
rect -1750 14965 -1710 14969
rect -1674 14964 -1663 14970
rect -2307 14946 -2306 14954
rect -2149 14957 -2135 14958
rect -2149 14953 -2119 14957
rect -2024 14948 -2021 14957
rect -2325 14934 -2317 14942
rect -2325 14886 -2320 14934
rect -2317 14926 -2306 14934
rect -2185 14932 -2169 14944
rect -2056 14941 -2040 14945
rect -2021 14941 -2008 14948
rect -2056 14930 -2054 14940
rect -2056 14929 -2048 14930
rect -2307 14890 -2306 14898
rect -2111 14897 -2054 14903
rect -2325 14878 -2314 14886
rect -2104 14879 -2101 14883
rect -2325 14858 -2320 14878
rect -2314 14870 -2306 14878
rect -2104 14876 -2101 14878
rect -2084 14876 -2054 14877
rect -2000 14876 -1992 14959
rect -1758 14958 -1750 14959
rect -1758 14957 -1749 14958
rect -1758 14956 -1710 14957
rect -1663 14954 -1658 14964
rect -1831 14946 -1783 14950
rect -1784 14933 -1783 14946
rect -1674 14936 -1663 14942
rect -1826 14931 -1796 14932
rect -1663 14926 -1658 14936
rect -1654 14932 -1647 14942
rect -1644 14918 -1637 14932
rect -1758 14900 -1750 14903
rect -1758 14897 -1710 14900
rect -1844 14885 -1828 14887
rect -1844 14884 -1792 14885
rect -1828 14883 -1792 14884
rect -1772 14883 -1758 14891
rect -1750 14888 -1702 14895
rect -1750 14880 -1710 14884
rect -1700 14880 -1692 14900
rect -1674 14892 -1665 14900
rect -1674 14880 -1666 14888
rect -1758 14876 -1710 14877
rect -2307 14862 -2306 14870
rect -2139 14866 -2123 14875
rect -2111 14870 -2016 14876
rect -2139 14859 -2111 14866
rect -2325 14850 -2314 14858
rect -2177 14852 -2161 14853
rect -2141 14852 -2119 14854
rect -2104 14852 -2101 14870
rect -2076 14859 -2046 14864
rect -2325 14842 -2320 14850
rect -2314 14842 -2306 14850
rect -2076 14848 -2054 14854
rect -2021 14851 -2016 14870
rect -2000 14870 -1818 14876
rect -1802 14870 -1776 14876
rect -1760 14870 -1710 14876
rect -1666 14872 -1658 14880
rect -2189 14842 -2175 14847
rect -2373 14840 -2175 14842
rect -2373 14839 -2359 14840
rect -2371 14702 -2366 14839
rect -2348 14787 -2343 14840
rect -2325 14830 -2320 14840
rect -2307 14834 -2306 14840
rect -2189 14839 -2175 14840
rect -2149 14838 -2119 14847
rect -2084 14846 -2036 14847
rect -2000 14846 -1992 14870
rect -1758 14868 -1710 14870
rect -1758 14866 -1755 14868
rect -1828 14859 -1792 14866
rect -1768 14857 -1760 14864
rect -1758 14859 -1757 14866
rect -1710 14865 -1702 14866
rect -1750 14859 -1702 14865
rect -1674 14864 -1665 14872
rect -1768 14854 -1764 14857
rect -1758 14854 -1755 14859
rect -1818 14846 -1789 14854
rect -1758 14847 -1754 14854
rect -1750 14849 -1710 14854
rect -1674 14852 -1666 14860
rect -1758 14846 -1692 14847
rect -2084 14844 -1692 14846
rect -1666 14844 -1658 14852
rect -2084 14841 -1690 14844
rect -2084 14838 -2054 14841
rect -2046 14839 -1710 14841
rect -2325 14822 -2314 14830
rect -2076 14829 -2046 14836
rect -2325 14802 -2320 14822
rect -2314 14814 -2306 14822
rect -2076 14821 -2054 14827
rect -2084 14817 -2054 14819
rect -2104 14814 -2054 14817
rect -2307 14806 -2306 14814
rect -2084 14811 -2054 14814
rect -2325 14788 -2314 14802
rect -2348 14763 -2341 14787
rect -2325 14772 -2320 14788
rect -2314 14786 -2309 14788
rect -2309 14774 -2298 14786
rect -2092 14783 -2060 14784
rect -2062 14778 -2060 14783
rect -2314 14772 -2309 14774
rect -2348 14702 -2343 14763
rect -2325 14760 -2314 14772
rect -2076 14768 -2062 14778
rect -2076 14762 -2046 14766
rect -2014 14765 -2003 14774
rect -2062 14760 -2046 14762
rect -2325 14744 -2320 14760
rect -2314 14758 -2309 14760
rect -2076 14759 -2062 14760
rect -2309 14746 -2298 14758
rect -2092 14753 -2076 14759
rect -2046 14753 -2026 14754
rect -2314 14744 -2309 14746
rect -2046 14744 -2042 14745
rect -2325 14732 -2314 14744
rect -2141 14740 -2134 14742
rect -2052 14740 -2046 14744
rect -2292 14735 -2111 14740
rect -2096 14738 -2046 14740
rect -2076 14735 -2046 14738
rect -2325 14702 -2320 14732
rect -2314 14730 -2309 14732
rect -2092 14718 -2062 14720
rect -2094 14714 -2062 14718
rect -2000 14702 -1992 14839
rect -1758 14838 -1710 14839
rect -1680 14836 -1665 14844
rect -1750 14829 -1702 14836
rect -1680 14832 -1672 14836
rect -1680 14827 -1666 14832
rect -1836 14823 -1820 14824
rect -1837 14819 -1820 14823
rect -1750 14821 -1710 14827
rect -1674 14824 -1666 14827
rect -1837 14812 -1789 14819
rect -1758 14818 -1710 14819
rect -1760 14815 -1692 14818
rect -1666 14816 -1658 14824
rect -1837 14811 -1820 14812
rect -1764 14811 -1692 14815
rect -1674 14811 -1665 14816
rect -1680 14808 -1665 14811
rect -1750 14792 -1702 14794
rect -1680 14784 -1672 14808
rect -1671 14788 -1666 14804
rect -1854 14783 -1806 14784
rect -1829 14768 -1806 14778
rect -1655 14776 -1650 14788
rect -1666 14772 -1655 14776
rect -1829 14762 -1798 14766
rect -1680 14765 -1672 14768
rect -1806 14760 -1798 14762
rect -1671 14760 -1666 14772
rect -1829 14759 -1806 14760
rect -1854 14757 -1829 14759
rect -1854 14753 -1806 14757
rect -1829 14741 -1806 14751
rect -1655 14748 -1650 14760
rect -1666 14744 -1655 14748
rect -1829 14735 -1680 14740
rect -1671 14732 -1666 14744
rect -1854 14718 -1806 14720
rect -1854 14714 -1680 14718
rect -1642 14702 -1637 14918
rect -1619 14916 -1614 15226
rect -1619 14842 -1612 14866
rect -1619 14702 -1614 14842
rect -1530 14702 -1526 15468
rect -1506 14702 -1502 15468
rect -1499 15467 -1485 15468
rect -1482 15467 -1475 15491
rect -1482 14702 -1478 15467
rect -1458 14702 -1454 15492
rect -1434 14702 -1430 15492
rect -1410 14702 -1406 15492
rect -1386 14702 -1382 15492
rect -1362 14702 -1358 15492
rect -1338 14702 -1334 15492
rect -1314 14702 -1310 15492
rect -1290 14702 -1286 15492
rect -1266 14702 -1262 15492
rect -1242 14702 -1238 15492
rect -1218 14702 -1214 15492
rect -1194 14702 -1190 15492
rect -1170 14702 -1166 15492
rect -1146 14702 -1142 15492
rect -1122 14702 -1118 15492
rect -1098 14702 -1094 15492
rect -1074 14702 -1070 15492
rect -1050 14702 -1046 15492
rect -1026 14702 -1022 15492
rect -1002 14702 -998 15492
rect -978 14702 -974 15492
rect -954 14702 -950 15492
rect -930 14702 -926 15492
rect -906 14702 -902 15492
rect -882 14702 -878 15492
rect -858 14702 -854 15492
rect -845 15461 -840 15471
rect -834 15461 -830 15492
rect -835 15447 -830 15461
rect -834 14702 -830 15447
rect -810 15395 -806 15492
rect -810 15371 -803 15395
rect -810 14702 -806 15371
rect -786 14702 -782 15492
rect -762 14702 -758 15492
rect -749 15317 -744 15327
rect -738 15317 -734 15492
rect -739 15303 -734 15317
rect -738 14702 -734 15303
rect -714 15251 -710 15492
rect -714 15227 -707 15251
rect -714 14702 -710 15227
rect -690 14702 -686 15492
rect -666 14702 -662 15492
rect -642 14702 -638 15492
rect -618 14702 -614 15492
rect -594 14702 -590 15492
rect -570 14702 -566 15492
rect -546 14702 -542 15492
rect -522 14702 -518 15492
rect -498 14702 -494 15492
rect -474 14702 -470 15492
rect -450 14702 -446 15492
rect -426 14702 -422 15492
rect -402 14702 -398 15492
rect -378 14702 -374 15492
rect -354 14702 -350 15492
rect -330 14702 -326 15492
rect -306 14702 -302 15492
rect -293 14741 -288 14751
rect -282 14741 -278 15492
rect -283 14727 -278 14741
rect -293 14717 -288 14727
rect -283 14703 -278 14717
rect -282 14702 -278 14703
rect -258 14702 -254 15492
rect -234 14702 -230 15492
rect -210 14702 -206 15492
rect -186 14702 -182 15492
rect -179 15491 -165 15492
rect -162 15467 -155 15515
rect -162 14702 -158 15467
rect -138 14702 -134 15564
rect -114 14702 -110 15564
rect -90 14702 -86 15564
rect -66 14702 -62 15564
rect -42 14702 -38 15564
rect -18 14702 -14 15564
rect 6 14702 10 15564
rect 30 14702 34 15564
rect 54 14702 58 15564
rect 78 14702 82 15564
rect 102 14702 106 15564
rect 126 14702 130 15564
rect 150 14702 154 15564
rect 174 14702 178 15564
rect 198 14702 202 15564
rect 222 14702 226 15564
rect 246 14702 250 15564
rect 270 14702 274 15564
rect 294 14702 298 15564
rect 307 15269 312 15279
rect 318 15269 322 15564
rect 317 15255 322 15269
rect 318 14702 322 15255
rect 342 15203 346 15564
rect 342 15179 349 15203
rect 342 14702 346 15179
rect 366 14702 370 15564
rect 390 14702 394 15564
rect 414 14702 418 15564
rect 438 14702 442 15564
rect 462 14702 466 15564
rect 486 14702 490 15564
rect 510 14702 514 15564
rect 534 14702 538 15564
rect 558 14702 562 15564
rect 582 14702 586 15564
rect 606 14702 610 15564
rect 630 14702 634 15564
rect 654 14702 658 15564
rect 678 14702 682 15564
rect 702 14702 706 15564
rect 726 14702 730 15564
rect 750 14702 754 15564
rect 774 14702 778 15564
rect 798 14702 802 15564
rect 822 14702 826 15564
rect 846 14702 850 15564
rect 870 14702 874 15564
rect 894 14702 898 15564
rect 918 14702 922 15564
rect 942 14702 946 15564
rect 966 14702 970 15564
rect 990 14702 994 15564
rect 1014 14702 1018 15564
rect 1038 14702 1042 15564
rect 1062 14702 1066 15564
rect 1086 14702 1090 15564
rect 1110 14702 1114 15564
rect 1134 14702 1138 15564
rect 1158 14702 1162 15564
rect 1182 14702 1186 15564
rect 1206 14702 1210 15564
rect 1230 14702 1234 15564
rect 1254 14702 1258 15564
rect 1278 14702 1282 15564
rect 1302 14702 1306 15564
rect 1326 14702 1330 15564
rect 1350 14702 1354 15564
rect 1374 14702 1378 15564
rect 1398 14702 1402 15564
rect 1422 14702 1426 15564
rect 1446 14702 1450 15564
rect 1470 14702 1474 15564
rect 1494 14702 1498 15564
rect 1518 14702 1522 15564
rect 1542 14702 1546 15564
rect 1566 14702 1570 15564
rect 1590 14702 1594 15564
rect 1614 14702 1618 15564
rect 1638 14702 1642 15564
rect 1662 14702 1666 15564
rect 1686 14702 1690 15564
rect 1710 14702 1714 15564
rect 1734 14702 1738 15564
rect 1758 14702 1762 15564
rect 1782 14702 1786 15564
rect 1806 14702 1810 15564
rect 1830 14702 1834 15564
rect 1854 14702 1858 15564
rect 1878 14702 1882 15564
rect 1902 14702 1906 15564
rect 1926 14702 1930 15564
rect 1950 14702 1954 15564
rect 1974 14702 1978 15564
rect 1998 14702 2002 15564
rect 2011 14909 2016 14919
rect 2022 14909 2026 15564
rect 2035 15485 2040 15495
rect 2046 15485 2050 15564
rect 2045 15471 2050 15485
rect 2021 14895 2026 14909
rect 2011 14885 2016 14895
rect 2021 14871 2026 14885
rect 2022 14702 2026 14871
rect 2046 14843 2050 15471
rect 2070 15419 2074 15564
rect 2070 15395 2077 15419
rect 2046 14798 2053 14843
rect 2070 14798 2074 15395
rect 2094 14798 2098 15564
rect 2118 14798 2122 15564
rect 2142 14798 2146 15564
rect 2166 14798 2170 15564
rect 2190 14798 2194 15564
rect 2214 14798 2218 15564
rect 2238 14798 2242 15564
rect 2262 14798 2266 15564
rect 2286 14798 2290 15564
rect 2310 14798 2314 15564
rect 2334 14798 2338 15564
rect 2358 14798 2362 15564
rect 2382 14798 2386 15564
rect 2406 14798 2410 15564
rect 2430 14798 2434 15564
rect 2454 14798 2458 15564
rect 2478 14798 2482 15564
rect 2502 14798 2506 15564
rect 2526 14798 2530 15564
rect 2550 14798 2554 15564
rect 2574 14798 2578 15564
rect 2598 14798 2602 15564
rect 2622 14798 2626 15564
rect 2646 14798 2650 15564
rect 2670 14798 2674 15564
rect 2694 14798 2698 15564
rect 2718 14798 2722 15564
rect 2742 14798 2746 15564
rect 2766 14798 2770 15564
rect 2790 14798 2794 15564
rect 2814 14798 2818 15564
rect 2838 14798 2842 15564
rect 2862 14798 2866 15564
rect 2886 14798 2890 15564
rect 2910 14798 2914 15564
rect 2934 14798 2938 15564
rect 2958 14798 2962 15564
rect 2982 14798 2986 15564
rect 3006 14798 3010 15564
rect 3030 14798 3034 15564
rect 3054 14798 3058 15564
rect 3078 14798 3082 15564
rect 3102 14798 3106 15564
rect 3126 14798 3130 15564
rect 3150 14798 3154 15564
rect 3174 14798 3178 15564
rect 3198 14798 3202 15564
rect 3222 14798 3226 15564
rect 3246 14798 3250 15564
rect 3270 14798 3274 15564
rect 3294 14798 3298 15564
rect 3318 14798 3322 15564
rect 3342 14798 3346 15564
rect 3366 14798 3370 15564
rect 3390 14798 3394 15564
rect 3414 14798 3418 15564
rect 3438 14798 3442 15564
rect 3462 14798 3466 15564
rect 3486 14798 3490 15564
rect 3510 14798 3514 15564
rect 3534 14798 3538 15564
rect 3558 14798 3562 15564
rect 3582 14798 3586 15564
rect 3606 14798 3610 15564
rect 3619 15557 3624 15564
rect 3630 15557 3634 15564
rect 3629 15543 3634 15557
rect 3619 15509 3624 15519
rect 3629 15495 3634 15509
rect 3619 14885 3624 14895
rect 3630 14885 3634 15495
rect 3629 14871 3634 14885
rect 3619 14798 3651 14799
rect 2029 14796 3651 14798
rect 2029 14795 2043 14796
rect 2046 14795 2053 14796
rect 2035 14765 2040 14775
rect 2046 14765 2050 14795
rect 2045 14751 2050 14765
rect 2046 14702 2050 14751
rect 2070 14702 2074 14796
rect 2094 14702 2098 14796
rect 2118 14702 2122 14796
rect 2142 14702 2146 14796
rect 2166 14702 2170 14796
rect 2190 14702 2194 14796
rect 2214 14702 2218 14796
rect 2238 14702 2242 14796
rect 2262 14702 2266 14796
rect 2286 14702 2290 14796
rect 2310 14702 2314 14796
rect 2334 14702 2338 14796
rect 2358 14702 2362 14796
rect 2382 14702 2386 14796
rect 2406 14702 2410 14796
rect 2430 14702 2434 14796
rect 2454 14702 2458 14796
rect 2478 14702 2482 14796
rect 2502 14702 2506 14796
rect 2526 14702 2530 14796
rect 2550 14702 2554 14796
rect 2574 14702 2578 14796
rect 2598 14702 2602 14796
rect 2622 14702 2626 14796
rect 2646 14702 2650 14796
rect 2670 14702 2674 14796
rect 2694 14702 2698 14796
rect 2718 14702 2722 14796
rect 2742 14702 2746 14796
rect 2766 14702 2770 14796
rect 2790 14702 2794 14796
rect 2814 14702 2818 14796
rect 2838 14702 2842 14796
rect 2862 14702 2866 14796
rect 2886 14702 2890 14796
rect 2910 14702 2914 14796
rect 2934 14702 2938 14796
rect 2958 14702 2962 14796
rect 2982 14702 2986 14796
rect 3006 14702 3010 14796
rect 3030 14702 3034 14796
rect 3054 14702 3058 14796
rect 3078 14702 3082 14796
rect 3102 14702 3106 14796
rect 3126 14702 3130 14796
rect 3150 14702 3154 14796
rect 3174 14702 3178 14796
rect 3198 14702 3202 14796
rect 3222 14702 3226 14796
rect 3246 14702 3250 14796
rect 3270 14702 3274 14796
rect 3294 14702 3298 14796
rect 3318 14702 3322 14796
rect 3342 14702 3346 14796
rect 3366 14702 3370 14796
rect 3390 14702 3394 14796
rect 3414 14702 3418 14796
rect 3438 14702 3442 14796
rect 3462 14702 3466 14796
rect 3486 14702 3490 14796
rect 3510 14702 3514 14796
rect 3534 14702 3538 14796
rect 3558 14702 3562 14796
rect 3582 14702 3586 14796
rect 3606 14702 3610 14796
rect 3619 14789 3624 14796
rect 3637 14795 3651 14796
rect 3629 14775 3634 14789
rect 3619 14717 3624 14727
rect 3630 14717 3634 14775
rect 3629 14703 3634 14717
rect 3643 14713 3651 14717
rect 3637 14703 3643 14713
rect 3619 14702 3651 14703
rect -2393 14700 3651 14702
rect -2371 14678 -2366 14700
rect -2348 14678 -2343 14700
rect -2325 14678 -2320 14700
rect -2072 14698 -2036 14699
rect -2072 14692 -2054 14698
rect -2309 14684 -2301 14692
rect -2317 14678 -2309 14684
rect -2092 14683 -2062 14688
rect -2000 14679 -1992 14700
rect -1938 14699 -1906 14700
rect -1920 14698 -1906 14699
rect -1806 14692 -1680 14698
rect -1854 14683 -1806 14688
rect -1655 14684 -1647 14692
rect -1982 14679 -1966 14680
rect -2000 14678 -1966 14679
rect -1846 14678 -1806 14681
rect -1663 14678 -1655 14684
rect -1642 14678 -1637 14700
rect -1619 14678 -1614 14700
rect -1530 14678 -1526 14700
rect -1506 14678 -1502 14700
rect -1482 14678 -1478 14700
rect -1458 14678 -1454 14700
rect -1434 14678 -1430 14700
rect -1410 14678 -1406 14700
rect -1386 14678 -1382 14700
rect -1362 14678 -1358 14700
rect -1338 14678 -1334 14700
rect -1314 14678 -1310 14700
rect -1290 14678 -1286 14700
rect -1266 14678 -1262 14700
rect -1242 14678 -1238 14700
rect -1218 14678 -1214 14700
rect -1194 14678 -1190 14700
rect -1170 14678 -1166 14700
rect -1146 14678 -1142 14700
rect -1122 14678 -1118 14700
rect -1098 14678 -1094 14700
rect -1074 14678 -1070 14700
rect -1050 14678 -1046 14700
rect -1026 14678 -1022 14700
rect -1002 14678 -998 14700
rect -978 14678 -974 14700
rect -954 14678 -950 14700
rect -930 14678 -926 14700
rect -906 14678 -902 14700
rect -882 14678 -878 14700
rect -858 14678 -854 14700
rect -834 14678 -830 14700
rect -810 14678 -806 14700
rect -786 14678 -782 14700
rect -762 14678 -758 14700
rect -738 14678 -734 14700
rect -714 14678 -710 14700
rect -690 14678 -686 14700
rect -666 14678 -662 14700
rect -642 14678 -638 14700
rect -618 14678 -614 14700
rect -594 14678 -590 14700
rect -570 14678 -566 14700
rect -546 14678 -542 14700
rect -522 14678 -518 14700
rect -498 14678 -494 14700
rect -474 14678 -470 14700
rect -450 14678 -446 14700
rect -426 14678 -422 14700
rect -402 14678 -398 14700
rect -378 14678 -374 14700
rect -354 14678 -350 14700
rect -330 14678 -326 14700
rect -306 14678 -302 14700
rect -282 14678 -278 14700
rect -258 14678 -254 14700
rect -234 14678 -230 14700
rect -210 14678 -206 14700
rect -186 14678 -182 14700
rect -162 14678 -158 14700
rect -138 14678 -134 14700
rect -114 14678 -110 14700
rect -90 14678 -86 14700
rect -66 14678 -62 14700
rect -42 14678 -38 14700
rect -18 14678 -14 14700
rect 6 14678 10 14700
rect 30 14678 34 14700
rect 54 14678 58 14700
rect 78 14678 82 14700
rect 102 14678 106 14700
rect 126 14678 130 14700
rect 150 14678 154 14700
rect 174 14678 178 14700
rect 198 14678 202 14700
rect 222 14678 226 14700
rect 246 14678 250 14700
rect 270 14678 274 14700
rect 294 14678 298 14700
rect 318 14678 322 14700
rect 342 14678 346 14700
rect 366 14678 370 14700
rect 390 14678 394 14700
rect 414 14678 418 14700
rect 438 14678 442 14700
rect 462 14678 466 14700
rect 486 14678 490 14700
rect 510 14678 514 14700
rect 534 14678 538 14700
rect 558 14678 562 14700
rect 582 14678 586 14700
rect 606 14678 610 14700
rect 630 14678 634 14700
rect 654 14678 658 14700
rect 678 14678 682 14700
rect 702 14678 706 14700
rect 726 14678 730 14700
rect 750 14678 754 14700
rect 774 14678 778 14700
rect 798 14678 802 14700
rect 822 14678 826 14700
rect 846 14678 850 14700
rect 870 14678 874 14700
rect 894 14678 898 14700
rect 918 14678 922 14700
rect 942 14678 946 14700
rect 966 14678 970 14700
rect 990 14678 994 14700
rect 1014 14678 1018 14700
rect 1038 14678 1042 14700
rect 1062 14678 1066 14700
rect 1086 14678 1090 14700
rect 1110 14678 1114 14700
rect 1134 14678 1138 14700
rect 1158 14678 1162 14700
rect 1182 14678 1186 14700
rect 1206 14678 1210 14700
rect 1230 14678 1234 14700
rect 1254 14678 1258 14700
rect 1278 14678 1282 14700
rect 1302 14678 1306 14700
rect 1326 14678 1330 14700
rect 1350 14678 1354 14700
rect 1374 14678 1378 14700
rect 1398 14678 1402 14700
rect 1422 14678 1426 14700
rect 1446 14678 1450 14700
rect 1470 14678 1474 14700
rect 1494 14678 1498 14700
rect 1518 14678 1522 14700
rect 1542 14678 1546 14700
rect 1566 14678 1570 14700
rect 1590 14678 1594 14700
rect 1614 14678 1618 14700
rect 1638 14678 1642 14700
rect 1662 14678 1666 14700
rect 1686 14678 1690 14700
rect 1710 14678 1714 14700
rect 1734 14678 1738 14700
rect 1758 14678 1762 14700
rect 1782 14678 1786 14700
rect 1806 14678 1810 14700
rect 1830 14678 1834 14700
rect 1854 14678 1858 14700
rect 1878 14679 1882 14700
rect 1867 14678 1901 14679
rect -2393 14676 1901 14678
rect -2371 14654 -2366 14676
rect -2348 14654 -2343 14676
rect -2325 14654 -2320 14676
rect -2000 14674 -1966 14676
rect -2309 14656 -2301 14664
rect -2062 14663 -2054 14670
rect -2092 14656 -2084 14663
rect -2062 14656 -2026 14658
rect -2317 14654 -2309 14656
rect -2062 14654 -2012 14656
rect -2000 14654 -1992 14674
rect -1982 14673 -1966 14674
rect -1846 14672 -1806 14676
rect -1846 14665 -1798 14670
rect -1806 14663 -1798 14665
rect -1854 14661 -1846 14663
rect -1854 14656 -1806 14661
rect -1655 14656 -1647 14664
rect -1864 14654 -1796 14655
rect -1663 14654 -1655 14656
rect -1642 14654 -1637 14676
rect -1619 14654 -1614 14676
rect -1530 14654 -1526 14676
rect -1506 14654 -1502 14676
rect -1482 14654 -1478 14676
rect -1458 14654 -1454 14676
rect -1434 14654 -1430 14676
rect -1410 14654 -1406 14676
rect -1386 14654 -1382 14676
rect -1362 14654 -1358 14676
rect -1338 14654 -1334 14676
rect -1314 14654 -1310 14676
rect -1290 14654 -1286 14676
rect -1266 14654 -1262 14676
rect -1242 14654 -1238 14676
rect -1218 14654 -1214 14676
rect -1194 14654 -1190 14676
rect -1170 14654 -1166 14676
rect -1146 14654 -1142 14676
rect -1122 14654 -1118 14676
rect -1098 14654 -1094 14676
rect -1074 14654 -1070 14676
rect -1050 14654 -1046 14676
rect -1026 14654 -1022 14676
rect -1002 14654 -998 14676
rect -978 14654 -974 14676
rect -954 14654 -950 14676
rect -930 14654 -926 14676
rect -906 14654 -902 14676
rect -882 14654 -878 14676
rect -858 14654 -854 14676
rect -834 14654 -830 14676
rect -810 14654 -806 14676
rect -786 14654 -782 14676
rect -762 14654 -758 14676
rect -738 14654 -734 14676
rect -714 14654 -710 14676
rect -690 14654 -686 14676
rect -666 14654 -662 14676
rect -642 14654 -638 14676
rect -618 14654 -614 14676
rect -594 14654 -590 14676
rect -570 14654 -566 14676
rect -546 14654 -542 14676
rect -522 14654 -518 14676
rect -498 14654 -494 14676
rect -474 14654 -470 14676
rect -450 14654 -446 14676
rect -426 14654 -422 14676
rect -402 14654 -398 14676
rect -378 14654 -374 14676
rect -354 14654 -350 14676
rect -330 14654 -326 14676
rect -306 14654 -302 14676
rect -282 14654 -278 14676
rect -258 14675 -254 14676
rect -2393 14652 -261 14654
rect -2371 14606 -2366 14652
rect -2348 14606 -2343 14652
rect -2325 14606 -2320 14652
rect -2317 14648 -2309 14652
rect -2062 14648 -2054 14652
rect -2154 14644 -2138 14646
rect -2057 14644 -2054 14648
rect -2292 14638 -2054 14644
rect -2052 14638 -2044 14648
rect -2092 14622 -2062 14624
rect -2094 14618 -2062 14622
rect -2000 14606 -1992 14652
rect -1846 14645 -1806 14652
rect -1663 14648 -1655 14652
rect -1846 14638 -1680 14644
rect -1854 14622 -1806 14624
rect -1854 14618 -1680 14622
rect -1979 14606 -1945 14608
rect -1642 14606 -1637 14652
rect -1619 14606 -1614 14652
rect -1530 14606 -1526 14652
rect -1506 14606 -1502 14652
rect -1482 14606 -1478 14652
rect -1458 14606 -1454 14652
rect -1434 14606 -1430 14652
rect -1410 14606 -1406 14652
rect -1386 14606 -1382 14652
rect -1362 14606 -1358 14652
rect -1338 14606 -1334 14652
rect -1314 14606 -1310 14652
rect -1290 14606 -1286 14652
rect -1266 14606 -1262 14652
rect -1242 14606 -1238 14652
rect -1218 14606 -1214 14652
rect -1194 14606 -1190 14652
rect -1170 14606 -1166 14652
rect -1146 14606 -1142 14652
rect -1122 14606 -1118 14652
rect -1098 14606 -1094 14652
rect -1074 14606 -1070 14652
rect -1050 14606 -1046 14652
rect -1026 14606 -1022 14652
rect -1002 14606 -998 14652
rect -978 14606 -974 14652
rect -954 14606 -950 14652
rect -930 14606 -926 14652
rect -906 14606 -902 14652
rect -882 14606 -878 14652
rect -858 14606 -854 14652
rect -834 14606 -830 14652
rect -810 14606 -806 14652
rect -786 14606 -782 14652
rect -762 14606 -758 14652
rect -738 14606 -734 14652
rect -714 14606 -710 14652
rect -690 14606 -686 14652
rect -666 14606 -662 14652
rect -642 14606 -638 14652
rect -618 14606 -614 14652
rect -594 14606 -590 14652
rect -570 14606 -566 14652
rect -546 14606 -542 14652
rect -522 14606 -518 14652
rect -498 14606 -494 14652
rect -474 14606 -470 14652
rect -450 14606 -446 14652
rect -426 14606 -422 14652
rect -402 14606 -398 14652
rect -378 14606 -374 14652
rect -354 14606 -350 14652
rect -330 14606 -326 14652
rect -306 14606 -302 14652
rect -282 14606 -278 14652
rect -275 14651 -261 14652
rect -258 14627 -251 14675
rect -258 14606 -254 14627
rect -234 14606 -230 14676
rect -210 14606 -206 14676
rect -186 14606 -182 14676
rect -162 14606 -158 14676
rect -138 14606 -134 14676
rect -114 14606 -110 14676
rect -90 14606 -86 14676
rect -66 14606 -62 14676
rect -42 14606 -38 14676
rect -18 14606 -14 14676
rect 6 14606 10 14676
rect 30 14606 34 14676
rect 54 14606 58 14676
rect 78 14606 82 14676
rect 102 14606 106 14676
rect 126 14606 130 14676
rect 150 14606 154 14676
rect 174 14606 178 14676
rect 198 14606 202 14676
rect 222 14606 226 14676
rect 246 14606 250 14676
rect 270 14606 274 14676
rect 294 14606 298 14676
rect 318 14606 322 14676
rect 342 14606 346 14676
rect 366 14606 370 14676
rect 390 14606 394 14676
rect 414 14606 418 14676
rect 438 14606 442 14676
rect 462 14606 466 14676
rect 486 14606 490 14676
rect 510 14606 514 14676
rect 534 14606 538 14676
rect 558 14606 562 14676
rect 582 14606 586 14676
rect 606 14606 610 14676
rect 630 14606 634 14676
rect 654 14606 658 14676
rect 678 14606 682 14676
rect 702 14606 706 14676
rect 726 14606 730 14676
rect 750 14606 754 14676
rect 774 14606 778 14676
rect 798 14606 802 14676
rect 822 14606 826 14676
rect 846 14606 850 14676
rect 870 14606 874 14676
rect 894 14606 898 14676
rect 918 14606 922 14676
rect 942 14606 946 14676
rect 966 14606 970 14676
rect 990 14606 994 14676
rect 1014 14606 1018 14676
rect 1038 14606 1042 14676
rect 1062 14606 1066 14676
rect 1086 14606 1090 14676
rect 1110 14606 1114 14676
rect 1123 14645 1128 14655
rect 1134 14645 1138 14676
rect 1133 14631 1138 14645
rect 1123 14630 1157 14631
rect 1158 14630 1162 14676
rect 1182 14630 1186 14676
rect 1206 14630 1210 14676
rect 1230 14630 1234 14676
rect 1254 14630 1258 14676
rect 1278 14630 1282 14676
rect 1302 14630 1306 14676
rect 1326 14630 1330 14676
rect 1350 14630 1354 14676
rect 1374 14630 1378 14676
rect 1398 14630 1402 14676
rect 1422 14630 1426 14676
rect 1446 14630 1450 14676
rect 1470 14630 1474 14676
rect 1494 14630 1498 14676
rect 1518 14630 1522 14676
rect 1542 14630 1546 14676
rect 1566 14630 1570 14676
rect 1590 14630 1594 14676
rect 1614 14630 1618 14676
rect 1638 14630 1642 14676
rect 1662 14630 1666 14676
rect 1686 14630 1690 14676
rect 1710 14630 1714 14676
rect 1734 14630 1738 14676
rect 1758 14630 1762 14676
rect 1782 14630 1786 14676
rect 1806 14630 1810 14676
rect 1830 14630 1834 14676
rect 1854 14630 1858 14676
rect 1867 14669 1872 14676
rect 1878 14669 1882 14676
rect 1877 14655 1882 14669
rect 1878 14630 1882 14655
rect 1902 14630 1906 14700
rect 1926 14630 1930 14700
rect 1950 14630 1954 14700
rect 1974 14630 1978 14700
rect 1998 14630 2002 14700
rect 2022 14630 2026 14700
rect 2046 14630 2050 14700
rect 2070 14699 2074 14700
rect 2070 14675 2077 14699
rect 2070 14630 2074 14675
rect 2094 14630 2098 14700
rect 2118 14630 2122 14700
rect 2142 14630 2146 14700
rect 2166 14630 2170 14700
rect 2190 14630 2194 14700
rect 2214 14630 2218 14700
rect 2238 14630 2242 14700
rect 2262 14630 2266 14700
rect 2286 14630 2290 14700
rect 2310 14630 2314 14700
rect 2334 14630 2338 14700
rect 2358 14630 2362 14700
rect 2382 14630 2386 14700
rect 2406 14630 2410 14700
rect 2430 14630 2434 14700
rect 2454 14630 2458 14700
rect 2478 14630 2482 14700
rect 2502 14630 2506 14700
rect 2526 14630 2530 14700
rect 2550 14630 2554 14700
rect 2574 14630 2578 14700
rect 2598 14630 2602 14700
rect 2622 14630 2626 14700
rect 2646 14630 2650 14700
rect 2670 14630 2674 14700
rect 2694 14630 2698 14700
rect 2718 14630 2722 14700
rect 2742 14630 2746 14700
rect 2766 14630 2770 14700
rect 2790 14630 2794 14700
rect 2814 14630 2818 14700
rect 2838 14630 2842 14700
rect 2862 14630 2866 14700
rect 2886 14630 2890 14700
rect 2910 14630 2914 14700
rect 2934 14630 2938 14700
rect 2958 14630 2962 14700
rect 2982 14630 2986 14700
rect 3006 14630 3010 14700
rect 3030 14630 3034 14700
rect 3054 14630 3058 14700
rect 3078 14630 3082 14700
rect 3102 14630 3106 14700
rect 3126 14630 3130 14700
rect 3150 14630 3154 14700
rect 3174 14630 3178 14700
rect 3198 14630 3202 14700
rect 3222 14630 3226 14700
rect 3246 14630 3250 14700
rect 3270 14630 3274 14700
rect 3294 14630 3298 14700
rect 3318 14630 3322 14700
rect 3342 14630 3346 14700
rect 3366 14630 3370 14700
rect 3390 14630 3394 14700
rect 3414 14630 3418 14700
rect 3438 14630 3442 14700
rect 3462 14630 3466 14700
rect 3486 14630 3490 14700
rect 3510 14630 3514 14700
rect 3534 14630 3538 14700
rect 3558 14630 3562 14700
rect 3582 14630 3586 14700
rect 3606 14630 3610 14700
rect 3619 14693 3624 14700
rect 3637 14699 3651 14700
rect 3629 14679 3634 14693
rect 3630 14631 3634 14679
rect 3619 14630 3651 14631
rect 1123 14628 3651 14630
rect 1123 14621 1128 14628
rect 1133 14607 1138 14621
rect 1134 14606 1138 14607
rect 1158 14606 1162 14628
rect 1182 14606 1186 14628
rect 1206 14606 1210 14628
rect 1230 14606 1234 14628
rect 1254 14606 1258 14628
rect 1278 14606 1282 14628
rect 1302 14606 1306 14628
rect 1326 14606 1330 14628
rect 1350 14606 1354 14628
rect 1374 14606 1378 14628
rect 1398 14606 1402 14628
rect 1422 14606 1426 14628
rect 1446 14606 1450 14628
rect 1470 14606 1474 14628
rect 1494 14606 1498 14628
rect 1518 14606 1522 14628
rect 1542 14606 1546 14628
rect 1566 14606 1570 14628
rect 1590 14606 1594 14628
rect 1614 14606 1618 14628
rect 1638 14606 1642 14628
rect 1662 14606 1666 14628
rect 1686 14606 1690 14628
rect 1710 14606 1714 14628
rect 1734 14606 1738 14628
rect 1758 14606 1762 14628
rect 1782 14606 1786 14628
rect 1806 14606 1810 14628
rect 1830 14606 1834 14628
rect 1854 14606 1858 14628
rect 1878 14606 1882 14628
rect 1902 14606 1906 14628
rect 1926 14606 1930 14628
rect 1950 14606 1954 14628
rect 1974 14606 1978 14628
rect 1998 14606 2002 14628
rect 2022 14606 2026 14628
rect 2046 14606 2050 14628
rect 2070 14606 2074 14628
rect 2094 14606 2098 14628
rect 2118 14606 2122 14628
rect 2142 14606 2146 14628
rect 2166 14606 2170 14628
rect 2190 14606 2194 14628
rect 2214 14606 2218 14628
rect 2238 14606 2242 14628
rect 2262 14606 2266 14628
rect 2286 14606 2290 14628
rect 2310 14606 2314 14628
rect 2334 14606 2338 14628
rect 2358 14606 2362 14628
rect 2382 14606 2386 14628
rect 2406 14606 2410 14628
rect 2430 14606 2434 14628
rect 2454 14606 2458 14628
rect 2478 14606 2482 14628
rect 2502 14606 2506 14628
rect 2526 14606 2530 14628
rect 2550 14606 2554 14628
rect 2574 14606 2578 14628
rect 2598 14606 2602 14628
rect 2622 14606 2626 14628
rect 2646 14606 2650 14628
rect 2670 14606 2674 14628
rect 2694 14606 2698 14628
rect 2718 14606 2722 14628
rect 2742 14606 2746 14628
rect 2766 14606 2770 14628
rect 2790 14606 2794 14628
rect 2814 14606 2818 14628
rect 2838 14606 2842 14628
rect 2862 14606 2866 14628
rect 2886 14606 2890 14628
rect 2910 14606 2914 14628
rect 2934 14606 2938 14628
rect 2958 14606 2962 14628
rect 2982 14606 2986 14628
rect 3006 14606 3010 14628
rect 3030 14606 3034 14628
rect 3054 14606 3058 14628
rect 3078 14606 3082 14628
rect 3102 14606 3106 14628
rect 3126 14606 3130 14628
rect 3150 14606 3154 14628
rect 3174 14606 3178 14628
rect 3198 14606 3202 14628
rect 3222 14606 3226 14628
rect 3246 14606 3250 14628
rect 3270 14606 3274 14628
rect 3294 14606 3298 14628
rect 3318 14606 3322 14628
rect 3342 14606 3346 14628
rect 3366 14606 3370 14628
rect 3390 14606 3394 14628
rect 3414 14606 3418 14628
rect 3438 14606 3442 14628
rect 3462 14606 3466 14628
rect 3486 14606 3490 14628
rect 3510 14606 3514 14628
rect 3534 14606 3538 14628
rect 3558 14606 3562 14628
rect 3582 14606 3586 14628
rect 3606 14606 3610 14628
rect 3619 14621 3624 14628
rect 3630 14621 3634 14628
rect 3637 14627 3651 14628
rect 3629 14607 3634 14621
rect 3643 14617 3651 14621
rect 3637 14607 3643 14617
rect 3619 14606 3651 14607
rect -2393 14604 3651 14606
rect -2371 14558 -2366 14604
rect -2348 14558 -2343 14604
rect -2325 14558 -2320 14604
rect -2080 14603 -1906 14604
rect -2080 14602 -2036 14603
rect -2080 14596 -2054 14602
rect -2309 14588 -2301 14594
rect -2317 14578 -2309 14588
rect -2070 14587 -2040 14594
rect -2054 14579 -2040 14582
rect -2000 14577 -1992 14603
rect -1920 14602 -1906 14603
rect -1850 14596 -1846 14604
rect -1840 14596 -1792 14604
rect -1969 14584 -1966 14593
rect -1850 14589 -1802 14594
rect -1906 14587 -1802 14589
rect -1655 14588 -1647 14594
rect -1906 14586 -1850 14587
rect -1846 14579 -1802 14585
rect -1663 14578 -1655 14588
rect -1860 14577 -1798 14578
rect -2078 14570 -2070 14577
rect -2309 14560 -2301 14566
rect -2317 14558 -2309 14560
rect -2154 14558 -2145 14568
rect -2044 14567 -2040 14572
rect -2028 14570 -1945 14577
rect -1929 14570 -1794 14577
rect -2070 14560 -2040 14567
rect -2044 14558 -2028 14560
rect -2000 14558 -1992 14570
rect -1860 14569 -1798 14570
rect -1850 14560 -1802 14567
rect -1655 14560 -1647 14566
rect -1978 14558 -1942 14559
rect -1663 14558 -1655 14560
rect -1642 14558 -1637 14604
rect -1619 14558 -1614 14604
rect -1530 14558 -1526 14604
rect -1506 14558 -1502 14604
rect -1482 14558 -1478 14604
rect -1458 14558 -1454 14604
rect -1434 14558 -1430 14604
rect -1410 14558 -1406 14604
rect -1386 14558 -1382 14604
rect -1362 14558 -1358 14604
rect -1338 14558 -1334 14604
rect -1314 14558 -1310 14604
rect -1290 14558 -1286 14604
rect -1266 14558 -1262 14604
rect -1242 14558 -1238 14604
rect -1218 14558 -1214 14604
rect -1194 14558 -1190 14604
rect -1170 14558 -1166 14604
rect -1146 14558 -1142 14604
rect -1122 14558 -1118 14604
rect -1098 14558 -1094 14604
rect -1074 14558 -1070 14604
rect -1050 14558 -1046 14604
rect -1026 14558 -1022 14604
rect -1002 14558 -998 14604
rect -978 14558 -974 14604
rect -954 14558 -950 14604
rect -930 14558 -926 14604
rect -906 14558 -902 14604
rect -882 14558 -878 14604
rect -858 14558 -854 14604
rect -834 14558 -830 14604
rect -810 14558 -806 14604
rect -786 14558 -782 14604
rect -762 14558 -758 14604
rect -738 14558 -734 14604
rect -714 14558 -710 14604
rect -690 14558 -686 14604
rect -666 14558 -662 14604
rect -642 14558 -638 14604
rect -618 14558 -614 14604
rect -594 14558 -590 14604
rect -570 14558 -566 14604
rect -546 14558 -542 14604
rect -522 14558 -518 14604
rect -498 14558 -494 14604
rect -474 14558 -470 14604
rect -450 14558 -446 14604
rect -426 14558 -422 14604
rect -402 14558 -398 14604
rect -378 14558 -374 14604
rect -354 14558 -350 14604
rect -330 14558 -326 14604
rect -306 14558 -302 14604
rect -282 14558 -278 14604
rect -258 14558 -254 14604
rect -234 14558 -230 14604
rect -210 14558 -206 14604
rect -186 14558 -182 14604
rect -162 14558 -158 14604
rect -138 14558 -134 14604
rect -114 14558 -110 14604
rect -90 14558 -86 14604
rect -66 14558 -62 14604
rect -42 14558 -38 14604
rect -18 14558 -14 14604
rect 6 14558 10 14604
rect 30 14558 34 14604
rect 54 14558 58 14604
rect 78 14558 82 14604
rect 102 14558 106 14604
rect 126 14558 130 14604
rect 150 14558 154 14604
rect 174 14558 178 14604
rect 198 14558 202 14604
rect 222 14558 226 14604
rect 246 14558 250 14604
rect 270 14558 274 14604
rect 294 14558 298 14604
rect 318 14558 322 14604
rect 342 14558 346 14604
rect 366 14558 370 14604
rect 390 14558 394 14604
rect 414 14558 418 14604
rect 438 14558 442 14604
rect 462 14558 466 14604
rect 486 14558 490 14604
rect 510 14558 514 14604
rect 534 14558 538 14604
rect 558 14558 562 14604
rect 582 14558 586 14604
rect 606 14558 610 14604
rect 630 14558 634 14604
rect 654 14558 658 14604
rect 678 14558 682 14604
rect 702 14558 706 14604
rect 726 14558 730 14604
rect 750 14558 754 14604
rect 774 14558 778 14604
rect 798 14558 802 14604
rect 822 14558 826 14604
rect 846 14558 850 14604
rect 870 14558 874 14604
rect 894 14558 898 14604
rect 918 14558 922 14604
rect 942 14558 946 14604
rect 966 14558 970 14604
rect 990 14558 994 14604
rect 1014 14558 1018 14604
rect 1038 14558 1042 14604
rect 1062 14558 1066 14604
rect 1086 14558 1090 14604
rect 1110 14558 1114 14604
rect 1134 14558 1138 14604
rect 1158 14579 1162 14604
rect -2393 14556 1155 14558
rect -2371 14462 -2366 14556
rect -2348 14462 -2343 14556
rect -2325 14518 -2320 14556
rect -2317 14550 -2309 14556
rect -2145 14552 -2138 14556
rect -2070 14552 -2054 14556
rect -2078 14543 -2054 14550
rect -2062 14518 -2032 14519
rect -2000 14518 -1992 14556
rect -1846 14552 -1802 14556
rect -1846 14542 -1792 14551
rect -1663 14550 -1655 14556
rect -1942 14520 -1937 14532
rect -1850 14529 -1822 14530
rect -1850 14525 -1802 14529
rect -2325 14510 -2317 14518
rect -2062 14516 -1961 14518
rect -2325 14490 -2320 14510
rect -2317 14502 -2309 14510
rect -2062 14503 -2040 14514
rect -2032 14509 -1961 14516
rect -1947 14510 -1942 14518
rect -1842 14516 -1794 14519
rect -2070 14498 -2022 14502
rect -2325 14476 -2317 14490
rect -2072 14482 -2032 14483
rect -2102 14476 -2032 14482
rect -2325 14462 -2320 14476
rect -2317 14474 -2309 14476
rect -2309 14462 -2301 14474
rect -2070 14467 -2062 14472
rect -2000 14462 -1992 14509
rect -1942 14508 -1937 14510
rect -1932 14500 -1927 14508
rect -1912 14505 -1896 14511
rect -1842 14503 -1802 14514
rect -1671 14510 -1663 14518
rect -1663 14502 -1655 14510
rect -1850 14498 -1680 14502
rect -1924 14484 -1921 14486
rect -1806 14476 -1680 14482
rect -1671 14476 -1663 14490
rect -1663 14474 -1655 14476
rect -1854 14467 -1806 14472
rect -1974 14462 -1964 14463
rect -1960 14462 -1944 14464
rect -1842 14462 -1806 14465
rect -1655 14462 -1647 14474
rect -1642 14462 -1637 14556
rect -1619 14462 -1614 14556
rect -1530 14462 -1526 14556
rect -1506 14462 -1502 14556
rect -1482 14462 -1478 14556
rect -1458 14462 -1454 14556
rect -1434 14462 -1430 14556
rect -1410 14462 -1406 14556
rect -1386 14462 -1382 14556
rect -1362 14462 -1358 14556
rect -1338 14462 -1334 14556
rect -1314 14462 -1310 14556
rect -1290 14462 -1286 14556
rect -1266 14462 -1262 14556
rect -1242 14462 -1238 14556
rect -1218 14462 -1214 14556
rect -1194 14462 -1190 14556
rect -1170 14462 -1166 14556
rect -1146 14462 -1142 14556
rect -1122 14462 -1118 14556
rect -1098 14462 -1094 14556
rect -1074 14462 -1070 14556
rect -1050 14462 -1046 14556
rect -1026 14462 -1022 14556
rect -1002 14462 -998 14556
rect -978 14462 -974 14556
rect -954 14462 -950 14556
rect -930 14462 -926 14556
rect -906 14462 -902 14556
rect -882 14462 -878 14556
rect -858 14462 -854 14556
rect -834 14462 -830 14556
rect -810 14462 -806 14556
rect -786 14462 -782 14556
rect -762 14462 -758 14556
rect -738 14462 -734 14556
rect -725 14525 -720 14535
rect -714 14525 -710 14556
rect -715 14511 -710 14525
rect -725 14510 -691 14511
rect -690 14510 -686 14556
rect -666 14510 -662 14556
rect -642 14510 -638 14556
rect -618 14510 -614 14556
rect -594 14510 -590 14556
rect -570 14510 -566 14556
rect -546 14510 -542 14556
rect -522 14510 -518 14556
rect -498 14510 -494 14556
rect -474 14510 -470 14556
rect -450 14510 -446 14556
rect -426 14510 -422 14556
rect -402 14510 -398 14556
rect -378 14510 -374 14556
rect -354 14510 -350 14556
rect -330 14510 -326 14556
rect -306 14510 -302 14556
rect -282 14510 -278 14556
rect -258 14510 -254 14556
rect -234 14510 -230 14556
rect -210 14510 -206 14556
rect -186 14510 -182 14556
rect -162 14510 -158 14556
rect -138 14510 -134 14556
rect -114 14510 -110 14556
rect -90 14510 -86 14556
rect -66 14510 -62 14556
rect -42 14510 -38 14556
rect -18 14510 -14 14556
rect 6 14510 10 14556
rect 30 14510 34 14556
rect 54 14510 58 14556
rect 78 14510 82 14556
rect 102 14510 106 14556
rect 126 14510 130 14556
rect 150 14510 154 14556
rect 174 14510 178 14556
rect 198 14510 202 14556
rect 222 14510 226 14556
rect 246 14510 250 14556
rect 270 14510 274 14556
rect 294 14510 298 14556
rect 318 14510 322 14556
rect 342 14510 346 14556
rect 366 14510 370 14556
rect 390 14510 394 14556
rect 414 14510 418 14556
rect 438 14510 442 14556
rect 462 14510 466 14556
rect 486 14510 490 14556
rect 510 14510 514 14556
rect 534 14510 538 14556
rect 558 14510 562 14556
rect 582 14510 586 14556
rect 606 14510 610 14556
rect 630 14510 634 14556
rect 654 14510 658 14556
rect 678 14510 682 14556
rect 702 14510 706 14556
rect 726 14510 730 14556
rect 750 14510 754 14556
rect 774 14510 778 14556
rect 798 14510 802 14556
rect 822 14510 826 14556
rect 846 14510 850 14556
rect 870 14510 874 14556
rect 894 14510 898 14556
rect 918 14510 922 14556
rect 942 14510 946 14556
rect 966 14510 970 14556
rect 990 14510 994 14556
rect 1014 14510 1018 14556
rect 1038 14510 1042 14556
rect 1062 14510 1066 14556
rect 1086 14510 1090 14556
rect 1110 14510 1114 14556
rect 1134 14510 1138 14556
rect 1141 14555 1155 14556
rect 1158 14531 1165 14579
rect 1158 14510 1162 14531
rect 1182 14510 1186 14604
rect 1206 14510 1210 14604
rect 1230 14510 1234 14604
rect 1254 14510 1258 14604
rect 1278 14510 1282 14604
rect 1302 14510 1306 14604
rect 1326 14510 1330 14604
rect 1350 14510 1354 14604
rect 1374 14510 1378 14604
rect 1398 14510 1402 14604
rect 1422 14510 1426 14604
rect 1446 14510 1450 14604
rect 1470 14510 1474 14604
rect 1494 14510 1498 14604
rect 1518 14510 1522 14604
rect 1542 14510 1546 14604
rect 1566 14510 1570 14604
rect 1590 14510 1594 14604
rect 1614 14510 1618 14604
rect 1638 14510 1642 14604
rect 1662 14510 1666 14604
rect 1686 14510 1690 14604
rect 1710 14510 1714 14604
rect 1734 14510 1738 14604
rect 1758 14510 1762 14604
rect 1782 14510 1786 14604
rect 1806 14510 1810 14604
rect 1830 14510 1834 14604
rect 1854 14510 1858 14604
rect 1878 14510 1882 14604
rect 1902 14603 1906 14604
rect 1902 14579 1909 14603
rect 1902 14510 1906 14579
rect 1926 14510 1930 14604
rect 1950 14510 1954 14604
rect 1974 14510 1978 14604
rect 1998 14510 2002 14604
rect 2022 14510 2026 14604
rect 2046 14510 2050 14604
rect 2070 14510 2074 14604
rect 2094 14510 2098 14604
rect 2118 14510 2122 14604
rect 2142 14510 2146 14604
rect 2166 14510 2170 14604
rect 2190 14510 2194 14604
rect 2214 14510 2218 14604
rect 2238 14510 2242 14604
rect 2262 14510 2266 14604
rect 2286 14510 2290 14604
rect 2310 14510 2314 14604
rect 2334 14510 2338 14604
rect 2358 14510 2362 14604
rect 2382 14510 2386 14604
rect 2406 14510 2410 14604
rect 2430 14510 2434 14604
rect 2454 14510 2458 14604
rect 2478 14510 2482 14604
rect 2502 14510 2506 14604
rect 2526 14510 2530 14604
rect 2550 14510 2554 14604
rect 2574 14510 2578 14604
rect 2598 14510 2602 14604
rect 2622 14510 2626 14604
rect 2646 14510 2650 14604
rect 2670 14510 2674 14604
rect 2694 14510 2698 14604
rect 2718 14510 2722 14604
rect 2742 14510 2746 14604
rect 2766 14510 2770 14604
rect 2790 14510 2794 14604
rect 2814 14510 2818 14604
rect 2838 14510 2842 14604
rect 2862 14510 2866 14604
rect 2886 14510 2890 14604
rect 2910 14510 2914 14604
rect 2934 14510 2938 14604
rect 2958 14510 2962 14604
rect 2982 14510 2986 14604
rect 3006 14510 3010 14604
rect 3030 14510 3034 14604
rect 3054 14510 3058 14604
rect 3078 14510 3082 14604
rect 3102 14510 3106 14604
rect 3126 14510 3130 14604
rect 3150 14510 3154 14604
rect 3174 14510 3178 14604
rect 3198 14510 3202 14604
rect 3222 14510 3226 14604
rect 3246 14510 3250 14604
rect 3259 14549 3264 14559
rect 3270 14549 3274 14604
rect 3269 14535 3274 14549
rect 3270 14510 3274 14535
rect 3294 14510 3298 14604
rect 3318 14510 3322 14604
rect 3342 14510 3346 14604
rect 3366 14510 3370 14604
rect 3390 14510 3394 14604
rect 3414 14510 3418 14604
rect 3438 14510 3442 14604
rect 3462 14510 3466 14604
rect 3486 14510 3490 14604
rect 3510 14510 3514 14604
rect 3534 14510 3538 14604
rect 3558 14510 3562 14604
rect 3582 14510 3586 14604
rect 3606 14510 3610 14604
rect 3619 14597 3624 14604
rect 3637 14603 3651 14604
rect 3629 14583 3634 14597
rect 3630 14511 3634 14583
rect 3619 14510 3651 14511
rect -725 14508 3651 14510
rect -725 14501 -720 14508
rect -715 14487 -710 14501
rect -714 14462 -710 14487
rect -690 14462 -686 14508
rect -666 14462 -662 14508
rect -642 14462 -638 14508
rect -618 14462 -614 14508
rect -594 14462 -590 14508
rect -570 14462 -566 14508
rect -546 14462 -542 14508
rect -522 14462 -518 14508
rect -498 14462 -494 14508
rect -474 14462 -470 14508
rect -450 14462 -446 14508
rect -426 14462 -422 14508
rect -402 14462 -398 14508
rect -378 14462 -374 14508
rect -354 14462 -350 14508
rect -330 14462 -326 14508
rect -306 14462 -302 14508
rect -282 14462 -278 14508
rect -258 14462 -254 14508
rect -234 14462 -230 14508
rect -210 14462 -206 14508
rect -186 14462 -182 14508
rect -162 14462 -158 14508
rect -138 14462 -134 14508
rect -114 14462 -110 14508
rect -90 14462 -86 14508
rect -66 14462 -62 14508
rect -42 14462 -38 14508
rect -18 14462 -14 14508
rect 6 14462 10 14508
rect 30 14462 34 14508
rect 54 14462 58 14508
rect 78 14462 82 14508
rect 102 14462 106 14508
rect 126 14462 130 14508
rect 150 14462 154 14508
rect 174 14462 178 14508
rect 198 14462 202 14508
rect 222 14462 226 14508
rect 246 14462 250 14508
rect 270 14462 274 14508
rect 294 14462 298 14508
rect 318 14462 322 14508
rect 342 14462 346 14508
rect 366 14462 370 14508
rect 390 14462 394 14508
rect 414 14462 418 14508
rect 438 14462 442 14508
rect 462 14462 466 14508
rect 486 14462 490 14508
rect 510 14462 514 14508
rect 534 14462 538 14508
rect 558 14462 562 14508
rect 582 14462 586 14508
rect 606 14462 610 14508
rect 630 14462 634 14508
rect 654 14462 658 14508
rect 678 14462 682 14508
rect 702 14462 706 14508
rect 726 14462 730 14508
rect 750 14462 754 14508
rect 774 14462 778 14508
rect 798 14462 802 14508
rect 822 14462 826 14508
rect 846 14462 850 14508
rect 870 14462 874 14508
rect 894 14462 898 14508
rect 918 14462 922 14508
rect 942 14462 946 14508
rect 966 14462 970 14508
rect 990 14462 994 14508
rect 1014 14462 1018 14508
rect 1038 14462 1042 14508
rect 1062 14462 1066 14508
rect 1086 14462 1090 14508
rect 1110 14462 1114 14508
rect 1134 14462 1138 14508
rect 1158 14462 1162 14508
rect 1182 14462 1186 14508
rect 1206 14462 1210 14508
rect 1230 14462 1234 14508
rect 1254 14462 1258 14508
rect 1278 14462 1282 14508
rect 1302 14462 1306 14508
rect 1326 14462 1330 14508
rect 1350 14462 1354 14508
rect 1374 14462 1378 14508
rect 1398 14462 1402 14508
rect 1422 14462 1426 14508
rect 1446 14462 1450 14508
rect 1470 14462 1474 14508
rect 1494 14462 1498 14508
rect 1518 14462 1522 14508
rect 1542 14462 1546 14508
rect 1566 14462 1570 14508
rect 1590 14462 1594 14508
rect 1614 14462 1618 14508
rect 1638 14462 1642 14508
rect 1662 14462 1666 14508
rect 1686 14462 1690 14508
rect 1710 14462 1714 14508
rect 1734 14462 1738 14508
rect 1758 14462 1762 14508
rect 1782 14462 1786 14508
rect 1806 14462 1810 14508
rect 1830 14462 1834 14508
rect 1854 14462 1858 14508
rect 1878 14462 1882 14508
rect 1902 14462 1906 14508
rect 1926 14462 1930 14508
rect 1950 14462 1954 14508
rect 1974 14462 1978 14508
rect 1998 14462 2002 14508
rect 2022 14462 2026 14508
rect 2046 14463 2050 14508
rect 2035 14462 2069 14463
rect -2393 14460 2069 14462
rect -2371 14438 -2366 14460
rect -2348 14438 -2343 14460
rect -2325 14448 -2317 14460
rect -2325 14438 -2320 14448
rect -2317 14446 -2309 14448
rect -2062 14447 -2032 14454
rect -2309 14438 -2301 14446
rect -2070 14440 -2062 14447
rect -2000 14442 -1992 14460
rect -1974 14458 -1944 14460
rect -1960 14457 -1944 14458
rect -1842 14456 -1806 14460
rect -1842 14449 -1798 14454
rect -1806 14447 -1798 14449
rect -1671 14448 -1663 14460
rect -1854 14445 -1842 14447
rect -1663 14446 -1655 14448
rect -2062 14438 -2036 14440
rect -2393 14436 -2036 14438
rect -2032 14438 -2012 14440
rect -2004 14438 -1974 14442
rect -1854 14440 -1806 14445
rect -1864 14438 -1796 14439
rect -1655 14438 -1647 14446
rect -1642 14438 -1637 14460
rect -1619 14438 -1614 14460
rect -1530 14438 -1526 14460
rect -1506 14439 -1502 14460
rect -1517 14438 -1483 14439
rect -2032 14436 -1483 14438
rect -2371 14390 -2366 14436
rect -2348 14390 -2343 14436
rect -2325 14432 -2320 14436
rect -2309 14434 -2301 14436
rect -2317 14432 -2309 14434
rect -2325 14420 -2317 14432
rect -2052 14430 -2036 14432
rect -2052 14428 -2032 14430
rect -2062 14422 -2032 14428
rect -2325 14390 -2320 14420
rect -2317 14418 -2309 14420
rect -2092 14406 -2062 14408
rect -2094 14402 -2062 14406
rect -2000 14390 -1992 14436
rect -1904 14429 -1874 14436
rect -1842 14429 -1806 14436
rect -1655 14434 -1647 14436
rect -1663 14432 -1655 14434
rect -1842 14422 -1680 14428
rect -1671 14420 -1663 14432
rect -1663 14418 -1655 14420
rect -1854 14406 -1806 14408
rect -1854 14402 -1680 14406
rect -1642 14390 -1637 14436
rect -1619 14390 -1614 14436
rect -1530 14390 -1526 14436
rect -1517 14429 -1512 14436
rect -1506 14429 -1502 14436
rect -1507 14415 -1502 14429
rect -1506 14390 -1502 14415
rect -1482 14390 -1478 14460
rect -1458 14390 -1454 14460
rect -1434 14390 -1430 14460
rect -1410 14390 -1406 14460
rect -1386 14390 -1382 14460
rect -1362 14390 -1358 14460
rect -1338 14390 -1334 14460
rect -1314 14390 -1310 14460
rect -1290 14390 -1286 14460
rect -1266 14390 -1262 14460
rect -1242 14390 -1238 14460
rect -1218 14390 -1214 14460
rect -1194 14390 -1190 14460
rect -1170 14390 -1166 14460
rect -1146 14390 -1142 14460
rect -1122 14390 -1118 14460
rect -1098 14390 -1094 14460
rect -1074 14390 -1070 14460
rect -1050 14390 -1046 14460
rect -1026 14390 -1022 14460
rect -1002 14390 -998 14460
rect -978 14390 -974 14460
rect -954 14390 -950 14460
rect -930 14390 -926 14460
rect -906 14390 -902 14460
rect -882 14390 -878 14460
rect -858 14390 -854 14460
rect -834 14390 -830 14460
rect -810 14390 -806 14460
rect -786 14390 -782 14460
rect -762 14390 -758 14460
rect -738 14390 -734 14460
rect -714 14390 -710 14460
rect -690 14459 -686 14460
rect -690 14411 -683 14459
rect -690 14390 -686 14411
rect -666 14390 -662 14460
rect -642 14390 -638 14460
rect -618 14390 -614 14460
rect -594 14390 -590 14460
rect -570 14390 -566 14460
rect -546 14390 -542 14460
rect -522 14390 -518 14460
rect -498 14390 -494 14460
rect -474 14390 -470 14460
rect -450 14390 -446 14460
rect -426 14390 -422 14460
rect -402 14390 -398 14460
rect -378 14390 -374 14460
rect -354 14390 -350 14460
rect -330 14390 -326 14460
rect -306 14390 -302 14460
rect -282 14390 -278 14460
rect -258 14390 -254 14460
rect -234 14390 -230 14460
rect -210 14390 -206 14460
rect -186 14390 -182 14460
rect -162 14390 -158 14460
rect -138 14390 -134 14460
rect -114 14390 -110 14460
rect -90 14390 -86 14460
rect -66 14390 -62 14460
rect -42 14390 -38 14460
rect -18 14390 -14 14460
rect 6 14390 10 14460
rect 30 14390 34 14460
rect 54 14390 58 14460
rect 78 14390 82 14460
rect 102 14390 106 14460
rect 126 14390 130 14460
rect 150 14390 154 14460
rect 174 14390 178 14460
rect 198 14390 202 14460
rect 222 14390 226 14460
rect 246 14390 250 14460
rect 270 14390 274 14460
rect 294 14390 298 14460
rect 318 14390 322 14460
rect 342 14390 346 14460
rect 366 14390 370 14460
rect 390 14390 394 14460
rect 414 14390 418 14460
rect 438 14390 442 14460
rect 462 14390 466 14460
rect 486 14390 490 14460
rect 510 14390 514 14460
rect 534 14390 538 14460
rect 558 14390 562 14460
rect 582 14390 586 14460
rect 606 14390 610 14460
rect 630 14390 634 14460
rect 654 14390 658 14460
rect 678 14390 682 14460
rect 702 14390 706 14460
rect 726 14390 730 14460
rect 750 14390 754 14460
rect 774 14390 778 14460
rect 798 14390 802 14460
rect 822 14390 826 14460
rect 846 14390 850 14460
rect 870 14390 874 14460
rect 894 14390 898 14460
rect 918 14390 922 14460
rect 942 14390 946 14460
rect 966 14390 970 14460
rect 990 14390 994 14460
rect 1014 14390 1018 14460
rect 1038 14390 1042 14460
rect 1062 14390 1066 14460
rect 1086 14390 1090 14460
rect 1110 14390 1114 14460
rect 1134 14390 1138 14460
rect 1158 14390 1162 14460
rect 1182 14390 1186 14460
rect 1206 14390 1210 14460
rect 1230 14390 1234 14460
rect 1254 14390 1258 14460
rect 1278 14390 1282 14460
rect 1302 14390 1306 14460
rect 1326 14390 1330 14460
rect 1350 14390 1354 14460
rect 1374 14390 1378 14460
rect 1398 14390 1402 14460
rect 1422 14390 1426 14460
rect 1446 14390 1450 14460
rect 1470 14390 1474 14460
rect 1494 14390 1498 14460
rect 1518 14390 1522 14460
rect 1542 14390 1546 14460
rect 1566 14390 1570 14460
rect 1590 14390 1594 14460
rect 1614 14390 1618 14460
rect 1638 14390 1642 14460
rect 1662 14390 1666 14460
rect 1686 14390 1690 14460
rect 1710 14390 1714 14460
rect 1734 14390 1738 14460
rect 1758 14390 1762 14460
rect 1782 14390 1786 14460
rect 1806 14390 1810 14460
rect 1830 14390 1834 14460
rect 1854 14390 1858 14460
rect 1878 14390 1882 14460
rect 1902 14390 1906 14460
rect 1926 14390 1930 14460
rect 1950 14390 1954 14460
rect 1974 14390 1978 14460
rect 1998 14390 2002 14460
rect 2022 14390 2026 14460
rect 2035 14453 2040 14460
rect 2046 14453 2050 14460
rect 2045 14439 2050 14453
rect 2035 14429 2040 14439
rect 2045 14415 2050 14429
rect 2046 14390 2050 14415
rect 2070 14390 2074 14508
rect 2094 14390 2098 14508
rect 2118 14390 2122 14508
rect 2142 14390 2146 14508
rect 2166 14390 2170 14508
rect 2190 14390 2194 14508
rect 2214 14390 2218 14508
rect 2238 14390 2242 14508
rect 2262 14390 2266 14508
rect 2286 14390 2290 14508
rect 2310 14390 2314 14508
rect 2334 14390 2338 14508
rect 2358 14390 2362 14508
rect 2382 14390 2386 14508
rect 2406 14390 2410 14508
rect 2430 14390 2434 14508
rect 2454 14390 2458 14508
rect 2478 14390 2482 14508
rect 2502 14390 2506 14508
rect 2526 14390 2530 14508
rect 2550 14390 2554 14508
rect 2574 14390 2578 14508
rect 2598 14390 2602 14508
rect 2622 14390 2626 14508
rect 2646 14390 2650 14508
rect 2670 14390 2674 14508
rect 2694 14390 2698 14508
rect 2718 14390 2722 14508
rect 2742 14390 2746 14508
rect 2766 14390 2770 14508
rect 2790 14390 2794 14508
rect 2814 14390 2818 14508
rect 2838 14390 2842 14508
rect 2862 14390 2866 14508
rect 2886 14390 2890 14508
rect 2910 14390 2914 14508
rect 2934 14390 2938 14508
rect 2958 14390 2962 14508
rect 2982 14390 2986 14508
rect 3006 14390 3010 14508
rect 3030 14390 3034 14508
rect 3054 14390 3058 14508
rect 3078 14390 3082 14508
rect 3102 14390 3106 14508
rect 3126 14390 3130 14508
rect 3150 14390 3154 14508
rect 3174 14390 3178 14508
rect 3198 14390 3202 14508
rect 3222 14390 3226 14508
rect 3246 14390 3250 14508
rect 3270 14390 3274 14508
rect 3294 14483 3298 14508
rect 3294 14459 3301 14483
rect 3294 14390 3298 14459
rect 3318 14390 3322 14508
rect 3342 14390 3346 14508
rect 3366 14390 3370 14508
rect 3390 14390 3394 14508
rect 3414 14390 3418 14508
rect 3438 14390 3442 14508
rect 3462 14390 3466 14508
rect 3486 14390 3490 14508
rect 3510 14390 3514 14508
rect 3534 14390 3538 14508
rect 3558 14390 3562 14508
rect 3582 14390 3586 14508
rect 3606 14390 3610 14508
rect 3619 14501 3624 14508
rect 3630 14501 3634 14508
rect 3637 14507 3651 14508
rect 3629 14487 3634 14501
rect 3619 14477 3624 14487
rect 3629 14463 3634 14477
rect 3619 14429 3624 14439
rect 3630 14429 3634 14463
rect 3629 14415 3634 14429
rect 3643 14425 3651 14429
rect 3637 14415 3643 14425
rect 3619 14390 3651 14391
rect -2393 14388 3651 14390
rect -2371 14366 -2366 14388
rect -2348 14366 -2343 14388
rect -2325 14366 -2320 14388
rect -2072 14386 -2036 14387
rect -2072 14380 -2054 14386
rect -2309 14372 -2301 14380
rect -2317 14366 -2309 14372
rect -2092 14371 -2062 14376
rect -2000 14367 -1992 14388
rect -1938 14387 -1906 14388
rect -1920 14386 -1906 14387
rect -1806 14380 -1680 14386
rect -1854 14371 -1806 14376
rect -1655 14372 -1647 14380
rect -1982 14367 -1966 14368
rect -2000 14366 -1966 14367
rect -1846 14366 -1806 14369
rect -1663 14366 -1655 14372
rect -1642 14366 -1637 14388
rect -1619 14366 -1614 14388
rect -1530 14366 -1526 14388
rect -1506 14366 -1502 14388
rect -1482 14366 -1478 14388
rect -1458 14366 -1454 14388
rect -1434 14366 -1430 14388
rect -1410 14366 -1406 14388
rect -1386 14366 -1382 14388
rect -1362 14366 -1358 14388
rect -1338 14366 -1334 14388
rect -1314 14366 -1310 14388
rect -1290 14366 -1286 14388
rect -1266 14366 -1262 14388
rect -1242 14366 -1238 14388
rect -1218 14366 -1214 14388
rect -1194 14366 -1190 14388
rect -1170 14366 -1166 14388
rect -1146 14366 -1142 14388
rect -1122 14366 -1118 14388
rect -1098 14366 -1094 14388
rect -1074 14366 -1070 14388
rect -1050 14366 -1046 14388
rect -1026 14366 -1022 14388
rect -1002 14366 -998 14388
rect -978 14366 -974 14388
rect -954 14367 -950 14388
rect -965 14366 -931 14367
rect -2393 14364 -931 14366
rect -2371 14342 -2366 14364
rect -2348 14342 -2343 14364
rect -2325 14342 -2320 14364
rect -2000 14362 -1966 14364
rect -2309 14344 -2301 14352
rect -2062 14351 -2054 14358
rect -2092 14344 -2084 14351
rect -2062 14344 -2026 14346
rect -2317 14342 -2309 14344
rect -2062 14342 -2012 14344
rect -2000 14342 -1992 14362
rect -1982 14361 -1966 14362
rect -1846 14360 -1806 14364
rect -1846 14353 -1798 14358
rect -1806 14351 -1798 14353
rect -1854 14349 -1846 14351
rect -1854 14344 -1806 14349
rect -1655 14344 -1647 14352
rect -1864 14342 -1796 14343
rect -1663 14342 -1655 14344
rect -1642 14342 -1637 14364
rect -1619 14342 -1614 14364
rect -1530 14342 -1526 14364
rect -1506 14342 -1502 14364
rect -1482 14363 -1478 14364
rect -2393 14340 -1485 14342
rect -2371 14294 -2366 14340
rect -2348 14294 -2343 14340
rect -2325 14294 -2320 14340
rect -2317 14336 -2309 14340
rect -2062 14336 -2054 14340
rect -2154 14332 -2138 14334
rect -2057 14332 -2054 14336
rect -2292 14326 -2054 14332
rect -2052 14326 -2044 14336
rect -2092 14310 -2062 14312
rect -2094 14306 -2062 14310
rect -2000 14294 -1992 14340
rect -1846 14333 -1806 14340
rect -1663 14336 -1655 14340
rect -1846 14326 -1680 14332
rect -1854 14310 -1806 14312
rect -1854 14306 -1680 14310
rect -1642 14294 -1637 14340
rect -1619 14294 -1614 14340
rect -1530 14294 -1526 14340
rect -1506 14294 -1502 14340
rect -1499 14339 -1485 14340
rect -1482 14339 -1475 14363
rect -1482 14294 -1478 14339
rect -1458 14294 -1454 14364
rect -1434 14294 -1430 14364
rect -1410 14294 -1406 14364
rect -1386 14294 -1382 14364
rect -1362 14294 -1358 14364
rect -1338 14294 -1334 14364
rect -1314 14294 -1310 14364
rect -1290 14294 -1286 14364
rect -1266 14294 -1262 14364
rect -1242 14294 -1238 14364
rect -1218 14294 -1214 14364
rect -1194 14294 -1190 14364
rect -1170 14294 -1166 14364
rect -1146 14294 -1142 14364
rect -1122 14294 -1118 14364
rect -1098 14294 -1094 14364
rect -1074 14294 -1070 14364
rect -1050 14294 -1046 14364
rect -1026 14294 -1022 14364
rect -1002 14294 -998 14364
rect -978 14294 -974 14364
rect -965 14357 -960 14364
rect -954 14357 -950 14364
rect -955 14343 -950 14357
rect -954 14294 -950 14343
rect -930 14294 -926 14388
rect -906 14294 -902 14388
rect -882 14294 -878 14388
rect -858 14294 -854 14388
rect -834 14294 -830 14388
rect -810 14294 -806 14388
rect -786 14294 -782 14388
rect -762 14294 -758 14388
rect -738 14294 -734 14388
rect -714 14294 -710 14388
rect -690 14294 -686 14388
rect -666 14294 -662 14388
rect -642 14294 -638 14388
rect -618 14294 -614 14388
rect -594 14294 -590 14388
rect -570 14294 -566 14388
rect -546 14294 -542 14388
rect -522 14294 -518 14388
rect -498 14294 -494 14388
rect -474 14294 -470 14388
rect -450 14294 -446 14388
rect -426 14294 -422 14388
rect -402 14294 -398 14388
rect -378 14294 -374 14388
rect -354 14294 -350 14388
rect -330 14294 -326 14388
rect -306 14294 -302 14388
rect -282 14294 -278 14388
rect -258 14294 -254 14388
rect -234 14294 -230 14388
rect -210 14294 -206 14388
rect -186 14294 -182 14388
rect -162 14294 -158 14388
rect -138 14294 -134 14388
rect -114 14294 -110 14388
rect -90 14294 -86 14388
rect -66 14294 -62 14388
rect -42 14294 -38 14388
rect -18 14294 -14 14388
rect 6 14294 10 14388
rect 30 14294 34 14388
rect 54 14294 58 14388
rect 78 14294 82 14388
rect 102 14294 106 14388
rect 126 14294 130 14388
rect 150 14294 154 14388
rect 174 14294 178 14388
rect 198 14294 202 14388
rect 222 14294 226 14388
rect 246 14294 250 14388
rect 270 14294 274 14388
rect 294 14294 298 14388
rect 318 14294 322 14388
rect 342 14294 346 14388
rect 366 14294 370 14388
rect 390 14294 394 14388
rect 414 14294 418 14388
rect 438 14294 442 14388
rect 462 14294 466 14388
rect 486 14294 490 14388
rect 510 14294 514 14388
rect 534 14294 538 14388
rect 558 14294 562 14388
rect 582 14294 586 14388
rect 606 14294 610 14388
rect 630 14294 634 14388
rect 654 14294 658 14388
rect 678 14294 682 14388
rect 702 14294 706 14388
rect 726 14294 730 14388
rect 750 14294 754 14388
rect 774 14294 778 14388
rect 798 14294 802 14388
rect 822 14294 826 14388
rect 846 14294 850 14388
rect 870 14294 874 14388
rect 894 14294 898 14388
rect 918 14294 922 14388
rect 942 14294 946 14388
rect 955 14333 960 14343
rect 966 14333 970 14388
rect 965 14319 970 14333
rect 966 14294 970 14319
rect 990 14294 994 14388
rect 1014 14294 1018 14388
rect 1038 14294 1042 14388
rect 1062 14294 1066 14388
rect 1086 14294 1090 14388
rect 1110 14294 1114 14388
rect 1134 14294 1138 14388
rect 1158 14294 1162 14388
rect 1182 14294 1186 14388
rect 1206 14294 1210 14388
rect 1230 14294 1234 14388
rect 1254 14294 1258 14388
rect 1278 14294 1282 14388
rect 1302 14294 1306 14388
rect 1326 14294 1330 14388
rect 1350 14294 1354 14388
rect 1374 14294 1378 14388
rect 1398 14294 1402 14388
rect 1422 14294 1426 14388
rect 1446 14294 1450 14388
rect 1470 14294 1474 14388
rect 1494 14294 1498 14388
rect 1518 14294 1522 14388
rect 1542 14294 1546 14388
rect 1566 14294 1570 14388
rect 1590 14294 1594 14388
rect 1614 14294 1618 14388
rect 1638 14294 1642 14388
rect 1662 14294 1666 14388
rect 1686 14294 1690 14388
rect 1710 14294 1714 14388
rect 1734 14294 1738 14388
rect 1758 14294 1762 14388
rect 1782 14294 1786 14388
rect 1806 14294 1810 14388
rect 1830 14294 1834 14388
rect 1854 14294 1858 14388
rect 1878 14294 1882 14388
rect 1902 14294 1906 14388
rect 1926 14294 1930 14388
rect 1950 14294 1954 14388
rect 1974 14294 1978 14388
rect 1998 14294 2002 14388
rect 2022 14294 2026 14388
rect 2046 14294 2050 14388
rect 2070 14387 2074 14388
rect 2070 14339 2077 14387
rect 2070 14294 2074 14339
rect 2094 14294 2098 14388
rect 2118 14294 2122 14388
rect 2142 14294 2146 14388
rect 2166 14294 2170 14388
rect 2190 14294 2194 14388
rect 2214 14294 2218 14388
rect 2238 14294 2242 14388
rect 2262 14294 2266 14388
rect 2286 14294 2290 14388
rect 2310 14294 2314 14388
rect 2334 14294 2338 14388
rect 2358 14294 2362 14388
rect 2382 14294 2386 14388
rect 2406 14294 2410 14388
rect 2430 14294 2434 14388
rect 2454 14294 2458 14388
rect 2478 14294 2482 14388
rect 2502 14294 2506 14388
rect 2526 14294 2530 14388
rect 2550 14294 2554 14388
rect 2574 14294 2578 14388
rect 2598 14294 2602 14388
rect 2622 14294 2626 14388
rect 2646 14294 2650 14388
rect 2670 14294 2674 14388
rect 2694 14294 2698 14388
rect 2718 14294 2722 14388
rect 2742 14294 2746 14388
rect 2766 14294 2770 14388
rect 2790 14294 2794 14388
rect 2814 14294 2818 14388
rect 2838 14294 2842 14388
rect 2862 14294 2866 14388
rect 2886 14294 2890 14388
rect 2910 14294 2914 14388
rect 2934 14294 2938 14388
rect 2958 14294 2962 14388
rect 2982 14294 2986 14388
rect 3006 14294 3010 14388
rect 3030 14294 3034 14388
rect 3054 14294 3058 14388
rect 3078 14294 3082 14388
rect 3102 14294 3106 14388
rect 3126 14294 3130 14388
rect 3150 14294 3154 14388
rect 3174 14294 3178 14388
rect 3198 14294 3202 14388
rect 3222 14294 3226 14388
rect 3246 14294 3250 14388
rect 3270 14294 3274 14388
rect 3294 14294 3298 14388
rect 3318 14294 3322 14388
rect 3342 14294 3346 14388
rect 3366 14294 3370 14388
rect 3390 14294 3394 14388
rect 3414 14294 3418 14388
rect 3438 14294 3442 14388
rect 3462 14294 3466 14388
rect 3486 14294 3490 14388
rect 3510 14294 3514 14388
rect 3534 14294 3538 14388
rect 3558 14294 3562 14388
rect 3582 14294 3586 14388
rect 3606 14294 3610 14388
rect 3619 14381 3624 14388
rect 3637 14387 3651 14388
rect 3629 14367 3634 14381
rect 3630 14294 3634 14367
rect 3643 14294 3651 14295
rect -2393 14292 3651 14294
rect -2371 14270 -2366 14292
rect -2348 14270 -2343 14292
rect -2325 14270 -2320 14292
rect -2072 14290 -2036 14291
rect -2072 14284 -2054 14290
rect -2309 14276 -2301 14284
rect -2317 14270 -2309 14276
rect -2092 14275 -2062 14280
rect -2000 14271 -1992 14292
rect -1938 14291 -1906 14292
rect -1920 14290 -1906 14291
rect -1806 14284 -1680 14290
rect -1854 14275 -1806 14280
rect -1655 14276 -1647 14284
rect -1982 14271 -1966 14272
rect -2000 14270 -1966 14271
rect -1846 14270 -1806 14273
rect -1663 14270 -1655 14276
rect -1642 14270 -1637 14292
rect -1619 14270 -1614 14292
rect -1530 14270 -1526 14292
rect -1506 14270 -1502 14292
rect -1482 14270 -1478 14292
rect -1458 14270 -1454 14292
rect -1434 14270 -1430 14292
rect -1410 14270 -1406 14292
rect -1386 14270 -1382 14292
rect -1362 14270 -1358 14292
rect -1338 14270 -1334 14292
rect -1314 14270 -1310 14292
rect -1290 14270 -1286 14292
rect -1266 14270 -1262 14292
rect -1242 14270 -1238 14292
rect -1218 14270 -1214 14292
rect -1194 14270 -1190 14292
rect -1170 14270 -1166 14292
rect -1146 14270 -1142 14292
rect -1122 14270 -1118 14292
rect -1098 14270 -1094 14292
rect -1074 14270 -1070 14292
rect -1050 14270 -1046 14292
rect -1026 14270 -1022 14292
rect -1002 14270 -998 14292
rect -978 14270 -974 14292
rect -954 14270 -950 14292
rect -930 14291 -926 14292
rect -2393 14268 -933 14270
rect -2371 14246 -2366 14268
rect -2348 14246 -2343 14268
rect -2325 14246 -2320 14268
rect -2000 14266 -1966 14268
rect -2309 14248 -2301 14256
rect -2062 14255 -2054 14262
rect -2092 14248 -2084 14255
rect -2062 14248 -2026 14250
rect -2317 14246 -2309 14248
rect -2062 14246 -2012 14248
rect -2000 14246 -1992 14266
rect -1982 14265 -1966 14266
rect -1846 14264 -1806 14268
rect -1846 14257 -1798 14262
rect -1806 14255 -1798 14257
rect -1854 14253 -1846 14255
rect -1854 14248 -1806 14253
rect -1655 14248 -1647 14256
rect -1864 14246 -1796 14247
rect -1663 14246 -1655 14248
rect -1642 14246 -1637 14268
rect -1619 14246 -1614 14268
rect -1530 14246 -1526 14268
rect -1506 14246 -1502 14268
rect -1482 14246 -1478 14268
rect -1458 14246 -1454 14268
rect -1434 14246 -1430 14268
rect -1410 14246 -1406 14268
rect -1386 14246 -1382 14268
rect -1362 14246 -1358 14268
rect -1338 14246 -1334 14268
rect -1314 14246 -1310 14268
rect -1290 14246 -1286 14268
rect -1266 14246 -1262 14268
rect -1242 14246 -1238 14268
rect -1218 14246 -1214 14268
rect -1194 14246 -1190 14268
rect -1170 14246 -1166 14268
rect -1146 14246 -1142 14268
rect -1122 14246 -1118 14268
rect -1098 14246 -1094 14268
rect -1074 14246 -1070 14268
rect -1050 14246 -1046 14268
rect -1026 14246 -1022 14268
rect -1002 14246 -998 14268
rect -978 14246 -974 14268
rect -954 14246 -950 14268
rect -947 14267 -933 14268
rect -930 14267 -923 14291
rect -930 14246 -926 14267
rect -906 14246 -902 14292
rect -882 14246 -878 14292
rect -858 14246 -854 14292
rect -834 14246 -830 14292
rect -810 14246 -806 14292
rect -786 14246 -782 14292
rect -762 14246 -758 14292
rect -738 14246 -734 14292
rect -714 14246 -710 14292
rect -690 14246 -686 14292
rect -666 14246 -662 14292
rect -642 14246 -638 14292
rect -618 14246 -614 14292
rect -594 14246 -590 14292
rect -570 14246 -566 14292
rect -546 14246 -542 14292
rect -522 14246 -518 14292
rect -498 14246 -494 14292
rect -474 14246 -470 14292
rect -450 14246 -446 14292
rect -426 14246 -422 14292
rect -402 14246 -398 14292
rect -378 14246 -374 14292
rect -354 14246 -350 14292
rect -330 14246 -326 14292
rect -306 14246 -302 14292
rect -282 14246 -278 14292
rect -258 14246 -254 14292
rect -234 14246 -230 14292
rect -210 14246 -206 14292
rect -186 14246 -182 14292
rect -162 14246 -158 14292
rect -138 14246 -134 14292
rect -114 14246 -110 14292
rect -90 14246 -86 14292
rect -66 14246 -62 14292
rect -42 14246 -38 14292
rect -18 14246 -14 14292
rect 6 14246 10 14292
rect 30 14246 34 14292
rect 54 14246 58 14292
rect 78 14246 82 14292
rect 102 14246 106 14292
rect 126 14246 130 14292
rect 150 14246 154 14292
rect 174 14246 178 14292
rect 198 14246 202 14292
rect 222 14246 226 14292
rect 246 14246 250 14292
rect 270 14246 274 14292
rect 294 14246 298 14292
rect 318 14246 322 14292
rect 342 14246 346 14292
rect 366 14246 370 14292
rect 390 14246 394 14292
rect 414 14246 418 14292
rect 438 14246 442 14292
rect 462 14246 466 14292
rect 475 14261 480 14271
rect 486 14261 490 14292
rect 485 14247 490 14261
rect 475 14246 509 14247
rect 510 14246 514 14292
rect 534 14246 538 14292
rect 558 14246 562 14292
rect 582 14246 586 14292
rect 606 14246 610 14292
rect 630 14246 634 14292
rect 654 14246 658 14292
rect 678 14246 682 14292
rect 702 14246 706 14292
rect 726 14246 730 14292
rect 750 14246 754 14292
rect 774 14246 778 14292
rect 798 14246 802 14292
rect 822 14246 826 14292
rect 846 14246 850 14292
rect 870 14246 874 14292
rect 894 14246 898 14292
rect 918 14246 922 14292
rect 942 14246 946 14292
rect 966 14246 970 14292
rect 990 14267 994 14292
rect -2393 14244 987 14246
rect -2371 14198 -2366 14244
rect -2348 14198 -2343 14244
rect -2325 14198 -2320 14244
rect -2317 14240 -2309 14244
rect -2062 14240 -2054 14244
rect -2154 14236 -2138 14238
rect -2057 14236 -2054 14240
rect -2292 14230 -2054 14236
rect -2052 14230 -2044 14240
rect -2092 14214 -2062 14216
rect -2094 14210 -2062 14214
rect -2000 14198 -1992 14244
rect -1846 14237 -1806 14244
rect -1663 14240 -1655 14244
rect -1846 14230 -1680 14236
rect -1854 14214 -1806 14216
rect -1854 14210 -1680 14214
rect -1979 14198 -1945 14200
rect -1642 14198 -1637 14244
rect -1619 14198 -1614 14244
rect -1530 14198 -1526 14244
rect -1506 14198 -1502 14244
rect -1482 14198 -1478 14244
rect -1458 14198 -1454 14244
rect -1434 14198 -1430 14244
rect -1410 14198 -1406 14244
rect -1386 14198 -1382 14244
rect -1362 14198 -1358 14244
rect -1338 14198 -1334 14244
rect -1314 14198 -1310 14244
rect -1290 14198 -1286 14244
rect -1266 14198 -1262 14244
rect -1242 14198 -1238 14244
rect -1218 14198 -1214 14244
rect -1194 14198 -1190 14244
rect -1170 14198 -1166 14244
rect -1146 14198 -1142 14244
rect -1122 14198 -1118 14244
rect -1098 14198 -1094 14244
rect -1074 14198 -1070 14244
rect -1050 14198 -1046 14244
rect -1026 14198 -1022 14244
rect -1002 14198 -998 14244
rect -978 14198 -974 14244
rect -954 14198 -950 14244
rect -930 14198 -926 14244
rect -906 14198 -902 14244
rect -882 14198 -878 14244
rect -858 14198 -854 14244
rect -834 14198 -830 14244
rect -810 14198 -806 14244
rect -786 14198 -782 14244
rect -762 14198 -758 14244
rect -738 14198 -734 14244
rect -714 14198 -710 14244
rect -690 14198 -686 14244
rect -666 14198 -662 14244
rect -642 14198 -638 14244
rect -618 14198 -614 14244
rect -594 14198 -590 14244
rect -570 14198 -566 14244
rect -546 14198 -542 14244
rect -522 14198 -518 14244
rect -498 14198 -494 14244
rect -474 14198 -470 14244
rect -450 14198 -446 14244
rect -426 14198 -422 14244
rect -402 14198 -398 14244
rect -378 14198 -374 14244
rect -354 14198 -350 14244
rect -330 14198 -326 14244
rect -306 14198 -302 14244
rect -282 14198 -278 14244
rect -258 14198 -254 14244
rect -234 14198 -230 14244
rect -210 14198 -206 14244
rect -186 14198 -182 14244
rect -162 14198 -158 14244
rect -138 14198 -134 14244
rect -114 14198 -110 14244
rect -90 14198 -86 14244
rect -66 14198 -62 14244
rect -42 14198 -38 14244
rect -18 14198 -14 14244
rect 6 14198 10 14244
rect 30 14198 34 14244
rect 54 14198 58 14244
rect 78 14198 82 14244
rect 102 14198 106 14244
rect 126 14198 130 14244
rect 150 14198 154 14244
rect 174 14198 178 14244
rect 198 14198 202 14244
rect 222 14198 226 14244
rect 246 14198 250 14244
rect 270 14198 274 14244
rect 294 14198 298 14244
rect 318 14198 322 14244
rect 342 14198 346 14244
rect 366 14198 370 14244
rect 390 14198 394 14244
rect 414 14198 418 14244
rect 438 14198 442 14244
rect 462 14198 466 14244
rect 475 14237 480 14244
rect 485 14223 490 14237
rect 486 14198 490 14223
rect 510 14198 514 14244
rect 534 14198 538 14244
rect 558 14198 562 14244
rect 582 14198 586 14244
rect 606 14198 610 14244
rect 630 14198 634 14244
rect 654 14198 658 14244
rect 678 14198 682 14244
rect 702 14198 706 14244
rect 726 14198 730 14244
rect 750 14198 754 14244
rect 774 14198 778 14244
rect 798 14198 802 14244
rect 822 14198 826 14244
rect 846 14198 850 14244
rect 870 14198 874 14244
rect 894 14198 898 14244
rect 918 14198 922 14244
rect 942 14198 946 14244
rect 966 14198 970 14244
rect 973 14243 987 14244
rect 990 14243 997 14267
rect 990 14198 994 14243
rect 1014 14198 1018 14292
rect 1038 14198 1042 14292
rect 1062 14198 1066 14292
rect 1086 14198 1090 14292
rect 1110 14198 1114 14292
rect 1134 14198 1138 14292
rect 1158 14198 1162 14292
rect 1182 14198 1186 14292
rect 1206 14198 1210 14292
rect 1230 14198 1234 14292
rect 1254 14198 1258 14292
rect 1278 14198 1282 14292
rect 1302 14198 1306 14292
rect 1326 14198 1330 14292
rect 1350 14198 1354 14292
rect 1374 14198 1378 14292
rect 1398 14198 1402 14292
rect 1422 14198 1426 14292
rect 1446 14198 1450 14292
rect 1470 14198 1474 14292
rect 1494 14198 1498 14292
rect 1518 14198 1522 14292
rect 1542 14198 1546 14292
rect 1566 14198 1570 14292
rect 1590 14198 1594 14292
rect 1614 14198 1618 14292
rect 1638 14198 1642 14292
rect 1662 14198 1666 14292
rect 1686 14198 1690 14292
rect 1710 14198 1714 14292
rect 1734 14198 1738 14292
rect 1758 14198 1762 14292
rect 1782 14198 1786 14292
rect 1806 14198 1810 14292
rect 1830 14198 1834 14292
rect 1854 14198 1858 14292
rect 1878 14198 1882 14292
rect 1902 14198 1906 14292
rect 1926 14198 1930 14292
rect 1950 14198 1954 14292
rect 1974 14198 1978 14292
rect 1998 14198 2002 14292
rect 2022 14198 2026 14292
rect 2046 14198 2050 14292
rect 2070 14198 2074 14292
rect 2094 14198 2098 14292
rect 2118 14198 2122 14292
rect 2142 14198 2146 14292
rect 2166 14198 2170 14292
rect 2190 14198 2194 14292
rect 2214 14198 2218 14292
rect 2238 14198 2242 14292
rect 2262 14198 2266 14292
rect 2286 14198 2290 14292
rect 2310 14198 2314 14292
rect 2334 14198 2338 14292
rect 2358 14198 2362 14292
rect 2382 14198 2386 14292
rect 2406 14198 2410 14292
rect 2430 14198 2434 14292
rect 2454 14198 2458 14292
rect 2478 14198 2482 14292
rect 2502 14198 2506 14292
rect 2526 14198 2530 14292
rect 2550 14198 2554 14292
rect 2574 14198 2578 14292
rect 2598 14198 2602 14292
rect 2622 14198 2626 14292
rect 2646 14198 2650 14292
rect 2670 14198 2674 14292
rect 2694 14198 2698 14292
rect 2718 14198 2722 14292
rect 2742 14198 2746 14292
rect 2766 14198 2770 14292
rect 2790 14198 2794 14292
rect 2814 14198 2818 14292
rect 2838 14198 2842 14292
rect 2862 14198 2866 14292
rect 2886 14198 2890 14292
rect 2910 14198 2914 14292
rect 2934 14198 2938 14292
rect 2958 14198 2962 14292
rect 2982 14198 2986 14292
rect 3006 14198 3010 14292
rect 3030 14198 3034 14292
rect 3054 14198 3058 14292
rect 3078 14198 3082 14292
rect 3102 14198 3106 14292
rect 3126 14198 3130 14292
rect 3150 14198 3154 14292
rect 3174 14198 3178 14292
rect 3198 14198 3202 14292
rect 3222 14198 3226 14292
rect 3246 14198 3250 14292
rect 3259 14237 3264 14247
rect 3270 14237 3274 14292
rect 3269 14223 3274 14237
rect 3259 14213 3264 14223
rect 3269 14199 3274 14213
rect 3270 14198 3274 14199
rect 3294 14198 3298 14292
rect 3318 14198 3322 14292
rect 3342 14198 3346 14292
rect 3366 14198 3370 14292
rect 3390 14198 3394 14292
rect 3414 14198 3418 14292
rect 3438 14198 3442 14292
rect 3462 14198 3466 14292
rect 3486 14198 3490 14292
rect 3510 14198 3514 14292
rect 3534 14198 3538 14292
rect 3558 14198 3562 14292
rect 3582 14198 3586 14292
rect 3606 14198 3610 14292
rect 3630 14198 3634 14292
rect 3637 14291 3651 14292
rect 3643 14285 3648 14291
rect 3653 14271 3658 14285
rect 3643 14213 3648 14223
rect 3654 14213 3658 14271
rect 3653 14199 3658 14213
rect 3667 14209 3675 14213
rect 3661 14199 3667 14209
rect 3643 14198 3675 14199
rect -2393 14196 3675 14198
rect -2371 14150 -2366 14196
rect -2348 14150 -2343 14196
rect -2325 14150 -2320 14196
rect -2080 14195 -1906 14196
rect -2080 14194 -2036 14195
rect -2080 14188 -2054 14194
rect -2309 14180 -2301 14186
rect -2317 14170 -2309 14180
rect -2070 14179 -2040 14186
rect -2054 14171 -2040 14174
rect -2000 14169 -1992 14195
rect -1920 14194 -1906 14195
rect -1850 14188 -1846 14196
rect -1840 14188 -1792 14196
rect -1969 14176 -1966 14185
rect -1850 14181 -1802 14186
rect -1906 14179 -1802 14181
rect -1655 14180 -1647 14186
rect -1906 14178 -1850 14179
rect -1846 14171 -1802 14177
rect -1663 14170 -1655 14180
rect -1860 14169 -1798 14170
rect -2078 14162 -2070 14169
rect -2309 14152 -2301 14158
rect -2317 14150 -2309 14152
rect -2154 14150 -2145 14160
rect -2044 14159 -2040 14164
rect -2028 14162 -1945 14169
rect -1929 14162 -1794 14169
rect -2070 14152 -2040 14159
rect -2044 14150 -2028 14152
rect -2000 14150 -1992 14162
rect -1860 14161 -1798 14162
rect -1850 14152 -1802 14159
rect -1655 14152 -1647 14158
rect -1978 14150 -1942 14151
rect -1663 14150 -1655 14152
rect -1642 14150 -1637 14196
rect -1619 14150 -1614 14196
rect -1530 14150 -1526 14196
rect -1506 14150 -1502 14196
rect -1482 14150 -1478 14196
rect -1458 14150 -1454 14196
rect -1434 14150 -1430 14196
rect -1410 14150 -1406 14196
rect -1386 14150 -1382 14196
rect -1362 14150 -1358 14196
rect -1338 14150 -1334 14196
rect -1314 14150 -1310 14196
rect -1290 14150 -1286 14196
rect -1266 14150 -1262 14196
rect -1242 14150 -1238 14196
rect -1218 14150 -1214 14196
rect -1194 14150 -1190 14196
rect -1170 14150 -1166 14196
rect -1146 14150 -1142 14196
rect -1122 14150 -1118 14196
rect -1098 14150 -1094 14196
rect -1074 14150 -1070 14196
rect -1050 14150 -1046 14196
rect -1026 14150 -1022 14196
rect -1002 14150 -998 14196
rect -978 14150 -974 14196
rect -954 14150 -950 14196
rect -930 14150 -926 14196
rect -906 14150 -902 14196
rect -882 14150 -878 14196
rect -858 14150 -854 14196
rect -834 14150 -830 14196
rect -810 14150 -806 14196
rect -786 14150 -782 14196
rect -762 14150 -758 14196
rect -738 14150 -734 14196
rect -714 14150 -710 14196
rect -690 14150 -686 14196
rect -666 14150 -662 14196
rect -642 14150 -638 14196
rect -618 14150 -614 14196
rect -594 14150 -590 14196
rect -570 14150 -566 14196
rect -546 14150 -542 14196
rect -522 14150 -518 14196
rect -498 14150 -494 14196
rect -474 14150 -470 14196
rect -450 14150 -446 14196
rect -426 14150 -422 14196
rect -402 14150 -398 14196
rect -378 14150 -374 14196
rect -354 14150 -350 14196
rect -330 14150 -326 14196
rect -306 14150 -302 14196
rect -282 14150 -278 14196
rect -258 14150 -254 14196
rect -234 14150 -230 14196
rect -210 14150 -206 14196
rect -186 14150 -182 14196
rect -162 14150 -158 14196
rect -138 14150 -134 14196
rect -114 14150 -110 14196
rect -90 14150 -86 14196
rect -66 14150 -62 14196
rect -42 14150 -38 14196
rect -18 14150 -14 14196
rect 6 14150 10 14196
rect 30 14150 34 14196
rect 54 14150 58 14196
rect 78 14150 82 14196
rect 102 14150 106 14196
rect 126 14150 130 14196
rect 150 14150 154 14196
rect 174 14150 178 14196
rect 198 14150 202 14196
rect 222 14150 226 14196
rect 246 14150 250 14196
rect 270 14150 274 14196
rect 294 14150 298 14196
rect 318 14150 322 14196
rect 342 14150 346 14196
rect 366 14150 370 14196
rect 390 14150 394 14196
rect 414 14150 418 14196
rect 438 14150 442 14196
rect 462 14150 466 14196
rect 486 14151 490 14196
rect 510 14195 514 14196
rect 475 14150 509 14151
rect -2393 14148 509 14150
rect -2371 14054 -2366 14148
rect -2348 14054 -2343 14148
rect -2325 14110 -2320 14148
rect -2317 14142 -2309 14148
rect -2145 14144 -2138 14148
rect -2070 14144 -2054 14148
rect -2078 14135 -2054 14142
rect -2062 14110 -2032 14111
rect -2000 14110 -1992 14148
rect -1846 14144 -1802 14148
rect -1846 14134 -1792 14143
rect -1663 14142 -1655 14148
rect -1942 14112 -1937 14124
rect -1850 14121 -1822 14122
rect -1850 14117 -1802 14121
rect -2325 14102 -2317 14110
rect -2062 14108 -1961 14110
rect -2325 14082 -2320 14102
rect -2317 14094 -2309 14102
rect -2062 14095 -2040 14106
rect -2032 14101 -1961 14108
rect -1947 14102 -1942 14110
rect -1842 14108 -1794 14111
rect -2070 14090 -2022 14094
rect -2325 14068 -2317 14082
rect -2072 14074 -2032 14075
rect -2102 14068 -2032 14074
rect -2325 14054 -2320 14068
rect -2317 14066 -2309 14068
rect -2309 14054 -2301 14066
rect -2070 14059 -2062 14064
rect -2000 14054 -1992 14101
rect -1942 14100 -1937 14102
rect -1932 14092 -1927 14100
rect -1912 14097 -1896 14103
rect -1842 14095 -1802 14106
rect -1671 14102 -1663 14110
rect -1663 14094 -1655 14102
rect -1850 14090 -1680 14094
rect -1924 14076 -1921 14078
rect -1806 14068 -1680 14074
rect -1671 14068 -1663 14082
rect -1663 14066 -1655 14068
rect -1854 14059 -1806 14064
rect -1974 14054 -1964 14055
rect -1960 14054 -1944 14056
rect -1842 14054 -1806 14057
rect -1655 14054 -1647 14066
rect -1642 14054 -1637 14148
rect -1619 14054 -1614 14148
rect -1530 14054 -1526 14148
rect -1506 14054 -1502 14148
rect -1482 14054 -1478 14148
rect -1458 14054 -1454 14148
rect -1434 14054 -1430 14148
rect -1410 14054 -1406 14148
rect -1386 14055 -1382 14148
rect -1397 14054 -1363 14055
rect -2393 14052 -1363 14054
rect -2371 14030 -2366 14052
rect -2348 14030 -2343 14052
rect -2325 14040 -2317 14052
rect -2325 14030 -2320 14040
rect -2317 14038 -2309 14040
rect -2062 14039 -2032 14046
rect -2309 14030 -2301 14038
rect -2070 14032 -2062 14039
rect -2000 14034 -1992 14052
rect -1974 14050 -1944 14052
rect -1960 14049 -1944 14050
rect -1842 14048 -1806 14052
rect -1842 14041 -1798 14046
rect -1806 14039 -1798 14041
rect -1671 14040 -1663 14052
rect -1854 14037 -1842 14039
rect -1663 14038 -1655 14040
rect -2062 14030 -2036 14032
rect -2393 14028 -2036 14030
rect -2032 14030 -2012 14032
rect -2004 14030 -1974 14034
rect -1854 14032 -1806 14037
rect -1864 14030 -1796 14031
rect -1655 14030 -1647 14038
rect -1642 14030 -1637 14052
rect -1619 14030 -1614 14052
rect -1530 14030 -1526 14052
rect -1506 14030 -1502 14052
rect -1482 14030 -1478 14052
rect -1458 14030 -1454 14052
rect -1434 14030 -1430 14052
rect -1410 14030 -1406 14052
rect -1397 14045 -1392 14052
rect -1386 14045 -1382 14052
rect -1387 14031 -1382 14045
rect -1386 14030 -1382 14031
rect -1362 14030 -1358 14148
rect -1338 14030 -1334 14148
rect -1314 14030 -1310 14148
rect -1290 14030 -1286 14148
rect -1266 14030 -1262 14148
rect -1242 14030 -1238 14148
rect -1218 14030 -1214 14148
rect -1194 14030 -1190 14148
rect -1170 14030 -1166 14148
rect -1146 14030 -1142 14148
rect -1122 14030 -1118 14148
rect -1098 14030 -1094 14148
rect -1074 14030 -1070 14148
rect -1050 14030 -1046 14148
rect -1026 14030 -1022 14148
rect -1002 14030 -998 14148
rect -978 14030 -974 14148
rect -954 14030 -950 14148
rect -930 14030 -926 14148
rect -906 14030 -902 14148
rect -882 14030 -878 14148
rect -858 14030 -854 14148
rect -834 14030 -830 14148
rect -810 14030 -806 14148
rect -786 14030 -782 14148
rect -762 14030 -758 14148
rect -738 14030 -734 14148
rect -714 14030 -710 14148
rect -690 14030 -686 14148
rect -666 14030 -662 14148
rect -642 14030 -638 14148
rect -618 14030 -614 14148
rect -594 14030 -590 14148
rect -570 14030 -566 14148
rect -546 14030 -542 14148
rect -522 14030 -518 14148
rect -498 14030 -494 14148
rect -474 14030 -470 14148
rect -450 14030 -446 14148
rect -426 14030 -422 14148
rect -402 14030 -398 14148
rect -378 14030 -374 14148
rect -354 14030 -350 14148
rect -330 14030 -326 14148
rect -306 14030 -302 14148
rect -282 14030 -278 14148
rect -258 14030 -254 14148
rect -234 14030 -230 14148
rect -210 14030 -206 14148
rect -186 14030 -182 14148
rect -162 14030 -158 14148
rect -138 14030 -134 14148
rect -114 14030 -110 14148
rect -90 14030 -86 14148
rect -66 14030 -62 14148
rect -42 14030 -38 14148
rect -18 14030 -14 14148
rect 6 14030 10 14148
rect 30 14030 34 14148
rect 54 14030 58 14148
rect 78 14030 82 14148
rect 102 14030 106 14148
rect 126 14030 130 14148
rect 150 14030 154 14148
rect 174 14030 178 14148
rect 198 14030 202 14148
rect 222 14030 226 14148
rect 246 14030 250 14148
rect 270 14030 274 14148
rect 294 14030 298 14148
rect 318 14030 322 14148
rect 342 14030 346 14148
rect 366 14030 370 14148
rect 390 14030 394 14148
rect 414 14030 418 14148
rect 438 14030 442 14148
rect 462 14030 466 14148
rect 475 14141 480 14148
rect 486 14141 490 14148
rect 493 14147 507 14148
rect 510 14147 517 14195
rect 485 14127 490 14141
rect 486 14030 490 14127
rect 510 14075 514 14147
rect 510 14051 517 14075
rect 510 14030 514 14051
rect 534 14030 538 14196
rect 558 14030 562 14196
rect 582 14030 586 14196
rect 606 14030 610 14196
rect 630 14030 634 14196
rect 654 14030 658 14196
rect 678 14030 682 14196
rect 702 14030 706 14196
rect 726 14030 730 14196
rect 750 14030 754 14196
rect 774 14030 778 14196
rect 798 14030 802 14196
rect 822 14030 826 14196
rect 846 14030 850 14196
rect 870 14030 874 14196
rect 894 14030 898 14196
rect 918 14030 922 14196
rect 942 14030 946 14196
rect 966 14031 970 14196
rect 979 14117 984 14127
rect 990 14117 994 14196
rect 989 14103 994 14117
rect 979 14102 1013 14103
rect 1014 14102 1018 14196
rect 1038 14102 1042 14196
rect 1062 14102 1066 14196
rect 1086 14102 1090 14196
rect 1110 14102 1114 14196
rect 1134 14102 1138 14196
rect 1158 14102 1162 14196
rect 1182 14102 1186 14196
rect 1206 14102 1210 14196
rect 1230 14102 1234 14196
rect 1254 14102 1258 14196
rect 1278 14102 1282 14196
rect 1302 14102 1306 14196
rect 1326 14102 1330 14196
rect 1350 14102 1354 14196
rect 1374 14102 1378 14196
rect 1398 14102 1402 14196
rect 1422 14102 1426 14196
rect 1446 14102 1450 14196
rect 1470 14102 1474 14196
rect 1494 14102 1498 14196
rect 1518 14102 1522 14196
rect 1542 14102 1546 14196
rect 1566 14102 1570 14196
rect 1590 14102 1594 14196
rect 1614 14102 1618 14196
rect 1638 14102 1642 14196
rect 1662 14102 1666 14196
rect 1686 14102 1690 14196
rect 1710 14102 1714 14196
rect 1734 14102 1738 14196
rect 1758 14102 1762 14196
rect 1782 14102 1786 14196
rect 1806 14102 1810 14196
rect 1830 14102 1834 14196
rect 1854 14102 1858 14196
rect 1878 14102 1882 14196
rect 1902 14102 1906 14196
rect 1926 14102 1930 14196
rect 1950 14102 1954 14196
rect 1974 14102 1978 14196
rect 1998 14102 2002 14196
rect 2022 14102 2026 14196
rect 2046 14102 2050 14196
rect 2070 14102 2074 14196
rect 2094 14102 2098 14196
rect 2118 14102 2122 14196
rect 2142 14102 2146 14196
rect 2166 14102 2170 14196
rect 2190 14102 2194 14196
rect 2214 14102 2218 14196
rect 2238 14102 2242 14196
rect 2262 14102 2266 14196
rect 2286 14102 2290 14196
rect 2310 14102 2314 14196
rect 2334 14102 2338 14196
rect 2358 14102 2362 14196
rect 2382 14102 2386 14196
rect 2406 14102 2410 14196
rect 2430 14102 2434 14196
rect 2454 14102 2458 14196
rect 2478 14102 2482 14196
rect 2502 14102 2506 14196
rect 2526 14102 2530 14196
rect 2550 14102 2554 14196
rect 2574 14102 2578 14196
rect 2598 14102 2602 14196
rect 2622 14102 2626 14196
rect 2646 14102 2650 14196
rect 2670 14102 2674 14196
rect 2694 14102 2698 14196
rect 2718 14102 2722 14196
rect 2742 14102 2746 14196
rect 2766 14102 2770 14196
rect 2790 14102 2794 14196
rect 2814 14102 2818 14196
rect 2838 14102 2842 14196
rect 2862 14102 2866 14196
rect 2886 14102 2890 14196
rect 2910 14102 2914 14196
rect 2934 14102 2938 14196
rect 2958 14102 2962 14196
rect 2982 14102 2986 14196
rect 3006 14102 3010 14196
rect 3030 14102 3034 14196
rect 3054 14102 3058 14196
rect 3078 14102 3082 14196
rect 3102 14102 3106 14196
rect 3126 14102 3130 14196
rect 3150 14102 3154 14196
rect 3174 14102 3178 14196
rect 3198 14102 3202 14196
rect 3222 14102 3226 14196
rect 3246 14102 3250 14196
rect 3270 14102 3274 14196
rect 3294 14171 3298 14196
rect 3294 14123 3301 14171
rect 3294 14102 3298 14123
rect 3318 14102 3322 14196
rect 3342 14102 3346 14196
rect 3366 14102 3370 14196
rect 3390 14102 3394 14196
rect 3414 14102 3418 14196
rect 3438 14102 3442 14196
rect 3462 14102 3466 14196
rect 3486 14102 3490 14196
rect 3510 14102 3514 14196
rect 3534 14102 3538 14196
rect 3558 14102 3562 14196
rect 3582 14102 3586 14196
rect 3606 14102 3610 14196
rect 3630 14102 3634 14196
rect 3643 14189 3648 14196
rect 3661 14195 3675 14196
rect 3653 14175 3658 14189
rect 3654 14103 3658 14175
rect 3643 14102 3675 14103
rect 979 14100 3675 14102
rect 979 14093 984 14100
rect 989 14079 994 14093
rect 955 14030 989 14031
rect -2032 14028 989 14030
rect -2371 13958 -2366 14028
rect -2348 13958 -2343 14028
rect -2325 14024 -2320 14028
rect -2309 14026 -2301 14028
rect -2317 14024 -2309 14026
rect -2325 14012 -2317 14024
rect -2052 14022 -2036 14024
rect -2052 14020 -2032 14022
rect -2062 14014 -2032 14020
rect -2325 13958 -2320 14012
rect -2317 14010 -2309 14012
rect -2092 13998 -2062 14000
rect -2094 13994 -2062 13998
rect -2309 13964 -2301 13970
rect -2317 13958 -2309 13964
rect -2000 13958 -1992 14028
rect -1904 14021 -1874 14028
rect -1842 14021 -1806 14028
rect -1655 14026 -1647 14028
rect -1663 14024 -1655 14026
rect -1842 14014 -1680 14020
rect -1671 14012 -1663 14024
rect -1663 14010 -1655 14012
rect -1854 13998 -1806 14000
rect -1854 13994 -1680 13998
rect -1655 13964 -1647 13970
rect -1663 13958 -1655 13964
rect -1642 13958 -1637 14028
rect -1619 13958 -1614 14028
rect -1530 13958 -1526 14028
rect -1506 13958 -1502 14028
rect -1482 13958 -1478 14028
rect -1458 13958 -1454 14028
rect -1434 13958 -1430 14028
rect -1410 13958 -1406 14028
rect -1386 13958 -1382 14028
rect -1362 13979 -1358 14028
rect -2393 13956 -1365 13958
rect -2371 13862 -2366 13956
rect -2348 13862 -2343 13956
rect -2325 13894 -2320 13956
rect -2317 13954 -2309 13956
rect -2000 13955 -1966 13956
rect -2000 13954 -1982 13955
rect -1663 13954 -1655 13956
rect -2028 13946 -2018 13948
rect -2309 13936 -2301 13942
rect -2091 13936 -2061 13943
rect -2317 13926 -2309 13936
rect -2044 13934 -2028 13936
rect -2026 13934 -2014 13946
rect -2084 13928 -2061 13934
rect -2044 13932 -2014 13934
rect -2292 13918 -2054 13927
rect -2325 13886 -2317 13894
rect -2325 13866 -2320 13886
rect -2317 13878 -2309 13886
rect -2325 13862 -2317 13866
rect -2095 13864 -2083 13868
rect -2000 13865 -1992 13954
rect -1982 13953 -1966 13954
rect -1980 13936 -1932 13943
rect -1655 13936 -1647 13942
rect -1846 13918 -1680 13927
rect -1663 13926 -1655 13936
rect -1671 13886 -1663 13894
rect -1663 13878 -1655 13886
rect -2119 13862 -2069 13864
rect -2053 13862 -1972 13865
rect -1926 13862 -1892 13865
rect -1671 13862 -1663 13866
rect -1642 13862 -1637 13956
rect -1619 13862 -1614 13956
rect -1530 13862 -1526 13956
rect -1506 13862 -1502 13956
rect -1482 13862 -1478 13956
rect -1458 13862 -1454 13956
rect -1434 13862 -1430 13956
rect -1410 13862 -1406 13956
rect -1386 13862 -1382 13956
rect -1379 13955 -1365 13956
rect -1362 13955 -1355 13979
rect -1362 13862 -1358 13955
rect -1338 13862 -1334 14028
rect -1314 13862 -1310 14028
rect -1290 13862 -1286 14028
rect -1266 13862 -1262 14028
rect -1242 13862 -1238 14028
rect -1218 13862 -1214 14028
rect -1194 13862 -1190 14028
rect -1170 13862 -1166 14028
rect -1146 13862 -1142 14028
rect -1122 13862 -1118 14028
rect -1098 13862 -1094 14028
rect -1074 13862 -1070 14028
rect -1050 13862 -1046 14028
rect -1026 13862 -1022 14028
rect -1002 13862 -998 14028
rect -978 13862 -974 14028
rect -954 13862 -950 14028
rect -930 13862 -926 14028
rect -906 13862 -902 14028
rect -882 13862 -878 14028
rect -858 13862 -854 14028
rect -834 13862 -830 14028
rect -810 13862 -806 14028
rect -786 13862 -782 14028
rect -762 13862 -758 14028
rect -738 13862 -734 14028
rect -714 13862 -710 14028
rect -690 13862 -686 14028
rect -666 13862 -662 14028
rect -642 13862 -638 14028
rect -618 13862 -614 14028
rect -594 13862 -590 14028
rect -570 13862 -566 14028
rect -546 13862 -542 14028
rect -522 13862 -518 14028
rect -498 13862 -494 14028
rect -474 13862 -470 14028
rect -450 13862 -446 14028
rect -426 13862 -422 14028
rect -402 13862 -398 14028
rect -378 13862 -374 14028
rect -354 13862 -350 14028
rect -330 13862 -326 14028
rect -306 13862 -302 14028
rect -282 13862 -278 14028
rect -258 13862 -254 14028
rect -234 13862 -230 14028
rect -210 13862 -206 14028
rect -186 13862 -182 14028
rect -162 13862 -158 14028
rect -138 13862 -134 14028
rect -114 13862 -110 14028
rect -90 13862 -86 14028
rect -66 13862 -62 14028
rect -42 13862 -38 14028
rect -18 13862 -14 14028
rect 6 13862 10 14028
rect 30 13862 34 14028
rect 54 13862 58 14028
rect 78 13862 82 14028
rect 102 13862 106 14028
rect 126 13862 130 14028
rect 150 13862 154 14028
rect 174 13862 178 14028
rect 198 13862 202 14028
rect 222 13862 226 14028
rect 246 13862 250 14028
rect 270 13862 274 14028
rect 294 13862 298 14028
rect 318 13862 322 14028
rect 342 13862 346 14028
rect 366 13862 370 14028
rect 390 13862 394 14028
rect 414 13862 418 14028
rect 438 13862 442 14028
rect 462 13862 466 14028
rect 486 13862 490 14028
rect 510 13862 514 14028
rect 534 13862 538 14028
rect 558 13862 562 14028
rect 582 13862 586 14028
rect 606 13862 610 14028
rect 630 13862 634 14028
rect 654 13862 658 14028
rect 678 13862 682 14028
rect 702 13862 706 14028
rect 726 13862 730 14028
rect 750 13862 754 14028
rect 774 13862 778 14028
rect 798 13862 802 14028
rect 822 13862 826 14028
rect 846 13862 850 14028
rect 870 13862 874 14028
rect 894 13862 898 14028
rect 918 13862 922 14028
rect 942 13862 946 14028
rect 955 14021 960 14028
rect 966 14021 970 14028
rect 965 14007 970 14021
rect 966 13862 970 14007
rect 990 13955 994 14079
rect 1014 14051 1018 14100
rect 1014 14003 1021 14051
rect 990 13931 997 13955
rect 990 13862 994 13931
rect 1014 13862 1018 14003
rect 1038 13862 1042 14100
rect 1062 13862 1066 14100
rect 1086 13862 1090 14100
rect 1110 13862 1114 14100
rect 1134 13862 1138 14100
rect 1158 13862 1162 14100
rect 1182 13862 1186 14100
rect 1206 13862 1210 14100
rect 1230 13862 1234 14100
rect 1254 13862 1258 14100
rect 1278 13862 1282 14100
rect 1302 13862 1306 14100
rect 1326 13862 1330 14100
rect 1350 13862 1354 14100
rect 1374 13862 1378 14100
rect 1398 13862 1402 14100
rect 1422 13862 1426 14100
rect 1446 13862 1450 14100
rect 1470 13862 1474 14100
rect 1494 13862 1498 14100
rect 1518 13862 1522 14100
rect 1542 13862 1546 14100
rect 1566 13862 1570 14100
rect 1590 13862 1594 14100
rect 1614 13862 1618 14100
rect 1638 13862 1642 14100
rect 1662 13862 1666 14100
rect 1686 13862 1690 14100
rect 1710 13862 1714 14100
rect 1734 13862 1738 14100
rect 1758 13862 1762 14100
rect 1771 13901 1776 13911
rect 1782 13901 1786 14100
rect 1781 13887 1786 13901
rect 1782 13862 1786 13887
rect 1806 13862 1810 14100
rect 1830 13862 1834 14100
rect 1854 13862 1858 14100
rect 1878 13862 1882 14100
rect 1902 13862 1906 14100
rect 1926 13862 1930 14100
rect 1950 13862 1954 14100
rect 1974 13862 1978 14100
rect 1998 13862 2002 14100
rect 2022 13862 2026 14100
rect 2046 13862 2050 14100
rect 2070 13862 2074 14100
rect 2094 13862 2098 14100
rect 2118 13862 2122 14100
rect 2142 13862 2146 14100
rect 2166 13862 2170 14100
rect 2190 13862 2194 14100
rect 2214 13862 2218 14100
rect 2238 13862 2242 14100
rect 2262 13862 2266 14100
rect 2286 13862 2290 14100
rect 2310 13862 2314 14100
rect 2334 13862 2338 14100
rect 2358 13862 2362 14100
rect 2382 13862 2386 14100
rect 2406 13862 2410 14100
rect 2430 13862 2434 14100
rect 2454 13862 2458 14100
rect 2478 13862 2482 14100
rect 2502 13862 2506 14100
rect 2526 13862 2530 14100
rect 2550 13862 2554 14100
rect 2574 13862 2578 14100
rect 2598 13862 2602 14100
rect 2622 13862 2626 14100
rect 2646 13862 2650 14100
rect 2670 13862 2674 14100
rect 2694 13862 2698 14100
rect 2718 13862 2722 14100
rect 2742 13862 2746 14100
rect 2766 13862 2770 14100
rect 2790 13862 2794 14100
rect 2814 13862 2818 14100
rect 2838 13862 2842 14100
rect 2862 13862 2866 14100
rect 2886 13862 2890 14100
rect 2910 13862 2914 14100
rect 2934 13862 2938 14100
rect 2958 13862 2962 14100
rect 2982 13862 2986 14100
rect 3006 13862 3010 14100
rect 3030 13862 3034 14100
rect 3054 13862 3058 14100
rect 3078 13862 3082 14100
rect 3102 13862 3106 14100
rect 3126 13862 3130 14100
rect 3150 13862 3154 14100
rect 3174 13862 3178 14100
rect 3198 13862 3202 14100
rect 3222 13862 3226 14100
rect 3246 13862 3250 14100
rect 3270 13862 3274 14100
rect 3294 13862 3298 14100
rect 3318 13862 3322 14100
rect 3342 13862 3346 14100
rect 3366 13862 3370 14100
rect 3390 13862 3394 14100
rect 3414 13862 3418 14100
rect 3438 13862 3442 14100
rect 3462 13862 3466 14100
rect 3486 13862 3490 14100
rect 3510 13862 3514 14100
rect 3534 13862 3538 14100
rect 3558 13862 3562 14100
rect 3582 13862 3586 14100
rect 3606 13862 3610 14100
rect 3630 13862 3634 14100
rect 3643 14093 3648 14100
rect 3654 14093 3658 14100
rect 3661 14099 3675 14100
rect 3653 14079 3658 14093
rect 3643 14069 3648 14079
rect 3653 14055 3658 14069
rect 3654 13862 3658 14055
rect 3667 13949 3672 13959
rect 3677 13935 3682 13949
rect 3678 13862 3682 13935
rect 3691 13862 3699 13863
rect -2393 13860 3699 13862
rect -2371 13814 -2366 13860
rect -2348 13814 -2343 13860
rect -2325 13856 -2317 13860
rect -2325 13838 -2320 13856
rect -2317 13850 -2309 13856
rect -2095 13854 -2083 13860
rect -2053 13858 -1972 13860
rect -2083 13852 -2079 13854
rect -2079 13851 -2067 13852
rect -2079 13850 -2043 13851
rect -2091 13846 -2043 13850
rect -2000 13846 -1992 13858
rect -1671 13856 -1663 13860
rect -1982 13846 -1916 13851
rect -1663 13850 -1655 13856
rect -2091 13845 -2018 13846
rect -2091 13843 -2067 13845
rect -2053 13843 -2018 13845
rect -2002 13845 -1916 13846
rect -2002 13843 -1972 13845
rect -1924 13843 -1916 13845
rect -2079 13841 -2067 13843
rect -2000 13842 -1992 13843
rect -2325 13828 -2317 13838
rect -2112 13837 -2096 13841
rect -2083 13838 -2079 13841
rect -2027 13840 -1992 13842
rect -2109 13836 -2096 13837
rect -2112 13829 -2096 13836
rect -2083 13829 -2053 13836
rect -2018 13832 -2017 13840
rect -2023 13830 -2017 13832
rect -2009 13832 -2002 13835
rect -2009 13830 -2003 13832
rect -2109 13828 -2096 13829
rect -2325 13814 -2320 13828
rect -2317 13822 -2309 13828
rect -2112 13825 -2096 13828
rect -2017 13819 -2003 13830
rect -2017 13818 -2009 13819
rect -2074 13814 -2040 13816
rect -2000 13814 -1992 13840
rect -1972 13829 -1924 13836
rect -1671 13828 -1663 13838
rect -1663 13822 -1655 13828
rect -1642 13814 -1637 13860
rect -1619 13814 -1614 13860
rect -1530 13814 -1526 13860
rect -1506 13814 -1502 13860
rect -1482 13814 -1478 13860
rect -1458 13814 -1454 13860
rect -1434 13814 -1430 13860
rect -1410 13814 -1406 13860
rect -1386 13814 -1382 13860
rect -1362 13814 -1358 13860
rect -1338 13814 -1334 13860
rect -1314 13814 -1310 13860
rect -1290 13814 -1286 13860
rect -1266 13814 -1262 13860
rect -1242 13814 -1238 13860
rect -1218 13814 -1214 13860
rect -1194 13814 -1190 13860
rect -1170 13814 -1166 13860
rect -1146 13814 -1142 13860
rect -1122 13814 -1118 13860
rect -1098 13814 -1094 13860
rect -1074 13814 -1070 13860
rect -1050 13814 -1046 13860
rect -1026 13814 -1022 13860
rect -1002 13814 -998 13860
rect -978 13814 -974 13860
rect -954 13814 -950 13860
rect -930 13814 -926 13860
rect -906 13814 -902 13860
rect -882 13814 -878 13860
rect -858 13814 -854 13860
rect -834 13814 -830 13860
rect -810 13814 -806 13860
rect -786 13814 -782 13860
rect -762 13814 -758 13860
rect -738 13814 -734 13860
rect -714 13814 -710 13860
rect -690 13814 -686 13860
rect -666 13814 -662 13860
rect -642 13814 -638 13860
rect -618 13814 -614 13860
rect -594 13814 -590 13860
rect -570 13814 -566 13860
rect -546 13814 -542 13860
rect -522 13814 -518 13860
rect -498 13814 -494 13860
rect -474 13814 -470 13860
rect -450 13814 -446 13860
rect -426 13814 -422 13860
rect -402 13814 -398 13860
rect -378 13814 -374 13860
rect -354 13814 -350 13860
rect -330 13814 -326 13860
rect -306 13814 -302 13860
rect -282 13814 -278 13860
rect -258 13814 -254 13860
rect -234 13814 -230 13860
rect -210 13814 -206 13860
rect -186 13814 -182 13860
rect -162 13814 -158 13860
rect -138 13814 -134 13860
rect -114 13814 -110 13860
rect -90 13814 -86 13860
rect -66 13814 -62 13860
rect -42 13814 -38 13860
rect -18 13814 -14 13860
rect 6 13814 10 13860
rect 30 13814 34 13860
rect 54 13814 58 13860
rect 78 13814 82 13860
rect 102 13815 106 13860
rect 91 13814 125 13815
rect -2393 13812 125 13814
rect -2371 13766 -2366 13812
rect -2348 13766 -2343 13812
rect -2325 13810 -2320 13812
rect -2325 13800 -2317 13810
rect -2325 13780 -2320 13800
rect -2317 13794 -2309 13800
rect -2325 13772 -2317 13780
rect -2101 13775 -2071 13778
rect -2325 13766 -2320 13772
rect -2317 13766 -2309 13772
rect -2000 13770 -1992 13812
rect -1671 13800 -1663 13810
rect -1663 13794 -1655 13800
rect -1854 13784 -1680 13788
rect -1846 13775 -1798 13778
rect -2079 13769 -2043 13770
rect -2007 13769 -1991 13770
rect -2079 13768 -2071 13769
rect -2079 13766 -2029 13768
rect -2011 13766 -1991 13769
rect -1846 13767 -1806 13773
rect -1671 13772 -1663 13780
rect -1864 13766 -1796 13767
rect -1663 13766 -1655 13772
rect -1642 13766 -1637 13812
rect -1619 13766 -1614 13812
rect -1530 13766 -1526 13812
rect -1506 13766 -1502 13812
rect -1482 13766 -1478 13812
rect -1458 13766 -1454 13812
rect -1434 13766 -1430 13812
rect -1410 13766 -1406 13812
rect -1386 13766 -1382 13812
rect -1362 13766 -1358 13812
rect -1338 13766 -1334 13812
rect -1314 13766 -1310 13812
rect -1290 13766 -1286 13812
rect -1266 13766 -1262 13812
rect -1242 13766 -1238 13812
rect -1218 13766 -1214 13812
rect -1194 13766 -1190 13812
rect -1170 13766 -1166 13812
rect -1146 13766 -1142 13812
rect -1122 13766 -1118 13812
rect -1098 13766 -1094 13812
rect -1074 13766 -1070 13812
rect -1050 13766 -1046 13812
rect -1026 13766 -1022 13812
rect -1002 13766 -998 13812
rect -978 13766 -974 13812
rect -954 13766 -950 13812
rect -930 13766 -926 13812
rect -906 13766 -902 13812
rect -882 13766 -878 13812
rect -858 13766 -854 13812
rect -834 13766 -830 13812
rect -810 13766 -806 13812
rect -786 13766 -782 13812
rect -762 13766 -758 13812
rect -738 13766 -734 13812
rect -714 13766 -710 13812
rect -690 13766 -686 13812
rect -666 13766 -662 13812
rect -642 13766 -638 13812
rect -618 13766 -614 13812
rect -594 13766 -590 13812
rect -570 13766 -566 13812
rect -546 13766 -542 13812
rect -522 13766 -518 13812
rect -498 13766 -494 13812
rect -474 13767 -470 13812
rect -485 13766 -451 13767
rect -2393 13764 -451 13766
rect -2371 13718 -2366 13764
rect -2348 13718 -2343 13764
rect -2325 13752 -2320 13764
rect -2079 13762 -2071 13764
rect -2072 13760 -2071 13762
rect -2109 13755 -2101 13760
rect -2101 13753 -2079 13755
rect -2069 13753 -2068 13760
rect -2325 13744 -2317 13752
rect -2079 13748 -2071 13753
rect -2325 13724 -2320 13744
rect -2317 13736 -2309 13744
rect -2074 13739 -2071 13748
rect -2069 13744 -2068 13748
rect -2109 13730 -2079 13733
rect -2325 13718 -2317 13724
rect -2080 13718 -2071 13719
rect -2000 13718 -1992 13764
rect -1846 13762 -1806 13764
rect -1854 13757 -1806 13761
rect -1854 13755 -1846 13757
rect -1846 13753 -1806 13755
rect -1806 13751 -1798 13753
rect -1846 13748 -1798 13751
rect -1846 13735 -1806 13746
rect -1671 13744 -1663 13752
rect -1663 13736 -1655 13744
rect -1854 13730 -1680 13734
rect -1926 13718 -1892 13721
rect -1671 13718 -1663 13724
rect -1642 13718 -1637 13764
rect -1619 13718 -1614 13764
rect -1530 13718 -1526 13764
rect -1506 13718 -1502 13764
rect -1482 13718 -1478 13764
rect -1458 13718 -1454 13764
rect -1434 13718 -1430 13764
rect -1410 13718 -1406 13764
rect -1386 13718 -1382 13764
rect -1362 13718 -1358 13764
rect -1338 13718 -1334 13764
rect -1314 13718 -1310 13764
rect -1290 13718 -1286 13764
rect -1266 13718 -1262 13764
rect -1242 13718 -1238 13764
rect -1218 13718 -1214 13764
rect -1194 13718 -1190 13764
rect -1170 13718 -1166 13764
rect -1146 13718 -1142 13764
rect -1122 13718 -1118 13764
rect -1098 13718 -1094 13764
rect -1074 13718 -1070 13764
rect -1050 13718 -1046 13764
rect -1026 13718 -1022 13764
rect -1002 13718 -998 13764
rect -978 13718 -974 13764
rect -954 13718 -950 13764
rect -930 13718 -926 13764
rect -906 13718 -902 13764
rect -882 13718 -878 13764
rect -858 13718 -854 13764
rect -834 13718 -830 13764
rect -810 13718 -806 13764
rect -786 13718 -782 13764
rect -762 13718 -758 13764
rect -738 13718 -734 13764
rect -714 13718 -710 13764
rect -690 13718 -686 13764
rect -666 13718 -662 13764
rect -642 13718 -638 13764
rect -618 13718 -614 13764
rect -594 13718 -590 13764
rect -570 13718 -566 13764
rect -546 13718 -542 13764
rect -522 13718 -518 13764
rect -498 13718 -494 13764
rect -485 13757 -480 13764
rect -474 13757 -470 13764
rect -475 13743 -470 13757
rect -485 13742 -451 13743
rect -450 13742 -446 13812
rect -426 13742 -422 13812
rect -402 13742 -398 13812
rect -378 13742 -374 13812
rect -354 13742 -350 13812
rect -330 13742 -326 13812
rect -306 13742 -302 13812
rect -282 13742 -278 13812
rect -258 13742 -254 13812
rect -234 13742 -230 13812
rect -210 13742 -206 13812
rect -186 13742 -182 13812
rect -162 13742 -158 13812
rect -138 13742 -134 13812
rect -114 13742 -110 13812
rect -90 13742 -86 13812
rect -77 13781 -72 13791
rect -66 13781 -62 13812
rect -67 13767 -62 13781
rect -77 13766 -43 13767
rect -42 13766 -38 13812
rect -18 13766 -14 13812
rect 6 13766 10 13812
rect 30 13766 34 13812
rect 54 13766 58 13812
rect 78 13766 82 13812
rect 91 13805 96 13812
rect 102 13805 106 13812
rect 101 13791 106 13805
rect 91 13781 96 13791
rect 101 13767 106 13781
rect 102 13766 106 13767
rect 126 13766 130 13860
rect 150 13766 154 13860
rect 174 13766 178 13860
rect 198 13766 202 13860
rect 222 13766 226 13860
rect 246 13766 250 13860
rect 270 13766 274 13860
rect 294 13766 298 13860
rect 318 13766 322 13860
rect 342 13766 346 13860
rect 366 13766 370 13860
rect 390 13766 394 13860
rect 414 13766 418 13860
rect 438 13766 442 13860
rect 462 13766 466 13860
rect 486 13766 490 13860
rect 510 13766 514 13860
rect 534 13766 538 13860
rect 558 13766 562 13860
rect 571 13829 576 13839
rect 582 13829 586 13860
rect 581 13815 586 13829
rect 571 13814 605 13815
rect 606 13814 610 13860
rect 630 13814 634 13860
rect 654 13814 658 13860
rect 678 13814 682 13860
rect 702 13814 706 13860
rect 726 13814 730 13860
rect 750 13814 754 13860
rect 774 13814 778 13860
rect 798 13814 802 13860
rect 822 13814 826 13860
rect 846 13814 850 13860
rect 870 13814 874 13860
rect 894 13814 898 13860
rect 918 13814 922 13860
rect 942 13814 946 13860
rect 966 13814 970 13860
rect 990 13814 994 13860
rect 1014 13814 1018 13860
rect 1038 13814 1042 13860
rect 1062 13814 1066 13860
rect 1086 13814 1090 13860
rect 1110 13814 1114 13860
rect 1134 13814 1138 13860
rect 1158 13814 1162 13860
rect 1182 13814 1186 13860
rect 1206 13814 1210 13860
rect 1230 13814 1234 13860
rect 1254 13814 1258 13860
rect 1278 13814 1282 13860
rect 1302 13814 1306 13860
rect 1326 13814 1330 13860
rect 1350 13814 1354 13860
rect 1374 13814 1378 13860
rect 1398 13814 1402 13860
rect 1422 13814 1426 13860
rect 1446 13814 1450 13860
rect 1470 13814 1474 13860
rect 1494 13814 1498 13860
rect 1518 13814 1522 13860
rect 1542 13814 1546 13860
rect 1566 13814 1570 13860
rect 1590 13814 1594 13860
rect 1614 13814 1618 13860
rect 1638 13814 1642 13860
rect 1662 13814 1666 13860
rect 1686 13814 1690 13860
rect 1710 13814 1714 13860
rect 1734 13814 1738 13860
rect 1758 13814 1762 13860
rect 1782 13814 1786 13860
rect 1806 13835 1810 13860
rect 571 13812 1803 13814
rect 571 13805 576 13812
rect 581 13791 586 13805
rect 582 13766 586 13791
rect 606 13766 610 13812
rect 630 13766 634 13812
rect 654 13766 658 13812
rect 678 13766 682 13812
rect 702 13766 706 13812
rect 726 13766 730 13812
rect 750 13766 754 13812
rect 774 13766 778 13812
rect 798 13766 802 13812
rect 822 13766 826 13812
rect 846 13766 850 13812
rect 870 13766 874 13812
rect 894 13766 898 13812
rect 918 13766 922 13812
rect 942 13766 946 13812
rect 966 13766 970 13812
rect 990 13766 994 13812
rect 1014 13766 1018 13812
rect 1038 13766 1042 13812
rect 1062 13766 1066 13812
rect 1086 13766 1090 13812
rect 1110 13766 1114 13812
rect 1134 13766 1138 13812
rect 1158 13766 1162 13812
rect 1182 13766 1186 13812
rect 1206 13766 1210 13812
rect 1230 13766 1234 13812
rect 1254 13766 1258 13812
rect 1278 13766 1282 13812
rect 1302 13766 1306 13812
rect 1326 13766 1330 13812
rect 1350 13766 1354 13812
rect 1374 13766 1378 13812
rect 1398 13766 1402 13812
rect 1422 13766 1426 13812
rect 1446 13766 1450 13812
rect 1470 13766 1474 13812
rect 1494 13766 1498 13812
rect 1518 13766 1522 13812
rect 1542 13766 1546 13812
rect 1566 13766 1570 13812
rect 1590 13766 1594 13812
rect 1614 13766 1618 13812
rect 1638 13766 1642 13812
rect 1662 13766 1666 13812
rect 1686 13766 1690 13812
rect 1710 13766 1714 13812
rect 1734 13766 1738 13812
rect 1758 13766 1762 13812
rect 1782 13766 1786 13812
rect 1789 13811 1803 13812
rect 1806 13811 1813 13835
rect 1806 13766 1810 13811
rect 1830 13766 1834 13860
rect 1854 13766 1858 13860
rect 1878 13766 1882 13860
rect 1902 13766 1906 13860
rect 1926 13766 1930 13860
rect 1950 13766 1954 13860
rect 1974 13766 1978 13860
rect 1998 13766 2002 13860
rect 2022 13766 2026 13860
rect 2046 13766 2050 13860
rect 2070 13766 2074 13860
rect 2094 13766 2098 13860
rect 2118 13766 2122 13860
rect 2142 13766 2146 13860
rect 2166 13766 2170 13860
rect 2190 13766 2194 13860
rect 2214 13766 2218 13860
rect 2238 13766 2242 13860
rect 2262 13766 2266 13860
rect 2286 13766 2290 13860
rect 2310 13766 2314 13860
rect 2334 13766 2338 13860
rect 2358 13766 2362 13860
rect 2382 13766 2386 13860
rect 2406 13766 2410 13860
rect 2430 13766 2434 13860
rect 2454 13766 2458 13860
rect 2478 13766 2482 13860
rect 2502 13766 2506 13860
rect 2526 13766 2530 13860
rect 2550 13766 2554 13860
rect 2574 13766 2578 13860
rect 2598 13766 2602 13860
rect 2622 13766 2626 13860
rect 2646 13766 2650 13860
rect 2670 13766 2674 13860
rect 2694 13766 2698 13860
rect 2718 13766 2722 13860
rect 2742 13766 2746 13860
rect 2766 13766 2770 13860
rect 2790 13766 2794 13860
rect 2814 13766 2818 13860
rect 2838 13766 2842 13860
rect 2862 13766 2866 13860
rect 2886 13766 2890 13860
rect 2910 13766 2914 13860
rect 2934 13766 2938 13860
rect 2958 13766 2962 13860
rect 2982 13766 2986 13860
rect 3006 13766 3010 13860
rect 3030 13766 3034 13860
rect 3054 13766 3058 13860
rect 3078 13766 3082 13860
rect 3102 13766 3106 13860
rect 3126 13766 3130 13860
rect 3150 13766 3154 13860
rect 3174 13766 3178 13860
rect 3198 13766 3202 13860
rect 3222 13766 3226 13860
rect 3246 13766 3250 13860
rect 3270 13766 3274 13860
rect 3294 13766 3298 13860
rect 3318 13766 3322 13860
rect 3342 13766 3346 13860
rect 3366 13766 3370 13860
rect 3390 13766 3394 13860
rect 3414 13766 3418 13860
rect 3438 13766 3442 13860
rect 3462 13766 3466 13860
rect 3486 13766 3490 13860
rect 3510 13766 3514 13860
rect 3534 13766 3538 13860
rect 3558 13766 3562 13860
rect 3582 13766 3586 13860
rect 3606 13766 3610 13860
rect 3630 13766 3634 13860
rect 3654 13767 3658 13860
rect 3667 13781 3672 13791
rect 3678 13781 3682 13860
rect 3685 13859 3699 13860
rect 3691 13853 3696 13859
rect 3701 13839 3706 13853
rect 3691 13805 3696 13815
rect 3702 13805 3706 13839
rect 3701 13791 3706 13805
rect 3677 13767 3682 13781
rect 3643 13766 3677 13767
rect -77 13764 3677 13766
rect -77 13757 -72 13764
rect -67 13743 -62 13757
rect -66 13742 -62 13743
rect -42 13742 -38 13764
rect -18 13742 -14 13764
rect 6 13742 10 13764
rect 30 13742 34 13764
rect 54 13742 58 13764
rect 78 13742 82 13764
rect 102 13742 106 13764
rect 126 13742 130 13764
rect 150 13742 154 13764
rect 174 13742 178 13764
rect 198 13742 202 13764
rect 222 13742 226 13764
rect 246 13742 250 13764
rect 270 13742 274 13764
rect 294 13742 298 13764
rect 318 13742 322 13764
rect 342 13742 346 13764
rect 366 13742 370 13764
rect 390 13742 394 13764
rect 414 13742 418 13764
rect 438 13742 442 13764
rect 462 13742 466 13764
rect 486 13742 490 13764
rect 510 13742 514 13764
rect 534 13742 538 13764
rect 558 13742 562 13764
rect 582 13742 586 13764
rect 606 13763 610 13764
rect -485 13740 603 13742
rect -485 13733 -480 13740
rect -475 13719 -470 13733
rect -474 13718 -470 13719
rect -450 13718 -446 13740
rect -426 13718 -422 13740
rect -402 13718 -398 13740
rect -378 13718 -374 13740
rect -354 13718 -350 13740
rect -330 13718 -326 13740
rect -306 13718 -302 13740
rect -282 13718 -278 13740
rect -258 13718 -254 13740
rect -234 13718 -230 13740
rect -210 13718 -206 13740
rect -186 13718 -182 13740
rect -162 13718 -158 13740
rect -138 13718 -134 13740
rect -114 13718 -110 13740
rect -90 13718 -86 13740
rect -66 13718 -62 13740
rect -42 13718 -38 13740
rect -18 13718 -14 13740
rect 6 13718 10 13740
rect 30 13718 34 13740
rect 54 13718 58 13740
rect 78 13718 82 13740
rect 102 13718 106 13740
rect 126 13739 130 13740
rect -2393 13716 123 13718
rect -2371 13694 -2366 13716
rect -2348 13694 -2343 13716
rect -2325 13710 -2317 13716
rect -2325 13694 -2320 13710
rect -2317 13708 -2309 13710
rect -2309 13696 -2301 13708
rect -2080 13707 -2071 13716
rect -2068 13706 -2059 13707
rect -2068 13699 -2038 13706
rect -2317 13694 -2309 13696
rect -2068 13694 -2059 13699
rect -2000 13698 -1992 13716
rect -1846 13708 -1794 13716
rect -1671 13710 -1663 13716
rect -1663 13708 -1655 13710
rect -1852 13699 -1804 13706
rect -2011 13696 -1983 13698
rect -2025 13695 -1983 13696
rect -2025 13694 -1975 13695
rect -1846 13694 -1804 13697
rect -1655 13696 -1647 13708
rect -1663 13694 -1655 13696
rect -1642 13694 -1637 13716
rect -1619 13694 -1614 13716
rect -1530 13694 -1526 13716
rect -1506 13694 -1502 13716
rect -1482 13694 -1478 13716
rect -1458 13695 -1454 13716
rect -1469 13694 -1435 13695
rect -2393 13692 -1435 13694
rect -2371 13670 -2366 13692
rect -2348 13670 -2343 13692
rect -2325 13682 -2317 13692
rect -2068 13691 -2038 13692
rect -2068 13689 -2059 13691
rect -2013 13690 -1983 13692
rect -1846 13691 -1804 13692
rect -2000 13689 -1983 13690
rect -1862 13689 -1798 13690
rect -2076 13682 -2068 13689
rect -2061 13682 -2045 13684
rect -2038 13682 -2001 13689
rect -2325 13670 -2320 13682
rect -2317 13680 -2309 13682
rect -2309 13670 -2301 13680
rect -2068 13679 -2045 13682
rect -2015 13681 -2001 13682
rect -2068 13672 -2038 13679
rect -2068 13670 -2045 13672
rect -2000 13670 -1992 13689
rect -1985 13687 -1796 13689
rect -1985 13682 -1852 13687
rect -1846 13682 -1796 13687
rect -1671 13682 -1663 13692
rect -1846 13681 -1798 13682
rect -1663 13680 -1655 13682
rect -1852 13672 -1804 13679
rect -1976 13670 -1940 13671
rect -1655 13670 -1647 13680
rect -1642 13670 -1637 13692
rect -1619 13670 -1614 13692
rect -1530 13670 -1526 13692
rect -1506 13670 -1502 13692
rect -1482 13670 -1478 13692
rect -1469 13685 -1464 13692
rect -1458 13685 -1454 13692
rect -1459 13671 -1454 13685
rect -1469 13670 -1435 13671
rect -1434 13670 -1430 13716
rect -1410 13670 -1406 13716
rect -1386 13670 -1382 13716
rect -1362 13670 -1358 13716
rect -1338 13670 -1334 13716
rect -1314 13670 -1310 13716
rect -1290 13670 -1286 13716
rect -1266 13670 -1262 13716
rect -1242 13670 -1238 13716
rect -1218 13670 -1214 13716
rect -1194 13670 -1190 13716
rect -1170 13670 -1166 13716
rect -1146 13670 -1142 13716
rect -1122 13670 -1118 13716
rect -1098 13670 -1094 13716
rect -1074 13670 -1070 13716
rect -1050 13670 -1046 13716
rect -1026 13670 -1022 13716
rect -1002 13670 -998 13716
rect -978 13670 -974 13716
rect -954 13670 -950 13716
rect -930 13670 -926 13716
rect -906 13670 -902 13716
rect -882 13670 -878 13716
rect -858 13670 -854 13716
rect -834 13670 -830 13716
rect -810 13670 -806 13716
rect -786 13670 -782 13716
rect -762 13670 -758 13716
rect -738 13670 -734 13716
rect -714 13670 -710 13716
rect -690 13670 -686 13716
rect -666 13670 -662 13716
rect -642 13670 -638 13716
rect -618 13671 -614 13716
rect -629 13670 -595 13671
rect -2393 13668 -595 13670
rect -2371 13598 -2366 13668
rect -2348 13598 -2343 13668
rect -2325 13666 -2320 13668
rect -2317 13666 -2309 13668
rect -2325 13654 -2317 13666
rect -2068 13662 -2059 13668
rect -2076 13655 -2071 13662
rect -2068 13654 -2059 13655
rect -2325 13634 -2320 13654
rect -2317 13652 -2309 13654
rect -2325 13626 -2317 13634
rect -2060 13628 -2030 13631
rect -2325 13606 -2320 13626
rect -2317 13618 -2309 13626
rect -2060 13615 -2038 13626
rect -2033 13619 -2030 13628
rect -2028 13624 -2027 13628
rect -2068 13610 -2038 13613
rect -2325 13598 -2317 13606
rect -2000 13598 -1992 13668
rect -1846 13664 -1804 13668
rect -1663 13666 -1655 13668
rect -1846 13654 -1794 13663
rect -1671 13654 -1663 13666
rect -1663 13652 -1655 13654
rect -1912 13643 -1884 13645
rect -1852 13637 -1804 13641
rect -1844 13628 -1796 13631
rect -1671 13626 -1663 13634
rect -1844 13615 -1804 13626
rect -1663 13618 -1655 13626
rect -1852 13610 -1680 13614
rect -1926 13598 -1892 13601
rect -1671 13598 -1663 13606
rect -1642 13598 -1637 13668
rect -1619 13598 -1614 13668
rect -1530 13598 -1526 13668
rect -1506 13598 -1502 13668
rect -1482 13598 -1478 13668
rect -1469 13661 -1464 13668
rect -1459 13647 -1454 13661
rect -1458 13598 -1454 13647
rect -1434 13619 -1430 13668
rect -2393 13596 -1437 13598
rect -2371 13574 -2366 13596
rect -2348 13574 -2343 13596
rect -2325 13590 -2317 13596
rect -2325 13574 -2320 13590
rect -2309 13578 -2301 13590
rect -2068 13579 -2038 13586
rect -2317 13574 -2309 13578
rect -2000 13576 -1992 13596
rect -1844 13588 -1794 13596
rect -1671 13590 -1663 13596
rect -1852 13579 -1804 13586
rect -1655 13578 -1647 13590
rect -2025 13575 -1991 13576
rect -2025 13574 -1975 13575
rect -1844 13574 -1804 13577
rect -1663 13574 -1655 13578
rect -1642 13574 -1637 13596
rect -1619 13574 -1614 13596
rect -1530 13574 -1526 13596
rect -1506 13574 -1502 13596
rect -1482 13574 -1478 13596
rect -1458 13574 -1454 13596
rect -1451 13595 -1437 13596
rect -1434 13574 -1427 13619
rect -1410 13574 -1406 13668
rect -1386 13574 -1382 13668
rect -1362 13574 -1358 13668
rect -1338 13574 -1334 13668
rect -1314 13574 -1310 13668
rect -1290 13574 -1286 13668
rect -1266 13574 -1262 13668
rect -1242 13574 -1238 13668
rect -1218 13574 -1214 13668
rect -1194 13574 -1190 13668
rect -1170 13574 -1166 13668
rect -1146 13574 -1142 13668
rect -1122 13574 -1118 13668
rect -1098 13574 -1094 13668
rect -1074 13574 -1070 13668
rect -1050 13574 -1046 13668
rect -1026 13574 -1022 13668
rect -1002 13574 -998 13668
rect -978 13574 -974 13668
rect -965 13637 -960 13647
rect -954 13637 -950 13668
rect -955 13623 -950 13637
rect -965 13622 -931 13623
rect -930 13622 -926 13668
rect -906 13622 -902 13668
rect -882 13622 -878 13668
rect -858 13622 -854 13668
rect -834 13622 -830 13668
rect -810 13622 -806 13668
rect -786 13622 -782 13668
rect -762 13622 -758 13668
rect -738 13622 -734 13668
rect -714 13622 -710 13668
rect -690 13622 -686 13668
rect -666 13622 -662 13668
rect -642 13622 -638 13668
rect -629 13661 -624 13668
rect -618 13661 -614 13668
rect -619 13647 -614 13661
rect -629 13637 -624 13647
rect -619 13623 -614 13637
rect -618 13622 -614 13623
rect -594 13622 -590 13716
rect -570 13622 -566 13716
rect -546 13622 -542 13716
rect -522 13622 -518 13716
rect -498 13622 -494 13716
rect -474 13622 -470 13716
rect -450 13691 -446 13716
rect -450 13646 -443 13691
rect -426 13646 -422 13716
rect -402 13646 -398 13716
rect -378 13646 -374 13716
rect -354 13646 -350 13716
rect -330 13646 -326 13716
rect -306 13646 -302 13716
rect -282 13646 -278 13716
rect -258 13646 -254 13716
rect -234 13646 -230 13716
rect -210 13646 -206 13716
rect -186 13646 -182 13716
rect -162 13646 -158 13716
rect -138 13646 -134 13716
rect -114 13646 -110 13716
rect -90 13646 -86 13716
rect -66 13646 -62 13716
rect -42 13715 -38 13716
rect -42 13667 -35 13715
rect -42 13646 -38 13667
rect -18 13646 -14 13716
rect 6 13646 10 13716
rect 30 13646 34 13716
rect 54 13646 58 13716
rect 78 13646 82 13716
rect 102 13646 106 13716
rect 109 13715 123 13716
rect 126 13691 133 13739
rect 126 13646 130 13691
rect 150 13646 154 13740
rect 174 13646 178 13740
rect 198 13646 202 13740
rect 222 13646 226 13740
rect 246 13646 250 13740
rect 270 13646 274 13740
rect 294 13646 298 13740
rect 318 13646 322 13740
rect 342 13646 346 13740
rect 366 13646 370 13740
rect 390 13646 394 13740
rect 414 13646 418 13740
rect 438 13646 442 13740
rect 462 13646 466 13740
rect 486 13646 490 13740
rect 510 13646 514 13740
rect 534 13646 538 13740
rect 558 13646 562 13740
rect 582 13646 586 13740
rect 589 13739 603 13740
rect 606 13718 613 13763
rect 630 13718 634 13764
rect 654 13718 658 13764
rect 678 13718 682 13764
rect 702 13718 706 13764
rect 726 13718 730 13764
rect 750 13718 754 13764
rect 774 13718 778 13764
rect 798 13718 802 13764
rect 822 13718 826 13764
rect 846 13718 850 13764
rect 870 13718 874 13764
rect 894 13718 898 13764
rect 918 13718 922 13764
rect 942 13718 946 13764
rect 966 13718 970 13764
rect 990 13718 994 13764
rect 1014 13718 1018 13764
rect 1038 13718 1042 13764
rect 1062 13718 1066 13764
rect 1086 13718 1090 13764
rect 1110 13718 1114 13764
rect 1134 13718 1138 13764
rect 1158 13718 1162 13764
rect 1182 13718 1186 13764
rect 1206 13718 1210 13764
rect 1230 13718 1234 13764
rect 1254 13718 1258 13764
rect 1278 13718 1282 13764
rect 1302 13718 1306 13764
rect 1326 13718 1330 13764
rect 1350 13718 1354 13764
rect 1374 13718 1378 13764
rect 1398 13718 1402 13764
rect 1422 13718 1426 13764
rect 1446 13718 1450 13764
rect 1470 13718 1474 13764
rect 1494 13718 1498 13764
rect 1518 13718 1522 13764
rect 1542 13718 1546 13764
rect 1566 13718 1570 13764
rect 1590 13718 1594 13764
rect 1614 13718 1618 13764
rect 1638 13718 1642 13764
rect 1662 13718 1666 13764
rect 1686 13718 1690 13764
rect 1710 13718 1714 13764
rect 1734 13718 1738 13764
rect 1758 13718 1762 13764
rect 1782 13718 1786 13764
rect 1806 13718 1810 13764
rect 1830 13718 1834 13764
rect 1854 13718 1858 13764
rect 1878 13718 1882 13764
rect 1902 13718 1906 13764
rect 1926 13718 1930 13764
rect 1950 13718 1954 13764
rect 1974 13718 1978 13764
rect 1998 13718 2002 13764
rect 2022 13718 2026 13764
rect 2046 13718 2050 13764
rect 2070 13718 2074 13764
rect 2094 13718 2098 13764
rect 2118 13718 2122 13764
rect 2142 13718 2146 13764
rect 2166 13718 2170 13764
rect 2190 13718 2194 13764
rect 2214 13718 2218 13764
rect 2238 13718 2242 13764
rect 2262 13718 2266 13764
rect 2286 13718 2290 13764
rect 2310 13718 2314 13764
rect 2334 13718 2338 13764
rect 2358 13718 2362 13764
rect 2382 13718 2386 13764
rect 2406 13718 2410 13764
rect 2430 13718 2434 13764
rect 2454 13718 2458 13764
rect 2478 13718 2482 13764
rect 2502 13718 2506 13764
rect 2526 13718 2530 13764
rect 2550 13718 2554 13764
rect 2574 13718 2578 13764
rect 2598 13718 2602 13764
rect 2622 13718 2626 13764
rect 2646 13718 2650 13764
rect 2670 13718 2674 13764
rect 2694 13718 2698 13764
rect 2718 13718 2722 13764
rect 2742 13718 2746 13764
rect 2766 13718 2770 13764
rect 2790 13718 2794 13764
rect 2814 13718 2818 13764
rect 2838 13718 2842 13764
rect 2862 13718 2866 13764
rect 2886 13718 2890 13764
rect 2910 13718 2914 13764
rect 2934 13718 2938 13764
rect 2958 13718 2962 13764
rect 2982 13718 2986 13764
rect 3006 13718 3010 13764
rect 3030 13718 3034 13764
rect 3054 13718 3058 13764
rect 3078 13718 3082 13764
rect 3102 13718 3106 13764
rect 3126 13718 3130 13764
rect 3150 13718 3154 13764
rect 3174 13718 3178 13764
rect 3198 13718 3202 13764
rect 3222 13718 3226 13764
rect 3246 13718 3250 13764
rect 3270 13718 3274 13764
rect 3294 13718 3298 13764
rect 3318 13718 3322 13764
rect 3342 13718 3346 13764
rect 3366 13718 3370 13764
rect 3390 13718 3394 13764
rect 3414 13718 3418 13764
rect 3438 13718 3442 13764
rect 3462 13718 3466 13764
rect 3486 13718 3490 13764
rect 3510 13718 3514 13764
rect 3534 13718 3538 13764
rect 3558 13718 3562 13764
rect 3582 13718 3586 13764
rect 3606 13718 3610 13764
rect 3619 13733 3624 13743
rect 3630 13733 3634 13764
rect 3643 13757 3648 13764
rect 3654 13757 3658 13764
rect 3653 13743 3658 13757
rect 3629 13719 3634 13733
rect 3619 13718 3653 13719
rect 589 13716 3653 13718
rect 589 13715 603 13716
rect 606 13715 613 13716
rect 606 13646 610 13715
rect 630 13646 634 13716
rect 654 13646 658 13716
rect 678 13646 682 13716
rect 702 13646 706 13716
rect 726 13646 730 13716
rect 750 13646 754 13716
rect 774 13646 778 13716
rect 798 13646 802 13716
rect 822 13646 826 13716
rect 846 13646 850 13716
rect 870 13646 874 13716
rect 894 13646 898 13716
rect 918 13646 922 13716
rect 942 13646 946 13716
rect 966 13646 970 13716
rect 990 13646 994 13716
rect 1014 13646 1018 13716
rect 1038 13646 1042 13716
rect 1062 13646 1066 13716
rect 1086 13646 1090 13716
rect 1110 13646 1114 13716
rect 1134 13646 1138 13716
rect 1158 13646 1162 13716
rect 1182 13646 1186 13716
rect 1206 13646 1210 13716
rect 1230 13646 1234 13716
rect 1254 13646 1258 13716
rect 1278 13646 1282 13716
rect 1302 13646 1306 13716
rect 1326 13646 1330 13716
rect 1350 13646 1354 13716
rect 1374 13646 1378 13716
rect 1398 13646 1402 13716
rect 1422 13646 1426 13716
rect 1446 13646 1450 13716
rect 1470 13646 1474 13716
rect 1494 13646 1498 13716
rect 1518 13646 1522 13716
rect 1542 13646 1546 13716
rect 1566 13646 1570 13716
rect 1590 13646 1594 13716
rect 1614 13646 1618 13716
rect 1638 13646 1642 13716
rect 1662 13646 1666 13716
rect 1686 13646 1690 13716
rect 1710 13646 1714 13716
rect 1734 13646 1738 13716
rect 1758 13646 1762 13716
rect 1782 13646 1786 13716
rect 1806 13646 1810 13716
rect 1830 13646 1834 13716
rect 1854 13646 1858 13716
rect 1878 13646 1882 13716
rect 1902 13646 1906 13716
rect 1926 13646 1930 13716
rect 1950 13646 1954 13716
rect 1974 13646 1978 13716
rect 1998 13646 2002 13716
rect 2022 13646 2026 13716
rect 2046 13646 2050 13716
rect 2070 13646 2074 13716
rect 2094 13646 2098 13716
rect 2118 13646 2122 13716
rect 2142 13646 2146 13716
rect 2166 13646 2170 13716
rect 2190 13646 2194 13716
rect 2214 13646 2218 13716
rect 2238 13646 2242 13716
rect 2262 13646 2266 13716
rect 2286 13646 2290 13716
rect 2310 13646 2314 13716
rect 2334 13646 2338 13716
rect 2358 13646 2362 13716
rect 2382 13646 2386 13716
rect 2406 13646 2410 13716
rect 2430 13646 2434 13716
rect 2454 13646 2458 13716
rect 2478 13646 2482 13716
rect 2502 13646 2506 13716
rect 2526 13646 2530 13716
rect 2550 13646 2554 13716
rect 2574 13646 2578 13716
rect 2598 13646 2602 13716
rect 2622 13646 2626 13716
rect 2646 13646 2650 13716
rect 2670 13646 2674 13716
rect 2694 13646 2698 13716
rect 2718 13646 2722 13716
rect 2742 13646 2746 13716
rect 2766 13646 2770 13716
rect 2790 13646 2794 13716
rect 2814 13646 2818 13716
rect 2838 13646 2842 13716
rect 2862 13646 2866 13716
rect 2886 13646 2890 13716
rect 2910 13646 2914 13716
rect 2934 13646 2938 13716
rect 2958 13646 2962 13716
rect 2982 13646 2986 13716
rect 3006 13646 3010 13716
rect 3030 13646 3034 13716
rect 3054 13646 3058 13716
rect 3078 13646 3082 13716
rect 3102 13646 3106 13716
rect 3126 13646 3130 13716
rect 3150 13646 3154 13716
rect 3174 13646 3178 13716
rect 3198 13646 3202 13716
rect 3222 13646 3226 13716
rect 3246 13646 3250 13716
rect 3270 13646 3274 13716
rect 3294 13646 3298 13716
rect 3318 13646 3322 13716
rect 3342 13646 3346 13716
rect 3366 13646 3370 13716
rect 3390 13646 3394 13716
rect 3414 13646 3418 13716
rect 3438 13646 3442 13716
rect 3462 13646 3466 13716
rect 3486 13646 3490 13716
rect 3510 13646 3514 13716
rect 3534 13646 3538 13716
rect 3558 13646 3562 13716
rect 3582 13646 3586 13716
rect 3606 13646 3610 13716
rect 3619 13709 3624 13716
rect 3629 13695 3634 13709
rect 3630 13647 3634 13695
rect 3619 13646 3651 13647
rect -467 13644 3651 13646
rect -467 13643 -453 13644
rect -450 13643 -443 13644
rect -450 13622 -446 13643
rect -426 13622 -422 13644
rect -402 13622 -398 13644
rect -378 13622 -374 13644
rect -354 13622 -350 13644
rect -330 13622 -326 13644
rect -306 13622 -302 13644
rect -282 13622 -278 13644
rect -258 13622 -254 13644
rect -234 13622 -230 13644
rect -210 13622 -206 13644
rect -186 13622 -182 13644
rect -162 13622 -158 13644
rect -138 13622 -134 13644
rect -114 13622 -110 13644
rect -90 13622 -86 13644
rect -66 13622 -62 13644
rect -42 13622 -38 13644
rect -18 13622 -14 13644
rect 6 13622 10 13644
rect 30 13622 34 13644
rect 54 13622 58 13644
rect 78 13622 82 13644
rect 102 13622 106 13644
rect 126 13622 130 13644
rect 150 13622 154 13644
rect 174 13622 178 13644
rect 198 13622 202 13644
rect 222 13622 226 13644
rect 246 13622 250 13644
rect 270 13622 274 13644
rect 294 13622 298 13644
rect 318 13622 322 13644
rect 342 13622 346 13644
rect 366 13622 370 13644
rect 390 13622 394 13644
rect 414 13622 418 13644
rect 438 13622 442 13644
rect 462 13622 466 13644
rect 486 13622 490 13644
rect 510 13622 514 13644
rect 534 13622 538 13644
rect 558 13622 562 13644
rect 582 13622 586 13644
rect 606 13622 610 13644
rect 630 13622 634 13644
rect 654 13622 658 13644
rect 678 13622 682 13644
rect 702 13622 706 13644
rect 726 13622 730 13644
rect 750 13622 754 13644
rect 774 13622 778 13644
rect 798 13622 802 13644
rect 822 13622 826 13644
rect 846 13622 850 13644
rect 870 13622 874 13644
rect 894 13622 898 13644
rect 918 13622 922 13644
rect 942 13622 946 13644
rect 966 13622 970 13644
rect 990 13622 994 13644
rect 1014 13622 1018 13644
rect 1038 13622 1042 13644
rect 1062 13622 1066 13644
rect 1086 13622 1090 13644
rect 1110 13622 1114 13644
rect 1134 13622 1138 13644
rect 1158 13622 1162 13644
rect 1182 13622 1186 13644
rect 1206 13622 1210 13644
rect 1230 13622 1234 13644
rect 1254 13622 1258 13644
rect 1278 13622 1282 13644
rect 1302 13622 1306 13644
rect 1326 13622 1330 13644
rect 1350 13622 1354 13644
rect 1374 13622 1378 13644
rect 1398 13622 1402 13644
rect 1422 13622 1426 13644
rect 1446 13622 1450 13644
rect 1470 13622 1474 13644
rect 1494 13622 1498 13644
rect 1518 13622 1522 13644
rect 1542 13622 1546 13644
rect 1566 13622 1570 13644
rect 1590 13622 1594 13644
rect 1614 13622 1618 13644
rect 1638 13622 1642 13644
rect 1662 13622 1666 13644
rect 1686 13622 1690 13644
rect 1710 13622 1714 13644
rect 1734 13622 1738 13644
rect 1758 13622 1762 13644
rect 1782 13622 1786 13644
rect 1806 13622 1810 13644
rect 1830 13622 1834 13644
rect 1854 13622 1858 13644
rect 1878 13622 1882 13644
rect 1902 13622 1906 13644
rect 1926 13622 1930 13644
rect 1950 13622 1954 13644
rect 1974 13622 1978 13644
rect 1998 13622 2002 13644
rect 2022 13622 2026 13644
rect 2046 13622 2050 13644
rect 2070 13622 2074 13644
rect 2094 13622 2098 13644
rect 2118 13622 2122 13644
rect 2142 13622 2146 13644
rect 2166 13622 2170 13644
rect 2190 13622 2194 13644
rect 2214 13622 2218 13644
rect 2238 13622 2242 13644
rect 2262 13622 2266 13644
rect 2286 13622 2290 13644
rect 2310 13622 2314 13644
rect 2334 13622 2338 13644
rect 2358 13622 2362 13644
rect 2382 13622 2386 13644
rect 2406 13622 2410 13644
rect 2430 13622 2434 13644
rect 2454 13622 2458 13644
rect 2478 13622 2482 13644
rect 2502 13622 2506 13644
rect 2526 13622 2530 13644
rect 2550 13622 2554 13644
rect 2574 13622 2578 13644
rect 2598 13622 2602 13644
rect 2622 13622 2626 13644
rect 2646 13622 2650 13644
rect 2670 13622 2674 13644
rect 2694 13622 2698 13644
rect 2718 13622 2722 13644
rect 2742 13622 2746 13644
rect 2766 13622 2770 13644
rect 2790 13622 2794 13644
rect 2814 13622 2818 13644
rect 2838 13622 2842 13644
rect 2862 13622 2866 13644
rect 2886 13622 2890 13644
rect 2910 13622 2914 13644
rect 2934 13622 2938 13644
rect 2958 13622 2962 13644
rect 2982 13622 2986 13644
rect 3006 13622 3010 13644
rect 3030 13622 3034 13644
rect 3054 13622 3058 13644
rect 3078 13622 3082 13644
rect 3102 13622 3106 13644
rect 3126 13622 3130 13644
rect 3150 13622 3154 13644
rect 3174 13622 3178 13644
rect 3198 13622 3202 13644
rect 3222 13622 3226 13644
rect 3246 13622 3250 13644
rect 3270 13622 3274 13644
rect 3294 13622 3298 13644
rect 3318 13622 3322 13644
rect 3342 13622 3346 13644
rect 3366 13622 3370 13644
rect 3390 13622 3394 13644
rect 3414 13622 3418 13644
rect 3438 13622 3442 13644
rect 3462 13622 3466 13644
rect 3486 13622 3490 13644
rect 3510 13622 3514 13644
rect 3534 13622 3538 13644
rect 3558 13622 3562 13644
rect 3582 13622 3586 13644
rect 3606 13623 3610 13644
rect 3619 13637 3624 13644
rect 3630 13637 3634 13644
rect 3637 13643 3651 13644
rect 3629 13623 3634 13637
rect 3643 13633 3651 13637
rect 3637 13623 3643 13633
rect 3595 13622 3629 13623
rect -965 13620 3629 13622
rect -965 13613 -960 13620
rect -955 13599 -950 13613
rect -954 13574 -950 13599
rect -930 13574 -926 13620
rect -906 13574 -902 13620
rect -882 13574 -878 13620
rect -858 13574 -854 13620
rect -834 13574 -830 13620
rect -810 13574 -806 13620
rect -786 13574 -782 13620
rect -762 13574 -758 13620
rect -738 13574 -734 13620
rect -714 13574 -710 13620
rect -690 13574 -686 13620
rect -666 13574 -662 13620
rect -642 13574 -638 13620
rect -618 13574 -614 13620
rect -594 13595 -590 13620
rect -2393 13572 -597 13574
rect -2371 13550 -2366 13572
rect -2348 13550 -2343 13572
rect -2325 13562 -2317 13572
rect -2060 13562 -2020 13569
rect -2004 13564 -2001 13569
rect -2015 13562 -2001 13564
rect -2000 13562 -1992 13572
rect -1972 13570 -1958 13572
rect -1844 13571 -1804 13572
rect -1862 13569 -1796 13570
rect -1985 13567 -1796 13569
rect -1985 13562 -1852 13567
rect -2325 13550 -2320 13562
rect -2309 13550 -2301 13562
rect -2068 13552 -2060 13559
rect -2015 13552 -1990 13562
rect -1844 13561 -1796 13567
rect -1671 13562 -1663 13572
rect -1852 13552 -1804 13559
rect -2020 13550 -2004 13552
rect -2000 13550 -1992 13552
rect -1976 13550 -1940 13551
rect -1655 13550 -1647 13562
rect -1642 13550 -1637 13572
rect -1619 13550 -1614 13572
rect -1530 13550 -1526 13572
rect -1506 13550 -1502 13572
rect -1482 13550 -1478 13572
rect -1458 13550 -1454 13572
rect -1451 13571 -1437 13572
rect -1434 13571 -1427 13572
rect -1434 13550 -1430 13571
rect -1410 13550 -1406 13572
rect -1386 13550 -1382 13572
rect -1362 13550 -1358 13572
rect -1338 13550 -1334 13572
rect -1314 13550 -1310 13572
rect -1290 13550 -1286 13572
rect -1266 13550 -1262 13572
rect -1242 13550 -1238 13572
rect -1218 13550 -1214 13572
rect -1194 13550 -1190 13572
rect -1170 13550 -1166 13572
rect -1146 13550 -1142 13572
rect -1122 13550 -1118 13572
rect -1098 13550 -1094 13572
rect -1074 13550 -1070 13572
rect -1050 13550 -1046 13572
rect -1026 13550 -1022 13572
rect -1002 13550 -998 13572
rect -978 13550 -974 13572
rect -954 13550 -950 13572
rect -930 13571 -926 13572
rect -2393 13548 -933 13550
rect -2371 13478 -2366 13548
rect -2348 13478 -2343 13548
rect -2325 13546 -2320 13548
rect -2317 13546 -2309 13548
rect -2325 13534 -2317 13546
rect -2060 13535 -2030 13542
rect -2325 13514 -2320 13534
rect -2325 13506 -2317 13514
rect -2060 13508 -2030 13511
rect -2325 13486 -2320 13506
rect -2317 13498 -2309 13506
rect -2060 13495 -2038 13506
rect -2033 13499 -2030 13508
rect -2028 13504 -2027 13508
rect -2068 13490 -2038 13493
rect -2325 13478 -2317 13486
rect -2000 13478 -1992 13548
rect -1844 13544 -1804 13548
rect -1663 13546 -1655 13548
rect -1844 13534 -1794 13543
rect -1671 13534 -1663 13546
rect -1912 13523 -1884 13525
rect -1852 13517 -1804 13521
rect -1844 13508 -1796 13511
rect -1671 13506 -1663 13514
rect -1844 13495 -1804 13506
rect -1663 13498 -1655 13506
rect -1852 13490 -1680 13494
rect -1926 13478 -1892 13481
rect -1671 13478 -1663 13486
rect -1642 13478 -1637 13548
rect -1619 13478 -1614 13548
rect -1530 13478 -1526 13548
rect -1506 13478 -1502 13548
rect -1482 13478 -1478 13548
rect -1458 13478 -1454 13548
rect -1434 13478 -1430 13548
rect -1410 13478 -1406 13548
rect -1386 13478 -1382 13548
rect -1362 13478 -1358 13548
rect -1338 13478 -1334 13548
rect -1314 13478 -1310 13548
rect -1290 13478 -1286 13548
rect -1266 13478 -1262 13548
rect -1242 13478 -1238 13548
rect -1218 13478 -1214 13548
rect -1194 13478 -1190 13548
rect -1170 13478 -1166 13548
rect -1146 13478 -1142 13548
rect -1122 13478 -1118 13548
rect -1098 13478 -1094 13548
rect -1074 13478 -1070 13548
rect -1050 13478 -1046 13548
rect -1026 13478 -1022 13548
rect -1002 13478 -998 13548
rect -978 13478 -974 13548
rect -954 13478 -950 13548
rect -947 13547 -933 13548
rect -930 13526 -923 13571
rect -906 13526 -902 13572
rect -882 13526 -878 13572
rect -858 13526 -854 13572
rect -834 13526 -830 13572
rect -810 13526 -806 13572
rect -786 13526 -782 13572
rect -762 13526 -758 13572
rect -738 13526 -734 13572
rect -714 13526 -710 13572
rect -690 13526 -686 13572
rect -666 13526 -662 13572
rect -642 13526 -638 13572
rect -618 13526 -614 13572
rect -611 13571 -597 13572
rect -594 13550 -587 13595
rect -570 13550 -566 13620
rect -546 13550 -542 13620
rect -522 13550 -518 13620
rect -498 13550 -494 13620
rect -474 13550 -470 13620
rect -450 13550 -446 13620
rect -426 13550 -422 13620
rect -402 13550 -398 13620
rect -378 13550 -374 13620
rect -354 13550 -350 13620
rect -330 13550 -326 13620
rect -306 13550 -302 13620
rect -282 13550 -278 13620
rect -258 13550 -254 13620
rect -234 13550 -230 13620
rect -210 13550 -206 13620
rect -186 13550 -182 13620
rect -162 13550 -158 13620
rect -138 13550 -134 13620
rect -114 13550 -110 13620
rect -90 13550 -86 13620
rect -66 13550 -62 13620
rect -42 13550 -38 13620
rect -18 13550 -14 13620
rect 6 13550 10 13620
rect 30 13550 34 13620
rect 54 13550 58 13620
rect 78 13550 82 13620
rect 102 13550 106 13620
rect 126 13550 130 13620
rect 150 13550 154 13620
rect 174 13550 178 13620
rect 198 13550 202 13620
rect 222 13550 226 13620
rect 246 13550 250 13620
rect 270 13550 274 13620
rect 294 13550 298 13620
rect 318 13550 322 13620
rect 331 13565 336 13575
rect 342 13565 346 13620
rect 341 13551 346 13565
rect 366 13550 370 13620
rect 390 13550 394 13620
rect 414 13550 418 13620
rect 438 13550 442 13620
rect 462 13550 466 13620
rect 486 13550 490 13620
rect 510 13550 514 13620
rect 534 13550 538 13620
rect 558 13550 562 13620
rect 582 13550 586 13620
rect 606 13550 610 13620
rect 630 13550 634 13620
rect 654 13550 658 13620
rect 678 13550 682 13620
rect 702 13550 706 13620
rect 726 13550 730 13620
rect 750 13550 754 13620
rect 774 13550 778 13620
rect 798 13550 802 13620
rect 822 13550 826 13620
rect 846 13550 850 13620
rect 870 13550 874 13620
rect 894 13550 898 13620
rect 918 13550 922 13620
rect 942 13550 946 13620
rect 966 13550 970 13620
rect 990 13550 994 13620
rect 1014 13550 1018 13620
rect 1038 13550 1042 13620
rect 1062 13550 1066 13620
rect 1086 13550 1090 13620
rect 1110 13550 1114 13620
rect 1134 13550 1138 13620
rect 1158 13551 1162 13620
rect 1147 13550 1181 13551
rect -611 13548 1181 13550
rect -611 13547 -597 13548
rect -594 13547 -587 13548
rect -594 13526 -590 13547
rect -570 13526 -566 13548
rect -546 13526 -542 13548
rect -522 13526 -518 13548
rect -498 13526 -494 13548
rect -474 13526 -470 13548
rect -450 13526 -446 13548
rect -426 13526 -422 13548
rect -402 13526 -398 13548
rect -378 13526 -374 13548
rect -354 13526 -350 13548
rect -330 13526 -326 13548
rect -306 13526 -302 13548
rect -282 13526 -278 13548
rect -258 13526 -254 13548
rect -234 13526 -230 13548
rect -210 13526 -206 13548
rect -186 13526 -182 13548
rect -162 13526 -158 13548
rect -138 13526 -134 13548
rect -114 13526 -110 13548
rect -90 13526 -86 13548
rect -66 13526 -62 13548
rect -42 13526 -38 13548
rect -18 13526 -14 13548
rect 6 13526 10 13548
rect 30 13526 34 13548
rect 54 13526 58 13548
rect 78 13526 82 13548
rect 102 13526 106 13548
rect 126 13526 130 13548
rect 150 13526 154 13548
rect 174 13526 178 13548
rect 198 13526 202 13548
rect 222 13527 226 13548
rect 211 13526 245 13527
rect -947 13524 245 13526
rect -947 13523 -933 13524
rect -930 13523 -923 13524
rect -930 13478 -926 13523
rect -906 13478 -902 13524
rect -882 13478 -878 13524
rect -858 13478 -854 13524
rect -834 13478 -830 13524
rect -810 13478 -806 13524
rect -786 13478 -782 13524
rect -762 13478 -758 13524
rect -738 13478 -734 13524
rect -714 13478 -710 13524
rect -690 13478 -686 13524
rect -666 13478 -662 13524
rect -642 13478 -638 13524
rect -618 13478 -614 13524
rect -594 13478 -590 13524
rect -570 13478 -566 13524
rect -546 13478 -542 13524
rect -522 13478 -518 13524
rect -498 13478 -494 13524
rect -474 13478 -470 13524
rect -450 13478 -446 13524
rect -426 13478 -422 13524
rect -402 13478 -398 13524
rect -378 13478 -374 13524
rect -354 13478 -350 13524
rect -330 13478 -326 13524
rect -306 13478 -302 13524
rect -282 13478 -278 13524
rect -258 13478 -254 13524
rect -234 13478 -230 13524
rect -210 13478 -206 13524
rect -186 13478 -182 13524
rect -162 13478 -158 13524
rect -138 13478 -134 13524
rect -114 13478 -110 13524
rect -90 13478 -86 13524
rect -66 13478 -62 13524
rect -42 13478 -38 13524
rect -18 13478 -14 13524
rect 6 13478 10 13524
rect 30 13478 34 13524
rect 54 13478 58 13524
rect 78 13478 82 13524
rect 102 13478 106 13524
rect 126 13478 130 13524
rect 150 13478 154 13524
rect 174 13478 178 13524
rect 198 13478 202 13524
rect 211 13517 216 13524
rect 222 13517 226 13524
rect 221 13503 226 13517
rect 211 13502 245 13503
rect 246 13502 250 13548
rect 270 13502 274 13548
rect 294 13502 298 13548
rect 318 13502 322 13548
rect 331 13526 365 13527
rect 366 13526 370 13548
rect 390 13526 394 13548
rect 414 13526 418 13548
rect 438 13526 442 13548
rect 462 13526 466 13548
rect 486 13526 490 13548
rect 510 13526 514 13548
rect 534 13526 538 13548
rect 558 13526 562 13548
rect 582 13526 586 13548
rect 606 13526 610 13548
rect 630 13526 634 13548
rect 654 13526 658 13548
rect 678 13526 682 13548
rect 702 13526 706 13548
rect 726 13526 730 13548
rect 750 13526 754 13548
rect 774 13526 778 13548
rect 798 13526 802 13548
rect 822 13526 826 13548
rect 846 13526 850 13548
rect 870 13526 874 13548
rect 894 13526 898 13548
rect 918 13526 922 13548
rect 942 13526 946 13548
rect 966 13526 970 13548
rect 990 13526 994 13548
rect 1014 13526 1018 13548
rect 1038 13526 1042 13548
rect 1062 13526 1066 13548
rect 1086 13526 1090 13548
rect 1110 13526 1114 13548
rect 1134 13526 1138 13548
rect 1147 13541 1152 13548
rect 1158 13541 1162 13548
rect 1157 13527 1162 13541
rect 1182 13526 1186 13620
rect 1206 13526 1210 13620
rect 1230 13526 1234 13620
rect 1254 13526 1258 13620
rect 1278 13526 1282 13620
rect 1302 13526 1306 13620
rect 1326 13526 1330 13620
rect 1350 13526 1354 13620
rect 1374 13526 1378 13620
rect 1398 13526 1402 13620
rect 1422 13526 1426 13620
rect 1446 13526 1450 13620
rect 1470 13526 1474 13620
rect 1494 13526 1498 13620
rect 1518 13526 1522 13620
rect 1542 13526 1546 13620
rect 1566 13526 1570 13620
rect 1590 13526 1594 13620
rect 1614 13526 1618 13620
rect 1638 13526 1642 13620
rect 1662 13526 1666 13620
rect 1686 13526 1690 13620
rect 1710 13526 1714 13620
rect 1734 13526 1738 13620
rect 1758 13526 1762 13620
rect 1782 13526 1786 13620
rect 1806 13526 1810 13620
rect 1830 13526 1834 13620
rect 1854 13526 1858 13620
rect 1878 13526 1882 13620
rect 1902 13526 1906 13620
rect 1926 13526 1930 13620
rect 1950 13526 1954 13620
rect 1974 13526 1978 13620
rect 1998 13526 2002 13620
rect 2022 13526 2026 13620
rect 2046 13526 2050 13620
rect 2070 13526 2074 13620
rect 2094 13526 2098 13620
rect 2118 13526 2122 13620
rect 2142 13526 2146 13620
rect 2166 13526 2170 13620
rect 2190 13526 2194 13620
rect 2214 13526 2218 13620
rect 2238 13526 2242 13620
rect 2262 13526 2266 13620
rect 2286 13526 2290 13620
rect 2310 13526 2314 13620
rect 2334 13526 2338 13620
rect 2358 13526 2362 13620
rect 2382 13526 2386 13620
rect 2406 13526 2410 13620
rect 2430 13526 2434 13620
rect 2454 13526 2458 13620
rect 2478 13526 2482 13620
rect 2502 13526 2506 13620
rect 2526 13526 2530 13620
rect 2550 13526 2554 13620
rect 2574 13526 2578 13620
rect 2598 13526 2602 13620
rect 2622 13526 2626 13620
rect 2646 13526 2650 13620
rect 2670 13526 2674 13620
rect 2694 13526 2698 13620
rect 2718 13526 2722 13620
rect 2742 13526 2746 13620
rect 2766 13526 2770 13620
rect 2790 13526 2794 13620
rect 2814 13526 2818 13620
rect 2838 13526 2842 13620
rect 2862 13526 2866 13620
rect 2886 13526 2890 13620
rect 2910 13526 2914 13620
rect 2934 13526 2938 13620
rect 2958 13526 2962 13620
rect 2982 13526 2986 13620
rect 3006 13526 3010 13620
rect 3030 13526 3034 13620
rect 3054 13526 3058 13620
rect 3078 13526 3082 13620
rect 3102 13526 3106 13620
rect 3126 13526 3130 13620
rect 3150 13526 3154 13620
rect 3174 13526 3178 13620
rect 3198 13526 3202 13620
rect 3222 13526 3226 13620
rect 3246 13526 3250 13620
rect 3270 13526 3274 13620
rect 3294 13526 3298 13620
rect 3318 13526 3322 13620
rect 3342 13526 3346 13620
rect 3366 13526 3370 13620
rect 3390 13526 3394 13620
rect 3414 13526 3418 13620
rect 3438 13526 3442 13620
rect 3462 13526 3466 13620
rect 3486 13526 3490 13620
rect 3510 13526 3514 13620
rect 3534 13526 3538 13620
rect 3558 13526 3562 13620
rect 3582 13526 3586 13620
rect 3595 13613 3600 13620
rect 3606 13613 3610 13620
rect 3605 13599 3610 13613
rect 3595 13589 3600 13599
rect 3605 13575 3610 13589
rect 3606 13527 3610 13575
rect 3595 13526 3627 13527
rect 331 13524 3627 13526
rect 331 13517 336 13524
rect 341 13503 346 13517
rect 342 13502 346 13503
rect 366 13502 370 13524
rect 390 13502 394 13524
rect 414 13502 418 13524
rect 438 13502 442 13524
rect 462 13502 466 13524
rect 486 13502 490 13524
rect 510 13502 514 13524
rect 534 13502 538 13524
rect 558 13502 562 13524
rect 582 13502 586 13524
rect 606 13502 610 13524
rect 630 13502 634 13524
rect 654 13502 658 13524
rect 678 13502 682 13524
rect 702 13502 706 13524
rect 726 13502 730 13524
rect 750 13502 754 13524
rect 774 13502 778 13524
rect 798 13502 802 13524
rect 822 13502 826 13524
rect 846 13502 850 13524
rect 870 13502 874 13524
rect 894 13502 898 13524
rect 918 13502 922 13524
rect 942 13502 946 13524
rect 966 13502 970 13524
rect 990 13502 994 13524
rect 1014 13502 1018 13524
rect 1038 13502 1042 13524
rect 1062 13502 1066 13524
rect 1086 13502 1090 13524
rect 1110 13502 1114 13524
rect 1134 13502 1138 13524
rect 1182 13502 1186 13524
rect 1206 13502 1210 13524
rect 1230 13502 1234 13524
rect 1254 13502 1258 13524
rect 1278 13502 1282 13524
rect 1302 13502 1306 13524
rect 1326 13502 1330 13524
rect 1350 13502 1354 13524
rect 1374 13502 1378 13524
rect 1398 13502 1402 13524
rect 1422 13502 1426 13524
rect 1446 13502 1450 13524
rect 1470 13502 1474 13524
rect 1494 13502 1498 13524
rect 1518 13502 1522 13524
rect 1542 13502 1546 13524
rect 1566 13502 1570 13524
rect 1590 13502 1594 13524
rect 1614 13502 1618 13524
rect 1638 13502 1642 13524
rect 1662 13502 1666 13524
rect 1686 13502 1690 13524
rect 1710 13502 1714 13524
rect 1734 13502 1738 13524
rect 1758 13502 1762 13524
rect 1782 13502 1786 13524
rect 1806 13502 1810 13524
rect 1830 13502 1834 13524
rect 1854 13502 1858 13524
rect 1878 13502 1882 13524
rect 1902 13502 1906 13524
rect 1926 13502 1930 13524
rect 1950 13502 1954 13524
rect 1974 13502 1978 13524
rect 1998 13502 2002 13524
rect 2022 13502 2026 13524
rect 2046 13502 2050 13524
rect 2070 13502 2074 13524
rect 2094 13502 2098 13524
rect 2118 13502 2122 13524
rect 2142 13502 2146 13524
rect 2166 13502 2170 13524
rect 2190 13502 2194 13524
rect 2214 13502 2218 13524
rect 2238 13502 2242 13524
rect 2262 13502 2266 13524
rect 2286 13502 2290 13524
rect 2310 13502 2314 13524
rect 2334 13502 2338 13524
rect 2358 13502 2362 13524
rect 2382 13502 2386 13524
rect 2406 13502 2410 13524
rect 2430 13502 2434 13524
rect 2454 13502 2458 13524
rect 2478 13502 2482 13524
rect 2502 13502 2506 13524
rect 2526 13502 2530 13524
rect 2550 13502 2554 13524
rect 2574 13502 2578 13524
rect 2598 13502 2602 13524
rect 2622 13502 2626 13524
rect 2646 13502 2650 13524
rect 2670 13502 2674 13524
rect 2694 13502 2698 13524
rect 2718 13502 2722 13524
rect 2742 13502 2746 13524
rect 2766 13502 2770 13524
rect 2790 13502 2794 13524
rect 2814 13502 2818 13524
rect 2838 13502 2842 13524
rect 2862 13502 2866 13524
rect 2886 13502 2890 13524
rect 2910 13502 2914 13524
rect 2934 13502 2938 13524
rect 2958 13502 2962 13524
rect 2982 13502 2986 13524
rect 3006 13502 3010 13524
rect 3030 13502 3034 13524
rect 3054 13502 3058 13524
rect 3078 13502 3082 13524
rect 3102 13502 3106 13524
rect 3126 13502 3130 13524
rect 3150 13502 3154 13524
rect 3174 13502 3178 13524
rect 3198 13502 3202 13524
rect 3222 13502 3226 13524
rect 3246 13502 3250 13524
rect 3270 13502 3274 13524
rect 3294 13502 3298 13524
rect 3318 13502 3322 13524
rect 3342 13502 3346 13524
rect 3366 13502 3370 13524
rect 3390 13502 3394 13524
rect 3414 13502 3418 13524
rect 3438 13502 3442 13524
rect 3462 13502 3466 13524
rect 3486 13502 3490 13524
rect 3510 13502 3514 13524
rect 3534 13502 3538 13524
rect 3558 13502 3562 13524
rect 3582 13503 3586 13524
rect 3595 13517 3600 13524
rect 3606 13517 3610 13524
rect 3613 13523 3627 13524
rect 3605 13503 3610 13517
rect 3619 13513 3627 13517
rect 3613 13503 3619 13513
rect 3571 13502 3605 13503
rect 211 13500 3605 13502
rect 211 13493 216 13500
rect 221 13479 226 13493
rect 222 13478 226 13479
rect 246 13478 250 13500
rect 270 13478 274 13500
rect 294 13478 298 13500
rect 318 13478 322 13500
rect 342 13478 346 13500
rect 366 13499 370 13500
rect -2393 13476 363 13478
rect -2371 13454 -2366 13476
rect -2348 13454 -2343 13476
rect -2325 13470 -2317 13476
rect -2325 13454 -2320 13470
rect -2309 13458 -2301 13470
rect -2068 13459 -2038 13466
rect -2317 13454 -2309 13458
rect -2000 13456 -1992 13476
rect -1844 13468 -1794 13476
rect -1671 13470 -1663 13476
rect -1852 13459 -1804 13466
rect -1655 13458 -1647 13470
rect -2025 13455 -1991 13456
rect -2025 13454 -1975 13455
rect -1844 13454 -1804 13457
rect -1663 13454 -1655 13458
rect -1642 13454 -1637 13476
rect -1619 13454 -1614 13476
rect -1530 13454 -1526 13476
rect -1506 13454 -1502 13476
rect -1482 13454 -1478 13476
rect -1458 13454 -1454 13476
rect -1434 13454 -1430 13476
rect -1410 13454 -1406 13476
rect -1386 13454 -1382 13476
rect -1362 13454 -1358 13476
rect -1338 13454 -1334 13476
rect -1314 13454 -1310 13476
rect -1290 13454 -1286 13476
rect -1266 13454 -1262 13476
rect -1242 13454 -1238 13476
rect -1218 13454 -1214 13476
rect -1194 13454 -1190 13476
rect -1170 13454 -1166 13476
rect -1146 13454 -1142 13476
rect -1122 13454 -1118 13476
rect -1098 13454 -1094 13476
rect -1074 13454 -1070 13476
rect -1050 13454 -1046 13476
rect -1026 13454 -1022 13476
rect -1002 13454 -998 13476
rect -978 13454 -974 13476
rect -954 13454 -950 13476
rect -930 13454 -926 13476
rect -906 13454 -902 13476
rect -882 13454 -878 13476
rect -858 13454 -854 13476
rect -834 13454 -830 13476
rect -810 13454 -806 13476
rect -786 13454 -782 13476
rect -762 13454 -758 13476
rect -738 13454 -734 13476
rect -714 13454 -710 13476
rect -690 13454 -686 13476
rect -666 13454 -662 13476
rect -642 13454 -638 13476
rect -618 13454 -614 13476
rect -594 13454 -590 13476
rect -570 13454 -566 13476
rect -546 13454 -542 13476
rect -522 13454 -518 13476
rect -498 13454 -494 13476
rect -474 13454 -470 13476
rect -450 13454 -446 13476
rect -426 13454 -422 13476
rect -402 13454 -398 13476
rect -378 13454 -374 13476
rect -354 13454 -350 13476
rect -330 13454 -326 13476
rect -306 13454 -302 13476
rect -282 13454 -278 13476
rect -258 13454 -254 13476
rect -234 13454 -230 13476
rect -210 13454 -206 13476
rect -186 13454 -182 13476
rect -162 13454 -158 13476
rect -138 13454 -134 13476
rect -114 13454 -110 13476
rect -90 13454 -86 13476
rect -66 13454 -62 13476
rect -42 13454 -38 13476
rect -18 13454 -14 13476
rect 6 13454 10 13476
rect 30 13454 34 13476
rect 54 13454 58 13476
rect 78 13454 82 13476
rect 102 13454 106 13476
rect 126 13454 130 13476
rect 150 13454 154 13476
rect 174 13454 178 13476
rect 198 13454 202 13476
rect 222 13454 226 13476
rect 246 13454 250 13476
rect 270 13454 274 13476
rect 294 13454 298 13476
rect 318 13454 322 13476
rect 342 13454 346 13476
rect 349 13475 363 13476
rect 366 13475 373 13499
rect 390 13454 394 13500
rect 414 13454 418 13500
rect 438 13454 442 13500
rect 462 13454 466 13500
rect 486 13454 490 13500
rect 510 13454 514 13500
rect 534 13454 538 13500
rect 558 13454 562 13500
rect 582 13454 586 13500
rect 606 13454 610 13500
rect 630 13454 634 13500
rect 654 13455 658 13500
rect 643 13454 677 13455
rect -2393 13452 677 13454
rect -2371 13430 -2366 13452
rect -2348 13430 -2343 13452
rect -2325 13442 -2317 13452
rect -2060 13442 -2020 13449
rect -2004 13444 -2001 13449
rect -2015 13442 -2001 13444
rect -2000 13442 -1992 13452
rect -1972 13450 -1958 13452
rect -1844 13451 -1804 13452
rect -1862 13449 -1796 13450
rect -1985 13447 -1796 13449
rect -1985 13442 -1852 13447
rect -2325 13430 -2320 13442
rect -2309 13430 -2301 13442
rect -2068 13432 -2060 13439
rect -2015 13432 -1990 13442
rect -1844 13441 -1796 13447
rect -1671 13442 -1663 13452
rect -1852 13432 -1804 13439
rect -2020 13430 -2004 13432
rect -2000 13430 -1992 13432
rect -1976 13430 -1940 13431
rect -1655 13430 -1647 13442
rect -1642 13430 -1637 13452
rect -1619 13430 -1614 13452
rect -1530 13431 -1526 13452
rect -1541 13430 -1507 13431
rect -2393 13428 -1507 13430
rect -2371 13358 -2366 13428
rect -2348 13358 -2343 13428
rect -2325 13426 -2320 13428
rect -2317 13426 -2309 13428
rect -2325 13414 -2317 13426
rect -2060 13415 -2030 13422
rect -2325 13394 -2320 13414
rect -2325 13386 -2317 13394
rect -2060 13388 -2030 13391
rect -2325 13366 -2320 13386
rect -2317 13378 -2309 13386
rect -2060 13375 -2038 13386
rect -2033 13379 -2030 13388
rect -2028 13384 -2027 13388
rect -2068 13370 -2038 13373
rect -2325 13358 -2317 13366
rect -2000 13358 -1992 13428
rect -1844 13424 -1804 13428
rect -1663 13426 -1655 13428
rect -1844 13414 -1794 13423
rect -1671 13414 -1663 13426
rect -1912 13403 -1884 13405
rect -1852 13397 -1804 13401
rect -1844 13388 -1796 13391
rect -1671 13386 -1663 13394
rect -1844 13375 -1804 13386
rect -1663 13378 -1655 13386
rect -1852 13370 -1680 13374
rect -1926 13358 -1892 13361
rect -1671 13358 -1663 13366
rect -1642 13358 -1637 13428
rect -1619 13358 -1614 13428
rect -1541 13421 -1536 13428
rect -1530 13421 -1526 13428
rect -1531 13407 -1526 13421
rect -1541 13397 -1536 13407
rect -1531 13383 -1526 13397
rect -1530 13358 -1526 13383
rect -1506 13358 -1502 13452
rect -1482 13358 -1478 13452
rect -1458 13358 -1454 13452
rect -1434 13358 -1430 13452
rect -1410 13358 -1406 13452
rect -1386 13358 -1382 13452
rect -1362 13358 -1358 13452
rect -1338 13358 -1334 13452
rect -1314 13358 -1310 13452
rect -1290 13358 -1286 13452
rect -1277 13397 -1272 13407
rect -1266 13397 -1262 13452
rect -1267 13383 -1262 13397
rect -1277 13382 -1243 13383
rect -1242 13382 -1238 13452
rect -1218 13382 -1214 13452
rect -1194 13382 -1190 13452
rect -1170 13382 -1166 13452
rect -1146 13382 -1142 13452
rect -1122 13382 -1118 13452
rect -1098 13382 -1094 13452
rect -1074 13382 -1070 13452
rect -1050 13382 -1046 13452
rect -1026 13382 -1022 13452
rect -1002 13382 -998 13452
rect -978 13382 -974 13452
rect -954 13382 -950 13452
rect -930 13382 -926 13452
rect -906 13382 -902 13452
rect -882 13382 -878 13452
rect -858 13382 -854 13452
rect -834 13382 -830 13452
rect -810 13382 -806 13452
rect -786 13382 -782 13452
rect -762 13382 -758 13452
rect -738 13382 -734 13452
rect -714 13382 -710 13452
rect -690 13382 -686 13452
rect -666 13382 -662 13452
rect -642 13382 -638 13452
rect -618 13382 -614 13452
rect -594 13382 -590 13452
rect -570 13382 -566 13452
rect -546 13382 -542 13452
rect -522 13382 -518 13452
rect -498 13382 -494 13452
rect -474 13382 -470 13452
rect -450 13382 -446 13452
rect -426 13382 -422 13452
rect -402 13382 -398 13452
rect -378 13382 -374 13452
rect -354 13382 -350 13452
rect -330 13382 -326 13452
rect -306 13382 -302 13452
rect -282 13382 -278 13452
rect -258 13382 -254 13452
rect -234 13382 -230 13452
rect -210 13382 -206 13452
rect -186 13382 -182 13452
rect -162 13382 -158 13452
rect -138 13382 -134 13452
rect -114 13382 -110 13452
rect -90 13382 -86 13452
rect -66 13382 -62 13452
rect -42 13382 -38 13452
rect -18 13382 -14 13452
rect 6 13382 10 13452
rect 30 13382 34 13452
rect 54 13382 58 13452
rect 78 13382 82 13452
rect 102 13382 106 13452
rect 126 13382 130 13452
rect 150 13382 154 13452
rect 174 13382 178 13452
rect 198 13382 202 13452
rect 222 13382 226 13452
rect 246 13451 250 13452
rect 246 13403 253 13451
rect 246 13382 250 13403
rect 270 13382 274 13452
rect 294 13382 298 13452
rect 318 13382 322 13452
rect 342 13382 346 13452
rect 366 13427 373 13451
rect 366 13382 370 13427
rect 390 13382 394 13452
rect 414 13382 418 13452
rect 438 13382 442 13452
rect 462 13382 466 13452
rect 486 13382 490 13452
rect 510 13382 514 13452
rect 534 13382 538 13452
rect 558 13382 562 13452
rect 582 13382 586 13452
rect 606 13382 610 13452
rect 630 13382 634 13452
rect 643 13445 648 13452
rect 654 13445 658 13452
rect 653 13431 658 13445
rect 654 13382 658 13431
rect 678 13382 682 13500
rect 702 13382 706 13500
rect 726 13382 730 13500
rect 750 13382 754 13500
rect 774 13382 778 13500
rect 798 13382 802 13500
rect 822 13382 826 13500
rect 846 13382 850 13500
rect 870 13382 874 13500
rect 894 13382 898 13500
rect 918 13382 922 13500
rect 942 13382 946 13500
rect 966 13382 970 13500
rect 990 13382 994 13500
rect 1014 13382 1018 13500
rect 1038 13382 1042 13500
rect 1062 13382 1066 13500
rect 1086 13382 1090 13500
rect 1110 13382 1114 13500
rect 1134 13382 1138 13500
rect 1147 13469 1152 13479
rect 1182 13475 1186 13500
rect 1157 13455 1162 13469
rect 1171 13465 1179 13469
rect 1165 13455 1171 13465
rect 1158 13382 1162 13455
rect 1182 13451 1189 13475
rect -1277 13380 1179 13382
rect -1277 13373 -1272 13380
rect -1267 13359 -1262 13373
rect -1266 13358 -1262 13359
rect -1242 13358 -1238 13380
rect -1218 13358 -1214 13380
rect -1194 13358 -1190 13380
rect -1170 13358 -1166 13380
rect -1146 13358 -1142 13380
rect -1122 13358 -1118 13380
rect -1098 13358 -1094 13380
rect -1074 13358 -1070 13380
rect -1050 13358 -1046 13380
rect -1026 13358 -1022 13380
rect -1002 13358 -998 13380
rect -978 13358 -974 13380
rect -954 13358 -950 13380
rect -930 13358 -926 13380
rect -906 13358 -902 13380
rect -882 13358 -878 13380
rect -858 13358 -854 13380
rect -834 13358 -830 13380
rect -810 13358 -806 13380
rect -786 13358 -782 13380
rect -762 13358 -758 13380
rect -738 13358 -734 13380
rect -714 13358 -710 13380
rect -690 13358 -686 13380
rect -666 13358 -662 13380
rect -642 13358 -638 13380
rect -618 13358 -614 13380
rect -594 13358 -590 13380
rect -570 13358 -566 13380
rect -546 13358 -542 13380
rect -522 13358 -518 13380
rect -498 13358 -494 13380
rect -474 13358 -470 13380
rect -450 13358 -446 13380
rect -426 13358 -422 13380
rect -402 13358 -398 13380
rect -378 13358 -374 13380
rect -354 13358 -350 13380
rect -330 13358 -326 13380
rect -306 13358 -302 13380
rect -282 13358 -278 13380
rect -258 13358 -254 13380
rect -234 13358 -230 13380
rect -210 13358 -206 13380
rect -186 13358 -182 13380
rect -162 13358 -158 13380
rect -138 13358 -134 13380
rect -114 13358 -110 13380
rect -90 13358 -86 13380
rect -66 13358 -62 13380
rect -42 13358 -38 13380
rect -18 13358 -14 13380
rect 6 13358 10 13380
rect 30 13358 34 13380
rect 54 13358 58 13380
rect 78 13358 82 13380
rect 102 13358 106 13380
rect 126 13358 130 13380
rect 150 13358 154 13380
rect 174 13358 178 13380
rect 198 13358 202 13380
rect 222 13358 226 13380
rect 246 13358 250 13380
rect 270 13358 274 13380
rect 294 13358 298 13380
rect 318 13358 322 13380
rect 342 13358 346 13380
rect 366 13358 370 13380
rect 390 13358 394 13380
rect 414 13358 418 13380
rect 438 13358 442 13380
rect 462 13358 466 13380
rect 486 13358 490 13380
rect 510 13358 514 13380
rect 534 13358 538 13380
rect 558 13358 562 13380
rect 582 13358 586 13380
rect 606 13358 610 13380
rect 630 13358 634 13380
rect 654 13358 658 13380
rect 678 13379 682 13380
rect -2393 13356 675 13358
rect -2371 13334 -2366 13356
rect -2348 13334 -2343 13356
rect -2325 13350 -2317 13356
rect -2325 13334 -2320 13350
rect -2309 13338 -2301 13350
rect -2068 13339 -2038 13346
rect -2317 13334 -2309 13338
rect -2000 13336 -1992 13356
rect -1844 13348 -1794 13356
rect -1671 13350 -1663 13356
rect -1852 13339 -1804 13346
rect -1655 13338 -1647 13350
rect -2025 13335 -1991 13336
rect -2025 13334 -1975 13335
rect -1844 13334 -1804 13337
rect -1663 13334 -1655 13338
rect -1642 13334 -1637 13356
rect -1619 13334 -1614 13356
rect -1530 13334 -1526 13356
rect -1506 13355 -1502 13356
rect -2393 13332 -1509 13334
rect -2371 13310 -2366 13332
rect -2348 13310 -2343 13332
rect -2325 13322 -2317 13332
rect -2060 13322 -2020 13329
rect -2004 13324 -2001 13329
rect -2015 13322 -2001 13324
rect -2000 13322 -1992 13332
rect -1972 13330 -1958 13332
rect -1844 13331 -1804 13332
rect -1862 13329 -1796 13330
rect -1985 13327 -1796 13329
rect -1985 13322 -1852 13327
rect -2325 13310 -2320 13322
rect -2309 13310 -2301 13322
rect -2068 13312 -2060 13319
rect -2015 13312 -1990 13322
rect -1844 13321 -1796 13327
rect -1671 13322 -1663 13332
rect -1852 13312 -1804 13319
rect -2020 13310 -2004 13312
rect -2000 13310 -1992 13312
rect -1976 13310 -1940 13311
rect -1655 13310 -1647 13322
rect -1642 13310 -1637 13332
rect -1619 13310 -1614 13332
rect -1530 13310 -1526 13332
rect -1523 13331 -1509 13332
rect -1506 13310 -1499 13355
rect -1482 13310 -1478 13356
rect -1458 13310 -1454 13356
rect -1434 13310 -1430 13356
rect -1410 13310 -1406 13356
rect -1386 13310 -1382 13356
rect -1362 13310 -1358 13356
rect -1338 13310 -1334 13356
rect -1314 13310 -1310 13356
rect -1290 13310 -1286 13356
rect -1266 13310 -1262 13356
rect -1242 13331 -1238 13356
rect -2393 13308 -1245 13310
rect -2371 13238 -2366 13308
rect -2348 13238 -2343 13308
rect -2325 13306 -2320 13308
rect -2317 13306 -2309 13308
rect -2325 13294 -2317 13306
rect -2060 13295 -2030 13302
rect -2325 13274 -2320 13294
rect -2325 13266 -2317 13274
rect -2060 13268 -2030 13271
rect -2325 13246 -2320 13266
rect -2317 13258 -2309 13266
rect -2060 13255 -2038 13266
rect -2033 13259 -2030 13268
rect -2028 13264 -2027 13268
rect -2068 13250 -2038 13253
rect -2325 13238 -2317 13246
rect -2000 13238 -1992 13308
rect -1844 13304 -1804 13308
rect -1663 13306 -1655 13308
rect -1844 13294 -1794 13303
rect -1671 13294 -1663 13306
rect -1912 13283 -1884 13285
rect -1852 13277 -1804 13281
rect -1844 13268 -1796 13271
rect -1671 13266 -1663 13274
rect -1844 13255 -1804 13266
rect -1663 13258 -1655 13266
rect -1852 13250 -1680 13254
rect -1926 13238 -1892 13241
rect -1671 13238 -1663 13246
rect -1642 13238 -1637 13308
rect -1619 13238 -1614 13308
rect -1530 13238 -1526 13308
rect -1523 13307 -1509 13308
rect -1506 13307 -1499 13308
rect -1506 13238 -1502 13307
rect -1482 13238 -1478 13308
rect -1458 13238 -1454 13308
rect -1434 13238 -1430 13308
rect -1410 13238 -1406 13308
rect -1386 13238 -1382 13308
rect -1362 13238 -1358 13308
rect -1338 13238 -1334 13308
rect -1314 13238 -1310 13308
rect -1290 13238 -1286 13308
rect -1266 13238 -1262 13308
rect -1259 13307 -1245 13308
rect -1242 13286 -1235 13331
rect -1218 13286 -1214 13356
rect -1194 13286 -1190 13356
rect -1170 13286 -1166 13356
rect -1146 13286 -1142 13356
rect -1122 13286 -1118 13356
rect -1098 13286 -1094 13356
rect -1074 13286 -1070 13356
rect -1050 13286 -1046 13356
rect -1026 13286 -1022 13356
rect -1002 13286 -998 13356
rect -978 13286 -974 13356
rect -954 13286 -950 13356
rect -930 13286 -926 13356
rect -906 13286 -902 13356
rect -882 13286 -878 13356
rect -858 13286 -854 13356
rect -834 13286 -830 13356
rect -810 13286 -806 13356
rect -786 13286 -782 13356
rect -762 13286 -758 13356
rect -738 13286 -734 13356
rect -714 13286 -710 13356
rect -690 13286 -686 13356
rect -666 13286 -662 13356
rect -642 13286 -638 13356
rect -618 13286 -614 13356
rect -594 13286 -590 13356
rect -570 13286 -566 13356
rect -546 13286 -542 13356
rect -522 13286 -518 13356
rect -498 13286 -494 13356
rect -474 13286 -470 13356
rect -450 13286 -446 13356
rect -426 13286 -422 13356
rect -402 13286 -398 13356
rect -378 13286 -374 13356
rect -354 13286 -350 13356
rect -330 13286 -326 13356
rect -306 13286 -302 13356
rect -282 13286 -278 13356
rect -258 13286 -254 13356
rect -234 13286 -230 13356
rect -210 13286 -206 13356
rect -186 13286 -182 13356
rect -162 13286 -158 13356
rect -138 13286 -134 13356
rect -114 13286 -110 13356
rect -90 13286 -86 13356
rect -66 13286 -62 13356
rect -42 13286 -38 13356
rect -18 13286 -14 13356
rect 6 13286 10 13356
rect 30 13286 34 13356
rect 54 13286 58 13356
rect 78 13286 82 13356
rect 102 13286 106 13356
rect 126 13286 130 13356
rect 150 13286 154 13356
rect 174 13286 178 13356
rect 198 13286 202 13356
rect 222 13286 226 13356
rect 246 13286 250 13356
rect 270 13286 274 13356
rect 294 13286 298 13356
rect 318 13286 322 13356
rect 342 13286 346 13356
rect 366 13286 370 13356
rect 390 13286 394 13356
rect 414 13286 418 13356
rect 438 13286 442 13356
rect 462 13286 466 13356
rect 486 13286 490 13356
rect 510 13286 514 13356
rect 534 13286 538 13356
rect 558 13286 562 13356
rect 582 13286 586 13356
rect 606 13286 610 13356
rect 630 13286 634 13356
rect 654 13286 658 13356
rect 661 13355 675 13356
rect 678 13355 685 13379
rect 678 13286 682 13355
rect 702 13286 706 13380
rect 726 13286 730 13380
rect 750 13286 754 13380
rect 774 13286 778 13380
rect 798 13286 802 13380
rect 822 13286 826 13380
rect 846 13286 850 13380
rect 870 13286 874 13380
rect 894 13286 898 13380
rect 918 13286 922 13380
rect 942 13287 946 13380
rect 931 13286 965 13287
rect -1259 13284 965 13286
rect -1259 13283 -1245 13284
rect -1242 13283 -1235 13284
rect -1242 13238 -1238 13283
rect -1218 13238 -1214 13284
rect -1194 13238 -1190 13284
rect -1170 13238 -1166 13284
rect -1146 13238 -1142 13284
rect -1122 13238 -1118 13284
rect -1098 13238 -1094 13284
rect -1074 13238 -1070 13284
rect -1050 13238 -1046 13284
rect -1026 13238 -1022 13284
rect -1002 13238 -998 13284
rect -978 13238 -974 13284
rect -954 13238 -950 13284
rect -930 13238 -926 13284
rect -906 13238 -902 13284
rect -882 13238 -878 13284
rect -858 13238 -854 13284
rect -834 13238 -830 13284
rect -810 13238 -806 13284
rect -786 13238 -782 13284
rect -762 13238 -758 13284
rect -738 13238 -734 13284
rect -714 13238 -710 13284
rect -690 13238 -686 13284
rect -666 13238 -662 13284
rect -642 13238 -638 13284
rect -618 13238 -614 13284
rect -594 13238 -590 13284
rect -570 13238 -566 13284
rect -546 13238 -542 13284
rect -522 13238 -518 13284
rect -498 13238 -494 13284
rect -474 13238 -470 13284
rect -450 13238 -446 13284
rect -426 13238 -422 13284
rect -402 13238 -398 13284
rect -378 13238 -374 13284
rect -354 13238 -350 13284
rect -330 13238 -326 13284
rect -306 13238 -302 13284
rect -282 13238 -278 13284
rect -258 13238 -254 13284
rect -234 13238 -230 13284
rect -210 13238 -206 13284
rect -186 13238 -182 13284
rect -162 13238 -158 13284
rect -138 13238 -134 13284
rect -114 13238 -110 13284
rect -90 13238 -86 13284
rect -66 13238 -62 13284
rect -42 13238 -38 13284
rect -18 13238 -14 13284
rect 6 13238 10 13284
rect 30 13238 34 13284
rect 54 13238 58 13284
rect 78 13238 82 13284
rect 102 13238 106 13284
rect 126 13238 130 13284
rect 150 13238 154 13284
rect 174 13238 178 13284
rect 198 13238 202 13284
rect 222 13238 226 13284
rect 246 13238 250 13284
rect 270 13238 274 13284
rect 294 13238 298 13284
rect 318 13238 322 13284
rect 342 13238 346 13284
rect 366 13238 370 13284
rect 390 13238 394 13284
rect 414 13238 418 13284
rect 438 13238 442 13284
rect 462 13238 466 13284
rect 486 13238 490 13284
rect 510 13238 514 13284
rect 534 13238 538 13284
rect 558 13238 562 13284
rect 582 13238 586 13284
rect 606 13238 610 13284
rect 630 13238 634 13284
rect 654 13238 658 13284
rect 678 13238 682 13284
rect 702 13238 706 13284
rect 726 13238 730 13284
rect 750 13238 754 13284
rect 774 13238 778 13284
rect 798 13238 802 13284
rect 822 13238 826 13284
rect 846 13238 850 13284
rect 870 13238 874 13284
rect 894 13238 898 13284
rect 918 13238 922 13284
rect 931 13277 936 13284
rect 942 13277 946 13284
rect 941 13263 946 13277
rect 931 13262 965 13263
rect 966 13262 970 13380
rect 990 13262 994 13380
rect 1014 13262 1018 13380
rect 1038 13262 1042 13380
rect 1062 13262 1066 13380
rect 1086 13262 1090 13380
rect 1110 13262 1114 13380
rect 1134 13262 1138 13380
rect 1158 13262 1162 13380
rect 1165 13379 1179 13380
rect 1182 13379 1189 13403
rect 1182 13262 1186 13379
rect 1206 13262 1210 13500
rect 1230 13262 1234 13500
rect 1254 13262 1258 13500
rect 1278 13262 1282 13500
rect 1302 13262 1306 13500
rect 1326 13262 1330 13500
rect 1350 13262 1354 13500
rect 1374 13262 1378 13500
rect 1398 13262 1402 13500
rect 1422 13262 1426 13500
rect 1446 13262 1450 13500
rect 1470 13262 1474 13500
rect 1494 13262 1498 13500
rect 1518 13262 1522 13500
rect 1542 13262 1546 13500
rect 1566 13262 1570 13500
rect 1590 13262 1594 13500
rect 1614 13262 1618 13500
rect 1638 13262 1642 13500
rect 1662 13262 1666 13500
rect 1686 13262 1690 13500
rect 1710 13262 1714 13500
rect 1734 13262 1738 13500
rect 1758 13262 1762 13500
rect 1782 13262 1786 13500
rect 1806 13262 1810 13500
rect 1830 13262 1834 13500
rect 1854 13262 1858 13500
rect 1878 13262 1882 13500
rect 1902 13262 1906 13500
rect 1926 13262 1930 13500
rect 1950 13262 1954 13500
rect 1974 13262 1978 13500
rect 1998 13262 2002 13500
rect 2022 13262 2026 13500
rect 2046 13262 2050 13500
rect 2070 13262 2074 13500
rect 2094 13262 2098 13500
rect 2118 13262 2122 13500
rect 2142 13262 2146 13500
rect 2166 13262 2170 13500
rect 2190 13262 2194 13500
rect 2214 13262 2218 13500
rect 2238 13262 2242 13500
rect 2262 13262 2266 13500
rect 2286 13262 2290 13500
rect 2310 13262 2314 13500
rect 2334 13262 2338 13500
rect 2358 13262 2362 13500
rect 2382 13262 2386 13500
rect 2406 13262 2410 13500
rect 2430 13262 2434 13500
rect 2454 13262 2458 13500
rect 2478 13262 2482 13500
rect 2502 13262 2506 13500
rect 2526 13262 2530 13500
rect 2539 13325 2544 13335
rect 2550 13325 2554 13500
rect 2549 13311 2554 13325
rect 2539 13301 2544 13311
rect 2549 13287 2554 13301
rect 2550 13262 2554 13287
rect 2574 13262 2578 13500
rect 2598 13262 2602 13500
rect 2622 13262 2626 13500
rect 2646 13262 2650 13500
rect 2670 13262 2674 13500
rect 2694 13262 2698 13500
rect 2718 13262 2722 13500
rect 2742 13262 2746 13500
rect 2766 13262 2770 13500
rect 2779 13301 2784 13311
rect 2790 13301 2794 13500
rect 2789 13287 2794 13301
rect 2779 13286 2813 13287
rect 2814 13286 2818 13500
rect 2838 13286 2842 13500
rect 2862 13286 2866 13500
rect 2886 13286 2890 13500
rect 2910 13286 2914 13500
rect 2934 13286 2938 13500
rect 2958 13286 2962 13500
rect 2982 13286 2986 13500
rect 3006 13286 3010 13500
rect 3030 13286 3034 13500
rect 3054 13286 3058 13500
rect 3078 13286 3082 13500
rect 3102 13286 3106 13500
rect 3126 13286 3130 13500
rect 3150 13286 3154 13500
rect 3174 13286 3178 13500
rect 3198 13286 3202 13500
rect 3222 13286 3226 13500
rect 3246 13286 3250 13500
rect 3270 13286 3274 13500
rect 3294 13286 3298 13500
rect 3318 13286 3322 13500
rect 3342 13286 3346 13500
rect 3366 13286 3370 13500
rect 3390 13286 3394 13500
rect 3414 13286 3418 13500
rect 3438 13286 3442 13500
rect 3462 13286 3466 13500
rect 3486 13286 3490 13500
rect 3510 13286 3514 13500
rect 3534 13286 3538 13500
rect 3547 13373 3552 13383
rect 3558 13373 3562 13500
rect 3571 13493 3576 13500
rect 3582 13493 3586 13500
rect 3581 13479 3586 13493
rect 3557 13359 3562 13373
rect 3547 13349 3552 13359
rect 3557 13335 3562 13349
rect 3558 13287 3562 13335
rect 3547 13286 3579 13287
rect 2779 13284 3579 13286
rect 2779 13277 2784 13284
rect 2789 13263 2794 13277
rect 2790 13262 2794 13263
rect 2814 13262 2818 13284
rect 2838 13262 2842 13284
rect 2862 13262 2866 13284
rect 2886 13262 2890 13284
rect 2910 13262 2914 13284
rect 2934 13262 2938 13284
rect 2958 13262 2962 13284
rect 2982 13262 2986 13284
rect 3006 13262 3010 13284
rect 3030 13262 3034 13284
rect 3054 13262 3058 13284
rect 3078 13262 3082 13284
rect 3102 13262 3106 13284
rect 3126 13262 3130 13284
rect 3150 13262 3154 13284
rect 3174 13262 3178 13284
rect 3198 13262 3202 13284
rect 3222 13262 3226 13284
rect 3246 13262 3250 13284
rect 3270 13262 3274 13284
rect 3294 13262 3298 13284
rect 3318 13262 3322 13284
rect 3342 13262 3346 13284
rect 3366 13262 3370 13284
rect 3390 13262 3394 13284
rect 3414 13262 3418 13284
rect 3438 13262 3442 13284
rect 3462 13262 3466 13284
rect 3486 13262 3490 13284
rect 3510 13262 3514 13284
rect 3534 13263 3538 13284
rect 3547 13277 3552 13284
rect 3558 13277 3562 13284
rect 3565 13283 3579 13284
rect 3557 13263 3562 13277
rect 3571 13273 3579 13277
rect 3565 13263 3571 13273
rect 3523 13262 3557 13263
rect 931 13260 3557 13262
rect 931 13253 936 13260
rect 941 13239 946 13253
rect 942 13238 946 13239
rect 966 13238 970 13260
rect 990 13238 994 13260
rect 1014 13238 1018 13260
rect 1038 13238 1042 13260
rect 1062 13238 1066 13260
rect 1086 13238 1090 13260
rect 1110 13238 1114 13260
rect 1134 13238 1138 13260
rect 1158 13238 1162 13260
rect 1182 13238 1186 13260
rect 1206 13238 1210 13260
rect 1230 13238 1234 13260
rect 1254 13238 1258 13260
rect 1278 13238 1282 13260
rect 1302 13238 1306 13260
rect 1326 13238 1330 13260
rect 1350 13238 1354 13260
rect 1374 13238 1378 13260
rect 1398 13238 1402 13260
rect 1422 13238 1426 13260
rect 1446 13238 1450 13260
rect 1470 13238 1474 13260
rect 1494 13238 1498 13260
rect 1518 13238 1522 13260
rect 1542 13238 1546 13260
rect 1566 13238 1570 13260
rect 1590 13238 1594 13260
rect 1614 13238 1618 13260
rect 1638 13238 1642 13260
rect 1662 13238 1666 13260
rect 1686 13238 1690 13260
rect 1710 13238 1714 13260
rect 1734 13238 1738 13260
rect 1758 13238 1762 13260
rect 1782 13238 1786 13260
rect 1806 13238 1810 13260
rect 1830 13238 1834 13260
rect 1854 13238 1858 13260
rect 1878 13238 1882 13260
rect 1902 13238 1906 13260
rect 1926 13238 1930 13260
rect 1950 13238 1954 13260
rect 1974 13238 1978 13260
rect 1998 13238 2002 13260
rect 2022 13238 2026 13260
rect 2046 13238 2050 13260
rect 2070 13238 2074 13260
rect 2094 13238 2098 13260
rect 2118 13238 2122 13260
rect 2142 13238 2146 13260
rect 2166 13238 2170 13260
rect 2190 13238 2194 13260
rect 2214 13238 2218 13260
rect 2238 13238 2242 13260
rect 2262 13238 2266 13260
rect 2286 13238 2290 13260
rect 2310 13238 2314 13260
rect 2334 13238 2338 13260
rect 2358 13238 2362 13260
rect 2382 13238 2386 13260
rect 2406 13238 2410 13260
rect 2430 13238 2434 13260
rect 2454 13238 2458 13260
rect 2478 13238 2482 13260
rect 2502 13238 2506 13260
rect 2526 13238 2530 13260
rect 2550 13238 2554 13260
rect 2574 13259 2578 13260
rect -2393 13236 2571 13238
rect -2371 13214 -2366 13236
rect -2348 13214 -2343 13236
rect -2325 13230 -2317 13236
rect -2325 13214 -2320 13230
rect -2309 13218 -2301 13230
rect -2068 13219 -2038 13226
rect -2317 13214 -2309 13218
rect -2000 13216 -1992 13236
rect -1844 13228 -1794 13236
rect -1671 13230 -1663 13236
rect -1852 13219 -1804 13226
rect -1655 13218 -1647 13230
rect -2025 13215 -1991 13216
rect -2025 13214 -1975 13215
rect -1844 13214 -1804 13217
rect -1663 13214 -1655 13218
rect -1642 13214 -1637 13236
rect -1619 13214 -1614 13236
rect -1530 13214 -1526 13236
rect -1506 13214 -1502 13236
rect -1482 13214 -1478 13236
rect -1458 13214 -1454 13236
rect -1434 13214 -1430 13236
rect -1410 13214 -1406 13236
rect -1386 13215 -1382 13236
rect -1397 13214 -1363 13215
rect -2393 13212 -1363 13214
rect -2371 13190 -2366 13212
rect -2348 13190 -2343 13212
rect -2325 13202 -2317 13212
rect -2060 13202 -2020 13209
rect -2004 13204 -2001 13209
rect -2015 13202 -2001 13204
rect -2000 13202 -1992 13212
rect -1972 13210 -1958 13212
rect -1844 13211 -1804 13212
rect -1862 13209 -1796 13210
rect -1985 13207 -1796 13209
rect -1985 13202 -1852 13207
rect -2325 13190 -2320 13202
rect -2309 13190 -2301 13202
rect -2068 13192 -2060 13199
rect -2015 13192 -1990 13202
rect -1844 13201 -1796 13207
rect -1671 13202 -1663 13212
rect -1852 13192 -1804 13199
rect -2020 13190 -2004 13192
rect -2000 13190 -1992 13192
rect -1976 13190 -1940 13191
rect -1655 13190 -1647 13202
rect -1642 13190 -1637 13212
rect -1619 13190 -1614 13212
rect -1530 13190 -1526 13212
rect -1506 13190 -1502 13212
rect -1482 13190 -1478 13212
rect -1458 13190 -1454 13212
rect -1434 13190 -1430 13212
rect -1410 13190 -1406 13212
rect -1397 13205 -1392 13212
rect -1386 13205 -1382 13212
rect -1387 13191 -1382 13205
rect -1386 13190 -1382 13191
rect -1362 13190 -1358 13236
rect -1338 13190 -1334 13236
rect -1314 13190 -1310 13236
rect -1290 13190 -1286 13236
rect -1266 13190 -1262 13236
rect -1242 13190 -1238 13236
rect -1218 13190 -1214 13236
rect -1194 13190 -1190 13236
rect -1170 13190 -1166 13236
rect -1146 13190 -1142 13236
rect -1122 13190 -1118 13236
rect -1098 13190 -1094 13236
rect -1074 13190 -1070 13236
rect -1050 13190 -1046 13236
rect -1026 13190 -1022 13236
rect -1002 13190 -998 13236
rect -978 13190 -974 13236
rect -954 13190 -950 13236
rect -930 13190 -926 13236
rect -906 13190 -902 13236
rect -882 13190 -878 13236
rect -858 13190 -854 13236
rect -834 13190 -830 13236
rect -810 13190 -806 13236
rect -786 13190 -782 13236
rect -762 13190 -758 13236
rect -738 13190 -734 13236
rect -714 13190 -710 13236
rect -690 13190 -686 13236
rect -666 13190 -662 13236
rect -642 13190 -638 13236
rect -618 13190 -614 13236
rect -594 13190 -590 13236
rect -570 13190 -566 13236
rect -546 13190 -542 13236
rect -522 13190 -518 13236
rect -498 13190 -494 13236
rect -474 13190 -470 13236
rect -450 13190 -446 13236
rect -426 13190 -422 13236
rect -402 13190 -398 13236
rect -378 13190 -374 13236
rect -354 13190 -350 13236
rect -330 13190 -326 13236
rect -306 13190 -302 13236
rect -282 13190 -278 13236
rect -258 13190 -254 13236
rect -234 13190 -230 13236
rect -210 13190 -206 13236
rect -186 13190 -182 13236
rect -162 13190 -158 13236
rect -138 13190 -134 13236
rect -114 13190 -110 13236
rect -90 13190 -86 13236
rect -66 13190 -62 13236
rect -42 13190 -38 13236
rect -18 13190 -14 13236
rect 6 13190 10 13236
rect 30 13190 34 13236
rect 54 13190 58 13236
rect 78 13190 82 13236
rect 102 13190 106 13236
rect 126 13190 130 13236
rect 150 13190 154 13236
rect 174 13190 178 13236
rect 198 13190 202 13236
rect 222 13190 226 13236
rect 246 13190 250 13236
rect 270 13190 274 13236
rect 294 13190 298 13236
rect 318 13190 322 13236
rect 342 13190 346 13236
rect 366 13190 370 13236
rect 390 13190 394 13236
rect 414 13190 418 13236
rect 438 13190 442 13236
rect 462 13190 466 13236
rect 486 13190 490 13236
rect 510 13190 514 13236
rect 534 13190 538 13236
rect 558 13190 562 13236
rect 582 13190 586 13236
rect 606 13190 610 13236
rect 630 13190 634 13236
rect 654 13190 658 13236
rect 678 13190 682 13236
rect 702 13190 706 13236
rect 726 13190 730 13236
rect 750 13190 754 13236
rect 774 13190 778 13236
rect 798 13190 802 13236
rect 822 13190 826 13236
rect 846 13190 850 13236
rect 870 13190 874 13236
rect 894 13190 898 13236
rect 918 13190 922 13236
rect 942 13190 946 13236
rect 966 13211 970 13236
rect -2393 13188 963 13190
rect -2371 13118 -2366 13188
rect -2348 13118 -2343 13188
rect -2325 13186 -2320 13188
rect -2317 13186 -2309 13188
rect -2325 13174 -2317 13186
rect -2060 13175 -2030 13182
rect -2325 13154 -2320 13174
rect -2325 13146 -2317 13154
rect -2060 13148 -2030 13151
rect -2325 13126 -2320 13146
rect -2317 13138 -2309 13146
rect -2060 13135 -2038 13146
rect -2033 13139 -2030 13148
rect -2028 13144 -2027 13148
rect -2068 13130 -2038 13133
rect -2325 13118 -2317 13126
rect -2000 13118 -1992 13188
rect -1844 13184 -1804 13188
rect -1663 13186 -1655 13188
rect -1844 13174 -1794 13183
rect -1671 13174 -1663 13186
rect -1912 13163 -1884 13165
rect -1852 13157 -1804 13161
rect -1844 13148 -1796 13151
rect -1671 13146 -1663 13154
rect -1844 13135 -1804 13146
rect -1663 13138 -1655 13146
rect -1852 13130 -1680 13134
rect -1926 13118 -1892 13121
rect -1671 13118 -1663 13126
rect -1642 13118 -1637 13188
rect -1619 13118 -1614 13188
rect -1530 13118 -1526 13188
rect -1506 13118 -1502 13188
rect -1482 13118 -1478 13188
rect -1458 13118 -1454 13188
rect -1434 13118 -1430 13188
rect -1410 13118 -1406 13188
rect -1386 13118 -1382 13188
rect -1362 13139 -1358 13188
rect -2393 13116 -1365 13118
rect -2371 13094 -2366 13116
rect -2348 13094 -2343 13116
rect -2325 13110 -2317 13116
rect -2325 13094 -2320 13110
rect -2309 13098 -2301 13110
rect -2068 13099 -2038 13106
rect -2317 13094 -2309 13098
rect -2000 13096 -1992 13116
rect -1844 13108 -1794 13116
rect -1671 13110 -1663 13116
rect -1852 13099 -1804 13106
rect -1655 13098 -1647 13110
rect -2025 13095 -1991 13096
rect -2025 13094 -1975 13095
rect -1844 13094 -1804 13097
rect -1663 13094 -1655 13098
rect -1642 13094 -1637 13116
rect -1619 13094 -1614 13116
rect -1530 13094 -1526 13116
rect -1506 13094 -1502 13116
rect -1482 13094 -1478 13116
rect -1458 13094 -1454 13116
rect -1434 13094 -1430 13116
rect -1410 13094 -1406 13116
rect -1386 13094 -1382 13116
rect -1379 13115 -1365 13116
rect -1362 13115 -1355 13139
rect -1362 13094 -1358 13115
rect -1338 13094 -1334 13188
rect -1314 13094 -1310 13188
rect -1290 13094 -1286 13188
rect -1266 13094 -1262 13188
rect -1242 13094 -1238 13188
rect -1218 13094 -1214 13188
rect -1194 13094 -1190 13188
rect -1170 13094 -1166 13188
rect -1146 13094 -1142 13188
rect -1122 13094 -1118 13188
rect -1098 13094 -1094 13188
rect -1074 13094 -1070 13188
rect -1050 13094 -1046 13188
rect -1026 13094 -1022 13188
rect -1002 13094 -998 13188
rect -978 13094 -974 13188
rect -954 13094 -950 13188
rect -930 13094 -926 13188
rect -906 13094 -902 13188
rect -882 13094 -878 13188
rect -858 13094 -854 13188
rect -834 13094 -830 13188
rect -810 13094 -806 13188
rect -786 13094 -782 13188
rect -762 13094 -758 13188
rect -738 13094 -734 13188
rect -714 13094 -710 13188
rect -690 13094 -686 13188
rect -666 13094 -662 13188
rect -642 13094 -638 13188
rect -618 13094 -614 13188
rect -594 13094 -590 13188
rect -570 13094 -566 13188
rect -546 13094 -542 13188
rect -522 13094 -518 13188
rect -498 13094 -494 13188
rect -474 13094 -470 13188
rect -450 13094 -446 13188
rect -426 13094 -422 13188
rect -402 13094 -398 13188
rect -378 13094 -374 13188
rect -354 13094 -350 13188
rect -330 13094 -326 13188
rect -306 13094 -302 13188
rect -282 13094 -278 13188
rect -258 13094 -254 13188
rect -234 13094 -230 13188
rect -210 13094 -206 13188
rect -186 13094 -182 13188
rect -162 13094 -158 13188
rect -138 13094 -134 13188
rect -114 13094 -110 13188
rect -90 13094 -86 13188
rect -66 13094 -62 13188
rect -42 13094 -38 13188
rect -18 13094 -14 13188
rect 6 13094 10 13188
rect 30 13094 34 13188
rect 54 13094 58 13188
rect 78 13094 82 13188
rect 102 13094 106 13188
rect 126 13094 130 13188
rect 150 13094 154 13188
rect 174 13094 178 13188
rect 198 13094 202 13188
rect 222 13094 226 13188
rect 246 13094 250 13188
rect 270 13094 274 13188
rect 294 13094 298 13188
rect 318 13094 322 13188
rect 342 13094 346 13188
rect 366 13094 370 13188
rect 390 13094 394 13188
rect 414 13094 418 13188
rect 438 13094 442 13188
rect 462 13094 466 13188
rect 475 13157 480 13167
rect 486 13157 490 13188
rect 485 13143 490 13157
rect 475 13142 509 13143
rect 510 13142 514 13188
rect 534 13142 538 13188
rect 558 13142 562 13188
rect 582 13142 586 13188
rect 606 13142 610 13188
rect 630 13142 634 13188
rect 654 13142 658 13188
rect 678 13142 682 13188
rect 702 13142 706 13188
rect 726 13142 730 13188
rect 750 13142 754 13188
rect 774 13142 778 13188
rect 798 13142 802 13188
rect 822 13142 826 13188
rect 846 13142 850 13188
rect 870 13142 874 13188
rect 894 13142 898 13188
rect 918 13142 922 13188
rect 942 13142 946 13188
rect 949 13187 963 13188
rect 966 13163 973 13211
rect 966 13142 970 13163
rect 990 13142 994 13236
rect 1014 13142 1018 13236
rect 1038 13142 1042 13236
rect 1062 13142 1066 13236
rect 1086 13142 1090 13236
rect 1110 13142 1114 13236
rect 1134 13142 1138 13236
rect 1158 13142 1162 13236
rect 1182 13142 1186 13236
rect 1206 13142 1210 13236
rect 1230 13142 1234 13236
rect 1254 13142 1258 13236
rect 1278 13142 1282 13236
rect 1302 13142 1306 13236
rect 1326 13142 1330 13236
rect 1350 13142 1354 13236
rect 1374 13142 1378 13236
rect 1398 13142 1402 13236
rect 1422 13142 1426 13236
rect 1446 13142 1450 13236
rect 1470 13142 1474 13236
rect 1494 13142 1498 13236
rect 1518 13142 1522 13236
rect 1542 13142 1546 13236
rect 1566 13142 1570 13236
rect 1590 13142 1594 13236
rect 1614 13142 1618 13236
rect 1638 13142 1642 13236
rect 1662 13142 1666 13236
rect 1686 13142 1690 13236
rect 1710 13142 1714 13236
rect 1734 13142 1738 13236
rect 1758 13142 1762 13236
rect 1782 13142 1786 13236
rect 1806 13142 1810 13236
rect 1830 13142 1834 13236
rect 1854 13142 1858 13236
rect 1878 13142 1882 13236
rect 1902 13142 1906 13236
rect 1926 13142 1930 13236
rect 1950 13142 1954 13236
rect 1974 13142 1978 13236
rect 1998 13142 2002 13236
rect 2022 13142 2026 13236
rect 2046 13142 2050 13236
rect 2070 13142 2074 13236
rect 2094 13142 2098 13236
rect 2118 13142 2122 13236
rect 2142 13142 2146 13236
rect 2166 13142 2170 13236
rect 2190 13142 2194 13236
rect 2214 13142 2218 13236
rect 2238 13142 2242 13236
rect 2262 13142 2266 13236
rect 2286 13142 2290 13236
rect 2310 13142 2314 13236
rect 2334 13142 2338 13236
rect 2358 13142 2362 13236
rect 2382 13142 2386 13236
rect 2406 13142 2410 13236
rect 2430 13142 2434 13236
rect 2454 13142 2458 13236
rect 2478 13142 2482 13236
rect 2502 13142 2506 13236
rect 2526 13142 2530 13236
rect 2539 13181 2544 13191
rect 2550 13181 2554 13236
rect 2557 13235 2571 13236
rect 2549 13167 2554 13181
rect 2574 13211 2581 13259
rect 2539 13166 2573 13167
rect 2574 13166 2578 13211
rect 2598 13166 2602 13260
rect 2622 13166 2626 13260
rect 2646 13166 2650 13260
rect 2670 13166 2674 13260
rect 2694 13166 2698 13260
rect 2718 13166 2722 13260
rect 2742 13166 2746 13260
rect 2766 13166 2770 13260
rect 2790 13166 2794 13260
rect 2814 13235 2818 13260
rect 2814 13187 2821 13235
rect 2814 13166 2818 13187
rect 2838 13166 2842 13260
rect 2862 13166 2866 13260
rect 2886 13166 2890 13260
rect 2910 13166 2914 13260
rect 2934 13166 2938 13260
rect 2958 13166 2962 13260
rect 2982 13166 2986 13260
rect 3006 13166 3010 13260
rect 3030 13166 3034 13260
rect 3054 13166 3058 13260
rect 3078 13166 3082 13260
rect 3102 13166 3106 13260
rect 3126 13166 3130 13260
rect 3150 13166 3154 13260
rect 3174 13166 3178 13260
rect 3198 13166 3202 13260
rect 3222 13166 3226 13260
rect 3246 13166 3250 13260
rect 3270 13166 3274 13260
rect 3294 13166 3298 13260
rect 3318 13166 3322 13260
rect 3342 13166 3346 13260
rect 3366 13166 3370 13260
rect 3390 13166 3394 13260
rect 3414 13166 3418 13260
rect 3438 13166 3442 13260
rect 3462 13166 3466 13260
rect 3486 13166 3490 13260
rect 3510 13166 3514 13260
rect 3523 13253 3528 13260
rect 3534 13253 3538 13260
rect 3533 13239 3538 13253
rect 3523 13229 3528 13239
rect 3533 13215 3538 13229
rect 3534 13167 3538 13215
rect 3523 13166 3555 13167
rect 2539 13164 3555 13166
rect 2539 13157 2544 13164
rect 2549 13143 2554 13157
rect 2550 13142 2554 13143
rect 2574 13142 2578 13164
rect 2598 13142 2602 13164
rect 2622 13142 2626 13164
rect 2646 13142 2650 13164
rect 2670 13142 2674 13164
rect 2694 13142 2698 13164
rect 2718 13142 2722 13164
rect 2742 13142 2746 13164
rect 2766 13142 2770 13164
rect 2790 13142 2794 13164
rect 2814 13142 2818 13164
rect 2838 13142 2842 13164
rect 2862 13142 2866 13164
rect 2886 13142 2890 13164
rect 2910 13142 2914 13164
rect 2934 13142 2938 13164
rect 2958 13142 2962 13164
rect 2982 13142 2986 13164
rect 3006 13142 3010 13164
rect 3030 13142 3034 13164
rect 3054 13142 3058 13164
rect 3078 13142 3082 13164
rect 3102 13142 3106 13164
rect 3126 13142 3130 13164
rect 3150 13142 3154 13164
rect 3174 13142 3178 13164
rect 3198 13142 3202 13164
rect 3222 13142 3226 13164
rect 3246 13142 3250 13164
rect 3270 13142 3274 13164
rect 3294 13142 3298 13164
rect 3318 13142 3322 13164
rect 3342 13142 3346 13164
rect 3366 13142 3370 13164
rect 3390 13142 3394 13164
rect 3414 13142 3418 13164
rect 3438 13142 3442 13164
rect 3462 13142 3466 13164
rect 3486 13142 3490 13164
rect 3510 13143 3514 13164
rect 3523 13157 3528 13164
rect 3534 13157 3538 13164
rect 3541 13163 3555 13164
rect 3533 13143 3538 13157
rect 3547 13153 3555 13157
rect 3541 13143 3547 13153
rect 3499 13142 3533 13143
rect 475 13140 3533 13142
rect 475 13133 480 13140
rect 485 13119 490 13133
rect 486 13094 490 13119
rect 510 13094 514 13140
rect 534 13094 538 13140
rect 558 13094 562 13140
rect 582 13094 586 13140
rect 606 13094 610 13140
rect 630 13094 634 13140
rect 654 13095 658 13140
rect 643 13094 677 13095
rect -2393 13092 677 13094
rect -2371 13070 -2366 13092
rect -2348 13070 -2343 13092
rect -2325 13082 -2317 13092
rect -2060 13082 -2020 13089
rect -2004 13084 -2001 13089
rect -2015 13082 -2001 13084
rect -2000 13082 -1992 13092
rect -1972 13090 -1958 13092
rect -1844 13091 -1804 13092
rect -1862 13089 -1796 13090
rect -1985 13087 -1796 13089
rect -1985 13082 -1852 13087
rect -2325 13070 -2320 13082
rect -2309 13070 -2301 13082
rect -2068 13072 -2060 13079
rect -2015 13072 -1990 13082
rect -1844 13081 -1796 13087
rect -1671 13082 -1663 13092
rect -1852 13072 -1804 13079
rect -2020 13070 -2004 13072
rect -2000 13070 -1992 13072
rect -1976 13070 -1940 13071
rect -1655 13070 -1647 13082
rect -1642 13070 -1637 13092
rect -1619 13070 -1614 13092
rect -1530 13070 -1526 13092
rect -1506 13070 -1502 13092
rect -1482 13070 -1478 13092
rect -1458 13070 -1454 13092
rect -1434 13070 -1430 13092
rect -1410 13070 -1406 13092
rect -1386 13070 -1382 13092
rect -1362 13070 -1358 13092
rect -1338 13070 -1334 13092
rect -1314 13070 -1310 13092
rect -1290 13070 -1286 13092
rect -1266 13070 -1262 13092
rect -1242 13070 -1238 13092
rect -1218 13070 -1214 13092
rect -1194 13070 -1190 13092
rect -1170 13070 -1166 13092
rect -1146 13070 -1142 13092
rect -1122 13070 -1118 13092
rect -1098 13070 -1094 13092
rect -1074 13070 -1070 13092
rect -1050 13071 -1046 13092
rect -1061 13070 -1027 13071
rect -2393 13068 -1027 13070
rect -2371 12998 -2366 13068
rect -2348 12998 -2343 13068
rect -2325 13066 -2320 13068
rect -2317 13066 -2309 13068
rect -2325 13054 -2317 13066
rect -2060 13055 -2030 13062
rect -2325 13034 -2320 13054
rect -2325 13026 -2317 13034
rect -2060 13028 -2030 13031
rect -2325 13006 -2320 13026
rect -2317 13018 -2309 13026
rect -2060 13015 -2038 13026
rect -2033 13019 -2030 13028
rect -2028 13024 -2027 13028
rect -2068 13010 -2038 13013
rect -2325 12998 -2317 13006
rect -2000 12998 -1992 13068
rect -1844 13064 -1804 13068
rect -1663 13066 -1655 13068
rect -1844 13054 -1794 13063
rect -1671 13054 -1663 13066
rect -1912 13043 -1884 13045
rect -1852 13037 -1804 13041
rect -1844 13028 -1796 13031
rect -1671 13026 -1663 13034
rect -1844 13015 -1804 13026
rect -1663 13018 -1655 13026
rect -1852 13010 -1680 13014
rect -1926 12998 -1892 13001
rect -1671 12998 -1663 13006
rect -1642 12998 -1637 13068
rect -1619 12998 -1614 13068
rect -1530 12998 -1526 13068
rect -1506 12998 -1502 13068
rect -1482 12998 -1478 13068
rect -1458 12998 -1454 13068
rect -1434 12998 -1430 13068
rect -1410 12998 -1406 13068
rect -1386 12998 -1382 13068
rect -1362 12998 -1358 13068
rect -1338 12998 -1334 13068
rect -1314 12998 -1310 13068
rect -1290 12998 -1286 13068
rect -1266 12998 -1262 13068
rect -1242 12998 -1238 13068
rect -1218 12998 -1214 13068
rect -1194 12998 -1190 13068
rect -1170 12998 -1166 13068
rect -1146 12998 -1142 13068
rect -1122 12998 -1118 13068
rect -1098 12998 -1094 13068
rect -1074 12998 -1070 13068
rect -1061 13061 -1056 13068
rect -1050 13061 -1046 13068
rect -1051 13047 -1046 13061
rect -1050 12998 -1046 13047
rect -1026 12998 -1022 13092
rect -1002 12998 -998 13092
rect -978 12998 -974 13092
rect -954 12998 -950 13092
rect -930 12998 -926 13092
rect -906 12998 -902 13092
rect -882 12998 -878 13092
rect -858 12998 -854 13092
rect -834 12998 -830 13092
rect -810 12998 -806 13092
rect -786 12998 -782 13092
rect -762 12998 -758 13092
rect -738 12998 -734 13092
rect -714 12998 -710 13092
rect -690 12998 -686 13092
rect -666 12998 -662 13092
rect -642 12998 -638 13092
rect -618 12998 -614 13092
rect -594 12998 -590 13092
rect -570 12998 -566 13092
rect -546 12998 -542 13092
rect -522 12998 -518 13092
rect -498 12998 -494 13092
rect -474 12998 -470 13092
rect -450 12998 -446 13092
rect -426 12998 -422 13092
rect -402 12998 -398 13092
rect -378 12998 -374 13092
rect -354 12998 -350 13092
rect -330 12998 -326 13092
rect -306 12998 -302 13092
rect -282 12998 -278 13092
rect -258 12998 -254 13092
rect -234 12998 -230 13092
rect -210 12998 -206 13092
rect -186 12998 -182 13092
rect -162 12998 -158 13092
rect -138 12998 -134 13092
rect -114 12998 -110 13092
rect -90 12998 -86 13092
rect -66 12998 -62 13092
rect -42 12998 -38 13092
rect -18 12998 -14 13092
rect 6 12998 10 13092
rect 30 12998 34 13092
rect 54 12998 58 13092
rect 78 12998 82 13092
rect 102 12998 106 13092
rect 126 12998 130 13092
rect 150 12998 154 13092
rect 174 12998 178 13092
rect 198 12998 202 13092
rect 222 12998 226 13092
rect 246 12998 250 13092
rect 270 12998 274 13092
rect 294 12998 298 13092
rect 318 12998 322 13092
rect 342 12998 346 13092
rect 366 12998 370 13092
rect 390 12998 394 13092
rect 414 12998 418 13092
rect 438 12998 442 13092
rect 462 12998 466 13092
rect 486 12998 490 13092
rect 510 13091 514 13092
rect 510 13046 517 13091
rect 534 13046 538 13092
rect 558 13046 562 13092
rect 582 13046 586 13092
rect 606 13046 610 13092
rect 630 13046 634 13092
rect 643 13085 648 13092
rect 654 13085 658 13092
rect 653 13071 658 13085
rect 643 13061 648 13071
rect 653 13047 658 13061
rect 654 13046 658 13047
rect 678 13046 682 13140
rect 702 13046 706 13140
rect 726 13046 730 13140
rect 750 13046 754 13140
rect 774 13046 778 13140
rect 798 13046 802 13140
rect 822 13046 826 13140
rect 846 13046 850 13140
rect 870 13046 874 13140
rect 894 13046 898 13140
rect 918 13046 922 13140
rect 942 13046 946 13140
rect 966 13046 970 13140
rect 990 13046 994 13140
rect 1014 13046 1018 13140
rect 1038 13046 1042 13140
rect 1062 13046 1066 13140
rect 1086 13046 1090 13140
rect 1110 13046 1114 13140
rect 1134 13046 1138 13140
rect 1158 13046 1162 13140
rect 1182 13046 1186 13140
rect 1206 13046 1210 13140
rect 1230 13046 1234 13140
rect 1254 13046 1258 13140
rect 1278 13046 1282 13140
rect 1302 13046 1306 13140
rect 1326 13046 1330 13140
rect 1350 13046 1354 13140
rect 1374 13046 1378 13140
rect 1398 13046 1402 13140
rect 1422 13046 1426 13140
rect 1446 13046 1450 13140
rect 1470 13046 1474 13140
rect 1494 13046 1498 13140
rect 1518 13046 1522 13140
rect 1542 13046 1546 13140
rect 1566 13046 1570 13140
rect 1590 13046 1594 13140
rect 1614 13046 1618 13140
rect 1638 13046 1642 13140
rect 1662 13046 1666 13140
rect 1686 13046 1690 13140
rect 1710 13046 1714 13140
rect 1734 13046 1738 13140
rect 1758 13046 1762 13140
rect 1782 13046 1786 13140
rect 1806 13046 1810 13140
rect 1830 13046 1834 13140
rect 1854 13046 1858 13140
rect 1878 13046 1882 13140
rect 1902 13046 1906 13140
rect 1926 13046 1930 13140
rect 1950 13046 1954 13140
rect 1974 13046 1978 13140
rect 1998 13046 2002 13140
rect 2022 13046 2026 13140
rect 2046 13046 2050 13140
rect 2070 13046 2074 13140
rect 2094 13046 2098 13140
rect 2118 13046 2122 13140
rect 2142 13046 2146 13140
rect 2166 13046 2170 13140
rect 2190 13046 2194 13140
rect 2214 13046 2218 13140
rect 2238 13046 2242 13140
rect 2262 13046 2266 13140
rect 2286 13046 2290 13140
rect 2310 13046 2314 13140
rect 2334 13046 2338 13140
rect 2358 13046 2362 13140
rect 2382 13046 2386 13140
rect 2406 13046 2410 13140
rect 2430 13046 2434 13140
rect 2454 13046 2458 13140
rect 2478 13046 2482 13140
rect 2502 13046 2506 13140
rect 2526 13046 2530 13140
rect 2550 13046 2554 13140
rect 2574 13115 2578 13140
rect 2574 13070 2581 13115
rect 2598 13070 2602 13140
rect 2622 13070 2626 13140
rect 2646 13070 2650 13140
rect 2670 13070 2674 13140
rect 2694 13070 2698 13140
rect 2718 13070 2722 13140
rect 2742 13070 2746 13140
rect 2766 13070 2770 13140
rect 2790 13070 2794 13140
rect 2814 13070 2818 13140
rect 2838 13070 2842 13140
rect 2862 13070 2866 13140
rect 2886 13070 2890 13140
rect 2910 13070 2914 13140
rect 2934 13070 2938 13140
rect 2958 13070 2962 13140
rect 2982 13070 2986 13140
rect 3006 13070 3010 13140
rect 3030 13070 3034 13140
rect 3054 13070 3058 13140
rect 3078 13070 3082 13140
rect 3102 13070 3106 13140
rect 3126 13070 3130 13140
rect 3150 13070 3154 13140
rect 3174 13070 3178 13140
rect 3198 13070 3202 13140
rect 3222 13070 3226 13140
rect 3246 13070 3250 13140
rect 3270 13070 3274 13140
rect 3294 13070 3298 13140
rect 3318 13070 3322 13140
rect 3342 13070 3346 13140
rect 3366 13070 3370 13140
rect 3390 13070 3394 13140
rect 3414 13070 3418 13140
rect 3438 13070 3442 13140
rect 3462 13070 3466 13140
rect 3486 13070 3490 13140
rect 3499 13133 3504 13140
rect 3510 13133 3514 13140
rect 3509 13119 3514 13133
rect 3499 13109 3504 13119
rect 3509 13095 3514 13109
rect 3510 13071 3514 13095
rect 3499 13070 3533 13071
rect 2557 13068 3533 13070
rect 2557 13067 2571 13068
rect 2574 13067 2581 13068
rect 2574 13046 2578 13067
rect 2598 13046 2602 13068
rect 2622 13046 2626 13068
rect 2646 13046 2650 13068
rect 2670 13046 2674 13068
rect 2694 13046 2698 13068
rect 2718 13046 2722 13068
rect 2742 13046 2746 13068
rect 2766 13046 2770 13068
rect 2790 13046 2794 13068
rect 2814 13046 2818 13068
rect 2838 13046 2842 13068
rect 2862 13046 2866 13068
rect 2886 13046 2890 13068
rect 2910 13046 2914 13068
rect 2934 13046 2938 13068
rect 2958 13046 2962 13068
rect 2982 13046 2986 13068
rect 3006 13046 3010 13068
rect 3030 13046 3034 13068
rect 3054 13046 3058 13068
rect 3078 13046 3082 13068
rect 3102 13046 3106 13068
rect 3126 13046 3130 13068
rect 3150 13047 3154 13068
rect 3139 13046 3173 13047
rect 493 13044 3173 13046
rect 493 13043 507 13044
rect 510 13043 517 13044
rect 510 12998 514 13043
rect 534 12998 538 13044
rect 558 12998 562 13044
rect 582 12998 586 13044
rect 606 12998 610 13044
rect 630 12998 634 13044
rect 654 12998 658 13044
rect 678 13019 682 13044
rect -2393 12996 675 12998
rect -2371 12974 -2366 12996
rect -2348 12974 -2343 12996
rect -2325 12990 -2317 12996
rect -2325 12974 -2320 12990
rect -2309 12978 -2301 12990
rect -2068 12979 -2038 12986
rect -2317 12974 -2309 12978
rect -2000 12976 -1992 12996
rect -1844 12988 -1794 12996
rect -1671 12990 -1663 12996
rect -1852 12979 -1804 12986
rect -1655 12978 -1647 12990
rect -2025 12975 -1991 12976
rect -2025 12974 -1975 12975
rect -1844 12974 -1804 12977
rect -1663 12974 -1655 12978
rect -1642 12974 -1637 12996
rect -1619 12974 -1614 12996
rect -1530 12974 -1526 12996
rect -1506 12974 -1502 12996
rect -1482 12974 -1478 12996
rect -1458 12974 -1454 12996
rect -1434 12974 -1430 12996
rect -1410 12974 -1406 12996
rect -1386 12974 -1382 12996
rect -1362 12974 -1358 12996
rect -1338 12974 -1334 12996
rect -1314 12974 -1310 12996
rect -1290 12974 -1286 12996
rect -1266 12974 -1262 12996
rect -1242 12974 -1238 12996
rect -1218 12974 -1214 12996
rect -1194 12974 -1190 12996
rect -1170 12974 -1166 12996
rect -1146 12974 -1142 12996
rect -1122 12974 -1118 12996
rect -1098 12974 -1094 12996
rect -1074 12974 -1070 12996
rect -1050 12974 -1046 12996
rect -1026 12995 -1022 12996
rect -2393 12972 -1029 12974
rect -2371 12950 -2366 12972
rect -2348 12950 -2343 12972
rect -2325 12962 -2317 12972
rect -2060 12962 -2020 12969
rect -2004 12964 -2001 12969
rect -2015 12962 -2001 12964
rect -2000 12962 -1992 12972
rect -1972 12970 -1958 12972
rect -1844 12971 -1804 12972
rect -1862 12969 -1796 12970
rect -1985 12967 -1796 12969
rect -1985 12962 -1852 12967
rect -2325 12950 -2320 12962
rect -2309 12950 -2301 12962
rect -2068 12952 -2060 12959
rect -2015 12952 -1990 12962
rect -1844 12961 -1796 12967
rect -1671 12962 -1663 12972
rect -1852 12952 -1804 12959
rect -2020 12950 -2004 12952
rect -2000 12950 -1992 12952
rect -1976 12950 -1940 12951
rect -1655 12950 -1647 12962
rect -1642 12950 -1637 12972
rect -1619 12950 -1614 12972
rect -1530 12950 -1526 12972
rect -1506 12950 -1502 12972
rect -1482 12950 -1478 12972
rect -1458 12950 -1454 12972
rect -1434 12950 -1430 12972
rect -1410 12950 -1406 12972
rect -1386 12950 -1382 12972
rect -1362 12950 -1358 12972
rect -1338 12950 -1334 12972
rect -1314 12950 -1310 12972
rect -1290 12950 -1286 12972
rect -1266 12950 -1262 12972
rect -1242 12950 -1238 12972
rect -1218 12950 -1214 12972
rect -1194 12950 -1190 12972
rect -1170 12950 -1166 12972
rect -1146 12950 -1142 12972
rect -1122 12950 -1118 12972
rect -1098 12950 -1094 12972
rect -1074 12950 -1070 12972
rect -1050 12951 -1046 12972
rect -1043 12971 -1029 12972
rect -1026 12971 -1019 12995
rect -1061 12950 -1027 12951
rect -2393 12948 -1027 12950
rect -2371 12878 -2366 12948
rect -2348 12878 -2343 12948
rect -2325 12946 -2320 12948
rect -2317 12946 -2309 12948
rect -2325 12934 -2317 12946
rect -2060 12935 -2030 12942
rect -2325 12914 -2320 12934
rect -2325 12906 -2317 12914
rect -2060 12908 -2030 12911
rect -2325 12886 -2320 12906
rect -2317 12898 -2309 12906
rect -2060 12895 -2038 12906
rect -2033 12899 -2030 12908
rect -2028 12904 -2027 12908
rect -2068 12890 -2038 12893
rect -2325 12878 -2317 12886
rect -2000 12878 -1992 12948
rect -1844 12944 -1804 12948
rect -1663 12946 -1655 12948
rect -1844 12934 -1794 12943
rect -1671 12934 -1663 12946
rect -1912 12923 -1884 12925
rect -1852 12917 -1804 12921
rect -1844 12908 -1796 12911
rect -1671 12906 -1663 12914
rect -1844 12895 -1804 12906
rect -1663 12898 -1655 12906
rect -1852 12890 -1680 12894
rect -1926 12878 -1892 12881
rect -1671 12878 -1663 12886
rect -1642 12878 -1637 12948
rect -1619 12878 -1614 12948
rect -1530 12878 -1526 12948
rect -1506 12878 -1502 12948
rect -1482 12878 -1478 12948
rect -1458 12878 -1454 12948
rect -1434 12878 -1430 12948
rect -1410 12878 -1406 12948
rect -1386 12878 -1382 12948
rect -1362 12878 -1358 12948
rect -1338 12878 -1334 12948
rect -1314 12878 -1310 12948
rect -1290 12878 -1286 12948
rect -1266 12878 -1262 12948
rect -1242 12878 -1238 12948
rect -1218 12878 -1214 12948
rect -1194 12878 -1190 12948
rect -1170 12878 -1166 12948
rect -1146 12878 -1142 12948
rect -1122 12878 -1118 12948
rect -1098 12878 -1094 12948
rect -1074 12878 -1070 12948
rect -1061 12941 -1056 12948
rect -1050 12941 -1046 12948
rect -1051 12927 -1046 12941
rect -1061 12917 -1056 12927
rect -1051 12903 -1046 12917
rect -1050 12878 -1046 12903
rect -1026 12878 -1022 12971
rect -1002 12878 -998 12996
rect -978 12878 -974 12996
rect -954 12878 -950 12996
rect -930 12878 -926 12996
rect -906 12878 -902 12996
rect -882 12878 -878 12996
rect -858 12878 -854 12996
rect -834 12878 -830 12996
rect -810 12878 -806 12996
rect -786 12878 -782 12996
rect -762 12878 -758 12996
rect -738 12878 -734 12996
rect -714 12878 -710 12996
rect -690 12878 -686 12996
rect -666 12878 -662 12996
rect -642 12878 -638 12996
rect -618 12878 -614 12996
rect -594 12878 -590 12996
rect -581 12917 -576 12927
rect -570 12917 -566 12996
rect -571 12903 -566 12917
rect -581 12902 -547 12903
rect -546 12902 -542 12996
rect -522 12902 -518 12996
rect -498 12902 -494 12996
rect -474 12902 -470 12996
rect -450 12902 -446 12996
rect -426 12902 -422 12996
rect -402 12902 -398 12996
rect -378 12902 -374 12996
rect -354 12902 -350 12996
rect -330 12902 -326 12996
rect -306 12902 -302 12996
rect -282 12902 -278 12996
rect -258 12902 -254 12996
rect -234 12902 -230 12996
rect -210 12902 -206 12996
rect -186 12902 -182 12996
rect -162 12902 -158 12996
rect -138 12902 -134 12996
rect -114 12902 -110 12996
rect -90 12902 -86 12996
rect -66 12902 -62 12996
rect -42 12902 -38 12996
rect -18 12902 -14 12996
rect 6 12902 10 12996
rect 30 12902 34 12996
rect 54 12902 58 12996
rect 78 12902 82 12996
rect 102 12902 106 12996
rect 126 12902 130 12996
rect 150 12902 154 12996
rect 174 12902 178 12996
rect 198 12902 202 12996
rect 222 12902 226 12996
rect 246 12902 250 12996
rect 270 12902 274 12996
rect 294 12902 298 12996
rect 318 12902 322 12996
rect 342 12902 346 12996
rect 366 12902 370 12996
rect 390 12902 394 12996
rect 414 12902 418 12996
rect 438 12902 442 12996
rect 462 12902 466 12996
rect 486 12902 490 12996
rect 510 12902 514 12996
rect 534 12902 538 12996
rect 558 12902 562 12996
rect 582 12902 586 12996
rect 606 12902 610 12996
rect 630 12902 634 12996
rect 654 12902 658 12996
rect 661 12995 675 12996
rect 678 12974 685 13019
rect 702 12974 706 13044
rect 726 12974 730 13044
rect 750 12974 754 13044
rect 774 12974 778 13044
rect 798 12974 802 13044
rect 822 12974 826 13044
rect 846 12974 850 13044
rect 870 12974 874 13044
rect 894 12974 898 13044
rect 918 12974 922 13044
rect 942 12974 946 13044
rect 966 12974 970 13044
rect 990 12974 994 13044
rect 1014 12974 1018 13044
rect 1038 12974 1042 13044
rect 1062 12974 1066 13044
rect 1086 12974 1090 13044
rect 1110 12974 1114 13044
rect 1134 12974 1138 13044
rect 1158 12974 1162 13044
rect 1182 12974 1186 13044
rect 1206 12974 1210 13044
rect 1230 12974 1234 13044
rect 1254 12974 1258 13044
rect 1278 12974 1282 13044
rect 1302 12974 1306 13044
rect 1326 12974 1330 13044
rect 1350 12974 1354 13044
rect 1374 12974 1378 13044
rect 1398 12974 1402 13044
rect 1422 12974 1426 13044
rect 1446 12974 1450 13044
rect 1470 12974 1474 13044
rect 1494 12974 1498 13044
rect 1518 12974 1522 13044
rect 1542 12974 1546 13044
rect 1566 12974 1570 13044
rect 1590 12974 1594 13044
rect 1614 12974 1618 13044
rect 1638 12974 1642 13044
rect 1662 12974 1666 13044
rect 1686 12974 1690 13044
rect 1710 12974 1714 13044
rect 1734 12975 1738 13044
rect 1723 12974 1757 12975
rect 661 12972 1757 12974
rect 661 12971 675 12972
rect 678 12971 685 12972
rect 678 12902 682 12971
rect 702 12902 706 12972
rect 726 12902 730 12972
rect 750 12902 754 12972
rect 774 12902 778 12972
rect 798 12902 802 12972
rect 822 12902 826 12972
rect 846 12902 850 12972
rect 870 12902 874 12972
rect 894 12902 898 12972
rect 918 12902 922 12972
rect 942 12902 946 12972
rect 966 12902 970 12972
rect 990 12902 994 12972
rect 1014 12902 1018 12972
rect 1038 12902 1042 12972
rect 1062 12902 1066 12972
rect 1086 12902 1090 12972
rect 1110 12902 1114 12972
rect 1134 12902 1138 12972
rect 1158 12902 1162 12972
rect 1182 12902 1186 12972
rect 1206 12902 1210 12972
rect 1230 12902 1234 12972
rect 1254 12902 1258 12972
rect 1278 12902 1282 12972
rect 1302 12902 1306 12972
rect 1326 12902 1330 12972
rect 1350 12902 1354 12972
rect 1374 12902 1378 12972
rect 1398 12902 1402 12972
rect 1422 12902 1426 12972
rect 1446 12902 1450 12972
rect 1470 12902 1474 12972
rect 1494 12902 1498 12972
rect 1518 12902 1522 12972
rect 1542 12902 1546 12972
rect 1566 12902 1570 12972
rect 1590 12902 1594 12972
rect 1614 12902 1618 12972
rect 1638 12902 1642 12972
rect 1662 12902 1666 12972
rect 1686 12902 1690 12972
rect 1710 12902 1714 12972
rect 1723 12965 1728 12972
rect 1734 12965 1738 12972
rect 1733 12951 1738 12965
rect 1723 12950 1757 12951
rect 1758 12950 1762 13044
rect 1782 12950 1786 13044
rect 1806 12950 1810 13044
rect 1830 12950 1834 13044
rect 1854 12950 1858 13044
rect 1878 12950 1882 13044
rect 1902 12950 1906 13044
rect 1926 12950 1930 13044
rect 1950 12950 1954 13044
rect 1974 12950 1978 13044
rect 1998 12950 2002 13044
rect 2022 12950 2026 13044
rect 2046 12950 2050 13044
rect 2070 12950 2074 13044
rect 2094 12950 2098 13044
rect 2118 12950 2122 13044
rect 2142 12950 2146 13044
rect 2166 12950 2170 13044
rect 2190 12950 2194 13044
rect 2214 12950 2218 13044
rect 2238 12950 2242 13044
rect 2262 12950 2266 13044
rect 2286 12950 2290 13044
rect 2310 12950 2314 13044
rect 2334 12950 2338 13044
rect 2358 12950 2362 13044
rect 2382 12950 2386 13044
rect 2406 12950 2410 13044
rect 2430 12950 2434 13044
rect 2454 12950 2458 13044
rect 2478 12950 2482 13044
rect 2502 12950 2506 13044
rect 2526 12950 2530 13044
rect 2550 12950 2554 13044
rect 2574 12950 2578 13044
rect 2598 12950 2602 13044
rect 2622 12950 2626 13044
rect 2646 12950 2650 13044
rect 2670 12950 2674 13044
rect 2694 12950 2698 13044
rect 2718 12950 2722 13044
rect 2742 12950 2746 13044
rect 2766 12950 2770 13044
rect 2790 12950 2794 13044
rect 2814 12950 2818 13044
rect 2838 12950 2842 13044
rect 2862 12950 2866 13044
rect 2886 12950 2890 13044
rect 2910 12950 2914 13044
rect 2934 12950 2938 13044
rect 2958 12950 2962 13044
rect 2982 12950 2986 13044
rect 3006 12950 3010 13044
rect 3030 12950 3034 13044
rect 3054 12950 3058 13044
rect 3078 12950 3082 13044
rect 3102 12950 3106 13044
rect 3126 12950 3130 13044
rect 3139 13037 3144 13044
rect 3150 13037 3154 13044
rect 3149 13023 3154 13037
rect 3150 12950 3154 13023
rect 3174 12971 3178 13068
rect 1723 12948 3171 12950
rect 1723 12941 1728 12948
rect 1733 12927 1738 12941
rect 1734 12902 1738 12927
rect 1758 12902 1762 12948
rect 1782 12902 1786 12948
rect 1806 12902 1810 12948
rect 1830 12902 1834 12948
rect 1854 12902 1858 12948
rect 1878 12902 1882 12948
rect 1902 12902 1906 12948
rect 1926 12902 1930 12948
rect 1950 12902 1954 12948
rect 1974 12902 1978 12948
rect 1998 12902 2002 12948
rect 2022 12902 2026 12948
rect 2046 12902 2050 12948
rect 2070 12902 2074 12948
rect 2094 12902 2098 12948
rect 2118 12902 2122 12948
rect 2142 12902 2146 12948
rect 2166 12902 2170 12948
rect 2190 12902 2194 12948
rect 2214 12902 2218 12948
rect 2238 12902 2242 12948
rect 2262 12902 2266 12948
rect 2286 12902 2290 12948
rect 2310 12902 2314 12948
rect 2334 12902 2338 12948
rect 2358 12902 2362 12948
rect 2382 12902 2386 12948
rect 2406 12902 2410 12948
rect 2430 12902 2434 12948
rect 2454 12902 2458 12948
rect 2478 12902 2482 12948
rect 2502 12902 2506 12948
rect 2526 12902 2530 12948
rect 2550 12902 2554 12948
rect 2574 12902 2578 12948
rect 2598 12902 2602 12948
rect 2622 12902 2626 12948
rect 2646 12902 2650 12948
rect 2670 12902 2674 12948
rect 2694 12902 2698 12948
rect 2718 12902 2722 12948
rect 2742 12902 2746 12948
rect 2766 12902 2770 12948
rect 2790 12902 2794 12948
rect 2814 12902 2818 12948
rect 2838 12902 2842 12948
rect 2862 12902 2866 12948
rect 2886 12902 2890 12948
rect 2910 12902 2914 12948
rect 2934 12902 2938 12948
rect 2958 12902 2962 12948
rect 2982 12902 2986 12948
rect 3006 12902 3010 12948
rect 3030 12902 3034 12948
rect 3054 12902 3058 12948
rect 3078 12902 3082 12948
rect 3102 12902 3106 12948
rect 3126 12902 3130 12948
rect 3150 12902 3154 12948
rect 3157 12947 3171 12948
rect 3174 12947 3181 12971
rect 3174 12902 3178 12947
rect 3198 12902 3202 13068
rect 3222 12902 3226 13068
rect 3246 12902 3250 13068
rect 3270 12902 3274 13068
rect 3294 12902 3298 13068
rect 3318 12902 3322 13068
rect 3342 12902 3346 13068
rect 3366 12902 3370 13068
rect 3390 12902 3394 13068
rect 3414 12902 3418 13068
rect 3438 12902 3442 13068
rect 3462 12902 3466 13068
rect 3486 12903 3490 13068
rect 3499 13061 3504 13068
rect 3510 13061 3514 13068
rect 3509 13047 3514 13061
rect 3523 13057 3531 13061
rect 3517 13047 3523 13057
rect 3499 12989 3504 12999
rect 3509 12975 3514 12989
rect 3523 12985 3531 12989
rect 3517 12975 3523 12985
rect 3499 12941 3504 12951
rect 3510 12941 3514 12975
rect 3509 12927 3514 12941
rect 3475 12902 3509 12903
rect -581 12900 3509 12902
rect -581 12893 -576 12900
rect -571 12879 -566 12893
rect -570 12878 -566 12879
rect -546 12878 -542 12900
rect -522 12878 -518 12900
rect -498 12878 -494 12900
rect -474 12878 -470 12900
rect -450 12878 -446 12900
rect -426 12878 -422 12900
rect -402 12878 -398 12900
rect -378 12878 -374 12900
rect -354 12878 -350 12900
rect -330 12878 -326 12900
rect -306 12878 -302 12900
rect -282 12878 -278 12900
rect -258 12878 -254 12900
rect -234 12878 -230 12900
rect -210 12878 -206 12900
rect -186 12878 -182 12900
rect -162 12878 -158 12900
rect -138 12878 -134 12900
rect -114 12878 -110 12900
rect -90 12878 -86 12900
rect -66 12878 -62 12900
rect -42 12878 -38 12900
rect -18 12878 -14 12900
rect 6 12878 10 12900
rect 30 12878 34 12900
rect 54 12878 58 12900
rect 78 12878 82 12900
rect 102 12878 106 12900
rect 126 12878 130 12900
rect 150 12878 154 12900
rect 174 12878 178 12900
rect 198 12878 202 12900
rect 222 12878 226 12900
rect 246 12878 250 12900
rect 270 12878 274 12900
rect 294 12878 298 12900
rect 318 12878 322 12900
rect 342 12878 346 12900
rect 366 12878 370 12900
rect 390 12878 394 12900
rect 414 12878 418 12900
rect 438 12878 442 12900
rect 462 12878 466 12900
rect 486 12878 490 12900
rect 510 12878 514 12900
rect 534 12878 538 12900
rect 558 12878 562 12900
rect 582 12878 586 12900
rect 606 12878 610 12900
rect 630 12878 634 12900
rect 654 12878 658 12900
rect 678 12878 682 12900
rect 702 12878 706 12900
rect 726 12878 730 12900
rect 750 12878 754 12900
rect 774 12878 778 12900
rect 798 12878 802 12900
rect 822 12878 826 12900
rect 846 12878 850 12900
rect 870 12878 874 12900
rect 894 12878 898 12900
rect 918 12878 922 12900
rect 942 12878 946 12900
rect 966 12878 970 12900
rect 990 12878 994 12900
rect 1014 12878 1018 12900
rect 1038 12878 1042 12900
rect 1062 12878 1066 12900
rect 1086 12878 1090 12900
rect 1110 12878 1114 12900
rect 1134 12878 1138 12900
rect 1158 12878 1162 12900
rect 1182 12878 1186 12900
rect 1206 12878 1210 12900
rect 1230 12878 1234 12900
rect 1254 12878 1258 12900
rect 1278 12878 1282 12900
rect 1302 12878 1306 12900
rect 1326 12878 1330 12900
rect 1350 12878 1354 12900
rect 1374 12878 1378 12900
rect 1398 12878 1402 12900
rect 1422 12878 1426 12900
rect 1446 12878 1450 12900
rect 1470 12878 1474 12900
rect 1494 12878 1498 12900
rect 1518 12878 1522 12900
rect 1542 12878 1546 12900
rect 1566 12878 1570 12900
rect 1590 12878 1594 12900
rect 1614 12878 1618 12900
rect 1638 12878 1642 12900
rect 1662 12878 1666 12900
rect 1686 12878 1690 12900
rect 1710 12878 1714 12900
rect 1734 12878 1738 12900
rect 1758 12899 1762 12900
rect -2393 12876 1755 12878
rect -2371 12854 -2366 12876
rect -2348 12854 -2343 12876
rect -2325 12870 -2317 12876
rect -2325 12854 -2320 12870
rect -2309 12858 -2301 12870
rect -2068 12859 -2038 12866
rect -2317 12854 -2309 12858
rect -2000 12856 -1992 12876
rect -1844 12868 -1794 12876
rect -1671 12870 -1663 12876
rect -1852 12859 -1804 12866
rect -1655 12858 -1647 12870
rect -2025 12855 -1991 12856
rect -2025 12854 -1975 12855
rect -1844 12854 -1804 12857
rect -1663 12854 -1655 12858
rect -1642 12854 -1637 12876
rect -1619 12854 -1614 12876
rect -1530 12854 -1526 12876
rect -1506 12854 -1502 12876
rect -1482 12854 -1478 12876
rect -1458 12854 -1454 12876
rect -1434 12854 -1430 12876
rect -1410 12854 -1406 12876
rect -1386 12854 -1382 12876
rect -1362 12854 -1358 12876
rect -1338 12854 -1334 12876
rect -1314 12854 -1310 12876
rect -1290 12854 -1286 12876
rect -1266 12854 -1262 12876
rect -1242 12854 -1238 12876
rect -1218 12854 -1214 12876
rect -1194 12854 -1190 12876
rect -1170 12854 -1166 12876
rect -1146 12854 -1142 12876
rect -1122 12854 -1118 12876
rect -1098 12854 -1094 12876
rect -1074 12854 -1070 12876
rect -1050 12855 -1046 12876
rect -1026 12875 -1022 12876
rect -1061 12854 -1029 12855
rect -2393 12852 -1029 12854
rect -2371 12830 -2366 12852
rect -2348 12830 -2343 12852
rect -2325 12842 -2317 12852
rect -2060 12842 -2020 12849
rect -2004 12844 -2001 12849
rect -2015 12842 -2001 12844
rect -2000 12842 -1992 12852
rect -1972 12850 -1958 12852
rect -1844 12851 -1804 12852
rect -1862 12849 -1796 12850
rect -1985 12847 -1796 12849
rect -1985 12842 -1852 12847
rect -2325 12830 -2320 12842
rect -2309 12830 -2301 12842
rect -2068 12832 -2060 12839
rect -2015 12832 -1990 12842
rect -1844 12841 -1796 12847
rect -1671 12842 -1663 12852
rect -1852 12832 -1804 12839
rect -2020 12830 -2004 12832
rect -2000 12830 -1992 12832
rect -1976 12830 -1940 12831
rect -1655 12830 -1647 12842
rect -1642 12830 -1637 12852
rect -1619 12830 -1614 12852
rect -1530 12830 -1526 12852
rect -1506 12830 -1502 12852
rect -1482 12830 -1478 12852
rect -1458 12830 -1454 12852
rect -1434 12830 -1430 12852
rect -1410 12830 -1406 12852
rect -1386 12830 -1382 12852
rect -1362 12830 -1358 12852
rect -1338 12830 -1334 12852
rect -1314 12830 -1310 12852
rect -1290 12830 -1286 12852
rect -1266 12830 -1262 12852
rect -1242 12830 -1238 12852
rect -1218 12830 -1214 12852
rect -1194 12830 -1190 12852
rect -1170 12830 -1166 12852
rect -1146 12830 -1142 12852
rect -1122 12830 -1118 12852
rect -1098 12830 -1094 12852
rect -1074 12830 -1070 12852
rect -1061 12845 -1056 12852
rect -1050 12845 -1046 12852
rect -1043 12851 -1029 12852
rect -1051 12831 -1046 12845
rect -1037 12841 -1029 12845
rect -1043 12831 -1037 12841
rect -1050 12830 -1046 12831
rect -1026 12830 -1019 12875
rect -1002 12830 -998 12876
rect -978 12830 -974 12876
rect -954 12830 -950 12876
rect -930 12830 -926 12876
rect -906 12830 -902 12876
rect -882 12830 -878 12876
rect -858 12830 -854 12876
rect -834 12831 -830 12876
rect -845 12830 -811 12831
rect -2393 12828 -811 12830
rect -2371 12734 -2366 12828
rect -2348 12734 -2343 12828
rect -2325 12826 -2320 12828
rect -2317 12826 -2309 12828
rect -2325 12814 -2317 12826
rect -2060 12815 -2030 12822
rect -2325 12794 -2320 12814
rect -2325 12786 -2317 12794
rect -2060 12788 -2030 12791
rect -2325 12734 -2320 12786
rect -2317 12778 -2309 12786
rect -2060 12775 -2038 12786
rect -2033 12779 -2030 12788
rect -2028 12784 -2027 12788
rect -2068 12770 -2038 12773
rect -2309 12738 -2301 12746
rect -2317 12734 -2309 12738
rect -2000 12734 -1992 12828
rect -1844 12824 -1804 12828
rect -1663 12826 -1655 12828
rect -1844 12814 -1794 12823
rect -1671 12814 -1663 12826
rect -1912 12803 -1884 12805
rect -1852 12797 -1804 12801
rect -1844 12788 -1796 12791
rect -1671 12786 -1663 12794
rect -1844 12775 -1804 12786
rect -1663 12778 -1655 12786
rect -1852 12770 -1680 12774
rect -1655 12738 -1647 12746
rect -1663 12734 -1655 12738
rect -1642 12734 -1637 12828
rect -1619 12734 -1614 12828
rect -1541 12797 -1536 12807
rect -1530 12797 -1526 12828
rect -1531 12783 -1526 12797
rect -1541 12782 -1507 12783
rect -1506 12782 -1502 12828
rect -1482 12782 -1478 12828
rect -1458 12782 -1454 12828
rect -1434 12782 -1430 12828
rect -1410 12782 -1406 12828
rect -1386 12782 -1382 12828
rect -1362 12782 -1358 12828
rect -1338 12782 -1334 12828
rect -1314 12782 -1310 12828
rect -1290 12782 -1286 12828
rect -1266 12782 -1262 12828
rect -1242 12782 -1238 12828
rect -1218 12782 -1214 12828
rect -1194 12782 -1190 12828
rect -1170 12782 -1166 12828
rect -1146 12782 -1142 12828
rect -1122 12782 -1118 12828
rect -1098 12782 -1094 12828
rect -1074 12782 -1070 12828
rect -1050 12782 -1046 12828
rect -1043 12827 -1029 12828
rect -1026 12827 -1019 12828
rect -1026 12782 -1022 12827
rect -1002 12782 -998 12828
rect -978 12782 -974 12828
rect -954 12782 -950 12828
rect -930 12782 -926 12828
rect -906 12782 -902 12828
rect -882 12782 -878 12828
rect -858 12782 -854 12828
rect -845 12821 -840 12828
rect -834 12821 -830 12828
rect -835 12807 -830 12821
rect -845 12797 -840 12807
rect -835 12783 -830 12797
rect -834 12782 -830 12783
rect -810 12782 -806 12876
rect -786 12782 -782 12876
rect -762 12782 -758 12876
rect -738 12782 -734 12876
rect -714 12782 -710 12876
rect -690 12782 -686 12876
rect -666 12782 -662 12876
rect -642 12782 -638 12876
rect -618 12782 -614 12876
rect -594 12782 -590 12876
rect -570 12782 -566 12876
rect -546 12851 -542 12876
rect -546 12806 -539 12851
rect -522 12806 -518 12876
rect -498 12806 -494 12876
rect -474 12806 -470 12876
rect -450 12806 -446 12876
rect -426 12806 -422 12876
rect -402 12806 -398 12876
rect -378 12806 -374 12876
rect -354 12806 -350 12876
rect -330 12806 -326 12876
rect -306 12806 -302 12876
rect -282 12806 -278 12876
rect -258 12806 -254 12876
rect -234 12806 -230 12876
rect -210 12806 -206 12876
rect -186 12806 -182 12876
rect -162 12806 -158 12876
rect -138 12806 -134 12876
rect -114 12806 -110 12876
rect -90 12806 -86 12876
rect -66 12806 -62 12876
rect -42 12806 -38 12876
rect -18 12806 -14 12876
rect 6 12806 10 12876
rect 30 12806 34 12876
rect 54 12806 58 12876
rect 78 12806 82 12876
rect 102 12806 106 12876
rect 126 12806 130 12876
rect 150 12806 154 12876
rect 174 12806 178 12876
rect 198 12806 202 12876
rect 222 12806 226 12876
rect 246 12806 250 12876
rect 270 12806 274 12876
rect 294 12806 298 12876
rect 318 12806 322 12876
rect 342 12806 346 12876
rect 366 12806 370 12876
rect 390 12806 394 12876
rect 414 12806 418 12876
rect 438 12806 442 12876
rect 462 12806 466 12876
rect 486 12806 490 12876
rect 510 12806 514 12876
rect 534 12806 538 12876
rect 558 12806 562 12876
rect 582 12806 586 12876
rect 606 12806 610 12876
rect 630 12806 634 12876
rect 654 12806 658 12876
rect 678 12806 682 12876
rect 702 12806 706 12876
rect 726 12806 730 12876
rect 750 12806 754 12876
rect 774 12806 778 12876
rect 798 12806 802 12876
rect 822 12806 826 12876
rect 846 12806 850 12876
rect 870 12806 874 12876
rect 894 12806 898 12876
rect 918 12806 922 12876
rect 942 12806 946 12876
rect 966 12806 970 12876
rect 990 12806 994 12876
rect 1014 12806 1018 12876
rect 1038 12806 1042 12876
rect 1062 12806 1066 12876
rect 1086 12806 1090 12876
rect 1110 12806 1114 12876
rect 1134 12806 1138 12876
rect 1158 12806 1162 12876
rect 1182 12806 1186 12876
rect 1206 12806 1210 12876
rect 1230 12806 1234 12876
rect 1254 12806 1258 12876
rect 1278 12806 1282 12876
rect 1302 12806 1306 12876
rect 1326 12806 1330 12876
rect 1350 12806 1354 12876
rect 1374 12806 1378 12876
rect 1398 12806 1402 12876
rect 1422 12806 1426 12876
rect 1446 12806 1450 12876
rect 1470 12806 1474 12876
rect 1494 12806 1498 12876
rect 1518 12806 1522 12876
rect 1542 12806 1546 12876
rect 1566 12806 1570 12876
rect 1590 12806 1594 12876
rect 1614 12806 1618 12876
rect 1638 12806 1642 12876
rect 1662 12806 1666 12876
rect 1686 12806 1690 12876
rect 1710 12806 1714 12876
rect 1734 12806 1738 12876
rect 1741 12875 1755 12876
rect 1758 12851 1765 12899
rect 1758 12806 1762 12851
rect 1782 12806 1786 12900
rect 1806 12806 1810 12900
rect 1830 12806 1834 12900
rect 1854 12806 1858 12900
rect 1878 12806 1882 12900
rect 1902 12806 1906 12900
rect 1926 12806 1930 12900
rect 1950 12806 1954 12900
rect 1974 12806 1978 12900
rect 1998 12806 2002 12900
rect 2022 12806 2026 12900
rect 2046 12806 2050 12900
rect 2070 12806 2074 12900
rect 2094 12806 2098 12900
rect 2118 12806 2122 12900
rect 2142 12806 2146 12900
rect 2166 12806 2170 12900
rect 2190 12806 2194 12900
rect 2214 12806 2218 12900
rect 2238 12806 2242 12900
rect 2262 12806 2266 12900
rect 2286 12806 2290 12900
rect 2310 12806 2314 12900
rect 2334 12806 2338 12900
rect 2358 12806 2362 12900
rect 2382 12806 2386 12900
rect 2406 12806 2410 12900
rect 2430 12806 2434 12900
rect 2454 12806 2458 12900
rect 2478 12806 2482 12900
rect 2502 12806 2506 12900
rect 2526 12806 2530 12900
rect 2550 12806 2554 12900
rect 2574 12806 2578 12900
rect 2598 12806 2602 12900
rect 2622 12806 2626 12900
rect 2646 12806 2650 12900
rect 2670 12806 2674 12900
rect 2694 12806 2698 12900
rect 2718 12806 2722 12900
rect 2742 12806 2746 12900
rect 2766 12806 2770 12900
rect 2790 12806 2794 12900
rect 2814 12806 2818 12900
rect 2838 12806 2842 12900
rect 2862 12806 2866 12900
rect 2886 12806 2890 12900
rect 2910 12806 2914 12900
rect 2934 12806 2938 12900
rect 2958 12806 2962 12900
rect 2982 12806 2986 12900
rect 3006 12806 3010 12900
rect 3030 12806 3034 12900
rect 3054 12806 3058 12900
rect 3078 12806 3082 12900
rect 3102 12806 3106 12900
rect 3126 12806 3130 12900
rect 3150 12806 3154 12900
rect 3174 12806 3178 12900
rect 3198 12806 3202 12900
rect 3222 12806 3226 12900
rect 3246 12806 3250 12900
rect 3270 12806 3274 12900
rect 3294 12806 3298 12900
rect 3318 12806 3322 12900
rect 3342 12806 3346 12900
rect 3366 12806 3370 12900
rect 3390 12806 3394 12900
rect 3414 12806 3418 12900
rect 3438 12806 3442 12900
rect 3462 12806 3466 12900
rect 3475 12893 3480 12900
rect 3486 12893 3490 12900
rect 3485 12879 3490 12893
rect 3475 12869 3480 12879
rect 3485 12855 3490 12869
rect 3486 12807 3490 12855
rect 3475 12806 3507 12807
rect -563 12804 3507 12806
rect -563 12803 -549 12804
rect -546 12803 -539 12804
rect -546 12782 -542 12803
rect -522 12782 -518 12804
rect -498 12782 -494 12804
rect -474 12782 -470 12804
rect -450 12782 -446 12804
rect -426 12782 -422 12804
rect -402 12782 -398 12804
rect -378 12782 -374 12804
rect -354 12782 -350 12804
rect -330 12782 -326 12804
rect -306 12782 -302 12804
rect -282 12782 -278 12804
rect -258 12782 -254 12804
rect -234 12782 -230 12804
rect -210 12782 -206 12804
rect -186 12782 -182 12804
rect -162 12782 -158 12804
rect -138 12782 -134 12804
rect -114 12782 -110 12804
rect -90 12782 -86 12804
rect -66 12782 -62 12804
rect -42 12782 -38 12804
rect -18 12782 -14 12804
rect 6 12782 10 12804
rect 30 12782 34 12804
rect 54 12782 58 12804
rect 78 12782 82 12804
rect 102 12782 106 12804
rect 126 12782 130 12804
rect 150 12782 154 12804
rect 174 12782 178 12804
rect 198 12782 202 12804
rect 222 12782 226 12804
rect 246 12782 250 12804
rect 270 12782 274 12804
rect 294 12782 298 12804
rect 318 12782 322 12804
rect 342 12782 346 12804
rect 366 12782 370 12804
rect 390 12782 394 12804
rect 414 12782 418 12804
rect 438 12782 442 12804
rect 462 12782 466 12804
rect 486 12782 490 12804
rect 510 12782 514 12804
rect 534 12782 538 12804
rect 558 12782 562 12804
rect 582 12782 586 12804
rect 606 12782 610 12804
rect 630 12782 634 12804
rect 654 12782 658 12804
rect 678 12782 682 12804
rect 702 12782 706 12804
rect 726 12782 730 12804
rect 750 12782 754 12804
rect 774 12782 778 12804
rect 798 12782 802 12804
rect 822 12782 826 12804
rect 846 12782 850 12804
rect 870 12782 874 12804
rect 894 12782 898 12804
rect 918 12782 922 12804
rect 942 12782 946 12804
rect 966 12782 970 12804
rect 990 12782 994 12804
rect 1014 12782 1018 12804
rect 1038 12782 1042 12804
rect 1062 12782 1066 12804
rect 1086 12782 1090 12804
rect 1110 12782 1114 12804
rect 1134 12782 1138 12804
rect 1158 12782 1162 12804
rect 1182 12782 1186 12804
rect 1206 12782 1210 12804
rect 1230 12782 1234 12804
rect 1254 12782 1258 12804
rect 1278 12782 1282 12804
rect 1302 12782 1306 12804
rect 1326 12782 1330 12804
rect 1350 12782 1354 12804
rect 1374 12782 1378 12804
rect 1398 12782 1402 12804
rect 1422 12782 1426 12804
rect 1446 12782 1450 12804
rect 1470 12782 1474 12804
rect 1494 12782 1498 12804
rect 1518 12782 1522 12804
rect 1542 12782 1546 12804
rect 1566 12782 1570 12804
rect 1590 12782 1594 12804
rect 1614 12782 1618 12804
rect 1638 12782 1642 12804
rect 1662 12782 1666 12804
rect 1686 12782 1690 12804
rect 1710 12782 1714 12804
rect 1734 12782 1738 12804
rect 1758 12782 1762 12804
rect 1782 12782 1786 12804
rect 1806 12782 1810 12804
rect 1830 12782 1834 12804
rect 1854 12782 1858 12804
rect 1878 12782 1882 12804
rect 1902 12782 1906 12804
rect 1926 12782 1930 12804
rect 1950 12782 1954 12804
rect 1974 12782 1978 12804
rect 1998 12782 2002 12804
rect 2022 12782 2026 12804
rect 2046 12782 2050 12804
rect 2070 12782 2074 12804
rect 2094 12782 2098 12804
rect 2118 12782 2122 12804
rect 2142 12782 2146 12804
rect 2166 12782 2170 12804
rect 2190 12782 2194 12804
rect 2214 12782 2218 12804
rect 2238 12782 2242 12804
rect 2262 12782 2266 12804
rect 2286 12782 2290 12804
rect 2310 12782 2314 12804
rect 2334 12782 2338 12804
rect 2358 12782 2362 12804
rect 2382 12782 2386 12804
rect 2406 12782 2410 12804
rect 2430 12782 2434 12804
rect 2454 12782 2458 12804
rect 2478 12782 2482 12804
rect 2502 12782 2506 12804
rect 2526 12782 2530 12804
rect 2550 12782 2554 12804
rect 2574 12782 2578 12804
rect 2598 12782 2602 12804
rect 2622 12782 2626 12804
rect 2646 12782 2650 12804
rect 2670 12782 2674 12804
rect 2694 12782 2698 12804
rect 2718 12782 2722 12804
rect 2742 12782 2746 12804
rect 2766 12782 2770 12804
rect 2790 12782 2794 12804
rect 2814 12782 2818 12804
rect 2838 12782 2842 12804
rect 2862 12782 2866 12804
rect 2886 12782 2890 12804
rect 2910 12782 2914 12804
rect 2934 12782 2938 12804
rect 2958 12782 2962 12804
rect 2982 12782 2986 12804
rect 3006 12782 3010 12804
rect 3030 12782 3034 12804
rect 3054 12782 3058 12804
rect 3078 12782 3082 12804
rect 3102 12782 3106 12804
rect 3126 12782 3130 12804
rect 3150 12782 3154 12804
rect 3174 12782 3178 12804
rect 3198 12782 3202 12804
rect 3222 12782 3226 12804
rect 3246 12782 3250 12804
rect 3270 12782 3274 12804
rect 3294 12782 3298 12804
rect 3318 12782 3322 12804
rect 3342 12782 3346 12804
rect 3366 12782 3370 12804
rect 3390 12782 3394 12804
rect 3414 12782 3418 12804
rect 3438 12782 3442 12804
rect 3462 12783 3466 12804
rect 3475 12797 3480 12804
rect 3486 12797 3490 12804
rect 3493 12803 3507 12804
rect 3485 12783 3490 12797
rect 3499 12793 3507 12797
rect 3493 12783 3499 12793
rect 3451 12782 3485 12783
rect -1541 12780 3485 12782
rect -1541 12773 -1536 12780
rect -1531 12759 -1526 12773
rect -1530 12734 -1526 12759
rect -1506 12734 -1502 12780
rect -1482 12734 -1478 12780
rect -1458 12734 -1454 12780
rect -1434 12734 -1430 12780
rect -1410 12734 -1406 12780
rect -1386 12734 -1382 12780
rect -1362 12734 -1358 12780
rect -1338 12734 -1334 12780
rect -1314 12734 -1310 12780
rect -1290 12734 -1286 12780
rect -1266 12734 -1262 12780
rect -1242 12734 -1238 12780
rect -1218 12734 -1214 12780
rect -1194 12734 -1190 12780
rect -1170 12734 -1166 12780
rect -1146 12734 -1142 12780
rect -1122 12734 -1118 12780
rect -1098 12735 -1094 12780
rect -1109 12734 -1075 12735
rect -2393 12732 -2020 12734
rect -2012 12732 -1075 12734
rect -2371 12638 -2366 12732
rect -2348 12638 -2343 12732
rect -2325 12670 -2320 12732
rect -2317 12730 -2309 12732
rect -2062 12719 -2061 12720
rect -2060 12719 -2049 12732
rect -2309 12710 -2301 12718
rect -2068 12712 -2061 12719
rect -2020 12712 -2012 12724
rect -2317 12702 -2309 12710
rect -2124 12703 -2108 12705
rect -2060 12703 -2049 12712
rect -2020 12710 -2004 12712
rect -2000 12710 -1992 12732
rect -1972 12730 -1958 12732
rect -1663 12730 -1655 12732
rect -1958 12729 -1942 12730
rect -1980 12712 -1932 12719
rect -1655 12710 -1647 12718
rect -2292 12702 -2049 12703
rect -2036 12702 -2030 12710
rect -2020 12708 -1992 12710
rect -2292 12695 -2030 12702
rect -2292 12694 -2049 12695
rect -2031 12694 -2030 12695
rect -2026 12694 -2020 12700
rect -2325 12662 -2317 12670
rect -2325 12642 -2320 12662
rect -2317 12654 -2309 12662
rect -2325 12638 -2317 12642
rect -2095 12640 -2083 12644
rect -2000 12641 -1992 12708
rect -1844 12694 -1680 12703
rect -1663 12702 -1655 12710
rect -1671 12662 -1663 12670
rect -1663 12654 -1655 12662
rect -2119 12638 -2069 12640
rect -2053 12638 -1972 12641
rect -1926 12638 -1892 12641
rect -1671 12638 -1663 12642
rect -1642 12638 -1637 12732
rect -1619 12638 -1614 12732
rect -1530 12638 -1526 12732
rect -1506 12731 -1502 12732
rect -1506 12686 -1499 12731
rect -1482 12686 -1478 12732
rect -1458 12686 -1454 12732
rect -1434 12686 -1430 12732
rect -1410 12686 -1406 12732
rect -1386 12686 -1382 12732
rect -1362 12686 -1358 12732
rect -1338 12686 -1334 12732
rect -1314 12686 -1310 12732
rect -1290 12686 -1286 12732
rect -1266 12686 -1262 12732
rect -1242 12686 -1238 12732
rect -1218 12686 -1214 12732
rect -1194 12686 -1190 12732
rect -1170 12686 -1166 12732
rect -1146 12686 -1142 12732
rect -1122 12686 -1118 12732
rect -1109 12725 -1104 12732
rect -1098 12725 -1094 12732
rect -1099 12711 -1094 12725
rect -1098 12686 -1094 12711
rect -1074 12686 -1070 12780
rect -1050 12686 -1046 12780
rect -1026 12779 -1022 12780
rect -1026 12755 -1019 12779
rect -1026 12686 -1022 12755
rect -1002 12686 -998 12780
rect -978 12687 -974 12780
rect -989 12686 -955 12687
rect -1523 12684 -955 12686
rect -1523 12683 -1509 12684
rect -1506 12683 -1499 12684
rect -1506 12638 -1502 12683
rect -1482 12638 -1478 12684
rect -1458 12638 -1454 12684
rect -1434 12638 -1430 12684
rect -1410 12638 -1406 12684
rect -1386 12638 -1382 12684
rect -1362 12638 -1358 12684
rect -1338 12638 -1334 12684
rect -1314 12638 -1310 12684
rect -1290 12638 -1286 12684
rect -1266 12638 -1262 12684
rect -1242 12638 -1238 12684
rect -1218 12638 -1214 12684
rect -1194 12638 -1190 12684
rect -1170 12638 -1166 12684
rect -1146 12638 -1142 12684
rect -1122 12638 -1118 12684
rect -1098 12638 -1094 12684
rect -1074 12659 -1070 12684
rect -2393 12636 -1077 12638
rect -2371 12590 -2366 12636
rect -2348 12590 -2343 12636
rect -2325 12632 -2317 12636
rect -2325 12614 -2320 12632
rect -2317 12626 -2309 12632
rect -2095 12630 -2083 12636
rect -2053 12634 -1972 12636
rect -2083 12628 -2079 12630
rect -2079 12627 -2067 12628
rect -2079 12626 -2043 12627
rect -2091 12622 -2043 12626
rect -2000 12622 -1992 12634
rect -1671 12632 -1663 12636
rect -1982 12622 -1916 12627
rect -1663 12626 -1655 12632
rect -2091 12621 -2018 12622
rect -2091 12619 -2067 12621
rect -2053 12619 -2018 12621
rect -2002 12621 -1916 12622
rect -2002 12619 -1972 12621
rect -1924 12619 -1916 12621
rect -2079 12617 -2067 12619
rect -2000 12618 -1992 12619
rect -2325 12604 -2317 12614
rect -2112 12613 -2096 12617
rect -2083 12614 -2079 12617
rect -2027 12616 -1992 12618
rect -2109 12612 -2096 12613
rect -2112 12605 -2096 12612
rect -2083 12605 -2053 12612
rect -2018 12608 -2017 12616
rect -2023 12606 -2017 12608
rect -2009 12608 -2002 12611
rect -2009 12606 -2003 12608
rect -2109 12604 -2096 12605
rect -2325 12590 -2320 12604
rect -2317 12598 -2309 12604
rect -2112 12601 -2096 12604
rect -2017 12595 -2003 12606
rect -2017 12594 -2009 12595
rect -2074 12590 -2040 12592
rect -2000 12590 -1992 12616
rect -1972 12605 -1924 12612
rect -1671 12604 -1663 12614
rect -1663 12598 -1655 12604
rect -1642 12590 -1637 12636
rect -1619 12590 -1614 12636
rect -1530 12590 -1526 12636
rect -1506 12590 -1502 12636
rect -1482 12590 -1478 12636
rect -1458 12590 -1454 12636
rect -1434 12590 -1430 12636
rect -1410 12590 -1406 12636
rect -1386 12590 -1382 12636
rect -1362 12590 -1358 12636
rect -1338 12590 -1334 12636
rect -1314 12590 -1310 12636
rect -1290 12590 -1286 12636
rect -1266 12590 -1262 12636
rect -1242 12590 -1238 12636
rect -1218 12590 -1214 12636
rect -1194 12590 -1190 12636
rect -1170 12590 -1166 12636
rect -1146 12590 -1142 12636
rect -1122 12590 -1118 12636
rect -1098 12590 -1094 12636
rect -1091 12635 -1077 12636
rect -1074 12635 -1067 12659
rect -1074 12590 -1070 12635
rect -1050 12590 -1046 12684
rect -1026 12590 -1022 12684
rect -1002 12590 -998 12684
rect -989 12677 -984 12684
rect -978 12677 -974 12684
rect -979 12663 -974 12677
rect -989 12653 -984 12663
rect -979 12639 -974 12653
rect -978 12590 -974 12639
rect -954 12611 -950 12780
rect -2393 12588 -957 12590
rect -2371 12542 -2366 12588
rect -2348 12542 -2343 12588
rect -2325 12586 -2320 12588
rect -2325 12576 -2317 12586
rect -2325 12556 -2320 12576
rect -2317 12570 -2309 12576
rect -2325 12548 -2317 12556
rect -2101 12551 -2071 12554
rect -2325 12542 -2320 12548
rect -2317 12542 -2309 12548
rect -2000 12546 -1992 12588
rect -1671 12576 -1663 12586
rect -1663 12570 -1655 12576
rect -1854 12560 -1680 12564
rect -1846 12551 -1798 12554
rect -2079 12545 -2043 12546
rect -2007 12545 -1991 12546
rect -2079 12544 -2071 12545
rect -2079 12542 -2029 12544
rect -2011 12542 -1991 12545
rect -1846 12543 -1806 12549
rect -1671 12548 -1663 12556
rect -1864 12542 -1796 12543
rect -1663 12542 -1655 12548
rect -1642 12542 -1637 12588
rect -1619 12542 -1614 12588
rect -1530 12542 -1526 12588
rect -1506 12542 -1502 12588
rect -1482 12542 -1478 12588
rect -1458 12542 -1454 12588
rect -1434 12542 -1430 12588
rect -1410 12542 -1406 12588
rect -1386 12542 -1382 12588
rect -1362 12542 -1358 12588
rect -1338 12542 -1334 12588
rect -1314 12542 -1310 12588
rect -1290 12542 -1286 12588
rect -1266 12542 -1262 12588
rect -1242 12542 -1238 12588
rect -1218 12542 -1214 12588
rect -1194 12542 -1190 12588
rect -1170 12542 -1166 12588
rect -1146 12542 -1142 12588
rect -1122 12542 -1118 12588
rect -1098 12542 -1094 12588
rect -1074 12542 -1070 12588
rect -1050 12542 -1046 12588
rect -1026 12542 -1022 12588
rect -1002 12542 -998 12588
rect -978 12542 -974 12588
rect -971 12587 -957 12588
rect -954 12566 -947 12611
rect -930 12566 -926 12780
rect -906 12566 -902 12780
rect -882 12566 -878 12780
rect -858 12566 -854 12780
rect -834 12566 -830 12780
rect -810 12755 -806 12780
rect -810 12707 -803 12755
rect -810 12566 -806 12707
rect -786 12566 -782 12780
rect -762 12566 -758 12780
rect -738 12566 -734 12780
rect -714 12566 -710 12780
rect -690 12566 -686 12780
rect -666 12566 -662 12780
rect -642 12566 -638 12780
rect -618 12566 -614 12780
rect -594 12566 -590 12780
rect -570 12566 -566 12780
rect -546 12566 -542 12780
rect -522 12566 -518 12780
rect -498 12566 -494 12780
rect -474 12566 -470 12780
rect -450 12566 -446 12780
rect -426 12566 -422 12780
rect -402 12566 -398 12780
rect -378 12566 -374 12780
rect -354 12566 -350 12780
rect -330 12566 -326 12780
rect -306 12566 -302 12780
rect -282 12566 -278 12780
rect -258 12566 -254 12780
rect -234 12566 -230 12780
rect -210 12566 -206 12780
rect -186 12566 -182 12780
rect -162 12566 -158 12780
rect -138 12566 -134 12780
rect -114 12566 -110 12780
rect -90 12566 -86 12780
rect -66 12566 -62 12780
rect -42 12566 -38 12780
rect -18 12566 -14 12780
rect 6 12566 10 12780
rect 30 12566 34 12780
rect 54 12566 58 12780
rect 78 12566 82 12780
rect 102 12566 106 12780
rect 126 12566 130 12780
rect 150 12566 154 12780
rect 174 12566 178 12780
rect 198 12566 202 12780
rect 222 12566 226 12780
rect 246 12566 250 12780
rect 270 12566 274 12780
rect 294 12566 298 12780
rect 318 12566 322 12780
rect 342 12566 346 12780
rect 366 12566 370 12780
rect 390 12566 394 12780
rect 414 12566 418 12780
rect 438 12566 442 12780
rect 462 12566 466 12780
rect 486 12566 490 12780
rect 510 12566 514 12780
rect 534 12566 538 12780
rect 558 12566 562 12780
rect 582 12566 586 12780
rect 606 12566 610 12780
rect 630 12566 634 12780
rect 654 12566 658 12780
rect 678 12566 682 12780
rect 691 12629 696 12639
rect 702 12629 706 12780
rect 701 12615 706 12629
rect 726 12566 730 12780
rect 750 12566 754 12780
rect 774 12566 778 12780
rect 798 12566 802 12780
rect 822 12566 826 12780
rect 846 12566 850 12780
rect 870 12566 874 12780
rect 894 12566 898 12780
rect 918 12566 922 12780
rect 942 12566 946 12780
rect 966 12566 970 12780
rect 990 12566 994 12780
rect 1014 12566 1018 12780
rect 1038 12566 1042 12780
rect 1062 12566 1066 12780
rect 1086 12566 1090 12780
rect 1110 12566 1114 12780
rect 1134 12566 1138 12780
rect 1158 12566 1162 12780
rect 1182 12566 1186 12780
rect 1206 12566 1210 12780
rect 1230 12566 1234 12780
rect 1254 12566 1258 12780
rect 1278 12566 1282 12780
rect 1302 12566 1306 12780
rect 1326 12566 1330 12780
rect 1350 12566 1354 12780
rect 1374 12566 1378 12780
rect 1398 12566 1402 12780
rect 1422 12566 1426 12780
rect 1446 12566 1450 12780
rect 1470 12566 1474 12780
rect 1494 12566 1498 12780
rect 1518 12566 1522 12780
rect 1542 12566 1546 12780
rect 1566 12566 1570 12780
rect 1590 12566 1594 12780
rect 1614 12566 1618 12780
rect 1638 12566 1642 12780
rect 1662 12566 1666 12780
rect 1686 12566 1690 12780
rect 1710 12566 1714 12780
rect 1734 12566 1738 12780
rect 1758 12566 1762 12780
rect 1782 12566 1786 12780
rect 1806 12566 1810 12780
rect 1830 12566 1834 12780
rect 1854 12566 1858 12780
rect 1878 12566 1882 12780
rect 1902 12566 1906 12780
rect 1926 12566 1930 12780
rect 1950 12566 1954 12780
rect 1974 12566 1978 12780
rect 1998 12566 2002 12780
rect 2022 12566 2026 12780
rect 2046 12566 2050 12780
rect 2070 12566 2074 12780
rect 2094 12566 2098 12780
rect 2118 12566 2122 12780
rect 2142 12566 2146 12780
rect 2166 12566 2170 12780
rect 2190 12567 2194 12780
rect 2179 12566 2213 12567
rect -971 12564 2213 12566
rect -971 12563 -957 12564
rect -954 12563 -947 12564
rect -954 12542 -950 12563
rect -930 12542 -926 12564
rect -906 12542 -902 12564
rect -882 12542 -878 12564
rect -858 12543 -854 12564
rect -869 12542 -835 12543
rect -2393 12540 -835 12542
rect -2371 12494 -2366 12540
rect -2348 12494 -2343 12540
rect -2325 12528 -2320 12540
rect -2079 12538 -2071 12540
rect -2072 12536 -2071 12538
rect -2109 12531 -2101 12536
rect -2101 12529 -2079 12531
rect -2069 12529 -2068 12536
rect -2325 12520 -2317 12528
rect -2079 12524 -2071 12529
rect -2325 12500 -2320 12520
rect -2317 12512 -2309 12520
rect -2074 12515 -2071 12524
rect -2069 12520 -2068 12524
rect -2109 12506 -2079 12509
rect -2325 12494 -2317 12500
rect -2119 12494 -2069 12496
rect -2056 12494 -2026 12497
rect -2000 12494 -1992 12540
rect -1846 12538 -1806 12540
rect -1854 12533 -1806 12537
rect -1854 12531 -1846 12533
rect -1846 12529 -1806 12531
rect -1806 12527 -1798 12529
rect -1846 12524 -1798 12527
rect -1846 12511 -1806 12522
rect -1671 12520 -1663 12528
rect -1663 12512 -1655 12520
rect -1854 12506 -1680 12510
rect -1926 12494 -1892 12497
rect -1671 12494 -1663 12500
rect -1642 12494 -1637 12540
rect -1619 12494 -1614 12540
rect -1530 12494 -1526 12540
rect -1506 12494 -1502 12540
rect -1482 12494 -1478 12540
rect -1458 12494 -1454 12540
rect -1434 12494 -1430 12540
rect -1410 12494 -1406 12540
rect -1386 12494 -1382 12540
rect -1362 12494 -1358 12540
rect -1338 12494 -1334 12540
rect -1314 12494 -1310 12540
rect -1290 12494 -1286 12540
rect -1266 12494 -1262 12540
rect -1242 12494 -1238 12540
rect -1218 12494 -1214 12540
rect -1194 12494 -1190 12540
rect -1170 12494 -1166 12540
rect -1146 12494 -1142 12540
rect -1122 12494 -1118 12540
rect -1098 12494 -1094 12540
rect -1074 12494 -1070 12540
rect -1050 12494 -1046 12540
rect -1026 12494 -1022 12540
rect -1002 12494 -998 12540
rect -978 12494 -974 12540
rect -954 12494 -950 12540
rect -930 12494 -926 12540
rect -906 12494 -902 12540
rect -882 12494 -878 12540
rect -869 12533 -864 12540
rect -858 12533 -854 12540
rect -859 12519 -854 12533
rect -858 12494 -854 12519
rect -834 12494 -830 12564
rect -810 12494 -806 12564
rect -786 12494 -782 12564
rect -762 12494 -758 12564
rect -738 12494 -734 12564
rect -714 12494 -710 12564
rect -690 12494 -686 12564
rect -666 12494 -662 12564
rect -642 12494 -638 12564
rect -618 12494 -614 12564
rect -594 12494 -590 12564
rect -570 12494 -566 12564
rect -546 12494 -542 12564
rect -522 12494 -518 12564
rect -498 12494 -494 12564
rect -474 12494 -470 12564
rect -450 12494 -446 12564
rect -426 12494 -422 12564
rect -402 12494 -398 12564
rect -378 12494 -374 12564
rect -354 12494 -350 12564
rect -330 12494 -326 12564
rect -306 12494 -302 12564
rect -282 12494 -278 12564
rect -258 12494 -254 12564
rect -234 12494 -230 12564
rect -210 12494 -206 12564
rect -186 12494 -182 12564
rect -162 12494 -158 12564
rect -138 12494 -134 12564
rect -114 12494 -110 12564
rect -90 12494 -86 12564
rect -66 12494 -62 12564
rect -42 12494 -38 12564
rect -18 12494 -14 12564
rect 6 12494 10 12564
rect 30 12494 34 12564
rect 54 12494 58 12564
rect 78 12494 82 12564
rect 102 12494 106 12564
rect 126 12494 130 12564
rect 150 12494 154 12564
rect 174 12494 178 12564
rect 198 12494 202 12564
rect 222 12494 226 12564
rect 246 12494 250 12564
rect 270 12494 274 12564
rect 294 12494 298 12564
rect 318 12494 322 12564
rect 342 12494 346 12564
rect 366 12494 370 12564
rect 390 12494 394 12564
rect 414 12494 418 12564
rect 438 12494 442 12564
rect 462 12494 466 12564
rect 486 12494 490 12564
rect 510 12494 514 12564
rect 534 12494 538 12564
rect 558 12494 562 12564
rect 582 12494 586 12564
rect 606 12494 610 12564
rect 630 12494 634 12564
rect 654 12494 658 12564
rect 678 12494 682 12564
rect 726 12563 730 12564
rect 691 12540 723 12543
rect 691 12533 696 12540
rect 709 12539 723 12540
rect 726 12539 733 12563
rect 701 12519 706 12533
rect 702 12494 706 12519
rect 750 12494 754 12564
rect 774 12494 778 12564
rect 798 12494 802 12564
rect 822 12494 826 12564
rect 846 12494 850 12564
rect 870 12494 874 12564
rect 894 12494 898 12564
rect 918 12494 922 12564
rect 942 12494 946 12564
rect 966 12494 970 12564
rect 990 12494 994 12564
rect 1014 12494 1018 12564
rect 1038 12494 1042 12564
rect 1062 12494 1066 12564
rect 1086 12494 1090 12564
rect 1110 12494 1114 12564
rect 1134 12494 1138 12564
rect 1158 12494 1162 12564
rect 1182 12494 1186 12564
rect 1206 12494 1210 12564
rect 1230 12494 1234 12564
rect 1254 12494 1258 12564
rect 1278 12494 1282 12564
rect 1302 12494 1306 12564
rect 1326 12494 1330 12564
rect 1350 12494 1354 12564
rect 1374 12494 1378 12564
rect 1398 12494 1402 12564
rect 1422 12494 1426 12564
rect 1446 12494 1450 12564
rect 1470 12494 1474 12564
rect 1494 12494 1498 12564
rect 1518 12494 1522 12564
rect 1542 12494 1546 12564
rect 1566 12494 1570 12564
rect 1590 12494 1594 12564
rect 1614 12494 1618 12564
rect 1638 12494 1642 12564
rect 1662 12494 1666 12564
rect 1686 12494 1690 12564
rect 1710 12494 1714 12564
rect 1734 12494 1738 12564
rect 1758 12494 1762 12564
rect 1782 12494 1786 12564
rect 1806 12494 1810 12564
rect 1830 12494 1834 12564
rect 1854 12494 1858 12564
rect 1878 12494 1882 12564
rect 1902 12494 1906 12564
rect 1926 12494 1930 12564
rect 1950 12494 1954 12564
rect 1974 12494 1978 12564
rect 1998 12494 2002 12564
rect 2022 12494 2026 12564
rect 2046 12494 2050 12564
rect 2070 12494 2074 12564
rect 2094 12494 2098 12564
rect 2118 12494 2122 12564
rect 2142 12494 2146 12564
rect 2166 12494 2170 12564
rect 2179 12557 2184 12564
rect 2190 12557 2194 12564
rect 2189 12543 2194 12557
rect 2179 12518 2213 12519
rect 2214 12518 2218 12780
rect 2238 12518 2242 12780
rect 2251 12605 2256 12615
rect 2262 12605 2266 12780
rect 2261 12591 2266 12605
rect 2251 12566 2285 12567
rect 2286 12566 2290 12780
rect 2310 12566 2314 12780
rect 2334 12566 2338 12780
rect 2358 12566 2362 12780
rect 2382 12566 2386 12780
rect 2395 12581 2400 12591
rect 2406 12581 2410 12780
rect 2405 12567 2410 12581
rect 2430 12566 2434 12780
rect 2454 12566 2458 12780
rect 2478 12566 2482 12780
rect 2502 12566 2506 12780
rect 2526 12566 2530 12780
rect 2550 12566 2554 12780
rect 2574 12566 2578 12780
rect 2598 12566 2602 12780
rect 2622 12566 2626 12780
rect 2646 12566 2650 12780
rect 2670 12566 2674 12780
rect 2694 12566 2698 12780
rect 2718 12566 2722 12780
rect 2742 12566 2746 12780
rect 2766 12566 2770 12780
rect 2790 12566 2794 12780
rect 2814 12566 2818 12780
rect 2838 12566 2842 12780
rect 2862 12566 2866 12780
rect 2886 12566 2890 12780
rect 2910 12566 2914 12780
rect 2934 12566 2938 12780
rect 2958 12566 2962 12780
rect 2982 12566 2986 12780
rect 3006 12566 3010 12780
rect 3030 12566 3034 12780
rect 3054 12566 3058 12780
rect 3078 12566 3082 12780
rect 3102 12566 3106 12780
rect 3126 12566 3130 12780
rect 3150 12566 3154 12780
rect 3174 12566 3178 12780
rect 3198 12566 3202 12780
rect 3222 12566 3226 12780
rect 3246 12566 3250 12780
rect 3270 12566 3274 12780
rect 3294 12566 3298 12780
rect 3318 12566 3322 12780
rect 3342 12566 3346 12780
rect 3366 12566 3370 12780
rect 3390 12566 3394 12780
rect 3414 12567 3418 12780
rect 3427 12653 3432 12663
rect 3438 12653 3442 12780
rect 3451 12773 3456 12780
rect 3462 12773 3466 12780
rect 3461 12759 3466 12773
rect 3437 12639 3442 12653
rect 3403 12566 3437 12567
rect 2251 12564 3437 12566
rect 2251 12557 2256 12564
rect 2261 12543 2266 12557
rect 2262 12518 2266 12543
rect 2286 12539 2290 12564
rect 2179 12516 2283 12518
rect 2179 12509 2184 12516
rect 2189 12495 2194 12509
rect 2190 12494 2194 12495
rect 2214 12494 2218 12516
rect 2238 12494 2242 12516
rect 2262 12494 2266 12516
rect 2269 12515 2283 12516
rect 2286 12515 2293 12539
rect 2310 12494 2314 12564
rect 2334 12494 2338 12564
rect 2358 12494 2362 12564
rect 2382 12494 2386 12564
rect 2430 12515 2434 12564
rect 2395 12494 2427 12495
rect -2393 12492 2427 12494
rect -2371 12470 -2366 12492
rect -2348 12470 -2343 12492
rect -2325 12488 -2317 12492
rect -2325 12472 -2320 12488
rect -2317 12484 -2309 12488
rect -2309 12472 -2301 12484
rect -2109 12475 -2079 12482
rect -2000 12481 -1992 12492
rect -1671 12488 -1663 12492
rect -1846 12484 -1806 12486
rect -1663 12484 -1655 12488
rect -2009 12478 -1992 12481
rect -1854 12478 -1806 12482
rect -2071 12475 -1992 12478
rect -1983 12475 -1806 12478
rect -2009 12472 -1992 12475
rect -2325 12470 -2317 12472
rect -2033 12470 -1992 12472
rect -1846 12471 -1806 12473
rect -1655 12472 -1647 12484
rect -1864 12470 -1796 12471
rect -1671 12470 -1663 12472
rect -1642 12470 -1637 12492
rect -1619 12470 -1614 12492
rect -1530 12470 -1526 12492
rect -1506 12470 -1502 12492
rect -1482 12470 -1478 12492
rect -1458 12470 -1454 12492
rect -1434 12470 -1430 12492
rect -1410 12470 -1406 12492
rect -1386 12470 -1382 12492
rect -1362 12470 -1358 12492
rect -1338 12470 -1334 12492
rect -1314 12470 -1310 12492
rect -1290 12470 -1286 12492
rect -1266 12470 -1262 12492
rect -1242 12470 -1238 12492
rect -1218 12470 -1214 12492
rect -1194 12470 -1190 12492
rect -1170 12470 -1166 12492
rect -1146 12470 -1142 12492
rect -1122 12470 -1118 12492
rect -1098 12470 -1094 12492
rect -1074 12470 -1070 12492
rect -1050 12471 -1046 12492
rect -1061 12470 -1027 12471
rect -2393 12468 -1027 12470
rect -2371 12446 -2366 12468
rect -2348 12446 -2343 12468
rect -2325 12460 -2317 12468
rect -2079 12465 -2035 12468
rect -2013 12466 -1992 12468
rect -2000 12465 -1992 12466
rect -1904 12465 -1798 12468
rect -2101 12461 -2009 12465
rect -2023 12460 -2009 12461
rect -2000 12463 -1798 12465
rect -2000 12461 -1854 12463
rect -1846 12461 -1798 12463
rect -2325 12446 -2320 12460
rect -2317 12456 -2309 12460
rect -2309 12446 -2301 12456
rect -2109 12448 -2101 12455
rect -2023 12451 -2021 12460
rect -2000 12451 -1992 12461
rect -1671 12460 -1663 12468
rect -1846 12457 -1806 12459
rect -1663 12456 -1655 12460
rect -1854 12451 -1806 12455
rect -2071 12448 -1806 12451
rect -2074 12446 -2031 12448
rect -2000 12446 -1992 12448
rect -1655 12446 -1647 12456
rect -1642 12446 -1637 12468
rect -1619 12446 -1614 12468
rect -1530 12446 -1526 12468
rect -1506 12446 -1502 12468
rect -1482 12446 -1478 12468
rect -1458 12446 -1454 12468
rect -1434 12446 -1430 12468
rect -1410 12446 -1406 12468
rect -1386 12446 -1382 12468
rect -1362 12446 -1358 12468
rect -1338 12446 -1334 12468
rect -1314 12446 -1310 12468
rect -1290 12446 -1286 12468
rect -1266 12446 -1262 12468
rect -1242 12446 -1238 12468
rect -1218 12446 -1214 12468
rect -1194 12446 -1190 12468
rect -1170 12446 -1166 12468
rect -1146 12446 -1142 12468
rect -1122 12446 -1118 12468
rect -1098 12446 -1094 12468
rect -1074 12446 -1070 12468
rect -1061 12461 -1056 12468
rect -1050 12461 -1046 12468
rect -1051 12447 -1046 12461
rect -1050 12446 -1046 12447
rect -1026 12446 -1022 12492
rect -1002 12446 -998 12492
rect -978 12446 -974 12492
rect -954 12446 -950 12492
rect -930 12446 -926 12492
rect -906 12446 -902 12492
rect -882 12446 -878 12492
rect -858 12446 -854 12492
rect -834 12467 -830 12492
rect -2393 12444 -837 12446
rect -2371 12398 -2366 12444
rect -2348 12398 -2343 12444
rect -2325 12432 -2317 12444
rect -2074 12441 -2071 12444
rect -2101 12434 -2071 12441
rect -2325 12412 -2320 12432
rect -2317 12428 -2309 12432
rect -2064 12430 -2061 12438
rect -2325 12404 -2317 12412
rect -2101 12407 -2071 12410
rect -2325 12398 -2320 12404
rect -2317 12398 -2309 12404
rect -2000 12402 -1992 12444
rect -1846 12443 -1806 12444
rect -1846 12434 -1798 12441
rect -1671 12432 -1663 12444
rect -1846 12430 -1806 12432
rect -1663 12428 -1655 12432
rect -1854 12416 -1680 12420
rect -1846 12407 -1798 12410
rect -2079 12401 -2043 12402
rect -2007 12401 -1991 12402
rect -2079 12400 -2071 12401
rect -2079 12398 -2029 12400
rect -2011 12398 -1991 12401
rect -1846 12399 -1806 12405
rect -1671 12404 -1663 12412
rect -1864 12398 -1796 12399
rect -1663 12398 -1655 12404
rect -1642 12398 -1637 12444
rect -1619 12398 -1614 12444
rect -1530 12398 -1526 12444
rect -1506 12398 -1502 12444
rect -1482 12398 -1478 12444
rect -1458 12398 -1454 12444
rect -1434 12398 -1430 12444
rect -1410 12398 -1406 12444
rect -1386 12398 -1382 12444
rect -1362 12398 -1358 12444
rect -1338 12398 -1334 12444
rect -1314 12398 -1310 12444
rect -1290 12398 -1286 12444
rect -1266 12398 -1262 12444
rect -1242 12398 -1238 12444
rect -1218 12398 -1214 12444
rect -1194 12398 -1190 12444
rect -1170 12398 -1166 12444
rect -1146 12398 -1142 12444
rect -1122 12398 -1118 12444
rect -1098 12398 -1094 12444
rect -1074 12399 -1070 12444
rect -1085 12398 -1051 12399
rect -2393 12396 -1051 12398
rect -2371 12350 -2366 12396
rect -2348 12350 -2343 12396
rect -2325 12384 -2320 12396
rect -2079 12394 -2071 12396
rect -2072 12392 -2071 12394
rect -2109 12387 -2101 12392
rect -2101 12385 -2079 12387
rect -2069 12385 -2068 12392
rect -2325 12376 -2317 12384
rect -2079 12380 -2071 12385
rect -2325 12356 -2320 12376
rect -2317 12368 -2309 12376
rect -2074 12371 -2071 12380
rect -2069 12376 -2068 12380
rect -2109 12362 -2079 12365
rect -2325 12350 -2317 12356
rect -2000 12350 -1992 12396
rect -1846 12394 -1806 12396
rect -1854 12389 -1806 12393
rect -1854 12387 -1846 12389
rect -1846 12385 -1806 12387
rect -1806 12383 -1798 12385
rect -1846 12380 -1798 12383
rect -1846 12367 -1806 12378
rect -1671 12376 -1663 12384
rect -1663 12368 -1655 12376
rect -1854 12362 -1680 12366
rect -1671 12350 -1663 12356
rect -1642 12350 -1637 12396
rect -1619 12350 -1614 12396
rect -1530 12350 -1526 12396
rect -1506 12350 -1502 12396
rect -1482 12350 -1478 12396
rect -1458 12350 -1454 12396
rect -1434 12350 -1430 12396
rect -1410 12350 -1406 12396
rect -1386 12350 -1382 12396
rect -1362 12350 -1358 12396
rect -1338 12350 -1334 12396
rect -1314 12350 -1310 12396
rect -1290 12350 -1286 12396
rect -1266 12350 -1262 12396
rect -1242 12350 -1238 12396
rect -1218 12350 -1214 12396
rect -1194 12350 -1190 12396
rect -1170 12350 -1166 12396
rect -1146 12350 -1142 12396
rect -1122 12350 -1118 12396
rect -1098 12350 -1094 12396
rect -1085 12389 -1080 12396
rect -1074 12389 -1070 12396
rect -1075 12375 -1070 12389
rect -1085 12374 -1051 12375
rect -1050 12374 -1046 12444
rect -1026 12395 -1022 12444
rect -1085 12372 -1029 12374
rect -1085 12365 -1080 12372
rect -1075 12351 -1070 12365
rect -1074 12350 -1070 12351
rect -1050 12350 -1046 12372
rect -1043 12371 -1029 12372
rect -1026 12371 -1019 12395
rect -1026 12350 -1022 12371
rect -1002 12350 -998 12444
rect -978 12350 -974 12444
rect -954 12350 -950 12444
rect -930 12350 -926 12444
rect -906 12350 -902 12444
rect -882 12350 -878 12444
rect -858 12350 -854 12444
rect -851 12443 -837 12444
rect -834 12443 -827 12467
rect -834 12350 -830 12443
rect -810 12350 -806 12492
rect -786 12350 -782 12492
rect -762 12350 -758 12492
rect -738 12350 -734 12492
rect -714 12350 -710 12492
rect -690 12350 -686 12492
rect -666 12350 -662 12492
rect -653 12413 -648 12423
rect -642 12413 -638 12492
rect -643 12399 -638 12413
rect -653 12398 -619 12399
rect -618 12398 -614 12492
rect -594 12398 -590 12492
rect -570 12398 -566 12492
rect -546 12398 -542 12492
rect -522 12398 -518 12492
rect -498 12398 -494 12492
rect -474 12398 -470 12492
rect -450 12398 -446 12492
rect -426 12398 -422 12492
rect -402 12398 -398 12492
rect -378 12398 -374 12492
rect -354 12398 -350 12492
rect -330 12398 -326 12492
rect -306 12398 -302 12492
rect -282 12398 -278 12492
rect -258 12398 -254 12492
rect -234 12398 -230 12492
rect -210 12398 -206 12492
rect -186 12398 -182 12492
rect -162 12398 -158 12492
rect -138 12398 -134 12492
rect -114 12398 -110 12492
rect -90 12398 -86 12492
rect -66 12398 -62 12492
rect -42 12398 -38 12492
rect -18 12398 -14 12492
rect 6 12398 10 12492
rect 30 12398 34 12492
rect 54 12398 58 12492
rect 78 12398 82 12492
rect 102 12398 106 12492
rect 126 12398 130 12492
rect 150 12398 154 12492
rect 174 12398 178 12492
rect 198 12398 202 12492
rect 222 12398 226 12492
rect 246 12398 250 12492
rect 270 12398 274 12492
rect 294 12398 298 12492
rect 318 12398 322 12492
rect 342 12398 346 12492
rect 366 12398 370 12492
rect 390 12398 394 12492
rect 414 12398 418 12492
rect 438 12398 442 12492
rect 462 12398 466 12492
rect 486 12398 490 12492
rect 510 12398 514 12492
rect 534 12398 538 12492
rect 558 12398 562 12492
rect 582 12398 586 12492
rect 606 12398 610 12492
rect 630 12398 634 12492
rect 654 12398 658 12492
rect 678 12398 682 12492
rect 702 12398 706 12492
rect 726 12446 733 12467
rect 750 12446 754 12492
rect 774 12446 778 12492
rect 798 12446 802 12492
rect 822 12446 826 12492
rect 846 12446 850 12492
rect 870 12446 874 12492
rect 894 12446 898 12492
rect 918 12446 922 12492
rect 942 12446 946 12492
rect 966 12446 970 12492
rect 990 12446 994 12492
rect 1014 12446 1018 12492
rect 1038 12446 1042 12492
rect 1062 12446 1066 12492
rect 1086 12446 1090 12492
rect 1110 12446 1114 12492
rect 1134 12446 1138 12492
rect 1158 12446 1162 12492
rect 1182 12446 1186 12492
rect 1206 12446 1210 12492
rect 1230 12446 1234 12492
rect 1254 12446 1258 12492
rect 1278 12446 1282 12492
rect 1302 12446 1306 12492
rect 1326 12446 1330 12492
rect 1350 12446 1354 12492
rect 1374 12446 1378 12492
rect 1398 12446 1402 12492
rect 1422 12446 1426 12492
rect 1446 12446 1450 12492
rect 1470 12446 1474 12492
rect 1494 12446 1498 12492
rect 1518 12446 1522 12492
rect 1542 12446 1546 12492
rect 1566 12446 1570 12492
rect 1590 12446 1594 12492
rect 1614 12446 1618 12492
rect 1638 12446 1642 12492
rect 1662 12446 1666 12492
rect 1686 12446 1690 12492
rect 1710 12446 1714 12492
rect 1734 12446 1738 12492
rect 1758 12446 1762 12492
rect 1782 12446 1786 12492
rect 1806 12446 1810 12492
rect 1830 12446 1834 12492
rect 1854 12446 1858 12492
rect 1878 12446 1882 12492
rect 1902 12446 1906 12492
rect 1926 12446 1930 12492
rect 1950 12446 1954 12492
rect 1974 12446 1978 12492
rect 1998 12446 2002 12492
rect 2022 12446 2026 12492
rect 2046 12446 2050 12492
rect 2070 12446 2074 12492
rect 2094 12446 2098 12492
rect 2118 12446 2122 12492
rect 2142 12446 2146 12492
rect 2166 12446 2170 12492
rect 2190 12446 2194 12492
rect 2214 12491 2218 12492
rect 2214 12467 2221 12491
rect 2238 12446 2242 12492
rect 2262 12446 2266 12492
rect 2286 12467 2293 12491
rect 2286 12446 2290 12467
rect 2310 12446 2314 12492
rect 2334 12446 2338 12492
rect 2358 12446 2362 12492
rect 2382 12446 2386 12492
rect 2395 12485 2400 12492
rect 2413 12491 2427 12492
rect 2430 12491 2437 12515
rect 2405 12471 2410 12485
rect 2406 12446 2410 12471
rect 2454 12446 2458 12564
rect 2478 12446 2482 12564
rect 2502 12446 2506 12564
rect 2526 12446 2530 12564
rect 2550 12446 2554 12564
rect 2574 12446 2578 12564
rect 2598 12446 2602 12564
rect 2622 12446 2626 12564
rect 2646 12446 2650 12564
rect 2670 12446 2674 12564
rect 2694 12446 2698 12564
rect 2718 12446 2722 12564
rect 2742 12446 2746 12564
rect 2766 12446 2770 12564
rect 2790 12446 2794 12564
rect 2814 12446 2818 12564
rect 2838 12446 2842 12564
rect 2862 12446 2866 12564
rect 2886 12446 2890 12564
rect 2910 12446 2914 12564
rect 2934 12446 2938 12564
rect 2958 12446 2962 12564
rect 2982 12446 2986 12564
rect 3006 12446 3010 12564
rect 3030 12447 3034 12564
rect 3019 12446 3053 12447
rect 709 12444 3053 12446
rect 709 12443 723 12444
rect 726 12443 733 12444
rect 726 12398 730 12443
rect 750 12398 754 12444
rect 774 12398 778 12444
rect 798 12398 802 12444
rect 822 12398 826 12444
rect 846 12398 850 12444
rect 870 12398 874 12444
rect 894 12398 898 12444
rect 918 12398 922 12444
rect 942 12398 946 12444
rect 966 12398 970 12444
rect 990 12398 994 12444
rect 1014 12398 1018 12444
rect 1038 12398 1042 12444
rect 1062 12398 1066 12444
rect 1086 12398 1090 12444
rect 1110 12398 1114 12444
rect 1134 12398 1138 12444
rect 1158 12398 1162 12444
rect 1182 12398 1186 12444
rect 1206 12398 1210 12444
rect 1230 12398 1234 12444
rect 1254 12398 1258 12444
rect 1278 12398 1282 12444
rect 1302 12398 1306 12444
rect 1326 12398 1330 12444
rect 1350 12398 1354 12444
rect 1374 12398 1378 12444
rect 1398 12398 1402 12444
rect 1422 12398 1426 12444
rect 1446 12398 1450 12444
rect 1470 12398 1474 12444
rect 1494 12398 1498 12444
rect 1518 12398 1522 12444
rect 1542 12398 1546 12444
rect 1566 12398 1570 12444
rect 1590 12398 1594 12444
rect 1614 12398 1618 12444
rect 1638 12398 1642 12444
rect 1662 12398 1666 12444
rect 1686 12398 1690 12444
rect 1710 12398 1714 12444
rect 1734 12398 1738 12444
rect 1758 12398 1762 12444
rect 1782 12398 1786 12444
rect 1806 12398 1810 12444
rect 1830 12398 1834 12444
rect 1854 12398 1858 12444
rect 1878 12398 1882 12444
rect 1902 12398 1906 12444
rect 1926 12398 1930 12444
rect 1950 12398 1954 12444
rect 1974 12398 1978 12444
rect 1998 12398 2002 12444
rect 2022 12398 2026 12444
rect 2046 12398 2050 12444
rect 2070 12398 2074 12444
rect 2094 12398 2098 12444
rect 2118 12398 2122 12444
rect 2142 12398 2146 12444
rect 2166 12398 2170 12444
rect 2190 12398 2194 12444
rect 2214 12419 2221 12443
rect 2214 12398 2218 12419
rect 2238 12398 2242 12444
rect 2262 12398 2266 12444
rect 2286 12398 2290 12444
rect 2310 12398 2314 12444
rect 2334 12398 2338 12444
rect 2358 12398 2362 12444
rect 2382 12398 2386 12444
rect 2406 12398 2410 12444
rect -653 12396 2427 12398
rect -653 12389 -648 12396
rect -643 12375 -638 12389
rect -642 12350 -638 12375
rect -618 12350 -614 12396
rect -594 12350 -590 12396
rect -570 12350 -566 12396
rect -546 12350 -542 12396
rect -522 12350 -518 12396
rect -498 12350 -494 12396
rect -474 12350 -470 12396
rect -450 12350 -446 12396
rect -426 12350 -422 12396
rect -402 12350 -398 12396
rect -378 12350 -374 12396
rect -354 12350 -350 12396
rect -330 12350 -326 12396
rect -306 12350 -302 12396
rect -282 12350 -278 12396
rect -258 12350 -254 12396
rect -234 12350 -230 12396
rect -210 12350 -206 12396
rect -186 12350 -182 12396
rect -162 12350 -158 12396
rect -138 12350 -134 12396
rect -114 12350 -110 12396
rect -90 12350 -86 12396
rect -66 12350 -62 12396
rect -42 12350 -38 12396
rect -18 12350 -14 12396
rect 6 12350 10 12396
rect 30 12350 34 12396
rect 54 12350 58 12396
rect 78 12350 82 12396
rect 102 12350 106 12396
rect 126 12350 130 12396
rect 150 12350 154 12396
rect 174 12350 178 12396
rect 198 12350 202 12396
rect 222 12350 226 12396
rect 246 12350 250 12396
rect 270 12350 274 12396
rect 294 12350 298 12396
rect 318 12350 322 12396
rect 342 12350 346 12396
rect 366 12350 370 12396
rect 390 12350 394 12396
rect 414 12350 418 12396
rect 438 12350 442 12396
rect 462 12350 466 12396
rect 486 12350 490 12396
rect 510 12350 514 12396
rect 534 12350 538 12396
rect 558 12350 562 12396
rect 582 12350 586 12396
rect 606 12350 610 12396
rect 630 12350 634 12396
rect 654 12350 658 12396
rect 678 12350 682 12396
rect 702 12350 706 12396
rect 726 12350 730 12396
rect 750 12350 754 12396
rect 774 12350 778 12396
rect 798 12350 802 12396
rect 822 12350 826 12396
rect 846 12350 850 12396
rect 870 12350 874 12396
rect 894 12350 898 12396
rect 918 12350 922 12396
rect 942 12350 946 12396
rect 966 12350 970 12396
rect 990 12350 994 12396
rect 1014 12350 1018 12396
rect 1038 12350 1042 12396
rect 1062 12350 1066 12396
rect 1086 12350 1090 12396
rect 1110 12350 1114 12396
rect 1134 12350 1138 12396
rect 1158 12350 1162 12396
rect 1182 12350 1186 12396
rect 1206 12350 1210 12396
rect 1230 12350 1234 12396
rect 1254 12350 1258 12396
rect 1278 12350 1282 12396
rect 1302 12350 1306 12396
rect 1326 12350 1330 12396
rect 1350 12350 1354 12396
rect 1374 12350 1378 12396
rect 1398 12350 1402 12396
rect 1422 12350 1426 12396
rect 1446 12350 1450 12396
rect 1470 12350 1474 12396
rect 1494 12350 1498 12396
rect 1518 12350 1522 12396
rect 1542 12350 1546 12396
rect 1566 12350 1570 12396
rect 1590 12350 1594 12396
rect 1614 12350 1618 12396
rect 1638 12350 1642 12396
rect 1662 12350 1666 12396
rect 1686 12350 1690 12396
rect 1710 12350 1714 12396
rect 1734 12350 1738 12396
rect 1758 12350 1762 12396
rect 1782 12350 1786 12396
rect 1806 12350 1810 12396
rect 1830 12350 1834 12396
rect 1854 12350 1858 12396
rect 1878 12350 1882 12396
rect 1902 12350 1906 12396
rect 1926 12350 1930 12396
rect 1950 12350 1954 12396
rect 1974 12350 1978 12396
rect 1998 12350 2002 12396
rect 2022 12350 2026 12396
rect 2046 12350 2050 12396
rect 2070 12350 2074 12396
rect 2094 12350 2098 12396
rect 2118 12350 2122 12396
rect 2142 12350 2146 12396
rect 2166 12350 2170 12396
rect 2190 12350 2194 12396
rect 2214 12350 2218 12396
rect 2238 12350 2242 12396
rect 2262 12350 2266 12396
rect 2286 12350 2290 12396
rect 2310 12350 2314 12396
rect 2334 12350 2338 12396
rect 2358 12350 2362 12396
rect 2382 12350 2386 12396
rect 2406 12350 2410 12396
rect 2413 12395 2427 12396
rect 2430 12395 2437 12419
rect 2430 12350 2434 12395
rect 2454 12350 2458 12444
rect 2478 12350 2482 12444
rect 2502 12350 2506 12444
rect 2526 12350 2530 12444
rect 2550 12350 2554 12444
rect 2574 12350 2578 12444
rect 2598 12350 2602 12444
rect 2622 12350 2626 12444
rect 2646 12350 2650 12444
rect 2670 12350 2674 12444
rect 2694 12350 2698 12444
rect 2718 12350 2722 12444
rect 2742 12350 2746 12444
rect 2766 12350 2770 12444
rect 2790 12350 2794 12444
rect 2814 12350 2818 12444
rect 2838 12350 2842 12444
rect 2862 12350 2866 12444
rect 2886 12350 2890 12444
rect 2910 12350 2914 12444
rect 2934 12350 2938 12444
rect 2958 12350 2962 12444
rect 2982 12350 2986 12444
rect 3006 12350 3010 12444
rect 3019 12437 3024 12444
rect 3030 12437 3034 12444
rect 3029 12423 3034 12437
rect 3019 12422 3053 12423
rect 3054 12422 3058 12564
rect 3078 12422 3082 12564
rect 3102 12422 3106 12564
rect 3126 12422 3130 12564
rect 3150 12422 3154 12564
rect 3174 12422 3178 12564
rect 3198 12422 3202 12564
rect 3222 12422 3226 12564
rect 3246 12422 3250 12564
rect 3270 12422 3274 12564
rect 3294 12422 3298 12564
rect 3318 12422 3322 12564
rect 3342 12423 3346 12564
rect 3355 12509 3360 12519
rect 3366 12509 3370 12564
rect 3379 12533 3384 12543
rect 3390 12533 3394 12564
rect 3403 12557 3408 12564
rect 3414 12557 3418 12564
rect 3413 12543 3418 12557
rect 3389 12519 3394 12533
rect 3365 12495 3370 12509
rect 3331 12422 3365 12423
rect 3019 12420 3365 12422
rect 3019 12413 3024 12420
rect 3029 12399 3034 12413
rect 3030 12350 3034 12399
rect 3054 12371 3058 12420
rect -2393 12348 3051 12350
rect -2371 12326 -2366 12348
rect -2348 12326 -2343 12348
rect -2325 12340 -2317 12348
rect -2325 12326 -2320 12340
rect -2309 12328 -2301 12340
rect -2092 12331 -2062 12336
rect -2000 12328 -1992 12348
rect -2317 12326 -2309 12328
rect -2000 12326 -1983 12328
rect -1906 12326 -1904 12348
rect -1806 12340 -1680 12346
rect -1671 12340 -1663 12348
rect -1854 12331 -1806 12336
rect -1846 12326 -1806 12329
rect -1655 12328 -1647 12340
rect -1663 12326 -1655 12328
rect -1642 12326 -1637 12348
rect -1619 12326 -1614 12348
rect -1530 12326 -1526 12348
rect -1506 12326 -1502 12348
rect -1482 12326 -1478 12348
rect -1458 12326 -1454 12348
rect -1434 12326 -1430 12348
rect -1410 12326 -1406 12348
rect -1386 12326 -1382 12348
rect -1362 12326 -1358 12348
rect -1338 12327 -1334 12348
rect -1349 12326 -1315 12327
rect -2393 12324 -1315 12326
rect -2371 12302 -2366 12324
rect -2348 12302 -2343 12324
rect -2325 12312 -2317 12324
rect -2071 12320 -2062 12324
rect -2013 12322 -1983 12324
rect -2000 12321 -1983 12322
rect -2325 12302 -2320 12312
rect -2309 12302 -2301 12312
rect -2100 12311 -2092 12318
rect -2064 12316 -2062 12319
rect -2061 12311 -2059 12316
rect -2071 12306 -2062 12311
rect -2071 12304 -2026 12306
rect -2066 12302 -2012 12304
rect -2000 12302 -1992 12321
rect -1906 12319 -1904 12324
rect -1846 12320 -1806 12324
rect -1846 12313 -1798 12318
rect -1806 12311 -1798 12313
rect -1671 12312 -1663 12324
rect -1854 12309 -1846 12311
rect -1854 12304 -1806 12309
rect -1864 12302 -1796 12303
rect -1655 12302 -1647 12312
rect -1642 12302 -1637 12324
rect -1619 12302 -1614 12324
rect -1530 12302 -1526 12324
rect -1506 12302 -1502 12324
rect -1482 12302 -1478 12324
rect -1458 12302 -1454 12324
rect -1434 12302 -1430 12324
rect -1410 12302 -1406 12324
rect -1386 12302 -1382 12324
rect -1362 12302 -1358 12324
rect -1349 12317 -1344 12324
rect -1338 12317 -1334 12324
rect -1339 12303 -1334 12317
rect -1314 12302 -1310 12348
rect -1290 12302 -1286 12348
rect -1266 12302 -1262 12348
rect -1242 12302 -1238 12348
rect -1218 12302 -1214 12348
rect -1194 12302 -1190 12348
rect -1170 12302 -1166 12348
rect -1146 12302 -1142 12348
rect -1122 12302 -1118 12348
rect -1098 12302 -1094 12348
rect -1074 12302 -1070 12348
rect -1050 12323 -1046 12348
rect -2393 12300 -1053 12302
rect -2371 12254 -2366 12300
rect -2348 12254 -2343 12300
rect -2325 12296 -2320 12300
rect -2317 12296 -2309 12300
rect -2325 12284 -2317 12296
rect -2066 12295 -2062 12300
rect -2147 12292 -2134 12294
rect -2292 12286 -2071 12292
rect -2325 12254 -2320 12284
rect -2092 12270 -2062 12272
rect -2094 12266 -2062 12270
rect -2000 12254 -1992 12300
rect -1846 12293 -1806 12300
rect -1663 12296 -1655 12300
rect -1846 12286 -1680 12292
rect -1671 12284 -1663 12296
rect -1854 12270 -1806 12272
rect -1854 12266 -1680 12270
rect -1642 12254 -1637 12300
rect -1619 12254 -1614 12300
rect -1530 12254 -1526 12300
rect -1506 12254 -1502 12300
rect -1482 12254 -1478 12300
rect -1458 12254 -1454 12300
rect -1434 12254 -1430 12300
rect -1410 12254 -1406 12300
rect -1386 12254 -1382 12300
rect -1362 12254 -1358 12300
rect -1349 12269 -1344 12279
rect -1339 12255 -1334 12269
rect -1338 12254 -1334 12255
rect -1314 12254 -1310 12300
rect -1290 12254 -1286 12300
rect -1266 12254 -1262 12300
rect -1242 12254 -1238 12300
rect -1218 12254 -1214 12300
rect -1194 12254 -1190 12300
rect -1170 12254 -1166 12300
rect -1146 12254 -1142 12300
rect -1122 12254 -1118 12300
rect -1098 12254 -1094 12300
rect -1074 12254 -1070 12300
rect -1067 12299 -1053 12300
rect -1050 12278 -1043 12323
rect -1026 12278 -1022 12348
rect -1002 12278 -998 12348
rect -978 12278 -974 12348
rect -954 12278 -950 12348
rect -930 12278 -926 12348
rect -906 12278 -902 12348
rect -882 12278 -878 12348
rect -858 12278 -854 12348
rect -834 12278 -830 12348
rect -810 12278 -806 12348
rect -786 12278 -782 12348
rect -762 12278 -758 12348
rect -738 12278 -734 12348
rect -714 12278 -710 12348
rect -690 12278 -686 12348
rect -666 12278 -662 12348
rect -642 12278 -638 12348
rect -618 12347 -614 12348
rect -618 12302 -611 12347
rect -594 12302 -590 12348
rect -570 12302 -566 12348
rect -546 12302 -542 12348
rect -522 12302 -518 12348
rect -498 12302 -494 12348
rect -474 12302 -470 12348
rect -450 12302 -446 12348
rect -426 12302 -422 12348
rect -402 12302 -398 12348
rect -378 12302 -374 12348
rect -354 12302 -350 12348
rect -330 12302 -326 12348
rect -306 12302 -302 12348
rect -282 12302 -278 12348
rect -258 12302 -254 12348
rect -234 12302 -230 12348
rect -210 12302 -206 12348
rect -186 12302 -182 12348
rect -162 12302 -158 12348
rect -138 12302 -134 12348
rect -114 12302 -110 12348
rect -90 12302 -86 12348
rect -66 12302 -62 12348
rect -42 12302 -38 12348
rect -18 12302 -14 12348
rect 6 12302 10 12348
rect 30 12302 34 12348
rect 54 12302 58 12348
rect 78 12302 82 12348
rect 102 12302 106 12348
rect 126 12302 130 12348
rect 150 12302 154 12348
rect 174 12302 178 12348
rect 198 12302 202 12348
rect 222 12302 226 12348
rect 246 12302 250 12348
rect 270 12302 274 12348
rect 294 12302 298 12348
rect 318 12302 322 12348
rect 342 12302 346 12348
rect 366 12302 370 12348
rect 390 12302 394 12348
rect 414 12302 418 12348
rect 438 12302 442 12348
rect 462 12302 466 12348
rect 486 12302 490 12348
rect 510 12302 514 12348
rect 534 12302 538 12348
rect 558 12302 562 12348
rect 582 12302 586 12348
rect 606 12302 610 12348
rect 630 12302 634 12348
rect 654 12302 658 12348
rect 678 12302 682 12348
rect 702 12302 706 12348
rect 726 12302 730 12348
rect 750 12302 754 12348
rect 774 12302 778 12348
rect 798 12302 802 12348
rect 822 12302 826 12348
rect 846 12302 850 12348
rect 870 12302 874 12348
rect 894 12302 898 12348
rect 918 12302 922 12348
rect 942 12302 946 12348
rect 966 12302 970 12348
rect 990 12302 994 12348
rect 1014 12302 1018 12348
rect 1038 12302 1042 12348
rect 1062 12302 1066 12348
rect 1086 12302 1090 12348
rect 1110 12302 1114 12348
rect 1134 12302 1138 12348
rect 1158 12302 1162 12348
rect 1182 12302 1186 12348
rect 1206 12302 1210 12348
rect 1230 12302 1234 12348
rect 1254 12302 1258 12348
rect 1278 12302 1282 12348
rect 1302 12302 1306 12348
rect 1326 12302 1330 12348
rect 1350 12302 1354 12348
rect 1374 12302 1378 12348
rect 1398 12302 1402 12348
rect 1422 12302 1426 12348
rect 1446 12302 1450 12348
rect 1470 12302 1474 12348
rect 1494 12302 1498 12348
rect 1518 12302 1522 12348
rect 1542 12302 1546 12348
rect 1566 12302 1570 12348
rect 1590 12302 1594 12348
rect 1614 12302 1618 12348
rect 1638 12302 1642 12348
rect 1662 12302 1666 12348
rect 1686 12302 1690 12348
rect 1710 12302 1714 12348
rect 1734 12302 1738 12348
rect 1758 12302 1762 12348
rect 1782 12302 1786 12348
rect 1806 12302 1810 12348
rect 1830 12302 1834 12348
rect 1854 12302 1858 12348
rect 1878 12302 1882 12348
rect 1902 12302 1906 12348
rect 1926 12302 1930 12348
rect 1950 12302 1954 12348
rect 1974 12302 1978 12348
rect 1998 12302 2002 12348
rect 2022 12302 2026 12348
rect 2046 12302 2050 12348
rect 2070 12302 2074 12348
rect 2094 12302 2098 12348
rect 2118 12302 2122 12348
rect 2142 12302 2146 12348
rect 2166 12302 2170 12348
rect 2190 12302 2194 12348
rect 2214 12302 2218 12348
rect 2238 12302 2242 12348
rect 2262 12302 2266 12348
rect 2286 12302 2290 12348
rect 2310 12302 2314 12348
rect 2334 12302 2338 12348
rect 2358 12302 2362 12348
rect 2382 12302 2386 12348
rect 2406 12302 2410 12348
rect 2430 12302 2434 12348
rect 2454 12302 2458 12348
rect 2478 12302 2482 12348
rect 2502 12302 2506 12348
rect 2526 12302 2530 12348
rect 2550 12302 2554 12348
rect 2574 12302 2578 12348
rect 2598 12302 2602 12348
rect 2622 12302 2626 12348
rect 2646 12302 2650 12348
rect 2670 12302 2674 12348
rect 2694 12302 2698 12348
rect 2718 12302 2722 12348
rect 2742 12302 2746 12348
rect 2766 12302 2770 12348
rect 2790 12302 2794 12348
rect 2814 12302 2818 12348
rect 2838 12302 2842 12348
rect 2862 12302 2866 12348
rect 2886 12302 2890 12348
rect 2910 12302 2914 12348
rect 2934 12302 2938 12348
rect 2958 12302 2962 12348
rect 2982 12302 2986 12348
rect 3006 12302 3010 12348
rect 3030 12302 3034 12348
rect 3037 12347 3051 12348
rect 3054 12323 3061 12371
rect 3054 12302 3058 12323
rect 3078 12302 3082 12420
rect 3102 12302 3106 12420
rect 3126 12302 3130 12420
rect 3150 12302 3154 12420
rect 3174 12303 3178 12420
rect 3163 12302 3197 12303
rect -635 12300 3197 12302
rect -635 12299 -621 12300
rect -618 12299 -611 12300
rect -618 12278 -614 12299
rect -594 12278 -590 12300
rect -570 12278 -566 12300
rect -546 12278 -542 12300
rect -522 12278 -518 12300
rect -498 12278 -494 12300
rect -474 12278 -470 12300
rect -450 12278 -446 12300
rect -426 12278 -422 12300
rect -402 12278 -398 12300
rect -378 12278 -374 12300
rect -354 12278 -350 12300
rect -330 12278 -326 12300
rect -306 12278 -302 12300
rect -282 12278 -278 12300
rect -258 12278 -254 12300
rect -234 12278 -230 12300
rect -210 12278 -206 12300
rect -186 12278 -182 12300
rect -162 12278 -158 12300
rect -138 12278 -134 12300
rect -114 12278 -110 12300
rect -90 12278 -86 12300
rect -66 12278 -62 12300
rect -42 12278 -38 12300
rect -18 12278 -14 12300
rect 6 12278 10 12300
rect 30 12278 34 12300
rect 54 12278 58 12300
rect 78 12278 82 12300
rect 102 12278 106 12300
rect 126 12278 130 12300
rect 150 12278 154 12300
rect 174 12278 178 12300
rect 198 12278 202 12300
rect 222 12278 226 12300
rect 246 12278 250 12300
rect 270 12278 274 12300
rect 294 12278 298 12300
rect 318 12278 322 12300
rect 342 12278 346 12300
rect 366 12278 370 12300
rect 390 12278 394 12300
rect 414 12278 418 12300
rect 438 12278 442 12300
rect 462 12278 466 12300
rect 486 12278 490 12300
rect 510 12278 514 12300
rect 534 12278 538 12300
rect 558 12278 562 12300
rect 582 12278 586 12300
rect 606 12278 610 12300
rect 630 12278 634 12300
rect 654 12278 658 12300
rect 678 12278 682 12300
rect 702 12278 706 12300
rect 726 12278 730 12300
rect 750 12278 754 12300
rect 774 12278 778 12300
rect 798 12278 802 12300
rect 822 12278 826 12300
rect 846 12278 850 12300
rect 870 12278 874 12300
rect 894 12278 898 12300
rect 918 12278 922 12300
rect 942 12278 946 12300
rect 966 12278 970 12300
rect 990 12278 994 12300
rect 1014 12278 1018 12300
rect 1038 12278 1042 12300
rect 1062 12278 1066 12300
rect 1086 12278 1090 12300
rect 1110 12278 1114 12300
rect 1134 12278 1138 12300
rect 1158 12278 1162 12300
rect 1182 12278 1186 12300
rect 1206 12278 1210 12300
rect 1230 12278 1234 12300
rect 1254 12278 1258 12300
rect 1278 12278 1282 12300
rect 1302 12278 1306 12300
rect 1326 12278 1330 12300
rect 1350 12278 1354 12300
rect 1374 12278 1378 12300
rect 1398 12278 1402 12300
rect 1422 12278 1426 12300
rect 1446 12278 1450 12300
rect 1470 12278 1474 12300
rect 1494 12278 1498 12300
rect 1518 12278 1522 12300
rect 1542 12278 1546 12300
rect 1566 12278 1570 12300
rect 1590 12278 1594 12300
rect 1614 12278 1618 12300
rect 1638 12278 1642 12300
rect 1662 12278 1666 12300
rect 1686 12278 1690 12300
rect 1710 12278 1714 12300
rect 1734 12278 1738 12300
rect 1758 12278 1762 12300
rect 1782 12278 1786 12300
rect 1806 12278 1810 12300
rect 1830 12278 1834 12300
rect 1854 12278 1858 12300
rect 1878 12278 1882 12300
rect 1902 12278 1906 12300
rect 1926 12278 1930 12300
rect 1950 12278 1954 12300
rect 1974 12278 1978 12300
rect 1998 12278 2002 12300
rect 2022 12278 2026 12300
rect 2046 12278 2050 12300
rect 2070 12278 2074 12300
rect 2094 12278 2098 12300
rect 2118 12278 2122 12300
rect 2142 12278 2146 12300
rect 2166 12278 2170 12300
rect 2190 12278 2194 12300
rect 2214 12278 2218 12300
rect 2238 12278 2242 12300
rect 2262 12278 2266 12300
rect 2286 12278 2290 12300
rect 2310 12278 2314 12300
rect 2334 12278 2338 12300
rect 2358 12278 2362 12300
rect 2382 12278 2386 12300
rect 2406 12278 2410 12300
rect 2430 12278 2434 12300
rect 2454 12278 2458 12300
rect 2478 12278 2482 12300
rect 2502 12278 2506 12300
rect 2526 12278 2530 12300
rect 2550 12278 2554 12300
rect 2574 12278 2578 12300
rect 2598 12278 2602 12300
rect 2622 12278 2626 12300
rect 2646 12278 2650 12300
rect 2670 12278 2674 12300
rect 2694 12278 2698 12300
rect 2718 12278 2722 12300
rect 2742 12278 2746 12300
rect 2766 12278 2770 12300
rect 2790 12278 2794 12300
rect 2814 12278 2818 12300
rect 2838 12278 2842 12300
rect 2862 12278 2866 12300
rect 2886 12278 2890 12300
rect 2910 12278 2914 12300
rect 2934 12278 2938 12300
rect 2958 12278 2962 12300
rect 2982 12278 2986 12300
rect 3006 12278 3010 12300
rect 3030 12278 3034 12300
rect 3054 12278 3058 12300
rect 3078 12278 3082 12300
rect 3102 12278 3106 12300
rect 3126 12278 3130 12300
rect 3150 12278 3154 12300
rect 3163 12293 3168 12300
rect 3174 12293 3178 12300
rect 3173 12279 3178 12293
rect 3198 12278 3202 12420
rect 3222 12278 3226 12420
rect 3246 12278 3250 12420
rect 3270 12278 3274 12420
rect 3283 12365 3288 12375
rect 3294 12365 3298 12420
rect 3307 12389 3312 12399
rect 3318 12389 3322 12420
rect 3331 12413 3336 12420
rect 3342 12413 3346 12420
rect 3341 12399 3346 12413
rect 3317 12375 3322 12389
rect 3293 12351 3298 12365
rect 3283 12341 3288 12351
rect 3293 12327 3298 12341
rect 3294 12279 3298 12327
rect 3283 12278 3315 12279
rect -1067 12276 3315 12278
rect -1067 12275 -1053 12276
rect -1050 12275 -1043 12276
rect -1050 12254 -1046 12275
rect -1026 12254 -1022 12276
rect -1002 12254 -998 12276
rect -978 12254 -974 12276
rect -954 12254 -950 12276
rect -930 12254 -926 12276
rect -906 12254 -902 12276
rect -882 12254 -878 12276
rect -858 12254 -854 12276
rect -834 12254 -830 12276
rect -810 12254 -806 12276
rect -786 12254 -782 12276
rect -762 12254 -758 12276
rect -738 12254 -734 12276
rect -714 12254 -710 12276
rect -690 12254 -686 12276
rect -666 12254 -662 12276
rect -642 12254 -638 12276
rect -618 12254 -614 12276
rect -594 12254 -590 12276
rect -570 12254 -566 12276
rect -546 12254 -542 12276
rect -522 12254 -518 12276
rect -498 12254 -494 12276
rect -474 12254 -470 12276
rect -450 12254 -446 12276
rect -426 12254 -422 12276
rect -402 12254 -398 12276
rect -378 12254 -374 12276
rect -354 12254 -350 12276
rect -330 12254 -326 12276
rect -306 12254 -302 12276
rect -282 12254 -278 12276
rect -258 12254 -254 12276
rect -234 12254 -230 12276
rect -210 12254 -206 12276
rect -186 12254 -182 12276
rect -162 12254 -158 12276
rect -138 12254 -134 12276
rect -114 12254 -110 12276
rect -90 12254 -86 12276
rect -66 12254 -62 12276
rect -42 12254 -38 12276
rect -18 12254 -14 12276
rect 6 12254 10 12276
rect 30 12254 34 12276
rect 54 12254 58 12276
rect 78 12254 82 12276
rect 102 12254 106 12276
rect 126 12254 130 12276
rect 150 12254 154 12276
rect 174 12254 178 12276
rect 198 12254 202 12276
rect 222 12254 226 12276
rect 246 12254 250 12276
rect 270 12254 274 12276
rect 294 12254 298 12276
rect 318 12254 322 12276
rect 342 12254 346 12276
rect 366 12254 370 12276
rect 390 12254 394 12276
rect 414 12254 418 12276
rect 438 12254 442 12276
rect 462 12254 466 12276
rect 486 12254 490 12276
rect 510 12254 514 12276
rect 534 12254 538 12276
rect 558 12254 562 12276
rect 582 12254 586 12276
rect 606 12254 610 12276
rect 630 12254 634 12276
rect 654 12254 658 12276
rect 678 12254 682 12276
rect 702 12254 706 12276
rect 726 12254 730 12276
rect 750 12254 754 12276
rect 774 12254 778 12276
rect 798 12254 802 12276
rect 822 12254 826 12276
rect 846 12254 850 12276
rect 870 12254 874 12276
rect 894 12254 898 12276
rect 918 12254 922 12276
rect 942 12254 946 12276
rect 966 12254 970 12276
rect 990 12254 994 12276
rect 1014 12254 1018 12276
rect 1038 12254 1042 12276
rect 1062 12254 1066 12276
rect 1086 12254 1090 12276
rect 1110 12254 1114 12276
rect 1134 12254 1138 12276
rect 1158 12254 1162 12276
rect 1182 12254 1186 12276
rect 1206 12254 1210 12276
rect 1230 12254 1234 12276
rect 1254 12254 1258 12276
rect 1278 12254 1282 12276
rect 1302 12254 1306 12276
rect 1326 12254 1330 12276
rect 1350 12254 1354 12276
rect 1374 12254 1378 12276
rect 1398 12254 1402 12276
rect 1422 12254 1426 12276
rect 1446 12254 1450 12276
rect 1470 12254 1474 12276
rect 1494 12254 1498 12276
rect 1518 12254 1522 12276
rect 1542 12254 1546 12276
rect 1566 12254 1570 12276
rect 1590 12254 1594 12276
rect 1614 12254 1618 12276
rect 1638 12254 1642 12276
rect 1662 12254 1666 12276
rect 1686 12254 1690 12276
rect 1710 12254 1714 12276
rect 1734 12254 1738 12276
rect 1758 12254 1762 12276
rect 1782 12254 1786 12276
rect 1806 12254 1810 12276
rect 1830 12254 1834 12276
rect 1854 12254 1858 12276
rect 1878 12254 1882 12276
rect 1902 12254 1906 12276
rect 1926 12254 1930 12276
rect 1950 12254 1954 12276
rect 1974 12254 1978 12276
rect 1998 12254 2002 12276
rect 2022 12254 2026 12276
rect 2046 12254 2050 12276
rect 2070 12254 2074 12276
rect 2094 12254 2098 12276
rect 2118 12254 2122 12276
rect 2142 12254 2146 12276
rect 2166 12254 2170 12276
rect 2190 12254 2194 12276
rect 2214 12254 2218 12276
rect 2238 12254 2242 12276
rect 2262 12254 2266 12276
rect 2286 12254 2290 12276
rect 2310 12254 2314 12276
rect 2334 12254 2338 12276
rect 2358 12254 2362 12276
rect 2382 12254 2386 12276
rect 2406 12254 2410 12276
rect 2430 12254 2434 12276
rect 2454 12254 2458 12276
rect 2478 12254 2482 12276
rect 2502 12254 2506 12276
rect 2526 12254 2530 12276
rect 2550 12254 2554 12276
rect 2574 12254 2578 12276
rect 2598 12254 2602 12276
rect 2622 12254 2626 12276
rect 2646 12254 2650 12276
rect 2670 12254 2674 12276
rect 2694 12254 2698 12276
rect 2718 12254 2722 12276
rect 2742 12254 2746 12276
rect 2766 12254 2770 12276
rect 2790 12254 2794 12276
rect 2814 12254 2818 12276
rect 2838 12254 2842 12276
rect 2862 12254 2866 12276
rect 2886 12254 2890 12276
rect 2910 12254 2914 12276
rect 2934 12254 2938 12276
rect 2958 12254 2962 12276
rect 2982 12254 2986 12276
rect 3006 12254 3010 12276
rect 3030 12254 3034 12276
rect 3054 12254 3058 12276
rect 3078 12254 3082 12276
rect 3102 12254 3106 12276
rect 3126 12254 3130 12276
rect 3150 12254 3154 12276
rect 3163 12254 3197 12255
rect -2393 12252 3197 12254
rect -2371 12230 -2366 12252
rect -2348 12230 -2343 12252
rect -2325 12230 -2320 12252
rect -2072 12250 -2036 12251
rect -2072 12244 -2054 12250
rect -2309 12236 -2301 12244
rect -2317 12230 -2309 12236
rect -2092 12235 -2062 12240
rect -2000 12231 -1992 12252
rect -1938 12251 -1906 12252
rect -1920 12250 -1906 12251
rect -1806 12244 -1680 12250
rect -1854 12235 -1806 12240
rect -1655 12236 -1647 12244
rect -1982 12231 -1966 12232
rect -2000 12230 -1966 12231
rect -1846 12230 -1806 12233
rect -1663 12230 -1655 12236
rect -1642 12230 -1637 12252
rect -1619 12230 -1614 12252
rect -1530 12230 -1526 12252
rect -1506 12230 -1502 12252
rect -1482 12230 -1478 12252
rect -1458 12230 -1454 12252
rect -1434 12230 -1430 12252
rect -1410 12230 -1406 12252
rect -1386 12230 -1382 12252
rect -1362 12230 -1358 12252
rect -1338 12230 -1334 12252
rect -1314 12251 -1310 12252
rect -2393 12228 -1317 12230
rect -2371 12206 -2366 12228
rect -2348 12206 -2343 12228
rect -2325 12206 -2320 12228
rect -2000 12226 -1966 12228
rect -2309 12208 -2301 12216
rect -2062 12215 -2054 12222
rect -2092 12208 -2084 12215
rect -2062 12208 -2026 12210
rect -2317 12206 -2309 12208
rect -2062 12206 -2012 12208
rect -2000 12206 -1992 12226
rect -1982 12225 -1966 12226
rect -1846 12224 -1806 12228
rect -1846 12217 -1798 12222
rect -1806 12215 -1798 12217
rect -1854 12213 -1846 12215
rect -1854 12208 -1806 12213
rect -1655 12208 -1647 12216
rect -1864 12206 -1796 12207
rect -1663 12206 -1655 12208
rect -1642 12206 -1637 12228
rect -1619 12206 -1614 12228
rect -1530 12206 -1526 12228
rect -1506 12206 -1502 12228
rect -1482 12206 -1478 12228
rect -1458 12206 -1454 12228
rect -1434 12206 -1430 12228
rect -1410 12206 -1406 12228
rect -1386 12206 -1382 12228
rect -1362 12206 -1358 12228
rect -1338 12206 -1334 12228
rect -1331 12227 -1317 12228
rect -1314 12227 -1307 12251
rect -1290 12206 -1286 12252
rect -1266 12206 -1262 12252
rect -1242 12206 -1238 12252
rect -1218 12206 -1214 12252
rect -1194 12206 -1190 12252
rect -1170 12206 -1166 12252
rect -1146 12206 -1142 12252
rect -1122 12206 -1118 12252
rect -1098 12206 -1094 12252
rect -1074 12206 -1070 12252
rect -1050 12206 -1046 12252
rect -1026 12206 -1022 12252
rect -1002 12206 -998 12252
rect -978 12206 -974 12252
rect -954 12206 -950 12252
rect -930 12206 -926 12252
rect -906 12206 -902 12252
rect -882 12206 -878 12252
rect -858 12206 -854 12252
rect -834 12206 -830 12252
rect -810 12206 -806 12252
rect -786 12206 -782 12252
rect -762 12206 -758 12252
rect -738 12206 -734 12252
rect -714 12206 -710 12252
rect -690 12206 -686 12252
rect -666 12206 -662 12252
rect -642 12207 -638 12252
rect -653 12206 -619 12207
rect -2393 12204 -619 12206
rect -2371 12158 -2366 12204
rect -2348 12158 -2343 12204
rect -2325 12168 -2320 12204
rect -2317 12200 -2309 12204
rect -2062 12200 -2054 12204
rect -2154 12196 -2138 12198
rect -2057 12196 -2054 12200
rect -2292 12190 -2054 12196
rect -2052 12190 -2044 12200
rect -2092 12174 -2062 12176
rect -2094 12170 -2062 12174
rect -2325 12158 -2317 12168
rect -2095 12160 -2084 12164
rect -2000 12161 -1992 12204
rect -1846 12197 -1806 12204
rect -1663 12200 -1655 12204
rect -1846 12190 -1680 12196
rect -1854 12174 -1806 12176
rect -1854 12170 -1680 12174
rect -2119 12158 -2069 12160
rect -2054 12158 -1892 12161
rect -1671 12158 -1663 12168
rect -1642 12158 -1637 12204
rect -1619 12158 -1614 12204
rect -1530 12158 -1526 12204
rect -1506 12158 -1502 12204
rect -1482 12158 -1478 12204
rect -1458 12158 -1454 12204
rect -1434 12158 -1430 12204
rect -1410 12158 -1406 12204
rect -1386 12158 -1382 12204
rect -1362 12158 -1358 12204
rect -1338 12158 -1334 12204
rect -1314 12179 -1307 12203
rect -1314 12158 -1310 12179
rect -1290 12158 -1286 12204
rect -1266 12158 -1262 12204
rect -1242 12158 -1238 12204
rect -1218 12158 -1214 12204
rect -1194 12158 -1190 12204
rect -1170 12158 -1166 12204
rect -1146 12158 -1142 12204
rect -1122 12158 -1118 12204
rect -1098 12158 -1094 12204
rect -1074 12158 -1070 12204
rect -1050 12158 -1046 12204
rect -1026 12158 -1022 12204
rect -1002 12158 -998 12204
rect -978 12158 -974 12204
rect -954 12158 -950 12204
rect -930 12158 -926 12204
rect -906 12158 -902 12204
rect -882 12158 -878 12204
rect -858 12158 -854 12204
rect -834 12158 -830 12204
rect -810 12158 -806 12204
rect -786 12158 -782 12204
rect -762 12158 -758 12204
rect -738 12158 -734 12204
rect -714 12158 -710 12204
rect -690 12158 -686 12204
rect -666 12158 -662 12204
rect -653 12197 -648 12204
rect -642 12197 -638 12204
rect -643 12183 -638 12197
rect -642 12158 -638 12183
rect -618 12158 -614 12252
rect -594 12158 -590 12252
rect -570 12158 -566 12252
rect -546 12158 -542 12252
rect -522 12158 -518 12252
rect -498 12158 -494 12252
rect -474 12158 -470 12252
rect -450 12158 -446 12252
rect -426 12158 -422 12252
rect -402 12158 -398 12252
rect -378 12158 -374 12252
rect -354 12158 -350 12252
rect -330 12158 -326 12252
rect -306 12158 -302 12252
rect -282 12158 -278 12252
rect -258 12158 -254 12252
rect -234 12158 -230 12252
rect -210 12158 -206 12252
rect -186 12158 -182 12252
rect -162 12158 -158 12252
rect -138 12158 -134 12252
rect -114 12158 -110 12252
rect -90 12158 -86 12252
rect -66 12158 -62 12252
rect -42 12158 -38 12252
rect -18 12158 -14 12252
rect 6 12158 10 12252
rect 30 12158 34 12252
rect 54 12158 58 12252
rect 78 12158 82 12252
rect 102 12158 106 12252
rect 126 12158 130 12252
rect 150 12158 154 12252
rect 174 12158 178 12252
rect 198 12158 202 12252
rect 222 12158 226 12252
rect 246 12158 250 12252
rect 270 12158 274 12252
rect 294 12158 298 12252
rect 318 12158 322 12252
rect 342 12158 346 12252
rect 366 12158 370 12252
rect 390 12158 394 12252
rect 414 12158 418 12252
rect 427 12221 432 12231
rect 438 12221 442 12252
rect 437 12207 442 12221
rect 427 12206 461 12207
rect 462 12206 466 12252
rect 486 12206 490 12252
rect 510 12206 514 12252
rect 534 12206 538 12252
rect 558 12206 562 12252
rect 582 12206 586 12252
rect 606 12206 610 12252
rect 630 12206 634 12252
rect 654 12206 658 12252
rect 678 12206 682 12252
rect 702 12206 706 12252
rect 726 12206 730 12252
rect 750 12206 754 12252
rect 774 12206 778 12252
rect 798 12206 802 12252
rect 822 12206 826 12252
rect 846 12206 850 12252
rect 870 12206 874 12252
rect 894 12206 898 12252
rect 918 12206 922 12252
rect 942 12206 946 12252
rect 966 12206 970 12252
rect 990 12206 994 12252
rect 1014 12206 1018 12252
rect 1038 12206 1042 12252
rect 1062 12206 1066 12252
rect 1086 12206 1090 12252
rect 1110 12206 1114 12252
rect 1134 12206 1138 12252
rect 1158 12206 1162 12252
rect 1182 12206 1186 12252
rect 1206 12206 1210 12252
rect 1230 12206 1234 12252
rect 1254 12206 1258 12252
rect 1278 12206 1282 12252
rect 1302 12206 1306 12252
rect 1326 12206 1330 12252
rect 1350 12206 1354 12252
rect 1374 12206 1378 12252
rect 1398 12206 1402 12252
rect 1422 12206 1426 12252
rect 1446 12206 1450 12252
rect 1470 12206 1474 12252
rect 1494 12206 1498 12252
rect 1518 12206 1522 12252
rect 1542 12206 1546 12252
rect 1566 12206 1570 12252
rect 1590 12206 1594 12252
rect 1614 12206 1618 12252
rect 1638 12206 1642 12252
rect 1662 12206 1666 12252
rect 1686 12206 1690 12252
rect 1710 12206 1714 12252
rect 1734 12206 1738 12252
rect 1758 12206 1762 12252
rect 1782 12206 1786 12252
rect 1806 12206 1810 12252
rect 1830 12206 1834 12252
rect 1854 12206 1858 12252
rect 1878 12206 1882 12252
rect 1902 12206 1906 12252
rect 1926 12206 1930 12252
rect 1950 12206 1954 12252
rect 1974 12206 1978 12252
rect 1998 12206 2002 12252
rect 2022 12206 2026 12252
rect 2046 12206 2050 12252
rect 2070 12206 2074 12252
rect 2094 12206 2098 12252
rect 2118 12206 2122 12252
rect 2142 12206 2146 12252
rect 2166 12206 2170 12252
rect 2190 12206 2194 12252
rect 2214 12206 2218 12252
rect 2238 12206 2242 12252
rect 2262 12206 2266 12252
rect 2286 12206 2290 12252
rect 2310 12206 2314 12252
rect 2334 12206 2338 12252
rect 2358 12206 2362 12252
rect 2382 12206 2386 12252
rect 2406 12206 2410 12252
rect 2430 12206 2434 12252
rect 2454 12206 2458 12252
rect 2478 12206 2482 12252
rect 2502 12206 2506 12252
rect 2526 12206 2530 12252
rect 2550 12206 2554 12252
rect 2574 12206 2578 12252
rect 2598 12206 2602 12252
rect 2622 12206 2626 12252
rect 2646 12206 2650 12252
rect 2670 12206 2674 12252
rect 2694 12206 2698 12252
rect 2718 12206 2722 12252
rect 2742 12206 2746 12252
rect 2766 12206 2770 12252
rect 2790 12206 2794 12252
rect 2814 12206 2818 12252
rect 2838 12206 2842 12252
rect 2862 12206 2866 12252
rect 2886 12206 2890 12252
rect 2910 12206 2914 12252
rect 2934 12206 2938 12252
rect 2958 12206 2962 12252
rect 2982 12206 2986 12252
rect 3006 12206 3010 12252
rect 3030 12206 3034 12252
rect 3054 12206 3058 12252
rect 3078 12206 3082 12252
rect 3102 12206 3106 12252
rect 3126 12206 3130 12252
rect 3150 12206 3154 12252
rect 3163 12245 3168 12252
rect 3173 12231 3178 12245
rect 3174 12206 3178 12231
rect 3198 12227 3202 12276
rect 427 12204 3195 12206
rect 427 12197 432 12204
rect 437 12183 442 12197
rect 438 12158 442 12183
rect 462 12158 466 12204
rect 486 12158 490 12204
rect 510 12158 514 12204
rect 534 12158 538 12204
rect 558 12158 562 12204
rect 582 12158 586 12204
rect 606 12158 610 12204
rect 630 12158 634 12204
rect 654 12158 658 12204
rect 678 12158 682 12204
rect 702 12158 706 12204
rect 726 12158 730 12204
rect 750 12158 754 12204
rect 774 12158 778 12204
rect 798 12158 802 12204
rect 822 12158 826 12204
rect 846 12158 850 12204
rect 870 12158 874 12204
rect 894 12158 898 12204
rect 918 12158 922 12204
rect 942 12158 946 12204
rect 966 12158 970 12204
rect 990 12158 994 12204
rect 1014 12158 1018 12204
rect 1038 12158 1042 12204
rect 1062 12158 1066 12204
rect 1086 12158 1090 12204
rect 1110 12158 1114 12204
rect 1134 12158 1138 12204
rect 1158 12158 1162 12204
rect 1182 12158 1186 12204
rect 1206 12158 1210 12204
rect 1230 12158 1234 12204
rect 1254 12158 1258 12204
rect 1278 12158 1282 12204
rect 1302 12158 1306 12204
rect 1326 12158 1330 12204
rect 1350 12158 1354 12204
rect 1374 12158 1378 12204
rect 1398 12158 1402 12204
rect 1422 12158 1426 12204
rect 1446 12158 1450 12204
rect 1470 12158 1474 12204
rect 1494 12158 1498 12204
rect 1518 12158 1522 12204
rect 1542 12158 1546 12204
rect 1566 12158 1570 12204
rect 1590 12158 1594 12204
rect 1614 12158 1618 12204
rect 1638 12158 1642 12204
rect 1662 12158 1666 12204
rect 1686 12158 1690 12204
rect 1710 12158 1714 12204
rect 1734 12158 1738 12204
rect 1758 12158 1762 12204
rect 1782 12158 1786 12204
rect 1806 12158 1810 12204
rect 1830 12158 1834 12204
rect 1854 12158 1858 12204
rect 1878 12158 1882 12204
rect 1902 12158 1906 12204
rect 1926 12158 1930 12204
rect 1950 12158 1954 12204
rect 1974 12158 1978 12204
rect 1998 12158 2002 12204
rect 2022 12158 2026 12204
rect 2046 12158 2050 12204
rect 2070 12158 2074 12204
rect 2094 12158 2098 12204
rect 2118 12158 2122 12204
rect 2142 12158 2146 12204
rect 2166 12158 2170 12204
rect 2190 12158 2194 12204
rect 2214 12158 2218 12204
rect 2238 12158 2242 12204
rect 2262 12158 2266 12204
rect 2286 12158 2290 12204
rect 2310 12158 2314 12204
rect 2334 12158 2338 12204
rect 2358 12158 2362 12204
rect 2382 12158 2386 12204
rect 2406 12158 2410 12204
rect 2430 12158 2434 12204
rect 2454 12158 2458 12204
rect 2478 12158 2482 12204
rect 2502 12158 2506 12204
rect 2526 12158 2530 12204
rect 2550 12158 2554 12204
rect 2574 12158 2578 12204
rect 2598 12158 2602 12204
rect 2622 12158 2626 12204
rect 2646 12158 2650 12204
rect 2670 12158 2674 12204
rect 2694 12158 2698 12204
rect 2718 12158 2722 12204
rect 2742 12158 2746 12204
rect 2766 12158 2770 12204
rect 2790 12158 2794 12204
rect 2814 12158 2818 12204
rect 2838 12158 2842 12204
rect 2862 12158 2866 12204
rect 2886 12158 2890 12204
rect 2910 12158 2914 12204
rect 2934 12158 2938 12204
rect 2958 12158 2962 12204
rect 2982 12158 2986 12204
rect 3006 12158 3010 12204
rect 3030 12158 3034 12204
rect 3054 12158 3058 12204
rect 3078 12158 3082 12204
rect 3102 12158 3106 12204
rect 3126 12158 3130 12204
rect 3150 12158 3154 12204
rect 3174 12158 3178 12204
rect 3181 12203 3195 12204
rect 3198 12203 3205 12227
rect -2393 12156 3195 12158
rect -2371 12134 -2366 12156
rect -2348 12134 -2343 12156
rect -2325 12152 -2317 12156
rect -2325 12136 -2320 12152
rect -2309 12140 -2301 12152
rect -2095 12150 -2084 12156
rect -2054 12155 -1906 12156
rect -2054 12154 -2036 12155
rect -2084 12148 -2079 12150
rect -2317 12136 -2309 12140
rect -2092 12139 -2079 12146
rect -2000 12142 -1992 12155
rect -1920 12154 -1906 12155
rect -1671 12152 -1663 12156
rect -1846 12148 -1806 12150
rect -1854 12142 -1806 12146
rect -2054 12139 -1982 12142
rect -1966 12139 -1806 12142
rect -1655 12140 -1647 12152
rect -2003 12136 -1992 12139
rect -1904 12137 -1902 12139
rect -1854 12137 -1846 12139
rect -2325 12134 -2317 12136
rect -2033 12134 -1992 12136
rect -1854 12135 -1806 12137
rect -1663 12136 -1655 12140
rect -1864 12134 -1796 12135
rect -1671 12134 -1663 12136
rect -1642 12134 -1637 12156
rect -1619 12134 -1614 12156
rect -1530 12134 -1526 12156
rect -1506 12134 -1502 12156
rect -1482 12134 -1478 12156
rect -1458 12134 -1454 12156
rect -1434 12134 -1430 12156
rect -1410 12134 -1406 12156
rect -1386 12134 -1382 12156
rect -1362 12134 -1358 12156
rect -1338 12134 -1334 12156
rect -1314 12134 -1310 12156
rect -1290 12134 -1286 12156
rect -1266 12134 -1262 12156
rect -1242 12134 -1238 12156
rect -1218 12134 -1214 12156
rect -1194 12134 -1190 12156
rect -1170 12134 -1166 12156
rect -1146 12134 -1142 12156
rect -1122 12134 -1118 12156
rect -1098 12134 -1094 12156
rect -1074 12134 -1070 12156
rect -1050 12134 -1046 12156
rect -1026 12134 -1022 12156
rect -1002 12134 -998 12156
rect -978 12134 -974 12156
rect -954 12134 -950 12156
rect -930 12134 -926 12156
rect -906 12134 -902 12156
rect -882 12134 -878 12156
rect -858 12134 -854 12156
rect -834 12134 -830 12156
rect -810 12134 -806 12156
rect -786 12134 -782 12156
rect -762 12134 -758 12156
rect -738 12134 -734 12156
rect -714 12134 -710 12156
rect -690 12134 -686 12156
rect -666 12134 -662 12156
rect -642 12134 -638 12156
rect -618 12134 -614 12156
rect -594 12134 -590 12156
rect -570 12134 -566 12156
rect -546 12134 -542 12156
rect -522 12134 -518 12156
rect -498 12134 -494 12156
rect -474 12134 -470 12156
rect -450 12134 -446 12156
rect -426 12134 -422 12156
rect -402 12134 -398 12156
rect -378 12134 -374 12156
rect -354 12134 -350 12156
rect -330 12134 -326 12156
rect -306 12134 -302 12156
rect -282 12134 -278 12156
rect -258 12134 -254 12156
rect -234 12134 -230 12156
rect -210 12134 -206 12156
rect -186 12134 -182 12156
rect -162 12134 -158 12156
rect -138 12134 -134 12156
rect -114 12134 -110 12156
rect -90 12134 -86 12156
rect -66 12134 -62 12156
rect -42 12134 -38 12156
rect -18 12134 -14 12156
rect 6 12134 10 12156
rect 30 12134 34 12156
rect 54 12134 58 12156
rect 78 12134 82 12156
rect 102 12134 106 12156
rect 126 12134 130 12156
rect 150 12134 154 12156
rect 174 12134 178 12156
rect 198 12134 202 12156
rect 222 12134 226 12156
rect 246 12134 250 12156
rect 270 12134 274 12156
rect 294 12134 298 12156
rect 318 12134 322 12156
rect 342 12134 346 12156
rect 366 12134 370 12156
rect 390 12134 394 12156
rect 414 12134 418 12156
rect 438 12134 442 12156
rect 462 12155 466 12156
rect -2393 12132 459 12134
rect -2371 12110 -2366 12132
rect -2348 12110 -2343 12132
rect -2325 12124 -2317 12132
rect -2079 12129 -2018 12132
rect -2003 12131 -1966 12132
rect -2000 12130 -1982 12131
rect -2000 12129 -1992 12130
rect -2084 12125 -2009 12129
rect -2028 12124 -2009 12125
rect -2000 12125 -1854 12129
rect -1846 12125 -1798 12132
rect -2325 12110 -2320 12124
rect -2309 12112 -2301 12124
rect -2028 12122 -2018 12124
rect -2092 12112 -2084 12119
rect -2023 12115 -2014 12122
rect -2000 12115 -1992 12125
rect -1671 12124 -1663 12132
rect -1846 12121 -1806 12123
rect -1854 12115 -1806 12119
rect -2054 12112 -1806 12115
rect -1655 12112 -1647 12124
rect -2317 12110 -2309 12112
rect -2054 12110 -2024 12112
rect -2000 12110 -1992 12112
rect -1663 12110 -1655 12112
rect -1642 12110 -1637 12132
rect -1619 12110 -1614 12132
rect -1530 12110 -1526 12132
rect -1506 12110 -1502 12132
rect -1482 12110 -1478 12132
rect -1458 12110 -1454 12132
rect -1434 12110 -1430 12132
rect -1410 12110 -1406 12132
rect -1386 12110 -1382 12132
rect -1362 12110 -1358 12132
rect -1338 12110 -1334 12132
rect -1314 12110 -1310 12132
rect -1290 12110 -1286 12132
rect -1266 12110 -1262 12132
rect -1242 12110 -1238 12132
rect -1218 12110 -1214 12132
rect -1194 12110 -1190 12132
rect -1170 12110 -1166 12132
rect -1146 12110 -1142 12132
rect -1122 12110 -1118 12132
rect -1098 12110 -1094 12132
rect -1074 12110 -1070 12132
rect -1050 12110 -1046 12132
rect -1026 12110 -1022 12132
rect -1002 12110 -998 12132
rect -978 12110 -974 12132
rect -954 12110 -950 12132
rect -930 12110 -926 12132
rect -906 12110 -902 12132
rect -882 12110 -878 12132
rect -858 12110 -854 12132
rect -834 12110 -830 12132
rect -810 12110 -806 12132
rect -786 12110 -782 12132
rect -762 12110 -758 12132
rect -738 12110 -734 12132
rect -714 12110 -710 12132
rect -690 12110 -686 12132
rect -666 12110 -662 12132
rect -642 12110 -638 12132
rect -618 12131 -614 12132
rect -2393 12108 -2064 12110
rect -2060 12108 -621 12110
rect -2371 12062 -2366 12108
rect -2348 12062 -2343 12108
rect -2325 12096 -2317 12108
rect -2060 12105 -2054 12108
rect -2084 12098 -2054 12105
rect -2050 12102 -2044 12104
rect -2325 12076 -2320 12096
rect -2064 12094 -2054 12098
rect -2325 12068 -2317 12076
rect -2101 12071 -2071 12074
rect -2325 12062 -2320 12068
rect -2317 12062 -2309 12068
rect -2000 12066 -1992 12108
rect -1846 12107 -1806 12108
rect -1846 12098 -1798 12105
rect -1671 12096 -1663 12108
rect -1846 12094 -1806 12096
rect -1854 12080 -1680 12084
rect -1846 12071 -1798 12074
rect -2079 12065 -2043 12066
rect -2007 12065 -1991 12066
rect -2079 12064 -2071 12065
rect -2079 12062 -2029 12064
rect -2011 12062 -1991 12065
rect -1846 12063 -1806 12069
rect -1671 12068 -1663 12076
rect -1864 12062 -1796 12063
rect -1663 12062 -1655 12068
rect -1642 12062 -1637 12108
rect -1619 12062 -1614 12108
rect -1530 12062 -1526 12108
rect -1506 12062 -1502 12108
rect -1482 12062 -1478 12108
rect -1458 12062 -1454 12108
rect -1434 12062 -1430 12108
rect -1410 12062 -1406 12108
rect -1386 12062 -1382 12108
rect -1362 12062 -1358 12108
rect -1338 12062 -1334 12108
rect -1314 12062 -1310 12108
rect -1290 12062 -1286 12108
rect -1266 12062 -1262 12108
rect -1242 12062 -1238 12108
rect -1218 12062 -1214 12108
rect -1194 12062 -1190 12108
rect -1170 12062 -1166 12108
rect -1146 12062 -1142 12108
rect -1122 12062 -1118 12108
rect -1098 12062 -1094 12108
rect -1074 12062 -1070 12108
rect -1050 12062 -1046 12108
rect -1026 12062 -1022 12108
rect -1002 12062 -998 12108
rect -978 12062 -974 12108
rect -954 12062 -950 12108
rect -930 12062 -926 12108
rect -906 12062 -902 12108
rect -882 12062 -878 12108
rect -858 12062 -854 12108
rect -834 12062 -830 12108
rect -810 12062 -806 12108
rect -786 12062 -782 12108
rect -762 12062 -758 12108
rect -738 12062 -734 12108
rect -714 12062 -710 12108
rect -690 12062 -686 12108
rect -666 12062 -662 12108
rect -642 12062 -638 12108
rect -635 12107 -621 12108
rect -618 12107 -611 12131
rect -618 12062 -614 12107
rect -594 12062 -590 12132
rect -570 12062 -566 12132
rect -546 12062 -542 12132
rect -522 12062 -518 12132
rect -498 12062 -494 12132
rect -474 12062 -470 12132
rect -450 12062 -446 12132
rect -426 12062 -422 12132
rect -402 12062 -398 12132
rect -378 12062 -374 12132
rect -354 12062 -350 12132
rect -330 12062 -326 12132
rect -306 12062 -302 12132
rect -282 12062 -278 12132
rect -258 12062 -254 12132
rect -234 12062 -230 12132
rect -210 12062 -206 12132
rect -186 12062 -182 12132
rect -162 12062 -158 12132
rect -138 12062 -134 12132
rect -114 12062 -110 12132
rect -90 12062 -86 12132
rect -66 12062 -62 12132
rect -42 12062 -38 12132
rect -18 12062 -14 12132
rect 6 12062 10 12132
rect 30 12062 34 12132
rect 54 12062 58 12132
rect 78 12062 82 12132
rect 102 12062 106 12132
rect 126 12062 130 12132
rect 150 12062 154 12132
rect 174 12062 178 12132
rect 198 12062 202 12132
rect 222 12062 226 12132
rect 246 12062 250 12132
rect 270 12062 274 12132
rect 294 12062 298 12132
rect 318 12062 322 12132
rect 342 12062 346 12132
rect 366 12062 370 12132
rect 390 12062 394 12132
rect 414 12062 418 12132
rect 438 12062 442 12132
rect 445 12131 459 12132
rect 462 12110 469 12155
rect 486 12110 490 12156
rect 510 12110 514 12156
rect 534 12110 538 12156
rect 558 12110 562 12156
rect 582 12110 586 12156
rect 606 12110 610 12156
rect 630 12110 634 12156
rect 654 12110 658 12156
rect 678 12110 682 12156
rect 702 12110 706 12156
rect 726 12110 730 12156
rect 750 12110 754 12156
rect 774 12110 778 12156
rect 798 12110 802 12156
rect 822 12110 826 12156
rect 835 12125 840 12135
rect 846 12125 850 12156
rect 845 12111 850 12125
rect 846 12110 850 12111
rect 870 12110 874 12156
rect 894 12110 898 12156
rect 918 12110 922 12156
rect 942 12110 946 12156
rect 966 12110 970 12156
rect 990 12110 994 12156
rect 1014 12110 1018 12156
rect 1038 12110 1042 12156
rect 1062 12110 1066 12156
rect 1086 12110 1090 12156
rect 1110 12110 1114 12156
rect 1134 12110 1138 12156
rect 1158 12110 1162 12156
rect 1182 12110 1186 12156
rect 1206 12110 1210 12156
rect 1230 12110 1234 12156
rect 1254 12110 1258 12156
rect 1278 12110 1282 12156
rect 1302 12110 1306 12156
rect 1326 12110 1330 12156
rect 1350 12110 1354 12156
rect 1374 12110 1378 12156
rect 1398 12110 1402 12156
rect 1422 12110 1426 12156
rect 1446 12110 1450 12156
rect 1470 12110 1474 12156
rect 1494 12110 1498 12156
rect 1518 12110 1522 12156
rect 1542 12110 1546 12156
rect 1566 12110 1570 12156
rect 1590 12110 1594 12156
rect 1614 12110 1618 12156
rect 1638 12110 1642 12156
rect 1662 12110 1666 12156
rect 1686 12110 1690 12156
rect 1710 12110 1714 12156
rect 1734 12110 1738 12156
rect 1758 12110 1762 12156
rect 1782 12110 1786 12156
rect 1806 12110 1810 12156
rect 1830 12110 1834 12156
rect 1854 12111 1858 12156
rect 1843 12110 1877 12111
rect 445 12108 1877 12110
rect 445 12107 459 12108
rect 462 12107 469 12108
rect 462 12062 466 12107
rect 486 12062 490 12108
rect 510 12062 514 12108
rect 534 12062 538 12108
rect 558 12062 562 12108
rect 582 12062 586 12108
rect 606 12062 610 12108
rect 630 12062 634 12108
rect 654 12062 658 12108
rect 678 12062 682 12108
rect 702 12062 706 12108
rect 726 12062 730 12108
rect 750 12062 754 12108
rect 774 12062 778 12108
rect 798 12062 802 12108
rect 822 12062 826 12108
rect 846 12062 850 12108
rect 870 12062 874 12108
rect 894 12062 898 12108
rect 918 12062 922 12108
rect 942 12062 946 12108
rect 966 12062 970 12108
rect 990 12062 994 12108
rect 1014 12062 1018 12108
rect 1038 12062 1042 12108
rect 1062 12062 1066 12108
rect 1086 12062 1090 12108
rect 1110 12062 1114 12108
rect 1134 12062 1138 12108
rect 1158 12062 1162 12108
rect 1182 12062 1186 12108
rect 1206 12062 1210 12108
rect 1230 12062 1234 12108
rect 1254 12062 1258 12108
rect 1278 12062 1282 12108
rect 1302 12062 1306 12108
rect 1326 12062 1330 12108
rect 1350 12062 1354 12108
rect 1374 12062 1378 12108
rect 1398 12062 1402 12108
rect 1422 12062 1426 12108
rect 1446 12062 1450 12108
rect 1470 12062 1474 12108
rect 1494 12062 1498 12108
rect 1518 12062 1522 12108
rect 1542 12062 1546 12108
rect 1566 12062 1570 12108
rect 1590 12063 1594 12108
rect 1579 12062 1613 12063
rect -2393 12060 1613 12062
rect -2371 12014 -2366 12060
rect -2348 12014 -2343 12060
rect -2325 12048 -2320 12060
rect -2079 12058 -2071 12060
rect -2072 12056 -2071 12058
rect -2109 12051 -2101 12056
rect -2101 12049 -2079 12051
rect -2069 12049 -2068 12056
rect -2325 12040 -2317 12048
rect -2079 12044 -2071 12049
rect -2325 12020 -2320 12040
rect -2317 12032 -2309 12040
rect -2074 12035 -2071 12044
rect -2069 12040 -2068 12044
rect -2109 12026 -2079 12029
rect -2325 12014 -2317 12020
rect -2000 12014 -1992 12060
rect -1846 12058 -1806 12060
rect -1854 12053 -1806 12057
rect -1854 12051 -1846 12053
rect -1846 12049 -1806 12051
rect -1806 12047 -1798 12049
rect -1846 12044 -1798 12047
rect -1846 12031 -1806 12042
rect -1671 12040 -1663 12048
rect -1663 12032 -1655 12040
rect -1854 12026 -1680 12030
rect -1671 12014 -1663 12020
rect -1642 12014 -1637 12060
rect -1619 12014 -1614 12060
rect -1530 12014 -1526 12060
rect -1506 12014 -1502 12060
rect -1482 12014 -1478 12060
rect -1458 12014 -1454 12060
rect -1434 12014 -1430 12060
rect -1410 12014 -1406 12060
rect -1386 12014 -1382 12060
rect -1362 12014 -1358 12060
rect -1338 12014 -1334 12060
rect -1314 12014 -1310 12060
rect -1290 12014 -1286 12060
rect -1266 12014 -1262 12060
rect -1242 12014 -1238 12060
rect -1218 12014 -1214 12060
rect -1194 12014 -1190 12060
rect -1170 12014 -1166 12060
rect -1146 12014 -1142 12060
rect -1122 12014 -1118 12060
rect -1098 12014 -1094 12060
rect -1074 12014 -1070 12060
rect -1050 12014 -1046 12060
rect -1026 12014 -1022 12060
rect -1002 12014 -998 12060
rect -978 12014 -974 12060
rect -954 12014 -950 12060
rect -930 12014 -926 12060
rect -906 12014 -902 12060
rect -882 12014 -878 12060
rect -858 12014 -854 12060
rect -834 12014 -830 12060
rect -810 12014 -806 12060
rect -786 12014 -782 12060
rect -762 12014 -758 12060
rect -738 12014 -734 12060
rect -714 12014 -710 12060
rect -690 12014 -686 12060
rect -666 12014 -662 12060
rect -642 12014 -638 12060
rect -618 12014 -614 12060
rect -594 12014 -590 12060
rect -570 12014 -566 12060
rect -546 12014 -542 12060
rect -522 12014 -518 12060
rect -498 12014 -494 12060
rect -474 12014 -470 12060
rect -450 12014 -446 12060
rect -426 12014 -422 12060
rect -402 12014 -398 12060
rect -378 12014 -374 12060
rect -354 12014 -350 12060
rect -330 12014 -326 12060
rect -306 12014 -302 12060
rect -282 12014 -278 12060
rect -258 12014 -254 12060
rect -234 12014 -230 12060
rect -210 12014 -206 12060
rect -186 12014 -182 12060
rect -162 12014 -158 12060
rect -138 12014 -134 12060
rect -114 12014 -110 12060
rect -90 12014 -86 12060
rect -66 12014 -62 12060
rect -42 12014 -38 12060
rect -18 12014 -14 12060
rect 6 12014 10 12060
rect 30 12014 34 12060
rect 54 12014 58 12060
rect 78 12014 82 12060
rect 102 12014 106 12060
rect 126 12014 130 12060
rect 150 12014 154 12060
rect 174 12014 178 12060
rect 198 12014 202 12060
rect 222 12014 226 12060
rect 246 12014 250 12060
rect 270 12014 274 12060
rect 294 12014 298 12060
rect 318 12014 322 12060
rect 342 12014 346 12060
rect 366 12014 370 12060
rect 390 12014 394 12060
rect 414 12014 418 12060
rect 438 12014 442 12060
rect 462 12014 466 12060
rect 486 12014 490 12060
rect 510 12014 514 12060
rect 534 12014 538 12060
rect 558 12014 562 12060
rect 582 12014 586 12060
rect 606 12014 610 12060
rect 630 12014 634 12060
rect 654 12014 658 12060
rect 678 12014 682 12060
rect 702 12014 706 12060
rect 726 12014 730 12060
rect 750 12014 754 12060
rect 774 12014 778 12060
rect 798 12014 802 12060
rect 822 12014 826 12060
rect 846 12014 850 12060
rect 870 12059 874 12060
rect 870 12035 877 12059
rect 870 12014 874 12035
rect 894 12014 898 12060
rect 918 12014 922 12060
rect 942 12014 946 12060
rect 966 12014 970 12060
rect 990 12014 994 12060
rect 1014 12014 1018 12060
rect 1038 12014 1042 12060
rect 1062 12014 1066 12060
rect 1086 12014 1090 12060
rect 1110 12014 1114 12060
rect 1134 12014 1138 12060
rect 1158 12014 1162 12060
rect 1182 12014 1186 12060
rect 1206 12014 1210 12060
rect 1230 12014 1234 12060
rect 1254 12014 1258 12060
rect 1278 12014 1282 12060
rect 1302 12014 1306 12060
rect 1326 12014 1330 12060
rect 1350 12014 1354 12060
rect 1374 12014 1378 12060
rect 1398 12014 1402 12060
rect 1422 12014 1426 12060
rect 1446 12014 1450 12060
rect 1470 12014 1474 12060
rect 1494 12014 1498 12060
rect 1518 12014 1522 12060
rect 1542 12014 1546 12060
rect 1566 12014 1570 12060
rect 1579 12053 1584 12060
rect 1590 12053 1594 12060
rect 1589 12039 1594 12053
rect 1579 12029 1584 12039
rect 1589 12015 1594 12029
rect 1590 12014 1594 12015
rect 1614 12014 1618 12108
rect 1638 12014 1642 12108
rect 1662 12014 1666 12108
rect 1686 12014 1690 12108
rect 1710 12014 1714 12108
rect 1734 12014 1738 12108
rect 1758 12014 1762 12108
rect 1782 12014 1786 12108
rect 1806 12014 1810 12108
rect 1830 12014 1834 12108
rect 1843 12101 1848 12108
rect 1854 12101 1858 12108
rect 1853 12087 1858 12101
rect 1843 12062 1877 12063
rect 1878 12062 1882 12156
rect 1902 12062 1906 12156
rect 1926 12062 1930 12156
rect 1950 12062 1954 12156
rect 1974 12062 1978 12156
rect 1998 12062 2002 12156
rect 2022 12062 2026 12156
rect 2046 12062 2050 12156
rect 2070 12062 2074 12156
rect 2094 12062 2098 12156
rect 2118 12062 2122 12156
rect 2142 12062 2146 12156
rect 2166 12062 2170 12156
rect 2190 12062 2194 12156
rect 2214 12062 2218 12156
rect 2238 12062 2242 12156
rect 2262 12062 2266 12156
rect 2286 12062 2290 12156
rect 2310 12062 2314 12156
rect 2334 12062 2338 12156
rect 2358 12062 2362 12156
rect 2382 12062 2386 12156
rect 2406 12062 2410 12156
rect 2430 12062 2434 12156
rect 2454 12062 2458 12156
rect 2478 12062 2482 12156
rect 2491 12077 2496 12087
rect 2502 12077 2506 12156
rect 2501 12063 2506 12077
rect 2526 12062 2530 12156
rect 2550 12062 2554 12156
rect 2574 12062 2578 12156
rect 2598 12062 2602 12156
rect 2622 12062 2626 12156
rect 2646 12062 2650 12156
rect 2670 12062 2674 12156
rect 2694 12062 2698 12156
rect 2718 12062 2722 12156
rect 2742 12062 2746 12156
rect 2766 12062 2770 12156
rect 2790 12062 2794 12156
rect 2814 12062 2818 12156
rect 2838 12062 2842 12156
rect 2862 12062 2866 12156
rect 2886 12062 2890 12156
rect 2910 12062 2914 12156
rect 2934 12062 2938 12156
rect 2958 12062 2962 12156
rect 2982 12062 2986 12156
rect 3006 12062 3010 12156
rect 3030 12062 3034 12156
rect 3054 12062 3058 12156
rect 3078 12062 3082 12156
rect 3102 12062 3106 12156
rect 3126 12062 3130 12156
rect 3150 12062 3154 12156
rect 3174 12062 3178 12156
rect 3181 12155 3195 12156
rect 3198 12155 3205 12179
rect 3198 12062 3202 12155
rect 3222 12062 3226 12276
rect 3246 12062 3250 12276
rect 3259 12197 3264 12207
rect 3270 12197 3274 12276
rect 3283 12269 3288 12276
rect 3294 12269 3298 12276
rect 3301 12275 3315 12276
rect 3293 12255 3298 12269
rect 3307 12265 3315 12269
rect 3301 12255 3307 12265
rect 3269 12183 3274 12197
rect 3259 12149 3264 12159
rect 3269 12135 3274 12149
rect 3270 12063 3274 12135
rect 3259 12062 3291 12063
rect 1843 12060 3291 12062
rect 1843 12053 1848 12060
rect 1853 12039 1858 12053
rect 1854 12014 1858 12039
rect 1878 12035 1882 12060
rect -2393 12012 1875 12014
rect -2371 11990 -2366 12012
rect -2348 11990 -2343 12012
rect -2325 12004 -2317 12012
rect -2325 11990 -2320 12004
rect -2309 11992 -2301 12004
rect -2092 11995 -2062 12000
rect -2000 11992 -1992 12012
rect -2317 11990 -2309 11992
rect -2000 11990 -1983 11992
rect -1906 11990 -1904 12012
rect -1806 12004 -1680 12010
rect -1671 12004 -1663 12012
rect -1854 11995 -1806 12000
rect -1846 11990 -1806 11993
rect -1655 11992 -1647 12004
rect -1663 11990 -1655 11992
rect -1642 11990 -1637 12012
rect -1619 11990 -1614 12012
rect -1530 11990 -1526 12012
rect -1506 11990 -1502 12012
rect -1482 11990 -1478 12012
rect -1458 11990 -1454 12012
rect -1434 11990 -1430 12012
rect -1410 11990 -1406 12012
rect -1386 11990 -1382 12012
rect -1362 11990 -1358 12012
rect -1338 11990 -1334 12012
rect -1314 11990 -1310 12012
rect -1290 11990 -1286 12012
rect -1266 11990 -1262 12012
rect -1242 11990 -1238 12012
rect -1218 11990 -1214 12012
rect -1194 11990 -1190 12012
rect -1170 11990 -1166 12012
rect -1146 11990 -1142 12012
rect -1122 11990 -1118 12012
rect -1098 11990 -1094 12012
rect -1074 11990 -1070 12012
rect -1050 11990 -1046 12012
rect -1026 11990 -1022 12012
rect -1002 11990 -998 12012
rect -978 11990 -974 12012
rect -954 11990 -950 12012
rect -930 11990 -926 12012
rect -906 11990 -902 12012
rect -882 11990 -878 12012
rect -858 11990 -854 12012
rect -834 11990 -830 12012
rect -810 11990 -806 12012
rect -786 11990 -782 12012
rect -762 11990 -758 12012
rect -738 11990 -734 12012
rect -714 11990 -710 12012
rect -690 11990 -686 12012
rect -666 11990 -662 12012
rect -642 11990 -638 12012
rect -618 11990 -614 12012
rect -594 11990 -590 12012
rect -570 11990 -566 12012
rect -546 11990 -542 12012
rect -522 11990 -518 12012
rect -498 11990 -494 12012
rect -474 11990 -470 12012
rect -450 11990 -446 12012
rect -426 11990 -422 12012
rect -402 11990 -398 12012
rect -378 11990 -374 12012
rect -354 11990 -350 12012
rect -330 11990 -326 12012
rect -306 11990 -302 12012
rect -282 11990 -278 12012
rect -258 11990 -254 12012
rect -234 11990 -230 12012
rect -210 11990 -206 12012
rect -186 11990 -182 12012
rect -162 11990 -158 12012
rect -138 11990 -134 12012
rect -114 11990 -110 12012
rect -90 11990 -86 12012
rect -66 11990 -62 12012
rect -42 11990 -38 12012
rect -18 11990 -14 12012
rect 6 11990 10 12012
rect 30 11990 34 12012
rect 54 11990 58 12012
rect 78 11990 82 12012
rect 102 11990 106 12012
rect 126 11990 130 12012
rect 150 11990 154 12012
rect 174 11990 178 12012
rect 198 11990 202 12012
rect 222 11990 226 12012
rect 246 11990 250 12012
rect 270 11990 274 12012
rect 294 11990 298 12012
rect 318 11990 322 12012
rect 342 11990 346 12012
rect 366 11990 370 12012
rect 390 11990 394 12012
rect 414 11990 418 12012
rect 438 11990 442 12012
rect 462 11991 466 12012
rect 451 11990 485 11991
rect -2393 11988 485 11990
rect -2371 11966 -2366 11988
rect -2348 11966 -2343 11988
rect -2325 11976 -2317 11988
rect -2071 11984 -2062 11988
rect -2013 11986 -1983 11988
rect -2000 11985 -1983 11986
rect -2325 11966 -2320 11976
rect -2309 11966 -2301 11976
rect -2100 11975 -2092 11982
rect -2064 11980 -2062 11983
rect -2061 11975 -2059 11980
rect -2071 11970 -2062 11975
rect -2071 11968 -2026 11970
rect -2066 11966 -2012 11968
rect -2000 11966 -1992 11985
rect -1906 11983 -1904 11988
rect -1846 11984 -1806 11988
rect -1846 11977 -1798 11982
rect -1806 11975 -1798 11977
rect -1671 11976 -1663 11988
rect -1854 11973 -1846 11975
rect -1854 11968 -1806 11973
rect -1864 11966 -1796 11967
rect -1655 11966 -1647 11976
rect -1642 11966 -1637 11988
rect -1619 11966 -1614 11988
rect -1530 11966 -1526 11988
rect -1506 11966 -1502 11988
rect -1482 11966 -1478 11988
rect -1458 11966 -1454 11988
rect -1434 11966 -1430 11988
rect -1410 11966 -1406 11988
rect -1386 11966 -1382 11988
rect -1362 11966 -1358 11988
rect -1338 11966 -1334 11988
rect -1314 11966 -1310 11988
rect -1290 11966 -1286 11988
rect -1266 11966 -1262 11988
rect -1242 11966 -1238 11988
rect -1218 11966 -1214 11988
rect -1194 11966 -1190 11988
rect -1170 11966 -1166 11988
rect -1146 11966 -1142 11988
rect -1122 11966 -1118 11988
rect -1098 11966 -1094 11988
rect -1074 11966 -1070 11988
rect -1050 11966 -1046 11988
rect -1026 11966 -1022 11988
rect -1002 11966 -998 11988
rect -978 11966 -974 11988
rect -954 11966 -950 11988
rect -930 11966 -926 11988
rect -906 11966 -902 11988
rect -882 11966 -878 11988
rect -858 11966 -854 11988
rect -834 11966 -830 11988
rect -810 11966 -806 11988
rect -786 11966 -782 11988
rect -762 11966 -758 11988
rect -738 11966 -734 11988
rect -714 11966 -710 11988
rect -690 11966 -686 11988
rect -666 11966 -662 11988
rect -642 11966 -638 11988
rect -618 11966 -614 11988
rect -594 11966 -590 11988
rect -570 11966 -566 11988
rect -546 11966 -542 11988
rect -522 11966 -518 11988
rect -498 11966 -494 11988
rect -474 11966 -470 11988
rect -450 11966 -446 11988
rect -426 11966 -422 11988
rect -402 11966 -398 11988
rect -378 11966 -374 11988
rect -354 11966 -350 11988
rect -330 11966 -326 11988
rect -306 11966 -302 11988
rect -282 11966 -278 11988
rect -258 11966 -254 11988
rect -234 11966 -230 11988
rect -210 11966 -206 11988
rect -186 11966 -182 11988
rect -162 11966 -158 11988
rect -138 11966 -134 11988
rect -114 11966 -110 11988
rect -90 11966 -86 11988
rect -66 11966 -62 11988
rect -42 11966 -38 11988
rect -18 11966 -14 11988
rect 6 11966 10 11988
rect 30 11966 34 11988
rect 54 11966 58 11988
rect 78 11966 82 11988
rect 102 11966 106 11988
rect 126 11966 130 11988
rect 150 11966 154 11988
rect 174 11966 178 11988
rect 198 11966 202 11988
rect 222 11966 226 11988
rect 246 11966 250 11988
rect 270 11966 274 11988
rect 294 11966 298 11988
rect 318 11966 322 11988
rect 342 11966 346 11988
rect 366 11966 370 11988
rect 390 11966 394 11988
rect 414 11966 418 11988
rect 438 11966 442 11988
rect 451 11981 456 11988
rect 462 11981 466 11988
rect 461 11967 466 11981
rect 462 11966 466 11967
rect 486 11966 490 12012
rect 510 11966 514 12012
rect 534 11966 538 12012
rect 558 11966 562 12012
rect 582 11966 586 12012
rect 606 11966 610 12012
rect 630 11966 634 12012
rect 654 11966 658 12012
rect 678 11966 682 12012
rect 702 11966 706 12012
rect 726 11966 730 12012
rect 750 11966 754 12012
rect 774 11966 778 12012
rect 798 11966 802 12012
rect 822 11966 826 12012
rect 846 11966 850 12012
rect 870 11966 874 12012
rect 894 11966 898 12012
rect 918 11966 922 12012
rect 942 11966 946 12012
rect 966 11966 970 12012
rect 990 11966 994 12012
rect 1014 11966 1018 12012
rect 1038 11966 1042 12012
rect 1062 11966 1066 12012
rect 1086 11966 1090 12012
rect 1110 11966 1114 12012
rect 1134 11966 1138 12012
rect 1158 11966 1162 12012
rect 1182 11966 1186 12012
rect 1206 11966 1210 12012
rect 1230 11966 1234 12012
rect 1254 11966 1258 12012
rect 1278 11966 1282 12012
rect 1302 11966 1306 12012
rect 1326 11966 1330 12012
rect 1350 11966 1354 12012
rect 1374 11966 1378 12012
rect 1398 11966 1402 12012
rect 1422 11966 1426 12012
rect 1446 11967 1450 12012
rect 1435 11966 1469 11967
rect -2393 11964 1469 11966
rect -2371 11894 -2366 11964
rect -2348 11894 -2343 11964
rect -2325 11960 -2320 11964
rect -2317 11960 -2309 11964
rect -2325 11948 -2317 11960
rect -2066 11959 -2062 11964
rect -2147 11956 -2134 11958
rect -2292 11950 -2071 11956
rect -2325 11894 -2320 11948
rect -2092 11934 -2062 11936
rect -2094 11930 -2062 11934
rect -2309 11900 -2301 11906
rect -2317 11894 -2309 11900
rect -2000 11894 -1992 11964
rect -1846 11957 -1806 11964
rect -1663 11960 -1655 11964
rect -1846 11950 -1680 11956
rect -1671 11948 -1663 11960
rect -1854 11934 -1806 11936
rect -1854 11930 -1680 11934
rect -1655 11900 -1647 11906
rect -1663 11894 -1655 11900
rect -1642 11894 -1637 11964
rect -1619 11894 -1614 11964
rect -1530 11894 -1526 11964
rect -1506 11894 -1502 11964
rect -1482 11894 -1478 11964
rect -1458 11894 -1454 11964
rect -1434 11894 -1430 11964
rect -1410 11894 -1406 11964
rect -1386 11894 -1382 11964
rect -1362 11894 -1358 11964
rect -1338 11894 -1334 11964
rect -1314 11894 -1310 11964
rect -1290 11894 -1286 11964
rect -1266 11894 -1262 11964
rect -1242 11894 -1238 11964
rect -1218 11894 -1214 11964
rect -1194 11894 -1190 11964
rect -1170 11894 -1166 11964
rect -1146 11894 -1142 11964
rect -1122 11894 -1118 11964
rect -1098 11894 -1094 11964
rect -1074 11894 -1070 11964
rect -1050 11894 -1046 11964
rect -1026 11894 -1022 11964
rect -1002 11894 -998 11964
rect -978 11894 -974 11964
rect -954 11894 -950 11964
rect -930 11894 -926 11964
rect -906 11894 -902 11964
rect -882 11894 -878 11964
rect -858 11894 -854 11964
rect -834 11894 -830 11964
rect -810 11894 -806 11964
rect -786 11894 -782 11964
rect -762 11894 -758 11964
rect -738 11894 -734 11964
rect -714 11894 -710 11964
rect -690 11894 -686 11964
rect -666 11894 -662 11964
rect -642 11894 -638 11964
rect -618 11894 -614 11964
rect -594 11894 -590 11964
rect -570 11894 -566 11964
rect -546 11894 -542 11964
rect -522 11894 -518 11964
rect -498 11894 -494 11964
rect -474 11894 -470 11964
rect -450 11894 -446 11964
rect -426 11894 -422 11964
rect -402 11894 -398 11964
rect -378 11894 -374 11964
rect -354 11894 -350 11964
rect -330 11894 -326 11964
rect -306 11894 -302 11964
rect -282 11894 -278 11964
rect -258 11894 -254 11964
rect -234 11894 -230 11964
rect -210 11894 -206 11964
rect -186 11894 -182 11964
rect -162 11894 -158 11964
rect -138 11894 -134 11964
rect -114 11894 -110 11964
rect -90 11894 -86 11964
rect -66 11894 -62 11964
rect -42 11894 -38 11964
rect -18 11894 -14 11964
rect 6 11894 10 11964
rect 30 11894 34 11964
rect 54 11894 58 11964
rect 78 11894 82 11964
rect 102 11894 106 11964
rect 126 11894 130 11964
rect 150 11894 154 11964
rect 174 11894 178 11964
rect 198 11894 202 11964
rect 222 11894 226 11964
rect 246 11894 250 11964
rect 270 11894 274 11964
rect 294 11894 298 11964
rect 318 11894 322 11964
rect 342 11894 346 11964
rect 366 11894 370 11964
rect 390 11894 394 11964
rect 414 11894 418 11964
rect 438 11894 442 11964
rect 462 11894 466 11964
rect 486 11915 490 11964
rect -2393 11892 483 11894
rect -2371 11798 -2366 11892
rect -2348 11798 -2343 11892
rect -2325 11830 -2320 11892
rect -2317 11890 -2309 11892
rect -2000 11891 -1966 11892
rect -2000 11890 -1982 11891
rect -1663 11890 -1655 11892
rect -2028 11882 -2018 11884
rect -2309 11872 -2301 11878
rect -2091 11872 -2061 11879
rect -2317 11862 -2309 11872
rect -2044 11870 -2028 11872
rect -2026 11870 -2014 11882
rect -2084 11864 -2061 11870
rect -2044 11868 -2014 11870
rect -2292 11854 -2054 11863
rect -2325 11822 -2317 11830
rect -2325 11802 -2320 11822
rect -2317 11814 -2309 11822
rect -2325 11798 -2317 11802
rect -2095 11800 -2083 11804
rect -2000 11801 -1992 11890
rect -1982 11889 -1966 11890
rect -1980 11872 -1932 11879
rect -1655 11872 -1647 11878
rect -1846 11854 -1680 11863
rect -1663 11862 -1655 11872
rect -1671 11822 -1663 11830
rect -1663 11814 -1655 11822
rect -2119 11798 -2069 11800
rect -2053 11798 -1972 11801
rect -1926 11798 -1892 11801
rect -1671 11798 -1663 11802
rect -1642 11798 -1637 11892
rect -1619 11798 -1614 11892
rect -1530 11798 -1526 11892
rect -1506 11798 -1502 11892
rect -1482 11798 -1478 11892
rect -1458 11798 -1454 11892
rect -1434 11798 -1430 11892
rect -1410 11798 -1406 11892
rect -1386 11798 -1382 11892
rect -1362 11798 -1358 11892
rect -1338 11798 -1334 11892
rect -1314 11798 -1310 11892
rect -1290 11798 -1286 11892
rect -1266 11798 -1262 11892
rect -1242 11798 -1238 11892
rect -1218 11798 -1214 11892
rect -1194 11798 -1190 11892
rect -1170 11798 -1166 11892
rect -1146 11798 -1142 11892
rect -1122 11798 -1118 11892
rect -1098 11798 -1094 11892
rect -1074 11798 -1070 11892
rect -1050 11798 -1046 11892
rect -1026 11798 -1022 11892
rect -1002 11798 -998 11892
rect -978 11798 -974 11892
rect -954 11798 -950 11892
rect -930 11798 -926 11892
rect -906 11798 -902 11892
rect -882 11798 -878 11892
rect -858 11798 -854 11892
rect -834 11798 -830 11892
rect -810 11798 -806 11892
rect -786 11798 -782 11892
rect -762 11798 -758 11892
rect -738 11798 -734 11892
rect -714 11798 -710 11892
rect -690 11798 -686 11892
rect -666 11798 -662 11892
rect -642 11798 -638 11892
rect -618 11798 -614 11892
rect -594 11798 -590 11892
rect -570 11798 -566 11892
rect -546 11798 -542 11892
rect -522 11798 -518 11892
rect -498 11798 -494 11892
rect -474 11798 -470 11892
rect -450 11798 -446 11892
rect -426 11798 -422 11892
rect -402 11798 -398 11892
rect -378 11798 -374 11892
rect -354 11798 -350 11892
rect -330 11798 -326 11892
rect -306 11798 -302 11892
rect -282 11798 -278 11892
rect -258 11798 -254 11892
rect -234 11798 -230 11892
rect -210 11798 -206 11892
rect -186 11798 -182 11892
rect -162 11798 -158 11892
rect -138 11798 -134 11892
rect -114 11798 -110 11892
rect -90 11798 -86 11892
rect -66 11798 -62 11892
rect -42 11798 -38 11892
rect -18 11798 -14 11892
rect 6 11798 10 11892
rect 30 11798 34 11892
rect 43 11837 48 11847
rect 54 11837 58 11892
rect 53 11823 58 11837
rect 43 11813 48 11823
rect 53 11799 58 11813
rect 54 11798 58 11799
rect 78 11798 82 11892
rect 102 11798 106 11892
rect 126 11798 130 11892
rect 150 11798 154 11892
rect 174 11798 178 11892
rect 198 11798 202 11892
rect 222 11798 226 11892
rect 246 11798 250 11892
rect 270 11798 274 11892
rect 294 11798 298 11892
rect 318 11798 322 11892
rect 342 11798 346 11892
rect 366 11798 370 11892
rect 390 11798 394 11892
rect 414 11798 418 11892
rect 438 11798 442 11892
rect 462 11798 466 11892
rect 469 11891 483 11892
rect 486 11891 493 11915
rect 486 11798 490 11891
rect 510 11798 514 11964
rect 534 11798 538 11964
rect 558 11798 562 11964
rect 582 11798 586 11964
rect 606 11798 610 11964
rect 630 11798 634 11964
rect 654 11798 658 11964
rect 678 11798 682 11964
rect 702 11798 706 11964
rect 726 11798 730 11964
rect 750 11798 754 11964
rect 774 11798 778 11964
rect 798 11798 802 11964
rect 822 11798 826 11964
rect 846 11798 850 11964
rect 870 11798 874 11964
rect 894 11798 898 11964
rect 918 11798 922 11964
rect 942 11798 946 11964
rect 966 11798 970 11964
rect 990 11798 994 11964
rect 1014 11798 1018 11964
rect 1038 11798 1042 11964
rect 1062 11798 1066 11964
rect 1086 11798 1090 11964
rect 1110 11798 1114 11964
rect 1134 11798 1138 11964
rect 1158 11798 1162 11964
rect 1182 11798 1186 11964
rect 1206 11798 1210 11964
rect 1230 11798 1234 11964
rect 1254 11798 1258 11964
rect 1278 11798 1282 11964
rect 1302 11798 1306 11964
rect 1326 11798 1330 11964
rect 1350 11798 1354 11964
rect 1374 11798 1378 11964
rect 1398 11798 1402 11964
rect 1422 11798 1426 11964
rect 1435 11957 1440 11964
rect 1446 11957 1450 11964
rect 1445 11943 1450 11957
rect 1435 11933 1440 11943
rect 1445 11919 1450 11933
rect 1446 11798 1450 11919
rect 1470 11891 1474 12012
rect 1470 11843 1477 11891
rect 1470 11798 1474 11843
rect 1494 11798 1498 12012
rect 1518 11798 1522 12012
rect 1542 11798 1546 12012
rect 1566 11798 1570 12012
rect 1590 11798 1594 12012
rect 1614 11987 1618 12012
rect 1614 11942 1621 11987
rect 1638 11942 1642 12012
rect 1662 11942 1666 12012
rect 1686 11942 1690 12012
rect 1710 11942 1714 12012
rect 1734 11942 1738 12012
rect 1758 11942 1762 12012
rect 1782 11942 1786 12012
rect 1806 11942 1810 12012
rect 1830 11942 1834 12012
rect 1854 11942 1858 12012
rect 1861 12011 1875 12012
rect 1878 12011 1885 12035
rect 1878 11963 1885 11987
rect 1878 11942 1882 11963
rect 1902 11942 1906 12060
rect 1926 11942 1930 12060
rect 1950 11942 1954 12060
rect 1974 11942 1978 12060
rect 1998 11942 2002 12060
rect 2022 11942 2026 12060
rect 2046 11942 2050 12060
rect 2070 11942 2074 12060
rect 2094 11942 2098 12060
rect 2118 11942 2122 12060
rect 2142 11942 2146 12060
rect 2166 11942 2170 12060
rect 2190 11942 2194 12060
rect 2214 11942 2218 12060
rect 2238 11942 2242 12060
rect 2262 11942 2266 12060
rect 2286 11942 2290 12060
rect 2310 11942 2314 12060
rect 2334 11942 2338 12060
rect 2358 11942 2362 12060
rect 2382 11942 2386 12060
rect 2406 11942 2410 12060
rect 2430 11942 2434 12060
rect 2454 11942 2458 12060
rect 2478 11942 2482 12060
rect 2491 12005 2496 12015
rect 2526 12011 2530 12060
rect 2501 11991 2506 12005
rect 2515 12001 2523 12005
rect 2509 11991 2515 12001
rect 2502 11942 2506 11991
rect 2526 11987 2533 12011
rect 2550 11942 2554 12060
rect 2574 11942 2578 12060
rect 2598 11942 2602 12060
rect 2622 11942 2626 12060
rect 2646 11942 2650 12060
rect 2670 11942 2674 12060
rect 2694 11942 2698 12060
rect 2718 11942 2722 12060
rect 2742 11942 2746 12060
rect 2766 11942 2770 12060
rect 2790 11942 2794 12060
rect 2814 11942 2818 12060
rect 2838 11942 2842 12060
rect 2862 11942 2866 12060
rect 2886 11942 2890 12060
rect 2910 11942 2914 12060
rect 2934 11942 2938 12060
rect 2958 11942 2962 12060
rect 2982 11942 2986 12060
rect 3006 11942 3010 12060
rect 3030 11942 3034 12060
rect 3054 11942 3058 12060
rect 3078 11942 3082 12060
rect 3102 11942 3106 12060
rect 3126 11942 3130 12060
rect 3150 11942 3154 12060
rect 3174 11942 3178 12060
rect 3198 11942 3202 12060
rect 3222 11943 3226 12060
rect 3235 12029 3240 12039
rect 3246 12029 3250 12060
rect 3259 12053 3264 12060
rect 3270 12053 3274 12060
rect 3277 12059 3291 12060
rect 3269 12039 3274 12053
rect 3245 12015 3250 12029
rect 3211 11942 3245 11943
rect 1597 11940 3245 11942
rect 1597 11939 1611 11940
rect 1614 11939 1621 11940
rect 1614 11798 1618 11939
rect 1638 11798 1642 11940
rect 1662 11798 1666 11940
rect 1686 11798 1690 11940
rect 1710 11798 1714 11940
rect 1734 11798 1738 11940
rect 1758 11798 1762 11940
rect 1782 11798 1786 11940
rect 1806 11798 1810 11940
rect 1830 11798 1834 11940
rect 1854 11798 1858 11940
rect 1878 11798 1882 11940
rect 1902 11798 1906 11940
rect 1926 11798 1930 11940
rect 1950 11798 1954 11940
rect 1974 11798 1978 11940
rect 1998 11798 2002 11940
rect 2022 11798 2026 11940
rect 2046 11798 2050 11940
rect 2070 11798 2074 11940
rect 2094 11798 2098 11940
rect 2118 11798 2122 11940
rect 2142 11798 2146 11940
rect 2166 11798 2170 11940
rect 2190 11798 2194 11940
rect 2214 11798 2218 11940
rect 2238 11798 2242 11940
rect 2262 11798 2266 11940
rect 2286 11798 2290 11940
rect 2310 11798 2314 11940
rect 2334 11798 2338 11940
rect 2358 11798 2362 11940
rect 2382 11798 2386 11940
rect 2406 11798 2410 11940
rect 2430 11798 2434 11940
rect 2454 11798 2458 11940
rect 2478 11798 2482 11940
rect 2502 11798 2506 11940
rect 2526 11915 2533 11939
rect 2526 11798 2530 11915
rect 2550 11798 2554 11940
rect 2574 11798 2578 11940
rect 2598 11798 2602 11940
rect 2622 11798 2626 11940
rect 2646 11798 2650 11940
rect 2670 11798 2674 11940
rect 2694 11798 2698 11940
rect 2718 11798 2722 11940
rect 2742 11798 2746 11940
rect 2766 11798 2770 11940
rect 2790 11798 2794 11940
rect 2814 11798 2818 11940
rect 2838 11798 2842 11940
rect 2862 11798 2866 11940
rect 2886 11798 2890 11940
rect 2910 11798 2914 11940
rect 2934 11798 2938 11940
rect 2958 11798 2962 11940
rect 2982 11798 2986 11940
rect 3006 11798 3010 11940
rect 3030 11798 3034 11940
rect 3054 11798 3058 11940
rect 3078 11798 3082 11940
rect 3102 11798 3106 11940
rect 3126 11798 3130 11940
rect 3150 11798 3154 11940
rect 3174 11798 3178 11940
rect 3198 11798 3202 11940
rect 3211 11933 3216 11940
rect 3222 11933 3226 11940
rect 3221 11919 3226 11933
rect 3211 11885 3216 11895
rect 3221 11871 3226 11885
rect 3211 11813 3216 11823
rect 3222 11813 3226 11871
rect 3221 11799 3226 11813
rect 3235 11809 3243 11813
rect 3229 11799 3235 11809
rect 3211 11798 3243 11799
rect -2393 11796 3243 11798
rect -2371 11750 -2366 11796
rect -2348 11750 -2343 11796
rect -2325 11792 -2317 11796
rect -2325 11774 -2320 11792
rect -2317 11786 -2309 11792
rect -2095 11790 -2083 11796
rect -2053 11794 -1972 11796
rect -2083 11788 -2079 11790
rect -2079 11787 -2067 11788
rect -2079 11786 -2043 11787
rect -2091 11782 -2043 11786
rect -2000 11782 -1992 11794
rect -1671 11792 -1663 11796
rect -1982 11782 -1916 11787
rect -1663 11786 -1655 11792
rect -2091 11781 -2018 11782
rect -2091 11779 -2067 11781
rect -2053 11779 -2018 11781
rect -2002 11781 -1916 11782
rect -2002 11779 -1972 11781
rect -1924 11779 -1916 11781
rect -2079 11777 -2067 11779
rect -2000 11778 -1992 11779
rect -2325 11764 -2317 11774
rect -2112 11773 -2096 11777
rect -2083 11774 -2079 11777
rect -2027 11776 -1992 11778
rect -2109 11772 -2096 11773
rect -2112 11765 -2096 11772
rect -2083 11765 -2053 11772
rect -2018 11768 -2017 11776
rect -2023 11766 -2017 11768
rect -2009 11768 -2002 11771
rect -2009 11766 -2003 11768
rect -2109 11764 -2096 11765
rect -2325 11750 -2320 11764
rect -2317 11758 -2309 11764
rect -2112 11761 -2096 11764
rect -2017 11755 -2003 11766
rect -2017 11754 -2009 11755
rect -2074 11750 -2040 11752
rect -2000 11750 -1992 11776
rect -1972 11765 -1924 11772
rect -1671 11764 -1663 11774
rect -1663 11758 -1655 11764
rect -1642 11750 -1637 11796
rect -1619 11750 -1614 11796
rect -1530 11750 -1526 11796
rect -1506 11750 -1502 11796
rect -1482 11750 -1478 11796
rect -1458 11750 -1454 11796
rect -1434 11750 -1430 11796
rect -1410 11750 -1406 11796
rect -1386 11750 -1382 11796
rect -1362 11750 -1358 11796
rect -1338 11750 -1334 11796
rect -1314 11750 -1310 11796
rect -1290 11750 -1286 11796
rect -1266 11750 -1262 11796
rect -1242 11750 -1238 11796
rect -1218 11750 -1214 11796
rect -1194 11750 -1190 11796
rect -1170 11750 -1166 11796
rect -1146 11750 -1142 11796
rect -1122 11750 -1118 11796
rect -1098 11750 -1094 11796
rect -1074 11750 -1070 11796
rect -1050 11750 -1046 11796
rect -1026 11750 -1022 11796
rect -1002 11750 -998 11796
rect -978 11750 -974 11796
rect -954 11750 -950 11796
rect -930 11750 -926 11796
rect -906 11750 -902 11796
rect -882 11750 -878 11796
rect -858 11750 -854 11796
rect -834 11750 -830 11796
rect -810 11750 -806 11796
rect -786 11750 -782 11796
rect -762 11750 -758 11796
rect -738 11750 -734 11796
rect -714 11750 -710 11796
rect -690 11750 -686 11796
rect -666 11750 -662 11796
rect -642 11750 -638 11796
rect -618 11750 -614 11796
rect -594 11750 -590 11796
rect -570 11750 -566 11796
rect -546 11750 -542 11796
rect -522 11750 -518 11796
rect -498 11750 -494 11796
rect -474 11750 -470 11796
rect -450 11750 -446 11796
rect -426 11750 -422 11796
rect -402 11750 -398 11796
rect -378 11750 -374 11796
rect -354 11750 -350 11796
rect -330 11750 -326 11796
rect -306 11750 -302 11796
rect -282 11750 -278 11796
rect -258 11750 -254 11796
rect -234 11750 -230 11796
rect -210 11750 -206 11796
rect -186 11750 -182 11796
rect -162 11750 -158 11796
rect -138 11750 -134 11796
rect -114 11750 -110 11796
rect -101 11765 -96 11775
rect -90 11765 -86 11796
rect -91 11751 -86 11765
rect -90 11750 -86 11751
rect -66 11750 -62 11796
rect -42 11750 -38 11796
rect -18 11750 -14 11796
rect 6 11750 10 11796
rect 30 11750 34 11796
rect 54 11750 58 11796
rect 78 11771 82 11796
rect -2393 11748 75 11750
rect -2371 11702 -2366 11748
rect -2348 11702 -2343 11748
rect -2325 11746 -2320 11748
rect -2325 11736 -2317 11746
rect -2325 11716 -2320 11736
rect -2317 11730 -2309 11736
rect -2325 11708 -2317 11716
rect -2101 11711 -2071 11714
rect -2325 11702 -2320 11708
rect -2317 11702 -2309 11708
rect -2000 11706 -1992 11748
rect -1671 11736 -1663 11746
rect -1663 11730 -1655 11736
rect -1854 11720 -1680 11724
rect -1846 11711 -1798 11714
rect -2079 11705 -2043 11706
rect -2007 11705 -1991 11706
rect -2079 11704 -2071 11705
rect -2079 11702 -2029 11704
rect -2011 11702 -1991 11705
rect -1846 11703 -1806 11709
rect -1671 11708 -1663 11716
rect -1864 11702 -1796 11703
rect -1663 11702 -1655 11708
rect -1642 11702 -1637 11748
rect -1619 11702 -1614 11748
rect -1530 11702 -1526 11748
rect -1506 11702 -1502 11748
rect -1482 11702 -1478 11748
rect -1458 11702 -1454 11748
rect -1434 11702 -1430 11748
rect -1410 11702 -1406 11748
rect -1386 11702 -1382 11748
rect -1362 11702 -1358 11748
rect -1338 11702 -1334 11748
rect -1314 11702 -1310 11748
rect -1290 11702 -1286 11748
rect -1266 11702 -1262 11748
rect -1242 11702 -1238 11748
rect -1218 11702 -1214 11748
rect -1194 11702 -1190 11748
rect -1170 11702 -1166 11748
rect -1146 11702 -1142 11748
rect -1122 11702 -1118 11748
rect -1098 11702 -1094 11748
rect -1074 11702 -1070 11748
rect -1050 11702 -1046 11748
rect -1026 11702 -1022 11748
rect -1002 11702 -998 11748
rect -978 11702 -974 11748
rect -954 11702 -950 11748
rect -930 11702 -926 11748
rect -906 11702 -902 11748
rect -882 11702 -878 11748
rect -858 11702 -854 11748
rect -834 11702 -830 11748
rect -810 11702 -806 11748
rect -786 11702 -782 11748
rect -762 11702 -758 11748
rect -749 11717 -744 11727
rect -738 11717 -734 11748
rect -739 11703 -734 11717
rect -714 11702 -710 11748
rect -690 11702 -686 11748
rect -666 11702 -662 11748
rect -642 11702 -638 11748
rect -618 11702 -614 11748
rect -594 11702 -590 11748
rect -570 11702 -566 11748
rect -546 11702 -542 11748
rect -522 11702 -518 11748
rect -498 11702 -494 11748
rect -474 11702 -470 11748
rect -450 11702 -446 11748
rect -426 11702 -422 11748
rect -402 11702 -398 11748
rect -378 11702 -374 11748
rect -354 11702 -350 11748
rect -330 11702 -326 11748
rect -306 11702 -302 11748
rect -282 11702 -278 11748
rect -258 11702 -254 11748
rect -234 11702 -230 11748
rect -210 11702 -206 11748
rect -186 11702 -182 11748
rect -162 11702 -158 11748
rect -138 11702 -134 11748
rect -114 11702 -110 11748
rect -90 11702 -86 11748
rect -66 11702 -62 11748
rect -42 11702 -38 11748
rect -18 11702 -14 11748
rect 6 11702 10 11748
rect 30 11702 34 11748
rect 54 11702 58 11748
rect 61 11747 75 11748
rect 78 11723 85 11771
rect 78 11702 82 11723
rect 102 11702 106 11796
rect 126 11702 130 11796
rect 150 11702 154 11796
rect 174 11702 178 11796
rect 198 11702 202 11796
rect 222 11702 226 11796
rect 246 11702 250 11796
rect 270 11702 274 11796
rect 294 11703 298 11796
rect 283 11702 317 11703
rect -2393 11700 317 11702
rect -2371 11654 -2366 11700
rect -2348 11654 -2343 11700
rect -2325 11688 -2320 11700
rect -2079 11698 -2071 11700
rect -2072 11696 -2071 11698
rect -2109 11691 -2101 11696
rect -2101 11689 -2079 11691
rect -2069 11689 -2068 11696
rect -2325 11680 -2317 11688
rect -2079 11684 -2071 11689
rect -2325 11660 -2320 11680
rect -2317 11672 -2309 11680
rect -2074 11675 -2071 11684
rect -2069 11680 -2068 11684
rect -2109 11666 -2079 11669
rect -2325 11654 -2317 11660
rect -2000 11654 -1992 11700
rect -1846 11698 -1806 11700
rect -1854 11693 -1806 11697
rect -1854 11691 -1846 11693
rect -1846 11689 -1806 11691
rect -1806 11687 -1798 11689
rect -1846 11684 -1798 11687
rect -1846 11671 -1806 11682
rect -1671 11680 -1663 11688
rect -1663 11672 -1655 11680
rect -1854 11666 -1680 11670
rect -1671 11654 -1663 11660
rect -1642 11654 -1637 11700
rect -1619 11654 -1614 11700
rect -1530 11654 -1526 11700
rect -1506 11654 -1502 11700
rect -1482 11654 -1478 11700
rect -1458 11654 -1454 11700
rect -1434 11654 -1430 11700
rect -1410 11654 -1406 11700
rect -1386 11654 -1382 11700
rect -1362 11654 -1358 11700
rect -1338 11654 -1334 11700
rect -1314 11654 -1310 11700
rect -1290 11654 -1286 11700
rect -1266 11654 -1262 11700
rect -1242 11654 -1238 11700
rect -1218 11654 -1214 11700
rect -1194 11654 -1190 11700
rect -1170 11654 -1166 11700
rect -1146 11654 -1142 11700
rect -1122 11654 -1118 11700
rect -1098 11654 -1094 11700
rect -1074 11654 -1070 11700
rect -1050 11654 -1046 11700
rect -1026 11654 -1022 11700
rect -1002 11654 -998 11700
rect -978 11654 -974 11700
rect -954 11654 -950 11700
rect -930 11654 -926 11700
rect -906 11654 -902 11700
rect -882 11654 -878 11700
rect -858 11654 -854 11700
rect -834 11654 -830 11700
rect -810 11654 -806 11700
rect -786 11654 -782 11700
rect -762 11654 -758 11700
rect -749 11678 -715 11679
rect -714 11678 -710 11700
rect -690 11678 -686 11700
rect -666 11678 -662 11700
rect -642 11678 -638 11700
rect -618 11678 -614 11700
rect -594 11678 -590 11700
rect -570 11678 -566 11700
rect -546 11678 -542 11700
rect -522 11678 -518 11700
rect -498 11678 -494 11700
rect -474 11678 -470 11700
rect -450 11678 -446 11700
rect -426 11678 -422 11700
rect -402 11678 -398 11700
rect -378 11678 -374 11700
rect -354 11678 -350 11700
rect -330 11678 -326 11700
rect -306 11678 -302 11700
rect -282 11678 -278 11700
rect -258 11678 -254 11700
rect -234 11678 -230 11700
rect -210 11678 -206 11700
rect -186 11678 -182 11700
rect -162 11678 -158 11700
rect -138 11678 -134 11700
rect -114 11678 -110 11700
rect -90 11678 -86 11700
rect -66 11699 -62 11700
rect -749 11676 -69 11678
rect -749 11669 -744 11676
rect -739 11655 -734 11669
rect -738 11654 -734 11655
rect -714 11654 -710 11676
rect -690 11654 -686 11676
rect -666 11654 -662 11676
rect -642 11654 -638 11676
rect -618 11654 -614 11676
rect -594 11654 -590 11676
rect -570 11654 -566 11676
rect -546 11654 -542 11676
rect -522 11654 -518 11676
rect -498 11654 -494 11676
rect -474 11654 -470 11676
rect -450 11654 -446 11676
rect -426 11654 -422 11676
rect -402 11654 -398 11676
rect -378 11654 -374 11676
rect -354 11654 -350 11676
rect -330 11654 -326 11676
rect -306 11654 -302 11676
rect -282 11654 -278 11676
rect -258 11654 -254 11676
rect -234 11654 -230 11676
rect -210 11654 -206 11676
rect -186 11654 -182 11676
rect -162 11654 -158 11676
rect -138 11654 -134 11676
rect -114 11654 -110 11676
rect -90 11654 -86 11676
rect -83 11675 -69 11676
rect -66 11675 -59 11699
rect -66 11654 -62 11675
rect -42 11654 -38 11700
rect -18 11654 -14 11700
rect 6 11654 10 11700
rect 30 11654 34 11700
rect 54 11654 58 11700
rect 78 11654 82 11700
rect 102 11654 106 11700
rect 126 11654 130 11700
rect 150 11654 154 11700
rect 174 11654 178 11700
rect 198 11654 202 11700
rect 222 11654 226 11700
rect 246 11654 250 11700
rect 270 11654 274 11700
rect 283 11693 288 11700
rect 294 11693 298 11700
rect 293 11679 298 11693
rect 283 11654 317 11655
rect -2393 11652 317 11654
rect -2371 11630 -2366 11652
rect -2348 11630 -2343 11652
rect -2325 11644 -2317 11652
rect -2325 11630 -2320 11644
rect -2309 11632 -2301 11644
rect -2092 11635 -2062 11640
rect -2000 11632 -1992 11652
rect -2317 11630 -2309 11632
rect -2000 11630 -1983 11632
rect -1906 11630 -1904 11652
rect -1806 11644 -1680 11650
rect -1671 11644 -1663 11652
rect -1854 11635 -1806 11640
rect -1846 11630 -1806 11633
rect -1655 11632 -1647 11644
rect -1663 11630 -1655 11632
rect -1642 11630 -1637 11652
rect -1619 11630 -1614 11652
rect -1530 11630 -1526 11652
rect -1506 11630 -1502 11652
rect -1482 11630 -1478 11652
rect -1458 11630 -1454 11652
rect -1434 11630 -1430 11652
rect -1410 11630 -1406 11652
rect -1386 11630 -1382 11652
rect -1362 11630 -1358 11652
rect -1338 11630 -1334 11652
rect -1314 11630 -1310 11652
rect -1290 11630 -1286 11652
rect -1266 11630 -1262 11652
rect -1242 11630 -1238 11652
rect -1218 11630 -1214 11652
rect -1194 11630 -1190 11652
rect -1170 11630 -1166 11652
rect -1146 11630 -1142 11652
rect -1122 11630 -1118 11652
rect -1098 11630 -1094 11652
rect -1074 11630 -1070 11652
rect -1050 11630 -1046 11652
rect -1026 11630 -1022 11652
rect -1002 11630 -998 11652
rect -978 11630 -974 11652
rect -954 11630 -950 11652
rect -930 11630 -926 11652
rect -906 11630 -902 11652
rect -882 11630 -878 11652
rect -858 11630 -854 11652
rect -834 11630 -830 11652
rect -810 11630 -806 11652
rect -786 11630 -782 11652
rect -762 11630 -758 11652
rect -738 11630 -734 11652
rect -714 11651 -710 11652
rect -2393 11628 -717 11630
rect -2371 11606 -2366 11628
rect -2348 11606 -2343 11628
rect -2325 11616 -2317 11628
rect -2071 11624 -2062 11628
rect -2013 11626 -1983 11628
rect -2000 11625 -1983 11626
rect -2325 11606 -2320 11616
rect -2309 11606 -2301 11616
rect -2100 11615 -2092 11622
rect -2064 11620 -2062 11623
rect -2061 11615 -2059 11620
rect -2071 11610 -2062 11615
rect -2071 11608 -2026 11610
rect -2066 11606 -2012 11608
rect -2000 11606 -1992 11625
rect -1906 11623 -1904 11628
rect -1846 11624 -1806 11628
rect -1846 11617 -1798 11622
rect -1806 11615 -1798 11617
rect -1671 11616 -1663 11628
rect -1854 11613 -1846 11615
rect -1854 11608 -1806 11613
rect -1864 11606 -1796 11607
rect -1655 11606 -1647 11616
rect -1642 11606 -1637 11628
rect -1619 11606 -1614 11628
rect -1530 11606 -1526 11628
rect -1506 11606 -1502 11628
rect -1482 11606 -1478 11628
rect -1458 11606 -1454 11628
rect -1434 11606 -1430 11628
rect -1410 11606 -1406 11628
rect -1386 11606 -1382 11628
rect -1362 11606 -1358 11628
rect -1338 11606 -1334 11628
rect -1314 11606 -1310 11628
rect -1290 11606 -1286 11628
rect -1266 11606 -1262 11628
rect -1242 11606 -1238 11628
rect -1218 11606 -1214 11628
rect -1194 11606 -1190 11628
rect -1170 11606 -1166 11628
rect -1146 11606 -1142 11628
rect -1122 11606 -1118 11628
rect -1098 11606 -1094 11628
rect -1074 11606 -1070 11628
rect -1050 11606 -1046 11628
rect -1026 11606 -1022 11628
rect -1002 11606 -998 11628
rect -978 11606 -974 11628
rect -954 11606 -950 11628
rect -930 11606 -926 11628
rect -906 11606 -902 11628
rect -882 11606 -878 11628
rect -858 11606 -854 11628
rect -834 11606 -830 11628
rect -810 11606 -806 11628
rect -786 11606 -782 11628
rect -762 11606 -758 11628
rect -738 11606 -734 11628
rect -731 11627 -717 11628
rect -714 11627 -707 11651
rect -690 11606 -686 11652
rect -666 11606 -662 11652
rect -642 11606 -638 11652
rect -618 11606 -614 11652
rect -594 11606 -590 11652
rect -570 11606 -566 11652
rect -546 11606 -542 11652
rect -522 11606 -518 11652
rect -498 11606 -494 11652
rect -474 11606 -470 11652
rect -450 11607 -446 11652
rect -461 11606 -427 11607
rect -2393 11604 -427 11606
rect -2371 11558 -2366 11604
rect -2348 11558 -2343 11604
rect -2325 11600 -2320 11604
rect -2317 11600 -2309 11604
rect -2325 11588 -2317 11600
rect -2066 11599 -2062 11604
rect -2147 11596 -2134 11598
rect -2292 11590 -2071 11596
rect -2325 11568 -2320 11588
rect -2092 11574 -2062 11576
rect -2094 11570 -2062 11574
rect -2325 11558 -2317 11568
rect -2095 11560 -2084 11564
rect -2000 11561 -1992 11604
rect -1846 11597 -1806 11604
rect -1663 11600 -1655 11604
rect -1846 11590 -1680 11596
rect -1671 11588 -1663 11600
rect -1854 11574 -1806 11576
rect -1854 11570 -1680 11574
rect -2119 11558 -2069 11560
rect -2054 11558 -1892 11561
rect -1671 11558 -1663 11568
rect -1642 11558 -1637 11604
rect -1619 11558 -1614 11604
rect -1530 11558 -1526 11604
rect -1506 11558 -1502 11604
rect -1482 11558 -1478 11604
rect -1458 11558 -1454 11604
rect -1434 11558 -1430 11604
rect -1410 11558 -1406 11604
rect -1386 11558 -1382 11604
rect -1362 11558 -1358 11604
rect -1338 11558 -1334 11604
rect -1314 11558 -1310 11604
rect -1290 11558 -1286 11604
rect -1266 11558 -1262 11604
rect -1242 11558 -1238 11604
rect -1218 11558 -1214 11604
rect -1194 11558 -1190 11604
rect -1170 11558 -1166 11604
rect -1146 11558 -1142 11604
rect -1122 11558 -1118 11604
rect -1098 11558 -1094 11604
rect -1074 11558 -1070 11604
rect -1050 11558 -1046 11604
rect -1026 11558 -1022 11604
rect -1002 11558 -998 11604
rect -978 11558 -974 11604
rect -954 11558 -950 11604
rect -930 11558 -926 11604
rect -906 11558 -902 11604
rect -882 11558 -878 11604
rect -858 11558 -854 11604
rect -834 11558 -830 11604
rect -810 11558 -806 11604
rect -786 11558 -782 11604
rect -762 11558 -758 11604
rect -738 11558 -734 11604
rect -714 11579 -707 11603
rect -714 11558 -710 11579
rect -690 11558 -686 11604
rect -666 11558 -662 11604
rect -642 11558 -638 11604
rect -618 11558 -614 11604
rect -594 11558 -590 11604
rect -570 11558 -566 11604
rect -546 11558 -542 11604
rect -522 11558 -518 11604
rect -498 11558 -494 11604
rect -474 11558 -470 11604
rect -461 11597 -456 11604
rect -450 11597 -446 11604
rect -451 11583 -446 11597
rect -461 11582 -427 11583
rect -426 11582 -422 11652
rect -402 11582 -398 11652
rect -378 11582 -374 11652
rect -354 11582 -350 11652
rect -330 11582 -326 11652
rect -306 11582 -302 11652
rect -282 11582 -278 11652
rect -258 11582 -254 11652
rect -234 11582 -230 11652
rect -210 11582 -206 11652
rect -186 11582 -182 11652
rect -162 11582 -158 11652
rect -138 11582 -134 11652
rect -114 11582 -110 11652
rect -90 11582 -86 11652
rect -66 11582 -62 11652
rect -42 11582 -38 11652
rect -18 11582 -14 11652
rect 6 11582 10 11652
rect 30 11582 34 11652
rect 54 11582 58 11652
rect 78 11582 82 11652
rect 102 11582 106 11652
rect 126 11582 130 11652
rect 150 11582 154 11652
rect 174 11582 178 11652
rect 198 11582 202 11652
rect 222 11582 226 11652
rect 246 11582 250 11652
rect 270 11582 274 11652
rect 283 11645 288 11652
rect 293 11631 298 11645
rect 294 11582 298 11631
rect 318 11627 322 11796
rect 318 11603 325 11627
rect 342 11582 346 11796
rect 366 11582 370 11796
rect 390 11582 394 11796
rect 414 11582 418 11796
rect 438 11582 442 11796
rect 462 11582 466 11796
rect 486 11582 490 11796
rect 510 11582 514 11796
rect 534 11582 538 11796
rect 558 11582 562 11796
rect 582 11582 586 11796
rect 606 11582 610 11796
rect 630 11582 634 11796
rect 654 11582 658 11796
rect 678 11582 682 11796
rect 702 11582 706 11796
rect 726 11582 730 11796
rect 750 11582 754 11796
rect 774 11582 778 11796
rect 798 11582 802 11796
rect 822 11582 826 11796
rect 846 11582 850 11796
rect 870 11582 874 11796
rect 894 11582 898 11796
rect 918 11582 922 11796
rect 942 11582 946 11796
rect 955 11741 960 11751
rect 966 11741 970 11796
rect 965 11727 970 11741
rect 966 11582 970 11727
rect 990 11675 994 11796
rect 990 11651 997 11675
rect 990 11582 994 11651
rect 1014 11582 1018 11796
rect 1038 11582 1042 11796
rect 1062 11582 1066 11796
rect 1086 11582 1090 11796
rect 1110 11582 1114 11796
rect 1134 11582 1138 11796
rect 1158 11582 1162 11796
rect 1182 11582 1186 11796
rect 1206 11582 1210 11796
rect 1230 11582 1234 11796
rect 1254 11582 1258 11796
rect 1278 11582 1282 11796
rect 1302 11582 1306 11796
rect 1326 11582 1330 11796
rect 1350 11582 1354 11796
rect 1374 11582 1378 11796
rect 1398 11582 1402 11796
rect 1422 11582 1426 11796
rect 1446 11582 1450 11796
rect 1470 11582 1474 11796
rect 1494 11582 1498 11796
rect 1518 11582 1522 11796
rect 1542 11582 1546 11796
rect 1566 11582 1570 11796
rect 1590 11582 1594 11796
rect 1614 11582 1618 11796
rect 1627 11621 1632 11631
rect 1638 11621 1642 11796
rect 1637 11607 1642 11621
rect 1627 11597 1632 11607
rect 1637 11583 1642 11597
rect 1638 11582 1642 11583
rect 1662 11582 1666 11796
rect 1686 11582 1690 11796
rect 1710 11582 1714 11796
rect 1734 11582 1738 11796
rect 1758 11582 1762 11796
rect 1782 11582 1786 11796
rect 1806 11582 1810 11796
rect 1830 11582 1834 11796
rect 1854 11582 1858 11796
rect 1878 11582 1882 11796
rect 1902 11582 1906 11796
rect 1926 11582 1930 11796
rect 1950 11582 1954 11796
rect 1974 11582 1978 11796
rect 1998 11582 2002 11796
rect 2022 11582 2026 11796
rect 2046 11582 2050 11796
rect 2070 11582 2074 11796
rect 2094 11582 2098 11796
rect 2118 11582 2122 11796
rect 2142 11582 2146 11796
rect 2166 11582 2170 11796
rect 2190 11582 2194 11796
rect 2214 11582 2218 11796
rect 2238 11582 2242 11796
rect 2262 11582 2266 11796
rect 2286 11582 2290 11796
rect 2310 11582 2314 11796
rect 2334 11582 2338 11796
rect 2358 11582 2362 11796
rect 2382 11582 2386 11796
rect 2406 11582 2410 11796
rect 2430 11582 2434 11796
rect 2454 11582 2458 11796
rect 2478 11582 2482 11796
rect 2502 11582 2506 11796
rect 2526 11582 2530 11796
rect 2550 11582 2554 11796
rect 2574 11582 2578 11796
rect 2598 11582 2602 11796
rect 2622 11582 2626 11796
rect 2646 11582 2650 11796
rect 2670 11582 2674 11796
rect 2694 11582 2698 11796
rect 2718 11582 2722 11796
rect 2742 11582 2746 11796
rect 2766 11582 2770 11796
rect 2790 11582 2794 11796
rect 2814 11582 2818 11796
rect 2838 11582 2842 11796
rect 2862 11582 2866 11796
rect 2886 11582 2890 11796
rect 2910 11582 2914 11796
rect 2934 11582 2938 11796
rect 2958 11582 2962 11796
rect 2982 11582 2986 11796
rect 3006 11582 3010 11796
rect 3030 11582 3034 11796
rect 3054 11582 3058 11796
rect 3078 11582 3082 11796
rect 3102 11582 3106 11796
rect 3126 11582 3130 11796
rect 3150 11582 3154 11796
rect 3174 11583 3178 11796
rect 3187 11597 3192 11607
rect 3198 11597 3202 11796
rect 3211 11789 3216 11796
rect 3229 11795 3243 11796
rect 3221 11775 3226 11789
rect 3211 11669 3216 11679
rect 3222 11669 3226 11775
rect 3221 11655 3226 11669
rect 3197 11583 3202 11597
rect 3163 11582 3197 11583
rect -461 11580 3197 11582
rect -461 11573 -456 11580
rect -451 11559 -446 11573
rect -450 11558 -446 11559
rect -426 11558 -422 11580
rect -402 11558 -398 11580
rect -378 11558 -374 11580
rect -354 11558 -350 11580
rect -330 11558 -326 11580
rect -306 11558 -302 11580
rect -282 11558 -278 11580
rect -258 11558 -254 11580
rect -234 11558 -230 11580
rect -210 11558 -206 11580
rect -186 11558 -182 11580
rect -162 11558 -158 11580
rect -138 11558 -134 11580
rect -114 11558 -110 11580
rect -90 11558 -86 11580
rect -66 11558 -62 11580
rect -42 11558 -38 11580
rect -18 11558 -14 11580
rect 6 11558 10 11580
rect 30 11558 34 11580
rect 54 11558 58 11580
rect 78 11558 82 11580
rect 102 11558 106 11580
rect 126 11558 130 11580
rect 150 11558 154 11580
rect 174 11558 178 11580
rect 198 11558 202 11580
rect 222 11558 226 11580
rect 246 11558 250 11580
rect 270 11558 274 11580
rect 294 11558 298 11580
rect -2393 11556 315 11558
rect -2371 11534 -2366 11556
rect -2348 11534 -2343 11556
rect -2325 11552 -2317 11556
rect -2325 11536 -2320 11552
rect -2309 11540 -2301 11552
rect -2095 11550 -2084 11556
rect -2054 11555 -1906 11556
rect -2054 11554 -2036 11555
rect -2084 11548 -2079 11550
rect -2317 11536 -2309 11540
rect -2092 11539 -2079 11546
rect -2000 11542 -1992 11555
rect -1920 11554 -1906 11555
rect -1671 11552 -1663 11556
rect -1846 11548 -1806 11550
rect -1854 11542 -1806 11546
rect -2054 11539 -1982 11542
rect -1966 11539 -1806 11542
rect -1655 11540 -1647 11552
rect -2003 11536 -1992 11539
rect -1904 11537 -1902 11539
rect -1854 11537 -1846 11539
rect -2325 11534 -2317 11536
rect -2033 11534 -1992 11536
rect -1854 11535 -1806 11537
rect -1663 11536 -1655 11540
rect -1864 11534 -1796 11535
rect -1671 11534 -1663 11536
rect -1642 11534 -1637 11556
rect -1619 11534 -1614 11556
rect -1530 11534 -1526 11556
rect -1506 11534 -1502 11556
rect -1482 11534 -1478 11556
rect -1458 11534 -1454 11556
rect -1434 11534 -1430 11556
rect -1410 11534 -1406 11556
rect -1386 11534 -1382 11556
rect -1362 11534 -1358 11556
rect -1338 11534 -1334 11556
rect -1314 11534 -1310 11556
rect -1290 11534 -1286 11556
rect -1266 11534 -1262 11556
rect -1242 11534 -1238 11556
rect -1218 11534 -1214 11556
rect -1194 11534 -1190 11556
rect -1170 11534 -1166 11556
rect -1146 11534 -1142 11556
rect -1122 11534 -1118 11556
rect -1098 11534 -1094 11556
rect -1074 11534 -1070 11556
rect -1050 11534 -1046 11556
rect -1026 11534 -1022 11556
rect -1002 11534 -998 11556
rect -978 11534 -974 11556
rect -954 11534 -950 11556
rect -930 11534 -926 11556
rect -906 11534 -902 11556
rect -882 11534 -878 11556
rect -858 11534 -854 11556
rect -834 11534 -830 11556
rect -810 11534 -806 11556
rect -786 11534 -782 11556
rect -762 11534 -758 11556
rect -738 11534 -734 11556
rect -714 11534 -710 11556
rect -690 11534 -686 11556
rect -666 11534 -662 11556
rect -642 11534 -638 11556
rect -618 11534 -614 11556
rect -594 11534 -590 11556
rect -570 11534 -566 11556
rect -546 11534 -542 11556
rect -522 11534 -518 11556
rect -498 11534 -494 11556
rect -474 11534 -470 11556
rect -450 11534 -446 11556
rect -426 11534 -422 11556
rect -402 11534 -398 11556
rect -378 11534 -374 11556
rect -354 11534 -350 11556
rect -330 11534 -326 11556
rect -306 11534 -302 11556
rect -282 11534 -278 11556
rect -258 11534 -254 11556
rect -234 11534 -230 11556
rect -210 11534 -206 11556
rect -186 11534 -182 11556
rect -162 11534 -158 11556
rect -138 11534 -134 11556
rect -114 11534 -110 11556
rect -90 11534 -86 11556
rect -66 11534 -62 11556
rect -42 11534 -38 11556
rect -18 11534 -14 11556
rect 6 11534 10 11556
rect 30 11534 34 11556
rect 54 11534 58 11556
rect 78 11534 82 11556
rect 102 11534 106 11556
rect 126 11534 130 11556
rect 150 11534 154 11556
rect 174 11534 178 11556
rect 198 11534 202 11556
rect 222 11534 226 11556
rect 246 11534 250 11556
rect 270 11534 274 11556
rect 294 11534 298 11556
rect 301 11555 315 11556
rect 318 11555 325 11579
rect 318 11534 322 11555
rect 342 11534 346 11580
rect 366 11534 370 11580
rect 390 11534 394 11580
rect 414 11534 418 11580
rect 438 11534 442 11580
rect 462 11534 466 11580
rect 486 11534 490 11580
rect 510 11534 514 11580
rect 534 11534 538 11580
rect 558 11534 562 11580
rect 582 11534 586 11580
rect 606 11534 610 11580
rect 630 11534 634 11580
rect 654 11534 658 11580
rect 678 11534 682 11580
rect 702 11534 706 11580
rect 726 11534 730 11580
rect 750 11534 754 11580
rect 774 11534 778 11580
rect 798 11534 802 11580
rect 822 11534 826 11580
rect 846 11535 850 11580
rect 835 11534 869 11535
rect -2393 11532 869 11534
rect -2371 11510 -2366 11532
rect -2348 11510 -2343 11532
rect -2325 11524 -2317 11532
rect -2079 11529 -2018 11532
rect -2003 11531 -1966 11532
rect -2000 11530 -1982 11531
rect -2000 11529 -1992 11530
rect -2084 11525 -2009 11529
rect -2028 11524 -2009 11525
rect -2000 11525 -1854 11529
rect -1846 11525 -1798 11532
rect -2325 11510 -2320 11524
rect -2309 11512 -2301 11524
rect -2028 11522 -2018 11524
rect -2092 11512 -2084 11519
rect -2023 11515 -2014 11522
rect -2000 11515 -1992 11525
rect -1671 11524 -1663 11532
rect -1846 11521 -1806 11523
rect -1854 11515 -1806 11519
rect -2054 11512 -1806 11515
rect -1655 11512 -1647 11524
rect -2317 11510 -2309 11512
rect -2054 11510 -2024 11512
rect -2000 11510 -1992 11512
rect -1663 11510 -1655 11512
rect -1642 11510 -1637 11532
rect -1619 11510 -1614 11532
rect -1530 11510 -1526 11532
rect -1506 11510 -1502 11532
rect -1482 11510 -1478 11532
rect -1458 11510 -1454 11532
rect -1434 11510 -1430 11532
rect -1410 11510 -1406 11532
rect -1386 11510 -1382 11532
rect -1362 11510 -1358 11532
rect -1338 11510 -1334 11532
rect -1314 11510 -1310 11532
rect -1290 11510 -1286 11532
rect -1266 11510 -1262 11532
rect -1242 11510 -1238 11532
rect -1218 11510 -1214 11532
rect -1194 11510 -1190 11532
rect -1170 11510 -1166 11532
rect -1146 11510 -1142 11532
rect -1122 11510 -1118 11532
rect -1098 11510 -1094 11532
rect -1074 11510 -1070 11532
rect -1050 11510 -1046 11532
rect -1026 11510 -1022 11532
rect -1002 11510 -998 11532
rect -978 11510 -974 11532
rect -954 11510 -950 11532
rect -930 11510 -926 11532
rect -906 11510 -902 11532
rect -882 11510 -878 11532
rect -858 11510 -854 11532
rect -834 11510 -830 11532
rect -810 11510 -806 11532
rect -786 11510 -782 11532
rect -762 11510 -758 11532
rect -738 11510 -734 11532
rect -714 11510 -710 11532
rect -690 11510 -686 11532
rect -666 11510 -662 11532
rect -642 11510 -638 11532
rect -618 11510 -614 11532
rect -594 11510 -590 11532
rect -570 11510 -566 11532
rect -546 11510 -542 11532
rect -522 11510 -518 11532
rect -498 11510 -494 11532
rect -474 11510 -470 11532
rect -450 11510 -446 11532
rect -426 11531 -422 11532
rect -2393 11508 -2064 11510
rect -2060 11508 -429 11510
rect -2371 11462 -2366 11508
rect -2348 11462 -2343 11508
rect -2325 11496 -2317 11508
rect -2060 11505 -2054 11508
rect -2084 11498 -2054 11505
rect -2050 11502 -2044 11504
rect -2325 11476 -2320 11496
rect -2064 11494 -2054 11498
rect -2325 11468 -2317 11476
rect -2101 11471 -2071 11474
rect -2325 11462 -2320 11468
rect -2317 11462 -2309 11468
rect -2000 11466 -1992 11508
rect -1846 11507 -1806 11508
rect -1846 11498 -1798 11505
rect -1671 11496 -1663 11508
rect -1846 11494 -1806 11496
rect -1854 11480 -1680 11484
rect -1846 11471 -1798 11474
rect -2079 11465 -2043 11466
rect -2007 11465 -1991 11466
rect -2079 11464 -2071 11465
rect -2079 11462 -2029 11464
rect -2011 11462 -1991 11465
rect -1846 11463 -1806 11469
rect -1671 11468 -1663 11476
rect -1864 11462 -1796 11463
rect -1663 11462 -1655 11468
rect -1642 11462 -1637 11508
rect -1619 11462 -1614 11508
rect -1530 11462 -1526 11508
rect -1506 11462 -1502 11508
rect -1482 11462 -1478 11508
rect -1458 11462 -1454 11508
rect -1434 11462 -1430 11508
rect -1410 11462 -1406 11508
rect -1386 11462 -1382 11508
rect -1362 11462 -1358 11508
rect -1338 11462 -1334 11508
rect -1314 11462 -1310 11508
rect -1290 11462 -1286 11508
rect -1266 11462 -1262 11508
rect -1242 11462 -1238 11508
rect -1218 11462 -1214 11508
rect -1194 11462 -1190 11508
rect -1170 11462 -1166 11508
rect -1146 11462 -1142 11508
rect -1122 11462 -1118 11508
rect -1098 11462 -1094 11508
rect -1074 11462 -1070 11508
rect -1050 11462 -1046 11508
rect -1026 11462 -1022 11508
rect -1002 11462 -998 11508
rect -978 11462 -974 11508
rect -954 11462 -950 11508
rect -930 11462 -926 11508
rect -906 11462 -902 11508
rect -882 11462 -878 11508
rect -858 11462 -854 11508
rect -834 11462 -830 11508
rect -810 11462 -806 11508
rect -786 11462 -782 11508
rect -762 11462 -758 11508
rect -738 11462 -734 11508
rect -714 11462 -710 11508
rect -690 11462 -686 11508
rect -666 11462 -662 11508
rect -642 11462 -638 11508
rect -618 11462 -614 11508
rect -594 11462 -590 11508
rect -570 11462 -566 11508
rect -546 11462 -542 11508
rect -522 11462 -518 11508
rect -498 11462 -494 11508
rect -474 11462 -470 11508
rect -450 11462 -446 11508
rect -443 11507 -429 11508
rect -426 11486 -419 11531
rect -402 11486 -398 11532
rect -378 11486 -374 11532
rect -354 11486 -350 11532
rect -330 11486 -326 11532
rect -306 11486 -302 11532
rect -282 11486 -278 11532
rect -258 11486 -254 11532
rect -234 11486 -230 11532
rect -210 11486 -206 11532
rect -186 11486 -182 11532
rect -162 11486 -158 11532
rect -138 11486 -134 11532
rect -114 11486 -110 11532
rect -90 11486 -86 11532
rect -66 11486 -62 11532
rect -42 11486 -38 11532
rect -18 11486 -14 11532
rect 6 11486 10 11532
rect 30 11486 34 11532
rect 54 11486 58 11532
rect 78 11486 82 11532
rect 102 11486 106 11532
rect 126 11486 130 11532
rect 150 11486 154 11532
rect 174 11486 178 11532
rect 198 11486 202 11532
rect 222 11486 226 11532
rect 246 11486 250 11532
rect 270 11486 274 11532
rect 294 11486 298 11532
rect 318 11486 322 11532
rect 342 11486 346 11532
rect 366 11486 370 11532
rect 390 11486 394 11532
rect 414 11486 418 11532
rect 438 11486 442 11532
rect 462 11486 466 11532
rect 486 11486 490 11532
rect 510 11486 514 11532
rect 534 11486 538 11532
rect 558 11486 562 11532
rect 582 11486 586 11532
rect 595 11501 600 11511
rect 606 11501 610 11532
rect 605 11487 610 11501
rect 630 11486 634 11532
rect 654 11486 658 11532
rect 678 11486 682 11532
rect 702 11486 706 11532
rect 726 11486 730 11532
rect 750 11486 754 11532
rect 774 11486 778 11532
rect 798 11486 802 11532
rect 822 11486 826 11532
rect 835 11525 840 11532
rect 846 11525 850 11532
rect 845 11511 850 11525
rect 835 11501 840 11511
rect 845 11487 850 11501
rect 846 11486 850 11487
rect 870 11486 874 11580
rect 894 11486 898 11580
rect 918 11486 922 11580
rect 942 11486 946 11580
rect 966 11486 970 11580
rect 990 11486 994 11580
rect 1014 11486 1018 11580
rect 1038 11486 1042 11580
rect 1062 11486 1066 11580
rect 1086 11486 1090 11580
rect 1110 11486 1114 11580
rect 1134 11486 1138 11580
rect 1158 11486 1162 11580
rect 1182 11486 1186 11580
rect 1206 11486 1210 11580
rect 1230 11486 1234 11580
rect 1254 11486 1258 11580
rect 1278 11486 1282 11580
rect 1302 11486 1306 11580
rect 1326 11486 1330 11580
rect 1350 11486 1354 11580
rect 1374 11486 1378 11580
rect 1398 11487 1402 11580
rect 1387 11486 1421 11487
rect -443 11484 1421 11486
rect -443 11483 -429 11484
rect -426 11483 -419 11484
rect -426 11462 -422 11483
rect -402 11462 -398 11484
rect -378 11462 -374 11484
rect -354 11462 -350 11484
rect -330 11462 -326 11484
rect -306 11462 -302 11484
rect -282 11462 -278 11484
rect -258 11462 -254 11484
rect -234 11462 -230 11484
rect -210 11462 -206 11484
rect -186 11462 -182 11484
rect -162 11462 -158 11484
rect -138 11462 -134 11484
rect -114 11462 -110 11484
rect -90 11462 -86 11484
rect -66 11462 -62 11484
rect -42 11462 -38 11484
rect -18 11462 -14 11484
rect 6 11462 10 11484
rect 30 11462 34 11484
rect 54 11462 58 11484
rect 78 11462 82 11484
rect 102 11462 106 11484
rect 126 11462 130 11484
rect 150 11463 154 11484
rect 139 11462 173 11463
rect -2393 11460 173 11462
rect -2371 11390 -2366 11460
rect -2348 11390 -2343 11460
rect -2325 11448 -2320 11460
rect -2079 11458 -2071 11460
rect -2072 11456 -2071 11458
rect -2109 11451 -2101 11456
rect -2101 11449 -2079 11451
rect -2069 11449 -2068 11456
rect -2325 11440 -2317 11448
rect -2079 11444 -2071 11449
rect -2325 11390 -2320 11440
rect -2317 11432 -2309 11440
rect -2074 11435 -2071 11444
rect -2069 11440 -2068 11444
rect -2109 11426 -2079 11429
rect -2309 11392 -2301 11402
rect -2317 11390 -2309 11392
rect -2000 11390 -1992 11460
rect -1846 11458 -1806 11460
rect -1854 11453 -1806 11457
rect -1854 11451 -1846 11453
rect -1846 11449 -1806 11451
rect -1806 11447 -1798 11449
rect -1846 11444 -1798 11447
rect -1846 11431 -1806 11442
rect -1671 11440 -1663 11448
rect -1663 11432 -1655 11440
rect -1854 11426 -1680 11430
rect -1655 11392 -1647 11402
rect -1663 11390 -1655 11392
rect -1642 11390 -1637 11460
rect -1619 11390 -1614 11460
rect -1530 11390 -1526 11460
rect -1506 11390 -1502 11460
rect -1482 11390 -1478 11460
rect -1458 11390 -1454 11460
rect -1434 11390 -1430 11460
rect -1410 11390 -1406 11460
rect -1386 11390 -1382 11460
rect -1362 11390 -1358 11460
rect -1338 11390 -1334 11460
rect -1314 11390 -1310 11460
rect -1290 11390 -1286 11460
rect -1266 11390 -1262 11460
rect -1242 11390 -1238 11460
rect -1218 11390 -1214 11460
rect -1194 11390 -1190 11460
rect -1170 11390 -1166 11460
rect -1146 11390 -1142 11460
rect -1122 11390 -1118 11460
rect -1098 11390 -1094 11460
rect -1074 11390 -1070 11460
rect -1050 11390 -1046 11460
rect -1026 11390 -1022 11460
rect -1002 11390 -998 11460
rect -978 11390 -974 11460
rect -954 11390 -950 11460
rect -930 11390 -926 11460
rect -906 11390 -902 11460
rect -882 11390 -878 11460
rect -858 11390 -854 11460
rect -834 11390 -830 11460
rect -810 11390 -806 11460
rect -786 11390 -782 11460
rect -762 11390 -758 11460
rect -738 11390 -734 11460
rect -714 11390 -710 11460
rect -690 11390 -686 11460
rect -666 11390 -662 11460
rect -642 11390 -638 11460
rect -618 11390 -614 11460
rect -594 11390 -590 11460
rect -570 11390 -566 11460
rect -546 11390 -542 11460
rect -522 11390 -518 11460
rect -498 11390 -494 11460
rect -474 11390 -470 11460
rect -450 11390 -446 11460
rect -426 11390 -422 11460
rect -402 11390 -398 11460
rect -378 11390 -374 11460
rect -354 11390 -350 11460
rect -330 11390 -326 11460
rect -306 11390 -302 11460
rect -282 11390 -278 11460
rect -258 11390 -254 11460
rect -234 11390 -230 11460
rect -210 11390 -206 11460
rect -186 11390 -182 11460
rect -162 11390 -158 11460
rect -138 11390 -134 11460
rect -114 11390 -110 11460
rect -90 11390 -86 11460
rect -66 11390 -62 11460
rect -42 11390 -38 11460
rect -18 11390 -14 11460
rect 6 11390 10 11460
rect 30 11390 34 11460
rect 54 11390 58 11460
rect 78 11390 82 11460
rect 102 11390 106 11460
rect 126 11390 130 11460
rect 139 11453 144 11460
rect 150 11453 154 11460
rect 149 11439 154 11453
rect 150 11390 154 11439
rect 174 11390 178 11484
rect 198 11390 202 11484
rect 222 11390 226 11484
rect 246 11390 250 11484
rect 270 11390 274 11484
rect 294 11390 298 11484
rect 318 11390 322 11484
rect 342 11390 346 11484
rect 366 11390 370 11484
rect 390 11390 394 11484
rect 414 11390 418 11484
rect 438 11390 442 11484
rect 462 11390 466 11484
rect 486 11390 490 11484
rect 510 11390 514 11484
rect 534 11390 538 11484
rect 558 11390 562 11484
rect 582 11390 586 11484
rect 595 11462 629 11463
rect 630 11462 634 11484
rect 654 11462 658 11484
rect 678 11462 682 11484
rect 702 11462 706 11484
rect 726 11462 730 11484
rect 750 11462 754 11484
rect 774 11462 778 11484
rect 798 11462 802 11484
rect 822 11462 826 11484
rect 846 11462 850 11484
rect 870 11462 874 11484
rect 894 11462 898 11484
rect 918 11462 922 11484
rect 942 11462 946 11484
rect 966 11462 970 11484
rect 990 11462 994 11484
rect 1014 11462 1018 11484
rect 1038 11462 1042 11484
rect 1062 11462 1066 11484
rect 1086 11462 1090 11484
rect 1110 11462 1114 11484
rect 1134 11462 1138 11484
rect 1158 11462 1162 11484
rect 1182 11462 1186 11484
rect 1206 11462 1210 11484
rect 1230 11462 1234 11484
rect 1254 11462 1258 11484
rect 1278 11462 1282 11484
rect 1302 11462 1306 11484
rect 1326 11462 1330 11484
rect 1350 11462 1354 11484
rect 1374 11462 1378 11484
rect 1387 11477 1392 11484
rect 1398 11477 1402 11484
rect 1397 11463 1402 11477
rect 1422 11462 1426 11580
rect 1446 11462 1450 11580
rect 1470 11462 1474 11580
rect 1494 11462 1498 11580
rect 1518 11462 1522 11580
rect 1542 11462 1546 11580
rect 1566 11462 1570 11580
rect 1590 11462 1594 11580
rect 1614 11462 1618 11580
rect 1638 11462 1642 11580
rect 1662 11555 1666 11580
rect 1662 11510 1669 11555
rect 1686 11510 1690 11580
rect 1710 11510 1714 11580
rect 1734 11510 1738 11580
rect 1758 11510 1762 11580
rect 1782 11510 1786 11580
rect 1806 11510 1810 11580
rect 1830 11510 1834 11580
rect 1854 11510 1858 11580
rect 1878 11510 1882 11580
rect 1902 11510 1906 11580
rect 1926 11510 1930 11580
rect 1950 11510 1954 11580
rect 1974 11510 1978 11580
rect 1998 11510 2002 11580
rect 2022 11510 2026 11580
rect 2046 11510 2050 11580
rect 2070 11510 2074 11580
rect 2094 11510 2098 11580
rect 2118 11510 2122 11580
rect 2142 11510 2146 11580
rect 2166 11510 2170 11580
rect 2190 11510 2194 11580
rect 2214 11510 2218 11580
rect 2238 11510 2242 11580
rect 2262 11510 2266 11580
rect 2286 11510 2290 11580
rect 2310 11510 2314 11580
rect 2334 11510 2338 11580
rect 2358 11510 2362 11580
rect 2382 11510 2386 11580
rect 2406 11510 2410 11580
rect 2430 11510 2434 11580
rect 2454 11510 2458 11580
rect 2478 11510 2482 11580
rect 2502 11510 2506 11580
rect 2526 11510 2530 11580
rect 2550 11510 2554 11580
rect 2574 11510 2578 11580
rect 2598 11510 2602 11580
rect 2622 11510 2626 11580
rect 2646 11510 2650 11580
rect 2670 11510 2674 11580
rect 2694 11510 2698 11580
rect 2718 11510 2722 11580
rect 2742 11510 2746 11580
rect 2766 11510 2770 11580
rect 2790 11510 2794 11580
rect 2814 11510 2818 11580
rect 2838 11510 2842 11580
rect 2862 11510 2866 11580
rect 2886 11510 2890 11580
rect 2910 11510 2914 11580
rect 2934 11510 2938 11580
rect 2958 11510 2962 11580
rect 2982 11510 2986 11580
rect 3006 11510 3010 11580
rect 3030 11510 3034 11580
rect 3054 11510 3058 11580
rect 3078 11510 3082 11580
rect 3102 11510 3106 11580
rect 3126 11510 3130 11580
rect 3150 11510 3154 11580
rect 3163 11573 3168 11580
rect 3174 11573 3178 11580
rect 3173 11559 3178 11573
rect 3163 11549 3168 11559
rect 3173 11535 3178 11549
rect 3174 11511 3178 11535
rect 3163 11510 3197 11511
rect 1645 11508 3197 11510
rect 1645 11507 1659 11508
rect 1662 11507 1669 11508
rect 1662 11462 1666 11507
rect 1686 11462 1690 11508
rect 1710 11462 1714 11508
rect 1734 11462 1738 11508
rect 1758 11462 1762 11508
rect 1782 11462 1786 11508
rect 1806 11462 1810 11508
rect 1830 11462 1834 11508
rect 1854 11462 1858 11508
rect 1878 11462 1882 11508
rect 1902 11462 1906 11508
rect 1926 11462 1930 11508
rect 1950 11462 1954 11508
rect 1974 11462 1978 11508
rect 1998 11462 2002 11508
rect 2022 11462 2026 11508
rect 2046 11462 2050 11508
rect 2070 11462 2074 11508
rect 2094 11462 2098 11508
rect 2118 11462 2122 11508
rect 2142 11462 2146 11508
rect 2166 11462 2170 11508
rect 2190 11462 2194 11508
rect 2214 11462 2218 11508
rect 2238 11462 2242 11508
rect 2262 11462 2266 11508
rect 2286 11462 2290 11508
rect 2310 11462 2314 11508
rect 2334 11462 2338 11508
rect 2358 11462 2362 11508
rect 2382 11462 2386 11508
rect 2406 11462 2410 11508
rect 2430 11462 2434 11508
rect 2454 11462 2458 11508
rect 2478 11462 2482 11508
rect 2502 11462 2506 11508
rect 2526 11462 2530 11508
rect 2550 11462 2554 11508
rect 2574 11462 2578 11508
rect 2598 11462 2602 11508
rect 2622 11462 2626 11508
rect 2646 11462 2650 11508
rect 2670 11462 2674 11508
rect 2694 11462 2698 11508
rect 2718 11462 2722 11508
rect 2742 11462 2746 11508
rect 2766 11462 2770 11508
rect 2790 11462 2794 11508
rect 2814 11462 2818 11508
rect 2838 11462 2842 11508
rect 2862 11462 2866 11508
rect 2886 11462 2890 11508
rect 2910 11462 2914 11508
rect 2934 11462 2938 11508
rect 2958 11462 2962 11508
rect 2982 11462 2986 11508
rect 3006 11462 3010 11508
rect 3030 11462 3034 11508
rect 3054 11462 3058 11508
rect 3078 11462 3082 11508
rect 3102 11462 3106 11508
rect 3126 11462 3130 11508
rect 3150 11463 3154 11508
rect 3163 11501 3168 11508
rect 3174 11501 3178 11508
rect 3173 11487 3178 11501
rect 3187 11497 3195 11501
rect 3181 11487 3187 11497
rect 3139 11462 3173 11463
rect 595 11460 3173 11462
rect 595 11453 600 11460
rect 605 11439 610 11453
rect 606 11390 610 11439
rect 630 11435 634 11460
rect 630 11411 637 11435
rect 654 11390 658 11460
rect 678 11390 682 11460
rect 702 11390 706 11460
rect 726 11390 730 11460
rect 750 11390 754 11460
rect 774 11390 778 11460
rect 798 11390 802 11460
rect 822 11390 826 11460
rect 846 11390 850 11460
rect 870 11459 874 11460
rect 870 11411 877 11459
rect 870 11390 874 11411
rect 894 11390 898 11460
rect 918 11390 922 11460
rect 942 11390 946 11460
rect 966 11390 970 11460
rect 990 11390 994 11460
rect 1014 11390 1018 11460
rect 1038 11390 1042 11460
rect 1062 11390 1066 11460
rect 1086 11390 1090 11460
rect 1110 11390 1114 11460
rect 1134 11390 1138 11460
rect 1158 11390 1162 11460
rect 1182 11390 1186 11460
rect 1206 11390 1210 11460
rect 1230 11390 1234 11460
rect 1254 11390 1258 11460
rect 1278 11390 1282 11460
rect 1302 11390 1306 11460
rect 1326 11390 1330 11460
rect 1350 11390 1354 11460
rect 1374 11390 1378 11460
rect 1387 11429 1392 11439
rect 1397 11415 1402 11429
rect 1398 11390 1402 11415
rect 1422 11411 1426 11460
rect -2393 11388 1419 11390
rect -2371 11294 -2366 11388
rect -2348 11294 -2343 11388
rect -2325 11326 -2320 11388
rect -2317 11386 -2309 11388
rect -2013 11386 -1992 11388
rect -1663 11386 -1655 11388
rect -2000 11385 -1983 11386
rect -2026 11376 -2021 11380
rect -2062 11375 -2061 11376
rect -2309 11364 -2301 11374
rect -2091 11368 -2061 11375
rect -2317 11358 -2309 11364
rect -2132 11359 -2131 11361
rect -2101 11359 -2092 11361
rect -2091 11360 -2071 11366
rect -2062 11364 -2045 11368
rect -2036 11364 -2031 11366
rect -2292 11350 -2071 11359
rect -2107 11345 -2104 11349
rect -2325 11318 -2317 11326
rect -2325 11298 -2320 11318
rect -2317 11310 -2309 11318
rect -2325 11294 -2317 11298
rect -2000 11294 -1992 11385
rect -1980 11368 -1932 11375
rect -1655 11364 -1647 11374
rect -1846 11350 -1680 11359
rect -1663 11358 -1655 11364
rect -1671 11318 -1663 11326
rect -1663 11310 -1655 11318
rect -1671 11294 -1663 11298
rect -1642 11294 -1637 11388
rect -1619 11294 -1614 11388
rect -1530 11294 -1526 11388
rect -1506 11294 -1502 11388
rect -1482 11294 -1478 11388
rect -1458 11294 -1454 11388
rect -1434 11294 -1430 11388
rect -1410 11294 -1406 11388
rect -1386 11294 -1382 11388
rect -1362 11294 -1358 11388
rect -1338 11294 -1334 11388
rect -1314 11294 -1310 11388
rect -1290 11294 -1286 11388
rect -1266 11294 -1262 11388
rect -1242 11294 -1238 11388
rect -1218 11294 -1214 11388
rect -1194 11294 -1190 11388
rect -1170 11294 -1166 11388
rect -1146 11294 -1142 11388
rect -1122 11294 -1118 11388
rect -1098 11294 -1094 11388
rect -1074 11294 -1070 11388
rect -1050 11294 -1046 11388
rect -1026 11294 -1022 11388
rect -1002 11294 -998 11388
rect -978 11294 -974 11388
rect -954 11294 -950 11388
rect -930 11294 -926 11388
rect -906 11294 -902 11388
rect -882 11294 -878 11388
rect -858 11294 -854 11388
rect -834 11294 -830 11388
rect -810 11294 -806 11388
rect -786 11294 -782 11388
rect -762 11294 -758 11388
rect -738 11294 -734 11388
rect -714 11294 -710 11388
rect -690 11294 -686 11388
rect -666 11294 -662 11388
rect -642 11294 -638 11388
rect -618 11294 -614 11388
rect -594 11294 -590 11388
rect -570 11294 -566 11388
rect -546 11294 -542 11388
rect -522 11294 -518 11388
rect -498 11294 -494 11388
rect -474 11294 -470 11388
rect -450 11294 -446 11388
rect -426 11294 -422 11388
rect -402 11294 -398 11388
rect -378 11294 -374 11388
rect -354 11294 -350 11388
rect -330 11294 -326 11388
rect -306 11294 -302 11388
rect -282 11294 -278 11388
rect -258 11294 -254 11388
rect -234 11294 -230 11388
rect -210 11294 -206 11388
rect -186 11294 -182 11388
rect -162 11294 -158 11388
rect -138 11294 -134 11388
rect -114 11294 -110 11388
rect -90 11294 -86 11388
rect -66 11294 -62 11388
rect -42 11294 -38 11388
rect -18 11294 -14 11388
rect 6 11294 10 11388
rect 30 11294 34 11388
rect 54 11294 58 11388
rect 78 11294 82 11388
rect 102 11294 106 11388
rect 126 11294 130 11388
rect 150 11294 154 11388
rect 174 11387 178 11388
rect 174 11363 181 11387
rect 174 11294 178 11363
rect 198 11294 202 11388
rect 222 11294 226 11388
rect 246 11294 250 11388
rect 270 11294 274 11388
rect 294 11294 298 11388
rect 318 11294 322 11388
rect 342 11294 346 11388
rect 366 11294 370 11388
rect 390 11294 394 11388
rect 414 11294 418 11388
rect 438 11294 442 11388
rect 462 11294 466 11388
rect 486 11294 490 11388
rect 510 11294 514 11388
rect 534 11294 538 11388
rect 558 11294 562 11388
rect 582 11294 586 11388
rect 606 11294 610 11388
rect 630 11363 637 11387
rect 630 11294 634 11363
rect 654 11294 658 11388
rect 678 11294 682 11388
rect 702 11294 706 11388
rect 726 11294 730 11388
rect 750 11294 754 11388
rect 774 11294 778 11388
rect 798 11294 802 11388
rect 822 11294 826 11388
rect 846 11294 850 11388
rect 870 11294 874 11388
rect 894 11294 898 11388
rect 918 11294 922 11388
rect 942 11294 946 11388
rect 966 11294 970 11388
rect 990 11294 994 11388
rect 1014 11294 1018 11388
rect 1038 11294 1042 11388
rect 1062 11294 1066 11388
rect 1086 11294 1090 11388
rect 1110 11294 1114 11388
rect 1134 11294 1138 11388
rect 1158 11294 1162 11388
rect 1182 11294 1186 11388
rect 1206 11294 1210 11388
rect 1230 11294 1234 11388
rect 1254 11294 1258 11388
rect 1278 11294 1282 11388
rect 1302 11294 1306 11388
rect 1326 11294 1330 11388
rect 1350 11294 1354 11388
rect 1374 11294 1378 11388
rect 1398 11294 1402 11388
rect 1405 11387 1419 11388
rect 1422 11387 1429 11411
rect 1422 11342 1429 11363
rect 1446 11342 1450 11460
rect 1470 11342 1474 11460
rect 1494 11342 1498 11460
rect 1518 11342 1522 11460
rect 1542 11342 1546 11460
rect 1566 11342 1570 11460
rect 1590 11342 1594 11460
rect 1614 11342 1618 11460
rect 1638 11342 1642 11460
rect 1662 11342 1666 11460
rect 1686 11342 1690 11460
rect 1710 11342 1714 11460
rect 1734 11342 1738 11460
rect 1758 11342 1762 11460
rect 1782 11342 1786 11460
rect 1806 11342 1810 11460
rect 1830 11342 1834 11460
rect 1854 11342 1858 11460
rect 1878 11342 1882 11460
rect 1902 11342 1906 11460
rect 1926 11342 1930 11460
rect 1950 11342 1954 11460
rect 1974 11342 1978 11460
rect 1998 11342 2002 11460
rect 2022 11342 2026 11460
rect 2046 11342 2050 11460
rect 2070 11342 2074 11460
rect 2094 11342 2098 11460
rect 2118 11342 2122 11460
rect 2142 11342 2146 11460
rect 2166 11342 2170 11460
rect 2190 11342 2194 11460
rect 2214 11342 2218 11460
rect 2238 11342 2242 11460
rect 2262 11342 2266 11460
rect 2286 11342 2290 11460
rect 2310 11342 2314 11460
rect 2334 11342 2338 11460
rect 2358 11342 2362 11460
rect 2382 11342 2386 11460
rect 2406 11342 2410 11460
rect 2430 11342 2434 11460
rect 2454 11342 2458 11460
rect 2478 11342 2482 11460
rect 2502 11342 2506 11460
rect 2526 11342 2530 11460
rect 2550 11343 2554 11460
rect 2539 11342 2573 11343
rect 1405 11340 2573 11342
rect 1405 11339 1419 11340
rect 1422 11339 1429 11340
rect 1422 11294 1426 11339
rect 1446 11294 1450 11340
rect 1470 11294 1474 11340
rect 1494 11294 1498 11340
rect 1518 11294 1522 11340
rect 1542 11294 1546 11340
rect 1566 11294 1570 11340
rect 1590 11294 1594 11340
rect 1614 11294 1618 11340
rect 1638 11294 1642 11340
rect 1662 11294 1666 11340
rect 1686 11294 1690 11340
rect 1710 11294 1714 11340
rect 1734 11294 1738 11340
rect 1758 11294 1762 11340
rect 1782 11294 1786 11340
rect 1806 11294 1810 11340
rect 1830 11294 1834 11340
rect 1854 11294 1858 11340
rect 1878 11294 1882 11340
rect 1902 11294 1906 11340
rect 1926 11294 1930 11340
rect 1950 11294 1954 11340
rect 1974 11294 1978 11340
rect 1998 11294 2002 11340
rect 2022 11294 2026 11340
rect 2046 11294 2050 11340
rect 2070 11294 2074 11340
rect 2094 11294 2098 11340
rect 2118 11294 2122 11340
rect 2142 11294 2146 11340
rect 2166 11294 2170 11340
rect 2190 11294 2194 11340
rect 2214 11294 2218 11340
rect 2238 11294 2242 11340
rect 2262 11294 2266 11340
rect 2286 11294 2290 11340
rect 2310 11294 2314 11340
rect 2334 11294 2338 11340
rect 2358 11294 2362 11340
rect 2382 11294 2386 11340
rect 2406 11294 2410 11340
rect 2430 11294 2434 11340
rect 2454 11294 2458 11340
rect 2478 11294 2482 11340
rect 2502 11294 2506 11340
rect 2526 11294 2530 11340
rect 2539 11333 2544 11340
rect 2550 11333 2554 11340
rect 2549 11319 2554 11333
rect 2539 11309 2544 11319
rect 2549 11295 2554 11309
rect 2550 11294 2554 11295
rect 2574 11294 2578 11460
rect 2598 11294 2602 11460
rect 2622 11294 2626 11460
rect 2646 11294 2650 11460
rect 2670 11294 2674 11460
rect 2694 11294 2698 11460
rect 2718 11294 2722 11460
rect 2742 11294 2746 11460
rect 2766 11294 2770 11460
rect 2790 11294 2794 11460
rect 2814 11294 2818 11460
rect 2838 11294 2842 11460
rect 2862 11294 2866 11460
rect 2886 11294 2890 11460
rect 2910 11294 2914 11460
rect 2934 11294 2938 11460
rect 2958 11294 2962 11460
rect 2982 11294 2986 11460
rect 3006 11294 3010 11460
rect 3030 11294 3034 11460
rect 3054 11294 3058 11460
rect 3078 11294 3082 11460
rect 3102 11294 3106 11460
rect 3115 11429 3120 11439
rect 3126 11429 3130 11460
rect 3139 11453 3144 11460
rect 3150 11453 3154 11460
rect 3149 11439 3154 11453
rect 3125 11415 3130 11429
rect 3115 11381 3120 11391
rect 3125 11367 3130 11381
rect 3115 11309 3120 11319
rect 3126 11309 3130 11367
rect 3125 11295 3130 11309
rect 3139 11305 3147 11309
rect 3133 11295 3139 11305
rect 3115 11294 3147 11295
rect -2393 11292 -1969 11294
rect -1955 11292 3147 11294
rect -2371 11246 -2366 11292
rect -2348 11246 -2343 11292
rect -2325 11282 -2317 11292
rect -2080 11290 -1969 11292
rect -2080 11284 -2053 11290
rect -2325 11266 -2320 11282
rect -2309 11270 -2301 11282
rect -2070 11275 -2040 11282
rect -2000 11274 -1992 11290
rect -1972 11286 -1969 11290
rect -1972 11284 -1955 11286
rect -1955 11274 -1850 11283
rect -1671 11282 -1663 11292
rect -2317 11266 -2309 11270
rect -2070 11267 -2053 11273
rect -2027 11272 -1992 11274
rect -1969 11272 -1955 11273
rect -2325 11254 -2317 11266
rect -2292 11257 -2053 11266
rect -2325 11246 -2320 11254
rect -2309 11246 -2301 11254
rect -2000 11246 -1992 11272
rect -1655 11270 -1647 11282
rect -1663 11266 -1655 11270
rect -1972 11258 -1924 11265
rect -1945 11257 -1929 11258
rect -1860 11257 -1680 11266
rect -1671 11254 -1663 11266
rect -1978 11246 -1942 11247
rect -1655 11246 -1647 11254
rect -1642 11246 -1637 11292
rect -1619 11246 -1614 11292
rect -1530 11246 -1526 11292
rect -1506 11246 -1502 11292
rect -1482 11246 -1478 11292
rect -1458 11246 -1454 11292
rect -1434 11246 -1430 11292
rect -1410 11246 -1406 11292
rect -1386 11246 -1382 11292
rect -1362 11246 -1358 11292
rect -1338 11246 -1334 11292
rect -1314 11246 -1310 11292
rect -1290 11246 -1286 11292
rect -1266 11246 -1262 11292
rect -1242 11246 -1238 11292
rect -1218 11246 -1214 11292
rect -1194 11246 -1190 11292
rect -1170 11247 -1166 11292
rect -1181 11246 -1147 11247
rect -2393 11244 -1147 11246
rect -2371 11126 -2366 11244
rect -2348 11126 -2343 11244
rect -2325 11238 -2320 11244
rect -2309 11242 -2301 11244
rect -2317 11238 -2309 11242
rect -2325 11226 -2317 11238
rect -2325 11206 -2320 11226
rect -2062 11206 -2032 11207
rect -2000 11206 -1992 11244
rect -1655 11242 -1647 11244
rect -1663 11238 -1655 11242
rect -1671 11226 -1663 11238
rect -1942 11208 -1937 11220
rect -1850 11217 -1822 11218
rect -1850 11213 -1802 11217
rect -2325 11198 -2317 11206
rect -2062 11204 -1961 11206
rect -2325 11178 -2320 11198
rect -2317 11190 -2309 11198
rect -2062 11191 -2040 11202
rect -2032 11197 -1961 11204
rect -1947 11198 -1942 11206
rect -1842 11204 -1794 11207
rect -2070 11186 -2022 11190
rect -2325 11162 -2317 11178
rect -2080 11164 -2032 11173
rect -2325 11146 -2320 11162
rect -2309 11150 -2301 11162
rect -2070 11155 -2040 11162
rect -2317 11146 -2309 11150
rect -2325 11134 -2317 11146
rect -2000 11145 -1992 11197
rect -1942 11196 -1937 11198
rect -1932 11188 -1927 11196
rect -1912 11193 -1896 11199
rect -1842 11191 -1802 11202
rect -1671 11198 -1663 11206
rect -1663 11190 -1655 11198
rect -1850 11186 -1680 11190
rect -1937 11172 -1934 11174
rect -1924 11172 -1921 11174
rect -1850 11164 -1842 11174
rect -1840 11164 -1792 11173
rect -1924 11162 -1850 11163
rect -1671 11162 -1663 11178
rect -1960 11160 -1955 11161
rect -1969 11154 -1955 11160
rect -1924 11155 -1802 11162
rect -1924 11154 -1850 11155
rect -1969 11152 -1944 11154
rect -1955 11145 -1944 11152
rect -1842 11147 -1802 11153
rect -1655 11150 -1647 11162
rect -1663 11146 -1655 11150
rect -1860 11145 -1794 11146
rect -2040 11138 -1945 11145
rect -1929 11143 -1794 11145
rect -1929 11138 -1850 11143
rect -2325 11126 -2320 11134
rect -2309 11126 -2301 11134
rect -2070 11128 -2040 11135
rect -2000 11126 -1992 11138
rect -1842 11137 -1794 11143
rect -1945 11128 -1942 11130
rect -1850 11128 -1802 11135
rect -1671 11134 -1663 11146
rect -1978 11126 -1942 11127
rect -1655 11126 -1647 11134
rect -1642 11126 -1637 11244
rect -1619 11126 -1614 11244
rect -1530 11126 -1526 11244
rect -1506 11126 -1502 11244
rect -1482 11126 -1478 11244
rect -1458 11126 -1454 11244
rect -1434 11126 -1430 11244
rect -1410 11126 -1406 11244
rect -1386 11126 -1382 11244
rect -1362 11126 -1358 11244
rect -1338 11126 -1334 11244
rect -1314 11126 -1310 11244
rect -1290 11126 -1286 11244
rect -1266 11126 -1262 11244
rect -1242 11126 -1238 11244
rect -1218 11126 -1214 11244
rect -1194 11126 -1190 11244
rect -1181 11237 -1176 11244
rect -1170 11237 -1166 11244
rect -1171 11223 -1166 11237
rect -1170 11126 -1166 11223
rect -1146 11171 -1142 11292
rect -1146 11147 -1139 11171
rect -1146 11126 -1142 11147
rect -1122 11126 -1118 11292
rect -1098 11126 -1094 11292
rect -1074 11126 -1070 11292
rect -1050 11126 -1046 11292
rect -1026 11126 -1022 11292
rect -1002 11126 -998 11292
rect -978 11126 -974 11292
rect -954 11126 -950 11292
rect -930 11126 -926 11292
rect -906 11126 -902 11292
rect -882 11126 -878 11292
rect -858 11126 -854 11292
rect -834 11126 -830 11292
rect -810 11126 -806 11292
rect -786 11126 -782 11292
rect -762 11126 -758 11292
rect -738 11126 -734 11292
rect -714 11126 -710 11292
rect -690 11126 -686 11292
rect -666 11126 -662 11292
rect -642 11126 -638 11292
rect -618 11126 -614 11292
rect -594 11126 -590 11292
rect -570 11126 -566 11292
rect -546 11126 -542 11292
rect -522 11126 -518 11292
rect -498 11126 -494 11292
rect -474 11126 -470 11292
rect -450 11126 -446 11292
rect -426 11126 -422 11292
rect -402 11126 -398 11292
rect -378 11126 -374 11292
rect -354 11126 -350 11292
rect -330 11126 -326 11292
rect -306 11126 -302 11292
rect -282 11126 -278 11292
rect -258 11126 -254 11292
rect -234 11126 -230 11292
rect -210 11126 -206 11292
rect -186 11126 -182 11292
rect -162 11126 -158 11292
rect -138 11126 -134 11292
rect -114 11126 -110 11292
rect -90 11126 -86 11292
rect -66 11126 -62 11292
rect -42 11126 -38 11292
rect -18 11126 -14 11292
rect 6 11126 10 11292
rect 30 11126 34 11292
rect 54 11126 58 11292
rect 78 11126 82 11292
rect 102 11126 106 11292
rect 126 11126 130 11292
rect 150 11126 154 11292
rect 174 11126 178 11292
rect 198 11126 202 11292
rect 222 11126 226 11292
rect 246 11126 250 11292
rect 270 11126 274 11292
rect 294 11126 298 11292
rect 318 11126 322 11292
rect 342 11126 346 11292
rect 366 11126 370 11292
rect 390 11126 394 11292
rect 414 11126 418 11292
rect 438 11126 442 11292
rect 462 11126 466 11292
rect 486 11126 490 11292
rect 510 11126 514 11292
rect 534 11126 538 11292
rect 558 11126 562 11292
rect 582 11126 586 11292
rect 606 11126 610 11292
rect 630 11126 634 11292
rect 654 11126 658 11292
rect 678 11126 682 11292
rect 702 11126 706 11292
rect 726 11126 730 11292
rect 750 11126 754 11292
rect 774 11126 778 11292
rect 798 11126 802 11292
rect 822 11126 826 11292
rect 846 11126 850 11292
rect 870 11126 874 11292
rect 894 11126 898 11292
rect 918 11126 922 11292
rect 942 11126 946 11292
rect 966 11126 970 11292
rect 990 11126 994 11292
rect 1014 11126 1018 11292
rect 1038 11126 1042 11292
rect 1062 11126 1066 11292
rect 1086 11126 1090 11292
rect 1110 11126 1114 11292
rect 1134 11126 1138 11292
rect 1158 11126 1162 11292
rect 1182 11126 1186 11292
rect 1206 11126 1210 11292
rect 1230 11126 1234 11292
rect 1254 11126 1258 11292
rect 1278 11126 1282 11292
rect 1302 11126 1306 11292
rect 1326 11126 1330 11292
rect 1350 11126 1354 11292
rect 1374 11126 1378 11292
rect 1398 11126 1402 11292
rect 1422 11126 1426 11292
rect 1446 11126 1450 11292
rect 1470 11126 1474 11292
rect 1483 11213 1488 11223
rect 1494 11213 1498 11292
rect 1493 11199 1498 11213
rect 1483 11198 1517 11199
rect 1518 11198 1522 11292
rect 1542 11198 1546 11292
rect 1566 11198 1570 11292
rect 1590 11198 1594 11292
rect 1614 11198 1618 11292
rect 1638 11198 1642 11292
rect 1662 11198 1666 11292
rect 1686 11198 1690 11292
rect 1710 11198 1714 11292
rect 1734 11198 1738 11292
rect 1758 11198 1762 11292
rect 1782 11198 1786 11292
rect 1806 11198 1810 11292
rect 1830 11198 1834 11292
rect 1854 11198 1858 11292
rect 1878 11198 1882 11292
rect 1902 11198 1906 11292
rect 1926 11198 1930 11292
rect 1950 11198 1954 11292
rect 1974 11198 1978 11292
rect 1998 11198 2002 11292
rect 2022 11198 2026 11292
rect 2046 11198 2050 11292
rect 2070 11198 2074 11292
rect 2094 11198 2098 11292
rect 2118 11198 2122 11292
rect 2142 11198 2146 11292
rect 2166 11198 2170 11292
rect 2190 11198 2194 11292
rect 2214 11198 2218 11292
rect 2238 11198 2242 11292
rect 2262 11198 2266 11292
rect 2286 11198 2290 11292
rect 2310 11198 2314 11292
rect 2334 11198 2338 11292
rect 2358 11198 2362 11292
rect 2382 11198 2386 11292
rect 2406 11198 2410 11292
rect 2430 11198 2434 11292
rect 2454 11198 2458 11292
rect 2478 11198 2482 11292
rect 2502 11198 2506 11292
rect 2526 11198 2530 11292
rect 2550 11198 2554 11292
rect 2574 11267 2578 11292
rect 2574 11219 2581 11267
rect 2574 11198 2578 11219
rect 2598 11198 2602 11292
rect 2622 11198 2626 11292
rect 2646 11198 2650 11292
rect 2670 11198 2674 11292
rect 2694 11198 2698 11292
rect 2718 11198 2722 11292
rect 2742 11198 2746 11292
rect 2766 11198 2770 11292
rect 2790 11198 2794 11292
rect 2814 11198 2818 11292
rect 2838 11198 2842 11292
rect 2862 11198 2866 11292
rect 2886 11198 2890 11292
rect 2910 11198 2914 11292
rect 2934 11198 2938 11292
rect 2958 11198 2962 11292
rect 2982 11198 2986 11292
rect 3006 11198 3010 11292
rect 3030 11198 3034 11292
rect 3054 11198 3058 11292
rect 3078 11198 3082 11292
rect 3102 11198 3106 11292
rect 3115 11285 3120 11292
rect 3133 11291 3147 11292
rect 3125 11271 3130 11285
rect 3126 11199 3130 11271
rect 3115 11198 3147 11199
rect 1483 11196 3147 11198
rect 1483 11189 1488 11196
rect 1493 11175 1498 11189
rect 1494 11126 1498 11175
rect 1518 11147 1522 11196
rect -2393 11124 1515 11126
rect -2371 11030 -2366 11124
rect -2348 11030 -2343 11124
rect -2325 11118 -2320 11124
rect -2309 11122 -2301 11124
rect -2317 11118 -2309 11122
rect -2062 11120 -2040 11124
rect -2325 11106 -2317 11118
rect -2062 11111 -2032 11118
rect -2325 11086 -2320 11106
rect -2062 11086 -2032 11087
rect -2000 11086 -1992 11124
rect -1888 11119 -1874 11124
rect -1842 11120 -1802 11124
rect -1655 11122 -1647 11124
rect -1932 11110 -1924 11119
rect -1904 11117 -1874 11119
rect -1842 11110 -1792 11119
rect -1663 11118 -1655 11122
rect -1671 11106 -1663 11118
rect -1942 11088 -1937 11100
rect -1850 11097 -1822 11098
rect -1850 11093 -1802 11097
rect -2325 11078 -2317 11086
rect -2062 11084 -1961 11086
rect -2325 11058 -2320 11078
rect -2317 11070 -2309 11078
rect -2062 11071 -2040 11082
rect -2032 11077 -1961 11084
rect -1947 11078 -1942 11086
rect -1842 11084 -1794 11087
rect -2070 11066 -2022 11070
rect -2325 11046 -2317 11058
rect -2325 11030 -2320 11046
rect -2317 11042 -2309 11046
rect -2309 11030 -2301 11042
rect -2068 11035 -2038 11042
rect -2000 11032 -1992 11077
rect -1942 11076 -1937 11078
rect -1932 11068 -1927 11076
rect -1912 11073 -1896 11079
rect -1842 11071 -1802 11082
rect -1671 11078 -1663 11086
rect -1663 11070 -1655 11078
rect -1850 11066 -1680 11070
rect -1937 11052 -1934 11054
rect -1926 11052 -1921 11057
rect -1926 11047 -1924 11052
rect -1916 11044 -1914 11047
rect -1842 11044 -1794 11053
rect -1671 11046 -1663 11058
rect -1924 11034 -1916 11043
rect -1663 11042 -1655 11046
rect -1852 11035 -1804 11042
rect -1916 11033 -1914 11034
rect -2025 11031 -1991 11032
rect -2025 11030 -1975 11031
rect -1842 11030 -1804 11033
rect -1655 11030 -1647 11042
rect -1642 11030 -1637 11124
rect -1619 11030 -1614 11124
rect -1530 11030 -1526 11124
rect -1506 11030 -1502 11124
rect -1482 11030 -1478 11124
rect -1458 11030 -1454 11124
rect -1434 11030 -1430 11124
rect -1410 11030 -1406 11124
rect -1386 11031 -1382 11124
rect -1397 11030 -1363 11031
rect -2393 11028 -1363 11030
rect -2371 11006 -2366 11028
rect -2348 11006 -2343 11028
rect -2325 11018 -2317 11028
rect -2076 11018 -2068 11025
rect -2062 11018 -2001 11025
rect -2325 11006 -2320 11018
rect -2317 11014 -2309 11018
rect -2015 11017 -2001 11018
rect -2309 11006 -2301 11014
rect -2068 11008 -2062 11015
rect -2000 11010 -1992 11028
rect -1974 11026 -1960 11028
rect -1842 11027 -1804 11028
rect -1862 11025 -1794 11026
rect -1985 11023 -1794 11025
rect -1985 11018 -1852 11023
rect -1842 11017 -1794 11023
rect -1671 11018 -1663 11028
rect -2015 11008 -1985 11010
rect -1852 11008 -1804 11015
rect -1663 11014 -1655 11018
rect -2000 11006 -1992 11008
rect -1976 11006 -1940 11007
rect -1655 11006 -1647 11014
rect -1642 11006 -1637 11028
rect -1619 11006 -1614 11028
rect -1530 11006 -1526 11028
rect -1506 11006 -1502 11028
rect -1482 11006 -1478 11028
rect -1458 11006 -1454 11028
rect -1434 11006 -1430 11028
rect -1410 11006 -1406 11028
rect -1397 11021 -1392 11028
rect -1386 11021 -1382 11028
rect -1387 11007 -1382 11021
rect -1386 11006 -1382 11007
rect -1362 11006 -1358 11124
rect -1338 11006 -1334 11124
rect -1314 11006 -1310 11124
rect -1290 11006 -1286 11124
rect -1266 11006 -1262 11124
rect -1242 11006 -1238 11124
rect -1218 11006 -1214 11124
rect -1194 11006 -1190 11124
rect -1170 11006 -1166 11124
rect -1146 11006 -1142 11124
rect -1122 11006 -1118 11124
rect -1098 11006 -1094 11124
rect -1074 11006 -1070 11124
rect -1050 11006 -1046 11124
rect -1026 11006 -1022 11124
rect -1002 11006 -998 11124
rect -978 11006 -974 11124
rect -954 11006 -950 11124
rect -930 11006 -926 11124
rect -906 11006 -902 11124
rect -882 11006 -878 11124
rect -858 11006 -854 11124
rect -834 11006 -830 11124
rect -810 11006 -806 11124
rect -786 11006 -782 11124
rect -762 11006 -758 11124
rect -738 11006 -734 11124
rect -714 11006 -710 11124
rect -690 11006 -686 11124
rect -666 11006 -662 11124
rect -653 11093 -648 11103
rect -642 11093 -638 11124
rect -643 11079 -638 11093
rect -642 11006 -638 11079
rect -618 11027 -614 11124
rect -2393 11004 -621 11006
rect -2371 10934 -2366 11004
rect -2348 10934 -2343 11004
rect -2325 11002 -2320 11004
rect -2309 11002 -2301 11004
rect -2325 10990 -2317 11002
rect -2062 10991 -2032 10998
rect -2325 10970 -2320 10990
rect -2317 10986 -2309 10990
rect -2325 10962 -2317 10970
rect -2060 10964 -2030 10967
rect -2325 10942 -2320 10962
rect -2317 10954 -2309 10962
rect -2060 10951 -2038 10962
rect -2033 10955 -2030 10964
rect -2028 10960 -2027 10964
rect -2068 10946 -2038 10949
rect -2325 10934 -2317 10942
rect -2000 10937 -1992 11004
rect -1888 10999 -1874 11004
rect -1842 11000 -1804 11004
rect -1655 11002 -1647 11004
rect -1902 10997 -1874 10999
rect -1842 10990 -1794 10999
rect -1671 10990 -1663 11002
rect -1663 10986 -1655 10990
rect -1912 10979 -1884 10981
rect -1852 10973 -1804 10977
rect -1844 10964 -1796 10967
rect -1671 10962 -1663 10970
rect -1844 10951 -1804 10962
rect -1663 10954 -1655 10962
rect -1852 10946 -1680 10950
rect -2119 10934 -2069 10936
rect -2007 10934 -1977 10937
rect -1926 10934 -1892 10937
rect -1671 10934 -1663 10942
rect -1642 10934 -1637 11004
rect -1619 10934 -1614 11004
rect -1530 10934 -1526 11004
rect -1506 10934 -1502 11004
rect -1482 10934 -1478 11004
rect -1458 10934 -1454 11004
rect -1434 10934 -1430 11004
rect -1410 10934 -1406 11004
rect -1386 10934 -1382 11004
rect -1362 10955 -1358 11004
rect -2393 10932 -1365 10934
rect -2371 10910 -2366 10932
rect -2348 10910 -2343 10932
rect -2325 10928 -2317 10932
rect -2325 10912 -2320 10928
rect -2317 10926 -2309 10928
rect -2309 10914 -2301 10926
rect -2000 10918 -1992 10932
rect -1671 10928 -1663 10932
rect -1663 10926 -1655 10928
rect -1844 10924 -1806 10926
rect -1854 10918 -1806 10922
rect -2068 10915 -2060 10918
rect -2030 10915 -1958 10918
rect -1942 10915 -1806 10918
rect -2317 10912 -2309 10914
rect -2000 10912 -1992 10915
rect -1655 10914 -1647 10926
rect -2325 10910 -2317 10912
rect -2033 10910 -1992 10912
rect -1844 10911 -1806 10913
rect -1663 10912 -1655 10914
rect -1864 10910 -1796 10911
rect -1671 10910 -1663 10912
rect -1642 10910 -1637 10932
rect -1619 10910 -1614 10932
rect -1530 10910 -1526 10932
rect -1506 10910 -1502 10932
rect -1482 10910 -1478 10932
rect -1458 10910 -1454 10932
rect -1434 10910 -1430 10932
rect -1410 10910 -1406 10932
rect -1386 10910 -1382 10932
rect -1379 10931 -1365 10932
rect -1362 10931 -1355 10955
rect -1362 10910 -1358 10931
rect -1338 10910 -1334 11004
rect -1314 10910 -1310 11004
rect -1290 10910 -1286 11004
rect -1266 10910 -1262 11004
rect -1242 10910 -1238 11004
rect -1218 10910 -1214 11004
rect -1194 10910 -1190 11004
rect -1170 10910 -1166 11004
rect -1146 10910 -1142 11004
rect -1122 10910 -1118 11004
rect -1098 10910 -1094 11004
rect -1074 10910 -1070 11004
rect -1050 10910 -1046 11004
rect -1026 10910 -1022 11004
rect -1002 10910 -998 11004
rect -978 10910 -974 11004
rect -954 10910 -950 11004
rect -930 10910 -926 11004
rect -906 10910 -902 11004
rect -882 10910 -878 11004
rect -858 10910 -854 11004
rect -834 10910 -830 11004
rect -810 10910 -806 11004
rect -786 10910 -782 11004
rect -762 10910 -758 11004
rect -738 10910 -734 11004
rect -714 10910 -710 11004
rect -690 10910 -686 11004
rect -666 10910 -662 11004
rect -642 10910 -638 11004
rect -635 11003 -621 11004
rect -618 11003 -611 11027
rect -618 10910 -614 11003
rect -594 10910 -590 11124
rect -570 10910 -566 11124
rect -546 10910 -542 11124
rect -533 10973 -528 10983
rect -522 10973 -518 11124
rect -523 10959 -518 10973
rect -522 10910 -518 10959
rect -498 10910 -494 11124
rect -474 10910 -470 11124
rect -450 10910 -446 11124
rect -426 10910 -422 11124
rect -402 10910 -398 11124
rect -378 10910 -374 11124
rect -354 10910 -350 11124
rect -330 10910 -326 11124
rect -306 10910 -302 11124
rect -282 10910 -278 11124
rect -258 10910 -254 11124
rect -234 10910 -230 11124
rect -210 10910 -206 11124
rect -186 10910 -182 11124
rect -162 10910 -158 11124
rect -138 10910 -134 11124
rect -114 10910 -110 11124
rect -90 10910 -86 11124
rect -66 10910 -62 11124
rect -42 10910 -38 11124
rect -18 10911 -14 11124
rect -29 10910 5 10911
rect -2393 10908 5 10910
rect -2371 10886 -2366 10908
rect -2348 10886 -2343 10908
rect -2325 10900 -2317 10908
rect -2060 10905 -2030 10908
rect -2000 10905 -1992 10908
rect -1972 10906 -1958 10908
rect -1904 10905 -1798 10908
rect -2078 10901 -2020 10905
rect -2023 10900 -2020 10901
rect -2000 10903 -1798 10905
rect -2000 10901 -1854 10903
rect -1844 10901 -1798 10903
rect -2325 10886 -2320 10900
rect -2317 10898 -2309 10900
rect -2020 10898 -2004 10900
rect -2000 10898 -1992 10901
rect -1671 10900 -1663 10908
rect -2309 10886 -2301 10898
rect -2020 10896 -1992 10898
rect -1844 10897 -1806 10899
rect -1663 10898 -1655 10900
rect -2023 10891 -1992 10896
rect -1854 10891 -1806 10895
rect -2068 10888 -2060 10891
rect -2030 10888 -1806 10891
rect -2074 10886 -2060 10888
rect -2020 10886 -2004 10888
rect -2000 10886 -1992 10888
rect -1655 10886 -1647 10898
rect -1642 10886 -1637 10908
rect -1619 10886 -1614 10908
rect -1530 10886 -1526 10908
rect -1506 10886 -1502 10908
rect -1482 10886 -1478 10908
rect -1458 10886 -1454 10908
rect -1434 10886 -1430 10908
rect -1410 10886 -1406 10908
rect -1386 10886 -1382 10908
rect -1362 10886 -1358 10908
rect -1338 10886 -1334 10908
rect -1314 10886 -1310 10908
rect -1290 10886 -1286 10908
rect -1266 10886 -1262 10908
rect -1242 10886 -1238 10908
rect -1218 10886 -1214 10908
rect -1194 10886 -1190 10908
rect -1170 10886 -1166 10908
rect -1146 10886 -1142 10908
rect -1122 10886 -1118 10908
rect -1098 10886 -1094 10908
rect -1074 10886 -1070 10908
rect -1050 10886 -1046 10908
rect -1026 10886 -1022 10908
rect -1002 10886 -998 10908
rect -978 10887 -974 10908
rect -989 10886 -955 10887
rect -2393 10884 -2060 10886
rect -2050 10884 -955 10886
rect -2371 10838 -2366 10884
rect -2348 10838 -2343 10884
rect -2325 10872 -2317 10884
rect -2109 10881 -2108 10884
rect -2117 10874 -2108 10881
rect -2325 10852 -2320 10872
rect -2317 10870 -2309 10872
rect -2109 10870 -2108 10874
rect -2060 10874 -2030 10881
rect -2060 10870 -2034 10874
rect -2325 10844 -2317 10852
rect -2101 10847 -2071 10850
rect -2325 10838 -2320 10844
rect -2317 10838 -2309 10844
rect -2000 10842 -1992 10884
rect -1844 10883 -1806 10884
rect -1844 10874 -1798 10881
rect -1671 10872 -1663 10884
rect -1844 10870 -1806 10872
rect -1663 10870 -1655 10872
rect -1854 10856 -1680 10860
rect -1846 10847 -1798 10850
rect -2079 10841 -2043 10842
rect -2007 10841 -1991 10842
rect -2079 10840 -2071 10841
rect -2079 10838 -2029 10840
rect -2011 10838 -1991 10841
rect -1846 10839 -1806 10845
rect -1671 10844 -1663 10852
rect -1864 10838 -1796 10839
rect -1663 10838 -1655 10844
rect -1642 10838 -1637 10884
rect -1619 10838 -1614 10884
rect -1530 10838 -1526 10884
rect -1506 10838 -1502 10884
rect -1482 10838 -1478 10884
rect -1458 10838 -1454 10884
rect -1434 10838 -1430 10884
rect -1410 10838 -1406 10884
rect -1386 10838 -1382 10884
rect -1362 10838 -1358 10884
rect -1338 10838 -1334 10884
rect -1314 10838 -1310 10884
rect -1290 10838 -1286 10884
rect -1266 10838 -1262 10884
rect -1242 10838 -1238 10884
rect -1218 10838 -1214 10884
rect -1194 10838 -1190 10884
rect -1170 10838 -1166 10884
rect -1146 10838 -1142 10884
rect -1122 10838 -1118 10884
rect -1098 10838 -1094 10884
rect -1074 10838 -1070 10884
rect -1050 10838 -1046 10884
rect -1026 10838 -1022 10884
rect -1002 10838 -998 10884
rect -989 10877 -984 10884
rect -978 10877 -974 10884
rect -979 10863 -974 10877
rect -954 10838 -950 10908
rect -930 10838 -926 10908
rect -906 10838 -902 10908
rect -882 10839 -878 10908
rect -893 10838 -859 10839
rect -2393 10836 -859 10838
rect -2371 10790 -2366 10836
rect -2348 10790 -2343 10836
rect -2325 10824 -2320 10836
rect -2079 10834 -2071 10836
rect -2072 10832 -2071 10834
rect -2109 10827 -2101 10832
rect -2101 10825 -2079 10827
rect -2069 10825 -2068 10832
rect -2325 10816 -2317 10824
rect -2079 10820 -2071 10825
rect -2325 10796 -2320 10816
rect -2317 10808 -2309 10816
rect -2074 10811 -2071 10820
rect -2069 10816 -2068 10820
rect -2109 10802 -2079 10805
rect -2325 10790 -2317 10796
rect -2000 10790 -1992 10836
rect -1846 10834 -1806 10836
rect -1854 10829 -1806 10833
rect -1854 10827 -1846 10829
rect -1846 10825 -1806 10827
rect -1806 10823 -1798 10825
rect -1846 10820 -1798 10823
rect -1846 10807 -1806 10818
rect -1671 10816 -1663 10824
rect -1663 10808 -1655 10816
rect -1854 10802 -1680 10806
rect -1671 10790 -1663 10796
rect -1642 10790 -1637 10836
rect -1619 10790 -1614 10836
rect -1530 10790 -1526 10836
rect -1506 10790 -1502 10836
rect -1482 10790 -1478 10836
rect -1458 10790 -1454 10836
rect -1434 10790 -1430 10836
rect -1410 10790 -1406 10836
rect -1386 10790 -1382 10836
rect -1362 10790 -1358 10836
rect -1338 10790 -1334 10836
rect -1314 10790 -1310 10836
rect -1290 10790 -1286 10836
rect -1266 10790 -1262 10836
rect -1242 10790 -1238 10836
rect -1218 10790 -1214 10836
rect -1194 10790 -1190 10836
rect -1170 10790 -1166 10836
rect -1146 10790 -1142 10836
rect -1122 10790 -1118 10836
rect -1098 10790 -1094 10836
rect -1074 10790 -1070 10836
rect -1050 10790 -1046 10836
rect -1026 10790 -1022 10836
rect -1002 10790 -998 10836
rect -989 10814 -955 10815
rect -954 10814 -950 10836
rect -930 10814 -926 10836
rect -906 10814 -902 10836
rect -893 10829 -888 10836
rect -882 10829 -878 10836
rect -883 10815 -878 10829
rect -858 10814 -854 10908
rect -834 10814 -830 10908
rect -810 10814 -806 10908
rect -786 10814 -782 10908
rect -762 10814 -758 10908
rect -738 10814 -734 10908
rect -714 10814 -710 10908
rect -690 10814 -686 10908
rect -666 10814 -662 10908
rect -642 10814 -638 10908
rect -618 10814 -614 10908
rect -594 10814 -590 10908
rect -570 10814 -566 10908
rect -546 10814 -542 10908
rect -522 10814 -518 10908
rect -498 10907 -494 10908
rect -498 10883 -491 10907
rect -498 10814 -494 10883
rect -474 10814 -470 10908
rect -450 10814 -446 10908
rect -426 10814 -422 10908
rect -402 10814 -398 10908
rect -378 10814 -374 10908
rect -354 10814 -350 10908
rect -330 10814 -326 10908
rect -306 10814 -302 10908
rect -282 10814 -278 10908
rect -258 10814 -254 10908
rect -234 10814 -230 10908
rect -210 10814 -206 10908
rect -186 10814 -182 10908
rect -162 10814 -158 10908
rect -138 10814 -134 10908
rect -114 10814 -110 10908
rect -90 10814 -86 10908
rect -66 10814 -62 10908
rect -42 10814 -38 10908
rect -29 10901 -24 10908
rect -18 10901 -14 10908
rect -19 10887 -14 10901
rect -29 10877 -24 10887
rect -19 10863 -14 10877
rect -18 10814 -14 10863
rect 6 10835 10 11124
rect -989 10812 3 10814
rect -989 10805 -984 10812
rect -954 10811 -950 10812
rect -979 10791 -974 10805
rect -965 10801 -957 10805
rect -971 10791 -965 10801
rect -978 10790 -974 10791
rect -2393 10788 -957 10790
rect -2371 10766 -2366 10788
rect -2348 10766 -2343 10788
rect -2325 10780 -2317 10788
rect -2325 10766 -2320 10780
rect -2309 10768 -2301 10780
rect -2092 10771 -2062 10776
rect -2000 10768 -1992 10788
rect -2317 10766 -2309 10768
rect -2000 10766 -1983 10768
rect -1906 10766 -1904 10788
rect -1806 10780 -1680 10786
rect -1671 10780 -1663 10788
rect -1854 10771 -1806 10776
rect -1846 10766 -1806 10769
rect -1655 10768 -1647 10780
rect -1663 10766 -1655 10768
rect -1642 10766 -1637 10788
rect -1619 10766 -1614 10788
rect -1530 10766 -1526 10788
rect -1506 10766 -1502 10788
rect -1482 10766 -1478 10788
rect -1458 10766 -1454 10788
rect -1434 10766 -1430 10788
rect -1410 10766 -1406 10788
rect -1386 10766 -1382 10788
rect -1362 10766 -1358 10788
rect -1338 10766 -1334 10788
rect -1314 10766 -1310 10788
rect -1290 10766 -1286 10788
rect -1266 10766 -1262 10788
rect -1242 10766 -1238 10788
rect -1218 10766 -1214 10788
rect -1194 10766 -1190 10788
rect -1170 10766 -1166 10788
rect -1146 10766 -1142 10788
rect -1122 10766 -1118 10788
rect -1098 10766 -1094 10788
rect -1074 10766 -1070 10788
rect -1050 10766 -1046 10788
rect -1026 10766 -1022 10788
rect -1002 10766 -998 10788
rect -978 10766 -974 10788
rect -971 10787 -957 10788
rect -954 10787 -947 10811
rect -930 10766 -926 10812
rect -906 10766 -902 10812
rect -893 10781 -888 10791
rect -883 10767 -878 10781
rect -882 10766 -878 10767
rect -858 10766 -854 10812
rect -834 10766 -830 10812
rect -810 10766 -806 10812
rect -786 10766 -782 10812
rect -762 10766 -758 10812
rect -738 10766 -734 10812
rect -714 10766 -710 10812
rect -690 10766 -686 10812
rect -666 10766 -662 10812
rect -642 10766 -638 10812
rect -618 10766 -614 10812
rect -594 10766 -590 10812
rect -570 10766 -566 10812
rect -546 10766 -542 10812
rect -522 10766 -518 10812
rect -498 10766 -494 10812
rect -474 10766 -470 10812
rect -450 10766 -446 10812
rect -426 10766 -422 10812
rect -402 10766 -398 10812
rect -378 10766 -374 10812
rect -354 10766 -350 10812
rect -330 10766 -326 10812
rect -306 10766 -302 10812
rect -282 10766 -278 10812
rect -258 10766 -254 10812
rect -234 10766 -230 10812
rect -210 10766 -206 10812
rect -186 10766 -182 10812
rect -162 10766 -158 10812
rect -138 10766 -134 10812
rect -114 10766 -110 10812
rect -90 10766 -86 10812
rect -66 10766 -62 10812
rect -42 10766 -38 10812
rect -18 10766 -14 10812
rect -11 10811 3 10812
rect 6 10787 13 10835
rect 6 10766 10 10787
rect 30 10766 34 11124
rect 54 10766 58 11124
rect 78 10766 82 11124
rect 102 10766 106 11124
rect 126 10766 130 11124
rect 150 10766 154 11124
rect 174 10766 178 11124
rect 198 10766 202 11124
rect 222 10766 226 11124
rect 246 10766 250 11124
rect 270 10766 274 11124
rect 294 10766 298 11124
rect 318 10766 322 11124
rect 342 10766 346 11124
rect 366 10766 370 11124
rect 390 10766 394 11124
rect 414 10766 418 11124
rect 438 10766 442 11124
rect 462 10766 466 11124
rect 486 10766 490 11124
rect 510 10766 514 11124
rect 534 10766 538 11124
rect 558 10766 562 11124
rect 582 10766 586 11124
rect 606 10766 610 11124
rect 630 10766 634 11124
rect 654 10766 658 11124
rect 678 10766 682 11124
rect 702 10766 706 11124
rect 726 10766 730 11124
rect 750 10766 754 11124
rect 774 10766 778 11124
rect 798 10766 802 11124
rect 822 10766 826 11124
rect 846 10766 850 11124
rect 870 10766 874 11124
rect 894 10766 898 11124
rect 918 10766 922 11124
rect 942 10766 946 11124
rect 955 10997 960 11007
rect 966 10997 970 11124
rect 965 10983 970 10997
rect 955 10973 960 10983
rect 965 10959 970 10973
rect 966 10766 970 10959
rect 990 10931 994 11124
rect 990 10886 997 10931
rect 1014 10886 1018 11124
rect 1038 10886 1042 11124
rect 1062 10886 1066 11124
rect 1086 10886 1090 11124
rect 1110 10886 1114 11124
rect 1134 10886 1138 11124
rect 1158 10886 1162 11124
rect 1182 10886 1186 11124
rect 1206 10886 1210 11124
rect 1230 10886 1234 11124
rect 1254 10886 1258 11124
rect 1278 10886 1282 11124
rect 1302 10886 1306 11124
rect 1326 10886 1330 11124
rect 1350 10886 1354 11124
rect 1374 10886 1378 11124
rect 1398 10886 1402 11124
rect 1422 10886 1426 11124
rect 1446 10886 1450 11124
rect 1470 10886 1474 11124
rect 1494 10886 1498 11124
rect 1501 11123 1515 11124
rect 1518 11099 1525 11147
rect 1518 10886 1522 11099
rect 1542 10886 1546 11196
rect 1566 10886 1570 11196
rect 1590 10886 1594 11196
rect 1614 10886 1618 11196
rect 1638 10886 1642 11196
rect 1662 10886 1666 11196
rect 1686 10886 1690 11196
rect 1710 10886 1714 11196
rect 1734 10886 1738 11196
rect 1758 10886 1762 11196
rect 1782 10886 1786 11196
rect 1806 10886 1810 11196
rect 1830 10886 1834 11196
rect 1854 10886 1858 11196
rect 1878 10886 1882 11196
rect 1902 10886 1906 11196
rect 1926 10886 1930 11196
rect 1950 10886 1954 11196
rect 1974 10886 1978 11196
rect 1998 10886 2002 11196
rect 2022 10886 2026 11196
rect 2046 10886 2050 11196
rect 2070 10886 2074 11196
rect 2094 10886 2098 11196
rect 2118 10886 2122 11196
rect 2142 10886 2146 11196
rect 2166 10886 2170 11196
rect 2190 10886 2194 11196
rect 2214 10886 2218 11196
rect 2227 11117 2232 11127
rect 2238 11117 2242 11196
rect 2237 11103 2242 11117
rect 2227 11102 2261 11103
rect 2262 11102 2266 11196
rect 2286 11102 2290 11196
rect 2310 11102 2314 11196
rect 2334 11102 2338 11196
rect 2358 11102 2362 11196
rect 2382 11102 2386 11196
rect 2406 11102 2410 11196
rect 2430 11102 2434 11196
rect 2454 11102 2458 11196
rect 2478 11102 2482 11196
rect 2502 11102 2506 11196
rect 2526 11102 2530 11196
rect 2550 11102 2554 11196
rect 2574 11102 2578 11196
rect 2598 11102 2602 11196
rect 2622 11102 2626 11196
rect 2646 11102 2650 11196
rect 2670 11102 2674 11196
rect 2694 11102 2698 11196
rect 2718 11102 2722 11196
rect 2742 11102 2746 11196
rect 2766 11102 2770 11196
rect 2790 11102 2794 11196
rect 2814 11102 2818 11196
rect 2838 11102 2842 11196
rect 2862 11102 2866 11196
rect 2886 11102 2890 11196
rect 2910 11102 2914 11196
rect 2934 11102 2938 11196
rect 2958 11102 2962 11196
rect 2982 11102 2986 11196
rect 3006 11102 3010 11196
rect 3030 11102 3034 11196
rect 3054 11102 3058 11196
rect 3078 11102 3082 11196
rect 3102 11102 3106 11196
rect 3115 11189 3120 11196
rect 3126 11189 3130 11196
rect 3133 11195 3147 11196
rect 3125 11175 3130 11189
rect 3115 11165 3120 11175
rect 3125 11151 3130 11165
rect 3126 11103 3130 11151
rect 3115 11102 3147 11103
rect 2227 11100 3147 11102
rect 2227 11093 2232 11100
rect 2237 11079 2242 11093
rect 2238 10886 2242 11079
rect 2262 11051 2266 11100
rect 2262 11003 2269 11051
rect 2262 10886 2266 11003
rect 2286 10886 2290 11100
rect 2310 10886 2314 11100
rect 2334 10886 2338 11100
rect 2358 10886 2362 11100
rect 2382 10886 2386 11100
rect 2406 10886 2410 11100
rect 2430 10886 2434 11100
rect 2454 10886 2458 11100
rect 2478 10886 2482 11100
rect 2502 10886 2506 11100
rect 2526 10886 2530 11100
rect 2550 10886 2554 11100
rect 2574 10886 2578 11100
rect 2598 10886 2602 11100
rect 2622 10886 2626 11100
rect 2646 10886 2650 11100
rect 2670 10886 2674 11100
rect 2694 10886 2698 11100
rect 2718 10886 2722 11100
rect 2742 10886 2746 11100
rect 2766 10886 2770 11100
rect 2790 10886 2794 11100
rect 2814 10886 2818 11100
rect 2838 10886 2842 11100
rect 2862 10886 2866 11100
rect 2886 10886 2890 11100
rect 2910 10886 2914 11100
rect 2934 10886 2938 11100
rect 2958 10886 2962 11100
rect 2982 10886 2986 11100
rect 3006 10886 3010 11100
rect 3030 10886 3034 11100
rect 3054 10886 3058 11100
rect 3078 10886 3082 11100
rect 3102 10886 3106 11100
rect 3115 11093 3120 11100
rect 3126 11093 3130 11100
rect 3133 11099 3147 11100
rect 3125 11079 3130 11093
rect 3139 11089 3147 11093
rect 3133 11079 3139 11089
rect 3115 11045 3120 11055
rect 3125 11031 3130 11045
rect 3115 10973 3120 10983
rect 3126 10973 3130 11031
rect 3125 10959 3130 10973
rect 3139 10969 3147 10973
rect 3133 10959 3139 10969
rect 3115 10925 3120 10935
rect 3125 10911 3130 10925
rect 3126 10887 3130 10911
rect 3115 10886 3147 10887
rect 973 10884 3147 10886
rect 973 10883 987 10884
rect 990 10883 997 10884
rect 990 10766 994 10883
rect 1014 10766 1018 10884
rect 1038 10766 1042 10884
rect 1062 10766 1066 10884
rect 1086 10766 1090 10884
rect 1110 10766 1114 10884
rect 1134 10766 1138 10884
rect 1158 10766 1162 10884
rect 1182 10766 1186 10884
rect 1206 10766 1210 10884
rect 1230 10766 1234 10884
rect 1254 10766 1258 10884
rect 1278 10766 1282 10884
rect 1302 10766 1306 10884
rect 1326 10766 1330 10884
rect 1350 10766 1354 10884
rect 1374 10766 1378 10884
rect 1398 10766 1402 10884
rect 1422 10766 1426 10884
rect 1446 10766 1450 10884
rect 1470 10766 1474 10884
rect 1494 10766 1498 10884
rect 1518 10766 1522 10884
rect 1542 10766 1546 10884
rect 1566 10767 1570 10884
rect 1555 10766 1589 10767
rect -2393 10764 1589 10766
rect -2371 10742 -2366 10764
rect -2348 10742 -2343 10764
rect -2325 10752 -2317 10764
rect -2071 10760 -2062 10764
rect -2013 10762 -1983 10764
rect -2000 10761 -1983 10762
rect -2325 10742 -2320 10752
rect -2309 10742 -2301 10752
rect -2100 10751 -2092 10758
rect -2064 10756 -2062 10759
rect -2061 10751 -2059 10756
rect -2071 10746 -2062 10751
rect -2071 10744 -2026 10746
rect -2066 10742 -2012 10744
rect -2000 10742 -1992 10761
rect -1906 10759 -1904 10764
rect -1846 10760 -1806 10764
rect -1846 10753 -1798 10758
rect -1806 10751 -1798 10753
rect -1671 10752 -1663 10764
rect -1854 10749 -1846 10751
rect -1854 10744 -1806 10749
rect -1864 10742 -1796 10743
rect -1655 10742 -1647 10752
rect -1642 10742 -1637 10764
rect -1619 10742 -1614 10764
rect -1530 10742 -1526 10764
rect -1506 10742 -1502 10764
rect -1482 10742 -1478 10764
rect -1458 10742 -1454 10764
rect -1434 10742 -1430 10764
rect -1410 10742 -1406 10764
rect -1386 10742 -1382 10764
rect -1362 10742 -1358 10764
rect -1338 10742 -1334 10764
rect -1314 10742 -1310 10764
rect -1290 10742 -1286 10764
rect -1266 10742 -1262 10764
rect -1242 10743 -1238 10764
rect -1253 10742 -1219 10743
rect -2393 10740 -1219 10742
rect -2371 10694 -2366 10740
rect -2348 10694 -2343 10740
rect -2325 10736 -2320 10740
rect -2317 10736 -2309 10740
rect -2325 10724 -2317 10736
rect -2066 10735 -2062 10740
rect -2147 10732 -2134 10734
rect -2292 10726 -2071 10732
rect -2325 10694 -2320 10724
rect -2092 10710 -2062 10712
rect -2094 10706 -2062 10710
rect -2000 10694 -1992 10740
rect -1846 10733 -1806 10740
rect -1663 10736 -1655 10740
rect -1846 10726 -1680 10732
rect -1671 10724 -1663 10736
rect -1854 10710 -1806 10712
rect -1854 10706 -1680 10710
rect -1642 10694 -1637 10740
rect -1619 10694 -1614 10740
rect -1530 10694 -1526 10740
rect -1506 10694 -1502 10740
rect -1482 10694 -1478 10740
rect -1458 10694 -1454 10740
rect -1434 10694 -1430 10740
rect -1410 10694 -1406 10740
rect -1386 10694 -1382 10740
rect -1362 10694 -1358 10740
rect -1338 10694 -1334 10740
rect -1314 10694 -1310 10740
rect -1290 10694 -1286 10740
rect -1266 10694 -1262 10740
rect -1253 10733 -1248 10740
rect -1242 10733 -1238 10740
rect -1243 10719 -1238 10733
rect -1253 10709 -1248 10719
rect -1243 10695 -1238 10709
rect -1242 10694 -1238 10695
rect -1218 10694 -1214 10764
rect -1194 10694 -1190 10764
rect -1170 10694 -1166 10764
rect -1146 10694 -1142 10764
rect -1122 10694 -1118 10764
rect -1098 10694 -1094 10764
rect -1074 10694 -1070 10764
rect -1050 10694 -1046 10764
rect -1026 10694 -1022 10764
rect -1002 10694 -998 10764
rect -978 10694 -974 10764
rect -954 10718 -947 10739
rect -930 10718 -926 10764
rect -906 10718 -902 10764
rect -882 10718 -878 10764
rect -858 10763 -854 10764
rect -858 10739 -851 10763
rect -834 10718 -830 10764
rect -810 10718 -806 10764
rect -786 10718 -782 10764
rect -762 10718 -758 10764
rect -738 10718 -734 10764
rect -714 10718 -710 10764
rect -690 10718 -686 10764
rect -666 10718 -662 10764
rect -642 10718 -638 10764
rect -618 10718 -614 10764
rect -594 10718 -590 10764
rect -570 10718 -566 10764
rect -546 10718 -542 10764
rect -522 10718 -518 10764
rect -498 10718 -494 10764
rect -474 10718 -470 10764
rect -450 10718 -446 10764
rect -426 10718 -422 10764
rect -402 10718 -398 10764
rect -378 10718 -374 10764
rect -354 10718 -350 10764
rect -330 10718 -326 10764
rect -306 10718 -302 10764
rect -282 10718 -278 10764
rect -258 10718 -254 10764
rect -234 10718 -230 10764
rect -210 10718 -206 10764
rect -186 10718 -182 10764
rect -162 10718 -158 10764
rect -138 10718 -134 10764
rect -114 10718 -110 10764
rect -90 10718 -86 10764
rect -66 10718 -62 10764
rect -42 10718 -38 10764
rect -18 10718 -14 10764
rect 6 10718 10 10764
rect 30 10718 34 10764
rect 54 10718 58 10764
rect 78 10718 82 10764
rect 102 10718 106 10764
rect 126 10718 130 10764
rect 150 10718 154 10764
rect 174 10718 178 10764
rect 198 10718 202 10764
rect 222 10718 226 10764
rect 246 10718 250 10764
rect 270 10718 274 10764
rect 294 10718 298 10764
rect 318 10718 322 10764
rect 342 10718 346 10764
rect 366 10718 370 10764
rect 390 10718 394 10764
rect 414 10718 418 10764
rect 438 10718 442 10764
rect 462 10718 466 10764
rect 486 10718 490 10764
rect 510 10718 514 10764
rect 534 10718 538 10764
rect 558 10718 562 10764
rect 582 10718 586 10764
rect 606 10718 610 10764
rect 630 10718 634 10764
rect 654 10718 658 10764
rect 678 10718 682 10764
rect 702 10718 706 10764
rect 726 10718 730 10764
rect 750 10718 754 10764
rect 774 10718 778 10764
rect 798 10718 802 10764
rect 822 10718 826 10764
rect 846 10718 850 10764
rect 870 10718 874 10764
rect 894 10718 898 10764
rect 918 10718 922 10764
rect 942 10718 946 10764
rect 966 10718 970 10764
rect 990 10718 994 10764
rect 1014 10718 1018 10764
rect 1038 10718 1042 10764
rect 1062 10718 1066 10764
rect 1086 10718 1090 10764
rect 1110 10718 1114 10764
rect 1134 10718 1138 10764
rect 1158 10718 1162 10764
rect 1182 10718 1186 10764
rect 1206 10718 1210 10764
rect 1230 10718 1234 10764
rect 1254 10718 1258 10764
rect 1278 10718 1282 10764
rect 1302 10718 1306 10764
rect 1326 10718 1330 10764
rect 1350 10718 1354 10764
rect 1374 10718 1378 10764
rect 1398 10718 1402 10764
rect 1422 10718 1426 10764
rect 1446 10718 1450 10764
rect 1470 10718 1474 10764
rect 1494 10718 1498 10764
rect 1518 10718 1522 10764
rect 1542 10718 1546 10764
rect 1555 10757 1560 10764
rect 1566 10757 1570 10764
rect 1565 10743 1570 10757
rect 1555 10733 1560 10743
rect 1565 10719 1570 10733
rect 1566 10718 1570 10719
rect 1590 10718 1594 10884
rect 1614 10718 1618 10884
rect 1638 10718 1642 10884
rect 1662 10718 1666 10884
rect 1686 10718 1690 10884
rect 1710 10718 1714 10884
rect 1734 10718 1738 10884
rect 1758 10718 1762 10884
rect 1782 10718 1786 10884
rect 1806 10718 1810 10884
rect 1830 10718 1834 10884
rect 1854 10718 1858 10884
rect 1878 10718 1882 10884
rect 1902 10718 1906 10884
rect 1926 10718 1930 10884
rect 1950 10718 1954 10884
rect 1974 10718 1978 10884
rect 1998 10718 2002 10884
rect 2022 10718 2026 10884
rect 2046 10718 2050 10884
rect 2070 10718 2074 10884
rect 2094 10718 2098 10884
rect 2118 10718 2122 10884
rect 2142 10718 2146 10884
rect 2166 10718 2170 10884
rect 2190 10718 2194 10884
rect 2214 10718 2218 10884
rect 2238 10718 2242 10884
rect 2262 10718 2266 10884
rect 2286 10718 2290 10884
rect 2310 10718 2314 10884
rect 2334 10718 2338 10884
rect 2358 10718 2362 10884
rect 2382 10718 2386 10884
rect 2406 10718 2410 10884
rect 2430 10718 2434 10884
rect 2443 10853 2448 10863
rect 2454 10853 2458 10884
rect 2453 10839 2458 10853
rect 2443 10838 2477 10839
rect 2478 10838 2482 10884
rect 2502 10838 2506 10884
rect 2526 10838 2530 10884
rect 2550 10838 2554 10884
rect 2574 10838 2578 10884
rect 2598 10838 2602 10884
rect 2622 10838 2626 10884
rect 2646 10838 2650 10884
rect 2670 10838 2674 10884
rect 2694 10838 2698 10884
rect 2718 10838 2722 10884
rect 2742 10838 2746 10884
rect 2766 10838 2770 10884
rect 2790 10838 2794 10884
rect 2814 10838 2818 10884
rect 2838 10838 2842 10884
rect 2862 10838 2866 10884
rect 2886 10838 2890 10884
rect 2910 10838 2914 10884
rect 2934 10838 2938 10884
rect 2958 10838 2962 10884
rect 2982 10838 2986 10884
rect 3006 10838 3010 10884
rect 3030 10838 3034 10884
rect 3054 10838 3058 10884
rect 3078 10838 3082 10884
rect 3102 10839 3106 10884
rect 3115 10877 3120 10884
rect 3126 10877 3130 10884
rect 3133 10883 3147 10884
rect 3125 10863 3130 10877
rect 3091 10838 3125 10839
rect 2443 10836 3125 10838
rect 2443 10829 2448 10836
rect 2453 10815 2458 10829
rect 2454 10718 2458 10815
rect 2478 10787 2482 10836
rect 2478 10742 2485 10787
rect 2502 10742 2506 10836
rect 2526 10742 2530 10836
rect 2550 10742 2554 10836
rect 2574 10742 2578 10836
rect 2598 10742 2602 10836
rect 2622 10742 2626 10836
rect 2646 10742 2650 10836
rect 2670 10742 2674 10836
rect 2694 10742 2698 10836
rect 2718 10742 2722 10836
rect 2742 10742 2746 10836
rect 2766 10742 2770 10836
rect 2790 10742 2794 10836
rect 2814 10742 2818 10836
rect 2838 10742 2842 10836
rect 2862 10742 2866 10836
rect 2886 10742 2890 10836
rect 2910 10742 2914 10836
rect 2934 10742 2938 10836
rect 2958 10742 2962 10836
rect 2982 10742 2986 10836
rect 3006 10742 3010 10836
rect 3030 10742 3034 10836
rect 3054 10743 3058 10836
rect 3067 10805 3072 10815
rect 3078 10805 3082 10836
rect 3091 10829 3096 10836
rect 3102 10829 3106 10836
rect 3101 10815 3106 10829
rect 3077 10791 3082 10805
rect 3043 10742 3077 10743
rect 2461 10740 3077 10742
rect 2461 10739 2475 10740
rect 2478 10739 2485 10740
rect 2478 10718 2482 10739
rect 2502 10718 2506 10740
rect 2526 10718 2530 10740
rect 2550 10718 2554 10740
rect 2574 10718 2578 10740
rect 2598 10718 2602 10740
rect 2622 10718 2626 10740
rect 2646 10718 2650 10740
rect 2670 10718 2674 10740
rect 2694 10718 2698 10740
rect 2718 10718 2722 10740
rect 2742 10718 2746 10740
rect 2766 10718 2770 10740
rect 2790 10718 2794 10740
rect 2814 10718 2818 10740
rect 2838 10718 2842 10740
rect 2862 10718 2866 10740
rect 2886 10718 2890 10740
rect 2910 10718 2914 10740
rect 2934 10718 2938 10740
rect 2958 10718 2962 10740
rect 2982 10718 2986 10740
rect 3006 10718 3010 10740
rect 3030 10719 3034 10740
rect 3043 10733 3048 10740
rect 3054 10733 3058 10740
rect 3053 10719 3058 10733
rect 3019 10718 3053 10719
rect -971 10716 3053 10718
rect -971 10715 -957 10716
rect -954 10715 -947 10716
rect -954 10694 -950 10715
rect -930 10694 -926 10716
rect -906 10694 -902 10716
rect -882 10694 -878 10716
rect -2393 10692 -861 10694
rect -2371 10670 -2366 10692
rect -2348 10670 -2343 10692
rect -2325 10670 -2320 10692
rect -2072 10690 -2036 10691
rect -2072 10684 -2054 10690
rect -2309 10676 -2301 10684
rect -2317 10670 -2309 10676
rect -2092 10675 -2062 10680
rect -2000 10671 -1992 10692
rect -1938 10691 -1906 10692
rect -1920 10690 -1906 10691
rect -1806 10684 -1680 10690
rect -1854 10675 -1806 10680
rect -1655 10676 -1647 10684
rect -1982 10671 -1966 10672
rect -2000 10670 -1966 10671
rect -1846 10670 -1806 10673
rect -1663 10670 -1655 10676
rect -1642 10670 -1637 10692
rect -1619 10670 -1614 10692
rect -1530 10670 -1526 10692
rect -1506 10670 -1502 10692
rect -1482 10670 -1478 10692
rect -1458 10670 -1454 10692
rect -1434 10670 -1430 10692
rect -1410 10670 -1406 10692
rect -1386 10670 -1382 10692
rect -1362 10670 -1358 10692
rect -1338 10670 -1334 10692
rect -1314 10670 -1310 10692
rect -1290 10670 -1286 10692
rect -1266 10670 -1262 10692
rect -1242 10670 -1238 10692
rect -1218 10670 -1214 10692
rect -1194 10670 -1190 10692
rect -1170 10670 -1166 10692
rect -1146 10670 -1142 10692
rect -1122 10670 -1118 10692
rect -1098 10670 -1094 10692
rect -1074 10670 -1070 10692
rect -1050 10670 -1046 10692
rect -1026 10670 -1022 10692
rect -1002 10670 -998 10692
rect -978 10670 -974 10692
rect -954 10670 -950 10692
rect -930 10670 -926 10692
rect -906 10670 -902 10692
rect -882 10670 -878 10692
rect -875 10691 -861 10692
rect -858 10691 -851 10715
rect -858 10671 -854 10691
rect -869 10670 -835 10671
rect -2393 10668 -835 10670
rect -2371 10646 -2366 10668
rect -2348 10646 -2343 10668
rect -2325 10646 -2320 10668
rect -2000 10666 -1966 10668
rect -2309 10648 -2301 10656
rect -2062 10655 -2054 10662
rect -2092 10648 -2084 10655
rect -2062 10648 -2026 10650
rect -2317 10646 -2309 10648
rect -2062 10646 -2012 10648
rect -2000 10646 -1992 10666
rect -1982 10665 -1966 10666
rect -1846 10664 -1806 10668
rect -1846 10657 -1798 10662
rect -1806 10655 -1798 10657
rect -1854 10653 -1846 10655
rect -1854 10648 -1806 10653
rect -1655 10648 -1647 10656
rect -1864 10646 -1796 10647
rect -1663 10646 -1655 10648
rect -1642 10646 -1637 10668
rect -1619 10646 -1614 10668
rect -1530 10646 -1526 10668
rect -1506 10646 -1502 10668
rect -1482 10646 -1478 10668
rect -1458 10646 -1454 10668
rect -1434 10646 -1430 10668
rect -1410 10646 -1406 10668
rect -1386 10646 -1382 10668
rect -1362 10646 -1358 10668
rect -1338 10646 -1334 10668
rect -1314 10646 -1310 10668
rect -1290 10646 -1286 10668
rect -1266 10646 -1262 10668
rect -1242 10646 -1238 10668
rect -1218 10667 -1214 10668
rect -2393 10644 -1221 10646
rect -2371 10598 -2366 10644
rect -2348 10598 -2343 10644
rect -2325 10598 -2320 10644
rect -2317 10640 -2309 10644
rect -2062 10640 -2054 10644
rect -2154 10636 -2138 10638
rect -2057 10636 -2054 10640
rect -2292 10630 -2054 10636
rect -2052 10630 -2044 10640
rect -2092 10614 -2062 10616
rect -2094 10610 -2062 10614
rect -2000 10598 -1992 10644
rect -1846 10637 -1806 10644
rect -1663 10640 -1655 10644
rect -1846 10630 -1680 10636
rect -1854 10614 -1806 10616
rect -1854 10610 -1680 10614
rect -1642 10598 -1637 10644
rect -1619 10598 -1614 10644
rect -1530 10598 -1526 10644
rect -1506 10598 -1502 10644
rect -1482 10598 -1478 10644
rect -1458 10598 -1454 10644
rect -1434 10598 -1430 10644
rect -1410 10598 -1406 10644
rect -1386 10598 -1382 10644
rect -1362 10598 -1358 10644
rect -1338 10598 -1334 10644
rect -1314 10598 -1310 10644
rect -1290 10598 -1286 10644
rect -1266 10598 -1262 10644
rect -1242 10598 -1238 10644
rect -1235 10643 -1221 10644
rect -1218 10619 -1211 10667
rect -1218 10598 -1214 10619
rect -1194 10598 -1190 10668
rect -1170 10598 -1166 10668
rect -1146 10598 -1142 10668
rect -1122 10598 -1118 10668
rect -1098 10598 -1094 10668
rect -1074 10598 -1070 10668
rect -1050 10598 -1046 10668
rect -1026 10598 -1022 10668
rect -1002 10598 -998 10668
rect -978 10598 -974 10668
rect -954 10598 -950 10668
rect -930 10598 -926 10668
rect -906 10598 -902 10668
rect -882 10598 -878 10668
rect -869 10661 -864 10668
rect -858 10661 -854 10668
rect -859 10647 -854 10661
rect -858 10598 -854 10647
rect -834 10598 -830 10716
rect -810 10598 -806 10716
rect -786 10598 -782 10716
rect -762 10598 -758 10716
rect -738 10598 -734 10716
rect -714 10598 -710 10716
rect -690 10598 -686 10716
rect -666 10598 -662 10716
rect -642 10598 -638 10716
rect -618 10598 -614 10716
rect -594 10598 -590 10716
rect -570 10598 -566 10716
rect -546 10598 -542 10716
rect -522 10598 -518 10716
rect -498 10598 -494 10716
rect -474 10598 -470 10716
rect -450 10598 -446 10716
rect -426 10598 -422 10716
rect -402 10598 -398 10716
rect -378 10598 -374 10716
rect -354 10598 -350 10716
rect -330 10598 -326 10716
rect -306 10598 -302 10716
rect -282 10598 -278 10716
rect -258 10598 -254 10716
rect -234 10598 -230 10716
rect -210 10598 -206 10716
rect -186 10598 -182 10716
rect -162 10598 -158 10716
rect -138 10598 -134 10716
rect -114 10598 -110 10716
rect -90 10598 -86 10716
rect -66 10598 -62 10716
rect -42 10598 -38 10716
rect -18 10598 -14 10716
rect 6 10598 10 10716
rect 30 10598 34 10716
rect 54 10598 58 10716
rect 78 10598 82 10716
rect 102 10598 106 10716
rect 126 10598 130 10716
rect 150 10598 154 10716
rect 174 10598 178 10716
rect 198 10598 202 10716
rect 222 10598 226 10716
rect 246 10598 250 10716
rect 270 10598 274 10716
rect 294 10598 298 10716
rect 318 10598 322 10716
rect 342 10598 346 10716
rect 366 10598 370 10716
rect 390 10598 394 10716
rect 414 10598 418 10716
rect 438 10598 442 10716
rect 462 10598 466 10716
rect 486 10598 490 10716
rect 510 10598 514 10716
rect 534 10598 538 10716
rect 558 10598 562 10716
rect 582 10598 586 10716
rect 606 10598 610 10716
rect 630 10598 634 10716
rect 654 10598 658 10716
rect 678 10598 682 10716
rect 702 10598 706 10716
rect 726 10598 730 10716
rect 750 10598 754 10716
rect 774 10598 778 10716
rect 798 10598 802 10716
rect 822 10598 826 10716
rect 846 10598 850 10716
rect 870 10598 874 10716
rect 894 10598 898 10716
rect 918 10598 922 10716
rect 942 10598 946 10716
rect 966 10598 970 10716
rect 979 10637 984 10647
rect 990 10637 994 10716
rect 989 10623 994 10637
rect 990 10598 994 10623
rect 1014 10598 1018 10716
rect 1038 10598 1042 10716
rect 1062 10598 1066 10716
rect 1086 10598 1090 10716
rect 1110 10598 1114 10716
rect 1134 10598 1138 10716
rect 1158 10598 1162 10716
rect 1182 10598 1186 10716
rect 1206 10598 1210 10716
rect 1230 10598 1234 10716
rect 1254 10598 1258 10716
rect 1278 10598 1282 10716
rect 1302 10598 1306 10716
rect 1326 10598 1330 10716
rect 1350 10598 1354 10716
rect 1374 10598 1378 10716
rect 1398 10598 1402 10716
rect 1422 10598 1426 10716
rect 1446 10598 1450 10716
rect 1470 10598 1474 10716
rect 1494 10598 1498 10716
rect 1518 10598 1522 10716
rect 1542 10598 1546 10716
rect 1566 10598 1570 10716
rect 1590 10691 1594 10716
rect 1590 10643 1597 10691
rect 1590 10598 1594 10643
rect 1614 10598 1618 10716
rect 1638 10598 1642 10716
rect 1662 10598 1666 10716
rect 1686 10598 1690 10716
rect 1710 10598 1714 10716
rect 1734 10598 1738 10716
rect 1758 10598 1762 10716
rect 1782 10598 1786 10716
rect 1806 10598 1810 10716
rect 1830 10598 1834 10716
rect 1854 10598 1858 10716
rect 1878 10598 1882 10716
rect 1902 10598 1906 10716
rect 1926 10598 1930 10716
rect 1950 10598 1954 10716
rect 1974 10598 1978 10716
rect 1998 10598 2002 10716
rect 2022 10598 2026 10716
rect 2046 10598 2050 10716
rect 2070 10598 2074 10716
rect 2094 10598 2098 10716
rect 2118 10598 2122 10716
rect 2142 10598 2146 10716
rect 2166 10598 2170 10716
rect 2190 10598 2194 10716
rect 2214 10598 2218 10716
rect 2238 10598 2242 10716
rect 2262 10598 2266 10716
rect 2286 10598 2290 10716
rect 2310 10598 2314 10716
rect 2334 10598 2338 10716
rect 2358 10598 2362 10716
rect 2382 10598 2386 10716
rect 2406 10598 2410 10716
rect 2430 10598 2434 10716
rect 2454 10598 2458 10716
rect 2478 10598 2482 10716
rect 2502 10598 2506 10716
rect 2526 10598 2530 10716
rect 2550 10598 2554 10716
rect 2574 10598 2578 10716
rect 2598 10598 2602 10716
rect 2622 10598 2626 10716
rect 2646 10598 2650 10716
rect 2670 10598 2674 10716
rect 2694 10598 2698 10716
rect 2718 10598 2722 10716
rect 2742 10598 2746 10716
rect 2766 10598 2770 10716
rect 2790 10598 2794 10716
rect 2814 10598 2818 10716
rect 2838 10598 2842 10716
rect 2862 10598 2866 10716
rect 2886 10598 2890 10716
rect 2910 10598 2914 10716
rect 2934 10598 2938 10716
rect 2958 10598 2962 10716
rect 2982 10598 2986 10716
rect 3006 10598 3010 10716
rect 3019 10709 3024 10716
rect 3030 10709 3034 10716
rect 3029 10695 3034 10709
rect 3019 10685 3024 10695
rect 3029 10671 3034 10685
rect 3030 10598 3034 10671
rect 3043 10598 3051 10599
rect -2393 10596 3051 10598
rect -2371 10574 -2366 10596
rect -2348 10574 -2343 10596
rect -2325 10574 -2320 10596
rect -2072 10594 -2036 10595
rect -2072 10588 -2054 10594
rect -2309 10580 -2301 10588
rect -2317 10574 -2309 10580
rect -2092 10579 -2062 10584
rect -2000 10575 -1992 10596
rect -1938 10595 -1906 10596
rect -1920 10594 -1906 10595
rect -1806 10588 -1680 10594
rect -1854 10579 -1806 10584
rect -1655 10580 -1647 10588
rect -1982 10575 -1966 10576
rect -2000 10574 -1966 10575
rect -1846 10574 -1806 10577
rect -1663 10574 -1655 10580
rect -1642 10574 -1637 10596
rect -1619 10574 -1614 10596
rect -1530 10574 -1526 10596
rect -1506 10574 -1502 10596
rect -1482 10574 -1478 10596
rect -1458 10574 -1454 10596
rect -1434 10574 -1430 10596
rect -1410 10575 -1406 10596
rect -1421 10574 -1387 10575
rect -2393 10572 -1387 10574
rect -2371 10550 -2366 10572
rect -2348 10550 -2343 10572
rect -2325 10550 -2320 10572
rect -2000 10570 -1966 10572
rect -2309 10552 -2301 10560
rect -2062 10559 -2054 10566
rect -2092 10552 -2084 10559
rect -2062 10552 -2026 10554
rect -2317 10550 -2309 10552
rect -2062 10550 -2012 10552
rect -2000 10550 -1992 10570
rect -1982 10569 -1966 10570
rect -1846 10568 -1806 10572
rect -1846 10561 -1798 10566
rect -1806 10559 -1798 10561
rect -1854 10557 -1846 10559
rect -1854 10552 -1806 10557
rect -1655 10552 -1647 10560
rect -1864 10550 -1796 10551
rect -1663 10550 -1655 10552
rect -1642 10550 -1637 10572
rect -1619 10550 -1614 10572
rect -1530 10550 -1526 10572
rect -1506 10550 -1502 10572
rect -1482 10550 -1478 10572
rect -1458 10550 -1454 10572
rect -1434 10550 -1430 10572
rect -1421 10565 -1416 10572
rect -1410 10565 -1406 10572
rect -1411 10551 -1406 10565
rect -1421 10550 -1387 10551
rect -1386 10550 -1382 10596
rect -1362 10550 -1358 10596
rect -1338 10550 -1334 10596
rect -1314 10550 -1310 10596
rect -1290 10550 -1286 10596
rect -1266 10550 -1262 10596
rect -1242 10550 -1238 10596
rect -1218 10550 -1214 10596
rect -1194 10550 -1190 10596
rect -1170 10550 -1166 10596
rect -1146 10550 -1142 10596
rect -1122 10550 -1118 10596
rect -1098 10550 -1094 10596
rect -1074 10550 -1070 10596
rect -1050 10550 -1046 10596
rect -1026 10550 -1022 10596
rect -1002 10550 -998 10596
rect -978 10550 -974 10596
rect -954 10550 -950 10596
rect -930 10550 -926 10596
rect -906 10550 -902 10596
rect -882 10550 -878 10596
rect -858 10550 -854 10596
rect -834 10595 -830 10596
rect -834 10571 -827 10595
rect -834 10550 -830 10571
rect -810 10550 -806 10596
rect -786 10550 -782 10596
rect -762 10550 -758 10596
rect -738 10550 -734 10596
rect -714 10550 -710 10596
rect -690 10550 -686 10596
rect -666 10550 -662 10596
rect -642 10550 -638 10596
rect -618 10550 -614 10596
rect -594 10550 -590 10596
rect -570 10550 -566 10596
rect -546 10550 -542 10596
rect -522 10550 -518 10596
rect -498 10550 -494 10596
rect -474 10550 -470 10596
rect -450 10550 -446 10596
rect -426 10550 -422 10596
rect -402 10550 -398 10596
rect -378 10550 -374 10596
rect -354 10550 -350 10596
rect -330 10550 -326 10596
rect -306 10550 -302 10596
rect -282 10550 -278 10596
rect -258 10550 -254 10596
rect -234 10550 -230 10596
rect -210 10550 -206 10596
rect -186 10550 -182 10596
rect -162 10550 -158 10596
rect -138 10550 -134 10596
rect -114 10550 -110 10596
rect -90 10550 -86 10596
rect -66 10550 -62 10596
rect -42 10550 -38 10596
rect -18 10550 -14 10596
rect 6 10550 10 10596
rect 30 10550 34 10596
rect 54 10550 58 10596
rect 78 10550 82 10596
rect 102 10551 106 10596
rect 91 10550 125 10551
rect -2393 10548 125 10550
rect -2371 10502 -2366 10548
rect -2348 10502 -2343 10548
rect -2325 10502 -2320 10548
rect -2317 10544 -2309 10548
rect -2062 10544 -2054 10548
rect -2154 10540 -2138 10542
rect -2057 10540 -2054 10544
rect -2292 10534 -2054 10540
rect -2052 10534 -2044 10544
rect -2092 10518 -2062 10520
rect -2094 10514 -2062 10518
rect -2000 10502 -1992 10548
rect -1846 10541 -1806 10548
rect -1663 10544 -1655 10548
rect -1846 10534 -1680 10540
rect -1854 10518 -1806 10520
rect -1854 10514 -1680 10518
rect -1642 10502 -1637 10548
rect -1619 10502 -1614 10548
rect -1530 10502 -1526 10548
rect -1506 10502 -1502 10548
rect -1482 10502 -1478 10548
rect -1458 10502 -1454 10548
rect -1434 10502 -1430 10548
rect -1421 10541 -1416 10548
rect -1411 10527 -1406 10541
rect -1410 10502 -1406 10527
rect -1386 10502 -1382 10548
rect -1362 10502 -1358 10548
rect -1338 10502 -1334 10548
rect -1314 10502 -1310 10548
rect -1290 10502 -1286 10548
rect -1266 10502 -1262 10548
rect -1242 10502 -1238 10548
rect -1218 10502 -1214 10548
rect -1194 10502 -1190 10548
rect -1170 10502 -1166 10548
rect -1146 10502 -1142 10548
rect -1122 10502 -1118 10548
rect -1098 10502 -1094 10548
rect -1074 10502 -1070 10548
rect -1050 10502 -1046 10548
rect -1026 10502 -1022 10548
rect -1002 10502 -998 10548
rect -978 10502 -974 10548
rect -954 10502 -950 10548
rect -930 10502 -926 10548
rect -906 10502 -902 10548
rect -882 10502 -878 10548
rect -858 10502 -854 10548
rect -834 10502 -830 10548
rect -810 10502 -806 10548
rect -786 10502 -782 10548
rect -762 10502 -758 10548
rect -738 10502 -734 10548
rect -714 10502 -710 10548
rect -690 10502 -686 10548
rect -666 10502 -662 10548
rect -642 10502 -638 10548
rect -618 10502 -614 10548
rect -594 10502 -590 10548
rect -570 10502 -566 10548
rect -546 10502 -542 10548
rect -522 10502 -518 10548
rect -498 10502 -494 10548
rect -474 10502 -470 10548
rect -450 10502 -446 10548
rect -426 10502 -422 10548
rect -402 10502 -398 10548
rect -378 10502 -374 10548
rect -354 10502 -350 10548
rect -330 10502 -326 10548
rect -306 10502 -302 10548
rect -282 10502 -278 10548
rect -258 10502 -254 10548
rect -234 10502 -230 10548
rect -210 10502 -206 10548
rect -186 10502 -182 10548
rect -162 10502 -158 10548
rect -138 10502 -134 10548
rect -114 10502 -110 10548
rect -90 10502 -86 10548
rect -66 10502 -62 10548
rect -42 10502 -38 10548
rect -18 10502 -14 10548
rect 6 10502 10 10548
rect 30 10502 34 10548
rect 54 10502 58 10548
rect 78 10502 82 10548
rect 91 10541 96 10548
rect 102 10541 106 10548
rect 101 10527 106 10541
rect 91 10517 96 10527
rect 101 10503 106 10517
rect 102 10502 106 10503
rect 126 10502 130 10596
rect 150 10502 154 10596
rect 174 10502 178 10596
rect 198 10502 202 10596
rect 222 10502 226 10596
rect 246 10502 250 10596
rect 270 10502 274 10596
rect 294 10502 298 10596
rect 318 10502 322 10596
rect 342 10502 346 10596
rect 366 10502 370 10596
rect 390 10502 394 10596
rect 414 10502 418 10596
rect 438 10502 442 10596
rect 462 10502 466 10596
rect 486 10502 490 10596
rect 510 10502 514 10596
rect 534 10502 538 10596
rect 558 10502 562 10596
rect 582 10502 586 10596
rect 606 10502 610 10596
rect 630 10502 634 10596
rect 654 10502 658 10596
rect 678 10502 682 10596
rect 702 10502 706 10596
rect 726 10502 730 10596
rect 750 10502 754 10596
rect 774 10502 778 10596
rect 798 10502 802 10596
rect 822 10502 826 10596
rect 846 10502 850 10596
rect 870 10502 874 10596
rect 894 10502 898 10596
rect 918 10502 922 10596
rect 942 10502 946 10596
rect 966 10502 970 10596
rect 990 10502 994 10596
rect 1014 10571 1018 10596
rect 1014 10547 1021 10571
rect 1014 10502 1018 10547
rect 1038 10502 1042 10596
rect 1062 10502 1066 10596
rect 1086 10502 1090 10596
rect 1110 10502 1114 10596
rect 1134 10502 1138 10596
rect 1158 10502 1162 10596
rect 1182 10502 1186 10596
rect 1206 10502 1210 10596
rect 1230 10502 1234 10596
rect 1254 10502 1258 10596
rect 1278 10502 1282 10596
rect 1302 10502 1306 10596
rect 1326 10502 1330 10596
rect 1350 10502 1354 10596
rect 1374 10502 1378 10596
rect 1398 10502 1402 10596
rect 1422 10502 1426 10596
rect 1446 10502 1450 10596
rect 1470 10502 1474 10596
rect 1494 10502 1498 10596
rect 1518 10502 1522 10596
rect 1542 10502 1546 10596
rect 1566 10502 1570 10596
rect 1590 10502 1594 10596
rect 1614 10502 1618 10596
rect 1638 10502 1642 10596
rect 1662 10502 1666 10596
rect 1686 10502 1690 10596
rect 1710 10502 1714 10596
rect 1734 10502 1738 10596
rect 1758 10502 1762 10596
rect 1782 10502 1786 10596
rect 1806 10502 1810 10596
rect 1830 10502 1834 10596
rect 1854 10502 1858 10596
rect 1878 10502 1882 10596
rect 1902 10502 1906 10596
rect 1926 10502 1930 10596
rect 1950 10502 1954 10596
rect 1974 10502 1978 10596
rect 1998 10502 2002 10596
rect 2022 10502 2026 10596
rect 2046 10502 2050 10596
rect 2070 10502 2074 10596
rect 2094 10502 2098 10596
rect 2118 10502 2122 10596
rect 2142 10502 2146 10596
rect 2166 10502 2170 10596
rect 2190 10502 2194 10596
rect 2214 10502 2218 10596
rect 2238 10502 2242 10596
rect 2262 10502 2266 10596
rect 2286 10502 2290 10596
rect 2310 10502 2314 10596
rect 2334 10502 2338 10596
rect 2358 10502 2362 10596
rect 2382 10502 2386 10596
rect 2406 10502 2410 10596
rect 2430 10502 2434 10596
rect 2454 10502 2458 10596
rect 2478 10502 2482 10596
rect 2502 10502 2506 10596
rect 2526 10502 2530 10596
rect 2550 10502 2554 10596
rect 2574 10502 2578 10596
rect 2598 10502 2602 10596
rect 2622 10502 2626 10596
rect 2646 10502 2650 10596
rect 2670 10502 2674 10596
rect 2694 10502 2698 10596
rect 2718 10502 2722 10596
rect 2742 10502 2746 10596
rect 2766 10502 2770 10596
rect 2790 10502 2794 10596
rect 2814 10502 2818 10596
rect 2838 10502 2842 10596
rect 2862 10502 2866 10596
rect 2886 10502 2890 10596
rect 2910 10502 2914 10596
rect 2934 10502 2938 10596
rect 2958 10502 2962 10596
rect 2982 10502 2986 10596
rect 3006 10502 3010 10596
rect 3030 10502 3034 10596
rect 3037 10595 3051 10596
rect 3043 10589 3048 10595
rect 3053 10575 3058 10589
rect 3043 10517 3048 10527
rect 3054 10517 3058 10575
rect 3053 10503 3058 10517
rect 3067 10513 3075 10517
rect 3061 10503 3067 10513
rect 3043 10502 3075 10503
rect -2393 10500 3075 10502
rect -2371 10478 -2366 10500
rect -2348 10478 -2343 10500
rect -2325 10478 -2320 10500
rect -2072 10498 -2036 10499
rect -2072 10492 -2054 10498
rect -2309 10484 -2301 10492
rect -2317 10478 -2309 10484
rect -2092 10483 -2062 10488
rect -2000 10479 -1992 10500
rect -1938 10499 -1906 10500
rect -1920 10498 -1906 10499
rect -1806 10492 -1680 10498
rect -1854 10483 -1806 10488
rect -1655 10484 -1647 10492
rect -1982 10479 -1966 10480
rect -2000 10478 -1966 10479
rect -1846 10478 -1806 10481
rect -1663 10478 -1655 10484
rect -1642 10478 -1637 10500
rect -1619 10478 -1614 10500
rect -1530 10478 -1526 10500
rect -1506 10478 -1502 10500
rect -1482 10478 -1478 10500
rect -1458 10478 -1454 10500
rect -1434 10478 -1430 10500
rect -1410 10478 -1406 10500
rect -1386 10499 -1382 10500
rect -2393 10476 -1389 10478
rect -2371 10454 -2366 10476
rect -2348 10454 -2343 10476
rect -2325 10454 -2320 10476
rect -2000 10474 -1966 10476
rect -2309 10456 -2301 10464
rect -2062 10463 -2054 10470
rect -2092 10456 -2084 10463
rect -2062 10456 -2026 10458
rect -2317 10454 -2309 10456
rect -2062 10454 -2012 10456
rect -2000 10454 -1992 10474
rect -1982 10473 -1966 10474
rect -1846 10472 -1806 10476
rect -1846 10465 -1798 10470
rect -1806 10463 -1798 10465
rect -1854 10461 -1846 10463
rect -1854 10456 -1806 10461
rect -1655 10456 -1647 10464
rect -1864 10454 -1796 10455
rect -1663 10454 -1655 10456
rect -1642 10454 -1637 10476
rect -1619 10454 -1614 10476
rect -1530 10454 -1526 10476
rect -1506 10454 -1502 10476
rect -1482 10454 -1478 10476
rect -1458 10455 -1454 10476
rect -1469 10454 -1435 10455
rect -2393 10452 -1435 10454
rect -2371 10406 -2366 10452
rect -2348 10406 -2343 10452
rect -2325 10406 -2320 10452
rect -2317 10448 -2309 10452
rect -2062 10448 -2054 10452
rect -2154 10444 -2138 10446
rect -2057 10444 -2054 10448
rect -2292 10438 -2054 10444
rect -2052 10438 -2044 10448
rect -2092 10422 -2062 10424
rect -2094 10418 -2062 10422
rect -2000 10406 -1992 10452
rect -1846 10445 -1806 10452
rect -1663 10448 -1655 10452
rect -1846 10438 -1680 10444
rect -1854 10422 -1806 10424
rect -1854 10418 -1680 10422
rect -1642 10406 -1637 10452
rect -1619 10406 -1614 10452
rect -1530 10406 -1526 10452
rect -1506 10406 -1502 10452
rect -1482 10406 -1478 10452
rect -1469 10445 -1464 10452
rect -1458 10445 -1454 10452
rect -1459 10431 -1454 10445
rect -1458 10406 -1454 10431
rect -1434 10406 -1430 10476
rect -1410 10406 -1406 10476
rect -1403 10475 -1389 10476
rect -1386 10451 -1379 10499
rect -1386 10406 -1382 10451
rect -1362 10406 -1358 10500
rect -1338 10406 -1334 10500
rect -1314 10406 -1310 10500
rect -1290 10406 -1286 10500
rect -1266 10406 -1262 10500
rect -1242 10406 -1238 10500
rect -1218 10406 -1214 10500
rect -1194 10406 -1190 10500
rect -1170 10406 -1166 10500
rect -1146 10406 -1142 10500
rect -1122 10406 -1118 10500
rect -1098 10406 -1094 10500
rect -1074 10406 -1070 10500
rect -1050 10406 -1046 10500
rect -1026 10406 -1022 10500
rect -1002 10406 -998 10500
rect -978 10406 -974 10500
rect -954 10406 -950 10500
rect -930 10406 -926 10500
rect -906 10406 -902 10500
rect -882 10406 -878 10500
rect -858 10406 -854 10500
rect -834 10406 -830 10500
rect -810 10406 -806 10500
rect -786 10406 -782 10500
rect -762 10406 -758 10500
rect -738 10406 -734 10500
rect -725 10469 -720 10479
rect -714 10469 -710 10500
rect -715 10455 -710 10469
rect -714 10406 -710 10455
rect -690 10406 -686 10500
rect -666 10406 -662 10500
rect -642 10406 -638 10500
rect -618 10406 -614 10500
rect -594 10406 -590 10500
rect -570 10406 -566 10500
rect -546 10406 -542 10500
rect -522 10406 -518 10500
rect -498 10406 -494 10500
rect -474 10406 -470 10500
rect -450 10406 -446 10500
rect -426 10406 -422 10500
rect -402 10406 -398 10500
rect -378 10406 -374 10500
rect -354 10406 -350 10500
rect -330 10406 -326 10500
rect -306 10406 -302 10500
rect -282 10406 -278 10500
rect -258 10406 -254 10500
rect -234 10406 -230 10500
rect -210 10406 -206 10500
rect -186 10406 -182 10500
rect -162 10406 -158 10500
rect -138 10406 -134 10500
rect -114 10406 -110 10500
rect -90 10406 -86 10500
rect -66 10406 -62 10500
rect -42 10406 -38 10500
rect -18 10406 -14 10500
rect 6 10406 10 10500
rect 30 10406 34 10500
rect 54 10406 58 10500
rect 78 10406 82 10500
rect 102 10406 106 10500
rect 126 10475 130 10500
rect 126 10427 133 10475
rect 126 10406 130 10427
rect 150 10406 154 10500
rect 174 10406 178 10500
rect 198 10406 202 10500
rect 222 10406 226 10500
rect 246 10406 250 10500
rect 270 10406 274 10500
rect 294 10406 298 10500
rect 318 10406 322 10500
rect 342 10406 346 10500
rect 366 10406 370 10500
rect 390 10406 394 10500
rect 414 10406 418 10500
rect 438 10406 442 10500
rect 462 10406 466 10500
rect 486 10406 490 10500
rect 510 10406 514 10500
rect 534 10406 538 10500
rect 558 10406 562 10500
rect 582 10406 586 10500
rect 606 10406 610 10500
rect 630 10406 634 10500
rect 654 10406 658 10500
rect 678 10406 682 10500
rect 702 10406 706 10500
rect 726 10406 730 10500
rect 750 10406 754 10500
rect 774 10406 778 10500
rect 798 10406 802 10500
rect 822 10406 826 10500
rect 846 10406 850 10500
rect 870 10406 874 10500
rect 894 10406 898 10500
rect 918 10406 922 10500
rect 942 10406 946 10500
rect 966 10406 970 10500
rect 990 10406 994 10500
rect 1014 10406 1018 10500
rect 1038 10406 1042 10500
rect 1062 10406 1066 10500
rect 1086 10406 1090 10500
rect 1110 10406 1114 10500
rect 1134 10406 1138 10500
rect 1158 10406 1162 10500
rect 1182 10406 1186 10500
rect 1206 10406 1210 10500
rect 1230 10406 1234 10500
rect 1254 10406 1258 10500
rect 1278 10406 1282 10500
rect 1302 10406 1306 10500
rect 1326 10406 1330 10500
rect 1350 10406 1354 10500
rect 1374 10406 1378 10500
rect 1398 10406 1402 10500
rect 1422 10406 1426 10500
rect 1446 10406 1450 10500
rect 1470 10406 1474 10500
rect 1494 10406 1498 10500
rect 1518 10406 1522 10500
rect 1542 10406 1546 10500
rect 1566 10406 1570 10500
rect 1590 10406 1594 10500
rect 1614 10406 1618 10500
rect 1638 10406 1642 10500
rect 1662 10406 1666 10500
rect 1686 10406 1690 10500
rect 1710 10406 1714 10500
rect 1734 10406 1738 10500
rect 1758 10406 1762 10500
rect 1782 10406 1786 10500
rect 1806 10406 1810 10500
rect 1830 10406 1834 10500
rect 1854 10406 1858 10500
rect 1878 10406 1882 10500
rect 1902 10406 1906 10500
rect 1926 10406 1930 10500
rect 1950 10406 1954 10500
rect 1974 10406 1978 10500
rect 1998 10406 2002 10500
rect 2022 10406 2026 10500
rect 2046 10406 2050 10500
rect 2070 10406 2074 10500
rect 2094 10406 2098 10500
rect 2118 10406 2122 10500
rect 2142 10406 2146 10500
rect 2166 10406 2170 10500
rect 2190 10406 2194 10500
rect 2214 10406 2218 10500
rect 2238 10406 2242 10500
rect 2262 10406 2266 10500
rect 2286 10406 2290 10500
rect 2310 10406 2314 10500
rect 2334 10406 2338 10500
rect 2358 10406 2362 10500
rect 2382 10406 2386 10500
rect 2406 10406 2410 10500
rect 2430 10406 2434 10500
rect 2454 10406 2458 10500
rect 2478 10406 2482 10500
rect 2502 10406 2506 10500
rect 2526 10406 2530 10500
rect 2550 10406 2554 10500
rect 2574 10406 2578 10500
rect 2598 10406 2602 10500
rect 2622 10406 2626 10500
rect 2646 10406 2650 10500
rect 2670 10406 2674 10500
rect 2694 10406 2698 10500
rect 2718 10406 2722 10500
rect 2742 10406 2746 10500
rect 2766 10406 2770 10500
rect 2790 10406 2794 10500
rect 2814 10406 2818 10500
rect 2838 10406 2842 10500
rect 2862 10406 2866 10500
rect 2886 10406 2890 10500
rect 2910 10406 2914 10500
rect 2934 10406 2938 10500
rect 2958 10406 2962 10500
rect 2982 10406 2986 10500
rect 3006 10406 3010 10500
rect 3030 10406 3034 10500
rect 3043 10493 3048 10500
rect 3061 10499 3075 10500
rect 3053 10479 3058 10493
rect 3054 10406 3058 10479
rect 3067 10406 3075 10407
rect -2393 10404 3075 10406
rect -2371 10382 -2366 10404
rect -2348 10382 -2343 10404
rect -2325 10382 -2320 10404
rect -2072 10402 -2036 10403
rect -2072 10396 -2054 10402
rect -2309 10388 -2301 10396
rect -2317 10382 -2309 10388
rect -2092 10387 -2062 10392
rect -2000 10383 -1992 10404
rect -1938 10403 -1906 10404
rect -1920 10402 -1906 10403
rect -1806 10396 -1680 10402
rect -1854 10387 -1806 10392
rect -1655 10388 -1647 10396
rect -1982 10383 -1966 10384
rect -2000 10382 -1966 10383
rect -1846 10382 -1806 10385
rect -1663 10382 -1655 10388
rect -1642 10382 -1637 10404
rect -1619 10382 -1614 10404
rect -1530 10382 -1526 10404
rect -1506 10382 -1502 10404
rect -1482 10382 -1478 10404
rect -1458 10382 -1454 10404
rect -1434 10382 -1430 10404
rect -1410 10382 -1406 10404
rect -1386 10382 -1382 10404
rect -1362 10382 -1358 10404
rect -1338 10382 -1334 10404
rect -1314 10382 -1310 10404
rect -1290 10382 -1286 10404
rect -1266 10382 -1262 10404
rect -1242 10382 -1238 10404
rect -1218 10382 -1214 10404
rect -1194 10382 -1190 10404
rect -1170 10382 -1166 10404
rect -1146 10382 -1142 10404
rect -1122 10383 -1118 10404
rect -1133 10382 -1099 10383
rect -2393 10380 -1099 10382
rect -2371 10358 -2366 10380
rect -2348 10358 -2343 10380
rect -2325 10358 -2320 10380
rect -2000 10378 -1966 10380
rect -2309 10360 -2301 10368
rect -2062 10367 -2054 10374
rect -2092 10360 -2084 10367
rect -2062 10360 -2026 10362
rect -2317 10358 -2309 10360
rect -2062 10358 -2012 10360
rect -2000 10358 -1992 10378
rect -1982 10377 -1966 10378
rect -1846 10376 -1806 10380
rect -1846 10369 -1798 10374
rect -1806 10367 -1798 10369
rect -1854 10365 -1846 10367
rect -1854 10360 -1806 10365
rect -1655 10360 -1647 10368
rect -1864 10358 -1796 10359
rect -1663 10358 -1655 10360
rect -1642 10358 -1637 10380
rect -1619 10358 -1614 10380
rect -1530 10358 -1526 10380
rect -1506 10358 -1502 10380
rect -1482 10358 -1478 10380
rect -1458 10358 -1454 10380
rect -1434 10379 -1430 10380
rect -2393 10356 -1437 10358
rect -2371 10310 -2366 10356
rect -2348 10310 -2343 10356
rect -2325 10310 -2320 10356
rect -2317 10352 -2309 10356
rect -2062 10352 -2054 10356
rect -2154 10348 -2138 10350
rect -2057 10348 -2054 10352
rect -2292 10342 -2054 10348
rect -2052 10342 -2044 10352
rect -2092 10326 -2062 10328
rect -2094 10322 -2062 10326
rect -2000 10310 -1992 10356
rect -1846 10349 -1806 10356
rect -1663 10352 -1655 10356
rect -1846 10342 -1680 10348
rect -1854 10326 -1806 10328
rect -1854 10322 -1680 10326
rect -1642 10310 -1637 10356
rect -1619 10310 -1614 10356
rect -1530 10310 -1526 10356
rect -1506 10310 -1502 10356
rect -1482 10310 -1478 10356
rect -1458 10310 -1454 10356
rect -1451 10355 -1437 10356
rect -1434 10355 -1427 10379
rect -1434 10310 -1430 10355
rect -1410 10310 -1406 10380
rect -1386 10310 -1382 10380
rect -1362 10310 -1358 10380
rect -1338 10310 -1334 10380
rect -1314 10310 -1310 10380
rect -1290 10310 -1286 10380
rect -1266 10310 -1262 10380
rect -1242 10310 -1238 10380
rect -1218 10310 -1214 10380
rect -1194 10310 -1190 10380
rect -1170 10310 -1166 10380
rect -1146 10310 -1142 10380
rect -1133 10373 -1128 10380
rect -1122 10373 -1118 10380
rect -1123 10359 -1118 10373
rect -1133 10325 -1128 10335
rect -1123 10311 -1118 10325
rect -1122 10310 -1118 10311
rect -1098 10310 -1094 10404
rect -1074 10310 -1070 10404
rect -1050 10310 -1046 10404
rect -1026 10310 -1022 10404
rect -1002 10310 -998 10404
rect -978 10310 -974 10404
rect -954 10310 -950 10404
rect -930 10310 -926 10404
rect -906 10310 -902 10404
rect -882 10310 -878 10404
rect -858 10310 -854 10404
rect -834 10310 -830 10404
rect -810 10310 -806 10404
rect -786 10310 -782 10404
rect -762 10310 -758 10404
rect -738 10310 -734 10404
rect -725 10349 -720 10359
rect -714 10349 -710 10404
rect -715 10335 -710 10349
rect -690 10403 -686 10404
rect -690 10379 -683 10403
rect -725 10310 -691 10311
rect -2393 10308 -691 10310
rect -2371 10286 -2366 10308
rect -2348 10286 -2343 10308
rect -2325 10286 -2320 10308
rect -2072 10306 -2036 10307
rect -2072 10300 -2054 10306
rect -2309 10292 -2301 10300
rect -2317 10286 -2309 10292
rect -2092 10291 -2062 10296
rect -2000 10287 -1992 10308
rect -1938 10307 -1906 10308
rect -1920 10306 -1906 10307
rect -1806 10300 -1680 10306
rect -1854 10291 -1806 10296
rect -1655 10292 -1647 10300
rect -1982 10287 -1966 10288
rect -2000 10286 -1966 10287
rect -1846 10286 -1806 10289
rect -1663 10286 -1655 10292
rect -1642 10286 -1637 10308
rect -1619 10286 -1614 10308
rect -1530 10286 -1526 10308
rect -1506 10286 -1502 10308
rect -1482 10286 -1478 10308
rect -1458 10286 -1454 10308
rect -1434 10286 -1430 10308
rect -1410 10286 -1406 10308
rect -1386 10286 -1382 10308
rect -1362 10286 -1358 10308
rect -1338 10286 -1334 10308
rect -1314 10286 -1310 10308
rect -1290 10287 -1286 10308
rect -1301 10286 -1267 10287
rect -2393 10284 -1267 10286
rect -2371 10262 -2366 10284
rect -2348 10262 -2343 10284
rect -2325 10262 -2320 10284
rect -2000 10282 -1966 10284
rect -2309 10264 -2301 10272
rect -2062 10271 -2054 10278
rect -2092 10264 -2084 10271
rect -2062 10264 -2026 10266
rect -2317 10262 -2309 10264
rect -2062 10262 -2012 10264
rect -2000 10262 -1992 10282
rect -1982 10281 -1966 10282
rect -1846 10280 -1806 10284
rect -1846 10273 -1798 10278
rect -1806 10271 -1798 10273
rect -1854 10269 -1846 10271
rect -1854 10264 -1806 10269
rect -1655 10264 -1647 10272
rect -1864 10262 -1796 10263
rect -1663 10262 -1655 10264
rect -1642 10262 -1637 10284
rect -1619 10262 -1614 10284
rect -1530 10262 -1526 10284
rect -1506 10262 -1502 10284
rect -1482 10262 -1478 10284
rect -1458 10262 -1454 10284
rect -1434 10262 -1430 10284
rect -1410 10262 -1406 10284
rect -1386 10262 -1382 10284
rect -1362 10262 -1358 10284
rect -1338 10262 -1334 10284
rect -1314 10262 -1310 10284
rect -1301 10277 -1296 10284
rect -1290 10277 -1286 10284
rect -1291 10263 -1286 10277
rect -1266 10262 -1262 10308
rect -1242 10262 -1238 10308
rect -1218 10262 -1214 10308
rect -1194 10262 -1190 10308
rect -1170 10262 -1166 10308
rect -1146 10262 -1142 10308
rect -1122 10262 -1118 10308
rect -1098 10307 -1094 10308
rect -1098 10283 -1091 10307
rect -1074 10262 -1070 10308
rect -1050 10262 -1046 10308
rect -1026 10262 -1022 10308
rect -1002 10262 -998 10308
rect -978 10262 -974 10308
rect -954 10262 -950 10308
rect -930 10262 -926 10308
rect -906 10262 -902 10308
rect -882 10262 -878 10308
rect -858 10262 -854 10308
rect -834 10262 -830 10308
rect -810 10262 -806 10308
rect -786 10262 -782 10308
rect -762 10262 -758 10308
rect -738 10262 -734 10308
rect -725 10301 -720 10308
rect -715 10287 -710 10301
rect -714 10262 -710 10287
rect -690 10283 -686 10379
rect -2393 10260 -693 10262
rect -2371 10214 -2366 10260
rect -2348 10214 -2343 10260
rect -2325 10214 -2320 10260
rect -2317 10256 -2309 10260
rect -2062 10256 -2054 10260
rect -2154 10252 -2138 10254
rect -2057 10252 -2054 10256
rect -2292 10246 -2054 10252
rect -2052 10246 -2044 10256
rect -2092 10230 -2062 10232
rect -2094 10226 -2062 10230
rect -2000 10214 -1992 10260
rect -1846 10253 -1806 10260
rect -1663 10256 -1655 10260
rect -1846 10246 -1680 10252
rect -1854 10230 -1806 10232
rect -1854 10226 -1680 10230
rect -1642 10214 -1637 10260
rect -1619 10214 -1614 10260
rect -1530 10214 -1526 10260
rect -1506 10214 -1502 10260
rect -1482 10214 -1478 10260
rect -1458 10214 -1454 10260
rect -1434 10214 -1430 10260
rect -1410 10214 -1406 10260
rect -1386 10214 -1382 10260
rect -1362 10214 -1358 10260
rect -1338 10214 -1334 10260
rect -1314 10214 -1310 10260
rect -1301 10229 -1296 10239
rect -1291 10215 -1286 10229
rect -1290 10214 -1286 10215
rect -1266 10214 -1262 10260
rect -1242 10214 -1238 10260
rect -1218 10214 -1214 10260
rect -1194 10214 -1190 10260
rect -1170 10214 -1166 10260
rect -1146 10214 -1142 10260
rect -1122 10214 -1118 10260
rect -1098 10238 -1091 10259
rect -1074 10238 -1070 10260
rect -1050 10238 -1046 10260
rect -1026 10238 -1022 10260
rect -1002 10238 -998 10260
rect -978 10238 -974 10260
rect -954 10238 -950 10260
rect -930 10238 -926 10260
rect -906 10238 -902 10260
rect -882 10238 -878 10260
rect -858 10238 -854 10260
rect -834 10238 -830 10260
rect -810 10238 -806 10260
rect -786 10238 -782 10260
rect -762 10238 -758 10260
rect -738 10238 -734 10260
rect -714 10238 -710 10260
rect -707 10259 -693 10260
rect -690 10259 -683 10283
rect -666 10238 -662 10404
rect -642 10238 -638 10404
rect -618 10238 -614 10404
rect -594 10238 -590 10404
rect -570 10238 -566 10404
rect -546 10238 -542 10404
rect -522 10238 -518 10404
rect -498 10238 -494 10404
rect -474 10238 -470 10404
rect -450 10238 -446 10404
rect -426 10238 -422 10404
rect -402 10238 -398 10404
rect -378 10238 -374 10404
rect -354 10238 -350 10404
rect -330 10238 -326 10404
rect -306 10238 -302 10404
rect -282 10238 -278 10404
rect -258 10238 -254 10404
rect -234 10238 -230 10404
rect -210 10238 -206 10404
rect -186 10238 -182 10404
rect -162 10238 -158 10404
rect -138 10238 -134 10404
rect -114 10238 -110 10404
rect -90 10238 -86 10404
rect -66 10238 -62 10404
rect -42 10238 -38 10404
rect -18 10238 -14 10404
rect 6 10238 10 10404
rect 30 10238 34 10404
rect 54 10238 58 10404
rect 78 10238 82 10404
rect 102 10238 106 10404
rect 126 10238 130 10404
rect 150 10238 154 10404
rect 174 10238 178 10404
rect 198 10238 202 10404
rect 222 10238 226 10404
rect 246 10238 250 10404
rect 270 10238 274 10404
rect 294 10238 298 10404
rect 318 10238 322 10404
rect 342 10238 346 10404
rect 366 10238 370 10404
rect 390 10238 394 10404
rect 414 10238 418 10404
rect 427 10253 432 10263
rect 438 10253 442 10404
rect 437 10239 442 10253
rect 462 10238 466 10404
rect 486 10238 490 10404
rect 510 10238 514 10404
rect 534 10238 538 10404
rect 558 10238 562 10404
rect 582 10238 586 10404
rect 606 10238 610 10404
rect 630 10238 634 10404
rect 654 10238 658 10404
rect 678 10238 682 10404
rect 702 10238 706 10404
rect 726 10238 730 10404
rect 750 10238 754 10404
rect 774 10238 778 10404
rect 798 10238 802 10404
rect 822 10238 826 10404
rect 846 10238 850 10404
rect 870 10238 874 10404
rect 894 10238 898 10404
rect 918 10238 922 10404
rect 942 10238 946 10404
rect 966 10238 970 10404
rect 990 10238 994 10404
rect 1014 10238 1018 10404
rect 1038 10238 1042 10404
rect 1062 10238 1066 10404
rect 1086 10238 1090 10404
rect 1110 10238 1114 10404
rect 1134 10238 1138 10404
rect 1158 10238 1162 10404
rect 1182 10238 1186 10404
rect 1206 10238 1210 10404
rect 1230 10238 1234 10404
rect 1254 10238 1258 10404
rect 1278 10238 1282 10404
rect 1302 10238 1306 10404
rect 1326 10238 1330 10404
rect 1350 10238 1354 10404
rect 1374 10238 1378 10404
rect 1398 10238 1402 10404
rect 1422 10238 1426 10404
rect 1446 10238 1450 10404
rect 1470 10238 1474 10404
rect 1494 10238 1498 10404
rect 1518 10238 1522 10404
rect 1542 10238 1546 10404
rect 1566 10238 1570 10404
rect 1590 10238 1594 10404
rect 1614 10238 1618 10404
rect 1638 10238 1642 10404
rect 1662 10238 1666 10404
rect 1686 10238 1690 10404
rect 1710 10238 1714 10404
rect 1734 10238 1738 10404
rect 1758 10238 1762 10404
rect 1782 10238 1786 10404
rect 1806 10238 1810 10404
rect 1830 10238 1834 10404
rect 1854 10238 1858 10404
rect 1878 10238 1882 10404
rect 1902 10238 1906 10404
rect 1926 10238 1930 10404
rect 1950 10238 1954 10404
rect 1974 10238 1978 10404
rect 1998 10238 2002 10404
rect 2022 10238 2026 10404
rect 2046 10238 2050 10404
rect 2070 10238 2074 10404
rect 2094 10238 2098 10404
rect 2118 10238 2122 10404
rect 2142 10238 2146 10404
rect 2166 10238 2170 10404
rect 2190 10238 2194 10404
rect 2214 10238 2218 10404
rect 2238 10238 2242 10404
rect 2262 10238 2266 10404
rect 2286 10238 2290 10404
rect 2310 10238 2314 10404
rect 2334 10238 2338 10404
rect 2358 10238 2362 10404
rect 2382 10238 2386 10404
rect 2406 10238 2410 10404
rect 2430 10238 2434 10404
rect 2454 10238 2458 10404
rect 2478 10238 2482 10404
rect 2502 10238 2506 10404
rect 2526 10238 2530 10404
rect 2550 10238 2554 10404
rect 2574 10238 2578 10404
rect 2598 10238 2602 10404
rect 2622 10238 2626 10404
rect 2646 10238 2650 10404
rect 2670 10238 2674 10404
rect 2694 10238 2698 10404
rect 2718 10238 2722 10404
rect 2742 10238 2746 10404
rect 2766 10238 2770 10404
rect 2790 10238 2794 10404
rect 2814 10238 2818 10404
rect 2838 10238 2842 10404
rect 2862 10238 2866 10404
rect 2886 10238 2890 10404
rect 2910 10238 2914 10404
rect 2934 10238 2938 10404
rect 2958 10238 2962 10404
rect 2982 10238 2986 10404
rect 3006 10238 3010 10404
rect 3030 10238 3034 10404
rect 3054 10239 3058 10404
rect 3061 10403 3075 10404
rect 3067 10397 3072 10403
rect 3077 10383 3082 10397
rect 3067 10325 3072 10335
rect 3078 10325 3082 10383
rect 3077 10311 3082 10325
rect 3091 10321 3099 10325
rect 3085 10311 3091 10321
rect 3043 10238 3077 10239
rect -1115 10236 3077 10238
rect -1115 10235 -1101 10236
rect -1098 10235 -1091 10236
rect -1098 10214 -1094 10235
rect -1074 10214 -1070 10236
rect -1050 10214 -1046 10236
rect -1026 10214 -1022 10236
rect -1002 10214 -998 10236
rect -978 10214 -974 10236
rect -954 10214 -950 10236
rect -930 10214 -926 10236
rect -906 10214 -902 10236
rect -882 10214 -878 10236
rect -858 10214 -854 10236
rect -834 10214 -830 10236
rect -810 10214 -806 10236
rect -786 10214 -782 10236
rect -762 10214 -758 10236
rect -738 10214 -734 10236
rect -714 10214 -710 10236
rect -2393 10212 -693 10214
rect -2371 10190 -2366 10212
rect -2348 10190 -2343 10212
rect -2325 10190 -2320 10212
rect -2072 10210 -2036 10211
rect -2072 10204 -2054 10210
rect -2309 10196 -2301 10204
rect -2317 10190 -2309 10196
rect -2092 10195 -2062 10200
rect -2000 10191 -1992 10212
rect -1938 10211 -1906 10212
rect -1920 10210 -1906 10211
rect -1806 10204 -1680 10210
rect -1854 10195 -1806 10200
rect -1655 10196 -1647 10204
rect -1982 10191 -1966 10192
rect -2000 10190 -1966 10191
rect -1846 10190 -1806 10193
rect -1663 10190 -1655 10196
rect -1642 10190 -1637 10212
rect -1619 10190 -1614 10212
rect -1530 10190 -1526 10212
rect -1506 10190 -1502 10212
rect -1482 10190 -1478 10212
rect -1458 10190 -1454 10212
rect -1434 10190 -1430 10212
rect -1410 10190 -1406 10212
rect -1386 10190 -1382 10212
rect -1362 10190 -1358 10212
rect -1338 10190 -1334 10212
rect -1314 10190 -1310 10212
rect -1290 10190 -1286 10212
rect -1266 10211 -1262 10212
rect -2393 10188 -1269 10190
rect -2371 10166 -2366 10188
rect -2348 10166 -2343 10188
rect -2325 10166 -2320 10188
rect -2000 10186 -1966 10188
rect -2309 10168 -2301 10176
rect -2062 10175 -2054 10182
rect -2092 10168 -2084 10175
rect -2062 10168 -2026 10170
rect -2317 10166 -2309 10168
rect -2062 10166 -2012 10168
rect -2000 10166 -1992 10186
rect -1982 10185 -1966 10186
rect -1846 10184 -1806 10188
rect -1846 10177 -1798 10182
rect -1806 10175 -1798 10177
rect -1854 10173 -1846 10175
rect -1854 10168 -1806 10173
rect -1655 10168 -1647 10176
rect -1864 10166 -1796 10167
rect -1663 10166 -1655 10168
rect -1642 10166 -1637 10188
rect -1619 10166 -1614 10188
rect -1530 10166 -1526 10188
rect -1506 10166 -1502 10188
rect -1482 10167 -1478 10188
rect -1493 10166 -1459 10167
rect -2393 10164 -1459 10166
rect -2371 10118 -2366 10164
rect -2348 10118 -2343 10164
rect -2325 10118 -2320 10164
rect -2317 10160 -2309 10164
rect -2062 10160 -2054 10164
rect -2154 10156 -2138 10158
rect -2057 10156 -2054 10160
rect -2292 10150 -2054 10156
rect -2052 10150 -2044 10160
rect -2092 10134 -2062 10136
rect -2094 10130 -2062 10134
rect -2000 10118 -1992 10164
rect -1846 10157 -1806 10164
rect -1663 10160 -1655 10164
rect -1846 10150 -1680 10156
rect -1854 10134 -1806 10136
rect -1854 10130 -1680 10134
rect -1642 10118 -1637 10164
rect -1619 10118 -1614 10164
rect -1530 10118 -1526 10164
rect -1506 10118 -1502 10164
rect -1493 10157 -1488 10164
rect -1482 10157 -1478 10164
rect -1483 10143 -1478 10157
rect -1482 10118 -1478 10143
rect -1458 10118 -1454 10188
rect -1434 10118 -1430 10188
rect -1410 10118 -1406 10188
rect -1386 10118 -1382 10188
rect -1362 10118 -1358 10188
rect -1338 10118 -1334 10188
rect -1314 10118 -1310 10188
rect -1290 10118 -1286 10188
rect -1283 10187 -1269 10188
rect -1266 10187 -1259 10211
rect -1266 10139 -1259 10163
rect -1266 10118 -1262 10139
rect -1242 10118 -1238 10212
rect -1218 10118 -1214 10212
rect -1194 10118 -1190 10212
rect -1170 10118 -1166 10212
rect -1146 10118 -1142 10212
rect -1122 10118 -1118 10212
rect -1098 10118 -1094 10212
rect -1074 10118 -1070 10212
rect -1050 10118 -1046 10212
rect -1026 10118 -1022 10212
rect -1002 10118 -998 10212
rect -978 10118 -974 10212
rect -954 10118 -950 10212
rect -930 10118 -926 10212
rect -906 10118 -902 10212
rect -882 10118 -878 10212
rect -858 10118 -854 10212
rect -834 10118 -830 10212
rect -810 10118 -806 10212
rect -786 10118 -782 10212
rect -762 10118 -758 10212
rect -738 10118 -734 10212
rect -714 10118 -710 10212
rect -707 10211 -693 10212
rect -690 10211 -683 10235
rect -690 10118 -686 10211
rect -666 10118 -662 10236
rect -642 10118 -638 10236
rect -618 10118 -614 10236
rect -594 10118 -590 10236
rect -570 10118 -566 10236
rect -546 10118 -542 10236
rect -522 10118 -518 10236
rect -498 10118 -494 10236
rect -474 10118 -470 10236
rect -450 10118 -446 10236
rect -426 10118 -422 10236
rect -402 10118 -398 10236
rect -378 10118 -374 10236
rect -354 10118 -350 10236
rect -330 10118 -326 10236
rect -306 10118 -302 10236
rect -282 10118 -278 10236
rect -258 10118 -254 10236
rect -234 10118 -230 10236
rect -210 10118 -206 10236
rect -186 10118 -182 10236
rect -162 10118 -158 10236
rect -138 10118 -134 10236
rect -114 10118 -110 10236
rect -90 10118 -86 10236
rect -66 10118 -62 10236
rect -42 10118 -38 10236
rect -18 10118 -14 10236
rect 6 10118 10 10236
rect 30 10118 34 10236
rect 54 10118 58 10236
rect 78 10118 82 10236
rect 102 10118 106 10236
rect 126 10118 130 10236
rect 150 10118 154 10236
rect 174 10118 178 10236
rect 198 10118 202 10236
rect 222 10118 226 10236
rect 246 10118 250 10236
rect 270 10118 274 10236
rect 294 10118 298 10236
rect 318 10118 322 10236
rect 342 10118 346 10236
rect 366 10118 370 10236
rect 390 10118 394 10236
rect 414 10118 418 10236
rect 427 10205 432 10215
rect 437 10191 442 10205
rect 438 10118 442 10191
rect 462 10187 466 10236
rect 462 10163 469 10187
rect -2393 10116 459 10118
rect -2371 10094 -2366 10116
rect -2348 10094 -2343 10116
rect -2325 10094 -2320 10116
rect -2072 10114 -2036 10115
rect -2072 10108 -2054 10114
rect -2309 10100 -2301 10108
rect -2317 10094 -2309 10100
rect -2092 10099 -2062 10104
rect -2000 10095 -1992 10116
rect -1938 10115 -1906 10116
rect -1920 10114 -1906 10115
rect -1806 10108 -1680 10114
rect -1854 10099 -1806 10104
rect -1655 10100 -1647 10108
rect -1982 10095 -1966 10096
rect -2000 10094 -1966 10095
rect -1846 10094 -1806 10097
rect -1663 10094 -1655 10100
rect -1642 10094 -1637 10116
rect -1619 10094 -1614 10116
rect -1530 10094 -1526 10116
rect -1506 10094 -1502 10116
rect -1482 10094 -1478 10116
rect -1458 10094 -1454 10116
rect -1434 10094 -1430 10116
rect -1410 10094 -1406 10116
rect -1386 10094 -1382 10116
rect -1362 10094 -1358 10116
rect -1338 10094 -1334 10116
rect -1314 10094 -1310 10116
rect -1290 10094 -1286 10116
rect -1266 10094 -1262 10116
rect -1242 10094 -1238 10116
rect -1218 10094 -1214 10116
rect -1194 10094 -1190 10116
rect -1170 10094 -1166 10116
rect -1146 10094 -1142 10116
rect -1122 10094 -1118 10116
rect -1098 10094 -1094 10116
rect -1074 10094 -1070 10116
rect -1050 10095 -1046 10116
rect -1061 10094 -1027 10095
rect -2393 10092 -1027 10094
rect -2371 10070 -2366 10092
rect -2348 10070 -2343 10092
rect -2325 10070 -2320 10092
rect -2000 10090 -1966 10092
rect -2309 10072 -2301 10080
rect -2062 10079 -2054 10086
rect -2092 10072 -2084 10079
rect -2062 10072 -2026 10074
rect -2317 10070 -2309 10072
rect -2062 10070 -2012 10072
rect -2000 10070 -1992 10090
rect -1982 10089 -1966 10090
rect -1846 10088 -1806 10092
rect -1846 10081 -1798 10086
rect -1806 10079 -1798 10081
rect -1854 10077 -1846 10079
rect -1854 10072 -1806 10077
rect -1655 10072 -1647 10080
rect -1864 10070 -1796 10071
rect -1663 10070 -1655 10072
rect -1642 10070 -1637 10092
rect -1619 10070 -1614 10092
rect -1530 10070 -1526 10092
rect -1506 10070 -1502 10092
rect -1482 10070 -1478 10092
rect -1458 10091 -1454 10092
rect -2393 10068 -1461 10070
rect -2371 10022 -2366 10068
rect -2348 10022 -2343 10068
rect -2325 10022 -2320 10068
rect -2317 10064 -2309 10068
rect -2062 10064 -2054 10068
rect -2154 10060 -2138 10062
rect -2057 10060 -2054 10064
rect -2292 10054 -2054 10060
rect -2052 10054 -2044 10064
rect -2092 10038 -2062 10040
rect -2094 10034 -2062 10038
rect -2000 10022 -1992 10068
rect -1846 10061 -1806 10068
rect -1663 10064 -1655 10068
rect -1846 10054 -1680 10060
rect -1854 10038 -1806 10040
rect -1854 10034 -1680 10038
rect -1642 10022 -1637 10068
rect -1619 10022 -1614 10068
rect -1530 10022 -1526 10068
rect -1506 10022 -1502 10068
rect -1482 10022 -1478 10068
rect -1475 10067 -1461 10068
rect -1458 10067 -1451 10091
rect -1458 10022 -1454 10067
rect -1434 10022 -1430 10092
rect -1421 10061 -1416 10071
rect -1410 10061 -1406 10092
rect -1411 10047 -1406 10061
rect -1410 10022 -1406 10047
rect -1386 10022 -1382 10092
rect -1362 10022 -1358 10092
rect -1338 10022 -1334 10092
rect -1314 10022 -1310 10092
rect -1290 10022 -1286 10092
rect -1266 10022 -1262 10092
rect -1242 10022 -1238 10092
rect -1218 10022 -1214 10092
rect -1194 10022 -1190 10092
rect -1170 10022 -1166 10092
rect -1146 10022 -1142 10092
rect -1122 10022 -1118 10092
rect -1098 10022 -1094 10092
rect -1074 10022 -1070 10092
rect -1061 10085 -1056 10092
rect -1050 10085 -1046 10092
rect -1051 10071 -1046 10085
rect -1061 10061 -1056 10071
rect -1051 10047 -1046 10061
rect -1050 10022 -1046 10047
rect -1026 10022 -1022 10116
rect -1002 10022 -998 10116
rect -978 10022 -974 10116
rect -954 10022 -950 10116
rect -930 10022 -926 10116
rect -906 10022 -902 10116
rect -882 10022 -878 10116
rect -858 10022 -854 10116
rect -834 10022 -830 10116
rect -810 10022 -806 10116
rect -786 10022 -782 10116
rect -762 10022 -758 10116
rect -738 10022 -734 10116
rect -714 10022 -710 10116
rect -690 10022 -686 10116
rect -666 10022 -662 10116
rect -642 10022 -638 10116
rect -618 10022 -614 10116
rect -594 10022 -590 10116
rect -570 10022 -566 10116
rect -546 10022 -542 10116
rect -522 10022 -518 10116
rect -498 10022 -494 10116
rect -474 10022 -470 10116
rect -450 10022 -446 10116
rect -426 10022 -422 10116
rect -402 10022 -398 10116
rect -378 10022 -374 10116
rect -354 10022 -350 10116
rect -330 10022 -326 10116
rect -306 10022 -302 10116
rect -282 10022 -278 10116
rect -258 10022 -254 10116
rect -234 10022 -230 10116
rect -210 10022 -206 10116
rect -186 10022 -182 10116
rect -162 10022 -158 10116
rect -138 10022 -134 10116
rect -114 10022 -110 10116
rect -90 10022 -86 10116
rect -66 10022 -62 10116
rect -42 10022 -38 10116
rect -18 10022 -14 10116
rect 6 10022 10 10116
rect 30 10022 34 10116
rect 54 10022 58 10116
rect 78 10022 82 10116
rect 102 10022 106 10116
rect 126 10022 130 10116
rect 150 10022 154 10116
rect 174 10022 178 10116
rect 198 10022 202 10116
rect 222 10022 226 10116
rect 246 10022 250 10116
rect 270 10022 274 10116
rect 294 10022 298 10116
rect 318 10022 322 10116
rect 342 10022 346 10116
rect 366 10022 370 10116
rect 390 10022 394 10116
rect 414 10022 418 10116
rect 438 10022 442 10116
rect 445 10115 459 10116
rect 462 10115 469 10139
rect 462 10022 466 10115
rect 486 10022 490 10236
rect 510 10022 514 10236
rect 534 10022 538 10236
rect 558 10022 562 10236
rect 582 10022 586 10236
rect 606 10022 610 10236
rect 630 10022 634 10236
rect 654 10022 658 10236
rect 678 10022 682 10236
rect 702 10022 706 10236
rect 726 10022 730 10236
rect 750 10022 754 10236
rect 774 10022 778 10236
rect 798 10022 802 10236
rect 822 10022 826 10236
rect 846 10022 850 10236
rect 870 10022 874 10236
rect 894 10022 898 10236
rect 918 10022 922 10236
rect 942 10022 946 10236
rect 966 10022 970 10236
rect 990 10022 994 10236
rect 1014 10022 1018 10236
rect 1038 10022 1042 10236
rect 1062 10022 1066 10236
rect 1086 10022 1090 10236
rect 1110 10022 1114 10236
rect 1123 10181 1128 10191
rect 1134 10181 1138 10236
rect 1133 10167 1138 10181
rect 1134 10022 1138 10167
rect 1158 10115 1162 10236
rect 1158 10091 1165 10115
rect 1158 10022 1162 10091
rect 1182 10022 1186 10236
rect 1206 10022 1210 10236
rect 1230 10022 1234 10236
rect 1254 10022 1258 10236
rect 1278 10022 1282 10236
rect 1302 10022 1306 10236
rect 1326 10022 1330 10236
rect 1350 10022 1354 10236
rect 1374 10022 1378 10236
rect 1398 10022 1402 10236
rect 1422 10022 1426 10236
rect 1446 10022 1450 10236
rect 1470 10022 1474 10236
rect 1494 10022 1498 10236
rect 1518 10022 1522 10236
rect 1542 10022 1546 10236
rect 1566 10022 1570 10236
rect 1590 10022 1594 10236
rect 1614 10022 1618 10236
rect 1638 10022 1642 10236
rect 1662 10022 1666 10236
rect 1686 10022 1690 10236
rect 1710 10022 1714 10236
rect 1734 10022 1738 10236
rect 1758 10022 1762 10236
rect 1782 10022 1786 10236
rect 1806 10022 1810 10236
rect 1830 10022 1834 10236
rect 1854 10022 1858 10236
rect 1878 10022 1882 10236
rect 1902 10022 1906 10236
rect 1926 10022 1930 10236
rect 1950 10022 1954 10236
rect 1974 10022 1978 10236
rect 1998 10022 2002 10236
rect 2022 10022 2026 10236
rect 2046 10022 2050 10236
rect 2070 10022 2074 10236
rect 2094 10022 2098 10236
rect 2118 10022 2122 10236
rect 2142 10022 2146 10236
rect 2166 10022 2170 10236
rect 2190 10022 2194 10236
rect 2214 10022 2218 10236
rect 2238 10022 2242 10236
rect 2262 10022 2266 10236
rect 2286 10022 2290 10236
rect 2310 10022 2314 10236
rect 2334 10022 2338 10236
rect 2358 10022 2362 10236
rect 2382 10022 2386 10236
rect 2406 10022 2410 10236
rect 2430 10022 2434 10236
rect 2454 10022 2458 10236
rect 2478 10022 2482 10236
rect 2502 10022 2506 10236
rect 2526 10022 2530 10236
rect 2550 10022 2554 10236
rect 2574 10022 2578 10236
rect 2598 10022 2602 10236
rect 2622 10022 2626 10236
rect 2646 10022 2650 10236
rect 2670 10022 2674 10236
rect 2694 10022 2698 10236
rect 2718 10022 2722 10236
rect 2742 10022 2746 10236
rect 2766 10022 2770 10236
rect 2790 10022 2794 10236
rect 2814 10022 2818 10236
rect 2838 10022 2842 10236
rect 2862 10022 2866 10236
rect 2886 10022 2890 10236
rect 2910 10022 2914 10236
rect 2934 10022 2938 10236
rect 2958 10022 2962 10236
rect 2982 10022 2986 10236
rect 3006 10022 3010 10236
rect 3030 10022 3034 10236
rect 3043 10229 3048 10236
rect 3054 10229 3058 10236
rect 3053 10215 3058 10229
rect 3043 10109 3048 10119
rect 3053 10095 3058 10109
rect 3043 10061 3048 10071
rect 3054 10061 3058 10095
rect 3053 10047 3058 10061
rect 3043 10022 3075 10023
rect -2393 10020 3075 10022
rect -2371 9998 -2366 10020
rect -2348 9998 -2343 10020
rect -2325 9998 -2320 10020
rect -2072 10018 -2036 10019
rect -2072 10012 -2054 10018
rect -2309 10004 -2301 10012
rect -2317 9998 -2309 10004
rect -2092 10003 -2062 10008
rect -2000 9999 -1992 10020
rect -1938 10019 -1906 10020
rect -1920 10018 -1906 10019
rect -1806 10012 -1680 10018
rect -1854 10003 -1806 10008
rect -1655 10004 -1647 10012
rect -1982 9999 -1966 10000
rect -2000 9998 -1966 9999
rect -1846 9998 -1806 10001
rect -1663 9998 -1655 10004
rect -1642 9998 -1637 10020
rect -1619 9998 -1614 10020
rect -1530 9998 -1526 10020
rect -1506 9998 -1502 10020
rect -1482 9998 -1478 10020
rect -1458 9998 -1454 10020
rect -1434 9998 -1430 10020
rect -1410 9998 -1406 10020
rect -1386 9998 -1382 10020
rect -1362 9998 -1358 10020
rect -1338 9998 -1334 10020
rect -1314 9998 -1310 10020
rect -1290 9998 -1286 10020
rect -1266 9998 -1262 10020
rect -1242 9998 -1238 10020
rect -1218 9998 -1214 10020
rect -1194 9998 -1190 10020
rect -1170 9998 -1166 10020
rect -1146 9998 -1142 10020
rect -1122 9998 -1118 10020
rect -1098 9998 -1094 10020
rect -1074 9998 -1070 10020
rect -1050 9998 -1046 10020
rect -1026 10019 -1022 10020
rect -2393 9996 -1029 9998
rect -2371 9974 -2366 9996
rect -2348 9974 -2343 9996
rect -2325 9974 -2320 9996
rect -2000 9994 -1966 9996
rect -2309 9976 -2301 9984
rect -2062 9983 -2054 9990
rect -2092 9976 -2084 9983
rect -2062 9976 -2026 9978
rect -2317 9974 -2309 9976
rect -2062 9974 -2012 9976
rect -2000 9974 -1992 9994
rect -1982 9993 -1966 9994
rect -1846 9992 -1806 9996
rect -1846 9985 -1798 9990
rect -1806 9983 -1798 9985
rect -1854 9981 -1846 9983
rect -1854 9976 -1806 9981
rect -1655 9976 -1647 9984
rect -1864 9974 -1796 9975
rect -1663 9974 -1655 9976
rect -1642 9974 -1637 9996
rect -1619 9974 -1614 9996
rect -1530 9974 -1526 9996
rect -1506 9974 -1502 9996
rect -1482 9974 -1478 9996
rect -1458 9974 -1454 9996
rect -1434 9974 -1430 9996
rect -1410 9975 -1406 9996
rect -1386 9995 -1382 9996
rect -1421 9974 -1389 9975
rect -2393 9972 -1389 9974
rect -2371 9902 -2366 9972
rect -2348 9902 -2343 9972
rect -2325 9902 -2320 9972
rect -2317 9968 -2309 9972
rect -2062 9968 -2054 9972
rect -2154 9964 -2138 9966
rect -2057 9964 -2054 9968
rect -2292 9958 -2054 9964
rect -2052 9958 -2044 9968
rect -2092 9942 -2062 9944
rect -2094 9938 -2062 9942
rect -2309 9908 -2301 9914
rect -2317 9902 -2309 9908
rect -2000 9902 -1992 9972
rect -1846 9965 -1806 9972
rect -1663 9968 -1655 9972
rect -1846 9958 -1680 9964
rect -1854 9942 -1806 9944
rect -1854 9938 -1680 9942
rect -1655 9908 -1647 9914
rect -1663 9902 -1655 9908
rect -1642 9902 -1637 9972
rect -1619 9902 -1614 9972
rect -1530 9902 -1526 9972
rect -1506 9902 -1502 9972
rect -1482 9902 -1478 9972
rect -1458 9902 -1454 9972
rect -1434 9902 -1430 9972
rect -1421 9965 -1416 9972
rect -1410 9965 -1406 9972
rect -1403 9971 -1389 9972
rect -1386 9971 -1379 9995
rect -1411 9951 -1406 9965
rect -1410 9902 -1406 9951
rect -1386 9902 -1382 9971
rect -1362 9902 -1358 9996
rect -1338 9902 -1334 9996
rect -1314 9902 -1310 9996
rect -1290 9902 -1286 9996
rect -1266 9902 -1262 9996
rect -1242 9902 -1238 9996
rect -1218 9902 -1214 9996
rect -1194 9902 -1190 9996
rect -1170 9902 -1166 9996
rect -1146 9902 -1142 9996
rect -1122 9902 -1118 9996
rect -1098 9902 -1094 9996
rect -1074 9902 -1070 9996
rect -1050 9902 -1046 9996
rect -1043 9995 -1029 9996
rect -1026 9971 -1019 10019
rect -1026 9902 -1022 9971
rect -1002 9902 -998 10020
rect -978 9902 -974 10020
rect -954 9902 -950 10020
rect -930 9902 -926 10020
rect -906 9902 -902 10020
rect -882 9902 -878 10020
rect -858 9902 -854 10020
rect -834 9902 -830 10020
rect -810 9902 -806 10020
rect -786 9902 -782 10020
rect -762 9902 -758 10020
rect -738 9902 -734 10020
rect -714 9902 -710 10020
rect -690 9902 -686 10020
rect -666 9902 -662 10020
rect -642 9902 -638 10020
rect -618 9902 -614 10020
rect -594 9902 -590 10020
rect -570 9902 -566 10020
rect -546 9902 -542 10020
rect -522 9902 -518 10020
rect -498 9902 -494 10020
rect -474 9902 -470 10020
rect -450 9902 -446 10020
rect -426 9902 -422 10020
rect -402 9902 -398 10020
rect -378 9902 -374 10020
rect -354 9902 -350 10020
rect -330 9902 -326 10020
rect -306 9902 -302 10020
rect -282 9902 -278 10020
rect -258 9902 -254 10020
rect -234 9902 -230 10020
rect -210 9902 -206 10020
rect -186 9902 -182 10020
rect -162 9902 -158 10020
rect -138 9902 -134 10020
rect -114 9902 -110 10020
rect -90 9902 -86 10020
rect -66 9902 -62 10020
rect -42 9902 -38 10020
rect -18 9902 -14 10020
rect 6 9902 10 10020
rect 30 9902 34 10020
rect 54 9902 58 10020
rect 78 9902 82 10020
rect 102 9902 106 10020
rect 126 9902 130 10020
rect 150 9902 154 10020
rect 174 9902 178 10020
rect 198 9902 202 10020
rect 222 9902 226 10020
rect 246 9902 250 10020
rect 270 9902 274 10020
rect 294 9902 298 10020
rect 318 9902 322 10020
rect 342 9902 346 10020
rect 366 9902 370 10020
rect 390 9902 394 10020
rect 414 9902 418 10020
rect 438 9902 442 10020
rect 462 9902 466 10020
rect 486 9902 490 10020
rect 510 9902 514 10020
rect 534 9902 538 10020
rect 558 9902 562 10020
rect 582 9902 586 10020
rect 606 9902 610 10020
rect 630 9902 634 10020
rect 654 9902 658 10020
rect 678 9902 682 10020
rect 702 9902 706 10020
rect 726 9902 730 10020
rect 750 9902 754 10020
rect 774 9902 778 10020
rect 798 9902 802 10020
rect 822 9902 826 10020
rect 846 9902 850 10020
rect 870 9902 874 10020
rect 894 9902 898 10020
rect 918 9902 922 10020
rect 942 9902 946 10020
rect 966 9902 970 10020
rect 990 9902 994 10020
rect 1014 9902 1018 10020
rect 1038 9902 1042 10020
rect 1062 9902 1066 10020
rect 1086 9902 1090 10020
rect 1110 9902 1114 10020
rect 1134 9902 1138 10020
rect 1158 9902 1162 10020
rect 1182 9902 1186 10020
rect 1206 9902 1210 10020
rect 1230 9902 1234 10020
rect 1254 9902 1258 10020
rect 1278 9902 1282 10020
rect 1302 9902 1306 10020
rect 1326 9902 1330 10020
rect 1350 9902 1354 10020
rect 1374 9902 1378 10020
rect 1398 9902 1402 10020
rect 1422 9902 1426 10020
rect 1446 9902 1450 10020
rect 1470 9902 1474 10020
rect 1494 9902 1498 10020
rect 1507 9989 1512 9999
rect 1518 9989 1522 10020
rect 1517 9975 1522 9989
rect 1507 9974 1541 9975
rect 1542 9974 1546 10020
rect 1566 9974 1570 10020
rect 1590 9974 1594 10020
rect 1614 9974 1618 10020
rect 1638 9974 1642 10020
rect 1662 9974 1666 10020
rect 1686 9974 1690 10020
rect 1710 9974 1714 10020
rect 1734 9974 1738 10020
rect 1758 9974 1762 10020
rect 1782 9974 1786 10020
rect 1806 9974 1810 10020
rect 1830 9974 1834 10020
rect 1854 9974 1858 10020
rect 1878 9974 1882 10020
rect 1902 9974 1906 10020
rect 1926 9974 1930 10020
rect 1950 9974 1954 10020
rect 1974 9974 1978 10020
rect 1998 9974 2002 10020
rect 2022 9974 2026 10020
rect 2046 9974 2050 10020
rect 2070 9974 2074 10020
rect 2094 9974 2098 10020
rect 2118 9974 2122 10020
rect 2142 9974 2146 10020
rect 2166 9974 2170 10020
rect 2190 9974 2194 10020
rect 2214 9974 2218 10020
rect 2238 9974 2242 10020
rect 2262 9974 2266 10020
rect 2286 9974 2290 10020
rect 2310 9974 2314 10020
rect 2334 9974 2338 10020
rect 2358 9974 2362 10020
rect 2382 9974 2386 10020
rect 2406 9974 2410 10020
rect 2430 9974 2434 10020
rect 2454 9974 2458 10020
rect 2478 9974 2482 10020
rect 2502 9974 2506 10020
rect 2526 9974 2530 10020
rect 2550 9974 2554 10020
rect 2574 9974 2578 10020
rect 2598 9974 2602 10020
rect 2622 9974 2626 10020
rect 2646 9974 2650 10020
rect 2670 9974 2674 10020
rect 2694 9974 2698 10020
rect 2718 9974 2722 10020
rect 2742 9974 2746 10020
rect 2766 9974 2770 10020
rect 2790 9974 2794 10020
rect 2814 9974 2818 10020
rect 2838 9974 2842 10020
rect 2862 9974 2866 10020
rect 2886 9974 2890 10020
rect 2910 9974 2914 10020
rect 2934 9974 2938 10020
rect 2958 9974 2962 10020
rect 2982 9974 2986 10020
rect 3006 9974 3010 10020
rect 3030 9974 3034 10020
rect 3043 10013 3048 10020
rect 3061 10019 3075 10020
rect 3053 9999 3058 10013
rect 3054 9975 3058 9999
rect 3043 9974 3075 9975
rect 1507 9972 3075 9974
rect 1507 9965 1512 9972
rect 1517 9951 1522 9965
rect 1518 9902 1522 9951
rect 1542 9923 1546 9972
rect -2393 9900 1539 9902
rect -2371 9806 -2366 9900
rect -2348 9806 -2343 9900
rect -2325 9838 -2320 9900
rect -2317 9898 -2309 9900
rect -2000 9899 -1966 9900
rect -2000 9898 -1982 9899
rect -1663 9898 -1655 9900
rect -2028 9890 -2018 9892
rect -2309 9880 -2301 9886
rect -2091 9880 -2061 9887
rect -2317 9870 -2309 9880
rect -2044 9878 -2028 9880
rect -2026 9878 -2014 9890
rect -2084 9872 -2061 9878
rect -2044 9876 -2014 9878
rect -2292 9862 -2054 9871
rect -2325 9830 -2317 9838
rect -2325 9810 -2320 9830
rect -2317 9822 -2309 9830
rect -2325 9806 -2317 9810
rect -2000 9806 -1992 9898
rect -1982 9897 -1966 9898
rect -1980 9880 -1932 9887
rect -1655 9880 -1647 9886
rect -1846 9862 -1680 9871
rect -1663 9870 -1655 9880
rect -1671 9830 -1663 9838
rect -1663 9822 -1655 9830
rect -1926 9806 -1892 9809
rect -1671 9806 -1663 9810
rect -1642 9806 -1637 9900
rect -1619 9806 -1614 9900
rect -1530 9806 -1526 9900
rect -1506 9806 -1502 9900
rect -1482 9806 -1478 9900
rect -1458 9806 -1454 9900
rect -1434 9806 -1430 9900
rect -1410 9806 -1406 9900
rect -1386 9899 -1382 9900
rect -1386 9875 -1379 9899
rect -1386 9806 -1382 9875
rect -1362 9806 -1358 9900
rect -1338 9806 -1334 9900
rect -1314 9806 -1310 9900
rect -1290 9806 -1286 9900
rect -1266 9806 -1262 9900
rect -1242 9806 -1238 9900
rect -1218 9806 -1214 9900
rect -1194 9806 -1190 9900
rect -1170 9806 -1166 9900
rect -1146 9806 -1142 9900
rect -1122 9806 -1118 9900
rect -1098 9806 -1094 9900
rect -1074 9806 -1070 9900
rect -1050 9806 -1046 9900
rect -1026 9806 -1022 9900
rect -1002 9806 -998 9900
rect -978 9806 -974 9900
rect -954 9806 -950 9900
rect -930 9806 -926 9900
rect -906 9806 -902 9900
rect -882 9806 -878 9900
rect -858 9806 -854 9900
rect -834 9806 -830 9900
rect -810 9806 -806 9900
rect -786 9806 -782 9900
rect -762 9806 -758 9900
rect -738 9806 -734 9900
rect -714 9806 -710 9900
rect -690 9806 -686 9900
rect -666 9806 -662 9900
rect -642 9806 -638 9900
rect -618 9806 -614 9900
rect -594 9806 -590 9900
rect -570 9806 -566 9900
rect -546 9806 -542 9900
rect -522 9806 -518 9900
rect -498 9806 -494 9900
rect -474 9806 -470 9900
rect -450 9806 -446 9900
rect -426 9806 -422 9900
rect -402 9806 -398 9900
rect -378 9806 -374 9900
rect -354 9806 -350 9900
rect -330 9806 -326 9900
rect -306 9806 -302 9900
rect -282 9806 -278 9900
rect -258 9806 -254 9900
rect -234 9806 -230 9900
rect -210 9806 -206 9900
rect -186 9806 -182 9900
rect -162 9806 -158 9900
rect -138 9806 -134 9900
rect -114 9806 -110 9900
rect -90 9806 -86 9900
rect -66 9806 -62 9900
rect -42 9806 -38 9900
rect -18 9806 -14 9900
rect 6 9806 10 9900
rect 30 9806 34 9900
rect 54 9806 58 9900
rect 78 9806 82 9900
rect 102 9806 106 9900
rect 126 9806 130 9900
rect 150 9806 154 9900
rect 174 9806 178 9900
rect 198 9806 202 9900
rect 222 9806 226 9900
rect 246 9806 250 9900
rect 270 9806 274 9900
rect 294 9806 298 9900
rect 318 9806 322 9900
rect 342 9806 346 9900
rect 366 9806 370 9900
rect 390 9806 394 9900
rect 414 9806 418 9900
rect 438 9806 442 9900
rect 462 9806 466 9900
rect 486 9806 490 9900
rect 510 9806 514 9900
rect 534 9806 538 9900
rect 558 9806 562 9900
rect 582 9806 586 9900
rect 606 9806 610 9900
rect 630 9806 634 9900
rect 654 9806 658 9900
rect 678 9806 682 9900
rect 702 9806 706 9900
rect 726 9806 730 9900
rect 750 9806 754 9900
rect 774 9806 778 9900
rect 798 9806 802 9900
rect 822 9806 826 9900
rect 846 9806 850 9900
rect 870 9806 874 9900
rect 894 9806 898 9900
rect 918 9806 922 9900
rect 942 9806 946 9900
rect 966 9806 970 9900
rect 990 9806 994 9900
rect 1014 9806 1018 9900
rect 1038 9806 1042 9900
rect 1062 9806 1066 9900
rect 1086 9806 1090 9900
rect 1110 9806 1114 9900
rect 1134 9806 1138 9900
rect 1158 9806 1162 9900
rect 1182 9806 1186 9900
rect 1206 9806 1210 9900
rect 1230 9806 1234 9900
rect 1254 9806 1258 9900
rect 1278 9806 1282 9900
rect 1302 9806 1306 9900
rect 1326 9806 1330 9900
rect 1350 9806 1354 9900
rect 1374 9806 1378 9900
rect 1398 9806 1402 9900
rect 1422 9806 1426 9900
rect 1446 9806 1450 9900
rect 1470 9806 1474 9900
rect 1494 9806 1498 9900
rect 1518 9806 1522 9900
rect 1525 9899 1539 9900
rect 1542 9875 1549 9923
rect 1542 9806 1546 9875
rect 1566 9806 1570 9972
rect 1590 9806 1594 9972
rect 1614 9806 1618 9972
rect 1638 9806 1642 9972
rect 1662 9806 1666 9972
rect 1686 9806 1690 9972
rect 1710 9806 1714 9972
rect 1734 9806 1738 9972
rect 1758 9806 1762 9972
rect 1782 9806 1786 9972
rect 1806 9806 1810 9972
rect 1830 9806 1834 9972
rect 1843 9845 1848 9855
rect 1854 9845 1858 9972
rect 1853 9831 1858 9845
rect 1843 9821 1848 9831
rect 1853 9807 1858 9821
rect 1854 9806 1858 9807
rect 1878 9806 1882 9972
rect 1902 9806 1906 9972
rect 1926 9806 1930 9972
rect 1950 9806 1954 9972
rect 1974 9806 1978 9972
rect 1998 9806 2002 9972
rect 2022 9806 2026 9972
rect 2046 9806 2050 9972
rect 2070 9806 2074 9972
rect 2094 9806 2098 9972
rect 2118 9806 2122 9972
rect 2142 9806 2146 9972
rect 2166 9806 2170 9972
rect 2190 9806 2194 9972
rect 2214 9806 2218 9972
rect 2238 9806 2242 9972
rect 2262 9806 2266 9972
rect 2286 9806 2290 9972
rect 2310 9806 2314 9972
rect 2334 9806 2338 9972
rect 2358 9806 2362 9972
rect 2382 9806 2386 9972
rect 2406 9806 2410 9972
rect 2430 9806 2434 9972
rect 2454 9806 2458 9972
rect 2478 9806 2482 9972
rect 2502 9806 2506 9972
rect 2526 9806 2530 9972
rect 2550 9806 2554 9972
rect 2574 9806 2578 9972
rect 2598 9806 2602 9972
rect 2622 9806 2626 9972
rect 2646 9806 2650 9972
rect 2670 9806 2674 9972
rect 2694 9806 2698 9972
rect 2718 9806 2722 9972
rect 2742 9806 2746 9972
rect 2766 9806 2770 9972
rect 2790 9806 2794 9972
rect 2814 9806 2818 9972
rect 2838 9806 2842 9972
rect 2862 9806 2866 9972
rect 2886 9806 2890 9972
rect 2910 9806 2914 9972
rect 2934 9806 2938 9972
rect 2958 9806 2962 9972
rect 2982 9806 2986 9972
rect 3006 9806 3010 9972
rect 3030 9806 3034 9972
rect 3043 9965 3048 9972
rect 3054 9965 3058 9972
rect 3061 9971 3075 9972
rect 3053 9951 3058 9965
rect 3043 9893 3048 9903
rect 3053 9879 3058 9893
rect 3067 9889 3075 9893
rect 3061 9879 3067 9889
rect 3043 9821 3048 9831
rect 3054 9821 3058 9879
rect 3053 9807 3058 9821
rect 3067 9817 3075 9821
rect 3061 9807 3067 9817
rect 3043 9806 3075 9807
rect -2393 9804 3075 9806
rect -2371 9758 -2366 9804
rect -2348 9758 -2343 9804
rect -2325 9798 -2317 9804
rect -2053 9802 -1972 9804
rect -2325 9782 -2320 9798
rect -2317 9794 -2309 9798
rect -2069 9794 -2068 9795
rect -2309 9782 -2301 9794
rect -2069 9787 -2038 9794
rect -2069 9785 -2068 9787
rect -2000 9786 -1992 9802
rect -1926 9799 -1924 9804
rect -1916 9796 -1914 9799
rect -1671 9798 -1663 9804
rect -1982 9786 -1916 9795
rect -1663 9794 -1655 9798
rect -2325 9770 -2317 9782
rect -2068 9779 -2053 9785
rect -2027 9784 -1992 9786
rect -2076 9770 -2053 9777
rect -2011 9776 -2002 9784
rect -2000 9776 -1992 9784
rect -1655 9782 -1647 9794
rect -2003 9774 -1992 9776
rect -2325 9758 -2320 9770
rect -2317 9766 -2309 9770
rect -2309 9758 -2301 9766
rect -2015 9762 -2003 9774
rect -2000 9758 -1992 9774
rect -1972 9770 -1924 9777
rect -1862 9769 -1680 9778
rect -1671 9770 -1663 9782
rect -1663 9766 -1655 9770
rect -1976 9758 -1940 9759
rect -1655 9758 -1647 9766
rect -1642 9758 -1637 9804
rect -1619 9758 -1614 9804
rect -1589 9758 -1531 9759
rect -1530 9758 -1526 9804
rect -1506 9758 -1502 9804
rect -1482 9758 -1478 9804
rect -1458 9758 -1454 9804
rect -1434 9758 -1430 9804
rect -1410 9758 -1406 9804
rect -1386 9758 -1382 9804
rect -1362 9758 -1358 9804
rect -1338 9758 -1334 9804
rect -1314 9758 -1310 9804
rect -1290 9758 -1286 9804
rect -1266 9758 -1262 9804
rect -1242 9758 -1238 9804
rect -1218 9758 -1214 9804
rect -1194 9758 -1190 9804
rect -1170 9758 -1166 9804
rect -1146 9758 -1142 9804
rect -1122 9758 -1118 9804
rect -1098 9758 -1094 9804
rect -1074 9758 -1070 9804
rect -1050 9758 -1046 9804
rect -1026 9758 -1022 9804
rect -1002 9758 -998 9804
rect -978 9758 -974 9804
rect -954 9758 -950 9804
rect -930 9758 -926 9804
rect -906 9758 -902 9804
rect -882 9758 -878 9804
rect -858 9758 -854 9804
rect -834 9758 -830 9804
rect -810 9758 -806 9804
rect -786 9758 -782 9804
rect -762 9758 -758 9804
rect -738 9758 -734 9804
rect -714 9758 -710 9804
rect -690 9758 -686 9804
rect -666 9758 -662 9804
rect -642 9759 -638 9804
rect -653 9758 -619 9759
rect -2393 9756 -619 9758
rect -2371 9686 -2366 9756
rect -2348 9686 -2343 9756
rect -2325 9754 -2320 9756
rect -2309 9754 -2301 9756
rect -2325 9742 -2317 9754
rect -2325 9722 -2320 9742
rect -2317 9738 -2309 9742
rect -2325 9714 -2317 9722
rect -2060 9716 -2030 9719
rect -2325 9686 -2320 9714
rect -2317 9706 -2309 9714
rect -2060 9703 -2038 9714
rect -2033 9707 -2030 9716
rect -2028 9712 -2027 9716
rect -2068 9698 -2038 9701
rect -2000 9686 -1992 9756
rect -1655 9754 -1647 9756
rect -1671 9742 -1663 9754
rect -1663 9738 -1655 9742
rect -1912 9731 -1884 9733
rect -1852 9725 -1804 9729
rect -1844 9716 -1796 9719
rect -1671 9714 -1663 9722
rect -1844 9703 -1804 9714
rect -1663 9706 -1655 9714
rect -1852 9698 -1680 9702
rect -1642 9686 -1637 9756
rect -1619 9686 -1614 9756
rect -1565 9710 -1531 9711
rect -1530 9710 -1526 9756
rect -1506 9710 -1502 9756
rect -1482 9710 -1478 9756
rect -1458 9710 -1454 9756
rect -1434 9710 -1430 9756
rect -1410 9710 -1406 9756
rect -1386 9710 -1382 9756
rect -1362 9710 -1358 9756
rect -1338 9710 -1334 9756
rect -1314 9710 -1310 9756
rect -1290 9710 -1286 9756
rect -1266 9710 -1262 9756
rect -1242 9710 -1238 9756
rect -1218 9710 -1214 9756
rect -1194 9710 -1190 9756
rect -1170 9710 -1166 9756
rect -1146 9710 -1142 9756
rect -1122 9710 -1118 9756
rect -1098 9710 -1094 9756
rect -1074 9710 -1070 9756
rect -1050 9710 -1046 9756
rect -1026 9710 -1022 9756
rect -1002 9710 -998 9756
rect -978 9710 -974 9756
rect -954 9710 -950 9756
rect -930 9710 -926 9756
rect -906 9710 -902 9756
rect -882 9710 -878 9756
rect -858 9710 -854 9756
rect -834 9710 -830 9756
rect -810 9710 -806 9756
rect -786 9710 -782 9756
rect -762 9710 -758 9756
rect -738 9710 -734 9756
rect -714 9710 -710 9756
rect -690 9710 -686 9756
rect -666 9710 -662 9756
rect -653 9749 -648 9756
rect -642 9749 -638 9756
rect -643 9735 -638 9749
rect -618 9710 -614 9804
rect -594 9710 -590 9804
rect -570 9710 -566 9804
rect -546 9710 -542 9804
rect -522 9710 -518 9804
rect -498 9710 -494 9804
rect -474 9710 -470 9804
rect -450 9710 -446 9804
rect -426 9710 -422 9804
rect -402 9710 -398 9804
rect -378 9710 -374 9804
rect -354 9710 -350 9804
rect -330 9710 -326 9804
rect -306 9710 -302 9804
rect -282 9710 -278 9804
rect -258 9710 -254 9804
rect -234 9710 -230 9804
rect -210 9710 -206 9804
rect -186 9710 -182 9804
rect -162 9710 -158 9804
rect -138 9710 -134 9804
rect -114 9710 -110 9804
rect -90 9710 -86 9804
rect -66 9710 -62 9804
rect -42 9710 -38 9804
rect -18 9710 -14 9804
rect 6 9710 10 9804
rect 30 9710 34 9804
rect 54 9710 58 9804
rect 78 9710 82 9804
rect 102 9710 106 9804
rect 126 9710 130 9804
rect 150 9710 154 9804
rect 174 9710 178 9804
rect 198 9710 202 9804
rect 222 9710 226 9804
rect 246 9710 250 9804
rect 270 9710 274 9804
rect 294 9710 298 9804
rect 318 9710 322 9804
rect 342 9710 346 9804
rect 366 9710 370 9804
rect 390 9710 394 9804
rect 414 9710 418 9804
rect 438 9710 442 9804
rect 462 9710 466 9804
rect 486 9710 490 9804
rect 510 9710 514 9804
rect 534 9710 538 9804
rect 558 9710 562 9804
rect 582 9710 586 9804
rect 606 9710 610 9804
rect 630 9710 634 9804
rect 654 9710 658 9804
rect 678 9710 682 9804
rect 702 9710 706 9804
rect 726 9710 730 9804
rect 750 9710 754 9804
rect 774 9710 778 9804
rect 798 9710 802 9804
rect 822 9710 826 9804
rect 846 9710 850 9804
rect 870 9710 874 9804
rect 894 9710 898 9804
rect 918 9710 922 9804
rect 942 9710 946 9804
rect 966 9710 970 9804
rect 990 9710 994 9804
rect 1014 9710 1018 9804
rect 1038 9710 1042 9804
rect 1062 9710 1066 9804
rect 1086 9710 1090 9804
rect 1110 9710 1114 9804
rect 1134 9710 1138 9804
rect 1158 9710 1162 9804
rect 1182 9710 1186 9804
rect 1206 9710 1210 9804
rect 1230 9710 1234 9804
rect 1254 9710 1258 9804
rect 1278 9710 1282 9804
rect 1302 9710 1306 9804
rect 1326 9710 1330 9804
rect 1350 9710 1354 9804
rect 1374 9710 1378 9804
rect 1398 9710 1402 9804
rect 1422 9710 1426 9804
rect 1446 9710 1450 9804
rect 1470 9710 1474 9804
rect 1494 9710 1498 9804
rect 1518 9710 1522 9804
rect 1542 9710 1546 9804
rect 1566 9710 1570 9804
rect 1590 9710 1594 9804
rect 1614 9710 1618 9804
rect 1638 9710 1642 9804
rect 1662 9710 1666 9804
rect 1686 9710 1690 9804
rect 1710 9710 1714 9804
rect 1734 9710 1738 9804
rect 1758 9710 1762 9804
rect 1782 9710 1786 9804
rect 1806 9710 1810 9804
rect 1830 9710 1834 9804
rect 1854 9710 1858 9804
rect 1878 9779 1882 9804
rect 1878 9734 1885 9779
rect 1902 9734 1906 9804
rect 1926 9734 1930 9804
rect 1950 9734 1954 9804
rect 1974 9734 1978 9804
rect 1998 9734 2002 9804
rect 2022 9734 2026 9804
rect 2046 9734 2050 9804
rect 2070 9734 2074 9804
rect 2094 9734 2098 9804
rect 2118 9734 2122 9804
rect 2142 9734 2146 9804
rect 2166 9734 2170 9804
rect 2190 9734 2194 9804
rect 2214 9734 2218 9804
rect 2238 9734 2242 9804
rect 2262 9734 2266 9804
rect 2286 9734 2290 9804
rect 2310 9734 2314 9804
rect 2334 9734 2338 9804
rect 2358 9734 2362 9804
rect 2382 9734 2386 9804
rect 2406 9734 2410 9804
rect 2430 9734 2434 9804
rect 2454 9734 2458 9804
rect 2478 9734 2482 9804
rect 2502 9734 2506 9804
rect 2526 9734 2530 9804
rect 2550 9734 2554 9804
rect 2574 9734 2578 9804
rect 2598 9734 2602 9804
rect 2622 9734 2626 9804
rect 2646 9734 2650 9804
rect 2670 9734 2674 9804
rect 2694 9734 2698 9804
rect 2718 9734 2722 9804
rect 2742 9734 2746 9804
rect 2766 9734 2770 9804
rect 2790 9734 2794 9804
rect 2814 9735 2818 9804
rect 2803 9734 2837 9735
rect 1861 9732 2837 9734
rect 1861 9731 1875 9732
rect 1878 9731 1885 9732
rect 1878 9710 1882 9731
rect 1902 9710 1906 9732
rect 1926 9710 1930 9732
rect 1950 9710 1954 9732
rect 1974 9710 1978 9732
rect 1998 9710 2002 9732
rect 2022 9710 2026 9732
rect 2046 9710 2050 9732
rect 2070 9710 2074 9732
rect 2094 9710 2098 9732
rect 2118 9710 2122 9732
rect 2142 9710 2146 9732
rect 2166 9710 2170 9732
rect 2190 9710 2194 9732
rect 2214 9710 2218 9732
rect 2238 9710 2242 9732
rect 2262 9710 2266 9732
rect 2286 9710 2290 9732
rect 2310 9710 2314 9732
rect 2334 9710 2338 9732
rect 2358 9710 2362 9732
rect 2382 9710 2386 9732
rect 2406 9710 2410 9732
rect 2430 9710 2434 9732
rect 2454 9710 2458 9732
rect 2478 9710 2482 9732
rect 2502 9710 2506 9732
rect 2526 9710 2530 9732
rect 2550 9710 2554 9732
rect 2574 9710 2578 9732
rect 2598 9710 2602 9732
rect 2622 9710 2626 9732
rect 2646 9710 2650 9732
rect 2670 9710 2674 9732
rect 2694 9710 2698 9732
rect 2718 9710 2722 9732
rect 2742 9710 2746 9732
rect 2766 9710 2770 9732
rect 2790 9710 2794 9732
rect 2803 9725 2808 9732
rect 2814 9725 2818 9732
rect 2813 9711 2818 9725
rect 2838 9710 2842 9804
rect 2862 9710 2866 9804
rect 2886 9710 2890 9804
rect 2910 9710 2914 9804
rect 2934 9710 2938 9804
rect 2958 9710 2962 9804
rect 2982 9710 2986 9804
rect 3006 9710 3010 9804
rect 3030 9710 3034 9804
rect 3043 9797 3048 9804
rect 3061 9803 3075 9804
rect 3053 9783 3058 9797
rect 3054 9711 3058 9783
rect 3043 9710 3075 9711
rect -1565 9708 3075 9710
rect -1555 9687 -1547 9701
rect -2393 9684 -1557 9686
rect -1530 9684 -1526 9708
rect -2371 9662 -2366 9684
rect -2348 9662 -2343 9684
rect -2325 9662 -2320 9684
rect -2309 9666 -2301 9676
rect -2068 9667 -2062 9672
rect -2317 9662 -2309 9666
rect -2060 9662 -2050 9667
rect -2000 9662 -1992 9684
rect -1806 9676 -1680 9682
rect -1854 9667 -1806 9672
rect -1655 9666 -1647 9676
rect -1972 9662 -1964 9663
rect -1958 9662 -1942 9664
rect -1844 9662 -1806 9665
rect -1663 9662 -1655 9666
rect -1642 9662 -1637 9684
rect -1619 9662 -1614 9684
rect -1571 9683 -1557 9684
rect -1554 9670 -1547 9684
rect -1530 9662 -1523 9683
rect -1506 9662 -1502 9708
rect -1482 9662 -1478 9708
rect -1458 9662 -1454 9708
rect -1434 9662 -1430 9708
rect -1410 9662 -1406 9708
rect -1386 9662 -1382 9708
rect -1362 9662 -1358 9708
rect -1338 9662 -1334 9708
rect -1314 9662 -1310 9708
rect -1290 9662 -1286 9708
rect -1266 9662 -1262 9708
rect -1242 9662 -1238 9708
rect -1218 9662 -1214 9708
rect -1194 9662 -1190 9708
rect -1170 9662 -1166 9708
rect -1146 9662 -1142 9708
rect -1122 9662 -1118 9708
rect -1098 9662 -1094 9708
rect -1074 9662 -1070 9708
rect -1050 9662 -1046 9708
rect -1026 9662 -1022 9708
rect -1002 9662 -998 9708
rect -978 9662 -974 9708
rect -954 9662 -950 9708
rect -930 9662 -926 9708
rect -906 9662 -902 9708
rect -882 9662 -878 9708
rect -858 9662 -854 9708
rect -834 9662 -830 9708
rect -810 9662 -806 9708
rect -786 9662 -782 9708
rect -762 9662 -758 9708
rect -738 9662 -734 9708
rect -714 9662 -710 9708
rect -690 9662 -686 9708
rect -666 9662 -662 9708
rect -618 9683 -614 9708
rect -653 9662 -621 9663
rect -2393 9660 -1557 9662
rect -1547 9660 -621 9662
rect -2371 9638 -2366 9660
rect -2348 9638 -2343 9660
rect -2325 9638 -2320 9660
rect -2060 9654 -2050 9660
rect -2309 9638 -2301 9648
rect -2060 9647 -2030 9654
rect -2000 9650 -1992 9660
rect -1972 9658 -1942 9660
rect -1958 9657 -1942 9658
rect -1844 9656 -1806 9660
rect -2068 9640 -2062 9647
rect -2062 9638 -2036 9640
rect -2393 9636 -2036 9638
rect -2030 9638 -2012 9640
rect -2004 9638 -1990 9650
rect -1844 9649 -1798 9654
rect -1806 9647 -1798 9649
rect -1854 9645 -1844 9647
rect -1854 9640 -1806 9645
rect -1864 9638 -1796 9639
rect -1655 9638 -1647 9648
rect -1642 9638 -1637 9660
rect -1619 9638 -1614 9660
rect -1571 9659 -1557 9660
rect -1554 9659 -1533 9660
rect -1554 9646 -1547 9659
rect -1530 9638 -1523 9660
rect -1506 9638 -1502 9660
rect -1482 9638 -1478 9660
rect -1458 9638 -1454 9660
rect -1434 9638 -1430 9660
rect -1410 9638 -1406 9660
rect -1386 9638 -1382 9660
rect -1362 9638 -1358 9660
rect -1338 9638 -1334 9660
rect -1314 9638 -1310 9660
rect -1290 9638 -1286 9660
rect -1266 9638 -1262 9660
rect -1242 9638 -1238 9660
rect -1218 9638 -1214 9660
rect -1194 9638 -1190 9660
rect -1170 9638 -1166 9660
rect -1146 9638 -1142 9660
rect -1122 9638 -1118 9660
rect -1098 9638 -1094 9660
rect -1074 9638 -1070 9660
rect -1050 9638 -1046 9660
rect -1026 9638 -1022 9660
rect -1002 9638 -998 9660
rect -978 9638 -974 9660
rect -954 9638 -950 9660
rect -930 9638 -926 9660
rect -906 9638 -902 9660
rect -882 9638 -878 9660
rect -858 9638 -854 9660
rect -834 9638 -830 9660
rect -810 9638 -806 9660
rect -786 9638 -782 9660
rect -762 9638 -758 9660
rect -738 9638 -734 9660
rect -714 9638 -710 9660
rect -690 9638 -686 9660
rect -666 9638 -662 9660
rect -653 9653 -648 9660
rect -635 9659 -621 9660
rect -618 9659 -611 9683
rect -643 9639 -638 9653
rect -642 9638 -638 9639
rect -594 9638 -590 9708
rect -570 9638 -566 9708
rect -546 9638 -542 9708
rect -522 9638 -518 9708
rect -498 9638 -494 9708
rect -474 9638 -470 9708
rect -450 9638 -446 9708
rect -426 9638 -422 9708
rect -402 9638 -398 9708
rect -378 9638 -374 9708
rect -354 9638 -350 9708
rect -330 9638 -326 9708
rect -306 9638 -302 9708
rect -282 9638 -278 9708
rect -258 9638 -254 9708
rect -234 9638 -230 9708
rect -210 9638 -206 9708
rect -197 9677 -192 9687
rect -186 9677 -182 9708
rect -187 9663 -182 9677
rect -197 9638 -163 9639
rect -162 9638 -158 9708
rect -138 9638 -134 9708
rect -114 9638 -110 9708
rect -90 9638 -86 9708
rect -66 9638 -62 9708
rect -42 9638 -38 9708
rect -18 9638 -14 9708
rect 6 9638 10 9708
rect 30 9638 34 9708
rect 54 9638 58 9708
rect 78 9638 82 9708
rect 102 9638 106 9708
rect 126 9638 130 9708
rect 150 9638 154 9708
rect 174 9638 178 9708
rect 198 9638 202 9708
rect 222 9638 226 9708
rect 246 9638 250 9708
rect 270 9638 274 9708
rect 294 9638 298 9708
rect 318 9638 322 9708
rect 342 9638 346 9708
rect 366 9638 370 9708
rect 390 9638 394 9708
rect 414 9638 418 9708
rect 438 9638 442 9708
rect 462 9638 466 9708
rect 486 9638 490 9708
rect 510 9638 514 9708
rect 534 9638 538 9708
rect 558 9638 562 9708
rect 582 9638 586 9708
rect 606 9638 610 9708
rect 630 9638 634 9708
rect 654 9638 658 9708
rect 678 9638 682 9708
rect 702 9638 706 9708
rect 726 9638 730 9708
rect 739 9653 744 9663
rect 750 9653 754 9708
rect 749 9639 754 9653
rect 774 9638 778 9708
rect 798 9638 802 9708
rect 822 9638 826 9708
rect 846 9638 850 9708
rect 870 9638 874 9708
rect 894 9638 898 9708
rect 918 9638 922 9708
rect 942 9638 946 9708
rect 966 9638 970 9708
rect 990 9638 994 9708
rect 1014 9638 1018 9708
rect 1038 9638 1042 9708
rect 1062 9638 1066 9708
rect 1086 9638 1090 9708
rect 1110 9638 1114 9708
rect 1134 9638 1138 9708
rect 1158 9638 1162 9708
rect 1182 9638 1186 9708
rect 1206 9638 1210 9708
rect 1230 9638 1234 9708
rect 1254 9638 1258 9708
rect 1278 9638 1282 9708
rect 1302 9638 1306 9708
rect 1326 9638 1330 9708
rect 1350 9638 1354 9708
rect 1374 9638 1378 9708
rect 1398 9638 1402 9708
rect 1422 9638 1426 9708
rect 1446 9638 1450 9708
rect 1470 9638 1474 9708
rect 1494 9638 1498 9708
rect 1518 9638 1522 9708
rect 1542 9638 1546 9708
rect 1566 9638 1570 9708
rect 1590 9638 1594 9708
rect 1614 9638 1618 9708
rect 1638 9638 1642 9708
rect 1662 9638 1666 9708
rect 1686 9638 1690 9708
rect 1710 9638 1714 9708
rect 1734 9638 1738 9708
rect 1758 9638 1762 9708
rect 1782 9638 1786 9708
rect 1806 9638 1810 9708
rect 1830 9638 1834 9708
rect 1854 9638 1858 9708
rect 1878 9638 1882 9708
rect 1902 9638 1906 9708
rect 1926 9638 1930 9708
rect 1950 9638 1954 9708
rect 1974 9638 1978 9708
rect 1998 9638 2002 9708
rect 2022 9639 2026 9708
rect 2011 9638 2045 9639
rect -2030 9636 -1557 9638
rect -1547 9636 2045 9638
rect -2371 9219 -2366 9636
rect -2361 9239 -2353 9249
rect -2348 9239 -2343 9636
rect -2351 9223 -2343 9239
rect -2371 9193 -2363 9219
rect -2383 9021 -2376 9031
rect -2371 9021 -2366 9193
rect -2373 9010 -2366 9021
rect -2348 9010 -2343 9223
rect -2325 9505 -2320 9636
rect -2317 9632 -2309 9636
rect -2060 9632 -2050 9636
rect -2060 9630 -2036 9632
rect -2060 9628 -2030 9630
rect -2292 9622 -2030 9628
rect -2092 9606 -2062 9608
rect -2094 9602 -2062 9606
rect -2309 9572 -2301 9581
rect -2317 9565 -2309 9572
rect -2309 9544 -2301 9552
rect -2251 9546 -2093 9552
rect -2317 9536 -2309 9544
rect -2154 9539 -2138 9542
rect -2084 9539 -2054 9544
rect -2143 9526 -2138 9532
rect -2325 9495 -2317 9505
rect -2325 9476 -2320 9495
rect -2317 9489 -2309 9495
rect -2243 9478 -2221 9486
rect -2211 9478 -2201 9498
rect -2073 9478 -2065 9496
rect -2000 9478 -1992 9636
rect -1844 9629 -1806 9636
rect -1663 9632 -1655 9636
rect -1844 9622 -1680 9628
rect -1854 9606 -1806 9608
rect -1854 9602 -1680 9606
rect -1915 9572 -1906 9582
rect -1846 9580 -1837 9582
rect -1790 9580 -1680 9582
rect -1655 9572 -1647 9578
rect -1905 9563 -1896 9572
rect -1837 9571 -1790 9572
rect -1837 9556 -1798 9569
rect -1663 9562 -1655 9572
rect -1798 9546 -1790 9551
rect -1837 9544 -1798 9546
rect -1655 9544 -1647 9550
rect -1846 9542 -1837 9544
rect -1846 9539 -1798 9542
rect -1837 9526 -1798 9536
rect -1663 9534 -1655 9544
rect -1671 9494 -1663 9502
rect -1655 9494 -1647 9496
rect -1663 9486 -1647 9494
rect -1642 9486 -1637 9636
rect -1885 9478 -1877 9480
rect -1708 9478 -1672 9480
rect -2243 9477 -2213 9478
rect -2325 9467 -2317 9476
rect -2259 9471 -2211 9477
rect -2183 9471 -1877 9478
rect -1869 9471 -1758 9478
rect -1710 9472 -1672 9478
rect -1710 9471 -1692 9472
rect -2211 9467 -2201 9471
rect -2325 9447 -2320 9467
rect -2317 9460 -2309 9467
rect -2211 9460 -2198 9467
rect -2325 9439 -2317 9447
rect -2300 9440 -2292 9450
rect -2243 9441 -2228 9452
rect -2211 9444 -2181 9460
rect -2211 9441 -2201 9444
rect -2325 9419 -2320 9439
rect -2317 9431 -2309 9439
rect -2325 9411 -2317 9419
rect -2325 9391 -2320 9411
rect -2317 9403 -2309 9411
rect -2325 9382 -2317 9391
rect -2325 9363 -2320 9382
rect -2317 9375 -2309 9382
rect -2325 9354 -2317 9363
rect -2325 9334 -2320 9354
rect -2317 9347 -2309 9354
rect -2325 9326 -2317 9334
rect -2290 9327 -2282 9440
rect -2251 9430 -2240 9434
rect -2211 9430 -2181 9434
rect -2251 9427 -2181 9430
rect -2176 9420 -2173 9422
rect -2240 9413 -2173 9420
rect -2169 9415 -2163 9470
rect -2073 9434 -2065 9471
rect -2073 9430 -2043 9434
rect -2000 9430 -1992 9471
rect -1915 9440 -1907 9449
rect -1963 9434 -1955 9440
rect -1963 9430 -1915 9434
rect -1885 9430 -1877 9471
rect -1875 9466 -1869 9470
rect -1829 9448 -1781 9450
rect -1847 9444 -1781 9448
rect -1778 9444 -1771 9470
rect -1758 9463 -1710 9470
rect -1718 9456 -1710 9463
rect -1768 9446 -1760 9456
rect -1718 9454 -1700 9456
rect -2146 9427 -2135 9430
rect -2105 9427 -2043 9430
rect -2035 9427 -1989 9430
rect -1973 9427 -1915 9430
rect -1907 9427 -1854 9430
rect -2073 9425 -2043 9427
rect -2135 9413 -2105 9420
rect -2065 9418 -2043 9425
rect -2243 9402 -2240 9411
rect -2221 9405 -2213 9413
rect -2211 9405 -2208 9413
rect -2203 9406 -2173 9413
rect -2251 9395 -2240 9402
rect -2211 9402 -2203 9405
rect -2211 9395 -2181 9402
rect -2073 9395 -2043 9402
rect -2203 9372 -2173 9379
rect -2262 9354 -2240 9364
rect -2203 9363 -2176 9372
rect -2083 9361 -2075 9371
rect -2040 9361 -2035 9365
rect -2073 9349 -2043 9361
rect -2028 9349 -2023 9361
rect -2000 9354 -1992 9427
rect -1963 9424 -1955 9427
rect -1963 9423 -1915 9424
rect -1955 9413 -1907 9420
rect -1885 9416 -1877 9427
rect -1837 9422 -1828 9438
rect -1758 9431 -1750 9446
rect -1758 9430 -1692 9431
rect -1837 9420 -1833 9422
rect -1837 9418 -1835 9420
rect -1887 9413 -1851 9416
rect -1750 9413 -1702 9420
rect -1885 9408 -1877 9413
rect -1963 9395 -1915 9402
rect -1905 9363 -1897 9408
rect -1857 9390 -1851 9413
rect -1760 9405 -1758 9406
rect -1837 9395 -1789 9402
rect -1758 9396 -1750 9402
rect -1758 9395 -1710 9396
rect -1955 9360 -1915 9363
rect -1963 9354 -1962 9356
rect -2000 9351 -1981 9354
rect -1965 9351 -1962 9354
rect -1955 9354 -1907 9358
rect -1885 9354 -1877 9373
rect -1857 9360 -1851 9372
rect -1750 9368 -1702 9375
rect -1829 9360 -1789 9362
rect -1766 9358 -1760 9368
rect -1829 9354 -1781 9358
rect -1756 9354 -1740 9358
rect -1680 9354 -1672 9472
rect -1671 9466 -1663 9474
rect -1645 9470 -1637 9486
rect -1663 9458 -1655 9466
rect -1671 9438 -1663 9446
rect -1663 9430 -1655 9438
rect -1671 9410 -1663 9418
rect -1671 9394 -1669 9407
rect -1663 9402 -1655 9410
rect -1671 9382 -1663 9390
rect -1663 9374 -1655 9382
rect -1671 9354 -1663 9362
rect -1955 9351 -1837 9354
rect -1829 9351 -1740 9354
rect -2206 9341 -2176 9344
rect -2206 9338 -2203 9341
rect -2161 9339 -2145 9348
rect -2073 9346 -2065 9349
rect -2073 9345 -2043 9346
rect -2028 9345 -2012 9349
rect -2073 9338 -2065 9344
rect -2203 9337 -2176 9338
rect -2065 9337 -2043 9338
rect -2262 9331 -2232 9337
rect -2176 9331 -2173 9337
rect -2043 9331 -2035 9337
rect -2325 9306 -2320 9326
rect -2317 9318 -2309 9326
rect -2153 9325 -2146 9329
rect -2325 9298 -2317 9306
rect -2300 9302 -2292 9312
rect -2325 9278 -2320 9298
rect -2317 9290 -2309 9298
rect -2325 9270 -2317 9278
rect -2325 9250 -2320 9270
rect -2317 9262 -2309 9270
rect -2290 9269 -2282 9302
rect -2273 9298 -2264 9303
rect -2206 9298 -2176 9303
rect -2262 9291 -2232 9296
rect -2198 9287 -2176 9298
rect -2198 9273 -2176 9281
rect -2166 9265 -2158 9313
rect -2143 9309 -2136 9325
rect -2143 9298 -2113 9303
rect -2073 9298 -2065 9303
rect -2065 9296 -2043 9298
rect -2043 9291 -2035 9296
rect -2065 9270 -2043 9285
rect -2006 9269 -2004 9285
rect -2265 9255 -2260 9261
rect -2143 9255 -2113 9262
rect -2270 9254 -2240 9255
rect -2270 9251 -2265 9254
rect -2325 9242 -2317 9250
rect -2325 9222 -2320 9242
rect -2317 9234 -2309 9242
rect -2113 9239 -2105 9249
rect -2291 9227 -2270 9234
rect -2198 9232 -2168 9234
rect -2135 9233 -2105 9234
rect -2103 9233 -2095 9239
rect -2113 9232 -2105 9233
rect -2065 9232 -2035 9234
rect -2000 9232 -1992 9351
rect -1963 9344 -1960 9351
rect -1915 9347 -1905 9351
rect -1963 9343 -1955 9344
rect -1963 9337 -1915 9343
rect -1989 9310 -1973 9313
rect -1915 9310 -1907 9317
rect -1990 9275 -1989 9296
rect -1983 9232 -1981 9295
rect -1885 9286 -1877 9351
rect -1789 9346 -1778 9351
rect -1837 9343 -1829 9344
rect -1837 9337 -1789 9343
rect -1756 9342 -1740 9351
rect -1837 9327 -1829 9337
rect -1872 9308 -1867 9318
rect -1789 9310 -1781 9317
rect -1776 9310 -1769 9327
rect -1756 9320 -1750 9342
rect -1671 9338 -1669 9349
rect -1663 9346 -1655 9354
rect -1671 9326 -1663 9334
rect -1663 9318 -1655 9326
rect -1702 9308 -1696 9314
rect -1955 9284 -1915 9286
rect -1963 9282 -1955 9284
rect -1963 9275 -1915 9282
rect -1963 9267 -1955 9275
rect -1963 9266 -1915 9267
rect -1973 9260 -1965 9263
rect -1955 9260 -1907 9264
rect -1974 9257 -1907 9260
rect -1973 9253 -1965 9257
rect -1963 9253 -1960 9255
rect -1963 9249 -1915 9253
rect -1963 9241 -1955 9249
rect -1963 9237 -1915 9241
rect -1963 9234 -1955 9237
rect -2240 9227 -2206 9232
rect -2198 9227 -2143 9232
rect -2113 9227 -1981 9232
rect -1915 9227 -1907 9234
rect -2270 9222 -2266 9226
rect -2086 9223 -2070 9227
rect -2325 9214 -2317 9222
rect -2270 9215 -2240 9222
rect -2206 9215 -2176 9222
rect -2325 9194 -2320 9214
rect -2317 9206 -2309 9214
rect -2270 9210 -2266 9215
rect -2270 9206 -2266 9209
rect -2198 9206 -2176 9213
rect -2166 9206 -2158 9223
rect -2143 9215 -2113 9222
rect -2198 9197 -2168 9201
rect -2325 9186 -2317 9194
rect -2143 9192 -2136 9206
rect -2085 9201 -2060 9202
rect -2039 9201 -2035 9210
rect -2135 9194 -2105 9201
rect -2085 9194 -2035 9201
rect -2029 9194 -2025 9201
rect -2325 9173 -2320 9186
rect -2317 9178 -2309 9186
rect -2235 9176 -2232 9179
rect -2325 9147 -2317 9173
rect -2325 9138 -2320 9147
rect -2325 9130 -2317 9138
rect -2135 9130 -2119 9143
rect -2000 9135 -1992 9227
rect -1983 9209 -1981 9227
rect -1955 9209 -1915 9210
rect -1862 9206 -1857 9308
rect -1706 9304 -1702 9308
rect -1829 9292 -1789 9300
rect -1671 9298 -1663 9306
rect -1849 9284 -1842 9292
rect -1790 9284 -1781 9292
rect -1663 9290 -1655 9298
rect -1837 9275 -1829 9282
rect -1758 9275 -1732 9282
rect -1748 9266 -1732 9275
rect -1671 9270 -1663 9278
rect -1829 9257 -1781 9264
rect -1663 9262 -1655 9270
rect -1829 9251 -1789 9255
rect -1768 9252 -1760 9262
rect -1758 9251 -1750 9252
rect -1671 9242 -1663 9250
rect -1837 9239 -1780 9242
rect -1758 9236 -1748 9242
rect -1708 9236 -1690 9242
rect -1829 9227 -1781 9234
rect -1680 9225 -1672 9242
rect -1663 9234 -1655 9242
rect -1829 9216 -1791 9222
rect -1758 9216 -1710 9218
rect -1758 9209 -1692 9216
rect -1671 9214 -1663 9222
rect -1955 9198 -1907 9201
rect -1791 9198 -1781 9201
rect -1991 9194 -1839 9198
rect -1791 9194 -1780 9198
rect -1680 9191 -1672 9209
rect -1663 9206 -1655 9214
rect -1839 9181 -1791 9188
rect -1671 9186 -1663 9194
rect -1829 9175 -1791 9179
rect -1671 9176 -1669 9186
rect -1663 9178 -1655 9186
rect -1680 9160 -1672 9175
rect -1642 9160 -1637 9470
rect -1619 9420 -1614 9636
rect -1571 9635 -1557 9636
rect -1554 9635 -1533 9636
rect -1530 9611 -1523 9636
rect -1619 9394 -1611 9420
rect -1768 9144 -1760 9154
rect -1758 9137 -1710 9144
rect -2325 9110 -2320 9130
rect -2317 9122 -2306 9130
rect -2031 9127 -1992 9135
rect -1750 9133 -1710 9137
rect -1674 9132 -1663 9138
rect -2307 9114 -2306 9122
rect -2149 9125 -2135 9126
rect -2149 9121 -2119 9125
rect -2024 9116 -2021 9125
rect -2325 9102 -2317 9110
rect -2325 9054 -2320 9102
rect -2317 9094 -2306 9102
rect -2185 9100 -2169 9112
rect -2056 9109 -2040 9113
rect -2021 9109 -2008 9116
rect -2056 9098 -2054 9108
rect -2056 9097 -2048 9098
rect -2307 9058 -2306 9066
rect -2111 9065 -2054 9071
rect -2325 9046 -2314 9054
rect -2104 9047 -2101 9051
rect -2325 9026 -2320 9046
rect -2314 9038 -2306 9046
rect -2104 9044 -2101 9046
rect -2084 9044 -2054 9045
rect -2000 9044 -1992 9127
rect -1758 9126 -1750 9127
rect -1758 9125 -1749 9126
rect -1758 9124 -1710 9125
rect -1663 9122 -1658 9132
rect -1831 9114 -1783 9118
rect -1784 9101 -1783 9114
rect -1674 9104 -1663 9110
rect -1826 9099 -1796 9100
rect -1663 9094 -1658 9104
rect -1654 9100 -1647 9110
rect -1644 9086 -1637 9100
rect -1758 9068 -1750 9071
rect -1758 9065 -1710 9068
rect -1844 9053 -1828 9055
rect -1844 9052 -1792 9053
rect -1828 9051 -1792 9052
rect -1772 9051 -1758 9059
rect -1750 9056 -1702 9063
rect -1750 9048 -1710 9052
rect -1700 9048 -1692 9068
rect -1674 9060 -1665 9068
rect -1674 9048 -1666 9056
rect -1758 9044 -1710 9045
rect -2307 9030 -2306 9038
rect -2139 9034 -2123 9043
rect -2111 9038 -2016 9044
rect -2139 9027 -2111 9034
rect -2325 9018 -2314 9026
rect -2177 9020 -2161 9021
rect -2141 9020 -2119 9022
rect -2104 9020 -2101 9038
rect -2076 9027 -2046 9032
rect -2325 9010 -2320 9018
rect -2314 9010 -2306 9018
rect -2076 9016 -2054 9022
rect -2021 9019 -2016 9038
rect -2000 9038 -1818 9044
rect -1802 9038 -1776 9044
rect -1760 9038 -1710 9044
rect -1666 9040 -1658 9048
rect -2189 9010 -2175 9015
rect -2373 9008 -2175 9010
rect -2373 9007 -2359 9008
rect -2371 8822 -2366 9007
rect -2348 8955 -2343 9008
rect -2325 8998 -2320 9008
rect -2307 9002 -2306 9008
rect -2189 9007 -2175 9008
rect -2149 9006 -2119 9015
rect -2084 9014 -2036 9015
rect -2000 9014 -1992 9038
rect -1758 9036 -1710 9038
rect -1758 9034 -1755 9036
rect -1828 9027 -1792 9034
rect -1768 9025 -1760 9032
rect -1758 9027 -1757 9034
rect -1710 9033 -1702 9034
rect -1750 9027 -1702 9033
rect -1674 9032 -1665 9040
rect -1768 9022 -1764 9025
rect -1758 9022 -1755 9027
rect -1818 9014 -1789 9022
rect -1758 9015 -1754 9022
rect -1750 9017 -1710 9022
rect -1674 9020 -1666 9028
rect -1758 9014 -1692 9015
rect -2084 9012 -1692 9014
rect -1666 9012 -1658 9020
rect -2084 9009 -1690 9012
rect -2084 9006 -2054 9009
rect -2046 9007 -1710 9009
rect -2325 8990 -2314 8998
rect -2076 8997 -2046 9004
rect -2325 8970 -2320 8990
rect -2314 8982 -2306 8990
rect -2076 8989 -2054 8995
rect -2084 8985 -2054 8987
rect -2104 8982 -2054 8985
rect -2307 8974 -2306 8982
rect -2084 8979 -2054 8982
rect -2348 8931 -2341 8955
rect -2325 8954 -2314 8970
rect -2325 8938 -2320 8954
rect -2309 8942 -2298 8954
rect -2070 8953 -2040 8955
rect -2070 8951 -2013 8953
rect -2314 8938 -2309 8942
rect -2070 8939 -2046 8946
rect -2040 8945 -2013 8951
rect -2348 8822 -2343 8931
rect -2325 8926 -2314 8938
rect -2181 8931 -2151 8938
rect -2167 8929 -2151 8931
rect -2129 8930 -2111 8938
rect -2076 8937 -2070 8938
rect -2000 8937 -1992 9007
rect -1758 9006 -1710 9007
rect -1680 9004 -1665 9012
rect -1750 8997 -1702 9004
rect -1680 9000 -1672 9004
rect -1680 8995 -1666 9000
rect -1836 8991 -1820 8992
rect -1837 8987 -1820 8991
rect -1750 8989 -1710 8995
rect -1674 8992 -1666 8995
rect -1837 8980 -1789 8987
rect -1758 8986 -1710 8987
rect -1760 8983 -1692 8986
rect -1666 8984 -1658 8992
rect -1837 8979 -1820 8980
rect -1764 8979 -1692 8983
rect -1674 8979 -1665 8984
rect -1680 8976 -1665 8979
rect -1850 8951 -1802 8955
rect -1829 8939 -1802 8946
rect -1802 8937 -1781 8938
rect -2078 8930 -2046 8937
rect -2040 8930 -1945 8937
rect -1929 8930 -1850 8937
rect -1829 8930 -1781 8937
rect -1750 8933 -1682 8938
rect -1680 8933 -1672 8976
rect -1666 8956 -1665 8966
rect -1655 8944 -1650 8954
rect -1666 8938 -1655 8944
rect -1750 8930 -1702 8933
rect -2325 8910 -2320 8926
rect -2309 8914 -2298 8926
rect -2145 8921 -2129 8928
rect -2070 8921 -2040 8928
rect -2314 8910 -2309 8914
rect -2141 8912 -2129 8921
rect -2070 8912 -2046 8919
rect -2325 8898 -2314 8910
rect -2076 8903 -2046 8910
rect -2325 8878 -2320 8898
rect -2062 8878 -2032 8879
rect -2000 8878 -1992 8930
rect -1666 8928 -1665 8938
rect -1850 8921 -1802 8928
rect -1829 8912 -1802 8919
rect -1655 8916 -1650 8926
rect -1829 8903 -1792 8911
rect -1666 8910 -1655 8916
rect -1666 8900 -1665 8910
rect -1942 8880 -1937 8892
rect -1850 8889 -1822 8890
rect -1850 8885 -1802 8889
rect -2325 8870 -2317 8878
rect -2062 8876 -1961 8878
rect -2325 8850 -2320 8870
rect -2317 8862 -2309 8870
rect -2062 8863 -2040 8874
rect -2032 8869 -1961 8876
rect -1947 8870 -1942 8878
rect -1842 8876 -1794 8879
rect -2070 8858 -2022 8862
rect -2325 8834 -2317 8850
rect -2325 8822 -2320 8834
rect -2309 8822 -2301 8834
rect -2000 8822 -1992 8869
rect -1942 8868 -1937 8870
rect -1932 8860 -1927 8868
rect -1912 8865 -1896 8871
rect -1842 8863 -1802 8874
rect -1671 8870 -1663 8878
rect -1663 8862 -1655 8870
rect -1850 8858 -1680 8862
rect -1671 8834 -1663 8850
rect -1655 8822 -1647 8834
rect -1642 8822 -1637 9086
rect -1619 9084 -1614 9394
rect -1619 9010 -1612 9034
rect -1619 8822 -1614 9010
rect -1530 8822 -1526 9611
rect -1506 8822 -1502 9636
rect -1482 8822 -1478 9636
rect -1458 8822 -1454 9636
rect -1434 8822 -1430 9636
rect -1410 8822 -1406 9636
rect -1386 8822 -1382 9636
rect -1362 8822 -1358 9636
rect -1338 8822 -1334 9636
rect -1314 8822 -1310 9636
rect -1290 8822 -1286 9636
rect -1266 8822 -1262 9636
rect -1242 8822 -1238 9636
rect -1218 8822 -1214 9636
rect -1194 8822 -1190 9636
rect -1170 8822 -1166 9636
rect -1146 8822 -1142 9636
rect -1122 8822 -1118 9636
rect -1098 8822 -1094 9636
rect -1074 8822 -1070 9636
rect -1050 8822 -1046 9636
rect -1026 8822 -1022 9636
rect -1002 8822 -998 9636
rect -978 8822 -974 9636
rect -954 8822 -950 9636
rect -930 8822 -926 9636
rect -906 8822 -902 9636
rect -882 8822 -878 9636
rect -858 8822 -854 9636
rect -834 8822 -830 9636
rect -810 8822 -806 9636
rect -786 8822 -782 9636
rect -762 8822 -758 9636
rect -738 8822 -734 9636
rect -714 8822 -710 9636
rect -690 8822 -686 9636
rect -666 8822 -662 9636
rect -642 8822 -638 9636
rect -618 9563 -611 9587
rect -629 8909 -624 8919
rect -618 8909 -614 9563
rect -619 8895 -614 8909
rect -629 8885 -624 8895
rect -619 8871 -614 8885
rect -618 8822 -614 8871
rect -594 8843 -590 9636
rect -2393 8820 -597 8822
rect -2371 8726 -2366 8820
rect -2348 8726 -2343 8820
rect -2325 8818 -2320 8820
rect -2317 8818 -2309 8820
rect -2325 8806 -2317 8818
rect -2061 8807 -2046 8808
rect -2325 8790 -2320 8806
rect -2309 8794 -2301 8806
rect -2070 8800 -2046 8807
rect -2000 8802 -1992 8820
rect -1974 8818 -1960 8820
rect -1663 8818 -1655 8820
rect -1960 8817 -1944 8818
rect -1980 8802 -1932 8807
rect -1671 8806 -1663 8818
rect -2061 8798 -2046 8800
rect -2032 8800 -1932 8802
rect -2032 8798 -1980 8800
rect -2317 8790 -2309 8794
rect -2062 8792 -2061 8798
rect -2062 8790 -2051 8791
rect -2325 8778 -2317 8790
rect -2062 8783 -2032 8790
rect -2062 8782 -2051 8783
rect -2325 8758 -2320 8778
rect -2325 8750 -2317 8758
rect -2325 8730 -2320 8750
rect -2317 8742 -2309 8750
rect -2325 8726 -2317 8730
rect -2000 8726 -1992 8798
rect -1655 8794 -1647 8806
rect -1990 8782 -1924 8791
rect -1904 8789 -1874 8791
rect -1842 8782 -1680 8791
rect -1663 8790 -1655 8794
rect -1671 8778 -1663 8790
rect -1671 8750 -1663 8758
rect -1663 8742 -1655 8750
rect -1671 8726 -1663 8730
rect -1642 8726 -1637 8820
rect -1619 8726 -1614 8820
rect -1530 8726 -1526 8820
rect -1506 8726 -1502 8820
rect -1482 8726 -1478 8820
rect -1458 8726 -1454 8820
rect -1434 8726 -1430 8820
rect -1410 8726 -1406 8820
rect -1386 8726 -1382 8820
rect -1362 8726 -1358 8820
rect -1338 8726 -1334 8820
rect -1314 8726 -1310 8820
rect -1290 8726 -1286 8820
rect -1266 8726 -1262 8820
rect -1242 8726 -1238 8820
rect -1218 8726 -1214 8820
rect -1194 8726 -1190 8820
rect -1170 8726 -1166 8820
rect -1146 8726 -1142 8820
rect -1122 8726 -1118 8820
rect -1098 8726 -1094 8820
rect -1074 8726 -1070 8820
rect -1050 8726 -1046 8820
rect -1026 8726 -1022 8820
rect -1002 8726 -998 8820
rect -978 8726 -974 8820
rect -954 8726 -950 8820
rect -930 8726 -926 8820
rect -906 8726 -902 8820
rect -882 8726 -878 8820
rect -858 8726 -854 8820
rect -834 8726 -830 8820
rect -810 8726 -806 8820
rect -786 8726 -782 8820
rect -762 8726 -758 8820
rect -738 8726 -734 8820
rect -714 8726 -710 8820
rect -690 8726 -686 8820
rect -666 8726 -662 8820
rect -642 8726 -638 8820
rect -618 8726 -614 8820
rect -611 8819 -597 8820
rect -594 8795 -587 8843
rect -594 8726 -590 8795
rect -570 8726 -566 9636
rect -546 8726 -542 9636
rect -522 8726 -518 9636
rect -498 8726 -494 9636
rect -474 8726 -470 9636
rect -450 8726 -446 9636
rect -426 8726 -422 9636
rect -402 8726 -398 9636
rect -378 8726 -374 9636
rect -354 8726 -350 9636
rect -330 8726 -326 9636
rect -306 8726 -302 9636
rect -282 8726 -278 9636
rect -258 8726 -254 9636
rect -234 8726 -230 9636
rect -210 8726 -206 9636
rect -197 9629 -192 9636
rect -187 9615 -182 9629
rect -186 8726 -182 9615
rect -162 9611 -158 9636
rect -162 9587 -155 9611
rect -162 9539 -155 9563
rect -162 8726 -158 9539
rect -138 8726 -134 9636
rect -114 8726 -110 9636
rect -90 8726 -86 9636
rect -66 8726 -62 9636
rect -53 9437 -48 9447
rect -42 9437 -38 9636
rect -43 9423 -38 9437
rect -42 8726 -38 9423
rect -18 9371 -14 9636
rect -18 9347 -11 9371
rect -18 8726 -14 9347
rect 6 8726 10 9636
rect 30 8726 34 9636
rect 54 8726 58 9636
rect 78 8726 82 9636
rect 102 8726 106 9636
rect 115 9485 120 9495
rect 126 9485 130 9636
rect 125 9471 130 9485
rect 115 9461 120 9471
rect 125 9447 130 9461
rect 126 8726 130 9447
rect 150 9419 154 9636
rect 150 9371 157 9419
rect 150 8726 154 9371
rect 174 8726 178 9636
rect 198 8726 202 9636
rect 222 8726 226 9636
rect 246 8726 250 9636
rect 270 8726 274 9636
rect 294 8726 298 9636
rect 318 8726 322 9636
rect 331 9077 336 9087
rect 342 9077 346 9636
rect 341 9063 346 9077
rect 331 9053 336 9063
rect 341 9039 346 9053
rect 342 8726 346 9039
rect 366 9011 370 9636
rect 366 8966 373 9011
rect 390 8966 394 9636
rect 414 8966 418 9636
rect 438 8966 442 9636
rect 462 8966 466 9636
rect 486 8966 490 9636
rect 510 8966 514 9636
rect 534 8966 538 9636
rect 558 8966 562 9636
rect 582 8966 586 9636
rect 606 8966 610 9636
rect 630 8966 634 9636
rect 654 8966 658 9636
rect 678 8966 682 9636
rect 702 8966 706 9636
rect 726 8966 730 9636
rect 739 9614 773 9615
rect 774 9614 778 9636
rect 798 9614 802 9636
rect 822 9614 826 9636
rect 846 9614 850 9636
rect 870 9614 874 9636
rect 894 9614 898 9636
rect 918 9614 922 9636
rect 942 9614 946 9636
rect 966 9614 970 9636
rect 990 9614 994 9636
rect 1014 9614 1018 9636
rect 1038 9614 1042 9636
rect 1062 9614 1066 9636
rect 1086 9614 1090 9636
rect 1110 9614 1114 9636
rect 1134 9614 1138 9636
rect 1158 9614 1162 9636
rect 1182 9614 1186 9636
rect 1206 9614 1210 9636
rect 1230 9614 1234 9636
rect 1254 9614 1258 9636
rect 1278 9614 1282 9636
rect 1302 9614 1306 9636
rect 1326 9614 1330 9636
rect 1350 9614 1354 9636
rect 1374 9614 1378 9636
rect 1398 9614 1402 9636
rect 1422 9614 1426 9636
rect 1446 9614 1450 9636
rect 1470 9614 1474 9636
rect 1494 9614 1498 9636
rect 1518 9614 1522 9636
rect 1542 9614 1546 9636
rect 1566 9614 1570 9636
rect 1590 9614 1594 9636
rect 1614 9614 1618 9636
rect 1638 9614 1642 9636
rect 1662 9614 1666 9636
rect 1686 9614 1690 9636
rect 1710 9614 1714 9636
rect 1734 9614 1738 9636
rect 1758 9614 1762 9636
rect 1782 9614 1786 9636
rect 1806 9614 1810 9636
rect 1830 9614 1834 9636
rect 1854 9614 1858 9636
rect 1878 9614 1882 9636
rect 1902 9614 1906 9636
rect 1926 9614 1930 9636
rect 1950 9614 1954 9636
rect 1974 9614 1978 9636
rect 1998 9614 2002 9636
rect 2011 9629 2016 9636
rect 2022 9629 2026 9636
rect 2021 9615 2026 9629
rect 2046 9614 2050 9708
rect 2070 9614 2074 9708
rect 2094 9614 2098 9708
rect 2118 9614 2122 9708
rect 2142 9614 2146 9708
rect 2166 9614 2170 9708
rect 2190 9614 2194 9708
rect 2214 9614 2218 9708
rect 2238 9614 2242 9708
rect 2262 9614 2266 9708
rect 2286 9614 2290 9708
rect 2310 9614 2314 9708
rect 2334 9614 2338 9708
rect 2358 9614 2362 9708
rect 2382 9614 2386 9708
rect 2406 9614 2410 9708
rect 2430 9614 2434 9708
rect 2454 9614 2458 9708
rect 2478 9614 2482 9708
rect 2502 9614 2506 9708
rect 2526 9614 2530 9708
rect 2550 9614 2554 9708
rect 2574 9614 2578 9708
rect 2598 9614 2602 9708
rect 2622 9614 2626 9708
rect 2646 9614 2650 9708
rect 2670 9614 2674 9708
rect 2694 9614 2698 9708
rect 2718 9614 2722 9708
rect 2742 9614 2746 9708
rect 2766 9614 2770 9708
rect 2790 9614 2794 9708
rect 2803 9677 2808 9687
rect 2813 9663 2818 9677
rect 2814 9614 2818 9663
rect 2838 9659 2842 9708
rect 2838 9635 2845 9659
rect 2862 9614 2866 9708
rect 2886 9614 2890 9708
rect 2910 9614 2914 9708
rect 2934 9614 2938 9708
rect 2958 9614 2962 9708
rect 2982 9614 2986 9708
rect 3006 9615 3010 9708
rect 3019 9677 3024 9687
rect 3030 9677 3034 9708
rect 3043 9701 3048 9708
rect 3054 9701 3058 9708
rect 3061 9707 3075 9708
rect 3053 9687 3058 9701
rect 3029 9663 3034 9677
rect 2995 9614 3029 9615
rect 739 9612 3029 9614
rect 739 9605 744 9612
rect 749 9591 754 9605
rect 750 8966 754 9591
rect 774 9587 778 9612
rect 774 9563 781 9587
rect 774 9515 781 9539
rect 774 8966 778 9515
rect 798 8966 802 9612
rect 822 8966 826 9612
rect 846 8966 850 9612
rect 870 8966 874 9612
rect 894 8966 898 9612
rect 918 8966 922 9612
rect 942 8966 946 9612
rect 966 8966 970 9612
rect 990 8966 994 9612
rect 1014 8966 1018 9612
rect 1038 8966 1042 9612
rect 1062 8966 1066 9612
rect 1086 8966 1090 9612
rect 1110 8966 1114 9612
rect 1134 8966 1138 9612
rect 1158 8966 1162 9612
rect 1182 8966 1186 9612
rect 1206 8966 1210 9612
rect 1230 8966 1234 9612
rect 1254 8966 1258 9612
rect 1278 8966 1282 9612
rect 1302 8966 1306 9612
rect 1326 8966 1330 9612
rect 1350 8966 1354 9612
rect 1374 8966 1378 9612
rect 1398 8966 1402 9612
rect 1422 8966 1426 9612
rect 1446 8966 1450 9612
rect 1470 8966 1474 9612
rect 1494 8966 1498 9612
rect 1518 8966 1522 9612
rect 1542 8966 1546 9612
rect 1566 8966 1570 9612
rect 1590 8966 1594 9612
rect 1614 8966 1618 9612
rect 1638 8966 1642 9612
rect 1662 8966 1666 9612
rect 1686 8966 1690 9612
rect 1710 8966 1714 9612
rect 1734 8966 1738 9612
rect 1758 8966 1762 9612
rect 1782 8966 1786 9612
rect 1806 8966 1810 9612
rect 1830 8966 1834 9612
rect 1854 8966 1858 9612
rect 1878 8966 1882 9612
rect 1902 8966 1906 9612
rect 1926 8966 1930 9612
rect 1950 8966 1954 9612
rect 1974 8966 1978 9612
rect 1998 8966 2002 9612
rect 2011 9581 2016 9591
rect 2021 9567 2026 9581
rect 2022 8966 2026 9567
rect 2046 9563 2050 9612
rect 2046 9539 2053 9563
rect 2046 9491 2053 9515
rect 2046 8966 2050 9491
rect 2070 8966 2074 9612
rect 2094 8966 2098 9612
rect 2118 8966 2122 9612
rect 2142 8966 2146 9612
rect 2166 8966 2170 9612
rect 2190 8966 2194 9612
rect 2214 8966 2218 9612
rect 2238 8966 2242 9612
rect 2262 8966 2266 9612
rect 2286 8966 2290 9612
rect 2310 8966 2314 9612
rect 2334 8966 2338 9612
rect 2358 8966 2362 9612
rect 2382 8966 2386 9612
rect 2406 8966 2410 9612
rect 2430 8966 2434 9612
rect 2454 8966 2458 9612
rect 2478 8966 2482 9612
rect 2502 8966 2506 9612
rect 2526 8966 2530 9612
rect 2550 8966 2554 9612
rect 2574 8966 2578 9612
rect 2598 8966 2602 9612
rect 2622 8966 2626 9612
rect 2646 8966 2650 9612
rect 2670 8966 2674 9612
rect 2694 8966 2698 9612
rect 2718 8966 2722 9612
rect 2742 8966 2746 9612
rect 2766 8966 2770 9612
rect 2790 8966 2794 9612
rect 2814 8966 2818 9612
rect 2838 9590 2845 9611
rect 2862 9590 2866 9612
rect 2886 9590 2890 9612
rect 2910 9590 2914 9612
rect 2934 9590 2938 9612
rect 2958 9590 2962 9612
rect 2982 9591 2986 9612
rect 2995 9605 3000 9612
rect 3006 9605 3010 9612
rect 3005 9591 3010 9605
rect 2971 9590 3005 9591
rect 2821 9588 3005 9590
rect 2821 9587 2835 9588
rect 2838 9587 2845 9588
rect 2838 8966 2842 9587
rect 2862 8966 2866 9588
rect 2886 8966 2890 9588
rect 2910 8966 2914 9588
rect 2923 9053 2928 9063
rect 2934 9053 2938 9588
rect 2947 9461 2952 9471
rect 2958 9461 2962 9588
rect 2971 9581 2976 9588
rect 2982 9581 2986 9588
rect 2981 9567 2986 9581
rect 2957 9447 2962 9461
rect 2933 9039 2938 9053
rect 2923 8966 2955 8967
rect 349 8964 2955 8966
rect 349 8963 363 8964
rect 366 8963 373 8964
rect 366 8726 370 8963
rect 390 8726 394 8964
rect 414 8726 418 8964
rect 438 8726 442 8964
rect 462 8726 466 8964
rect 486 8726 490 8964
rect 510 8726 514 8964
rect 534 8726 538 8964
rect 558 8726 562 8964
rect 582 8726 586 8964
rect 606 8726 610 8964
rect 630 8726 634 8964
rect 654 8726 658 8964
rect 678 8726 682 8964
rect 702 8726 706 8964
rect 726 8726 730 8964
rect 750 8726 754 8964
rect 774 8726 778 8964
rect 798 8726 802 8964
rect 822 8726 826 8964
rect 835 8765 840 8775
rect 846 8765 850 8964
rect 845 8751 850 8765
rect 835 8741 840 8751
rect 845 8727 850 8741
rect 846 8726 850 8727
rect 870 8726 874 8964
rect 894 8726 898 8964
rect 918 8726 922 8964
rect 942 8726 946 8964
rect 966 8726 970 8964
rect 990 8726 994 8964
rect 1014 8726 1018 8964
rect 1038 8726 1042 8964
rect 1062 8726 1066 8964
rect 1086 8726 1090 8964
rect 1110 8726 1114 8964
rect 1134 8726 1138 8964
rect 1158 8726 1162 8964
rect 1182 8726 1186 8964
rect 1206 8726 1210 8964
rect 1230 8726 1234 8964
rect 1254 8726 1258 8964
rect 1278 8726 1282 8964
rect 1302 8726 1306 8964
rect 1326 8726 1330 8964
rect 1350 8726 1354 8964
rect 1374 8726 1378 8964
rect 1398 8726 1402 8964
rect 1422 8726 1426 8964
rect 1446 8726 1450 8964
rect 1470 8726 1474 8964
rect 1494 8726 1498 8964
rect 1518 8726 1522 8964
rect 1542 8726 1546 8964
rect 1566 8726 1570 8964
rect 1590 8726 1594 8964
rect 1614 8726 1618 8964
rect 1638 8726 1642 8964
rect 1662 8726 1666 8964
rect 1686 8726 1690 8964
rect 1710 8726 1714 8964
rect 1734 8726 1738 8964
rect 1758 8726 1762 8964
rect 1782 8726 1786 8964
rect 1806 8726 1810 8964
rect 1830 8726 1834 8964
rect 1854 8726 1858 8964
rect 1878 8726 1882 8964
rect 1902 8726 1906 8964
rect 1926 8726 1930 8964
rect 1950 8726 1954 8964
rect 1974 8726 1978 8964
rect 1998 8726 2002 8964
rect 2022 8726 2026 8964
rect 2046 8726 2050 8964
rect 2070 8726 2074 8964
rect 2094 8726 2098 8964
rect 2118 8726 2122 8964
rect 2142 8726 2146 8964
rect 2166 8726 2170 8964
rect 2190 8726 2194 8964
rect 2214 8726 2218 8964
rect 2238 8726 2242 8964
rect 2262 8726 2266 8964
rect 2275 8885 2280 8895
rect 2286 8885 2290 8964
rect 2285 8871 2290 8885
rect 2275 8870 2309 8871
rect 2310 8870 2314 8964
rect 2334 8870 2338 8964
rect 2358 8870 2362 8964
rect 2382 8870 2386 8964
rect 2406 8870 2410 8964
rect 2430 8870 2434 8964
rect 2454 8870 2458 8964
rect 2478 8870 2482 8964
rect 2502 8870 2506 8964
rect 2526 8870 2530 8964
rect 2550 8870 2554 8964
rect 2574 8870 2578 8964
rect 2598 8870 2602 8964
rect 2622 8870 2626 8964
rect 2646 8870 2650 8964
rect 2670 8870 2674 8964
rect 2694 8870 2698 8964
rect 2718 8870 2722 8964
rect 2742 8870 2746 8964
rect 2766 8870 2770 8964
rect 2790 8870 2794 8964
rect 2814 8870 2818 8964
rect 2838 8870 2842 8964
rect 2862 8870 2866 8964
rect 2886 8870 2890 8964
rect 2910 8870 2914 8964
rect 2923 8957 2928 8964
rect 2941 8963 2955 8964
rect 2933 8943 2938 8957
rect 2934 8871 2938 8943
rect 2923 8870 2955 8871
rect 2275 8868 2955 8870
rect 2275 8861 2280 8868
rect 2285 8847 2290 8861
rect 2286 8726 2290 8847
rect 2310 8819 2314 8868
rect 2310 8771 2317 8819
rect 2310 8726 2314 8771
rect 2334 8726 2338 8868
rect 2358 8726 2362 8868
rect 2382 8726 2386 8868
rect 2406 8726 2410 8868
rect 2430 8726 2434 8868
rect 2454 8726 2458 8868
rect 2478 8726 2482 8868
rect 2502 8726 2506 8868
rect 2526 8726 2530 8868
rect 2550 8726 2554 8868
rect 2574 8726 2578 8868
rect 2598 8726 2602 8868
rect 2622 8726 2626 8868
rect 2646 8726 2650 8868
rect 2670 8726 2674 8868
rect 2694 8726 2698 8868
rect 2718 8726 2722 8868
rect 2742 8726 2746 8868
rect 2766 8726 2770 8868
rect 2790 8726 2794 8868
rect 2814 8726 2818 8868
rect 2838 8726 2842 8868
rect 2862 8726 2866 8868
rect 2886 8726 2890 8868
rect 2910 8726 2914 8868
rect 2923 8861 2928 8868
rect 2934 8861 2938 8868
rect 2941 8867 2955 8868
rect 2933 8847 2938 8861
rect 2923 8813 2928 8823
rect 2933 8799 2938 8813
rect 2923 8741 2928 8751
rect 2934 8741 2938 8799
rect 2933 8727 2938 8741
rect 2947 8737 2955 8741
rect 2941 8727 2947 8737
rect 2923 8726 2955 8727
rect -2393 8724 2955 8726
rect -2371 8678 -2366 8724
rect -2348 8678 -2343 8724
rect -2325 8718 -2317 8724
rect -2018 8722 -2004 8724
rect -2325 8702 -2320 8718
rect -2317 8714 -2309 8718
rect -2069 8716 -2053 8718
rect -2309 8702 -2301 8714
rect -2096 8705 -2095 8711
rect -2000 8706 -1992 8724
rect -1671 8718 -1663 8724
rect -1663 8714 -1655 8718
rect -1977 8707 -1929 8713
rect -2112 8702 -2095 8705
rect -2325 8690 -2317 8702
rect -2325 8678 -2320 8690
rect -2317 8686 -2309 8690
rect -2112 8689 -2096 8702
rect -2059 8698 -2053 8705
rect -2027 8704 -1992 8706
rect -2059 8694 -2045 8698
rect -2018 8696 -2017 8698
rect -2083 8689 -2053 8690
rect -2019 8688 -2017 8692
rect -2309 8678 -2301 8686
rect -2017 8682 -2009 8688
rect -2000 8682 -1992 8704
rect -1972 8690 -1929 8705
rect -1655 8702 -1647 8714
rect -1671 8690 -1663 8702
rect -1972 8689 -1924 8690
rect -1663 8686 -1655 8690
rect -2033 8678 -1992 8682
rect -1655 8678 -1647 8686
rect -1642 8678 -1637 8724
rect -1619 8678 -1614 8724
rect -1530 8678 -1526 8724
rect -1506 8678 -1502 8724
rect -1482 8678 -1478 8724
rect -1458 8678 -1454 8724
rect -1434 8678 -1430 8724
rect -1410 8678 -1406 8724
rect -1386 8678 -1382 8724
rect -1362 8678 -1358 8724
rect -1338 8678 -1334 8724
rect -1314 8678 -1310 8724
rect -1290 8678 -1286 8724
rect -1266 8678 -1262 8724
rect -1242 8678 -1238 8724
rect -1218 8678 -1214 8724
rect -1194 8678 -1190 8724
rect -1170 8678 -1166 8724
rect -1146 8678 -1142 8724
rect -1122 8678 -1118 8724
rect -1098 8678 -1094 8724
rect -1074 8678 -1070 8724
rect -1050 8678 -1046 8724
rect -1026 8678 -1022 8724
rect -1002 8678 -998 8724
rect -978 8678 -974 8724
rect -954 8678 -950 8724
rect -930 8678 -926 8724
rect -906 8678 -902 8724
rect -882 8678 -878 8724
rect -858 8678 -854 8724
rect -834 8678 -830 8724
rect -810 8678 -806 8724
rect -786 8678 -782 8724
rect -762 8678 -758 8724
rect -738 8678 -734 8724
rect -714 8678 -710 8724
rect -690 8678 -686 8724
rect -666 8678 -662 8724
rect -642 8678 -638 8724
rect -618 8678 -614 8724
rect -594 8678 -590 8724
rect -570 8678 -566 8724
rect -546 8678 -542 8724
rect -522 8678 -518 8724
rect -498 8678 -494 8724
rect -474 8678 -470 8724
rect -450 8678 -446 8724
rect -426 8678 -422 8724
rect -402 8678 -398 8724
rect -378 8678 -374 8724
rect -354 8678 -350 8724
rect -330 8678 -326 8724
rect -306 8678 -302 8724
rect -282 8678 -278 8724
rect -258 8678 -254 8724
rect -234 8678 -230 8724
rect -210 8678 -206 8724
rect -186 8678 -182 8724
rect -162 8678 -158 8724
rect -138 8678 -134 8724
rect -114 8678 -110 8724
rect -90 8678 -86 8724
rect -66 8678 -62 8724
rect -42 8678 -38 8724
rect -18 8678 -14 8724
rect 6 8678 10 8724
rect 30 8678 34 8724
rect 54 8678 58 8724
rect 78 8678 82 8724
rect 102 8678 106 8724
rect 126 8678 130 8724
rect 150 8678 154 8724
rect 174 8678 178 8724
rect 198 8678 202 8724
rect 222 8678 226 8724
rect 246 8678 250 8724
rect 270 8678 274 8724
rect 294 8678 298 8724
rect 318 8678 322 8724
rect 342 8678 346 8724
rect 366 8678 370 8724
rect 390 8678 394 8724
rect 414 8678 418 8724
rect 438 8678 442 8724
rect 462 8678 466 8724
rect 486 8678 490 8724
rect 510 8678 514 8724
rect 534 8678 538 8724
rect 558 8678 562 8724
rect 582 8678 586 8724
rect 606 8678 610 8724
rect 630 8678 634 8724
rect 654 8678 658 8724
rect 678 8678 682 8724
rect 702 8678 706 8724
rect 726 8678 730 8724
rect 750 8678 754 8724
rect 774 8678 778 8724
rect 798 8678 802 8724
rect 822 8678 826 8724
rect 846 8678 850 8724
rect 870 8699 874 8724
rect -2393 8676 867 8678
rect -2371 8558 -2366 8676
rect -2348 8558 -2343 8676
rect -2325 8674 -2320 8676
rect -2309 8674 -2301 8676
rect -2325 8662 -2317 8674
rect -2325 8642 -2320 8662
rect -2317 8658 -2309 8662
rect -2325 8634 -2317 8642
rect -2325 8614 -2320 8634
rect -2317 8626 -2309 8634
rect -2117 8625 -2095 8635
rect -2045 8632 -2037 8646
rect -2325 8598 -2317 8614
rect -2325 8582 -2320 8598
rect -2309 8586 -2301 8598
rect -2317 8582 -2309 8586
rect -2117 8584 -2095 8591
rect -2069 8590 -2041 8598
rect -2017 8596 -2015 8598
rect -2325 8570 -2317 8582
rect -2125 8575 -2095 8582
rect -2047 8580 -2011 8582
rect -2059 8578 -2011 8580
rect -2000 8578 -1992 8676
rect -1655 8674 -1647 8676
rect -1671 8662 -1663 8674
rect -1663 8658 -1655 8662
rect -1969 8625 -1929 8637
rect -1671 8634 -1663 8642
rect -1663 8626 -1655 8634
rect -1671 8598 -1663 8614
rect -1655 8586 -1647 8598
rect -1663 8582 -1655 8586
rect -2125 8573 -2117 8575
rect -2059 8574 -2045 8578
rect -2021 8575 -1992 8578
rect -1977 8575 -1929 8582
rect -2325 8558 -2320 8570
rect -2309 8558 -2301 8570
rect -2131 8565 -2129 8570
rect -2125 8567 -2095 8573
rect -2021 8568 -2009 8572
rect -2125 8565 -2117 8567
rect -2133 8558 -2129 8565
rect -2117 8558 -2087 8565
rect -2025 8562 -2021 8568
rect -2000 8562 -1992 8575
rect -1969 8567 -1929 8573
rect -1671 8570 -1663 8582
rect -2033 8558 -1992 8562
rect -1969 8558 -1921 8565
rect -1655 8558 -1647 8570
rect -1642 8558 -1637 8676
rect -1619 8558 -1614 8676
rect -1530 8558 -1526 8676
rect -1506 8558 -1502 8676
rect -1482 8558 -1478 8676
rect -1458 8558 -1454 8676
rect -1434 8558 -1430 8676
rect -1410 8558 -1406 8676
rect -1386 8558 -1382 8676
rect -1362 8558 -1358 8676
rect -1338 8558 -1334 8676
rect -1314 8558 -1310 8676
rect -1290 8558 -1286 8676
rect -1266 8558 -1262 8676
rect -1242 8558 -1238 8676
rect -1218 8558 -1214 8676
rect -1194 8558 -1190 8676
rect -1170 8558 -1166 8676
rect -1146 8558 -1142 8676
rect -1122 8558 -1118 8676
rect -1098 8558 -1094 8676
rect -1074 8558 -1070 8676
rect -1050 8558 -1046 8676
rect -1026 8558 -1022 8676
rect -1002 8558 -998 8676
rect -978 8558 -974 8676
rect -954 8558 -950 8676
rect -930 8558 -926 8676
rect -906 8558 -902 8676
rect -882 8558 -878 8676
rect -858 8558 -854 8676
rect -834 8558 -830 8676
rect -810 8558 -806 8676
rect -786 8558 -782 8676
rect -762 8558 -758 8676
rect -738 8558 -734 8676
rect -714 8558 -710 8676
rect -690 8558 -686 8676
rect -666 8558 -662 8676
rect -642 8558 -638 8676
rect -618 8558 -614 8676
rect -594 8558 -590 8676
rect -570 8558 -566 8676
rect -546 8558 -542 8676
rect -522 8558 -518 8676
rect -498 8558 -494 8676
rect -474 8558 -470 8676
rect -450 8558 -446 8676
rect -426 8558 -422 8676
rect -402 8558 -398 8676
rect -378 8558 -374 8676
rect -354 8558 -350 8676
rect -330 8558 -326 8676
rect -306 8558 -302 8676
rect -282 8558 -278 8676
rect -258 8558 -254 8676
rect -234 8558 -230 8676
rect -210 8558 -206 8676
rect -186 8558 -182 8676
rect -162 8558 -158 8676
rect -138 8558 -134 8676
rect -114 8558 -110 8676
rect -90 8558 -86 8676
rect -66 8558 -62 8676
rect -42 8558 -38 8676
rect -18 8558 -14 8676
rect 6 8558 10 8676
rect 30 8558 34 8676
rect 54 8558 58 8676
rect 78 8558 82 8676
rect 102 8558 106 8676
rect 126 8558 130 8676
rect 150 8558 154 8676
rect 174 8558 178 8676
rect 198 8558 202 8676
rect 222 8558 226 8676
rect 246 8558 250 8676
rect 270 8558 274 8676
rect 294 8558 298 8676
rect 318 8558 322 8676
rect 342 8558 346 8676
rect 366 8559 370 8676
rect 355 8558 389 8559
rect -2393 8556 389 8558
rect -2371 8462 -2366 8556
rect -2348 8462 -2343 8556
rect -2325 8554 -2320 8556
rect -2317 8554 -2309 8556
rect -2131 8554 -2129 8556
rect -2125 8554 -2095 8556
rect -2325 8542 -2317 8554
rect -2117 8549 -2095 8554
rect -2325 8522 -2320 8542
rect -2325 8514 -2317 8522
rect -2325 8462 -2320 8514
rect -2317 8506 -2309 8514
rect -2117 8505 -2095 8515
rect -2045 8512 -2037 8526
rect -2309 8466 -2301 8476
rect -2087 8472 -2076 8480
rect -2017 8476 -2015 8483
rect -2317 8462 -2309 8466
rect -2092 8464 -2087 8472
rect -2092 8462 -2077 8463
rect -2000 8462 -1992 8556
rect -1663 8554 -1655 8556
rect -1671 8542 -1663 8554
rect -1969 8505 -1929 8517
rect -1671 8514 -1663 8522
rect -1663 8506 -1655 8514
rect -1655 8466 -1647 8476
rect -1928 8462 -1924 8463
rect -1854 8462 -1680 8463
rect -1663 8462 -1655 8466
rect -1642 8462 -1637 8556
rect -1619 8462 -1614 8556
rect -1530 8462 -1526 8556
rect -1506 8462 -1502 8556
rect -1482 8462 -1478 8556
rect -1458 8462 -1454 8556
rect -1434 8462 -1430 8556
rect -1410 8462 -1406 8556
rect -1386 8462 -1382 8556
rect -1362 8462 -1358 8556
rect -1338 8462 -1334 8556
rect -1314 8462 -1310 8556
rect -1290 8462 -1286 8556
rect -1266 8462 -1262 8556
rect -1242 8462 -1238 8556
rect -1218 8462 -1214 8556
rect -1194 8462 -1190 8556
rect -1170 8462 -1166 8556
rect -1146 8462 -1142 8556
rect -1122 8462 -1118 8556
rect -1098 8462 -1094 8556
rect -1074 8462 -1070 8556
rect -1050 8462 -1046 8556
rect -1026 8462 -1022 8556
rect -1002 8463 -998 8556
rect -1013 8462 -979 8463
rect -2393 8460 -979 8462
rect -2371 8438 -2366 8460
rect -2348 8438 -2343 8460
rect -2325 8438 -2320 8460
rect -2092 8455 -2037 8460
rect -2021 8455 -1969 8460
rect -1921 8455 -1913 8460
rect -1854 8456 -1680 8460
rect -2100 8453 -2092 8454
rect -2309 8438 -2301 8448
rect -2100 8447 -2087 8453
rect -2051 8440 -2026 8442
rect -2062 8438 -2012 8440
rect -2000 8438 -1992 8455
rect -1969 8447 -1921 8454
rect -1969 8438 -1964 8447
rect -1864 8438 -1796 8439
rect -1655 8438 -1647 8448
rect -1642 8438 -1637 8460
rect -1619 8438 -1614 8460
rect -1530 8438 -1526 8460
rect -1506 8438 -1502 8460
rect -1482 8438 -1478 8460
rect -1458 8438 -1454 8460
rect -1434 8438 -1430 8460
rect -1410 8438 -1406 8460
rect -1386 8438 -1382 8460
rect -1362 8438 -1358 8460
rect -1338 8438 -1334 8460
rect -1314 8438 -1310 8460
rect -1290 8438 -1286 8460
rect -1266 8438 -1262 8460
rect -1242 8438 -1238 8460
rect -1218 8438 -1214 8460
rect -1194 8438 -1190 8460
rect -1170 8438 -1166 8460
rect -1146 8438 -1142 8460
rect -1122 8438 -1118 8460
rect -1098 8438 -1094 8460
rect -1074 8438 -1070 8460
rect -1050 8438 -1046 8460
rect -1026 8438 -1022 8460
rect -1013 8453 -1008 8460
rect -1002 8453 -998 8460
rect -1003 8439 -998 8453
rect -978 8438 -974 8556
rect -954 8438 -950 8556
rect -930 8439 -926 8556
rect -941 8438 -907 8439
rect -2393 8436 -907 8438
rect -2371 8390 -2366 8436
rect -2348 8390 -2343 8436
rect -2325 8390 -2320 8436
rect -2317 8432 -2309 8436
rect -2105 8429 -2092 8432
rect -2092 8406 -2062 8408
rect -2094 8402 -2062 8406
rect -2000 8390 -1992 8436
rect -1663 8432 -1655 8436
rect -1969 8429 -1921 8432
rect -1854 8406 -1806 8408
rect -1854 8402 -1680 8406
rect -1642 8390 -1637 8436
rect -1619 8390 -1614 8436
rect -1530 8390 -1526 8436
rect -1506 8390 -1502 8436
rect -1482 8390 -1478 8436
rect -1458 8390 -1454 8436
rect -1434 8390 -1430 8436
rect -1410 8390 -1406 8436
rect -1386 8390 -1382 8436
rect -1362 8390 -1358 8436
rect -1338 8390 -1334 8436
rect -1314 8390 -1310 8436
rect -1290 8390 -1286 8436
rect -1266 8390 -1262 8436
rect -1242 8390 -1238 8436
rect -1218 8390 -1214 8436
rect -1194 8390 -1190 8436
rect -1170 8390 -1166 8436
rect -1146 8390 -1142 8436
rect -1122 8390 -1118 8436
rect -1098 8390 -1094 8436
rect -1074 8390 -1070 8436
rect -1050 8390 -1046 8436
rect -1026 8390 -1022 8436
rect -1013 8405 -1008 8415
rect -1003 8391 -998 8405
rect -1002 8390 -998 8391
rect -978 8390 -974 8436
rect -954 8390 -950 8436
rect -941 8429 -936 8436
rect -930 8429 -926 8436
rect -931 8415 -926 8429
rect -906 8390 -902 8556
rect -882 8390 -878 8556
rect -858 8390 -854 8556
rect -834 8390 -830 8556
rect -810 8390 -806 8556
rect -786 8390 -782 8556
rect -762 8390 -758 8556
rect -738 8390 -734 8556
rect -714 8390 -710 8556
rect -690 8390 -686 8556
rect -666 8390 -662 8556
rect -642 8390 -638 8556
rect -618 8390 -614 8556
rect -594 8390 -590 8556
rect -570 8390 -566 8556
rect -546 8390 -542 8556
rect -522 8390 -518 8556
rect -498 8390 -494 8556
rect -474 8390 -470 8556
rect -450 8390 -446 8556
rect -426 8390 -422 8556
rect -402 8390 -398 8556
rect -378 8390 -374 8556
rect -354 8390 -350 8556
rect -330 8390 -326 8556
rect -306 8390 -302 8556
rect -282 8390 -278 8556
rect -258 8390 -254 8556
rect -234 8390 -230 8556
rect -210 8390 -206 8556
rect -186 8390 -182 8556
rect -162 8390 -158 8556
rect -138 8390 -134 8556
rect -114 8390 -110 8556
rect -90 8390 -86 8556
rect -66 8390 -62 8556
rect -42 8390 -38 8556
rect -18 8390 -14 8556
rect 6 8390 10 8556
rect 30 8390 34 8556
rect 54 8390 58 8556
rect 78 8390 82 8556
rect 102 8390 106 8556
rect 126 8390 130 8556
rect 150 8390 154 8556
rect 174 8390 178 8556
rect 198 8390 202 8556
rect 222 8390 226 8556
rect 246 8390 250 8556
rect 270 8390 274 8556
rect 294 8390 298 8556
rect 318 8390 322 8556
rect 331 8525 336 8535
rect 342 8525 346 8556
rect 355 8549 360 8556
rect 366 8549 370 8556
rect 365 8535 370 8549
rect 355 8525 360 8535
rect 341 8511 346 8525
rect 365 8511 370 8525
rect 331 8510 365 8511
rect 366 8510 370 8511
rect 390 8510 394 8676
rect 414 8510 418 8676
rect 438 8510 442 8676
rect 462 8510 466 8676
rect 486 8510 490 8676
rect 510 8510 514 8676
rect 534 8510 538 8676
rect 558 8510 562 8676
rect 582 8510 586 8676
rect 606 8510 610 8676
rect 630 8510 634 8676
rect 654 8510 658 8676
rect 678 8510 682 8676
rect 702 8510 706 8676
rect 726 8510 730 8676
rect 750 8510 754 8676
rect 774 8510 778 8676
rect 798 8510 802 8676
rect 822 8510 826 8676
rect 846 8510 850 8676
rect 853 8675 867 8676
rect 870 8654 877 8699
rect 894 8654 898 8724
rect 918 8654 922 8724
rect 942 8654 946 8724
rect 966 8654 970 8724
rect 990 8654 994 8724
rect 1014 8654 1018 8724
rect 1038 8654 1042 8724
rect 1062 8654 1066 8724
rect 1086 8654 1090 8724
rect 1110 8654 1114 8724
rect 1134 8654 1138 8724
rect 1158 8654 1162 8724
rect 1182 8654 1186 8724
rect 1206 8655 1210 8724
rect 1195 8654 1229 8655
rect 853 8652 1229 8654
rect 853 8651 867 8652
rect 870 8651 877 8652
rect 870 8510 874 8651
rect 894 8510 898 8652
rect 918 8510 922 8652
rect 942 8510 946 8652
rect 966 8510 970 8652
rect 990 8510 994 8652
rect 1014 8510 1018 8652
rect 1038 8510 1042 8652
rect 1062 8510 1066 8652
rect 1086 8510 1090 8652
rect 1110 8510 1114 8652
rect 1134 8510 1138 8652
rect 1158 8510 1162 8652
rect 1182 8510 1186 8652
rect 1195 8645 1200 8652
rect 1206 8645 1210 8652
rect 1205 8631 1210 8645
rect 1195 8630 1229 8631
rect 1230 8630 1234 8724
rect 1254 8630 1258 8724
rect 1278 8630 1282 8724
rect 1302 8630 1306 8724
rect 1326 8630 1330 8724
rect 1350 8630 1354 8724
rect 1374 8630 1378 8724
rect 1398 8630 1402 8724
rect 1422 8630 1426 8724
rect 1446 8630 1450 8724
rect 1470 8630 1474 8724
rect 1494 8630 1498 8724
rect 1518 8630 1522 8724
rect 1542 8630 1546 8724
rect 1566 8630 1570 8724
rect 1590 8630 1594 8724
rect 1614 8630 1618 8724
rect 1638 8630 1642 8724
rect 1662 8630 1666 8724
rect 1686 8630 1690 8724
rect 1710 8630 1714 8724
rect 1734 8630 1738 8724
rect 1758 8630 1762 8724
rect 1782 8630 1786 8724
rect 1806 8630 1810 8724
rect 1830 8630 1834 8724
rect 1854 8630 1858 8724
rect 1878 8630 1882 8724
rect 1902 8630 1906 8724
rect 1926 8630 1930 8724
rect 1950 8630 1954 8724
rect 1974 8630 1978 8724
rect 1998 8630 2002 8724
rect 2022 8630 2026 8724
rect 2046 8630 2050 8724
rect 2059 8669 2064 8679
rect 2070 8669 2074 8724
rect 2069 8655 2074 8669
rect 2059 8654 2093 8655
rect 2094 8654 2098 8724
rect 2118 8654 2122 8724
rect 2142 8654 2146 8724
rect 2166 8654 2170 8724
rect 2190 8654 2194 8724
rect 2214 8654 2218 8724
rect 2238 8654 2242 8724
rect 2262 8654 2266 8724
rect 2286 8654 2290 8724
rect 2310 8654 2314 8724
rect 2334 8654 2338 8724
rect 2358 8654 2362 8724
rect 2382 8654 2386 8724
rect 2406 8654 2410 8724
rect 2430 8654 2434 8724
rect 2454 8654 2458 8724
rect 2478 8654 2482 8724
rect 2502 8654 2506 8724
rect 2526 8654 2530 8724
rect 2550 8654 2554 8724
rect 2574 8654 2578 8724
rect 2598 8654 2602 8724
rect 2622 8654 2626 8724
rect 2646 8654 2650 8724
rect 2670 8654 2674 8724
rect 2694 8654 2698 8724
rect 2718 8654 2722 8724
rect 2742 8654 2746 8724
rect 2766 8654 2770 8724
rect 2790 8654 2794 8724
rect 2814 8654 2818 8724
rect 2838 8654 2842 8724
rect 2862 8654 2866 8724
rect 2886 8654 2890 8724
rect 2910 8654 2914 8724
rect 2923 8717 2928 8724
rect 2941 8723 2955 8724
rect 2933 8703 2938 8717
rect 2934 8655 2938 8703
rect 2923 8654 2955 8655
rect 2059 8652 2955 8654
rect 2059 8645 2064 8652
rect 2069 8631 2074 8645
rect 2070 8630 2074 8631
rect 2094 8630 2098 8652
rect 2118 8630 2122 8652
rect 2142 8630 2146 8652
rect 2166 8630 2170 8652
rect 2190 8630 2194 8652
rect 2214 8630 2218 8652
rect 2238 8630 2242 8652
rect 2262 8630 2266 8652
rect 2286 8630 2290 8652
rect 2310 8630 2314 8652
rect 2334 8630 2338 8652
rect 2358 8630 2362 8652
rect 2382 8630 2386 8652
rect 2406 8630 2410 8652
rect 2430 8630 2434 8652
rect 2454 8630 2458 8652
rect 2478 8630 2482 8652
rect 2502 8630 2506 8652
rect 2526 8630 2530 8652
rect 2550 8630 2554 8652
rect 2574 8630 2578 8652
rect 2598 8630 2602 8652
rect 2622 8630 2626 8652
rect 2646 8630 2650 8652
rect 2670 8630 2674 8652
rect 2694 8630 2698 8652
rect 2718 8630 2722 8652
rect 2742 8630 2746 8652
rect 2766 8630 2770 8652
rect 2790 8630 2794 8652
rect 2814 8630 2818 8652
rect 2838 8630 2842 8652
rect 2862 8630 2866 8652
rect 2886 8630 2890 8652
rect 2910 8631 2914 8652
rect 2923 8645 2928 8652
rect 2934 8645 2938 8652
rect 2941 8651 2955 8652
rect 2933 8631 2938 8645
rect 2947 8641 2955 8645
rect 2941 8631 2947 8641
rect 2899 8630 2933 8631
rect 1195 8628 2933 8630
rect 1195 8621 1200 8628
rect 1205 8607 1210 8621
rect 1206 8510 1210 8607
rect 1230 8579 1234 8628
rect 1230 8534 1237 8579
rect 1254 8534 1258 8628
rect 1278 8534 1282 8628
rect 1302 8534 1306 8628
rect 1326 8534 1330 8628
rect 1350 8534 1354 8628
rect 1374 8534 1378 8628
rect 1398 8534 1402 8628
rect 1422 8534 1426 8628
rect 1446 8534 1450 8628
rect 1470 8534 1474 8628
rect 1494 8534 1498 8628
rect 1518 8534 1522 8628
rect 1542 8534 1546 8628
rect 1566 8534 1570 8628
rect 1590 8534 1594 8628
rect 1614 8534 1618 8628
rect 1638 8534 1642 8628
rect 1662 8534 1666 8628
rect 1686 8534 1690 8628
rect 1710 8534 1714 8628
rect 1734 8534 1738 8628
rect 1758 8534 1762 8628
rect 1782 8534 1786 8628
rect 1806 8534 1810 8628
rect 1830 8534 1834 8628
rect 1854 8534 1858 8628
rect 1878 8534 1882 8628
rect 1902 8534 1906 8628
rect 1926 8534 1930 8628
rect 1950 8534 1954 8628
rect 1974 8534 1978 8628
rect 1998 8534 2002 8628
rect 2022 8534 2026 8628
rect 2046 8534 2050 8628
rect 2070 8534 2074 8628
rect 2094 8603 2098 8628
rect 2094 8555 2101 8603
rect 2094 8534 2098 8555
rect 2118 8534 2122 8628
rect 2142 8534 2146 8628
rect 2166 8534 2170 8628
rect 2190 8534 2194 8628
rect 2214 8534 2218 8628
rect 2238 8534 2242 8628
rect 2262 8534 2266 8628
rect 2286 8534 2290 8628
rect 2310 8534 2314 8628
rect 2334 8534 2338 8628
rect 2358 8534 2362 8628
rect 2382 8534 2386 8628
rect 2406 8534 2410 8628
rect 2430 8534 2434 8628
rect 2454 8534 2458 8628
rect 2478 8534 2482 8628
rect 2502 8534 2506 8628
rect 2526 8534 2530 8628
rect 2550 8534 2554 8628
rect 2574 8534 2578 8628
rect 2598 8534 2602 8628
rect 2622 8534 2626 8628
rect 2646 8534 2650 8628
rect 2670 8534 2674 8628
rect 2694 8534 2698 8628
rect 2718 8534 2722 8628
rect 2742 8534 2746 8628
rect 2766 8534 2770 8628
rect 2790 8534 2794 8628
rect 2814 8534 2818 8628
rect 2838 8534 2842 8628
rect 2862 8534 2866 8628
rect 2886 8534 2890 8628
rect 2899 8621 2904 8628
rect 2910 8621 2914 8628
rect 2909 8607 2914 8621
rect 2899 8597 2904 8607
rect 2909 8583 2914 8597
rect 2910 8535 2914 8583
rect 2899 8534 2931 8535
rect 1213 8532 2931 8534
rect 1213 8531 1227 8532
rect 1230 8531 1237 8532
rect 1230 8510 1234 8531
rect 1254 8510 1258 8532
rect 1278 8510 1282 8532
rect 1302 8510 1306 8532
rect 1326 8510 1330 8532
rect 1350 8510 1354 8532
rect 1374 8510 1378 8532
rect 1398 8510 1402 8532
rect 1422 8510 1426 8532
rect 1446 8510 1450 8532
rect 1470 8510 1474 8532
rect 1494 8510 1498 8532
rect 1518 8510 1522 8532
rect 1542 8510 1546 8532
rect 1566 8510 1570 8532
rect 1590 8510 1594 8532
rect 1614 8510 1618 8532
rect 1638 8510 1642 8532
rect 1662 8510 1666 8532
rect 1686 8510 1690 8532
rect 1710 8510 1714 8532
rect 1734 8510 1738 8532
rect 1758 8510 1762 8532
rect 1782 8510 1786 8532
rect 1806 8510 1810 8532
rect 1830 8510 1834 8532
rect 1854 8510 1858 8532
rect 1878 8510 1882 8532
rect 1902 8510 1906 8532
rect 1926 8510 1930 8532
rect 1950 8510 1954 8532
rect 1974 8510 1978 8532
rect 1998 8510 2002 8532
rect 2022 8510 2026 8532
rect 2046 8510 2050 8532
rect 2070 8510 2074 8532
rect 2094 8510 2098 8532
rect 2118 8510 2122 8532
rect 2142 8510 2146 8532
rect 2166 8510 2170 8532
rect 2190 8510 2194 8532
rect 2214 8510 2218 8532
rect 2238 8510 2242 8532
rect 2262 8510 2266 8532
rect 2286 8510 2290 8532
rect 2310 8510 2314 8532
rect 2334 8510 2338 8532
rect 2358 8510 2362 8532
rect 2382 8510 2386 8532
rect 2406 8510 2410 8532
rect 2430 8510 2434 8532
rect 2454 8510 2458 8532
rect 2478 8510 2482 8532
rect 2502 8510 2506 8532
rect 2526 8510 2530 8532
rect 2550 8510 2554 8532
rect 2574 8510 2578 8532
rect 2598 8510 2602 8532
rect 2622 8510 2626 8532
rect 2646 8510 2650 8532
rect 2670 8510 2674 8532
rect 2694 8510 2698 8532
rect 2718 8510 2722 8532
rect 2742 8510 2746 8532
rect 2766 8510 2770 8532
rect 2790 8510 2794 8532
rect 2814 8510 2818 8532
rect 2838 8510 2842 8532
rect 2862 8510 2866 8532
rect 2886 8511 2890 8532
rect 2899 8525 2904 8532
rect 2910 8525 2914 8532
rect 2917 8531 2931 8532
rect 2909 8511 2914 8525
rect 2923 8521 2931 8525
rect 2917 8511 2923 8521
rect 2875 8510 2909 8511
rect 331 8508 2909 8510
rect 331 8501 336 8508
rect 341 8487 346 8501
rect 342 8390 346 8487
rect 366 8459 370 8508
rect 390 8483 394 8508
rect 366 8414 373 8459
rect 390 8435 397 8483
rect 390 8414 394 8435
rect 414 8414 418 8508
rect 438 8414 442 8508
rect 462 8414 466 8508
rect 486 8414 490 8508
rect 510 8414 514 8508
rect 534 8414 538 8508
rect 558 8414 562 8508
rect 582 8414 586 8508
rect 606 8414 610 8508
rect 630 8414 634 8508
rect 654 8414 658 8508
rect 678 8414 682 8508
rect 702 8414 706 8508
rect 726 8414 730 8508
rect 750 8414 754 8508
rect 774 8414 778 8508
rect 798 8414 802 8508
rect 822 8414 826 8508
rect 846 8414 850 8508
rect 870 8414 874 8508
rect 894 8414 898 8508
rect 918 8414 922 8508
rect 942 8414 946 8508
rect 966 8414 970 8508
rect 990 8414 994 8508
rect 1014 8414 1018 8508
rect 1038 8414 1042 8508
rect 1062 8414 1066 8508
rect 1086 8414 1090 8508
rect 1110 8414 1114 8508
rect 1134 8414 1138 8508
rect 1158 8414 1162 8508
rect 1182 8414 1186 8508
rect 1206 8414 1210 8508
rect 1230 8414 1234 8508
rect 1254 8414 1258 8508
rect 1278 8414 1282 8508
rect 1302 8414 1306 8508
rect 1326 8414 1330 8508
rect 1350 8414 1354 8508
rect 1374 8414 1378 8508
rect 1398 8414 1402 8508
rect 1422 8414 1426 8508
rect 1446 8414 1450 8508
rect 1470 8414 1474 8508
rect 1494 8414 1498 8508
rect 1518 8414 1522 8508
rect 1542 8414 1546 8508
rect 1566 8414 1570 8508
rect 1590 8414 1594 8508
rect 1614 8414 1618 8508
rect 1638 8414 1642 8508
rect 1662 8414 1666 8508
rect 1686 8414 1690 8508
rect 1710 8414 1714 8508
rect 1734 8414 1738 8508
rect 1758 8414 1762 8508
rect 1782 8414 1786 8508
rect 1806 8414 1810 8508
rect 1830 8414 1834 8508
rect 1854 8414 1858 8508
rect 1878 8414 1882 8508
rect 1902 8414 1906 8508
rect 1926 8414 1930 8508
rect 1950 8414 1954 8508
rect 1974 8414 1978 8508
rect 1998 8414 2002 8508
rect 2022 8414 2026 8508
rect 2046 8414 2050 8508
rect 2070 8414 2074 8508
rect 2094 8414 2098 8508
rect 2118 8414 2122 8508
rect 2142 8414 2146 8508
rect 2166 8414 2170 8508
rect 2190 8414 2194 8508
rect 2214 8414 2218 8508
rect 2238 8414 2242 8508
rect 2262 8414 2266 8508
rect 2286 8414 2290 8508
rect 2310 8414 2314 8508
rect 2334 8414 2338 8508
rect 2358 8414 2362 8508
rect 2382 8414 2386 8508
rect 2406 8414 2410 8508
rect 2430 8414 2434 8508
rect 2454 8414 2458 8508
rect 2478 8414 2482 8508
rect 2502 8414 2506 8508
rect 2526 8414 2530 8508
rect 2550 8414 2554 8508
rect 2574 8414 2578 8508
rect 2598 8414 2602 8508
rect 2622 8414 2626 8508
rect 2646 8414 2650 8508
rect 2670 8414 2674 8508
rect 2694 8414 2698 8508
rect 2718 8414 2722 8508
rect 2742 8414 2746 8508
rect 2766 8414 2770 8508
rect 2790 8414 2794 8508
rect 2814 8414 2818 8508
rect 2838 8414 2842 8508
rect 2862 8414 2866 8508
rect 2875 8501 2880 8508
rect 2886 8501 2890 8508
rect 2885 8487 2890 8501
rect 2875 8477 2880 8487
rect 2885 8463 2890 8477
rect 2886 8415 2890 8463
rect 2875 8414 2907 8415
rect 349 8412 2907 8414
rect 349 8411 363 8412
rect 366 8411 373 8412
rect 366 8390 370 8411
rect 390 8390 394 8412
rect 414 8390 418 8412
rect 438 8390 442 8412
rect 462 8390 466 8412
rect 486 8390 490 8412
rect 510 8390 514 8412
rect 534 8390 538 8412
rect 558 8390 562 8412
rect 582 8390 586 8412
rect 606 8390 610 8412
rect 630 8390 634 8412
rect 654 8390 658 8412
rect 678 8390 682 8412
rect 702 8390 706 8412
rect 726 8390 730 8412
rect 750 8390 754 8412
rect 774 8390 778 8412
rect 798 8390 802 8412
rect 822 8390 826 8412
rect 846 8390 850 8412
rect 870 8390 874 8412
rect 894 8390 898 8412
rect 918 8390 922 8412
rect 942 8390 946 8412
rect 966 8390 970 8412
rect 990 8390 994 8412
rect 1014 8390 1018 8412
rect 1038 8390 1042 8412
rect 1062 8390 1066 8412
rect 1086 8390 1090 8412
rect 1110 8390 1114 8412
rect 1134 8390 1138 8412
rect 1158 8390 1162 8412
rect 1182 8390 1186 8412
rect 1206 8390 1210 8412
rect 1230 8390 1234 8412
rect 1254 8390 1258 8412
rect 1278 8390 1282 8412
rect 1302 8390 1306 8412
rect 1326 8390 1330 8412
rect 1350 8390 1354 8412
rect 1374 8390 1378 8412
rect 1398 8390 1402 8412
rect 1422 8390 1426 8412
rect 1446 8390 1450 8412
rect 1470 8390 1474 8412
rect 1494 8390 1498 8412
rect 1518 8390 1522 8412
rect 1542 8390 1546 8412
rect 1566 8390 1570 8412
rect 1590 8390 1594 8412
rect 1614 8390 1618 8412
rect 1638 8390 1642 8412
rect 1662 8390 1666 8412
rect 1686 8390 1690 8412
rect 1710 8390 1714 8412
rect 1734 8390 1738 8412
rect 1758 8390 1762 8412
rect 1782 8390 1786 8412
rect 1806 8390 1810 8412
rect 1830 8390 1834 8412
rect 1854 8390 1858 8412
rect 1878 8390 1882 8412
rect 1902 8391 1906 8412
rect 1891 8390 1925 8391
rect -2393 8388 1925 8390
rect -2371 8366 -2366 8388
rect -2348 8366 -2343 8388
rect -2325 8366 -2320 8388
rect -2072 8386 -2036 8387
rect -2072 8380 -2054 8386
rect -2309 8372 -2301 8380
rect -2317 8366 -2309 8372
rect -2092 8371 -2062 8376
rect -2000 8367 -1992 8388
rect -1938 8387 -1906 8388
rect -1920 8386 -1906 8387
rect -1806 8380 -1680 8386
rect -1854 8371 -1806 8376
rect -1655 8372 -1647 8380
rect -1982 8367 -1966 8368
rect -2000 8366 -1966 8367
rect -1846 8366 -1806 8369
rect -1663 8366 -1655 8372
rect -1642 8366 -1637 8388
rect -1619 8366 -1614 8388
rect -1530 8366 -1526 8388
rect -1506 8366 -1502 8388
rect -1482 8366 -1478 8388
rect -1458 8366 -1454 8388
rect -1434 8366 -1430 8388
rect -1410 8366 -1406 8388
rect -1386 8366 -1382 8388
rect -1362 8366 -1358 8388
rect -1338 8366 -1334 8388
rect -1314 8366 -1310 8388
rect -1290 8366 -1286 8388
rect -1266 8366 -1262 8388
rect -1242 8366 -1238 8388
rect -1218 8366 -1214 8388
rect -1194 8366 -1190 8388
rect -1170 8366 -1166 8388
rect -1146 8366 -1142 8388
rect -1122 8366 -1118 8388
rect -1098 8366 -1094 8388
rect -1074 8366 -1070 8388
rect -1050 8366 -1046 8388
rect -1026 8366 -1022 8388
rect -1002 8366 -998 8388
rect -978 8387 -974 8388
rect -2393 8364 -981 8366
rect -2371 8342 -2366 8364
rect -2348 8342 -2343 8364
rect -2325 8342 -2320 8364
rect -2000 8362 -1966 8364
rect -2309 8344 -2301 8352
rect -2062 8351 -2054 8358
rect -2092 8344 -2084 8351
rect -2062 8344 -2026 8346
rect -2317 8342 -2309 8344
rect -2062 8342 -2012 8344
rect -2000 8342 -1992 8362
rect -1982 8361 -1966 8362
rect -1846 8360 -1806 8364
rect -1846 8353 -1798 8358
rect -1806 8351 -1798 8353
rect -1854 8349 -1846 8351
rect -1854 8344 -1806 8349
rect -1655 8344 -1647 8352
rect -1864 8342 -1796 8343
rect -1663 8342 -1655 8344
rect -1642 8342 -1637 8364
rect -1619 8342 -1614 8364
rect -1530 8342 -1526 8364
rect -1506 8342 -1502 8364
rect -1482 8342 -1478 8364
rect -1458 8342 -1454 8364
rect -1434 8342 -1430 8364
rect -1410 8342 -1406 8364
rect -1386 8342 -1382 8364
rect -1362 8342 -1358 8364
rect -1338 8342 -1334 8364
rect -1314 8342 -1310 8364
rect -1290 8342 -1286 8364
rect -1266 8342 -1262 8364
rect -1242 8342 -1238 8364
rect -1218 8342 -1214 8364
rect -1194 8342 -1190 8364
rect -1170 8342 -1166 8364
rect -1146 8342 -1142 8364
rect -1122 8342 -1118 8364
rect -1098 8342 -1094 8364
rect -1074 8342 -1070 8364
rect -1050 8342 -1046 8364
rect -1026 8342 -1022 8364
rect -1002 8342 -998 8364
rect -995 8363 -981 8364
rect -978 8363 -971 8387
rect -954 8342 -950 8388
rect -906 8363 -902 8388
rect -941 8342 -909 8343
rect -2393 8340 -909 8342
rect -2371 8294 -2366 8340
rect -2348 8294 -2343 8340
rect -2325 8294 -2320 8340
rect -2317 8336 -2309 8340
rect -2062 8336 -2054 8340
rect -2154 8332 -2138 8334
rect -2057 8332 -2054 8336
rect -2292 8326 -2054 8332
rect -2052 8326 -2044 8336
rect -2092 8310 -2062 8312
rect -2094 8306 -2062 8310
rect -2000 8294 -1992 8340
rect -1846 8333 -1806 8340
rect -1663 8336 -1655 8340
rect -1846 8326 -1680 8332
rect -1854 8310 -1806 8312
rect -1854 8306 -1680 8310
rect -1979 8294 -1945 8296
rect -1642 8294 -1637 8340
rect -1619 8294 -1614 8340
rect -1530 8294 -1526 8340
rect -1506 8294 -1502 8340
rect -1482 8294 -1478 8340
rect -1458 8294 -1454 8340
rect -1434 8294 -1430 8340
rect -1410 8294 -1406 8340
rect -1386 8294 -1382 8340
rect -1362 8294 -1358 8340
rect -1338 8294 -1334 8340
rect -1314 8294 -1310 8340
rect -1290 8294 -1286 8340
rect -1266 8294 -1262 8340
rect -1242 8294 -1238 8340
rect -1218 8294 -1214 8340
rect -1194 8294 -1190 8340
rect -1170 8294 -1166 8340
rect -1146 8294 -1142 8340
rect -1122 8294 -1118 8340
rect -1098 8294 -1094 8340
rect -1074 8294 -1070 8340
rect -1050 8294 -1046 8340
rect -1026 8294 -1022 8340
rect -1002 8294 -998 8340
rect -978 8315 -971 8339
rect -978 8294 -974 8315
rect -954 8294 -950 8340
rect -941 8333 -936 8340
rect -923 8339 -909 8340
rect -906 8339 -899 8363
rect -931 8319 -926 8333
rect -930 8294 -926 8319
rect -882 8294 -878 8388
rect -858 8294 -854 8388
rect -845 8333 -840 8343
rect -834 8333 -830 8388
rect -835 8319 -830 8333
rect -845 8318 -811 8319
rect -810 8318 -806 8388
rect -786 8318 -782 8388
rect -762 8318 -758 8388
rect -738 8318 -734 8388
rect -714 8318 -710 8388
rect -690 8318 -686 8388
rect -666 8318 -662 8388
rect -642 8318 -638 8388
rect -618 8318 -614 8388
rect -594 8318 -590 8388
rect -570 8318 -566 8388
rect -546 8318 -542 8388
rect -522 8318 -518 8388
rect -498 8318 -494 8388
rect -474 8318 -470 8388
rect -450 8318 -446 8388
rect -426 8318 -422 8388
rect -402 8318 -398 8388
rect -378 8318 -374 8388
rect -354 8318 -350 8388
rect -330 8318 -326 8388
rect -306 8318 -302 8388
rect -282 8318 -278 8388
rect -258 8318 -254 8388
rect -234 8318 -230 8388
rect -210 8318 -206 8388
rect -186 8318 -182 8388
rect -162 8318 -158 8388
rect -138 8318 -134 8388
rect -114 8318 -110 8388
rect -90 8318 -86 8388
rect -66 8318 -62 8388
rect -42 8318 -38 8388
rect -18 8318 -14 8388
rect 6 8318 10 8388
rect 30 8318 34 8388
rect 54 8318 58 8388
rect 78 8318 82 8388
rect 102 8318 106 8388
rect 126 8318 130 8388
rect 150 8318 154 8388
rect 174 8318 178 8388
rect 198 8318 202 8388
rect 222 8318 226 8388
rect 246 8318 250 8388
rect 270 8318 274 8388
rect 294 8318 298 8388
rect 318 8318 322 8388
rect 342 8318 346 8388
rect 366 8318 370 8388
rect 390 8318 394 8388
rect 414 8318 418 8388
rect 438 8318 442 8388
rect 462 8318 466 8388
rect 486 8318 490 8388
rect 510 8318 514 8388
rect 534 8318 538 8388
rect 558 8318 562 8388
rect 582 8318 586 8388
rect 606 8318 610 8388
rect 630 8318 634 8388
rect 654 8318 658 8388
rect 678 8318 682 8388
rect 702 8318 706 8388
rect 726 8318 730 8388
rect 750 8318 754 8388
rect 774 8318 778 8388
rect 798 8318 802 8388
rect 822 8318 826 8388
rect 846 8318 850 8388
rect 870 8318 874 8388
rect 894 8318 898 8388
rect 918 8318 922 8388
rect 942 8318 946 8388
rect 966 8318 970 8388
rect 990 8318 994 8388
rect 1014 8318 1018 8388
rect 1038 8318 1042 8388
rect 1062 8318 1066 8388
rect 1086 8318 1090 8388
rect 1110 8318 1114 8388
rect 1134 8318 1138 8388
rect 1158 8318 1162 8388
rect 1182 8318 1186 8388
rect 1206 8318 1210 8388
rect 1230 8318 1234 8388
rect 1254 8318 1258 8388
rect 1278 8318 1282 8388
rect 1302 8318 1306 8388
rect 1326 8318 1330 8388
rect 1350 8318 1354 8388
rect 1374 8318 1378 8388
rect 1398 8318 1402 8388
rect 1422 8318 1426 8388
rect 1446 8318 1450 8388
rect 1470 8318 1474 8388
rect 1494 8318 1498 8388
rect 1518 8318 1522 8388
rect 1542 8318 1546 8388
rect 1566 8318 1570 8388
rect 1590 8318 1594 8388
rect 1614 8318 1618 8388
rect 1638 8318 1642 8388
rect 1662 8318 1666 8388
rect 1686 8318 1690 8388
rect 1710 8318 1714 8388
rect 1734 8318 1738 8388
rect 1758 8318 1762 8388
rect 1782 8318 1786 8388
rect 1806 8318 1810 8388
rect 1830 8318 1834 8388
rect 1854 8318 1858 8388
rect 1878 8318 1882 8388
rect 1891 8381 1896 8388
rect 1902 8381 1906 8388
rect 1901 8367 1906 8381
rect 1891 8333 1896 8343
rect 1901 8319 1906 8333
rect 1902 8318 1906 8319
rect 1926 8318 1930 8412
rect 1950 8318 1954 8412
rect 1974 8318 1978 8412
rect 1998 8318 2002 8412
rect 2022 8318 2026 8412
rect 2046 8318 2050 8412
rect 2070 8318 2074 8412
rect 2094 8318 2098 8412
rect 2118 8318 2122 8412
rect 2142 8318 2146 8412
rect 2166 8318 2170 8412
rect 2179 8357 2184 8367
rect 2190 8357 2194 8412
rect 2189 8343 2194 8357
rect 2214 8318 2218 8412
rect 2238 8318 2242 8412
rect 2262 8318 2266 8412
rect 2286 8318 2290 8412
rect 2310 8318 2314 8412
rect 2334 8318 2338 8412
rect 2358 8318 2362 8412
rect 2382 8318 2386 8412
rect 2406 8318 2410 8412
rect 2430 8318 2434 8412
rect 2454 8318 2458 8412
rect 2478 8318 2482 8412
rect 2502 8318 2506 8412
rect 2526 8318 2530 8412
rect 2550 8318 2554 8412
rect 2574 8318 2578 8412
rect 2598 8318 2602 8412
rect 2622 8318 2626 8412
rect 2646 8318 2650 8412
rect 2670 8318 2674 8412
rect 2694 8318 2698 8412
rect 2718 8318 2722 8412
rect 2742 8318 2746 8412
rect 2766 8318 2770 8412
rect 2790 8318 2794 8412
rect 2814 8318 2818 8412
rect 2838 8319 2842 8412
rect 2851 8333 2856 8343
rect 2862 8333 2866 8412
rect 2875 8405 2880 8412
rect 2886 8405 2890 8412
rect 2893 8411 2907 8412
rect 2885 8391 2890 8405
rect 2899 8401 2907 8405
rect 2893 8391 2899 8401
rect 2861 8319 2866 8333
rect 2827 8318 2861 8319
rect -845 8316 2861 8318
rect -845 8309 -840 8316
rect -835 8295 -830 8309
rect -834 8294 -830 8295
rect -810 8294 -806 8316
rect -786 8294 -782 8316
rect -762 8294 -758 8316
rect -738 8294 -734 8316
rect -714 8294 -710 8316
rect -690 8294 -686 8316
rect -666 8294 -662 8316
rect -642 8294 -638 8316
rect -618 8294 -614 8316
rect -594 8294 -590 8316
rect -570 8294 -566 8316
rect -546 8294 -542 8316
rect -522 8294 -518 8316
rect -498 8294 -494 8316
rect -474 8294 -470 8316
rect -450 8294 -446 8316
rect -426 8294 -422 8316
rect -402 8294 -398 8316
rect -378 8294 -374 8316
rect -354 8294 -350 8316
rect -330 8294 -326 8316
rect -306 8294 -302 8316
rect -282 8294 -278 8316
rect -258 8294 -254 8316
rect -234 8294 -230 8316
rect -210 8294 -206 8316
rect -186 8294 -182 8316
rect -162 8294 -158 8316
rect -138 8294 -134 8316
rect -114 8294 -110 8316
rect -90 8294 -86 8316
rect -66 8294 -62 8316
rect -42 8294 -38 8316
rect -18 8294 -14 8316
rect 6 8294 10 8316
rect 30 8294 34 8316
rect 54 8294 58 8316
rect 78 8294 82 8316
rect 102 8294 106 8316
rect 126 8294 130 8316
rect 150 8294 154 8316
rect 174 8294 178 8316
rect 198 8294 202 8316
rect 222 8294 226 8316
rect 246 8294 250 8316
rect 270 8294 274 8316
rect 294 8294 298 8316
rect 318 8294 322 8316
rect 342 8294 346 8316
rect 366 8294 370 8316
rect 390 8294 394 8316
rect 414 8294 418 8316
rect 438 8294 442 8316
rect 462 8294 466 8316
rect 486 8294 490 8316
rect 510 8294 514 8316
rect 534 8294 538 8316
rect 558 8294 562 8316
rect 582 8294 586 8316
rect 606 8294 610 8316
rect 630 8294 634 8316
rect 654 8294 658 8316
rect 678 8294 682 8316
rect 702 8294 706 8316
rect 726 8294 730 8316
rect 750 8294 754 8316
rect 774 8294 778 8316
rect 798 8294 802 8316
rect 822 8294 826 8316
rect 846 8294 850 8316
rect 870 8294 874 8316
rect 894 8294 898 8316
rect 918 8294 922 8316
rect 942 8294 946 8316
rect 966 8294 970 8316
rect 990 8294 994 8316
rect 1014 8294 1018 8316
rect 1038 8294 1042 8316
rect 1062 8294 1066 8316
rect 1086 8294 1090 8316
rect 1110 8294 1114 8316
rect 1134 8294 1138 8316
rect 1158 8294 1162 8316
rect 1182 8294 1186 8316
rect 1206 8294 1210 8316
rect 1230 8294 1234 8316
rect 1254 8294 1258 8316
rect 1278 8294 1282 8316
rect 1302 8294 1306 8316
rect 1326 8294 1330 8316
rect 1350 8294 1354 8316
rect 1374 8294 1378 8316
rect 1398 8294 1402 8316
rect 1422 8294 1426 8316
rect 1446 8294 1450 8316
rect 1470 8294 1474 8316
rect 1494 8294 1498 8316
rect 1518 8294 1522 8316
rect 1542 8294 1546 8316
rect 1566 8294 1570 8316
rect 1590 8294 1594 8316
rect 1614 8294 1618 8316
rect 1638 8294 1642 8316
rect 1662 8294 1666 8316
rect 1686 8294 1690 8316
rect 1710 8294 1714 8316
rect 1734 8294 1738 8316
rect 1758 8294 1762 8316
rect 1782 8294 1786 8316
rect 1806 8294 1810 8316
rect 1830 8294 1834 8316
rect 1854 8294 1858 8316
rect 1878 8294 1882 8316
rect 1902 8294 1906 8316
rect 1926 8315 1930 8316
rect -2393 8292 1923 8294
rect -2371 8246 -2366 8292
rect -2348 8246 -2343 8292
rect -2325 8246 -2320 8292
rect -2080 8291 -1906 8292
rect -2080 8290 -2036 8291
rect -2080 8284 -2054 8290
rect -2309 8276 -2301 8282
rect -2317 8266 -2309 8276
rect -2070 8275 -2040 8282
rect -2054 8267 -2040 8270
rect -2000 8265 -1992 8291
rect -1920 8290 -1906 8291
rect -1850 8284 -1846 8292
rect -1840 8284 -1792 8292
rect -1969 8272 -1966 8281
rect -1850 8277 -1802 8282
rect -1906 8275 -1802 8277
rect -1655 8276 -1647 8282
rect -1906 8274 -1850 8275
rect -1846 8267 -1802 8273
rect -1663 8266 -1655 8276
rect -1860 8265 -1798 8266
rect -2078 8258 -2070 8265
rect -2309 8248 -2301 8254
rect -2317 8246 -2309 8248
rect -2154 8246 -2145 8256
rect -2044 8255 -2040 8260
rect -2028 8258 -1945 8265
rect -1929 8258 -1794 8265
rect -2070 8248 -2040 8255
rect -2044 8246 -2028 8248
rect -2000 8246 -1992 8258
rect -1860 8257 -1798 8258
rect -1850 8248 -1802 8255
rect -1655 8248 -1647 8254
rect -1978 8246 -1942 8247
rect -1663 8246 -1655 8248
rect -1642 8246 -1637 8292
rect -1619 8246 -1614 8292
rect -1530 8246 -1526 8292
rect -1506 8246 -1502 8292
rect -1482 8246 -1478 8292
rect -1458 8246 -1454 8292
rect -1434 8246 -1430 8292
rect -1410 8246 -1406 8292
rect -1386 8246 -1382 8292
rect -1362 8246 -1358 8292
rect -1338 8246 -1334 8292
rect -1314 8246 -1310 8292
rect -1290 8246 -1286 8292
rect -1266 8246 -1262 8292
rect -1242 8246 -1238 8292
rect -1218 8246 -1214 8292
rect -1194 8246 -1190 8292
rect -1170 8246 -1166 8292
rect -1146 8246 -1142 8292
rect -1122 8246 -1118 8292
rect -1098 8246 -1094 8292
rect -1074 8246 -1070 8292
rect -1050 8246 -1046 8292
rect -1026 8246 -1022 8292
rect -1002 8246 -998 8292
rect -978 8246 -974 8292
rect -954 8246 -950 8292
rect -930 8246 -926 8292
rect -906 8246 -899 8267
rect -882 8246 -878 8292
rect -858 8246 -854 8292
rect -834 8246 -830 8292
rect -810 8267 -806 8292
rect -2393 8244 -813 8246
rect -2371 8150 -2366 8244
rect -2348 8150 -2343 8244
rect -2325 8206 -2320 8244
rect -2317 8238 -2309 8244
rect -2145 8240 -2138 8244
rect -2070 8240 -2054 8244
rect -2078 8231 -2054 8238
rect -2062 8206 -2032 8207
rect -2000 8206 -1992 8244
rect -1846 8240 -1802 8244
rect -1846 8230 -1792 8239
rect -1663 8238 -1655 8244
rect -1942 8208 -1937 8220
rect -1850 8217 -1822 8218
rect -1850 8213 -1802 8217
rect -2325 8198 -2317 8206
rect -2062 8204 -1961 8206
rect -2325 8178 -2320 8198
rect -2317 8190 -2309 8198
rect -2062 8191 -2040 8202
rect -2032 8197 -1961 8204
rect -1947 8198 -1942 8206
rect -1842 8204 -1794 8207
rect -2070 8186 -2022 8190
rect -2325 8164 -2317 8178
rect -2072 8170 -2032 8171
rect -2102 8164 -2032 8170
rect -2325 8150 -2320 8164
rect -2317 8162 -2309 8164
rect -2309 8150 -2301 8162
rect -2070 8155 -2062 8160
rect -2000 8150 -1992 8197
rect -1942 8196 -1937 8198
rect -1932 8188 -1927 8196
rect -1912 8193 -1896 8199
rect -1842 8191 -1802 8202
rect -1671 8198 -1663 8206
rect -1663 8190 -1655 8198
rect -1850 8186 -1680 8190
rect -1924 8172 -1921 8174
rect -1806 8164 -1680 8170
rect -1671 8164 -1663 8178
rect -1663 8162 -1655 8164
rect -1854 8155 -1806 8160
rect -1974 8150 -1964 8151
rect -1960 8150 -1944 8152
rect -1842 8150 -1806 8153
rect -1655 8150 -1647 8162
rect -1642 8150 -1637 8244
rect -1619 8150 -1614 8244
rect -1530 8150 -1526 8244
rect -1506 8150 -1502 8244
rect -1482 8150 -1478 8244
rect -1458 8150 -1454 8244
rect -1434 8150 -1430 8244
rect -1410 8150 -1406 8244
rect -1386 8150 -1382 8244
rect -1362 8150 -1358 8244
rect -1338 8150 -1334 8244
rect -1314 8150 -1310 8244
rect -1290 8150 -1286 8244
rect -1266 8150 -1262 8244
rect -1242 8150 -1238 8244
rect -1218 8150 -1214 8244
rect -1194 8150 -1190 8244
rect -1170 8150 -1166 8244
rect -1146 8151 -1142 8244
rect -1157 8150 -1123 8151
rect -2393 8148 -1123 8150
rect -2371 8126 -2366 8148
rect -2348 8126 -2343 8148
rect -2325 8136 -2317 8148
rect -2325 8126 -2320 8136
rect -2317 8134 -2309 8136
rect -2062 8135 -2032 8142
rect -2309 8126 -2301 8134
rect -2070 8128 -2062 8135
rect -2000 8130 -1992 8148
rect -1974 8146 -1944 8148
rect -1960 8145 -1944 8146
rect -1842 8144 -1806 8148
rect -1842 8137 -1798 8142
rect -1806 8135 -1798 8137
rect -1671 8136 -1663 8148
rect -1854 8133 -1842 8135
rect -1663 8134 -1655 8136
rect -2062 8126 -2036 8128
rect -2393 8124 -2036 8126
rect -2032 8126 -2012 8128
rect -2004 8126 -1974 8130
rect -1854 8128 -1806 8133
rect -1864 8126 -1796 8127
rect -1655 8126 -1647 8134
rect -1642 8126 -1637 8148
rect -1619 8126 -1614 8148
rect -1530 8126 -1526 8148
rect -1506 8126 -1502 8148
rect -1482 8126 -1478 8148
rect -1458 8126 -1454 8148
rect -1434 8126 -1430 8148
rect -1410 8127 -1406 8148
rect -1421 8126 -1387 8127
rect -2032 8124 -1387 8126
rect -2371 8078 -2366 8124
rect -2348 8078 -2343 8124
rect -2325 8120 -2320 8124
rect -2309 8122 -2301 8124
rect -2317 8120 -2309 8122
rect -2325 8108 -2317 8120
rect -2052 8118 -2036 8120
rect -2052 8116 -2032 8118
rect -2062 8110 -2032 8116
rect -2325 8078 -2320 8108
rect -2317 8106 -2309 8108
rect -2092 8094 -2062 8096
rect -2094 8090 -2062 8094
rect -2000 8078 -1992 8124
rect -1904 8117 -1874 8124
rect -1842 8117 -1806 8124
rect -1655 8122 -1647 8124
rect -1663 8120 -1655 8122
rect -1842 8110 -1680 8116
rect -1671 8108 -1663 8120
rect -1663 8106 -1655 8108
rect -1854 8094 -1806 8096
rect -1854 8090 -1680 8094
rect -1642 8078 -1637 8124
rect -1619 8078 -1614 8124
rect -1530 8078 -1526 8124
rect -1506 8078 -1502 8124
rect -1482 8078 -1478 8124
rect -1458 8078 -1454 8124
rect -1434 8078 -1430 8124
rect -1421 8117 -1416 8124
rect -1410 8117 -1406 8124
rect -1411 8103 -1406 8117
rect -1410 8078 -1406 8103
rect -1386 8078 -1382 8148
rect -1362 8078 -1358 8148
rect -1338 8078 -1334 8148
rect -1314 8078 -1310 8148
rect -1290 8078 -1286 8148
rect -1266 8078 -1262 8148
rect -1242 8078 -1238 8148
rect -1218 8078 -1214 8148
rect -1194 8078 -1190 8148
rect -1170 8078 -1166 8148
rect -1157 8141 -1152 8148
rect -1146 8141 -1142 8148
rect -1147 8127 -1142 8141
rect -1157 8126 -1123 8127
rect -1122 8126 -1118 8244
rect -1098 8126 -1094 8244
rect -1074 8126 -1070 8244
rect -1050 8126 -1046 8244
rect -1026 8126 -1022 8244
rect -1002 8126 -998 8244
rect -978 8126 -974 8244
rect -954 8126 -950 8244
rect -930 8126 -926 8244
rect -923 8243 -909 8244
rect -906 8243 -899 8244
rect -906 8126 -902 8243
rect -882 8126 -878 8244
rect -858 8126 -854 8244
rect -834 8126 -830 8244
rect -827 8243 -813 8244
rect -810 8222 -803 8267
rect -786 8222 -782 8292
rect -762 8222 -758 8292
rect -738 8222 -734 8292
rect -714 8222 -710 8292
rect -690 8222 -686 8292
rect -666 8222 -662 8292
rect -642 8222 -638 8292
rect -618 8222 -614 8292
rect -594 8222 -590 8292
rect -570 8222 -566 8292
rect -546 8222 -542 8292
rect -522 8222 -518 8292
rect -509 8237 -504 8247
rect -498 8237 -494 8292
rect -499 8223 -494 8237
rect -474 8222 -470 8292
rect -450 8222 -446 8292
rect -426 8222 -422 8292
rect -402 8222 -398 8292
rect -378 8222 -374 8292
rect -354 8222 -350 8292
rect -330 8222 -326 8292
rect -306 8222 -302 8292
rect -282 8222 -278 8292
rect -258 8222 -254 8292
rect -234 8223 -230 8292
rect -245 8222 -211 8223
rect -827 8220 -211 8222
rect -827 8219 -813 8220
rect -810 8219 -803 8220
rect -810 8126 -806 8219
rect -786 8126 -782 8220
rect -762 8126 -758 8220
rect -738 8126 -734 8220
rect -714 8126 -710 8220
rect -690 8126 -686 8220
rect -666 8126 -662 8220
rect -642 8126 -638 8220
rect -618 8126 -614 8220
rect -594 8126 -590 8220
rect -570 8126 -566 8220
rect -546 8126 -542 8220
rect -522 8126 -518 8220
rect -509 8198 -475 8199
rect -474 8198 -470 8220
rect -450 8198 -446 8220
rect -426 8198 -422 8220
rect -402 8198 -398 8220
rect -378 8198 -374 8220
rect -354 8198 -350 8220
rect -330 8198 -326 8220
rect -306 8198 -302 8220
rect -282 8198 -278 8220
rect -258 8198 -254 8220
rect -245 8213 -240 8220
rect -234 8213 -230 8220
rect -235 8199 -230 8213
rect -210 8198 -206 8292
rect -186 8198 -182 8292
rect -162 8198 -158 8292
rect -138 8198 -134 8292
rect -114 8198 -110 8292
rect -90 8198 -86 8292
rect -66 8198 -62 8292
rect -42 8198 -38 8292
rect -18 8198 -14 8292
rect 6 8198 10 8292
rect 30 8198 34 8292
rect 54 8198 58 8292
rect 78 8198 82 8292
rect 102 8198 106 8292
rect 126 8198 130 8292
rect 150 8198 154 8292
rect 174 8198 178 8292
rect 198 8198 202 8292
rect 222 8198 226 8292
rect 246 8198 250 8292
rect 270 8198 274 8292
rect 294 8198 298 8292
rect 318 8198 322 8292
rect 342 8198 346 8292
rect 366 8198 370 8292
rect 390 8198 394 8292
rect 414 8198 418 8292
rect 438 8198 442 8292
rect 462 8198 466 8292
rect 486 8198 490 8292
rect 510 8198 514 8292
rect 534 8198 538 8292
rect 558 8198 562 8292
rect 582 8198 586 8292
rect 606 8198 610 8292
rect 630 8198 634 8292
rect 654 8198 658 8292
rect 678 8198 682 8292
rect 702 8198 706 8292
rect 726 8198 730 8292
rect 750 8198 754 8292
rect 774 8198 778 8292
rect 798 8198 802 8292
rect 822 8198 826 8292
rect 846 8198 850 8292
rect 870 8198 874 8292
rect 894 8198 898 8292
rect 918 8198 922 8292
rect 942 8198 946 8292
rect 966 8198 970 8292
rect 990 8198 994 8292
rect 1014 8198 1018 8292
rect 1038 8198 1042 8292
rect 1062 8198 1066 8292
rect 1086 8198 1090 8292
rect 1110 8198 1114 8292
rect 1134 8198 1138 8292
rect 1158 8198 1162 8292
rect 1182 8198 1186 8292
rect 1206 8198 1210 8292
rect 1230 8198 1234 8292
rect 1254 8198 1258 8292
rect 1278 8198 1282 8292
rect 1302 8198 1306 8292
rect 1326 8198 1330 8292
rect 1350 8198 1354 8292
rect 1374 8198 1378 8292
rect 1398 8198 1402 8292
rect 1422 8198 1426 8292
rect 1446 8198 1450 8292
rect 1470 8198 1474 8292
rect 1494 8198 1498 8292
rect 1518 8198 1522 8292
rect 1542 8198 1546 8292
rect 1566 8198 1570 8292
rect 1590 8198 1594 8292
rect 1614 8198 1618 8292
rect 1638 8198 1642 8292
rect 1662 8198 1666 8292
rect 1686 8198 1690 8292
rect 1710 8198 1714 8292
rect 1734 8198 1738 8292
rect 1758 8198 1762 8292
rect 1782 8198 1786 8292
rect 1806 8198 1810 8292
rect 1830 8198 1834 8292
rect 1854 8198 1858 8292
rect 1878 8198 1882 8292
rect 1902 8198 1906 8292
rect 1909 8291 1923 8292
rect 1926 8291 1933 8315
rect 1926 8243 1933 8267
rect 1926 8198 1930 8243
rect 1950 8198 1954 8316
rect 1974 8198 1978 8316
rect 1998 8198 2002 8316
rect 2022 8198 2026 8316
rect 2046 8198 2050 8316
rect 2070 8198 2074 8316
rect 2094 8198 2098 8316
rect 2118 8198 2122 8316
rect 2142 8198 2146 8316
rect 2166 8198 2170 8316
rect 2179 8285 2184 8295
rect 2214 8291 2218 8316
rect 2189 8271 2194 8285
rect 2203 8281 2211 8285
rect 2197 8271 2203 8281
rect 2190 8198 2194 8271
rect 2214 8267 2221 8291
rect -509 8196 2211 8198
rect -509 8189 -504 8196
rect -499 8175 -494 8189
rect -498 8126 -494 8175
rect -474 8171 -470 8196
rect -474 8147 -467 8171
rect -450 8126 -446 8196
rect -426 8126 -422 8196
rect -402 8126 -398 8196
rect -378 8126 -374 8196
rect -354 8126 -350 8196
rect -330 8126 -326 8196
rect -306 8126 -302 8196
rect -282 8126 -278 8196
rect -258 8126 -254 8196
rect -245 8165 -240 8175
rect -235 8151 -230 8165
rect -234 8126 -230 8151
rect -210 8147 -206 8196
rect -1157 8124 -213 8126
rect -1157 8117 -1152 8124
rect -1147 8103 -1142 8117
rect -1146 8078 -1142 8103
rect -1122 8078 -1118 8124
rect -1098 8078 -1094 8124
rect -1074 8078 -1070 8124
rect -1050 8078 -1046 8124
rect -1026 8078 -1022 8124
rect -1002 8078 -998 8124
rect -978 8078 -974 8124
rect -954 8078 -950 8124
rect -930 8078 -926 8124
rect -906 8078 -902 8124
rect -882 8078 -878 8124
rect -858 8078 -854 8124
rect -834 8078 -830 8124
rect -810 8078 -806 8124
rect -786 8078 -782 8124
rect -762 8078 -758 8124
rect -738 8078 -734 8124
rect -714 8078 -710 8124
rect -690 8078 -686 8124
rect -666 8078 -662 8124
rect -642 8078 -638 8124
rect -618 8078 -614 8124
rect -594 8078 -590 8124
rect -570 8078 -566 8124
rect -546 8078 -542 8124
rect -522 8078 -518 8124
rect -498 8078 -494 8124
rect -474 8099 -467 8123
rect -474 8078 -470 8099
rect -450 8078 -446 8124
rect -426 8078 -422 8124
rect -402 8078 -398 8124
rect -378 8078 -374 8124
rect -354 8078 -350 8124
rect -330 8078 -326 8124
rect -306 8078 -302 8124
rect -282 8078 -278 8124
rect -258 8078 -254 8124
rect -234 8078 -230 8124
rect -227 8123 -213 8124
rect -210 8123 -203 8147
rect -2393 8076 -213 8078
rect -2371 8054 -2366 8076
rect -2348 8054 -2343 8076
rect -2325 8054 -2320 8076
rect -2072 8074 -2036 8075
rect -2072 8068 -2054 8074
rect -2309 8060 -2301 8068
rect -2317 8054 -2309 8060
rect -2092 8059 -2062 8064
rect -2000 8055 -1992 8076
rect -1938 8075 -1906 8076
rect -1920 8074 -1906 8075
rect -1806 8068 -1680 8074
rect -1854 8059 -1806 8064
rect -1655 8060 -1647 8068
rect -1982 8055 -1966 8056
rect -2000 8054 -1966 8055
rect -1846 8054 -1806 8057
rect -1663 8054 -1655 8060
rect -1642 8054 -1637 8076
rect -1619 8054 -1614 8076
rect -1530 8054 -1526 8076
rect -1506 8054 -1502 8076
rect -1482 8054 -1478 8076
rect -1458 8054 -1454 8076
rect -1434 8054 -1430 8076
rect -1410 8054 -1406 8076
rect -1386 8054 -1382 8076
rect -1362 8054 -1358 8076
rect -1338 8054 -1334 8076
rect -1314 8054 -1310 8076
rect -1290 8054 -1286 8076
rect -1266 8054 -1262 8076
rect -1242 8054 -1238 8076
rect -1218 8054 -1214 8076
rect -1194 8054 -1190 8076
rect -1170 8054 -1166 8076
rect -1146 8054 -1142 8076
rect -1122 8075 -1118 8076
rect -2393 8052 -1125 8054
rect -2371 8030 -2366 8052
rect -2348 8030 -2343 8052
rect -2325 8030 -2320 8052
rect -2000 8050 -1966 8052
rect -2309 8032 -2301 8040
rect -2062 8039 -2054 8046
rect -2092 8032 -2084 8039
rect -2062 8032 -2026 8034
rect -2317 8030 -2309 8032
rect -2062 8030 -2012 8032
rect -2000 8030 -1992 8050
rect -1982 8049 -1966 8050
rect -1846 8048 -1806 8052
rect -1846 8041 -1798 8046
rect -1806 8039 -1798 8041
rect -1854 8037 -1846 8039
rect -1854 8032 -1806 8037
rect -1655 8032 -1647 8040
rect -1864 8030 -1796 8031
rect -1663 8030 -1655 8032
rect -1642 8030 -1637 8052
rect -1619 8030 -1614 8052
rect -1530 8030 -1526 8052
rect -1506 8031 -1502 8052
rect -1517 8030 -1483 8031
rect -2393 8028 -1483 8030
rect -2371 7982 -2366 8028
rect -2348 7982 -2343 8028
rect -2325 7982 -2320 8028
rect -2317 8024 -2309 8028
rect -2062 8024 -2054 8028
rect -2154 8020 -2138 8022
rect -2057 8020 -2054 8024
rect -2292 8014 -2054 8020
rect -2052 8014 -2044 8024
rect -2092 7998 -2062 8000
rect -2094 7994 -2062 7998
rect -2000 7982 -1992 8028
rect -1846 8021 -1806 8028
rect -1663 8024 -1655 8028
rect -1846 8014 -1680 8020
rect -1854 7998 -1806 8000
rect -1854 7994 -1680 7998
rect -1642 7982 -1637 8028
rect -1619 7982 -1614 8028
rect -1530 7982 -1526 8028
rect -1517 8021 -1512 8028
rect -1506 8021 -1502 8028
rect -1507 8007 -1502 8021
rect -1517 7997 -1512 8007
rect -1507 7983 -1502 7997
rect -1506 7982 -1502 7983
rect -1482 7982 -1478 8052
rect -1458 7982 -1454 8052
rect -1434 7982 -1430 8052
rect -1410 7982 -1406 8052
rect -1386 8051 -1382 8052
rect -1386 8027 -1379 8051
rect -1386 7982 -1382 8027
rect -1362 7982 -1358 8052
rect -1338 7982 -1334 8052
rect -1314 7982 -1310 8052
rect -1290 7982 -1286 8052
rect -1266 7982 -1262 8052
rect -1242 7982 -1238 8052
rect -1218 7982 -1214 8052
rect -1194 7982 -1190 8052
rect -1170 7982 -1166 8052
rect -1146 7982 -1142 8052
rect -1139 8051 -1125 8052
rect -1122 8027 -1115 8075
rect -1122 7982 -1118 8027
rect -1098 7982 -1094 8076
rect -1074 7982 -1070 8076
rect -1050 7982 -1046 8076
rect -1026 7982 -1022 8076
rect -1002 7982 -998 8076
rect -978 7982 -974 8076
rect -954 7982 -950 8076
rect -930 7982 -926 8076
rect -906 7982 -902 8076
rect -882 7982 -878 8076
rect -858 7982 -854 8076
rect -834 7982 -830 8076
rect -810 7982 -806 8076
rect -786 7982 -782 8076
rect -762 7982 -758 8076
rect -738 7982 -734 8076
rect -714 7982 -710 8076
rect -690 7982 -686 8076
rect -666 7982 -662 8076
rect -642 7982 -638 8076
rect -618 7982 -614 8076
rect -594 7982 -590 8076
rect -570 7982 -566 8076
rect -546 7982 -542 8076
rect -522 7982 -518 8076
rect -498 7982 -494 8076
rect -474 7982 -470 8076
rect -450 7982 -446 8076
rect -426 7982 -422 8076
rect -402 7982 -398 8076
rect -378 7982 -374 8076
rect -354 7982 -350 8076
rect -330 7982 -326 8076
rect -306 7982 -302 8076
rect -282 7982 -278 8076
rect -258 7982 -254 8076
rect -234 7982 -230 8076
rect -227 8075 -213 8076
rect -210 8075 -203 8099
rect -210 7982 -206 8075
rect -186 7982 -182 8196
rect -162 7982 -158 8196
rect -138 7982 -134 8196
rect -114 7982 -110 8196
rect -90 7982 -86 8196
rect -66 7982 -62 8196
rect -42 7982 -38 8196
rect -18 7982 -14 8196
rect 6 7982 10 8196
rect 30 7982 34 8196
rect 54 7982 58 8196
rect 78 7982 82 8196
rect 102 7982 106 8196
rect 126 7982 130 8196
rect 150 7982 154 8196
rect 174 7982 178 8196
rect 198 7982 202 8196
rect 222 7982 226 8196
rect 246 7982 250 8196
rect 270 7982 274 8196
rect 294 7982 298 8196
rect 318 7982 322 8196
rect 342 7982 346 8196
rect 366 7982 370 8196
rect 390 7982 394 8196
rect 414 7982 418 8196
rect 438 7982 442 8196
rect 462 7982 466 8196
rect 486 7982 490 8196
rect 510 7982 514 8196
rect 534 7982 538 8196
rect 558 7982 562 8196
rect 582 7982 586 8196
rect 606 7982 610 8196
rect 630 7982 634 8196
rect 654 7982 658 8196
rect 678 7982 682 8196
rect 702 7982 706 8196
rect 726 7982 730 8196
rect 750 7982 754 8196
rect 774 7982 778 8196
rect 798 7982 802 8196
rect 822 7982 826 8196
rect 846 7982 850 8196
rect 870 7982 874 8196
rect 894 7982 898 8196
rect 918 7982 922 8196
rect 942 7982 946 8196
rect 966 7982 970 8196
rect 990 7982 994 8196
rect 1014 7982 1018 8196
rect 1038 7982 1042 8196
rect 1062 7982 1066 8196
rect 1086 7982 1090 8196
rect 1110 7982 1114 8196
rect 1123 8045 1128 8055
rect 1134 8045 1138 8196
rect 1133 8031 1138 8045
rect 1123 8030 1157 8031
rect 1158 8030 1162 8196
rect 1182 8030 1186 8196
rect 1206 8030 1210 8196
rect 1230 8030 1234 8196
rect 1254 8030 1258 8196
rect 1278 8030 1282 8196
rect 1302 8030 1306 8196
rect 1326 8030 1330 8196
rect 1350 8030 1354 8196
rect 1374 8030 1378 8196
rect 1398 8030 1402 8196
rect 1422 8030 1426 8196
rect 1446 8030 1450 8196
rect 1470 8030 1474 8196
rect 1494 8030 1498 8196
rect 1518 8030 1522 8196
rect 1542 8030 1546 8196
rect 1566 8030 1570 8196
rect 1590 8030 1594 8196
rect 1614 8030 1618 8196
rect 1638 8030 1642 8196
rect 1662 8030 1666 8196
rect 1686 8030 1690 8196
rect 1710 8030 1714 8196
rect 1734 8030 1738 8196
rect 1758 8030 1762 8196
rect 1782 8030 1786 8196
rect 1806 8030 1810 8196
rect 1830 8030 1834 8196
rect 1854 8030 1858 8196
rect 1878 8030 1882 8196
rect 1902 8030 1906 8196
rect 1926 8030 1930 8196
rect 1950 8030 1954 8196
rect 1974 8030 1978 8196
rect 1998 8030 2002 8196
rect 2022 8030 2026 8196
rect 2046 8030 2050 8196
rect 2070 8030 2074 8196
rect 2094 8030 2098 8196
rect 2118 8030 2122 8196
rect 2142 8030 2146 8196
rect 2166 8030 2170 8196
rect 2190 8030 2194 8196
rect 2197 8195 2211 8196
rect 2214 8195 2221 8219
rect 2214 8030 2218 8195
rect 2238 8030 2242 8316
rect 2262 8030 2266 8316
rect 2286 8030 2290 8316
rect 2310 8030 2314 8316
rect 2334 8030 2338 8316
rect 2358 8030 2362 8316
rect 2382 8030 2386 8316
rect 2406 8030 2410 8316
rect 2430 8030 2434 8316
rect 2454 8030 2458 8316
rect 2478 8030 2482 8316
rect 2502 8030 2506 8316
rect 2526 8030 2530 8316
rect 2550 8030 2554 8316
rect 2574 8030 2578 8316
rect 2598 8030 2602 8316
rect 2622 8030 2626 8316
rect 2646 8030 2650 8316
rect 2670 8030 2674 8316
rect 2694 8030 2698 8316
rect 2718 8030 2722 8316
rect 2742 8030 2746 8316
rect 2766 8030 2770 8316
rect 2779 8117 2784 8127
rect 2790 8117 2794 8316
rect 2803 8189 2808 8199
rect 2814 8189 2818 8316
rect 2827 8309 2832 8316
rect 2838 8309 2842 8316
rect 2837 8295 2842 8309
rect 2813 8175 2818 8189
rect 2789 8103 2794 8117
rect 2779 8069 2784 8079
rect 2789 8055 2794 8069
rect 2790 8031 2794 8055
rect 2779 8030 2811 8031
rect 1123 8028 2811 8030
rect 1123 8021 1128 8028
rect 1133 8007 1138 8021
rect 1134 7982 1138 8007
rect 1158 7982 1162 8028
rect 1182 7982 1186 8028
rect 1206 7982 1210 8028
rect 1230 7982 1234 8028
rect 1254 7982 1258 8028
rect 1278 7982 1282 8028
rect 1302 7982 1306 8028
rect 1326 7982 1330 8028
rect 1350 7982 1354 8028
rect 1374 7982 1378 8028
rect 1398 7982 1402 8028
rect 1422 7982 1426 8028
rect 1446 7982 1450 8028
rect 1470 7982 1474 8028
rect 1494 7982 1498 8028
rect 1518 7982 1522 8028
rect 1542 7982 1546 8028
rect 1566 7982 1570 8028
rect 1590 7982 1594 8028
rect 1614 7982 1618 8028
rect 1638 7982 1642 8028
rect 1662 7982 1666 8028
rect 1686 7982 1690 8028
rect 1710 7982 1714 8028
rect 1734 7982 1738 8028
rect 1758 7982 1762 8028
rect 1782 7982 1786 8028
rect 1806 7982 1810 8028
rect 1830 7982 1834 8028
rect 1854 7982 1858 8028
rect 1878 7982 1882 8028
rect 1902 7982 1906 8028
rect 1926 7982 1930 8028
rect 1950 7982 1954 8028
rect 1974 7982 1978 8028
rect 1998 7982 2002 8028
rect 2022 7982 2026 8028
rect 2046 7982 2050 8028
rect 2070 7982 2074 8028
rect 2094 7982 2098 8028
rect 2118 7982 2122 8028
rect 2142 7982 2146 8028
rect 2166 7982 2170 8028
rect 2190 7982 2194 8028
rect 2214 7982 2218 8028
rect 2238 7982 2242 8028
rect 2262 7982 2266 8028
rect 2286 7982 2290 8028
rect 2310 7982 2314 8028
rect 2334 7982 2338 8028
rect 2358 7982 2362 8028
rect 2382 7982 2386 8028
rect 2406 7982 2410 8028
rect 2430 7982 2434 8028
rect 2454 7982 2458 8028
rect 2478 7982 2482 8028
rect 2502 7982 2506 8028
rect 2526 7982 2530 8028
rect 2550 7982 2554 8028
rect 2574 7982 2578 8028
rect 2598 7982 2602 8028
rect 2622 7982 2626 8028
rect 2646 7982 2650 8028
rect 2670 7982 2674 8028
rect 2694 7982 2698 8028
rect 2718 7982 2722 8028
rect 2742 7982 2746 8028
rect 2755 7997 2760 8007
rect 2766 7997 2770 8028
rect 2779 8021 2784 8028
rect 2790 8021 2794 8028
rect 2797 8027 2811 8028
rect 2789 8007 2794 8021
rect 2765 7983 2770 7997
rect 2755 7982 2789 7983
rect -2393 7980 2789 7982
rect -2371 7934 -2366 7980
rect -2348 7934 -2343 7980
rect -2325 7934 -2320 7980
rect -2309 7964 -2301 7974
rect -2317 7958 -2309 7964
rect -2097 7958 -2095 7967
rect -2309 7936 -2301 7946
rect -2097 7944 -2095 7948
rect -2292 7943 -2095 7944
rect -2097 7941 -2095 7943
rect -2084 7936 -2083 7979
rect -2069 7972 -2054 7974
rect -2054 7956 -2018 7958
rect -2054 7954 -2004 7956
rect -2059 7950 -2045 7954
rect -2054 7948 -2049 7950
rect -2317 7934 -2309 7936
rect -2084 7934 -2054 7936
rect -2044 7934 -2039 7948
rect -2025 7938 -2014 7944
rect -2000 7938 -1992 7980
rect -1920 7978 -1906 7980
rect -1977 7963 -1929 7969
rect -1655 7964 -1647 7974
rect -1977 7953 -1966 7963
rect -1663 7958 -1655 7964
rect -1977 7941 -1929 7943
rect -2033 7934 -1992 7938
rect -1655 7936 -1647 7946
rect -1663 7934 -1655 7936
rect -1642 7934 -1637 7980
rect -1619 7934 -1614 7980
rect -1530 7934 -1526 7980
rect -1506 7934 -1502 7980
rect -1482 7955 -1478 7980
rect -2393 7932 -1485 7934
rect -2371 7838 -2366 7932
rect -2348 7838 -2343 7932
rect -2325 7898 -2320 7932
rect -2317 7930 -2309 7932
rect -2084 7919 -2083 7932
rect -2084 7918 -2054 7919
rect -2325 7890 -2317 7898
rect -2325 7838 -2320 7890
rect -2317 7882 -2309 7890
rect -2117 7881 -2095 7891
rect -2045 7888 -2037 7902
rect -2309 7842 -2301 7852
rect -2087 7848 -2076 7856
rect -2017 7852 -2015 7859
rect -2317 7838 -2309 7842
rect -2092 7840 -2087 7848
rect -2092 7838 -2077 7839
rect -2000 7838 -1992 7932
rect -1663 7930 -1655 7932
rect -1969 7881 -1929 7893
rect -1671 7890 -1663 7898
rect -1663 7882 -1655 7890
rect -1655 7842 -1647 7852
rect -1928 7838 -1924 7839
rect -1854 7838 -1680 7839
rect -1663 7838 -1655 7842
rect -1642 7838 -1637 7932
rect -1619 7838 -1614 7932
rect -1530 7838 -1526 7932
rect -1506 7838 -1502 7932
rect -1499 7931 -1485 7932
rect -1482 7910 -1475 7955
rect -1458 7910 -1454 7980
rect -1434 7910 -1430 7980
rect -1410 7910 -1406 7980
rect -1386 7910 -1382 7980
rect -1362 7910 -1358 7980
rect -1338 7910 -1334 7980
rect -1314 7910 -1310 7980
rect -1290 7910 -1286 7980
rect -1266 7910 -1262 7980
rect -1242 7910 -1238 7980
rect -1218 7910 -1214 7980
rect -1194 7910 -1190 7980
rect -1170 7910 -1166 7980
rect -1146 7910 -1142 7980
rect -1122 7910 -1118 7980
rect -1098 7910 -1094 7980
rect -1074 7910 -1070 7980
rect -1050 7910 -1046 7980
rect -1026 7910 -1022 7980
rect -1002 7910 -998 7980
rect -978 7910 -974 7980
rect -954 7910 -950 7980
rect -930 7910 -926 7980
rect -906 7910 -902 7980
rect -882 7910 -878 7980
rect -858 7910 -854 7980
rect -834 7910 -830 7980
rect -810 7910 -806 7980
rect -786 7910 -782 7980
rect -762 7910 -758 7980
rect -738 7910 -734 7980
rect -714 7910 -710 7980
rect -690 7910 -686 7980
rect -666 7910 -662 7980
rect -642 7910 -638 7980
rect -618 7910 -614 7980
rect -594 7910 -590 7980
rect -570 7910 -566 7980
rect -546 7910 -542 7980
rect -522 7910 -518 7980
rect -498 7910 -494 7980
rect -474 7910 -470 7980
rect -450 7910 -446 7980
rect -426 7910 -422 7980
rect -402 7910 -398 7980
rect -378 7910 -374 7980
rect -354 7910 -350 7980
rect -330 7910 -326 7980
rect -306 7910 -302 7980
rect -282 7910 -278 7980
rect -258 7910 -254 7980
rect -234 7910 -230 7980
rect -210 7910 -206 7980
rect -186 7910 -182 7980
rect -162 7910 -158 7980
rect -138 7910 -134 7980
rect -114 7910 -110 7980
rect -90 7910 -86 7980
rect -66 7910 -62 7980
rect -42 7910 -38 7980
rect -18 7910 -14 7980
rect 6 7910 10 7980
rect 30 7910 34 7980
rect 54 7910 58 7980
rect 78 7910 82 7980
rect 102 7910 106 7980
rect 126 7910 130 7980
rect 150 7910 154 7980
rect 174 7910 178 7980
rect 198 7910 202 7980
rect 222 7910 226 7980
rect 246 7910 250 7980
rect 270 7910 274 7980
rect 294 7910 298 7980
rect 318 7910 322 7980
rect 342 7910 346 7980
rect 366 7910 370 7980
rect 390 7910 394 7980
rect 414 7910 418 7980
rect 438 7910 442 7980
rect 462 7910 466 7980
rect 475 7925 480 7935
rect 486 7925 490 7980
rect 485 7911 490 7925
rect 510 7910 514 7980
rect 534 7910 538 7980
rect 558 7910 562 7980
rect 582 7911 586 7980
rect 571 7910 605 7911
rect -1499 7908 605 7910
rect -1499 7907 -1485 7908
rect -1482 7907 -1475 7908
rect -1482 7838 -1478 7907
rect -1458 7838 -1454 7908
rect -1434 7838 -1430 7908
rect -1410 7838 -1406 7908
rect -1386 7838 -1382 7908
rect -1362 7838 -1358 7908
rect -1338 7838 -1334 7908
rect -1314 7838 -1310 7908
rect -1290 7838 -1286 7908
rect -1266 7838 -1262 7908
rect -1242 7838 -1238 7908
rect -1218 7838 -1214 7908
rect -1194 7838 -1190 7908
rect -1170 7838 -1166 7908
rect -1146 7838 -1142 7908
rect -1122 7838 -1118 7908
rect -1098 7838 -1094 7908
rect -1074 7838 -1070 7908
rect -1050 7838 -1046 7908
rect -1026 7838 -1022 7908
rect -1002 7838 -998 7908
rect -978 7838 -974 7908
rect -954 7838 -950 7908
rect -930 7838 -926 7908
rect -906 7838 -902 7908
rect -882 7838 -878 7908
rect -858 7838 -854 7908
rect -834 7838 -830 7908
rect -810 7838 -806 7908
rect -786 7838 -782 7908
rect -762 7838 -758 7908
rect -738 7838 -734 7908
rect -714 7838 -710 7908
rect -690 7838 -686 7908
rect -666 7838 -662 7908
rect -642 7838 -638 7908
rect -618 7838 -614 7908
rect -594 7838 -590 7908
rect -570 7838 -566 7908
rect -546 7838 -542 7908
rect -522 7838 -518 7908
rect -498 7838 -494 7908
rect -474 7838 -470 7908
rect -450 7838 -446 7908
rect -426 7838 -422 7908
rect -402 7838 -398 7908
rect -378 7838 -374 7908
rect -354 7838 -350 7908
rect -330 7838 -326 7908
rect -306 7838 -302 7908
rect -282 7838 -278 7908
rect -258 7838 -254 7908
rect -234 7838 -230 7908
rect -210 7838 -206 7908
rect -186 7838 -182 7908
rect -162 7838 -158 7908
rect -138 7838 -134 7908
rect -114 7838 -110 7908
rect -90 7838 -86 7908
rect -66 7838 -62 7908
rect -42 7838 -38 7908
rect -18 7838 -14 7908
rect 6 7838 10 7908
rect 30 7838 34 7908
rect 54 7838 58 7908
rect 78 7838 82 7908
rect 102 7838 106 7908
rect 126 7838 130 7908
rect 150 7838 154 7908
rect 174 7838 178 7908
rect 198 7838 202 7908
rect 222 7838 226 7908
rect 246 7838 250 7908
rect 270 7838 274 7908
rect 294 7839 298 7908
rect 283 7838 317 7839
rect -2393 7836 317 7838
rect -2371 7814 -2366 7836
rect -2348 7814 -2343 7836
rect -2325 7814 -2320 7836
rect -2092 7831 -2037 7836
rect -2021 7831 -1969 7836
rect -1921 7831 -1913 7836
rect -1854 7832 -1680 7836
rect -2100 7829 -2092 7830
rect -2309 7814 -2301 7824
rect -2100 7823 -2087 7829
rect -2051 7816 -2026 7818
rect -2062 7814 -2012 7816
rect -2000 7814 -1992 7831
rect -1969 7823 -1921 7830
rect -1969 7814 -1964 7823
rect -1864 7814 -1796 7815
rect -1655 7814 -1647 7824
rect -1642 7814 -1637 7836
rect -1619 7814 -1614 7836
rect -1530 7814 -1526 7836
rect -1506 7814 -1502 7836
rect -1482 7814 -1478 7836
rect -1458 7814 -1454 7836
rect -1434 7814 -1430 7836
rect -1410 7814 -1406 7836
rect -1386 7814 -1382 7836
rect -1362 7814 -1358 7836
rect -1338 7814 -1334 7836
rect -1314 7814 -1310 7836
rect -1290 7814 -1286 7836
rect -1266 7814 -1262 7836
rect -1242 7814 -1238 7836
rect -1218 7814 -1214 7836
rect -1194 7814 -1190 7836
rect -1170 7814 -1166 7836
rect -1146 7814 -1142 7836
rect -1122 7814 -1118 7836
rect -1098 7814 -1094 7836
rect -1074 7814 -1070 7836
rect -1050 7814 -1046 7836
rect -1026 7814 -1022 7836
rect -1002 7814 -998 7836
rect -978 7814 -974 7836
rect -954 7814 -950 7836
rect -930 7814 -926 7836
rect -906 7814 -902 7836
rect -882 7814 -878 7836
rect -858 7814 -854 7836
rect -834 7814 -830 7836
rect -810 7815 -806 7836
rect -821 7814 -787 7815
rect -2393 7812 -787 7814
rect -2371 7766 -2366 7812
rect -2348 7766 -2343 7812
rect -2325 7766 -2320 7812
rect -2317 7808 -2309 7812
rect -2105 7805 -2092 7808
rect -2092 7782 -2062 7784
rect -2094 7778 -2062 7782
rect -2000 7766 -1992 7812
rect -1663 7808 -1655 7812
rect -1969 7805 -1921 7808
rect -1854 7782 -1806 7784
rect -1854 7778 -1680 7782
rect -1926 7766 -1892 7769
rect -1642 7766 -1637 7812
rect -1619 7766 -1614 7812
rect -1530 7766 -1526 7812
rect -1506 7766 -1502 7812
rect -1482 7766 -1478 7812
rect -1458 7766 -1454 7812
rect -1434 7766 -1430 7812
rect -1410 7766 -1406 7812
rect -1386 7766 -1382 7812
rect -1362 7766 -1358 7812
rect -1338 7766 -1334 7812
rect -1314 7766 -1310 7812
rect -1290 7766 -1286 7812
rect -1266 7766 -1262 7812
rect -1242 7766 -1238 7812
rect -1218 7766 -1214 7812
rect -1194 7766 -1190 7812
rect -1170 7766 -1166 7812
rect -1146 7766 -1142 7812
rect -1122 7766 -1118 7812
rect -1098 7766 -1094 7812
rect -1074 7766 -1070 7812
rect -1050 7766 -1046 7812
rect -1026 7766 -1022 7812
rect -1002 7766 -998 7812
rect -978 7766 -974 7812
rect -954 7766 -950 7812
rect -930 7766 -926 7812
rect -906 7766 -902 7812
rect -882 7766 -878 7812
rect -858 7766 -854 7812
rect -834 7766 -830 7812
rect -821 7805 -816 7812
rect -810 7805 -806 7812
rect -811 7791 -806 7805
rect -821 7781 -816 7791
rect -811 7767 -806 7781
rect -810 7766 -806 7767
rect -786 7766 -782 7836
rect -762 7766 -758 7836
rect -738 7766 -734 7836
rect -714 7766 -710 7836
rect -690 7766 -686 7836
rect -666 7766 -662 7836
rect -642 7766 -638 7836
rect -618 7766 -614 7836
rect -594 7766 -590 7836
rect -570 7766 -566 7836
rect -546 7766 -542 7836
rect -522 7766 -518 7836
rect -498 7766 -494 7836
rect -474 7766 -470 7836
rect -450 7766 -446 7836
rect -426 7766 -422 7836
rect -402 7766 -398 7836
rect -378 7766 -374 7836
rect -354 7766 -350 7836
rect -330 7766 -326 7836
rect -306 7766 -302 7836
rect -282 7766 -278 7836
rect -258 7766 -254 7836
rect -234 7766 -230 7836
rect -210 7766 -206 7836
rect -186 7766 -182 7836
rect -162 7766 -158 7836
rect -138 7766 -134 7836
rect -114 7766 -110 7836
rect -90 7766 -86 7836
rect -66 7766 -62 7836
rect -42 7766 -38 7836
rect -18 7766 -14 7836
rect 6 7766 10 7836
rect 30 7766 34 7836
rect 54 7766 58 7836
rect 78 7766 82 7836
rect 102 7766 106 7836
rect 126 7766 130 7836
rect 150 7766 154 7836
rect 174 7766 178 7836
rect 198 7766 202 7836
rect 222 7766 226 7836
rect 246 7766 250 7836
rect 270 7766 274 7836
rect 283 7829 288 7836
rect 294 7829 298 7836
rect 293 7815 298 7829
rect 283 7814 317 7815
rect 318 7814 322 7908
rect 342 7814 346 7908
rect 366 7814 370 7908
rect 390 7814 394 7908
rect 414 7814 418 7908
rect 438 7814 442 7908
rect 462 7814 466 7908
rect 475 7886 509 7887
rect 510 7886 514 7908
rect 534 7886 538 7908
rect 558 7886 562 7908
rect 571 7901 576 7908
rect 582 7901 586 7908
rect 581 7887 586 7901
rect 606 7886 610 7980
rect 630 7886 634 7980
rect 654 7886 658 7980
rect 678 7886 682 7980
rect 702 7886 706 7980
rect 726 7886 730 7980
rect 750 7886 754 7980
rect 774 7886 778 7980
rect 798 7886 802 7980
rect 822 7886 826 7980
rect 846 7886 850 7980
rect 870 7886 874 7980
rect 894 7886 898 7980
rect 918 7886 922 7980
rect 942 7886 946 7980
rect 966 7886 970 7980
rect 990 7886 994 7980
rect 1014 7886 1018 7980
rect 1038 7886 1042 7980
rect 1062 7886 1066 7980
rect 1086 7886 1090 7980
rect 1110 7886 1114 7980
rect 1134 7886 1138 7980
rect 1158 7979 1162 7980
rect 1158 7931 1165 7979
rect 1158 7886 1162 7931
rect 1182 7886 1186 7980
rect 1206 7886 1210 7980
rect 1230 7886 1234 7980
rect 1254 7886 1258 7980
rect 1278 7886 1282 7980
rect 1302 7886 1306 7980
rect 1326 7886 1330 7980
rect 1350 7886 1354 7980
rect 1374 7886 1378 7980
rect 1398 7886 1402 7980
rect 1422 7886 1426 7980
rect 1446 7886 1450 7980
rect 1470 7886 1474 7980
rect 1494 7886 1498 7980
rect 1518 7886 1522 7980
rect 1542 7886 1546 7980
rect 1566 7886 1570 7980
rect 1590 7886 1594 7980
rect 1614 7886 1618 7980
rect 1638 7886 1642 7980
rect 1662 7886 1666 7980
rect 1686 7886 1690 7980
rect 1710 7886 1714 7980
rect 1734 7886 1738 7980
rect 1758 7886 1762 7980
rect 1782 7886 1786 7980
rect 1806 7886 1810 7980
rect 1830 7886 1834 7980
rect 1854 7886 1858 7980
rect 1878 7886 1882 7980
rect 1902 7886 1906 7980
rect 1926 7886 1930 7980
rect 1950 7886 1954 7980
rect 1974 7886 1978 7980
rect 1998 7886 2002 7980
rect 2022 7886 2026 7980
rect 2046 7886 2050 7980
rect 2070 7886 2074 7980
rect 2094 7886 2098 7980
rect 2118 7886 2122 7980
rect 2142 7886 2146 7980
rect 2166 7886 2170 7980
rect 2190 7886 2194 7980
rect 2214 7886 2218 7980
rect 2238 7886 2242 7980
rect 2262 7886 2266 7980
rect 2286 7886 2290 7980
rect 2310 7886 2314 7980
rect 2334 7886 2338 7980
rect 2358 7886 2362 7980
rect 2382 7886 2386 7980
rect 2406 7886 2410 7980
rect 2430 7886 2434 7980
rect 2454 7886 2458 7980
rect 2478 7886 2482 7980
rect 2502 7886 2506 7980
rect 2526 7886 2530 7980
rect 2550 7886 2554 7980
rect 2574 7886 2578 7980
rect 2598 7886 2602 7980
rect 2622 7886 2626 7980
rect 2646 7886 2650 7980
rect 2670 7886 2674 7980
rect 2694 7886 2698 7980
rect 2718 7886 2722 7980
rect 2742 7886 2746 7980
rect 2755 7973 2760 7980
rect 2765 7959 2770 7973
rect 2766 7887 2770 7959
rect 2755 7886 2787 7887
rect 475 7884 2787 7886
rect 475 7877 480 7884
rect 485 7863 490 7877
rect 486 7814 490 7863
rect 510 7859 514 7884
rect 510 7835 517 7859
rect 534 7814 538 7884
rect 558 7814 562 7884
rect 571 7853 576 7863
rect 581 7839 586 7853
rect 582 7814 586 7839
rect 606 7835 610 7884
rect 283 7812 603 7814
rect 283 7805 288 7812
rect 293 7791 298 7805
rect 294 7766 298 7791
rect 318 7766 322 7812
rect 342 7766 346 7812
rect 366 7766 370 7812
rect 390 7766 394 7812
rect 414 7766 418 7812
rect 438 7766 442 7812
rect 462 7766 466 7812
rect 486 7766 490 7812
rect 510 7790 517 7811
rect 534 7790 538 7812
rect 558 7790 562 7812
rect 582 7790 586 7812
rect 589 7811 603 7812
rect 606 7811 613 7835
rect 630 7790 634 7884
rect 654 7790 658 7884
rect 678 7790 682 7884
rect 702 7790 706 7884
rect 726 7790 730 7884
rect 750 7790 754 7884
rect 774 7790 778 7884
rect 798 7790 802 7884
rect 822 7790 826 7884
rect 846 7790 850 7884
rect 870 7790 874 7884
rect 894 7790 898 7884
rect 918 7790 922 7884
rect 942 7790 946 7884
rect 966 7790 970 7884
rect 990 7790 994 7884
rect 1014 7790 1018 7884
rect 1038 7790 1042 7884
rect 1062 7790 1066 7884
rect 1086 7790 1090 7884
rect 1110 7790 1114 7884
rect 1134 7790 1138 7884
rect 1158 7790 1162 7884
rect 1182 7790 1186 7884
rect 1206 7790 1210 7884
rect 1230 7790 1234 7884
rect 1254 7790 1258 7884
rect 1278 7790 1282 7884
rect 1302 7790 1306 7884
rect 1326 7790 1330 7884
rect 1350 7790 1354 7884
rect 1374 7790 1378 7884
rect 1398 7790 1402 7884
rect 1422 7790 1426 7884
rect 1446 7790 1450 7884
rect 1470 7790 1474 7884
rect 1494 7790 1498 7884
rect 1518 7790 1522 7884
rect 1542 7790 1546 7884
rect 1566 7790 1570 7884
rect 1590 7790 1594 7884
rect 1614 7790 1618 7884
rect 1638 7790 1642 7884
rect 1662 7790 1666 7884
rect 1686 7790 1690 7884
rect 1710 7790 1714 7884
rect 1734 7790 1738 7884
rect 1758 7790 1762 7884
rect 1782 7790 1786 7884
rect 1806 7790 1810 7884
rect 1830 7790 1834 7884
rect 1854 7790 1858 7884
rect 1878 7790 1882 7884
rect 1902 7790 1906 7884
rect 1926 7790 1930 7884
rect 1950 7790 1954 7884
rect 1974 7790 1978 7884
rect 1998 7790 2002 7884
rect 2022 7790 2026 7884
rect 2046 7790 2050 7884
rect 2070 7790 2074 7884
rect 2094 7790 2098 7884
rect 2118 7790 2122 7884
rect 2142 7790 2146 7884
rect 2166 7790 2170 7884
rect 2190 7790 2194 7884
rect 2214 7790 2218 7884
rect 2238 7790 2242 7884
rect 2262 7790 2266 7884
rect 2286 7790 2290 7884
rect 2310 7790 2314 7884
rect 2334 7790 2338 7884
rect 2358 7790 2362 7884
rect 2382 7790 2386 7884
rect 2406 7790 2410 7884
rect 2430 7790 2434 7884
rect 2454 7790 2458 7884
rect 2478 7790 2482 7884
rect 2502 7790 2506 7884
rect 2526 7790 2530 7884
rect 2550 7790 2554 7884
rect 2574 7790 2578 7884
rect 2598 7790 2602 7884
rect 2622 7790 2626 7884
rect 2646 7790 2650 7884
rect 2670 7790 2674 7884
rect 2694 7790 2698 7884
rect 2718 7791 2722 7884
rect 2731 7805 2736 7815
rect 2742 7805 2746 7884
rect 2755 7877 2760 7884
rect 2766 7877 2770 7884
rect 2773 7883 2787 7884
rect 2765 7863 2770 7877
rect 2741 7791 2746 7805
rect 2707 7790 2741 7791
rect 493 7788 2741 7790
rect 493 7787 507 7788
rect 510 7787 517 7788
rect 510 7766 514 7787
rect 534 7766 538 7788
rect 558 7766 562 7788
rect 582 7766 586 7788
rect -2393 7764 603 7766
rect -2371 7742 -2366 7764
rect -2348 7742 -2343 7764
rect -2325 7742 -2320 7764
rect -2054 7763 -1906 7764
rect -2054 7762 -2036 7763
rect -2309 7748 -2301 7758
rect -2317 7742 -2309 7748
rect -2068 7747 -2038 7754
rect -2000 7746 -1992 7763
rect -1920 7762 -1906 7763
rect -1846 7756 -1794 7764
rect -1852 7749 -1804 7754
rect -1902 7747 -1804 7749
rect -1655 7748 -1647 7758
rect -2000 7744 -1975 7746
rect -1902 7745 -1852 7747
rect -2025 7742 -1975 7744
rect -1846 7742 -1804 7745
rect -1663 7742 -1655 7748
rect -1642 7742 -1637 7764
rect -1619 7742 -1614 7764
rect -1530 7742 -1526 7764
rect -1506 7742 -1502 7764
rect -1482 7742 -1478 7764
rect -1458 7742 -1454 7764
rect -1434 7742 -1430 7764
rect -1410 7742 -1406 7764
rect -1386 7742 -1382 7764
rect -1362 7742 -1358 7764
rect -1338 7742 -1334 7764
rect -1314 7742 -1310 7764
rect -1290 7742 -1286 7764
rect -1266 7742 -1262 7764
rect -1242 7742 -1238 7764
rect -1218 7742 -1214 7764
rect -1194 7742 -1190 7764
rect -1170 7742 -1166 7764
rect -1146 7742 -1142 7764
rect -1122 7742 -1118 7764
rect -1098 7742 -1094 7764
rect -1074 7742 -1070 7764
rect -1050 7742 -1046 7764
rect -1026 7742 -1022 7764
rect -1002 7742 -998 7764
rect -978 7742 -974 7764
rect -954 7742 -950 7764
rect -930 7742 -926 7764
rect -906 7742 -902 7764
rect -882 7742 -878 7764
rect -858 7742 -854 7764
rect -834 7742 -830 7764
rect -810 7742 -806 7764
rect -786 7742 -782 7764
rect -762 7742 -758 7764
rect -738 7742 -734 7764
rect -714 7742 -710 7764
rect -690 7742 -686 7764
rect -666 7742 -662 7764
rect -642 7742 -638 7764
rect -618 7742 -614 7764
rect -594 7742 -590 7764
rect -570 7742 -566 7764
rect -546 7742 -542 7764
rect -522 7742 -518 7764
rect -498 7742 -494 7764
rect -474 7742 -470 7764
rect -450 7742 -446 7764
rect -426 7742 -422 7764
rect -402 7742 -398 7764
rect -378 7742 -374 7764
rect -354 7742 -350 7764
rect -330 7742 -326 7764
rect -306 7742 -302 7764
rect -282 7742 -278 7764
rect -258 7742 -254 7764
rect -234 7742 -230 7764
rect -210 7742 -206 7764
rect -186 7742 -182 7764
rect -162 7742 -158 7764
rect -138 7742 -134 7764
rect -114 7742 -110 7764
rect -90 7742 -86 7764
rect -66 7742 -62 7764
rect -42 7742 -38 7764
rect -18 7742 -14 7764
rect 6 7742 10 7764
rect 30 7742 34 7764
rect 54 7742 58 7764
rect 78 7742 82 7764
rect 102 7742 106 7764
rect 126 7742 130 7764
rect 150 7742 154 7764
rect 174 7742 178 7764
rect 198 7742 202 7764
rect 222 7742 226 7764
rect 246 7742 250 7764
rect 270 7742 274 7764
rect 294 7742 298 7764
rect 318 7763 322 7764
rect -2393 7740 315 7742
rect -2371 7718 -2366 7740
rect -2348 7718 -2343 7740
rect -2325 7718 -2320 7740
rect -2054 7739 -2038 7740
rect -2000 7739 -1966 7740
rect -1846 7739 -1804 7740
rect -2000 7738 -1975 7739
rect -2076 7730 -2054 7737
rect -2309 7720 -2301 7730
rect -2044 7727 -2038 7732
rect -2028 7730 -2001 7737
rect -2054 7720 -2038 7727
rect -2015 7729 -2001 7730
rect -2015 7720 -2014 7729
rect -2317 7718 -2309 7720
rect -2044 7718 -2028 7720
rect -2000 7718 -1992 7738
rect -1982 7737 -1975 7738
rect -1862 7737 -1798 7738
rect -1985 7730 -1796 7737
rect -1862 7729 -1798 7730
rect -1852 7720 -1804 7727
rect -1655 7720 -1647 7730
rect -1976 7718 -1940 7719
rect -1663 7718 -1655 7720
rect -1642 7718 -1637 7740
rect -1619 7718 -1614 7740
rect -1530 7718 -1526 7740
rect -1506 7718 -1502 7740
rect -1482 7718 -1478 7740
rect -1458 7718 -1454 7740
rect -1434 7718 -1430 7740
rect -1410 7718 -1406 7740
rect -1386 7718 -1382 7740
rect -1362 7718 -1358 7740
rect -1338 7718 -1334 7740
rect -1314 7718 -1310 7740
rect -1290 7718 -1286 7740
rect -1266 7718 -1262 7740
rect -1242 7718 -1238 7740
rect -1218 7718 -1214 7740
rect -1194 7718 -1190 7740
rect -1170 7718 -1166 7740
rect -1146 7718 -1142 7740
rect -1122 7718 -1118 7740
rect -1098 7718 -1094 7740
rect -1074 7718 -1070 7740
rect -1050 7718 -1046 7740
rect -1026 7718 -1022 7740
rect -1002 7718 -998 7740
rect -978 7718 -974 7740
rect -954 7718 -950 7740
rect -930 7718 -926 7740
rect -906 7718 -902 7740
rect -882 7718 -878 7740
rect -858 7718 -854 7740
rect -834 7718 -830 7740
rect -810 7718 -806 7740
rect -786 7739 -782 7740
rect -2393 7716 -789 7718
rect -2371 7646 -2366 7716
rect -2348 7646 -2343 7716
rect -2325 7682 -2320 7716
rect -2317 7714 -2309 7716
rect -2076 7703 -2054 7710
rect -2325 7674 -2317 7682
rect -2060 7676 -2030 7679
rect -2325 7654 -2320 7674
rect -2317 7666 -2309 7674
rect -2060 7663 -2038 7674
rect -2033 7667 -2030 7676
rect -2028 7672 -2027 7676
rect -2068 7658 -2038 7661
rect -2325 7646 -2317 7654
rect -2000 7646 -1992 7716
rect -1846 7712 -1804 7716
rect -1663 7714 -1655 7716
rect -1846 7702 -1794 7711
rect -1912 7691 -1884 7693
rect -1852 7685 -1804 7689
rect -1844 7676 -1796 7679
rect -1671 7674 -1663 7682
rect -1844 7663 -1804 7674
rect -1663 7666 -1655 7674
rect -1852 7658 -1680 7662
rect -1926 7646 -1892 7649
rect -1671 7646 -1663 7654
rect -1642 7646 -1637 7716
rect -1619 7646 -1614 7716
rect -1530 7646 -1526 7716
rect -1506 7646 -1502 7716
rect -1482 7646 -1478 7716
rect -1458 7646 -1454 7716
rect -1434 7646 -1430 7716
rect -1410 7646 -1406 7716
rect -1386 7646 -1382 7716
rect -1362 7646 -1358 7716
rect -1338 7646 -1334 7716
rect -1314 7646 -1310 7716
rect -1290 7646 -1286 7716
rect -1266 7646 -1262 7716
rect -1242 7646 -1238 7716
rect -1218 7646 -1214 7716
rect -1194 7646 -1190 7716
rect -1170 7646 -1166 7716
rect -1146 7646 -1142 7716
rect -1122 7646 -1118 7716
rect -1098 7646 -1094 7716
rect -1074 7646 -1070 7716
rect -1050 7646 -1046 7716
rect -1026 7646 -1022 7716
rect -1002 7646 -998 7716
rect -978 7646 -974 7716
rect -954 7646 -950 7716
rect -930 7646 -926 7716
rect -906 7646 -902 7716
rect -882 7646 -878 7716
rect -858 7646 -854 7716
rect -834 7646 -830 7716
rect -810 7646 -806 7716
rect -803 7715 -789 7716
rect -786 7694 -779 7739
rect -762 7694 -758 7740
rect -738 7694 -734 7740
rect -714 7694 -710 7740
rect -690 7694 -686 7740
rect -666 7694 -662 7740
rect -642 7694 -638 7740
rect -618 7694 -614 7740
rect -594 7694 -590 7740
rect -570 7694 -566 7740
rect -546 7694 -542 7740
rect -522 7694 -518 7740
rect -498 7694 -494 7740
rect -474 7694 -470 7740
rect -450 7694 -446 7740
rect -426 7694 -422 7740
rect -402 7694 -398 7740
rect -378 7694 -374 7740
rect -354 7694 -350 7740
rect -330 7694 -326 7740
rect -306 7694 -302 7740
rect -282 7694 -278 7740
rect -258 7694 -254 7740
rect -234 7694 -230 7740
rect -210 7694 -206 7740
rect -186 7694 -182 7740
rect -162 7695 -158 7740
rect -173 7694 -139 7695
rect -803 7692 -139 7694
rect -803 7691 -789 7692
rect -786 7691 -779 7692
rect -786 7646 -782 7691
rect -762 7646 -758 7692
rect -738 7646 -734 7692
rect -714 7646 -710 7692
rect -690 7646 -686 7692
rect -666 7646 -662 7692
rect -642 7646 -638 7692
rect -618 7646 -614 7692
rect -594 7646 -590 7692
rect -570 7646 -566 7692
rect -546 7646 -542 7692
rect -522 7646 -518 7692
rect -498 7646 -494 7692
rect -474 7646 -470 7692
rect -450 7646 -446 7692
rect -426 7646 -422 7692
rect -402 7646 -398 7692
rect -378 7646 -374 7692
rect -354 7646 -350 7692
rect -330 7646 -326 7692
rect -306 7646 -302 7692
rect -282 7646 -278 7692
rect -258 7646 -254 7692
rect -234 7646 -230 7692
rect -210 7646 -206 7692
rect -186 7646 -182 7692
rect -173 7685 -168 7692
rect -162 7685 -158 7692
rect -163 7671 -158 7685
rect -173 7670 -139 7671
rect -138 7670 -134 7740
rect -114 7670 -110 7740
rect -90 7670 -86 7740
rect -66 7670 -62 7740
rect -42 7670 -38 7740
rect -18 7670 -14 7740
rect 6 7670 10 7740
rect 30 7670 34 7740
rect 54 7670 58 7740
rect 78 7670 82 7740
rect 102 7670 106 7740
rect 126 7670 130 7740
rect 150 7670 154 7740
rect 174 7670 178 7740
rect 198 7670 202 7740
rect 222 7670 226 7740
rect 246 7670 250 7740
rect 270 7670 274 7740
rect 294 7670 298 7740
rect 301 7739 315 7740
rect 318 7718 325 7763
rect 342 7718 346 7764
rect 366 7718 370 7764
rect 390 7718 394 7764
rect 414 7718 418 7764
rect 438 7718 442 7764
rect 462 7718 466 7764
rect 486 7718 490 7764
rect 510 7718 514 7764
rect 534 7718 538 7764
rect 558 7718 562 7764
rect 582 7718 586 7764
rect 589 7763 603 7764
rect 606 7763 613 7787
rect 606 7718 610 7763
rect 630 7718 634 7788
rect 654 7718 658 7788
rect 678 7718 682 7788
rect 702 7718 706 7788
rect 726 7718 730 7788
rect 750 7718 754 7788
rect 774 7718 778 7788
rect 798 7718 802 7788
rect 822 7718 826 7788
rect 846 7718 850 7788
rect 870 7718 874 7788
rect 894 7718 898 7788
rect 918 7718 922 7788
rect 942 7718 946 7788
rect 966 7718 970 7788
rect 990 7718 994 7788
rect 1014 7718 1018 7788
rect 1038 7718 1042 7788
rect 1062 7718 1066 7788
rect 1086 7718 1090 7788
rect 1110 7718 1114 7788
rect 1134 7718 1138 7788
rect 1158 7718 1162 7788
rect 1182 7718 1186 7788
rect 1206 7718 1210 7788
rect 1230 7718 1234 7788
rect 1254 7718 1258 7788
rect 1278 7718 1282 7788
rect 1302 7718 1306 7788
rect 1326 7718 1330 7788
rect 1350 7718 1354 7788
rect 1374 7718 1378 7788
rect 1398 7718 1402 7788
rect 1422 7718 1426 7788
rect 1446 7718 1450 7788
rect 1470 7718 1474 7788
rect 1494 7718 1498 7788
rect 1518 7718 1522 7788
rect 1542 7718 1546 7788
rect 1566 7718 1570 7788
rect 1590 7718 1594 7788
rect 1614 7718 1618 7788
rect 1638 7718 1642 7788
rect 1662 7718 1666 7788
rect 1686 7718 1690 7788
rect 1710 7718 1714 7788
rect 1734 7718 1738 7788
rect 1758 7718 1762 7788
rect 1782 7718 1786 7788
rect 1806 7718 1810 7788
rect 1830 7718 1834 7788
rect 1854 7718 1858 7788
rect 1878 7718 1882 7788
rect 1902 7718 1906 7788
rect 1926 7718 1930 7788
rect 1950 7718 1954 7788
rect 1974 7718 1978 7788
rect 1998 7719 2002 7788
rect 1987 7718 2021 7719
rect 301 7716 2021 7718
rect 301 7715 315 7716
rect 318 7715 325 7716
rect 318 7670 322 7715
rect 342 7670 346 7716
rect 366 7670 370 7716
rect 390 7670 394 7716
rect 414 7670 418 7716
rect 438 7670 442 7716
rect 462 7670 466 7716
rect 486 7670 490 7716
rect 510 7670 514 7716
rect 534 7670 538 7716
rect 558 7670 562 7716
rect 582 7670 586 7716
rect 606 7670 610 7716
rect 630 7670 634 7716
rect 654 7670 658 7716
rect 678 7670 682 7716
rect 702 7670 706 7716
rect 726 7670 730 7716
rect 750 7670 754 7716
rect 774 7670 778 7716
rect 798 7670 802 7716
rect 822 7670 826 7716
rect 846 7670 850 7716
rect 870 7670 874 7716
rect 894 7670 898 7716
rect 918 7670 922 7716
rect 942 7670 946 7716
rect 966 7670 970 7716
rect 990 7670 994 7716
rect 1014 7670 1018 7716
rect 1038 7670 1042 7716
rect 1062 7670 1066 7716
rect 1086 7670 1090 7716
rect 1110 7670 1114 7716
rect 1134 7670 1138 7716
rect 1158 7670 1162 7716
rect 1182 7670 1186 7716
rect 1206 7670 1210 7716
rect 1230 7670 1234 7716
rect 1254 7670 1258 7716
rect 1278 7670 1282 7716
rect 1302 7670 1306 7716
rect 1326 7670 1330 7716
rect 1350 7670 1354 7716
rect 1374 7670 1378 7716
rect 1398 7670 1402 7716
rect 1422 7670 1426 7716
rect 1446 7670 1450 7716
rect 1470 7670 1474 7716
rect 1494 7670 1498 7716
rect 1518 7670 1522 7716
rect 1542 7670 1546 7716
rect 1566 7670 1570 7716
rect 1590 7670 1594 7716
rect 1614 7670 1618 7716
rect 1638 7670 1642 7716
rect 1662 7670 1666 7716
rect 1686 7670 1690 7716
rect 1710 7670 1714 7716
rect 1734 7670 1738 7716
rect 1758 7670 1762 7716
rect 1782 7670 1786 7716
rect 1806 7670 1810 7716
rect 1830 7670 1834 7716
rect 1854 7670 1858 7716
rect 1878 7670 1882 7716
rect 1902 7670 1906 7716
rect 1926 7670 1930 7716
rect 1950 7670 1954 7716
rect 1974 7670 1978 7716
rect 1987 7709 1992 7716
rect 1998 7709 2002 7716
rect 1997 7695 2002 7709
rect 1987 7694 2021 7695
rect 2022 7694 2026 7788
rect 2046 7694 2050 7788
rect 2070 7694 2074 7788
rect 2094 7694 2098 7788
rect 2118 7694 2122 7788
rect 2142 7694 2146 7788
rect 2155 7733 2160 7743
rect 2166 7733 2170 7788
rect 2165 7719 2170 7733
rect 2155 7718 2189 7719
rect 2190 7718 2194 7788
rect 2214 7718 2218 7788
rect 2238 7718 2242 7788
rect 2262 7718 2266 7788
rect 2286 7718 2290 7788
rect 2310 7718 2314 7788
rect 2334 7718 2338 7788
rect 2358 7718 2362 7788
rect 2382 7718 2386 7788
rect 2406 7718 2410 7788
rect 2430 7718 2434 7788
rect 2454 7718 2458 7788
rect 2478 7718 2482 7788
rect 2502 7718 2506 7788
rect 2526 7718 2530 7788
rect 2550 7718 2554 7788
rect 2574 7718 2578 7788
rect 2598 7718 2602 7788
rect 2622 7718 2626 7788
rect 2646 7718 2650 7788
rect 2670 7718 2674 7788
rect 2694 7718 2698 7788
rect 2707 7781 2712 7788
rect 2718 7781 2722 7788
rect 2717 7767 2722 7781
rect 2707 7757 2712 7767
rect 2717 7743 2722 7757
rect 2718 7719 2722 7743
rect 2707 7718 2741 7719
rect 2155 7716 2741 7718
rect 2155 7709 2160 7716
rect 2165 7695 2170 7709
rect 2166 7694 2170 7695
rect 2190 7694 2194 7716
rect 2214 7694 2218 7716
rect 2238 7694 2242 7716
rect 2262 7694 2266 7716
rect 2286 7694 2290 7716
rect 2310 7694 2314 7716
rect 2334 7694 2338 7716
rect 2358 7694 2362 7716
rect 2382 7694 2386 7716
rect 2406 7694 2410 7716
rect 2430 7694 2434 7716
rect 2454 7694 2458 7716
rect 2478 7694 2482 7716
rect 2502 7694 2506 7716
rect 2526 7694 2530 7716
rect 2550 7694 2554 7716
rect 2574 7694 2578 7716
rect 2598 7694 2602 7716
rect 2622 7694 2626 7716
rect 2646 7694 2650 7716
rect 2670 7694 2674 7716
rect 2694 7695 2698 7716
rect 2707 7709 2712 7716
rect 2718 7709 2722 7716
rect 2717 7695 2722 7709
rect 2731 7705 2739 7709
rect 2725 7695 2731 7705
rect 2683 7694 2717 7695
rect 1987 7692 2717 7694
rect 1987 7685 1992 7692
rect 1997 7671 2002 7685
rect 1998 7670 2002 7671
rect 2022 7670 2026 7692
rect 2046 7670 2050 7692
rect 2070 7670 2074 7692
rect 2094 7670 2098 7692
rect 2118 7670 2122 7692
rect 2142 7670 2146 7692
rect 2166 7670 2170 7692
rect 2190 7670 2194 7692
rect 2214 7670 2218 7692
rect 2238 7670 2242 7692
rect 2262 7670 2266 7692
rect 2286 7670 2290 7692
rect 2310 7670 2314 7692
rect 2334 7670 2338 7692
rect 2358 7670 2362 7692
rect 2382 7670 2386 7692
rect 2406 7670 2410 7692
rect 2430 7670 2434 7692
rect 2454 7670 2458 7692
rect 2478 7670 2482 7692
rect 2502 7670 2506 7692
rect 2526 7670 2530 7692
rect 2550 7670 2554 7692
rect 2574 7670 2578 7692
rect 2598 7670 2602 7692
rect 2622 7670 2626 7692
rect 2646 7670 2650 7692
rect 2670 7671 2674 7692
rect 2683 7685 2688 7692
rect 2694 7685 2698 7692
rect 2693 7671 2698 7685
rect 2659 7670 2693 7671
rect -173 7668 2693 7670
rect -173 7661 -168 7668
rect -163 7647 -158 7661
rect -162 7646 -158 7647
rect -138 7646 -134 7668
rect -114 7646 -110 7668
rect -90 7646 -86 7668
rect -66 7646 -62 7668
rect -42 7646 -38 7668
rect -18 7646 -14 7668
rect 6 7646 10 7668
rect 30 7646 34 7668
rect 54 7646 58 7668
rect 78 7646 82 7668
rect 102 7646 106 7668
rect 126 7646 130 7668
rect 150 7646 154 7668
rect 174 7646 178 7668
rect 198 7646 202 7668
rect 222 7646 226 7668
rect 246 7646 250 7668
rect 270 7646 274 7668
rect 294 7646 298 7668
rect 318 7646 322 7668
rect 342 7646 346 7668
rect 366 7646 370 7668
rect 390 7646 394 7668
rect 414 7646 418 7668
rect 438 7646 442 7668
rect 462 7646 466 7668
rect 486 7646 490 7668
rect 510 7646 514 7668
rect 534 7646 538 7668
rect 558 7646 562 7668
rect 582 7646 586 7668
rect 606 7646 610 7668
rect 630 7646 634 7668
rect 654 7646 658 7668
rect 678 7646 682 7668
rect 702 7646 706 7668
rect 726 7646 730 7668
rect 750 7646 754 7668
rect 774 7646 778 7668
rect 798 7646 802 7668
rect 822 7646 826 7668
rect 846 7646 850 7668
rect 870 7646 874 7668
rect 894 7646 898 7668
rect 918 7646 922 7668
rect 942 7646 946 7668
rect 966 7646 970 7668
rect 990 7646 994 7668
rect 1014 7646 1018 7668
rect 1038 7646 1042 7668
rect 1062 7646 1066 7668
rect 1086 7646 1090 7668
rect 1110 7646 1114 7668
rect 1134 7646 1138 7668
rect 1158 7646 1162 7668
rect 1182 7646 1186 7668
rect 1206 7646 1210 7668
rect 1230 7646 1234 7668
rect 1254 7646 1258 7668
rect 1278 7646 1282 7668
rect 1302 7646 1306 7668
rect 1326 7646 1330 7668
rect 1350 7646 1354 7668
rect 1374 7646 1378 7668
rect 1398 7646 1402 7668
rect 1422 7646 1426 7668
rect 1446 7646 1450 7668
rect 1470 7646 1474 7668
rect 1494 7646 1498 7668
rect 1518 7646 1522 7668
rect 1542 7646 1546 7668
rect 1566 7646 1570 7668
rect 1590 7646 1594 7668
rect 1614 7646 1618 7668
rect 1638 7646 1642 7668
rect 1662 7646 1666 7668
rect 1686 7646 1690 7668
rect 1710 7646 1714 7668
rect 1734 7646 1738 7668
rect 1758 7646 1762 7668
rect 1782 7646 1786 7668
rect 1806 7646 1810 7668
rect 1830 7646 1834 7668
rect 1854 7646 1858 7668
rect 1878 7646 1882 7668
rect 1902 7646 1906 7668
rect 1926 7646 1930 7668
rect 1950 7646 1954 7668
rect 1974 7646 1978 7668
rect 1998 7646 2002 7668
rect 2022 7646 2026 7668
rect 2046 7646 2050 7668
rect 2070 7646 2074 7668
rect 2094 7646 2098 7668
rect 2118 7646 2122 7668
rect 2142 7646 2146 7668
rect 2166 7646 2170 7668
rect 2190 7667 2194 7668
rect -2393 7644 2187 7646
rect -2371 7622 -2366 7644
rect -2348 7622 -2343 7644
rect -2325 7638 -2317 7644
rect -2325 7622 -2320 7638
rect -2309 7626 -2301 7638
rect -2068 7627 -2038 7634
rect -2317 7622 -2309 7626
rect -2000 7624 -1992 7644
rect -1844 7636 -1794 7644
rect -1671 7638 -1663 7644
rect -1852 7627 -1804 7634
rect -1655 7626 -1647 7638
rect -2025 7623 -1991 7624
rect -2025 7622 -1975 7623
rect -1844 7622 -1804 7625
rect -1663 7622 -1655 7626
rect -1642 7622 -1637 7644
rect -1619 7622 -1614 7644
rect -1530 7622 -1526 7644
rect -1506 7622 -1502 7644
rect -1482 7622 -1478 7644
rect -1458 7622 -1454 7644
rect -1434 7622 -1430 7644
rect -1410 7622 -1406 7644
rect -1386 7622 -1382 7644
rect -1362 7622 -1358 7644
rect -1338 7622 -1334 7644
rect -1314 7622 -1310 7644
rect -1290 7622 -1286 7644
rect -1266 7622 -1262 7644
rect -1242 7622 -1238 7644
rect -1218 7622 -1214 7644
rect -1194 7622 -1190 7644
rect -1170 7622 -1166 7644
rect -1146 7622 -1142 7644
rect -1122 7622 -1118 7644
rect -1098 7622 -1094 7644
rect -1074 7622 -1070 7644
rect -1050 7622 -1046 7644
rect -1026 7622 -1022 7644
rect -1002 7622 -998 7644
rect -978 7622 -974 7644
rect -954 7622 -950 7644
rect -930 7622 -926 7644
rect -906 7622 -902 7644
rect -882 7622 -878 7644
rect -858 7622 -854 7644
rect -834 7622 -830 7644
rect -810 7622 -806 7644
rect -786 7622 -782 7644
rect -762 7622 -758 7644
rect -738 7622 -734 7644
rect -714 7622 -710 7644
rect -690 7622 -686 7644
rect -666 7622 -662 7644
rect -642 7622 -638 7644
rect -618 7622 -614 7644
rect -594 7622 -590 7644
rect -570 7622 -566 7644
rect -546 7622 -542 7644
rect -522 7622 -518 7644
rect -498 7622 -494 7644
rect -474 7622 -470 7644
rect -450 7622 -446 7644
rect -426 7622 -422 7644
rect -402 7622 -398 7644
rect -378 7622 -374 7644
rect -354 7622 -350 7644
rect -330 7622 -326 7644
rect -306 7622 -302 7644
rect -282 7622 -278 7644
rect -258 7622 -254 7644
rect -234 7622 -230 7644
rect -210 7622 -206 7644
rect -186 7622 -182 7644
rect -162 7622 -158 7644
rect -138 7622 -134 7644
rect -114 7622 -110 7644
rect -90 7622 -86 7644
rect -66 7622 -62 7644
rect -42 7622 -38 7644
rect -18 7622 -14 7644
rect 6 7622 10 7644
rect 30 7622 34 7644
rect 54 7622 58 7644
rect 78 7622 82 7644
rect 102 7622 106 7644
rect 126 7622 130 7644
rect 150 7622 154 7644
rect 174 7623 178 7644
rect 163 7622 197 7623
rect -2393 7620 197 7622
rect -2371 7598 -2366 7620
rect -2348 7598 -2343 7620
rect -2325 7610 -2317 7620
rect -2060 7610 -2020 7617
rect -2004 7612 -2001 7617
rect -2015 7610 -2001 7612
rect -2000 7610 -1992 7620
rect -1972 7618 -1958 7620
rect -1844 7619 -1804 7620
rect -1862 7617 -1796 7618
rect -1985 7615 -1796 7617
rect -1985 7610 -1852 7615
rect -2325 7598 -2320 7610
rect -2309 7598 -2301 7610
rect -2068 7600 -2060 7607
rect -2015 7600 -1990 7610
rect -1844 7609 -1796 7615
rect -1671 7610 -1663 7620
rect -1852 7600 -1804 7607
rect -2020 7598 -2004 7600
rect -2000 7598 -1992 7600
rect -1976 7598 -1940 7599
rect -1655 7598 -1647 7610
rect -1642 7598 -1637 7620
rect -1619 7598 -1614 7620
rect -1530 7598 -1526 7620
rect -1506 7598 -1502 7620
rect -1482 7598 -1478 7620
rect -1458 7598 -1454 7620
rect -1434 7598 -1430 7620
rect -1410 7598 -1406 7620
rect -1386 7598 -1382 7620
rect -1362 7598 -1358 7620
rect -1338 7598 -1334 7620
rect -1314 7598 -1310 7620
rect -1290 7598 -1286 7620
rect -1266 7598 -1262 7620
rect -1242 7598 -1238 7620
rect -1218 7598 -1214 7620
rect -1194 7598 -1190 7620
rect -1170 7598 -1166 7620
rect -1146 7598 -1142 7620
rect -1122 7598 -1118 7620
rect -1098 7598 -1094 7620
rect -1074 7598 -1070 7620
rect -1050 7598 -1046 7620
rect -1026 7598 -1022 7620
rect -1002 7598 -998 7620
rect -978 7598 -974 7620
rect -954 7598 -950 7620
rect -930 7598 -926 7620
rect -906 7598 -902 7620
rect -882 7598 -878 7620
rect -858 7598 -854 7620
rect -834 7598 -830 7620
rect -810 7598 -806 7620
rect -786 7598 -782 7620
rect -762 7598 -758 7620
rect -738 7598 -734 7620
rect -714 7598 -710 7620
rect -690 7598 -686 7620
rect -666 7598 -662 7620
rect -642 7598 -638 7620
rect -618 7598 -614 7620
rect -594 7598 -590 7620
rect -570 7598 -566 7620
rect -546 7598 -542 7620
rect -522 7598 -518 7620
rect -498 7598 -494 7620
rect -474 7598 -470 7620
rect -450 7598 -446 7620
rect -426 7598 -422 7620
rect -402 7598 -398 7620
rect -378 7598 -374 7620
rect -354 7598 -350 7620
rect -330 7598 -326 7620
rect -306 7598 -302 7620
rect -282 7598 -278 7620
rect -258 7598 -254 7620
rect -234 7598 -230 7620
rect -210 7598 -206 7620
rect -186 7598 -182 7620
rect -162 7598 -158 7620
rect -138 7619 -134 7620
rect -2393 7596 -141 7598
rect -2371 7502 -2366 7596
rect -2348 7502 -2343 7596
rect -2325 7594 -2320 7596
rect -2317 7594 -2309 7596
rect -2325 7582 -2317 7594
rect -2060 7583 -2030 7590
rect -2325 7562 -2320 7582
rect -2325 7554 -2317 7562
rect -2060 7556 -2030 7559
rect -2325 7506 -2320 7554
rect -2317 7546 -2309 7554
rect -2060 7543 -2038 7554
rect -2033 7547 -2030 7556
rect -2028 7552 -2027 7556
rect -2068 7538 -2038 7541
rect -2325 7502 -2317 7506
rect -2000 7504 -1992 7596
rect -1844 7592 -1804 7596
rect -1663 7594 -1655 7596
rect -1844 7582 -1794 7591
rect -1671 7582 -1663 7594
rect -1912 7571 -1884 7573
rect -1852 7565 -1804 7569
rect -1844 7556 -1796 7559
rect -1671 7554 -1663 7562
rect -1844 7543 -1804 7554
rect -1663 7546 -1655 7554
rect -1852 7538 -1680 7542
rect -2000 7502 -1957 7504
rect -1671 7502 -1663 7506
rect -1642 7502 -1637 7596
rect -1619 7502 -1614 7596
rect -1530 7502 -1526 7596
rect -1506 7502 -1502 7596
rect -1482 7502 -1478 7596
rect -1458 7502 -1454 7596
rect -1434 7502 -1430 7596
rect -1410 7502 -1406 7596
rect -1386 7502 -1382 7596
rect -1362 7502 -1358 7596
rect -1338 7502 -1334 7596
rect -1314 7502 -1310 7596
rect -1290 7502 -1286 7596
rect -1266 7502 -1262 7596
rect -1242 7502 -1238 7596
rect -1218 7502 -1214 7596
rect -1194 7502 -1190 7596
rect -1170 7502 -1166 7596
rect -1146 7502 -1142 7596
rect -1122 7502 -1118 7596
rect -1098 7502 -1094 7596
rect -1074 7502 -1070 7596
rect -1050 7502 -1046 7596
rect -1026 7502 -1022 7596
rect -1002 7502 -998 7596
rect -978 7502 -974 7596
rect -954 7502 -950 7596
rect -930 7502 -926 7596
rect -906 7502 -902 7596
rect -882 7502 -878 7596
rect -858 7502 -854 7596
rect -834 7503 -830 7596
rect -845 7502 -811 7503
rect -2393 7500 -811 7502
rect -2371 4670 -2366 7500
rect -2348 4670 -2343 7500
rect -2325 7478 -2320 7500
rect -2317 7490 -2309 7500
rect -2325 7474 -2317 7478
rect -2325 7426 -2320 7474
rect -2317 7462 -2309 7474
rect -2163 7462 -2127 7465
rect -2124 7462 -2108 7466
rect -2060 7462 -2030 7466
rect -2325 7418 -2317 7426
rect -2325 7398 -2320 7418
rect -2317 7410 -2309 7418
rect -2325 7390 -2317 7398
rect -2325 7370 -2320 7390
rect -2317 7382 -2309 7390
rect -2127 7378 -2097 7379
rect -2325 7362 -2317 7370
rect -2325 7342 -2320 7362
rect -2317 7355 -2309 7362
rect -2127 7358 -2124 7367
rect -2119 7358 -2097 7371
rect -2092 7365 -2089 7371
rect -2087 7368 -2079 7381
rect -2127 7357 -2097 7358
rect -2317 7354 -2301 7355
rect -2309 7343 -2307 7354
rect -2145 7346 -2129 7353
rect -2066 7352 -2065 7353
rect -2325 7334 -2317 7342
rect -2325 7210 -2320 7334
rect -2317 7326 -2309 7334
rect -2297 7327 -2289 7343
rect -2150 7341 -2141 7343
rect -2129 7341 -2113 7343
rect -2119 7332 -2113 7341
rect -2125 7327 -2113 7332
rect -2101 7339 -2085 7343
rect -2101 7327 -2089 7339
rect -2317 7270 -2309 7286
rect -2317 7242 -2309 7258
rect -2193 7253 -2189 7263
rect -2199 7251 -2189 7253
rect -2177 7253 -2163 7263
rect -2177 7251 -2161 7253
rect -2325 7202 -2317 7210
rect -2325 7182 -2320 7202
rect -2317 7194 -2309 7202
rect -2325 7174 -2317 7182
rect -2325 7154 -2320 7174
rect -2317 7166 -2309 7174
rect -2127 7162 -2097 7163
rect -2325 7146 -2317 7154
rect -2325 7126 -2320 7146
rect -2317 7139 -2309 7146
rect -2127 7142 -2124 7151
rect -2119 7142 -2097 7155
rect -2092 7149 -2089 7155
rect -2087 7152 -2079 7165
rect -2127 7141 -2097 7142
rect -2317 7138 -2301 7139
rect -2309 7127 -2307 7138
rect -2145 7130 -2129 7137
rect -2066 7136 -2065 7137
rect -2325 7118 -2317 7126
rect -2325 6994 -2320 7118
rect -2317 7110 -2309 7118
rect -2297 7111 -2289 7127
rect -2150 7125 -2141 7127
rect -2129 7125 -2113 7127
rect -2119 7116 -2113 7125
rect -2125 7111 -2113 7116
rect -2101 7123 -2085 7127
rect -2101 7111 -2089 7123
rect -2317 7054 -2309 7070
rect -2317 7026 -2309 7042
rect -2193 7037 -2189 7047
rect -2199 7035 -2189 7037
rect -2177 7037 -2163 7047
rect -2177 7035 -2161 7037
rect -2325 6986 -2317 6994
rect -2325 6966 -2320 6986
rect -2317 6978 -2309 6986
rect -2325 6958 -2317 6966
rect -2325 6938 -2320 6958
rect -2317 6950 -2309 6958
rect -2127 6946 -2097 6947
rect -2325 6930 -2317 6938
rect -2325 6910 -2320 6930
rect -2317 6923 -2309 6930
rect -2127 6926 -2124 6935
rect -2119 6926 -2097 6939
rect -2092 6933 -2089 6939
rect -2087 6936 -2079 6949
rect -2127 6925 -2097 6926
rect -2317 6922 -2301 6923
rect -2309 6911 -2307 6922
rect -2145 6914 -2129 6921
rect -2066 6920 -2065 6921
rect -2325 6902 -2317 6910
rect -2325 6778 -2320 6902
rect -2317 6894 -2309 6902
rect -2297 6895 -2289 6911
rect -2150 6909 -2141 6911
rect -2129 6909 -2113 6911
rect -2119 6900 -2113 6909
rect -2125 6895 -2113 6900
rect -2101 6907 -2085 6911
rect -2101 6895 -2089 6907
rect -2317 6838 -2309 6854
rect -2317 6810 -2309 6826
rect -2193 6821 -2189 6831
rect -2199 6819 -2189 6821
rect -2177 6821 -2163 6831
rect -2177 6819 -2161 6821
rect -2325 6770 -2317 6778
rect -2325 6750 -2320 6770
rect -2317 6762 -2309 6770
rect -2325 6742 -2317 6750
rect -2325 6722 -2320 6742
rect -2317 6734 -2309 6742
rect -2127 6730 -2097 6731
rect -2325 6714 -2317 6722
rect -2325 6694 -2320 6714
rect -2317 6707 -2309 6714
rect -2127 6710 -2124 6719
rect -2119 6710 -2097 6723
rect -2092 6717 -2089 6723
rect -2087 6720 -2079 6733
rect -2127 6709 -2097 6710
rect -2317 6706 -2301 6707
rect -2309 6695 -2307 6706
rect -2145 6698 -2129 6705
rect -2066 6704 -2065 6705
rect -2325 6686 -2317 6694
rect -2325 6562 -2320 6686
rect -2317 6678 -2309 6686
rect -2297 6679 -2289 6695
rect -2150 6693 -2141 6695
rect -2129 6693 -2113 6695
rect -2119 6684 -2113 6693
rect -2125 6679 -2113 6684
rect -2101 6691 -2085 6695
rect -2101 6679 -2089 6691
rect -2317 6622 -2309 6638
rect -2317 6594 -2309 6610
rect -2193 6605 -2189 6615
rect -2199 6603 -2189 6605
rect -2177 6605 -2163 6615
rect -2177 6603 -2161 6605
rect -2325 6554 -2317 6562
rect -2325 6534 -2320 6554
rect -2317 6546 -2309 6554
rect -2325 6526 -2317 6534
rect -2325 6506 -2320 6526
rect -2317 6518 -2309 6526
rect -2127 6514 -2097 6515
rect -2325 6498 -2317 6506
rect -2325 6478 -2320 6498
rect -2317 6491 -2309 6498
rect -2127 6494 -2124 6503
rect -2119 6494 -2097 6507
rect -2092 6501 -2089 6507
rect -2087 6504 -2079 6517
rect -2127 6493 -2097 6494
rect -2317 6490 -2301 6491
rect -2309 6479 -2307 6490
rect -2145 6482 -2129 6489
rect -2066 6488 -2065 6489
rect -2325 6470 -2317 6478
rect -2325 6346 -2320 6470
rect -2317 6462 -2309 6470
rect -2297 6463 -2289 6479
rect -2150 6477 -2141 6479
rect -2129 6477 -2113 6479
rect -2119 6468 -2113 6477
rect -2125 6463 -2113 6468
rect -2101 6475 -2085 6479
rect -2101 6463 -2089 6475
rect -2317 6406 -2309 6422
rect -2317 6378 -2309 6394
rect -2193 6389 -2189 6399
rect -2199 6387 -2189 6389
rect -2177 6389 -2163 6399
rect -2177 6387 -2161 6389
rect -2325 6338 -2317 6346
rect -2325 6318 -2320 6338
rect -2317 6330 -2309 6338
rect -2325 6310 -2317 6318
rect -2325 6290 -2320 6310
rect -2317 6302 -2309 6310
rect -2127 6298 -2097 6299
rect -2325 6282 -2317 6290
rect -2325 6262 -2320 6282
rect -2317 6275 -2309 6282
rect -2127 6278 -2124 6287
rect -2119 6278 -2097 6291
rect -2092 6285 -2089 6291
rect -2087 6288 -2079 6301
rect -2127 6277 -2097 6278
rect -2317 6274 -2301 6275
rect -2309 6263 -2307 6274
rect -2145 6266 -2129 6273
rect -2066 6272 -2065 6273
rect -2325 6254 -2317 6262
rect -2325 6130 -2320 6254
rect -2317 6246 -2309 6254
rect -2297 6247 -2289 6263
rect -2150 6261 -2141 6263
rect -2129 6261 -2113 6263
rect -2119 6252 -2113 6261
rect -2125 6247 -2113 6252
rect -2101 6259 -2085 6263
rect -2101 6247 -2089 6259
rect -2317 6190 -2309 6206
rect -2317 6162 -2309 6178
rect -2193 6173 -2189 6183
rect -2199 6171 -2189 6173
rect -2177 6173 -2163 6183
rect -2177 6171 -2161 6173
rect -2325 6122 -2317 6130
rect -2325 6102 -2320 6122
rect -2317 6114 -2309 6122
rect -2325 6094 -2317 6102
rect -2325 6074 -2320 6094
rect -2317 6086 -2309 6094
rect -2127 6082 -2097 6083
rect -2325 6066 -2317 6074
rect -2325 6046 -2320 6066
rect -2317 6059 -2309 6066
rect -2127 6062 -2124 6071
rect -2119 6062 -2097 6075
rect -2092 6069 -2089 6075
rect -2087 6072 -2079 6085
rect -2127 6061 -2097 6062
rect -2317 6058 -2301 6059
rect -2309 6047 -2307 6058
rect -2145 6050 -2129 6057
rect -2066 6056 -2065 6057
rect -2325 6038 -2317 6046
rect -2325 5914 -2320 6038
rect -2317 6030 -2309 6038
rect -2297 6031 -2289 6047
rect -2150 6045 -2141 6047
rect -2129 6045 -2113 6047
rect -2119 6036 -2113 6045
rect -2125 6031 -2113 6036
rect -2101 6043 -2085 6047
rect -2101 6031 -2089 6043
rect -2317 5974 -2309 5990
rect -2317 5946 -2309 5962
rect -2193 5957 -2189 5967
rect -2199 5955 -2189 5957
rect -2177 5957 -2163 5967
rect -2177 5955 -2161 5957
rect -2325 5906 -2317 5914
rect -2325 5886 -2320 5906
rect -2317 5898 -2309 5906
rect -2325 5878 -2317 5886
rect -2325 5858 -2320 5878
rect -2317 5870 -2309 5878
rect -2127 5866 -2097 5867
rect -2325 5850 -2317 5858
rect -2325 5830 -2320 5850
rect -2317 5843 -2309 5850
rect -2127 5846 -2124 5855
rect -2119 5846 -2097 5859
rect -2092 5853 -2089 5859
rect -2087 5856 -2079 5869
rect -2127 5845 -2097 5846
rect -2317 5842 -2301 5843
rect -2309 5831 -2307 5842
rect -2145 5834 -2129 5841
rect -2066 5840 -2065 5841
rect -2325 5822 -2317 5830
rect -2325 5698 -2320 5822
rect -2317 5814 -2309 5822
rect -2297 5815 -2289 5831
rect -2150 5829 -2141 5831
rect -2129 5829 -2113 5831
rect -2119 5820 -2113 5829
rect -2125 5815 -2113 5820
rect -2101 5827 -2085 5831
rect -2101 5815 -2089 5827
rect -2317 5758 -2309 5774
rect -2317 5730 -2309 5746
rect -2193 5741 -2189 5751
rect -2199 5739 -2189 5741
rect -2177 5741 -2163 5751
rect -2177 5739 -2161 5741
rect -2325 5690 -2317 5698
rect -2325 5670 -2320 5690
rect -2317 5682 -2309 5690
rect -2325 5662 -2317 5670
rect -2325 5642 -2320 5662
rect -2317 5654 -2309 5662
rect -2127 5650 -2097 5651
rect -2325 5634 -2317 5642
rect -2325 5614 -2320 5634
rect -2317 5627 -2309 5634
rect -2127 5630 -2124 5639
rect -2119 5630 -2097 5643
rect -2092 5637 -2089 5643
rect -2087 5640 -2079 5653
rect -2127 5629 -2097 5630
rect -2317 5626 -2301 5627
rect -2309 5615 -2307 5626
rect -2145 5618 -2129 5625
rect -2066 5624 -2065 5625
rect -2325 5606 -2317 5614
rect -2325 5482 -2320 5606
rect -2317 5598 -2309 5606
rect -2297 5599 -2289 5615
rect -2150 5613 -2141 5615
rect -2129 5613 -2113 5615
rect -2119 5604 -2113 5613
rect -2125 5599 -2113 5604
rect -2101 5611 -2085 5615
rect -2101 5599 -2089 5611
rect -2317 5542 -2309 5558
rect -2317 5514 -2309 5530
rect -2193 5525 -2189 5535
rect -2199 5523 -2189 5525
rect -2177 5525 -2163 5535
rect -2177 5523 -2161 5525
rect -2325 5474 -2317 5482
rect -2325 5454 -2320 5474
rect -2317 5466 -2309 5474
rect -2325 5446 -2317 5454
rect -2325 5426 -2320 5446
rect -2317 5438 -2309 5446
rect -2127 5434 -2097 5435
rect -2325 5418 -2317 5426
rect -2325 5398 -2320 5418
rect -2317 5411 -2309 5418
rect -2127 5414 -2124 5423
rect -2119 5414 -2097 5427
rect -2092 5421 -2089 5427
rect -2087 5424 -2079 5437
rect -2127 5413 -2097 5414
rect -2317 5410 -2301 5411
rect -2309 5399 -2307 5410
rect -2145 5402 -2129 5409
rect -2066 5408 -2065 5409
rect -2325 5390 -2317 5398
rect -2325 5266 -2320 5390
rect -2317 5382 -2309 5390
rect -2297 5383 -2289 5399
rect -2150 5397 -2141 5399
rect -2129 5397 -2113 5399
rect -2119 5388 -2113 5397
rect -2125 5383 -2113 5388
rect -2101 5395 -2085 5399
rect -2101 5383 -2089 5395
rect -2317 5326 -2309 5342
rect -2317 5298 -2309 5314
rect -2193 5309 -2189 5319
rect -2199 5307 -2189 5309
rect -2177 5309 -2163 5319
rect -2177 5307 -2161 5309
rect -2325 5258 -2317 5266
rect -2325 5238 -2320 5258
rect -2317 5250 -2309 5258
rect -2325 5230 -2317 5238
rect -2325 5210 -2320 5230
rect -2317 5222 -2309 5230
rect -2127 5218 -2097 5219
rect -2325 5202 -2317 5210
rect -2325 5182 -2320 5202
rect -2317 5195 -2309 5202
rect -2127 5198 -2124 5207
rect -2119 5198 -2097 5211
rect -2092 5205 -2089 5211
rect -2087 5208 -2079 5221
rect -2127 5197 -2097 5198
rect -2317 5194 -2301 5195
rect -2309 5183 -2307 5194
rect -2145 5186 -2129 5193
rect -2066 5192 -2065 5193
rect -2325 5174 -2317 5182
rect -2325 5050 -2320 5174
rect -2317 5166 -2309 5174
rect -2297 5167 -2289 5183
rect -2150 5181 -2141 5183
rect -2129 5181 -2113 5183
rect -2119 5172 -2113 5181
rect -2125 5167 -2113 5172
rect -2101 5179 -2085 5183
rect -2101 5167 -2089 5179
rect -2317 5110 -2309 5126
rect -2317 5082 -2309 5098
rect -2193 5093 -2189 5103
rect -2199 5091 -2189 5093
rect -2177 5093 -2163 5103
rect -2177 5091 -2161 5093
rect -2325 5042 -2317 5050
rect -2325 5022 -2320 5042
rect -2317 5034 -2309 5042
rect -2325 5014 -2317 5022
rect -2325 4994 -2320 5014
rect -2317 5006 -2309 5014
rect -2127 5002 -2097 5003
rect -2325 4986 -2317 4994
rect -2325 4966 -2320 4986
rect -2317 4979 -2309 4986
rect -2127 4982 -2124 4991
rect -2119 4982 -2097 4995
rect -2092 4989 -2089 4995
rect -2087 4992 -2079 5005
rect -2127 4981 -2097 4982
rect -2317 4978 -2301 4979
rect -2309 4967 -2307 4978
rect -2145 4970 -2129 4977
rect -2066 4976 -2065 4977
rect -2325 4958 -2317 4966
rect -2325 4834 -2320 4958
rect -2317 4950 -2309 4958
rect -2297 4951 -2289 4967
rect -2150 4965 -2141 4967
rect -2129 4965 -2113 4967
rect -2119 4956 -2113 4965
rect -2125 4951 -2113 4956
rect -2101 4963 -2085 4967
rect -2101 4951 -2089 4963
rect -2317 4894 -2309 4910
rect -2317 4866 -2309 4882
rect -2193 4877 -2189 4887
rect -2199 4875 -2189 4877
rect -2177 4877 -2163 4887
rect -2177 4875 -2161 4877
rect -2325 4826 -2317 4834
rect -2325 4806 -2320 4826
rect -2317 4818 -2309 4826
rect -2325 4798 -2317 4806
rect -2325 4778 -2320 4798
rect -2317 4790 -2309 4798
rect -2127 4786 -2097 4787
rect -2325 4770 -2317 4778
rect -2325 4750 -2320 4770
rect -2317 4763 -2309 4770
rect -2127 4766 -2124 4775
rect -2119 4766 -2097 4779
rect -2092 4773 -2089 4779
rect -2087 4776 -2079 4789
rect -2127 4765 -2097 4766
rect -2317 4762 -2301 4763
rect -2309 4751 -2307 4762
rect -2145 4754 -2129 4761
rect -2066 4760 -2065 4761
rect -2325 4742 -2317 4750
rect -2325 4722 -2320 4742
rect -2317 4734 -2309 4742
rect -2297 4735 -2289 4751
rect -2150 4749 -2141 4751
rect -2129 4749 -2113 4751
rect -2119 4740 -2113 4749
rect -2125 4735 -2113 4740
rect -2101 4747 -2085 4751
rect -2101 4735 -2089 4747
rect -2325 4710 -2317 4722
rect -2325 4694 -2320 4710
rect -2317 4706 -2309 4710
rect -2068 4706 -2038 4707
rect -2309 4694 -2301 4706
rect -2068 4702 -2063 4706
rect -2000 4702 -1992 7500
rect -1972 7498 -1957 7500
rect -1958 7497 -1957 7498
rect -1984 7476 -1980 7494
rect -1663 7490 -1655 7500
rect -1832 7489 -1796 7490
rect -1824 7480 -1796 7482
rect -1954 7476 -1918 7480
rect -1796 7479 -1788 7480
rect -1822 7466 -1796 7478
rect -1671 7474 -1663 7478
rect -1857 7456 -1850 7466
rect -1844 7462 -1796 7466
rect -1663 7462 -1655 7474
rect -1847 7453 -1840 7456
rect -1671 7418 -1663 7426
rect -1663 7410 -1655 7418
rect -1946 7396 -1893 7404
rect -1927 7386 -1919 7394
rect -1901 7386 -1898 7396
rect -1671 7390 -1663 7398
rect -1927 7380 -1920 7386
rect -1936 7378 -1920 7380
rect -1919 7385 -1911 7386
rect -1919 7378 -1903 7385
rect -1901 7379 -1900 7386
rect -1663 7382 -1655 7390
rect -1901 7378 -1853 7379
rect -1893 7358 -1853 7371
rect -1671 7362 -1663 7370
rect -1901 7357 -1853 7358
rect -1663 7354 -1655 7362
rect -1915 7346 -1914 7353
rect -1767 7346 -1766 7353
rect -1671 7334 -1663 7342
rect -1663 7326 -1655 7334
rect -1977 7278 -1972 7288
rect -1663 7270 -1655 7286
rect -1972 7264 -1967 7267
rect -1944 7251 -1928 7254
rect -1927 7251 -1924 7254
rect -1663 7242 -1655 7258
rect -1671 7202 -1663 7210
rect -1663 7194 -1655 7202
rect -1946 7180 -1893 7188
rect -1927 7170 -1919 7178
rect -1901 7170 -1898 7180
rect -1671 7174 -1663 7182
rect -1927 7164 -1920 7170
rect -1936 7162 -1920 7164
rect -1919 7169 -1911 7170
rect -1919 7162 -1903 7169
rect -1901 7163 -1900 7170
rect -1663 7166 -1655 7174
rect -1901 7162 -1853 7163
rect -1893 7142 -1853 7155
rect -1671 7146 -1663 7154
rect -1901 7141 -1853 7142
rect -1663 7138 -1655 7146
rect -1915 7130 -1914 7137
rect -1767 7130 -1766 7137
rect -1671 7118 -1663 7126
rect -1663 7110 -1655 7118
rect -1977 7062 -1972 7072
rect -1663 7054 -1655 7070
rect -1972 7048 -1967 7051
rect -1944 7035 -1928 7038
rect -1927 7035 -1924 7038
rect -1663 7026 -1655 7042
rect -1671 6986 -1663 6994
rect -1663 6978 -1655 6986
rect -1946 6964 -1893 6972
rect -1927 6954 -1919 6962
rect -1901 6954 -1898 6964
rect -1671 6958 -1663 6966
rect -1927 6948 -1920 6954
rect -1936 6946 -1920 6948
rect -1919 6953 -1911 6954
rect -1919 6946 -1903 6953
rect -1901 6947 -1900 6954
rect -1663 6950 -1655 6958
rect -1901 6946 -1853 6947
rect -1893 6926 -1853 6939
rect -1671 6930 -1663 6938
rect -1901 6925 -1853 6926
rect -1663 6922 -1655 6930
rect -1915 6914 -1914 6921
rect -1767 6914 -1766 6921
rect -1671 6902 -1663 6910
rect -1663 6894 -1655 6902
rect -1977 6846 -1972 6856
rect -1663 6838 -1655 6854
rect -1972 6832 -1967 6835
rect -1944 6819 -1928 6822
rect -1927 6819 -1924 6822
rect -1663 6810 -1655 6826
rect -1671 6770 -1663 6778
rect -1663 6762 -1655 6770
rect -1946 6748 -1893 6756
rect -1927 6738 -1919 6746
rect -1901 6738 -1898 6748
rect -1671 6742 -1663 6750
rect -1927 6732 -1920 6738
rect -1936 6730 -1920 6732
rect -1919 6737 -1911 6738
rect -1919 6730 -1903 6737
rect -1901 6731 -1900 6738
rect -1663 6734 -1655 6742
rect -1901 6730 -1853 6731
rect -1893 6710 -1853 6723
rect -1671 6714 -1663 6722
rect -1901 6709 -1853 6710
rect -1663 6706 -1655 6714
rect -1915 6698 -1914 6705
rect -1767 6698 -1766 6705
rect -1671 6686 -1663 6694
rect -1663 6678 -1655 6686
rect -1977 6630 -1972 6640
rect -1663 6622 -1655 6638
rect -1972 6616 -1967 6619
rect -1944 6603 -1928 6606
rect -1927 6603 -1924 6606
rect -1663 6594 -1655 6610
rect -1671 6554 -1663 6562
rect -1663 6546 -1655 6554
rect -1946 6532 -1893 6540
rect -1927 6522 -1919 6530
rect -1901 6522 -1898 6532
rect -1671 6526 -1663 6534
rect -1927 6516 -1920 6522
rect -1936 6514 -1920 6516
rect -1919 6521 -1911 6522
rect -1919 6514 -1903 6521
rect -1901 6515 -1900 6522
rect -1663 6518 -1655 6526
rect -1901 6514 -1853 6515
rect -1893 6494 -1853 6507
rect -1671 6498 -1663 6506
rect -1901 6493 -1853 6494
rect -1663 6490 -1655 6498
rect -1915 6482 -1914 6489
rect -1767 6482 -1766 6489
rect -1671 6470 -1663 6478
rect -1663 6462 -1655 6470
rect -1977 6414 -1972 6424
rect -1663 6406 -1655 6422
rect -1972 6400 -1967 6403
rect -1944 6387 -1928 6390
rect -1927 6387 -1924 6390
rect -1663 6378 -1655 6394
rect -1671 6338 -1663 6346
rect -1663 6330 -1655 6338
rect -1946 6316 -1893 6324
rect -1927 6306 -1919 6314
rect -1901 6306 -1898 6316
rect -1671 6310 -1663 6318
rect -1927 6300 -1920 6306
rect -1936 6298 -1920 6300
rect -1919 6305 -1911 6306
rect -1919 6298 -1903 6305
rect -1901 6299 -1900 6306
rect -1663 6302 -1655 6310
rect -1901 6298 -1853 6299
rect -1893 6278 -1853 6291
rect -1671 6282 -1663 6290
rect -1901 6277 -1853 6278
rect -1663 6274 -1655 6282
rect -1915 6266 -1914 6273
rect -1767 6266 -1766 6273
rect -1671 6254 -1663 6262
rect -1663 6246 -1655 6254
rect -1977 6198 -1972 6208
rect -1663 6190 -1655 6206
rect -1972 6184 -1967 6187
rect -1944 6171 -1928 6174
rect -1927 6171 -1924 6174
rect -1663 6162 -1655 6178
rect -1671 6122 -1663 6130
rect -1663 6114 -1655 6122
rect -1946 6100 -1893 6108
rect -1927 6090 -1919 6098
rect -1901 6090 -1898 6100
rect -1671 6094 -1663 6102
rect -1927 6084 -1920 6090
rect -1936 6082 -1920 6084
rect -1919 6089 -1911 6090
rect -1919 6082 -1903 6089
rect -1901 6083 -1900 6090
rect -1663 6086 -1655 6094
rect -1901 6082 -1853 6083
rect -1893 6062 -1853 6075
rect -1671 6066 -1663 6074
rect -1901 6061 -1853 6062
rect -1663 6058 -1655 6066
rect -1915 6050 -1914 6057
rect -1767 6050 -1766 6057
rect -1671 6038 -1663 6046
rect -1663 6030 -1655 6038
rect -1977 5982 -1972 5992
rect -1663 5974 -1655 5990
rect -1972 5968 -1967 5971
rect -1944 5955 -1928 5958
rect -1927 5955 -1924 5958
rect -1663 5946 -1655 5962
rect -1671 5906 -1663 5914
rect -1663 5898 -1655 5906
rect -1946 5884 -1893 5892
rect -1927 5874 -1919 5882
rect -1901 5874 -1898 5884
rect -1671 5878 -1663 5886
rect -1927 5868 -1920 5874
rect -1936 5866 -1920 5868
rect -1919 5873 -1911 5874
rect -1919 5866 -1903 5873
rect -1901 5867 -1900 5874
rect -1663 5870 -1655 5878
rect -1901 5866 -1853 5867
rect -1893 5846 -1853 5859
rect -1671 5850 -1663 5858
rect -1901 5845 -1853 5846
rect -1663 5842 -1655 5850
rect -1915 5834 -1914 5841
rect -1767 5834 -1766 5841
rect -1671 5822 -1663 5830
rect -1663 5814 -1655 5822
rect -1977 5766 -1972 5776
rect -1663 5758 -1655 5774
rect -1972 5752 -1967 5755
rect -1944 5739 -1928 5742
rect -1927 5739 -1924 5742
rect -1663 5730 -1655 5746
rect -1671 5690 -1663 5698
rect -1663 5682 -1655 5690
rect -1946 5668 -1893 5676
rect -1927 5658 -1919 5666
rect -1901 5658 -1898 5668
rect -1671 5662 -1663 5670
rect -1927 5652 -1920 5658
rect -1936 5650 -1920 5652
rect -1919 5657 -1911 5658
rect -1919 5650 -1903 5657
rect -1901 5651 -1900 5658
rect -1663 5654 -1655 5662
rect -1901 5650 -1853 5651
rect -1893 5630 -1853 5643
rect -1671 5634 -1663 5642
rect -1901 5629 -1853 5630
rect -1663 5626 -1655 5634
rect -1915 5618 -1914 5625
rect -1767 5618 -1766 5625
rect -1671 5606 -1663 5614
rect -1663 5598 -1655 5606
rect -1977 5550 -1972 5560
rect -1663 5542 -1655 5558
rect -1972 5536 -1967 5539
rect -1944 5523 -1928 5526
rect -1927 5523 -1924 5526
rect -1663 5514 -1655 5530
rect -1671 5474 -1663 5482
rect -1663 5466 -1655 5474
rect -1946 5452 -1893 5460
rect -1927 5442 -1919 5450
rect -1901 5442 -1898 5452
rect -1671 5446 -1663 5454
rect -1927 5436 -1920 5442
rect -1936 5434 -1920 5436
rect -1919 5441 -1911 5442
rect -1919 5434 -1903 5441
rect -1901 5435 -1900 5442
rect -1663 5438 -1655 5446
rect -1901 5434 -1853 5435
rect -1893 5414 -1853 5427
rect -1671 5418 -1663 5426
rect -1901 5413 -1853 5414
rect -1663 5410 -1655 5418
rect -1915 5402 -1914 5409
rect -1767 5402 -1766 5409
rect -1671 5390 -1663 5398
rect -1663 5382 -1655 5390
rect -1977 5334 -1972 5344
rect -1663 5326 -1655 5342
rect -1972 5320 -1967 5323
rect -1944 5307 -1928 5310
rect -1927 5307 -1924 5310
rect -1663 5298 -1655 5314
rect -1671 5258 -1663 5266
rect -1663 5250 -1655 5258
rect -1946 5236 -1893 5244
rect -1927 5226 -1919 5234
rect -1901 5226 -1898 5236
rect -1671 5230 -1663 5238
rect -1927 5220 -1920 5226
rect -1936 5218 -1920 5220
rect -1919 5225 -1911 5226
rect -1919 5218 -1903 5225
rect -1901 5219 -1900 5226
rect -1663 5222 -1655 5230
rect -1901 5218 -1853 5219
rect -1893 5198 -1853 5211
rect -1671 5202 -1663 5210
rect -1901 5197 -1853 5198
rect -1663 5194 -1655 5202
rect -1915 5186 -1914 5193
rect -1767 5186 -1766 5193
rect -1671 5174 -1663 5182
rect -1663 5166 -1655 5174
rect -1977 5118 -1972 5128
rect -1663 5110 -1655 5126
rect -1972 5104 -1967 5107
rect -1944 5091 -1928 5094
rect -1927 5091 -1924 5094
rect -1663 5082 -1655 5098
rect -1671 5042 -1663 5050
rect -1663 5034 -1655 5042
rect -1946 5020 -1893 5028
rect -1927 5010 -1919 5018
rect -1901 5010 -1898 5020
rect -1671 5014 -1663 5022
rect -1927 5004 -1920 5010
rect -1936 5002 -1920 5004
rect -1919 5009 -1911 5010
rect -1919 5002 -1903 5009
rect -1901 5003 -1900 5010
rect -1663 5006 -1655 5014
rect -1901 5002 -1853 5003
rect -1893 4982 -1853 4995
rect -1671 4986 -1663 4994
rect -1901 4981 -1853 4982
rect -1663 4978 -1655 4986
rect -1915 4970 -1914 4977
rect -1767 4970 -1766 4977
rect -1671 4958 -1663 4966
rect -1663 4950 -1655 4958
rect -1977 4902 -1972 4912
rect -1663 4894 -1655 4910
rect -1972 4888 -1967 4891
rect -1944 4875 -1928 4878
rect -1927 4875 -1924 4878
rect -1663 4866 -1655 4882
rect -1671 4826 -1663 4834
rect -1663 4818 -1655 4826
rect -1946 4804 -1893 4812
rect -1927 4794 -1919 4802
rect -1901 4794 -1898 4804
rect -1671 4798 -1663 4806
rect -1927 4788 -1920 4794
rect -1936 4786 -1920 4788
rect -1919 4793 -1911 4794
rect -1919 4786 -1903 4793
rect -1901 4787 -1900 4794
rect -1663 4790 -1655 4798
rect -1901 4786 -1853 4787
rect -1893 4766 -1853 4779
rect -1671 4770 -1663 4778
rect -1901 4765 -1853 4766
rect -1663 4762 -1655 4770
rect -1915 4754 -1914 4761
rect -1767 4754 -1766 4761
rect -1671 4742 -1663 4750
rect -1663 4734 -1655 4742
rect -2325 4682 -2317 4694
rect -2058 4691 -2038 4702
rect -2028 4698 -1992 4702
rect -1916 4701 -1903 4711
rect -1671 4710 -1663 4722
rect -1852 4706 -1832 4707
rect -1663 4706 -1655 4710
rect -2068 4682 -2065 4687
rect -2058 4686 -2028 4689
rect -2011 4688 -2002 4692
rect -2000 4688 -1992 4698
rect -1893 4690 -1892 4697
rect -1852 4691 -1845 4706
rect -1655 4694 -1647 4706
rect -1854 4690 -1845 4691
rect -1893 4689 -1680 4690
rect -2001 4686 -1992 4688
rect -2038 4684 -2028 4686
rect -2058 4682 -2038 4684
rect -2325 4670 -2320 4682
rect -2317 4678 -2309 4682
rect -2309 4670 -2301 4678
rect -2068 4677 -2058 4682
rect -2068 4670 -2065 4677
rect -2016 4676 -2002 4686
rect -2000 4677 -1992 4686
rect -1972 4684 -1924 4689
rect -1671 4682 -1663 4694
rect -1663 4678 -1655 4682
rect -2001 4676 -1992 4677
rect -2015 4672 -2002 4676
rect -2000 4670 -1992 4676
rect -1976 4670 -1940 4671
rect -1655 4670 -1647 4678
rect -1642 4670 -1637 7500
rect -1619 4670 -1614 7500
rect -1530 4670 -1526 7500
rect -1506 4670 -1502 7500
rect -1482 4670 -1478 7500
rect -1458 4670 -1454 7500
rect -1434 4670 -1430 7500
rect -1410 4670 -1406 7500
rect -1386 4670 -1382 7500
rect -1362 4670 -1358 7500
rect -1338 4670 -1334 7500
rect -1314 4670 -1310 7500
rect -1290 4670 -1286 7500
rect -1277 4901 -1272 4911
rect -1266 4901 -1262 7500
rect -1267 4887 -1262 4901
rect -1277 4886 -1243 4887
rect -1242 4886 -1238 7500
rect -1218 4886 -1214 7500
rect -1194 4886 -1190 7500
rect -1170 4886 -1166 7500
rect -1146 4886 -1142 7500
rect -1122 4886 -1118 7500
rect -1098 4886 -1094 7500
rect -1074 4886 -1070 7500
rect -1050 4886 -1046 7500
rect -1026 4886 -1022 7500
rect -1002 4886 -998 7500
rect -978 4886 -974 7500
rect -954 4886 -950 7500
rect -930 4886 -926 7500
rect -906 4886 -902 7500
rect -882 4886 -878 7500
rect -858 4886 -854 7500
rect -845 7493 -840 7500
rect -834 7493 -830 7500
rect -835 7479 -830 7493
rect -834 4886 -830 7479
rect -810 7427 -806 7596
rect -810 7403 -803 7427
rect -810 4886 -806 7403
rect -786 4886 -782 7596
rect -762 4886 -758 7596
rect -738 4886 -734 7596
rect -714 4886 -710 7596
rect -701 7277 -696 7287
rect -690 7277 -686 7596
rect -691 7263 -686 7277
rect -690 4886 -686 7263
rect -666 7211 -662 7596
rect -666 7187 -659 7211
rect -666 4886 -662 7187
rect -642 4886 -638 7596
rect -618 4886 -614 7596
rect -594 4886 -590 7596
rect -570 4886 -566 7596
rect -546 4886 -542 7596
rect -522 4886 -518 7596
rect -498 4886 -494 7596
rect -474 4886 -470 7596
rect -450 4886 -446 7596
rect -426 4886 -422 7596
rect -402 4886 -398 7596
rect -378 4886 -374 7596
rect -354 4886 -350 7596
rect -330 4886 -326 7596
rect -306 4886 -302 7596
rect -282 4886 -278 7596
rect -258 4886 -254 7596
rect -234 4886 -230 7596
rect -210 4886 -206 7596
rect -186 4886 -182 7596
rect -162 4886 -158 7596
rect -155 7595 -141 7596
rect -138 7574 -131 7619
rect -114 7574 -110 7620
rect -90 7574 -86 7620
rect -77 7589 -72 7599
rect -66 7589 -62 7620
rect -67 7575 -62 7589
rect -42 7574 -38 7620
rect -18 7574 -14 7620
rect 6 7574 10 7620
rect 30 7574 34 7620
rect 54 7574 58 7620
rect 78 7574 82 7620
rect 102 7574 106 7620
rect 126 7574 130 7620
rect 150 7574 154 7620
rect 163 7613 168 7620
rect 174 7613 178 7620
rect 173 7599 178 7613
rect 163 7589 168 7599
rect 173 7575 178 7589
rect 174 7574 178 7575
rect 198 7574 202 7644
rect 222 7574 226 7644
rect 246 7574 250 7644
rect 270 7574 274 7644
rect 294 7574 298 7644
rect 318 7574 322 7644
rect 342 7574 346 7644
rect 366 7574 370 7644
rect 390 7574 394 7644
rect 414 7574 418 7644
rect 438 7574 442 7644
rect 462 7574 466 7644
rect 486 7574 490 7644
rect 510 7574 514 7644
rect 534 7574 538 7644
rect 558 7574 562 7644
rect 582 7574 586 7644
rect 606 7574 610 7644
rect 630 7574 634 7644
rect 654 7574 658 7644
rect 678 7574 682 7644
rect 702 7574 706 7644
rect 726 7574 730 7644
rect 750 7574 754 7644
rect 774 7575 778 7644
rect 763 7574 797 7575
rect -155 7572 797 7574
rect -155 7571 -141 7572
rect -138 7571 -131 7572
rect -138 4886 -134 7571
rect -114 4886 -110 7572
rect -90 4886 -86 7572
rect -77 7550 -43 7551
rect -42 7550 -38 7572
rect -18 7550 -14 7572
rect 6 7550 10 7572
rect 30 7550 34 7572
rect 54 7550 58 7572
rect 78 7550 82 7572
rect 102 7550 106 7572
rect 126 7550 130 7572
rect 150 7550 154 7572
rect 174 7550 178 7572
rect 198 7550 202 7572
rect 222 7550 226 7572
rect 246 7550 250 7572
rect 270 7550 274 7572
rect 294 7550 298 7572
rect 318 7550 322 7572
rect 342 7550 346 7572
rect 366 7550 370 7572
rect 390 7550 394 7572
rect 414 7550 418 7572
rect 438 7550 442 7572
rect 462 7550 466 7572
rect 486 7550 490 7572
rect 510 7550 514 7572
rect 534 7550 538 7572
rect 558 7550 562 7572
rect 582 7550 586 7572
rect 606 7550 610 7572
rect 630 7550 634 7572
rect 654 7550 658 7572
rect 678 7550 682 7572
rect 702 7550 706 7572
rect 726 7550 730 7572
rect 750 7550 754 7572
rect 763 7565 768 7572
rect 774 7565 778 7572
rect 773 7551 778 7565
rect 798 7550 802 7644
rect 822 7550 826 7644
rect 846 7550 850 7644
rect 870 7550 874 7644
rect 894 7550 898 7644
rect 918 7550 922 7644
rect 942 7550 946 7644
rect 966 7550 970 7644
rect 990 7550 994 7644
rect 1014 7550 1018 7644
rect 1038 7550 1042 7644
rect 1062 7550 1066 7644
rect 1086 7550 1090 7644
rect 1110 7550 1114 7644
rect 1134 7550 1138 7644
rect 1158 7550 1162 7644
rect 1182 7550 1186 7644
rect 1206 7550 1210 7644
rect 1230 7550 1234 7644
rect 1254 7550 1258 7644
rect 1278 7550 1282 7644
rect 1302 7550 1306 7644
rect 1326 7550 1330 7644
rect 1350 7550 1354 7644
rect 1374 7550 1378 7644
rect 1398 7550 1402 7644
rect 1422 7550 1426 7644
rect 1446 7550 1450 7644
rect 1470 7550 1474 7644
rect 1494 7550 1498 7644
rect 1518 7550 1522 7644
rect 1542 7550 1546 7644
rect 1566 7550 1570 7644
rect 1590 7550 1594 7644
rect 1614 7550 1618 7644
rect 1638 7550 1642 7644
rect 1662 7550 1666 7644
rect 1686 7550 1690 7644
rect 1710 7550 1714 7644
rect 1734 7550 1738 7644
rect 1758 7550 1762 7644
rect 1782 7550 1786 7644
rect 1806 7550 1810 7644
rect 1830 7550 1834 7644
rect 1854 7550 1858 7644
rect 1878 7550 1882 7644
rect 1902 7550 1906 7644
rect 1926 7550 1930 7644
rect 1950 7550 1954 7644
rect 1974 7550 1978 7644
rect 1998 7550 2002 7644
rect 2022 7643 2026 7644
rect 2022 7598 2029 7643
rect 2046 7598 2050 7644
rect 2070 7598 2074 7644
rect 2094 7598 2098 7644
rect 2118 7598 2122 7644
rect 2142 7598 2146 7644
rect 2166 7598 2170 7644
rect 2173 7643 2187 7644
rect 2190 7619 2197 7667
rect 2190 7598 2194 7619
rect 2214 7598 2218 7668
rect 2238 7598 2242 7668
rect 2262 7598 2266 7668
rect 2286 7598 2290 7668
rect 2310 7598 2314 7668
rect 2334 7598 2338 7668
rect 2358 7598 2362 7668
rect 2382 7598 2386 7668
rect 2406 7598 2410 7668
rect 2430 7598 2434 7668
rect 2454 7598 2458 7668
rect 2478 7598 2482 7668
rect 2502 7598 2506 7668
rect 2526 7598 2530 7668
rect 2550 7598 2554 7668
rect 2574 7598 2578 7668
rect 2598 7598 2602 7668
rect 2622 7598 2626 7668
rect 2646 7598 2650 7668
rect 2659 7661 2664 7668
rect 2670 7661 2674 7668
rect 2669 7647 2674 7661
rect 2659 7637 2664 7647
rect 2669 7623 2674 7637
rect 2670 7599 2674 7623
rect 2659 7598 2693 7599
rect 2005 7596 2693 7598
rect 2005 7595 2019 7596
rect 2022 7595 2029 7596
rect 2022 7550 2026 7595
rect 2046 7550 2050 7596
rect 2070 7550 2074 7596
rect 2094 7550 2098 7596
rect 2118 7550 2122 7596
rect 2142 7550 2146 7596
rect 2166 7550 2170 7596
rect 2190 7550 2194 7596
rect 2214 7550 2218 7596
rect 2238 7550 2242 7596
rect 2262 7550 2266 7596
rect 2286 7550 2290 7596
rect 2310 7550 2314 7596
rect 2334 7550 2338 7596
rect 2358 7550 2362 7596
rect 2382 7550 2386 7596
rect 2406 7550 2410 7596
rect 2430 7550 2434 7596
rect 2454 7550 2458 7596
rect 2478 7550 2482 7596
rect 2502 7550 2506 7596
rect 2526 7550 2530 7596
rect 2550 7550 2554 7596
rect 2574 7550 2578 7596
rect 2598 7550 2602 7596
rect 2622 7550 2626 7596
rect 2646 7551 2650 7596
rect 2659 7589 2664 7596
rect 2670 7589 2674 7596
rect 2669 7575 2674 7589
rect 2683 7585 2691 7589
rect 2677 7575 2683 7585
rect 2635 7550 2669 7551
rect -77 7548 2669 7550
rect -77 7541 -72 7548
rect -67 7527 -62 7541
rect -66 4886 -62 7527
rect -42 7523 -38 7548
rect -42 7499 -35 7523
rect -42 7451 -35 7475
rect -42 4886 -38 7451
rect -18 4886 -14 7548
rect 6 4886 10 7548
rect 30 4886 34 7548
rect 54 4886 58 7548
rect 78 4886 82 7548
rect 102 4886 106 7548
rect 126 4886 130 7548
rect 150 4886 154 7548
rect 174 4886 178 7548
rect 198 7547 202 7548
rect 198 7499 205 7547
rect 198 4886 202 7499
rect 222 4886 226 7548
rect 246 4886 250 7548
rect 270 4886 274 7548
rect 294 4886 298 7548
rect 318 4886 322 7548
rect 331 6197 336 6207
rect 342 6197 346 7548
rect 341 6183 346 6197
rect 331 6182 365 6183
rect 366 6182 370 7548
rect 379 6917 384 6927
rect 390 6917 394 7548
rect 403 7133 408 7143
rect 414 7133 418 7548
rect 413 7119 418 7133
rect 389 6903 394 6917
rect 390 6182 394 6903
rect 414 6851 418 7119
rect 438 7067 442 7548
rect 438 7043 445 7067
rect 414 6827 421 6851
rect 414 6182 418 6827
rect 438 6182 442 7043
rect 462 6182 466 7548
rect 486 6182 490 7548
rect 510 6182 514 7548
rect 534 6182 538 7548
rect 558 6182 562 7548
rect 582 6182 586 7548
rect 606 6182 610 7548
rect 630 6182 634 7548
rect 654 6182 658 7548
rect 667 6629 672 6639
rect 678 6629 682 7548
rect 677 6615 682 6629
rect 667 6614 701 6615
rect 702 6614 706 7548
rect 726 6614 730 7548
rect 750 6614 754 7548
rect 763 7517 768 7527
rect 773 7503 778 7517
rect 774 6614 778 7503
rect 798 7499 802 7548
rect 798 7475 805 7499
rect 798 7430 805 7451
rect 822 7430 826 7548
rect 846 7430 850 7548
rect 870 7430 874 7548
rect 894 7430 898 7548
rect 918 7430 922 7548
rect 942 7430 946 7548
rect 966 7430 970 7548
rect 990 7430 994 7548
rect 1014 7430 1018 7548
rect 1038 7430 1042 7548
rect 1062 7430 1066 7548
rect 1086 7430 1090 7548
rect 1110 7430 1114 7548
rect 1134 7430 1138 7548
rect 1158 7430 1162 7548
rect 1182 7430 1186 7548
rect 1206 7430 1210 7548
rect 1230 7430 1234 7548
rect 1254 7430 1258 7548
rect 1278 7430 1282 7548
rect 1302 7430 1306 7548
rect 1326 7430 1330 7548
rect 1350 7430 1354 7548
rect 1374 7430 1378 7548
rect 1398 7430 1402 7548
rect 1422 7430 1426 7548
rect 1446 7430 1450 7548
rect 1470 7430 1474 7548
rect 1494 7430 1498 7548
rect 1518 7430 1522 7548
rect 1542 7430 1546 7548
rect 1566 7430 1570 7548
rect 1590 7430 1594 7548
rect 1614 7430 1618 7548
rect 1638 7430 1642 7548
rect 1662 7430 1666 7548
rect 1686 7430 1690 7548
rect 1710 7430 1714 7548
rect 1734 7430 1738 7548
rect 1758 7430 1762 7548
rect 1782 7430 1786 7548
rect 1806 7430 1810 7548
rect 1830 7430 1834 7548
rect 1854 7430 1858 7548
rect 1878 7430 1882 7548
rect 1902 7430 1906 7548
rect 1926 7430 1930 7548
rect 1950 7430 1954 7548
rect 1974 7430 1978 7548
rect 1998 7430 2002 7548
rect 2022 7430 2026 7548
rect 2046 7430 2050 7548
rect 2070 7430 2074 7548
rect 2094 7430 2098 7548
rect 2118 7430 2122 7548
rect 2142 7430 2146 7548
rect 2166 7430 2170 7548
rect 2190 7430 2194 7548
rect 2214 7430 2218 7548
rect 2238 7430 2242 7548
rect 2262 7430 2266 7548
rect 2286 7430 2290 7548
rect 2310 7430 2314 7548
rect 2334 7430 2338 7548
rect 2358 7430 2362 7548
rect 2382 7430 2386 7548
rect 2406 7430 2410 7548
rect 2430 7430 2434 7548
rect 2454 7430 2458 7548
rect 2478 7430 2482 7548
rect 2502 7430 2506 7548
rect 2526 7430 2530 7548
rect 2550 7431 2554 7548
rect 2539 7430 2573 7431
rect 781 7428 2573 7430
rect 781 7427 795 7428
rect 798 7427 805 7428
rect 787 6845 792 6855
rect 798 6845 802 7427
rect 797 6831 802 6845
rect 787 6821 792 6831
rect 797 6807 802 6821
rect 798 6614 802 6807
rect 822 6779 826 7428
rect 822 6731 829 6779
rect 822 6614 826 6731
rect 846 6614 850 7428
rect 870 6614 874 7428
rect 894 6614 898 7428
rect 918 6614 922 7428
rect 942 6614 946 7428
rect 966 6614 970 7428
rect 990 6614 994 7428
rect 1014 6614 1018 7428
rect 1038 6614 1042 7428
rect 1062 6614 1066 7428
rect 1086 6614 1090 7428
rect 1110 6614 1114 7428
rect 1134 6614 1138 7428
rect 1158 6614 1162 7428
rect 1182 6614 1186 7428
rect 1206 6614 1210 7428
rect 1230 6614 1234 7428
rect 1254 6614 1258 7428
rect 1278 6614 1282 7428
rect 1302 6614 1306 7428
rect 1326 6614 1330 7428
rect 1350 6614 1354 7428
rect 1374 6614 1378 7428
rect 1398 6614 1402 7428
rect 1422 6614 1426 7428
rect 1446 6614 1450 7428
rect 1470 6614 1474 7428
rect 1494 6614 1498 7428
rect 1518 6614 1522 7428
rect 1542 6614 1546 7428
rect 1566 6614 1570 7428
rect 1590 6614 1594 7428
rect 1614 6614 1618 7428
rect 1638 6614 1642 7428
rect 1662 6614 1666 7428
rect 1686 6614 1690 7428
rect 1699 7349 1704 7359
rect 1710 7349 1714 7428
rect 1709 7335 1714 7349
rect 1710 6614 1714 7335
rect 1734 7283 1738 7428
rect 1734 7259 1741 7283
rect 1734 6614 1738 7259
rect 1758 6614 1762 7428
rect 1782 6614 1786 7428
rect 1806 6614 1810 7428
rect 1830 6614 1834 7428
rect 1854 6614 1858 7428
rect 1878 6614 1882 7428
rect 1902 6614 1906 7428
rect 1926 6614 1930 7428
rect 1950 6614 1954 7428
rect 1974 6614 1978 7428
rect 1998 6614 2002 7428
rect 2022 6614 2026 7428
rect 2046 6614 2050 7428
rect 2070 6614 2074 7428
rect 2094 6614 2098 7428
rect 2118 6614 2122 7428
rect 2142 6614 2146 7428
rect 2166 6614 2170 7428
rect 2190 6614 2194 7428
rect 2214 6614 2218 7428
rect 2238 6614 2242 7428
rect 2251 7061 2256 7071
rect 2262 7061 2266 7428
rect 2261 7047 2266 7061
rect 2262 6614 2266 7047
rect 2286 6995 2290 7428
rect 2286 6971 2293 6995
rect 2286 6614 2290 6971
rect 2310 6614 2314 7428
rect 2334 6614 2338 7428
rect 2358 6614 2362 7428
rect 2382 6614 2386 7428
rect 2406 6614 2410 7428
rect 2430 6614 2434 7428
rect 2454 6614 2458 7428
rect 2478 6614 2482 7428
rect 2502 6614 2506 7428
rect 2526 6614 2530 7428
rect 2539 7421 2544 7428
rect 2550 7421 2554 7428
rect 2549 7407 2554 7421
rect 2539 7205 2544 7215
rect 2550 7205 2554 7407
rect 2549 7191 2554 7205
rect 2539 6989 2544 6999
rect 2550 6989 2554 7191
rect 2549 6975 2554 6989
rect 2539 6773 2544 6783
rect 2550 6773 2554 6975
rect 2549 6759 2554 6773
rect 2550 6614 2554 6759
rect 2574 7355 2578 7548
rect 2574 7331 2581 7355
rect 2574 7139 2578 7331
rect 2574 7115 2581 7139
rect 2574 6923 2578 7115
rect 2574 6899 2581 6923
rect 2574 6707 2578 6899
rect 2587 6821 2592 6831
rect 2598 6821 2602 7548
rect 2611 7517 2616 7527
rect 2622 7517 2626 7548
rect 2635 7541 2640 7548
rect 2646 7541 2650 7548
rect 2645 7527 2650 7541
rect 2621 7503 2626 7517
rect 2597 6807 2602 6821
rect 2574 6683 2581 6707
rect 2587 6701 2592 6711
rect 2597 6687 2602 6701
rect 2574 6614 2578 6683
rect 2598 6615 2602 6687
rect 2587 6614 2619 6615
rect 667 6612 2619 6614
rect 667 6605 672 6612
rect 677 6591 682 6605
rect 667 6485 672 6495
rect 678 6485 682 6591
rect 677 6471 682 6485
rect 667 6269 672 6279
rect 678 6269 682 6471
rect 677 6255 682 6269
rect 678 6182 682 6255
rect 702 6563 706 6612
rect 702 6515 709 6563
rect 702 6419 706 6515
rect 702 6395 709 6419
rect 702 6203 706 6395
rect 331 6180 699 6182
rect 331 6173 336 6180
rect 341 6159 346 6173
rect 331 6125 336 6135
rect 342 6125 346 6159
rect 366 6131 370 6180
rect 341 6111 346 6125
rect 355 6121 363 6125
rect 349 6111 355 6121
rect 331 5909 336 5919
rect 342 5909 346 6111
rect 341 5895 346 5909
rect 331 5693 336 5703
rect 342 5693 346 5895
rect 341 5679 346 5693
rect 331 5477 336 5487
rect 342 5477 346 5679
rect 341 5463 346 5477
rect 331 5261 336 5271
rect 342 5261 346 5463
rect 341 5247 346 5261
rect 331 5045 336 5055
rect 342 5045 346 5247
rect 341 5031 346 5045
rect 342 4886 346 5031
rect 366 6083 373 6131
rect 366 6059 370 6083
rect 366 6035 373 6059
rect 366 5843 370 6035
rect 366 5819 373 5843
rect 366 5627 370 5819
rect 366 5603 373 5627
rect 366 5411 370 5603
rect 366 5387 373 5411
rect 366 5195 370 5387
rect 366 5171 373 5195
rect 366 4979 370 5171
rect 366 4955 373 4979
rect 366 4886 370 4955
rect 390 4886 394 6180
rect 414 4886 418 6180
rect 438 4886 442 6180
rect 462 4886 466 6180
rect 486 4886 490 6180
rect 510 4886 514 6180
rect 534 4886 538 6180
rect 558 4886 562 6180
rect 582 4886 586 6180
rect 606 4886 610 6180
rect 630 4886 634 6180
rect 654 4886 658 6180
rect 667 6053 672 6063
rect 678 6053 682 6180
rect 685 6179 699 6180
rect 702 6179 709 6203
rect 677 6039 682 6053
rect 667 5837 672 5847
rect 678 5837 682 6039
rect 677 5823 682 5837
rect 667 5621 672 5631
rect 678 5621 682 5823
rect 677 5607 682 5621
rect 667 5405 672 5415
rect 678 5405 682 5607
rect 677 5391 682 5405
rect 667 5189 672 5199
rect 678 5189 682 5391
rect 677 5175 682 5189
rect 667 4973 672 4983
rect 678 4973 682 5175
rect 677 4959 682 4973
rect 678 4886 682 4959
rect 702 5987 706 6179
rect 702 5963 709 5987
rect 702 5771 706 5963
rect 702 5747 709 5771
rect 702 5555 706 5747
rect 702 5531 709 5555
rect 702 5339 706 5531
rect 702 5315 709 5339
rect 702 5123 706 5315
rect 702 5099 709 5123
rect 702 4907 706 5099
rect -1277 4884 699 4886
rect -1277 4877 -1272 4884
rect -1267 4863 -1262 4877
rect -1266 4670 -1262 4863
rect -1242 4835 -1238 4884
rect -1242 4787 -1235 4835
rect -1242 4670 -1238 4787
rect -1218 4670 -1214 4884
rect -1194 4670 -1190 4884
rect -1170 4670 -1166 4884
rect -1146 4670 -1142 4884
rect -1122 4670 -1118 4884
rect -1098 4670 -1094 4884
rect -1074 4670 -1070 4884
rect -1050 4670 -1046 4884
rect -1026 4670 -1022 4884
rect -1002 4670 -998 4884
rect -978 4670 -974 4884
rect -954 4670 -950 4884
rect -930 4670 -926 4884
rect -906 4670 -902 4884
rect -882 4670 -878 4884
rect -858 4670 -854 4884
rect -834 4670 -830 4884
rect -810 4670 -806 4884
rect -786 4670 -782 4884
rect -762 4670 -758 4884
rect -738 4670 -734 4884
rect -714 4670 -710 4884
rect -690 4670 -686 4884
rect -666 4670 -662 4884
rect -642 4670 -638 4884
rect -618 4670 -614 4884
rect -594 4670 -590 4884
rect -570 4670 -566 4884
rect -546 4670 -542 4884
rect -522 4670 -518 4884
rect -498 4670 -494 4884
rect -474 4670 -470 4884
rect -450 4670 -446 4884
rect -426 4670 -422 4884
rect -402 4670 -398 4884
rect -378 4670 -374 4884
rect -354 4670 -350 4884
rect -330 4670 -326 4884
rect -306 4670 -302 4884
rect -282 4670 -278 4884
rect -258 4670 -254 4884
rect -234 4670 -230 4884
rect -210 4670 -206 4884
rect -186 4670 -182 4884
rect -162 4670 -158 4884
rect -138 4670 -134 4884
rect -114 4670 -110 4884
rect -101 4685 -96 4695
rect -90 4685 -86 4884
rect -91 4671 -86 4685
rect -90 4670 -86 4671
rect -66 4670 -62 4884
rect -42 4670 -38 4884
rect -18 4670 -14 4884
rect 6 4670 10 4884
rect 30 4670 34 4884
rect 54 4670 58 4884
rect 78 4670 82 4884
rect 102 4670 106 4884
rect 126 4670 130 4884
rect 150 4670 154 4884
rect 174 4670 178 4884
rect 198 4670 202 4884
rect 222 4670 226 4884
rect 246 4670 250 4884
rect 270 4670 274 4884
rect 294 4670 298 4884
rect 318 4670 322 4884
rect 331 4829 336 4839
rect 342 4829 346 4884
rect 341 4815 346 4829
rect 342 4670 346 4815
rect 366 4763 370 4884
rect 366 4739 373 4763
rect 366 4670 370 4739
rect 390 4670 394 4884
rect 414 4670 418 4884
rect 438 4670 442 4884
rect 462 4670 466 4884
rect 486 4670 490 4884
rect 510 4670 514 4884
rect 534 4670 538 4884
rect 558 4670 562 4884
rect 582 4670 586 4884
rect 606 4670 610 4884
rect 630 4670 634 4884
rect 654 4670 658 4884
rect 667 4757 672 4767
rect 678 4757 682 4884
rect 685 4883 699 4884
rect 702 4883 709 4907
rect 677 4743 682 4757
rect 678 4670 682 4743
rect 702 4691 706 4883
rect -2393 4668 -2018 4670
rect -2002 4668 699 4670
rect -2371 4574 -2366 4668
rect -2348 4574 -2343 4668
rect -2325 4666 -2320 4668
rect -2309 4666 -2301 4668
rect -2325 4654 -2317 4666
rect -2081 4659 -2077 4667
rect -2068 4659 -2065 4668
rect -2058 4659 -2028 4662
rect -2325 4634 -2320 4654
rect -2317 4650 -2309 4654
rect -2325 4626 -2317 4634
rect -2060 4628 -2030 4631
rect -2325 4578 -2320 4626
rect -2317 4618 -2309 4626
rect -2060 4615 -2038 4626
rect -2033 4619 -2030 4628
rect -2028 4624 -2027 4628
rect -2068 4610 -2038 4613
rect -2325 4574 -2317 4578
rect -2000 4576 -1992 4668
rect -1655 4666 -1647 4668
rect -1972 4659 -1924 4662
rect -1902 4659 -1794 4663
rect -1671 4654 -1663 4666
rect -1663 4650 -1655 4654
rect -1912 4643 -1884 4645
rect -1852 4637 -1804 4641
rect -1844 4628 -1796 4631
rect -1671 4626 -1663 4634
rect -1844 4615 -1804 4626
rect -1663 4618 -1655 4626
rect -1852 4610 -1680 4614
rect -2000 4574 -1957 4576
rect -1671 4574 -1663 4578
rect -1642 4574 -1637 4668
rect -1619 4574 -1614 4668
rect -1530 4574 -1526 4668
rect -1506 4574 -1502 4668
rect -1482 4574 -1478 4668
rect -1458 4574 -1454 4668
rect -1434 4574 -1430 4668
rect -1410 4574 -1406 4668
rect -1386 4574 -1382 4668
rect -1362 4574 -1358 4668
rect -1338 4574 -1334 4668
rect -1314 4574 -1310 4668
rect -1290 4574 -1286 4668
rect -1266 4574 -1262 4668
rect -1242 4574 -1238 4668
rect -1218 4574 -1214 4668
rect -1194 4574 -1190 4668
rect -1170 4574 -1166 4668
rect -1146 4574 -1142 4668
rect -1122 4574 -1118 4668
rect -1098 4574 -1094 4668
rect -1074 4574 -1070 4668
rect -1050 4574 -1046 4668
rect -1026 4574 -1022 4668
rect -1002 4574 -998 4668
rect -978 4574 -974 4668
rect -954 4574 -950 4668
rect -930 4574 -926 4668
rect -906 4574 -902 4668
rect -882 4574 -878 4668
rect -858 4574 -854 4668
rect -834 4574 -830 4668
rect -810 4574 -806 4668
rect -786 4574 -782 4668
rect -762 4574 -758 4668
rect -738 4574 -734 4668
rect -714 4574 -710 4668
rect -690 4574 -686 4668
rect -666 4574 -662 4668
rect -642 4574 -638 4668
rect -618 4574 -614 4668
rect -594 4574 -590 4668
rect -570 4574 -566 4668
rect -546 4574 -542 4668
rect -522 4574 -518 4668
rect -498 4574 -494 4668
rect -474 4574 -470 4668
rect -450 4574 -446 4668
rect -426 4574 -422 4668
rect -402 4574 -398 4668
rect -378 4574 -374 4668
rect -354 4574 -350 4668
rect -330 4574 -326 4668
rect -306 4574 -302 4668
rect -282 4574 -278 4668
rect -269 4637 -264 4647
rect -258 4637 -254 4668
rect -259 4623 -254 4637
rect -269 4622 -235 4623
rect -234 4622 -230 4668
rect -210 4622 -206 4668
rect -186 4622 -182 4668
rect -162 4622 -158 4668
rect -138 4622 -134 4668
rect -114 4622 -110 4668
rect -90 4622 -86 4668
rect -66 4622 -62 4668
rect -42 4622 -38 4668
rect -18 4622 -14 4668
rect 6 4622 10 4668
rect 30 4622 34 4668
rect 54 4622 58 4668
rect 78 4622 82 4668
rect 102 4622 106 4668
rect 126 4622 130 4668
rect 150 4622 154 4668
rect 174 4622 178 4668
rect 198 4622 202 4668
rect 222 4622 226 4668
rect 246 4622 250 4668
rect 270 4622 274 4668
rect 294 4622 298 4668
rect 318 4622 322 4668
rect 342 4622 346 4668
rect 366 4622 370 4668
rect 390 4622 394 4668
rect 414 4622 418 4668
rect 438 4622 442 4668
rect 462 4622 466 4668
rect 486 4622 490 4668
rect 510 4622 514 4668
rect 534 4622 538 4668
rect 558 4622 562 4668
rect 582 4622 586 4668
rect 606 4622 610 4668
rect 630 4622 634 4668
rect 654 4622 658 4668
rect 678 4622 682 4668
rect 685 4667 699 4668
rect 702 4667 709 4691
rect 702 4622 706 4667
rect 726 4622 730 6612
rect 750 4622 754 6612
rect 774 4622 778 6612
rect 798 4622 802 6612
rect 822 4622 826 6612
rect 846 4622 850 6612
rect 870 4622 874 6612
rect 894 4622 898 6612
rect 918 4622 922 6612
rect 931 5765 936 5775
rect 942 5765 946 6612
rect 941 5751 946 5765
rect 931 5741 936 5751
rect 941 5727 946 5741
rect 942 4622 946 5727
rect 966 5699 970 6612
rect 966 5651 973 5699
rect 966 4622 970 5651
rect 979 4661 984 4671
rect 990 4661 994 6612
rect 989 4647 994 4661
rect 979 4637 984 4647
rect 989 4623 994 4637
rect 990 4622 994 4623
rect 1014 4622 1018 6612
rect 1038 4622 1042 6612
rect 1062 4622 1066 6612
rect 1086 4622 1090 6612
rect 1110 4622 1114 6612
rect 1134 4622 1138 6612
rect 1158 4622 1162 6612
rect 1182 4622 1186 6612
rect 1206 4622 1210 6612
rect 1230 4622 1234 6612
rect 1254 4622 1258 6612
rect 1267 5549 1272 5559
rect 1278 5549 1282 6612
rect 1277 5535 1282 5549
rect 1267 5525 1272 5535
rect 1277 5511 1282 5525
rect 1278 4622 1282 5511
rect 1302 5483 1306 6612
rect 1302 5435 1309 5483
rect 1302 4622 1306 5435
rect 1326 4622 1330 6612
rect 1339 5333 1344 5343
rect 1350 5333 1354 6612
rect 1363 5981 1368 5991
rect 1374 5981 1378 6612
rect 1373 5967 1378 5981
rect 1363 5957 1368 5967
rect 1373 5943 1378 5957
rect 1349 5319 1354 5333
rect 1339 5309 1344 5319
rect 1349 5295 1354 5309
rect 1350 4622 1354 5295
rect 1374 5267 1378 5943
rect 1398 5915 1402 6612
rect 1398 5867 1405 5915
rect 1374 5219 1381 5267
rect 1374 4622 1378 5219
rect 1398 4622 1402 5867
rect 1422 4622 1426 6612
rect 1446 4622 1450 6612
rect 1459 6413 1464 6423
rect 1470 6413 1474 6612
rect 1469 6399 1474 6413
rect 1459 6389 1464 6399
rect 1469 6375 1474 6389
rect 1470 4622 1474 6375
rect 1494 6347 1498 6612
rect 1494 6299 1501 6347
rect 1494 4622 1498 6299
rect 1518 4622 1522 6612
rect 1542 4622 1546 6612
rect 1566 4622 1570 6612
rect 1590 4622 1594 6612
rect 1614 4622 1618 6612
rect 1638 4622 1642 6612
rect 1662 4622 1666 6612
rect 1686 4622 1690 6612
rect 1710 4622 1714 6612
rect 1734 4622 1738 6612
rect 1758 4622 1762 6612
rect 1782 4622 1786 6612
rect 1806 4622 1810 6612
rect 1830 4622 1834 6612
rect 1854 4622 1858 6612
rect 1878 4622 1882 6612
rect 1902 4622 1906 6612
rect 1926 4622 1930 6612
rect 1950 4622 1954 6612
rect 1974 4622 1978 6612
rect 1987 5117 1992 5127
rect 1998 5117 2002 6612
rect 1997 5103 2002 5117
rect 1987 5093 1992 5103
rect 1997 5079 2002 5093
rect 1998 4622 2002 5079
rect 2022 5051 2026 6612
rect 2022 5003 2029 5051
rect 2022 4622 2026 5003
rect 2046 4622 2050 6612
rect 2070 4622 2074 6612
rect 2094 4622 2098 6612
rect 2118 4622 2122 6612
rect 2142 4622 2146 6612
rect 2166 4622 2170 6612
rect 2190 4622 2194 6612
rect 2214 4622 2218 6612
rect 2238 4622 2242 6612
rect 2262 4622 2266 6612
rect 2286 4622 2290 6612
rect 2310 4622 2314 6612
rect 2334 4622 2338 6612
rect 2358 4622 2362 6612
rect 2382 4623 2386 6612
rect 2395 4877 2400 4887
rect 2406 4877 2410 6612
rect 2419 5093 2424 5103
rect 2430 5093 2434 6612
rect 2443 5309 2448 5319
rect 2454 5309 2458 6612
rect 2467 5525 2472 5535
rect 2478 5525 2482 6612
rect 2491 5741 2496 5751
rect 2502 5741 2506 6612
rect 2515 5957 2520 5967
rect 2526 5957 2530 6612
rect 2539 6557 2544 6567
rect 2550 6557 2554 6612
rect 2549 6543 2554 6557
rect 2539 6341 2544 6351
rect 2550 6341 2554 6543
rect 2574 6491 2578 6612
rect 2587 6605 2592 6612
rect 2598 6605 2602 6612
rect 2605 6611 2619 6612
rect 2597 6591 2602 6605
rect 2574 6467 2581 6491
rect 2563 6389 2568 6399
rect 2574 6389 2578 6467
rect 2573 6375 2578 6389
rect 2549 6327 2554 6341
rect 2539 6173 2544 6183
rect 2550 6173 2554 6327
rect 2549 6159 2554 6173
rect 2525 5943 2530 5957
rect 2501 5727 2506 5741
rect 2477 5511 2482 5525
rect 2453 5295 2458 5309
rect 2429 5079 2434 5093
rect 2405 4863 2410 4877
rect 2395 4709 2400 4719
rect 2405 4695 2410 4709
rect 2395 4637 2400 4647
rect 2406 4637 2410 4695
rect 2405 4623 2410 4637
rect 2419 4633 2427 4637
rect 2413 4623 2419 4633
rect 2371 4622 2405 4623
rect -269 4620 2405 4622
rect -269 4613 -264 4620
rect -259 4599 -254 4613
rect -258 4574 -254 4599
rect -234 4574 -230 4620
rect -210 4574 -206 4620
rect -186 4574 -182 4620
rect -162 4574 -158 4620
rect -138 4574 -134 4620
rect -114 4574 -110 4620
rect -90 4574 -86 4620
rect -66 4619 -62 4620
rect -66 4595 -59 4619
rect -66 4574 -62 4595
rect -42 4574 -38 4620
rect -18 4574 -14 4620
rect 6 4574 10 4620
rect 30 4574 34 4620
rect 54 4574 58 4620
rect 78 4574 82 4620
rect 102 4574 106 4620
rect 126 4574 130 4620
rect 150 4574 154 4620
rect 174 4574 178 4620
rect 198 4574 202 4620
rect 222 4574 226 4620
rect 246 4574 250 4620
rect 270 4574 274 4620
rect 294 4574 298 4620
rect 318 4574 322 4620
rect 342 4574 346 4620
rect 366 4574 370 4620
rect 390 4574 394 4620
rect 414 4574 418 4620
rect 438 4574 442 4620
rect 462 4574 466 4620
rect 486 4574 490 4620
rect 510 4574 514 4620
rect 534 4574 538 4620
rect 558 4574 562 4620
rect 582 4574 586 4620
rect 606 4574 610 4620
rect 630 4574 634 4620
rect 654 4574 658 4620
rect 678 4574 682 4620
rect 702 4574 706 4620
rect 726 4574 730 4620
rect 750 4574 754 4620
rect 774 4574 778 4620
rect 798 4574 802 4620
rect 822 4574 826 4620
rect 846 4574 850 4620
rect 870 4574 874 4620
rect 894 4574 898 4620
rect 918 4574 922 4620
rect 942 4574 946 4620
rect 966 4574 970 4620
rect 990 4574 994 4620
rect 1014 4595 1018 4620
rect -2393 4572 1011 4574
rect -2371 4334 -2366 4572
rect -2348 4334 -2343 4572
rect -2325 4550 -2320 4572
rect -2317 4562 -2309 4572
rect -2325 4546 -2317 4550
rect -2325 4498 -2320 4546
rect -2317 4534 -2309 4546
rect -2163 4534 -2127 4537
rect -2124 4534 -2108 4538
rect -2060 4534 -2030 4538
rect -2325 4490 -2317 4498
rect -2325 4470 -2320 4490
rect -2317 4482 -2309 4490
rect -2325 4462 -2317 4470
rect -2325 4442 -2320 4462
rect -2317 4454 -2309 4462
rect -2127 4450 -2097 4451
rect -2325 4434 -2317 4442
rect -2325 4414 -2320 4434
rect -2317 4427 -2309 4434
rect -2127 4430 -2124 4439
rect -2119 4430 -2097 4443
rect -2092 4437 -2089 4443
rect -2087 4440 -2079 4453
rect -2127 4429 -2097 4430
rect -2317 4426 -2301 4427
rect -2309 4415 -2307 4426
rect -2145 4418 -2129 4425
rect -2066 4424 -2065 4425
rect -2325 4406 -2317 4414
rect -2325 4386 -2320 4406
rect -2317 4398 -2309 4406
rect -2297 4399 -2289 4415
rect -2150 4413 -2141 4415
rect -2129 4413 -2113 4415
rect -2119 4404 -2113 4413
rect -2125 4399 -2113 4404
rect -2101 4411 -2085 4415
rect -2101 4399 -2089 4411
rect -2325 4374 -2317 4386
rect -2325 4358 -2320 4374
rect -2317 4370 -2309 4374
rect -2068 4370 -2038 4371
rect -2309 4358 -2301 4370
rect -2068 4366 -2063 4370
rect -2000 4366 -1992 4572
rect -1972 4570 -1957 4572
rect -1958 4569 -1957 4570
rect -1984 4548 -1980 4566
rect -1663 4562 -1655 4572
rect -1832 4561 -1796 4562
rect -1824 4552 -1796 4554
rect -1954 4548 -1918 4552
rect -1796 4551 -1788 4552
rect -1822 4538 -1796 4550
rect -1671 4546 -1663 4550
rect -1857 4528 -1850 4538
rect -1844 4534 -1796 4538
rect -1663 4534 -1655 4546
rect -1847 4525 -1840 4528
rect -1671 4490 -1663 4498
rect -1663 4482 -1655 4490
rect -1946 4468 -1893 4476
rect -1927 4458 -1919 4466
rect -1901 4458 -1898 4468
rect -1671 4462 -1663 4470
rect -1927 4452 -1920 4458
rect -1936 4450 -1920 4452
rect -1919 4457 -1911 4458
rect -1919 4450 -1903 4457
rect -1901 4451 -1900 4458
rect -1663 4454 -1655 4462
rect -1901 4450 -1853 4451
rect -1893 4430 -1853 4443
rect -1671 4434 -1663 4442
rect -1901 4429 -1853 4430
rect -1663 4426 -1655 4434
rect -1915 4418 -1914 4425
rect -1767 4418 -1766 4425
rect -1671 4406 -1663 4414
rect -1663 4398 -1655 4406
rect -2325 4346 -2317 4358
rect -2058 4355 -2038 4366
rect -2028 4362 -1992 4366
rect -1916 4365 -1903 4375
rect -1671 4374 -1663 4386
rect -1852 4370 -1832 4371
rect -1663 4370 -1655 4374
rect -2068 4346 -2065 4351
rect -2058 4350 -2028 4353
rect -2011 4352 -2002 4356
rect -2000 4352 -1992 4362
rect -1893 4354 -1892 4361
rect -1852 4355 -1845 4370
rect -1655 4358 -1647 4370
rect -1854 4354 -1845 4355
rect -1893 4353 -1680 4354
rect -2001 4350 -1992 4352
rect -2038 4348 -2028 4350
rect -2058 4346 -2038 4348
rect -2325 4334 -2320 4346
rect -2317 4342 -2309 4346
rect -2309 4334 -2301 4342
rect -2068 4341 -2058 4346
rect -2068 4334 -2065 4341
rect -2016 4340 -2002 4350
rect -2000 4341 -1992 4350
rect -1972 4348 -1924 4353
rect -1671 4346 -1663 4358
rect -1663 4342 -1655 4346
rect -2001 4340 -1992 4341
rect -2015 4336 -2002 4340
rect -2000 4334 -1992 4340
rect -1976 4334 -1940 4335
rect -1655 4334 -1647 4342
rect -1642 4334 -1637 4572
rect -1619 4334 -1614 4572
rect -1530 4334 -1526 4572
rect -1506 4334 -1502 4572
rect -1482 4334 -1478 4572
rect -1458 4334 -1454 4572
rect -1434 4334 -1430 4572
rect -1410 4335 -1406 4572
rect -1421 4334 -1387 4335
rect -2393 4332 -2018 4334
rect -2002 4332 -1387 4334
rect -2371 4262 -2366 4332
rect -2348 4262 -2343 4332
rect -2325 4330 -2320 4332
rect -2309 4330 -2301 4332
rect -2325 4318 -2317 4330
rect -2081 4323 -2077 4331
rect -2068 4323 -2065 4332
rect -2058 4323 -2028 4326
rect -2325 4298 -2320 4318
rect -2317 4314 -2309 4318
rect -2325 4290 -2317 4298
rect -2060 4292 -2030 4295
rect -2325 4262 -2320 4290
rect -2317 4282 -2309 4290
rect -2060 4279 -2038 4290
rect -2033 4283 -2030 4292
rect -2028 4288 -2027 4292
rect -2068 4274 -2038 4277
rect -2000 4262 -1992 4332
rect -1655 4330 -1647 4332
rect -1972 4323 -1924 4326
rect -1902 4323 -1794 4327
rect -1671 4318 -1663 4330
rect -1663 4314 -1655 4318
rect -1912 4307 -1884 4309
rect -1852 4301 -1804 4305
rect -1844 4292 -1796 4295
rect -1671 4290 -1663 4298
rect -1844 4279 -1804 4290
rect -1663 4282 -1655 4290
rect -1852 4274 -1680 4278
rect -1642 4262 -1637 4332
rect -1619 4262 -1614 4332
rect -1530 4262 -1526 4332
rect -1506 4262 -1502 4332
rect -1482 4262 -1478 4332
rect -1458 4262 -1454 4332
rect -1434 4262 -1430 4332
rect -1421 4325 -1416 4332
rect -1410 4325 -1406 4332
rect -1411 4311 -1406 4325
rect -1421 4286 -1387 4287
rect -1386 4286 -1382 4572
rect -1362 4286 -1358 4572
rect -1338 4286 -1334 4572
rect -1314 4286 -1310 4572
rect -1290 4286 -1286 4572
rect -1266 4286 -1262 4572
rect -1242 4286 -1238 4572
rect -1218 4286 -1214 4572
rect -1194 4286 -1190 4572
rect -1170 4286 -1166 4572
rect -1146 4286 -1142 4572
rect -1122 4286 -1118 4572
rect -1098 4286 -1094 4572
rect -1074 4286 -1070 4572
rect -1050 4286 -1046 4572
rect -1026 4286 -1022 4572
rect -1002 4286 -998 4572
rect -978 4286 -974 4572
rect -954 4286 -950 4572
rect -930 4286 -926 4572
rect -906 4286 -902 4572
rect -882 4286 -878 4572
rect -858 4286 -854 4572
rect -834 4286 -830 4572
rect -810 4286 -806 4572
rect -786 4286 -782 4572
rect -762 4286 -758 4572
rect -738 4286 -734 4572
rect -714 4286 -710 4572
rect -690 4286 -686 4572
rect -666 4286 -662 4572
rect -642 4286 -638 4572
rect -618 4286 -614 4572
rect -594 4286 -590 4572
rect -570 4286 -566 4572
rect -546 4286 -542 4572
rect -522 4286 -518 4572
rect -498 4286 -494 4572
rect -474 4286 -470 4572
rect -450 4286 -446 4572
rect -426 4286 -422 4572
rect -402 4286 -398 4572
rect -378 4286 -374 4572
rect -354 4286 -350 4572
rect -330 4286 -326 4572
rect -306 4286 -302 4572
rect -282 4286 -278 4572
rect -258 4286 -254 4572
rect -234 4571 -230 4572
rect -234 4523 -227 4571
rect -234 4286 -230 4523
rect -210 4286 -206 4572
rect -186 4286 -182 4572
rect -162 4286 -158 4572
rect -138 4286 -134 4572
rect -114 4286 -110 4572
rect -90 4286 -86 4572
rect -66 4286 -62 4572
rect -42 4286 -38 4572
rect -18 4286 -14 4572
rect 6 4286 10 4572
rect 30 4286 34 4572
rect 54 4286 58 4572
rect 78 4286 82 4572
rect 102 4286 106 4572
rect 126 4286 130 4572
rect 150 4286 154 4572
rect 174 4286 178 4572
rect 198 4286 202 4572
rect 222 4286 226 4572
rect 246 4286 250 4572
rect 270 4286 274 4572
rect 294 4286 298 4572
rect 318 4286 322 4572
rect 331 4493 336 4503
rect 342 4493 346 4572
rect 341 4479 346 4493
rect 342 4286 346 4479
rect 366 4427 370 4572
rect 366 4403 373 4427
rect 366 4286 370 4403
rect 390 4286 394 4572
rect 414 4286 418 4572
rect 438 4286 442 4572
rect 462 4286 466 4572
rect 486 4286 490 4572
rect 510 4286 514 4572
rect 534 4286 538 4572
rect 558 4286 562 4572
rect 582 4286 586 4572
rect 595 4301 600 4311
rect 606 4301 610 4572
rect 605 4287 610 4301
rect 630 4286 634 4572
rect 654 4286 658 4572
rect 667 4421 672 4431
rect 678 4421 682 4572
rect 677 4407 682 4421
rect 678 4286 682 4407
rect 702 4355 706 4572
rect 702 4331 709 4355
rect 702 4286 706 4331
rect 726 4286 730 4572
rect 750 4286 754 4572
rect 774 4286 778 4572
rect 798 4286 802 4572
rect 822 4286 826 4572
rect 846 4286 850 4572
rect 870 4286 874 4572
rect 894 4286 898 4572
rect 918 4286 922 4572
rect 942 4286 946 4572
rect 966 4286 970 4572
rect 990 4286 994 4572
rect 997 4571 1011 4572
rect 1014 4547 1021 4595
rect 1014 4286 1018 4547
rect 1038 4286 1042 4620
rect 1062 4286 1066 4620
rect 1086 4286 1090 4620
rect 1110 4286 1114 4620
rect 1134 4286 1138 4620
rect 1158 4286 1162 4620
rect 1182 4286 1186 4620
rect 1206 4286 1210 4620
rect 1230 4286 1234 4620
rect 1254 4286 1258 4620
rect 1278 4286 1282 4620
rect 1302 4286 1306 4620
rect 1326 4286 1330 4620
rect 1350 4286 1354 4620
rect 1374 4286 1378 4620
rect 1398 4286 1402 4620
rect 1422 4286 1426 4620
rect 1446 4286 1450 4620
rect 1470 4286 1474 4620
rect 1494 4286 1498 4620
rect 1518 4286 1522 4620
rect 1542 4286 1546 4620
rect 1566 4286 1570 4620
rect 1590 4286 1594 4620
rect 1614 4286 1618 4620
rect 1638 4286 1642 4620
rect 1651 4349 1656 4359
rect 1662 4349 1666 4620
rect 1661 4335 1666 4349
rect 1651 4325 1656 4335
rect 1661 4311 1666 4325
rect 1662 4286 1666 4311
rect 1686 4286 1690 4620
rect 1710 4286 1714 4620
rect 1734 4286 1738 4620
rect 1758 4286 1762 4620
rect 1782 4286 1786 4620
rect 1806 4286 1810 4620
rect 1830 4286 1834 4620
rect 1854 4286 1858 4620
rect 1878 4286 1882 4620
rect 1902 4286 1906 4620
rect 1926 4286 1930 4620
rect 1950 4286 1954 4620
rect 1974 4286 1978 4620
rect 1998 4286 2002 4620
rect 2022 4286 2026 4620
rect 2046 4286 2050 4620
rect 2070 4286 2074 4620
rect 2094 4286 2098 4620
rect 2118 4286 2122 4620
rect 2142 4286 2146 4620
rect 2166 4286 2170 4620
rect 2190 4286 2194 4620
rect 2214 4286 2218 4620
rect 2238 4286 2242 4620
rect 2262 4286 2266 4620
rect 2286 4286 2290 4620
rect 2310 4286 2314 4620
rect 2334 4287 2338 4620
rect 2347 4565 2352 4575
rect 2358 4565 2362 4620
rect 2371 4613 2376 4620
rect 2382 4613 2386 4620
rect 2381 4599 2386 4613
rect 2357 4551 2362 4565
rect 2347 4373 2352 4383
rect 2357 4359 2362 4373
rect 2347 4325 2352 4335
rect 2358 4325 2362 4359
rect 2357 4311 2362 4325
rect 2323 4286 2357 4287
rect -1421 4284 2357 4286
rect -1421 4277 -1416 4284
rect -1411 4263 -1406 4277
rect -1410 4262 -1406 4263
rect -1386 4262 -1382 4284
rect -1362 4262 -1358 4284
rect -1338 4262 -1334 4284
rect -1314 4262 -1310 4284
rect -1290 4262 -1286 4284
rect -1266 4262 -1262 4284
rect -1242 4262 -1238 4284
rect -1218 4262 -1214 4284
rect -1194 4262 -1190 4284
rect -1170 4262 -1166 4284
rect -1146 4262 -1142 4284
rect -1122 4262 -1118 4284
rect -1098 4262 -1094 4284
rect -1074 4262 -1070 4284
rect -1050 4262 -1046 4284
rect -1026 4262 -1022 4284
rect -1002 4262 -998 4284
rect -978 4262 -974 4284
rect -954 4262 -950 4284
rect -930 4262 -926 4284
rect -906 4262 -902 4284
rect -882 4262 -878 4284
rect -858 4262 -854 4284
rect -834 4262 -830 4284
rect -810 4262 -806 4284
rect -786 4262 -782 4284
rect -762 4262 -758 4284
rect -738 4262 -734 4284
rect -714 4262 -710 4284
rect -690 4262 -686 4284
rect -666 4262 -662 4284
rect -642 4262 -638 4284
rect -618 4262 -614 4284
rect -594 4262 -590 4284
rect -570 4262 -566 4284
rect -546 4262 -542 4284
rect -522 4262 -518 4284
rect -498 4262 -494 4284
rect -474 4262 -470 4284
rect -450 4262 -446 4284
rect -426 4262 -422 4284
rect -402 4262 -398 4284
rect -378 4262 -374 4284
rect -354 4262 -350 4284
rect -330 4262 -326 4284
rect -306 4262 -302 4284
rect -282 4262 -278 4284
rect -258 4262 -254 4284
rect -234 4262 -230 4284
rect -210 4262 -206 4284
rect -186 4262 -182 4284
rect -162 4262 -158 4284
rect -138 4262 -134 4284
rect -114 4262 -110 4284
rect -90 4262 -86 4284
rect -66 4262 -62 4284
rect -42 4262 -38 4284
rect -18 4262 -14 4284
rect 6 4262 10 4284
rect 30 4262 34 4284
rect 54 4262 58 4284
rect 78 4262 82 4284
rect 102 4262 106 4284
rect 126 4262 130 4284
rect 150 4262 154 4284
rect 174 4262 178 4284
rect 198 4262 202 4284
rect 222 4262 226 4284
rect 246 4262 250 4284
rect 270 4262 274 4284
rect 294 4262 298 4284
rect 318 4262 322 4284
rect 342 4262 346 4284
rect 366 4262 370 4284
rect 390 4262 394 4284
rect 414 4262 418 4284
rect 438 4262 442 4284
rect 462 4262 466 4284
rect 486 4262 490 4284
rect 510 4262 514 4284
rect 534 4262 538 4284
rect 558 4262 562 4284
rect 582 4262 586 4284
rect 595 4262 629 4263
rect -2393 4260 629 4262
rect -2371 4238 -2366 4260
rect -2348 4238 -2343 4260
rect -2325 4238 -2320 4260
rect -2309 4242 -2301 4252
rect -2068 4243 -2062 4248
rect -2317 4238 -2309 4242
rect -2060 4238 -2050 4243
rect -2000 4238 -1992 4260
rect -1806 4252 -1680 4258
rect -1854 4243 -1806 4248
rect -1655 4242 -1647 4252
rect -1972 4238 -1964 4239
rect -1958 4238 -1942 4240
rect -1844 4238 -1806 4241
rect -1663 4238 -1655 4242
rect -1642 4238 -1637 4260
rect -1619 4238 -1614 4260
rect -1530 4238 -1526 4260
rect -1506 4238 -1502 4260
rect -1482 4238 -1478 4260
rect -1458 4238 -1454 4260
rect -1434 4238 -1430 4260
rect -1410 4238 -1406 4260
rect -1386 4259 -1382 4260
rect -2393 4236 -1389 4238
rect -2371 4214 -2366 4236
rect -2348 4214 -2343 4236
rect -2325 4214 -2320 4236
rect -2060 4230 -2050 4236
rect -2309 4214 -2301 4224
rect -2060 4223 -2030 4230
rect -2000 4226 -1992 4236
rect -1972 4234 -1942 4236
rect -1958 4233 -1942 4234
rect -1844 4232 -1806 4236
rect -2068 4216 -2062 4223
rect -2062 4214 -2036 4216
rect -2393 4212 -2036 4214
rect -2030 4214 -2012 4216
rect -2004 4214 -1990 4226
rect -1844 4225 -1798 4230
rect -1806 4223 -1798 4225
rect -1854 4221 -1844 4223
rect -1854 4216 -1806 4221
rect -1864 4214 -1796 4215
rect -1655 4214 -1647 4224
rect -1642 4214 -1637 4236
rect -1619 4214 -1614 4236
rect -1530 4214 -1526 4236
rect -1506 4214 -1502 4236
rect -1482 4214 -1478 4236
rect -1458 4214 -1454 4236
rect -1434 4214 -1430 4236
rect -1410 4214 -1406 4236
rect -1403 4235 -1389 4236
rect -1386 4235 -1379 4259
rect -1362 4214 -1358 4260
rect -1338 4214 -1334 4260
rect -1314 4214 -1310 4260
rect -1290 4214 -1286 4260
rect -1277 4229 -1272 4239
rect -1266 4229 -1262 4260
rect -1267 4215 -1262 4229
rect -1277 4214 -1243 4215
rect -1242 4214 -1238 4260
rect -1218 4214 -1214 4260
rect -1194 4214 -1190 4260
rect -1170 4214 -1166 4260
rect -1146 4214 -1142 4260
rect -1122 4214 -1118 4260
rect -1098 4214 -1094 4260
rect -1074 4214 -1070 4260
rect -1050 4214 -1046 4260
rect -1026 4214 -1022 4260
rect -1002 4214 -998 4260
rect -978 4214 -974 4260
rect -954 4214 -950 4260
rect -930 4214 -926 4260
rect -906 4214 -902 4260
rect -882 4214 -878 4260
rect -858 4215 -854 4260
rect -869 4214 -835 4215
rect -2030 4212 -835 4214
rect -2371 4166 -2366 4212
rect -2348 4166 -2343 4212
rect -2325 4166 -2320 4212
rect -2317 4208 -2309 4212
rect -2060 4208 -2050 4212
rect -2060 4206 -2036 4208
rect -2060 4204 -2030 4206
rect -2292 4198 -2030 4204
rect -2092 4182 -2062 4184
rect -2094 4178 -2062 4182
rect -2000 4166 -1992 4212
rect -1844 4205 -1806 4212
rect -1663 4208 -1655 4212
rect -1844 4198 -1680 4204
rect -1854 4182 -1806 4184
rect -1854 4178 -1680 4182
rect -1642 4166 -1637 4212
rect -1619 4166 -1614 4212
rect -1530 4166 -1526 4212
rect -1506 4166 -1502 4212
rect -1482 4166 -1478 4212
rect -1458 4166 -1454 4212
rect -1434 4166 -1430 4212
rect -1410 4166 -1406 4212
rect -1386 4187 -1379 4211
rect -1386 4166 -1382 4187
rect -1362 4166 -1358 4212
rect -1338 4166 -1334 4212
rect -1314 4166 -1310 4212
rect -1290 4166 -1286 4212
rect -1277 4205 -1272 4212
rect -1267 4191 -1262 4205
rect -1266 4166 -1262 4191
rect -1242 4166 -1238 4212
rect -1218 4166 -1214 4212
rect -1194 4166 -1190 4212
rect -1170 4166 -1166 4212
rect -1146 4166 -1142 4212
rect -1122 4166 -1118 4212
rect -1098 4166 -1094 4212
rect -1074 4166 -1070 4212
rect -1050 4166 -1046 4212
rect -1026 4166 -1022 4212
rect -1002 4166 -998 4212
rect -978 4166 -974 4212
rect -954 4166 -950 4212
rect -930 4166 -926 4212
rect -906 4166 -902 4212
rect -882 4166 -878 4212
rect -869 4205 -864 4212
rect -858 4205 -854 4212
rect -859 4191 -854 4205
rect -869 4190 -835 4191
rect -834 4190 -830 4260
rect -810 4190 -806 4260
rect -786 4190 -782 4260
rect -762 4190 -758 4260
rect -738 4190 -734 4260
rect -714 4190 -710 4260
rect -690 4190 -686 4260
rect -666 4190 -662 4260
rect -642 4190 -638 4260
rect -618 4190 -614 4260
rect -594 4190 -590 4260
rect -570 4190 -566 4260
rect -546 4190 -542 4260
rect -522 4190 -518 4260
rect -498 4190 -494 4260
rect -474 4190 -470 4260
rect -450 4190 -446 4260
rect -426 4190 -422 4260
rect -402 4190 -398 4260
rect -378 4190 -374 4260
rect -354 4190 -350 4260
rect -330 4190 -326 4260
rect -306 4190 -302 4260
rect -282 4190 -278 4260
rect -258 4190 -254 4260
rect -234 4190 -230 4260
rect -210 4190 -206 4260
rect -186 4190 -182 4260
rect -162 4190 -158 4260
rect -138 4190 -134 4260
rect -114 4190 -110 4260
rect -90 4190 -86 4260
rect -66 4190 -62 4260
rect -42 4190 -38 4260
rect -18 4190 -14 4260
rect 6 4190 10 4260
rect 30 4190 34 4260
rect 54 4190 58 4260
rect 78 4190 82 4260
rect 102 4190 106 4260
rect 126 4190 130 4260
rect 150 4190 154 4260
rect 174 4190 178 4260
rect 198 4190 202 4260
rect 222 4190 226 4260
rect 246 4190 250 4260
rect 270 4190 274 4260
rect 294 4190 298 4260
rect 318 4190 322 4260
rect 342 4190 346 4260
rect 366 4190 370 4260
rect 390 4190 394 4260
rect 414 4190 418 4260
rect 438 4190 442 4260
rect 462 4190 466 4260
rect 486 4190 490 4260
rect 510 4190 514 4260
rect 534 4190 538 4260
rect 558 4190 562 4260
rect 582 4190 586 4260
rect 595 4253 600 4260
rect 605 4239 610 4253
rect 606 4190 610 4239
rect 630 4235 634 4284
rect 630 4211 637 4235
rect 654 4190 658 4284
rect 678 4190 682 4284
rect 702 4190 706 4284
rect 726 4190 730 4284
rect 750 4190 754 4284
rect 774 4190 778 4284
rect 798 4190 802 4284
rect 822 4190 826 4284
rect 846 4190 850 4284
rect 870 4190 874 4284
rect 894 4190 898 4284
rect 918 4190 922 4284
rect 942 4190 946 4284
rect 966 4190 970 4284
rect 990 4190 994 4284
rect 1014 4190 1018 4284
rect 1038 4190 1042 4284
rect 1062 4190 1066 4284
rect 1086 4190 1090 4284
rect 1110 4190 1114 4284
rect 1134 4190 1138 4284
rect 1158 4190 1162 4284
rect 1182 4190 1186 4284
rect 1206 4190 1210 4284
rect 1230 4190 1234 4284
rect 1254 4190 1258 4284
rect 1278 4190 1282 4284
rect 1302 4190 1306 4284
rect 1326 4190 1330 4284
rect 1350 4190 1354 4284
rect 1374 4190 1378 4284
rect 1398 4190 1402 4284
rect 1422 4190 1426 4284
rect 1446 4190 1450 4284
rect 1470 4190 1474 4284
rect 1494 4190 1498 4284
rect 1518 4190 1522 4284
rect 1542 4190 1546 4284
rect 1566 4190 1570 4284
rect 1590 4190 1594 4284
rect 1614 4190 1618 4284
rect 1638 4190 1642 4284
rect 1662 4190 1666 4284
rect 1686 4283 1690 4284
rect 1686 4235 1693 4283
rect 1686 4190 1690 4235
rect 1710 4190 1714 4284
rect 1734 4190 1738 4284
rect 1758 4190 1762 4284
rect 1782 4190 1786 4284
rect 1806 4190 1810 4284
rect 1830 4190 1834 4284
rect 1854 4190 1858 4284
rect 1878 4190 1882 4284
rect 1902 4190 1906 4284
rect 1926 4190 1930 4284
rect 1950 4190 1954 4284
rect 1974 4190 1978 4284
rect 1998 4190 2002 4284
rect 2022 4190 2026 4284
rect 2046 4190 2050 4284
rect 2070 4190 2074 4284
rect 2094 4190 2098 4284
rect 2118 4190 2122 4284
rect 2142 4190 2146 4284
rect 2166 4190 2170 4284
rect 2190 4190 2194 4284
rect 2214 4190 2218 4284
rect 2238 4190 2242 4284
rect 2262 4190 2266 4284
rect 2286 4190 2290 4284
rect 2310 4191 2314 4284
rect 2323 4277 2328 4284
rect 2334 4277 2338 4284
rect 2333 4263 2338 4277
rect 2299 4190 2333 4191
rect -869 4188 2333 4190
rect -869 4181 -864 4188
rect -859 4167 -854 4181
rect -858 4166 -854 4167
rect -834 4166 -830 4188
rect -810 4166 -806 4188
rect -786 4166 -782 4188
rect -762 4166 -758 4188
rect -738 4166 -734 4188
rect -714 4166 -710 4188
rect -690 4166 -686 4188
rect -666 4166 -662 4188
rect -642 4166 -638 4188
rect -618 4166 -614 4188
rect -594 4166 -590 4188
rect -570 4166 -566 4188
rect -546 4166 -542 4188
rect -522 4166 -518 4188
rect -498 4166 -494 4188
rect -474 4166 -470 4188
rect -450 4166 -446 4188
rect -426 4166 -422 4188
rect -402 4166 -398 4188
rect -378 4166 -374 4188
rect -354 4166 -350 4188
rect -330 4166 -326 4188
rect -306 4166 -302 4188
rect -282 4166 -278 4188
rect -258 4166 -254 4188
rect -234 4166 -230 4188
rect -210 4166 -206 4188
rect -186 4166 -182 4188
rect -162 4166 -158 4188
rect -138 4166 -134 4188
rect -114 4166 -110 4188
rect -90 4166 -86 4188
rect -66 4166 -62 4188
rect -42 4166 -38 4188
rect -18 4166 -14 4188
rect 6 4166 10 4188
rect 30 4166 34 4188
rect 54 4166 58 4188
rect 78 4166 82 4188
rect 102 4166 106 4188
rect 126 4166 130 4188
rect 150 4166 154 4188
rect 174 4166 178 4188
rect 198 4166 202 4188
rect 222 4166 226 4188
rect 246 4166 250 4188
rect 270 4166 274 4188
rect 294 4166 298 4188
rect 318 4166 322 4188
rect 342 4166 346 4188
rect 366 4166 370 4188
rect 390 4166 394 4188
rect 414 4166 418 4188
rect 438 4166 442 4188
rect 462 4166 466 4188
rect 486 4166 490 4188
rect 510 4166 514 4188
rect 534 4166 538 4188
rect 558 4166 562 4188
rect 582 4166 586 4188
rect 606 4166 610 4188
rect -2393 4164 627 4166
rect -2371 4142 -2366 4164
rect -2348 4142 -2343 4164
rect -2325 4142 -2320 4164
rect -2072 4162 -2036 4163
rect -2072 4156 -2054 4162
rect -2309 4148 -2301 4156
rect -2317 4142 -2309 4148
rect -2092 4147 -2062 4152
rect -2000 4143 -1992 4164
rect -1938 4163 -1906 4164
rect -1920 4162 -1906 4163
rect -1806 4156 -1680 4162
rect -1854 4147 -1806 4152
rect -1655 4148 -1647 4156
rect -1982 4143 -1966 4144
rect -2000 4142 -1966 4143
rect -1846 4142 -1806 4145
rect -1663 4142 -1655 4148
rect -1642 4142 -1637 4164
rect -1619 4142 -1614 4164
rect -1530 4142 -1526 4164
rect -1506 4142 -1502 4164
rect -1482 4142 -1478 4164
rect -1458 4142 -1454 4164
rect -1434 4142 -1430 4164
rect -1410 4142 -1406 4164
rect -1386 4143 -1382 4164
rect -1397 4142 -1363 4143
rect -2393 4140 -1363 4142
rect -2371 4118 -2366 4140
rect -2348 4118 -2343 4140
rect -2325 4118 -2320 4140
rect -2000 4138 -1966 4140
rect -2309 4120 -2301 4128
rect -2062 4127 -2054 4134
rect -2092 4120 -2084 4127
rect -2062 4120 -2026 4122
rect -2317 4118 -2309 4120
rect -2062 4118 -2012 4120
rect -2000 4118 -1992 4138
rect -1982 4137 -1966 4138
rect -1846 4136 -1806 4140
rect -1846 4129 -1798 4134
rect -1806 4127 -1798 4129
rect -1854 4125 -1846 4127
rect -1854 4120 -1806 4125
rect -1655 4120 -1647 4128
rect -1864 4118 -1796 4119
rect -1663 4118 -1655 4120
rect -1642 4118 -1637 4140
rect -1619 4118 -1614 4140
rect -1530 4118 -1526 4140
rect -1506 4118 -1502 4140
rect -1482 4118 -1478 4140
rect -1458 4118 -1454 4140
rect -1434 4118 -1430 4140
rect -1410 4118 -1406 4140
rect -1397 4133 -1392 4140
rect -1386 4133 -1382 4140
rect -1387 4119 -1382 4133
rect -1397 4118 -1363 4119
rect -1362 4118 -1358 4164
rect -1338 4118 -1334 4164
rect -1314 4118 -1310 4164
rect -1290 4118 -1286 4164
rect -1266 4118 -1262 4164
rect -1242 4163 -1238 4164
rect -1242 4118 -1235 4163
rect -1218 4118 -1214 4164
rect -1194 4118 -1190 4164
rect -1170 4118 -1166 4164
rect -1146 4118 -1142 4164
rect -1122 4118 -1118 4164
rect -1098 4118 -1094 4164
rect -1074 4118 -1070 4164
rect -1050 4118 -1046 4164
rect -1026 4118 -1022 4164
rect -1002 4118 -998 4164
rect -978 4118 -974 4164
rect -954 4118 -950 4164
rect -930 4118 -926 4164
rect -906 4118 -902 4164
rect -882 4118 -878 4164
rect -858 4118 -854 4164
rect -834 4139 -830 4164
rect -2393 4116 -837 4118
rect -2371 4070 -2366 4116
rect -2348 4070 -2343 4116
rect -2325 4070 -2320 4116
rect -2317 4112 -2309 4116
rect -2062 4112 -2054 4116
rect -2154 4108 -2138 4110
rect -2057 4108 -2054 4112
rect -2292 4102 -2054 4108
rect -2052 4102 -2044 4112
rect -2092 4086 -2062 4088
rect -2094 4082 -2062 4086
rect -2000 4070 -1992 4116
rect -1846 4109 -1806 4116
rect -1663 4112 -1655 4116
rect -1846 4102 -1680 4108
rect -1854 4086 -1806 4088
rect -1854 4082 -1680 4086
rect -1642 4070 -1637 4116
rect -1619 4070 -1614 4116
rect -1530 4070 -1526 4116
rect -1506 4070 -1502 4116
rect -1482 4070 -1478 4116
rect -1458 4070 -1454 4116
rect -1434 4070 -1430 4116
rect -1410 4070 -1406 4116
rect -1397 4109 -1392 4116
rect -1387 4095 -1382 4109
rect -1386 4070 -1382 4095
rect -1362 4070 -1358 4116
rect -1338 4070 -1334 4116
rect -1314 4070 -1310 4116
rect -1290 4070 -1286 4116
rect -1266 4070 -1262 4116
rect -1259 4115 -1245 4116
rect -1242 4115 -1235 4116
rect -1242 4070 -1238 4115
rect -1218 4070 -1214 4116
rect -1194 4070 -1190 4116
rect -1170 4070 -1166 4116
rect -1146 4070 -1142 4116
rect -1122 4070 -1118 4116
rect -1098 4070 -1094 4116
rect -1074 4070 -1070 4116
rect -1050 4070 -1046 4116
rect -1026 4070 -1022 4116
rect -1002 4070 -998 4116
rect -978 4070 -974 4116
rect -954 4070 -950 4116
rect -930 4070 -926 4116
rect -906 4070 -902 4116
rect -882 4070 -878 4116
rect -858 4070 -854 4116
rect -851 4115 -837 4116
rect -834 4091 -827 4139
rect -834 4070 -830 4091
rect -810 4070 -806 4164
rect -786 4070 -782 4164
rect -762 4070 -758 4164
rect -738 4070 -734 4164
rect -714 4070 -710 4164
rect -690 4070 -686 4164
rect -666 4070 -662 4164
rect -642 4070 -638 4164
rect -618 4070 -614 4164
rect -594 4070 -590 4164
rect -570 4070 -566 4164
rect -546 4070 -542 4164
rect -522 4070 -518 4164
rect -498 4070 -494 4164
rect -474 4070 -470 4164
rect -450 4070 -446 4164
rect -426 4070 -422 4164
rect -402 4070 -398 4164
rect -378 4070 -374 4164
rect -354 4070 -350 4164
rect -330 4070 -326 4164
rect -306 4070 -302 4164
rect -282 4070 -278 4164
rect -258 4070 -254 4164
rect -234 4070 -230 4164
rect -210 4070 -206 4164
rect -186 4070 -182 4164
rect -162 4070 -158 4164
rect -138 4070 -134 4164
rect -114 4070 -110 4164
rect -90 4070 -86 4164
rect -66 4070 -62 4164
rect -42 4070 -38 4164
rect -18 4070 -14 4164
rect 6 4070 10 4164
rect 30 4070 34 4164
rect 54 4070 58 4164
rect 78 4070 82 4164
rect 102 4070 106 4164
rect 126 4070 130 4164
rect 150 4070 154 4164
rect 174 4070 178 4164
rect 198 4070 202 4164
rect 222 4070 226 4164
rect 246 4070 250 4164
rect 270 4070 274 4164
rect 294 4070 298 4164
rect 318 4070 322 4164
rect 342 4070 346 4164
rect 366 4070 370 4164
rect 390 4070 394 4164
rect 414 4070 418 4164
rect 438 4070 442 4164
rect 462 4070 466 4164
rect 486 4070 490 4164
rect 510 4070 514 4164
rect 534 4070 538 4164
rect 558 4070 562 4164
rect 582 4070 586 4164
rect 606 4070 610 4164
rect 613 4163 627 4164
rect 630 4163 637 4187
rect 630 4070 634 4163
rect 654 4070 658 4188
rect 678 4070 682 4188
rect 702 4070 706 4188
rect 726 4070 730 4188
rect 750 4070 754 4188
rect 774 4070 778 4188
rect 798 4070 802 4188
rect 822 4070 826 4188
rect 846 4070 850 4188
rect 870 4070 874 4188
rect 894 4070 898 4188
rect 918 4070 922 4188
rect 942 4070 946 4188
rect 966 4070 970 4188
rect 990 4070 994 4188
rect 1014 4070 1018 4188
rect 1038 4070 1042 4188
rect 1062 4070 1066 4188
rect 1086 4070 1090 4188
rect 1110 4070 1114 4188
rect 1134 4070 1138 4188
rect 1158 4070 1162 4188
rect 1182 4070 1186 4188
rect 1206 4070 1210 4188
rect 1230 4070 1234 4188
rect 1254 4070 1258 4188
rect 1278 4070 1282 4188
rect 1302 4070 1306 4188
rect 1326 4070 1330 4188
rect 1350 4070 1354 4188
rect 1374 4070 1378 4188
rect 1398 4070 1402 4188
rect 1422 4070 1426 4188
rect 1446 4070 1450 4188
rect 1470 4070 1474 4188
rect 1494 4070 1498 4188
rect 1518 4070 1522 4188
rect 1542 4070 1546 4188
rect 1566 4070 1570 4188
rect 1590 4070 1594 4188
rect 1614 4070 1618 4188
rect 1638 4070 1642 4188
rect 1662 4070 1666 4188
rect 1686 4070 1690 4188
rect 1710 4070 1714 4188
rect 1734 4070 1738 4188
rect 1758 4070 1762 4188
rect 1782 4070 1786 4188
rect 1806 4070 1810 4188
rect 1830 4070 1834 4188
rect 1854 4070 1858 4188
rect 1878 4070 1882 4188
rect 1902 4070 1906 4188
rect 1926 4070 1930 4188
rect 1950 4070 1954 4188
rect 1974 4070 1978 4188
rect 1998 4070 2002 4188
rect 2022 4070 2026 4188
rect 2046 4070 2050 4188
rect 2070 4070 2074 4188
rect 2094 4070 2098 4188
rect 2118 4070 2122 4188
rect 2142 4070 2146 4188
rect 2166 4070 2170 4188
rect 2190 4070 2194 4188
rect 2214 4070 2218 4188
rect 2227 4109 2232 4119
rect 2238 4109 2242 4188
rect 2237 4095 2242 4109
rect 2227 4094 2261 4095
rect 2262 4094 2266 4188
rect 2286 4094 2290 4188
rect 2299 4181 2304 4188
rect 2310 4181 2314 4188
rect 2309 4167 2314 4181
rect 2299 4157 2304 4167
rect 2309 4143 2314 4157
rect 2310 4095 2314 4143
rect 2299 4094 2331 4095
rect 2227 4092 2331 4094
rect 2227 4085 2232 4092
rect 2237 4071 2242 4085
rect 2238 4070 2242 4071
rect 2262 4070 2266 4092
rect 2286 4070 2290 4092
rect 2299 4085 2304 4092
rect 2310 4085 2314 4092
rect 2317 4091 2331 4092
rect 2309 4071 2314 4085
rect 2323 4081 2331 4085
rect 2317 4071 2323 4081
rect 2299 4070 2331 4071
rect -2393 4068 2331 4070
rect -2371 4046 -2366 4068
rect -2348 4046 -2343 4068
rect -2325 4046 -2320 4068
rect -2072 4066 -2036 4067
rect -2072 4060 -2054 4066
rect -2309 4052 -2301 4060
rect -2317 4046 -2309 4052
rect -2092 4051 -2062 4056
rect -2000 4047 -1992 4068
rect -1938 4067 -1906 4068
rect -1920 4066 -1906 4067
rect -1806 4060 -1680 4066
rect -1854 4051 -1806 4056
rect -1655 4052 -1647 4060
rect -1982 4047 -1966 4048
rect -2000 4046 -1966 4047
rect -1846 4046 -1806 4049
rect -1663 4046 -1655 4052
rect -1642 4046 -1637 4068
rect -1619 4046 -1614 4068
rect -1530 4046 -1526 4068
rect -1506 4046 -1502 4068
rect -1482 4046 -1478 4068
rect -1458 4046 -1454 4068
rect -1434 4046 -1430 4068
rect -1410 4046 -1406 4068
rect -1386 4047 -1382 4068
rect -1362 4067 -1358 4068
rect -1397 4046 -1365 4047
rect -2393 4044 -1365 4046
rect -2371 4022 -2366 4044
rect -2348 4022 -2343 4044
rect -2325 4022 -2320 4044
rect -2000 4042 -1966 4044
rect -2309 4024 -2301 4032
rect -2062 4031 -2054 4038
rect -2092 4024 -2084 4031
rect -2062 4024 -2026 4026
rect -2317 4022 -2309 4024
rect -2062 4022 -2012 4024
rect -2000 4022 -1992 4042
rect -1982 4041 -1966 4042
rect -1846 4040 -1806 4044
rect -1846 4033 -1798 4038
rect -1806 4031 -1798 4033
rect -1854 4029 -1846 4031
rect -1854 4024 -1806 4029
rect -1655 4024 -1647 4032
rect -1864 4022 -1796 4023
rect -1663 4022 -1655 4024
rect -1642 4022 -1637 4044
rect -1619 4022 -1614 4044
rect -1530 4022 -1526 4044
rect -1506 4022 -1502 4044
rect -1482 4022 -1478 4044
rect -1458 4022 -1454 4044
rect -1434 4022 -1430 4044
rect -1410 4022 -1406 4044
rect -1397 4037 -1392 4044
rect -1386 4037 -1382 4044
rect -1379 4043 -1365 4044
rect -1387 4023 -1382 4037
rect -1373 4033 -1365 4037
rect -1379 4023 -1373 4033
rect -1386 4022 -1382 4023
rect -1362 4022 -1355 4067
rect -1338 4022 -1334 4068
rect -1314 4022 -1310 4068
rect -1290 4022 -1286 4068
rect -1266 4022 -1262 4068
rect -1242 4022 -1238 4068
rect -1218 4022 -1214 4068
rect -1194 4022 -1190 4068
rect -1170 4022 -1166 4068
rect -1146 4022 -1142 4068
rect -1122 4022 -1118 4068
rect -1098 4022 -1094 4068
rect -1074 4022 -1070 4068
rect -1050 4022 -1046 4068
rect -1026 4022 -1022 4068
rect -1002 4022 -998 4068
rect -978 4022 -974 4068
rect -954 4022 -950 4068
rect -930 4022 -926 4068
rect -906 4022 -902 4068
rect -882 4022 -878 4068
rect -858 4022 -854 4068
rect -834 4022 -830 4068
rect -810 4022 -806 4068
rect -786 4022 -782 4068
rect -762 4022 -758 4068
rect -738 4022 -734 4068
rect -714 4022 -710 4068
rect -690 4022 -686 4068
rect -666 4022 -662 4068
rect -642 4022 -638 4068
rect -618 4022 -614 4068
rect -594 4022 -590 4068
rect -570 4022 -566 4068
rect -546 4022 -542 4068
rect -522 4022 -518 4068
rect -498 4022 -494 4068
rect -474 4022 -470 4068
rect -450 4022 -446 4068
rect -426 4022 -422 4068
rect -402 4022 -398 4068
rect -378 4022 -374 4068
rect -354 4022 -350 4068
rect -330 4022 -326 4068
rect -306 4022 -302 4068
rect -282 4022 -278 4068
rect -258 4022 -254 4068
rect -234 4022 -230 4068
rect -210 4022 -206 4068
rect -186 4022 -182 4068
rect -162 4022 -158 4068
rect -138 4022 -134 4068
rect -114 4022 -110 4068
rect -90 4022 -86 4068
rect -66 4022 -62 4068
rect -42 4022 -38 4068
rect -18 4022 -14 4068
rect 6 4022 10 4068
rect 30 4022 34 4068
rect 54 4022 58 4068
rect 78 4022 82 4068
rect 102 4022 106 4068
rect 126 4022 130 4068
rect 150 4022 154 4068
rect 174 4022 178 4068
rect 198 4022 202 4068
rect 222 4022 226 4068
rect 246 4022 250 4068
rect 270 4022 274 4068
rect 294 4022 298 4068
rect 318 4022 322 4068
rect 342 4022 346 4068
rect 366 4022 370 4068
rect 390 4022 394 4068
rect 414 4022 418 4068
rect 438 4022 442 4068
rect 462 4022 466 4068
rect 486 4022 490 4068
rect 510 4022 514 4068
rect 534 4022 538 4068
rect 558 4022 562 4068
rect 582 4022 586 4068
rect 606 4022 610 4068
rect 630 4022 634 4068
rect 654 4022 658 4068
rect 678 4022 682 4068
rect 702 4022 706 4068
rect 726 4022 730 4068
rect 750 4022 754 4068
rect 774 4023 778 4068
rect 763 4022 797 4023
rect -2393 4020 797 4022
rect -2371 3974 -2366 4020
rect -2348 3974 -2343 4020
rect -2325 3974 -2320 4020
rect -2317 4016 -2309 4020
rect -2062 4016 -2054 4020
rect -2154 4012 -2138 4014
rect -2057 4012 -2054 4016
rect -2292 4006 -2054 4012
rect -2052 4006 -2044 4016
rect -2092 3990 -2062 3992
rect -2094 3986 -2062 3990
rect -2000 3974 -1992 4020
rect -1846 4013 -1806 4020
rect -1663 4016 -1655 4020
rect -1846 4006 -1680 4012
rect -1854 3990 -1806 3992
rect -1854 3986 -1680 3990
rect -1642 3974 -1637 4020
rect -1619 3974 -1614 4020
rect -1530 3974 -1526 4020
rect -1506 3974 -1502 4020
rect -1482 3974 -1478 4020
rect -1458 3974 -1454 4020
rect -1434 3974 -1430 4020
rect -1410 3974 -1406 4020
rect -1386 3974 -1382 4020
rect -1379 4019 -1365 4020
rect -1362 4019 -1355 4020
rect -1362 3974 -1358 4019
rect -1338 3974 -1334 4020
rect -1314 3974 -1310 4020
rect -1290 3974 -1286 4020
rect -1266 3974 -1262 4020
rect -1242 3974 -1238 4020
rect -1218 3974 -1214 4020
rect -1194 3974 -1190 4020
rect -1170 3974 -1166 4020
rect -1146 3974 -1142 4020
rect -1122 3974 -1118 4020
rect -1098 3974 -1094 4020
rect -1074 3974 -1070 4020
rect -1050 3974 -1046 4020
rect -1026 3974 -1022 4020
rect -1002 3974 -998 4020
rect -978 3974 -974 4020
rect -954 3974 -950 4020
rect -930 3974 -926 4020
rect -906 3974 -902 4020
rect -882 3974 -878 4020
rect -858 3974 -854 4020
rect -834 3974 -830 4020
rect -810 3974 -806 4020
rect -786 3974 -782 4020
rect -762 3974 -758 4020
rect -738 3974 -734 4020
rect -714 3974 -710 4020
rect -690 3974 -686 4020
rect -666 3974 -662 4020
rect -642 3974 -638 4020
rect -618 3974 -614 4020
rect -594 3974 -590 4020
rect -570 3974 -566 4020
rect -546 3974 -542 4020
rect -522 3974 -518 4020
rect -498 3974 -494 4020
rect -474 3974 -470 4020
rect -450 3974 -446 4020
rect -426 3974 -422 4020
rect -402 3974 -398 4020
rect -378 3974 -374 4020
rect -354 3974 -350 4020
rect -330 3974 -326 4020
rect -306 3974 -302 4020
rect -282 3974 -278 4020
rect -258 3974 -254 4020
rect -234 3974 -230 4020
rect -210 3974 -206 4020
rect -186 3974 -182 4020
rect -162 3974 -158 4020
rect -138 3974 -134 4020
rect -114 3974 -110 4020
rect -90 3974 -86 4020
rect -66 3974 -62 4020
rect -42 3974 -38 4020
rect -18 3974 -14 4020
rect 6 3974 10 4020
rect 30 3974 34 4020
rect 54 3974 58 4020
rect 78 3974 82 4020
rect 102 3974 106 4020
rect 126 3974 130 4020
rect 150 3974 154 4020
rect 174 3974 178 4020
rect 198 3974 202 4020
rect 222 3974 226 4020
rect 246 3974 250 4020
rect 270 3974 274 4020
rect 294 3974 298 4020
rect 318 3974 322 4020
rect 342 3974 346 4020
rect 366 3974 370 4020
rect 390 3974 394 4020
rect 414 3974 418 4020
rect 438 3974 442 4020
rect 462 3974 466 4020
rect 486 3974 490 4020
rect 510 3974 514 4020
rect 534 3974 538 4020
rect 558 3974 562 4020
rect 582 3974 586 4020
rect 606 3974 610 4020
rect 630 3974 634 4020
rect 654 3974 658 4020
rect 678 3974 682 4020
rect 702 3974 706 4020
rect 726 3974 730 4020
rect 750 3974 754 4020
rect 763 4013 768 4020
rect 774 4013 778 4020
rect 773 3999 778 4013
rect 763 3989 768 3999
rect 773 3975 778 3989
rect 774 3974 778 3975
rect 798 3974 802 4068
rect 822 3974 826 4068
rect 846 3974 850 4068
rect 870 3974 874 4068
rect 894 3974 898 4068
rect 918 3974 922 4068
rect 942 3974 946 4068
rect 966 3974 970 4068
rect 990 3974 994 4068
rect 1014 3974 1018 4068
rect 1038 3974 1042 4068
rect 1062 3974 1066 4068
rect 1086 3974 1090 4068
rect 1110 3974 1114 4068
rect 1134 3974 1138 4068
rect 1158 3974 1162 4068
rect 1182 3974 1186 4068
rect 1206 3974 1210 4068
rect 1230 3974 1234 4068
rect 1254 3974 1258 4068
rect 1278 3974 1282 4068
rect 1302 3974 1306 4068
rect 1326 3974 1330 4068
rect 1350 3974 1354 4068
rect 1374 3974 1378 4068
rect 1398 3974 1402 4068
rect 1422 3974 1426 4068
rect 1446 3974 1450 4068
rect 1470 3974 1474 4068
rect 1494 3974 1498 4068
rect 1518 3974 1522 4068
rect 1542 3974 1546 4068
rect 1566 3974 1570 4068
rect 1590 3974 1594 4068
rect 1614 3974 1618 4068
rect 1638 3974 1642 4068
rect 1662 3974 1666 4068
rect 1686 3974 1690 4068
rect 1710 3974 1714 4068
rect 1734 3974 1738 4068
rect 1758 3974 1762 4068
rect 1782 3974 1786 4068
rect 1806 3974 1810 4068
rect 1830 3974 1834 4068
rect 1854 3974 1858 4068
rect 1878 3974 1882 4068
rect 1902 3974 1906 4068
rect 1926 3974 1930 4068
rect 1950 3974 1954 4068
rect 1974 3974 1978 4068
rect 1998 3974 2002 4068
rect 2022 3974 2026 4068
rect 2046 3974 2050 4068
rect 2070 3974 2074 4068
rect 2094 3974 2098 4068
rect 2118 3974 2122 4068
rect 2142 3974 2146 4068
rect 2166 3974 2170 4068
rect 2190 3974 2194 4068
rect 2214 3974 2218 4068
rect 2238 3974 2242 4068
rect 2262 4043 2266 4068
rect 2262 3998 2269 4043
rect 2286 3998 2290 4068
rect 2299 4061 2304 4068
rect 2317 4067 2331 4068
rect 2309 4047 2314 4061
rect 2310 3999 2314 4047
rect 2299 3998 2331 3999
rect 2245 3996 2331 3998
rect 2245 3995 2259 3996
rect 2262 3995 2269 3996
rect 2262 3974 2266 3995
rect 2286 3974 2290 3996
rect 2299 3989 2304 3996
rect 2310 3989 2314 3996
rect 2317 3995 2331 3996
rect 2309 3975 2314 3989
rect 2323 3985 2331 3989
rect 2317 3975 2323 3985
rect 2299 3974 2331 3975
rect -2393 3972 2331 3974
rect -2371 3950 -2366 3972
rect -2348 3950 -2343 3972
rect -2325 3950 -2320 3972
rect -2072 3970 -2036 3971
rect -2072 3964 -2054 3970
rect -2309 3956 -2301 3964
rect -2317 3950 -2309 3956
rect -2092 3955 -2062 3960
rect -2000 3951 -1992 3972
rect -1938 3971 -1906 3972
rect -1920 3970 -1906 3971
rect -1806 3964 -1680 3970
rect -1854 3955 -1806 3960
rect -1655 3956 -1647 3964
rect -1982 3951 -1966 3952
rect -2000 3950 -1966 3951
rect -1846 3950 -1806 3953
rect -1663 3950 -1655 3956
rect -1642 3950 -1637 3972
rect -1619 3950 -1614 3972
rect -1530 3950 -1526 3972
rect -1506 3950 -1502 3972
rect -1482 3950 -1478 3972
rect -1458 3950 -1454 3972
rect -1434 3950 -1430 3972
rect -1410 3950 -1406 3972
rect -1386 3950 -1382 3972
rect -1362 3971 -1358 3972
rect -2393 3948 -1365 3950
rect -2371 3926 -2366 3948
rect -2348 3926 -2343 3948
rect -2325 3926 -2320 3948
rect -2000 3946 -1966 3948
rect -2309 3928 -2301 3936
rect -2062 3935 -2054 3942
rect -2092 3928 -2084 3935
rect -2062 3928 -2026 3930
rect -2317 3926 -2309 3928
rect -2062 3926 -2012 3928
rect -2000 3926 -1992 3946
rect -1982 3945 -1966 3946
rect -1846 3944 -1806 3948
rect -1846 3937 -1798 3942
rect -1806 3935 -1798 3937
rect -1854 3933 -1846 3935
rect -1854 3928 -1806 3933
rect -1655 3928 -1647 3936
rect -1864 3926 -1796 3927
rect -1663 3926 -1655 3928
rect -1642 3926 -1637 3948
rect -1619 3926 -1614 3948
rect -1530 3926 -1526 3948
rect -1506 3926 -1502 3948
rect -1482 3926 -1478 3948
rect -1458 3926 -1454 3948
rect -1434 3926 -1430 3948
rect -1410 3926 -1406 3948
rect -1386 3926 -1382 3948
rect -1379 3947 -1365 3948
rect -1362 3947 -1355 3971
rect -1362 3926 -1358 3947
rect -1338 3927 -1334 3972
rect -1349 3926 -1315 3927
rect -2393 3924 -1315 3926
rect -2371 3878 -2366 3924
rect -2348 3878 -2343 3924
rect -2325 3878 -2320 3924
rect -2317 3920 -2309 3924
rect -2062 3920 -2054 3924
rect -2154 3916 -2138 3918
rect -2057 3916 -2054 3920
rect -2292 3910 -2054 3916
rect -2052 3910 -2044 3920
rect -2092 3894 -2062 3896
rect -2094 3890 -2062 3894
rect -2000 3878 -1992 3924
rect -1846 3917 -1806 3924
rect -1663 3920 -1655 3924
rect -1846 3910 -1680 3916
rect -1854 3894 -1806 3896
rect -1854 3890 -1680 3894
rect -1642 3878 -1637 3924
rect -1619 3878 -1614 3924
rect -1530 3878 -1526 3924
rect -1506 3878 -1502 3924
rect -1482 3878 -1478 3924
rect -1458 3878 -1454 3924
rect -1434 3878 -1430 3924
rect -1410 3878 -1406 3924
rect -1386 3878 -1382 3924
rect -1362 3878 -1358 3924
rect -1349 3917 -1344 3924
rect -1338 3917 -1334 3924
rect -1339 3903 -1334 3917
rect -1349 3893 -1344 3903
rect -1339 3879 -1334 3893
rect -1338 3878 -1334 3879
rect -1314 3878 -1310 3972
rect -1290 3878 -1286 3972
rect -1266 3878 -1262 3972
rect -1242 3878 -1238 3972
rect -1218 3878 -1214 3972
rect -1194 3878 -1190 3972
rect -1170 3878 -1166 3972
rect -1146 3878 -1142 3972
rect -1122 3878 -1118 3972
rect -1098 3878 -1094 3972
rect -1074 3878 -1070 3972
rect -1050 3878 -1046 3972
rect -1026 3878 -1022 3972
rect -1002 3878 -998 3972
rect -978 3878 -974 3972
rect -954 3878 -950 3972
rect -930 3878 -926 3972
rect -906 3878 -902 3972
rect -882 3878 -878 3972
rect -858 3878 -854 3972
rect -834 3878 -830 3972
rect -810 3878 -806 3972
rect -786 3878 -782 3972
rect -762 3878 -758 3972
rect -738 3878 -734 3972
rect -714 3878 -710 3972
rect -690 3878 -686 3972
rect -666 3878 -662 3972
rect -642 3878 -638 3972
rect -618 3878 -614 3972
rect -594 3878 -590 3972
rect -570 3878 -566 3972
rect -546 3878 -542 3972
rect -522 3878 -518 3972
rect -498 3878 -494 3972
rect -474 3878 -470 3972
rect -450 3878 -446 3972
rect -426 3878 -422 3972
rect -402 3878 -398 3972
rect -378 3878 -374 3972
rect -354 3878 -350 3972
rect -330 3878 -326 3972
rect -306 3878 -302 3972
rect -282 3878 -278 3972
rect -258 3878 -254 3972
rect -234 3878 -230 3972
rect -210 3878 -206 3972
rect -186 3878 -182 3972
rect -162 3878 -158 3972
rect -138 3878 -134 3972
rect -114 3878 -110 3972
rect -90 3878 -86 3972
rect -66 3878 -62 3972
rect -42 3878 -38 3972
rect -18 3878 -14 3972
rect 6 3878 10 3972
rect 30 3878 34 3972
rect 54 3878 58 3972
rect 78 3878 82 3972
rect 102 3878 106 3972
rect 126 3878 130 3972
rect 150 3878 154 3972
rect 174 3878 178 3972
rect 198 3878 202 3972
rect 222 3878 226 3972
rect 246 3878 250 3972
rect 270 3878 274 3972
rect 294 3878 298 3972
rect 318 3878 322 3972
rect 342 3878 346 3972
rect 366 3878 370 3972
rect 390 3878 394 3972
rect 414 3878 418 3972
rect 438 3878 442 3972
rect 462 3878 466 3972
rect 486 3878 490 3972
rect 510 3878 514 3972
rect 523 3941 528 3951
rect 534 3941 538 3972
rect 533 3927 538 3941
rect 523 3926 557 3927
rect 558 3926 562 3972
rect 582 3926 586 3972
rect 606 3926 610 3972
rect 630 3926 634 3972
rect 654 3926 658 3972
rect 678 3926 682 3972
rect 702 3926 706 3972
rect 726 3926 730 3972
rect 750 3926 754 3972
rect 774 3926 778 3972
rect 798 3947 802 3972
rect 523 3924 795 3926
rect 523 3917 528 3924
rect 533 3903 538 3917
rect 534 3878 538 3903
rect 558 3878 562 3924
rect 582 3878 586 3924
rect 606 3878 610 3924
rect 630 3878 634 3924
rect 654 3878 658 3924
rect 678 3878 682 3924
rect 702 3878 706 3924
rect 726 3878 730 3924
rect 750 3878 754 3924
rect 774 3878 778 3924
rect 781 3923 795 3924
rect 798 3902 805 3947
rect 822 3902 826 3972
rect 846 3902 850 3972
rect 870 3902 874 3972
rect 894 3902 898 3972
rect 918 3902 922 3972
rect 942 3902 946 3972
rect 966 3902 970 3972
rect 990 3902 994 3972
rect 1014 3902 1018 3972
rect 1038 3902 1042 3972
rect 1062 3902 1066 3972
rect 1086 3902 1090 3972
rect 1110 3902 1114 3972
rect 1134 3902 1138 3972
rect 1158 3902 1162 3972
rect 1182 3902 1186 3972
rect 1206 3902 1210 3972
rect 1230 3902 1234 3972
rect 1254 3902 1258 3972
rect 1278 3902 1282 3972
rect 1302 3902 1306 3972
rect 1326 3902 1330 3972
rect 1350 3902 1354 3972
rect 1374 3902 1378 3972
rect 1398 3902 1402 3972
rect 1422 3902 1426 3972
rect 1446 3902 1450 3972
rect 1470 3902 1474 3972
rect 1494 3902 1498 3972
rect 1518 3902 1522 3972
rect 1542 3902 1546 3972
rect 1566 3902 1570 3972
rect 1590 3902 1594 3972
rect 1614 3902 1618 3972
rect 1638 3902 1642 3972
rect 1662 3902 1666 3972
rect 1686 3902 1690 3972
rect 1710 3902 1714 3972
rect 1734 3902 1738 3972
rect 1758 3902 1762 3972
rect 1782 3902 1786 3972
rect 1806 3902 1810 3972
rect 1830 3902 1834 3972
rect 1854 3902 1858 3972
rect 1878 3902 1882 3972
rect 1902 3902 1906 3972
rect 1926 3902 1930 3972
rect 1950 3902 1954 3972
rect 1974 3902 1978 3972
rect 1998 3902 2002 3972
rect 2022 3902 2026 3972
rect 2046 3902 2050 3972
rect 2070 3902 2074 3972
rect 2094 3902 2098 3972
rect 2118 3902 2122 3972
rect 2142 3902 2146 3972
rect 2166 3902 2170 3972
rect 2190 3902 2194 3972
rect 2214 3902 2218 3972
rect 2238 3902 2242 3972
rect 2262 3902 2266 3972
rect 2286 3903 2290 3972
rect 2299 3965 2304 3972
rect 2317 3971 2331 3972
rect 2309 3951 2314 3965
rect 2299 3917 2304 3927
rect 2310 3917 2314 3951
rect 2309 3903 2314 3917
rect 2323 3913 2331 3917
rect 2317 3903 2323 3913
rect 2275 3902 2309 3903
rect 781 3900 2309 3902
rect 781 3899 795 3900
rect 798 3899 805 3900
rect 798 3878 802 3899
rect 822 3878 826 3900
rect 846 3878 850 3900
rect 870 3878 874 3900
rect 894 3878 898 3900
rect 918 3878 922 3900
rect 942 3878 946 3900
rect 966 3878 970 3900
rect 990 3878 994 3900
rect 1014 3878 1018 3900
rect 1038 3878 1042 3900
rect 1062 3878 1066 3900
rect 1086 3878 1090 3900
rect 1110 3878 1114 3900
rect 1134 3878 1138 3900
rect 1158 3878 1162 3900
rect 1182 3878 1186 3900
rect 1206 3878 1210 3900
rect 1230 3878 1234 3900
rect 1254 3878 1258 3900
rect 1278 3878 1282 3900
rect 1302 3878 1306 3900
rect 1326 3878 1330 3900
rect 1350 3878 1354 3900
rect 1374 3878 1378 3900
rect 1398 3878 1402 3900
rect 1422 3878 1426 3900
rect 1446 3878 1450 3900
rect 1470 3878 1474 3900
rect 1494 3878 1498 3900
rect 1518 3878 1522 3900
rect 1542 3878 1546 3900
rect 1566 3878 1570 3900
rect 1590 3878 1594 3900
rect 1614 3878 1618 3900
rect 1638 3878 1642 3900
rect 1662 3878 1666 3900
rect 1686 3878 1690 3900
rect 1710 3878 1714 3900
rect 1734 3878 1738 3900
rect 1758 3878 1762 3900
rect 1782 3878 1786 3900
rect 1806 3878 1810 3900
rect 1830 3878 1834 3900
rect 1854 3878 1858 3900
rect 1878 3878 1882 3900
rect 1902 3878 1906 3900
rect 1926 3878 1930 3900
rect 1950 3878 1954 3900
rect 1974 3878 1978 3900
rect 1998 3878 2002 3900
rect 2022 3878 2026 3900
rect 2046 3878 2050 3900
rect 2070 3878 2074 3900
rect 2094 3878 2098 3900
rect 2118 3878 2122 3900
rect 2142 3878 2146 3900
rect 2166 3878 2170 3900
rect 2190 3878 2194 3900
rect 2214 3878 2218 3900
rect 2238 3878 2242 3900
rect 2262 3878 2266 3900
rect 2275 3893 2280 3900
rect 2286 3893 2290 3900
rect 2285 3879 2290 3893
rect 2275 3878 2309 3879
rect -2393 3876 2309 3878
rect -2371 3854 -2366 3876
rect -2348 3854 -2343 3876
rect -2325 3854 -2320 3876
rect -2072 3874 -2036 3875
rect -2072 3868 -2054 3874
rect -2309 3860 -2301 3868
rect -2317 3854 -2309 3860
rect -2092 3859 -2062 3864
rect -2000 3855 -1992 3876
rect -1938 3875 -1906 3876
rect -1920 3874 -1906 3875
rect -1806 3868 -1680 3874
rect -1854 3859 -1806 3864
rect -1655 3860 -1647 3868
rect -1982 3855 -1966 3856
rect -2000 3854 -1966 3855
rect -1846 3854 -1806 3857
rect -1663 3854 -1655 3860
rect -1642 3854 -1637 3876
rect -1619 3854 -1614 3876
rect -1530 3854 -1526 3876
rect -1506 3854 -1502 3876
rect -1482 3854 -1478 3876
rect -1458 3854 -1454 3876
rect -1434 3854 -1430 3876
rect -1410 3854 -1406 3876
rect -1386 3854 -1382 3876
rect -1362 3854 -1358 3876
rect -1338 3854 -1334 3876
rect -1314 3854 -1310 3876
rect -1290 3854 -1286 3876
rect -1266 3854 -1262 3876
rect -1242 3854 -1238 3876
rect -1218 3854 -1214 3876
rect -1194 3854 -1190 3876
rect -1170 3854 -1166 3876
rect -1146 3854 -1142 3876
rect -1122 3854 -1118 3876
rect -1098 3854 -1094 3876
rect -1074 3854 -1070 3876
rect -1050 3854 -1046 3876
rect -1026 3854 -1022 3876
rect -1002 3854 -998 3876
rect -978 3854 -974 3876
rect -954 3854 -950 3876
rect -930 3854 -926 3876
rect -906 3854 -902 3876
rect -882 3854 -878 3876
rect -858 3854 -854 3876
rect -834 3854 -830 3876
rect -810 3854 -806 3876
rect -786 3854 -782 3876
rect -762 3854 -758 3876
rect -738 3854 -734 3876
rect -714 3854 -710 3876
rect -690 3854 -686 3876
rect -666 3854 -662 3876
rect -642 3854 -638 3876
rect -618 3854 -614 3876
rect -594 3854 -590 3876
rect -570 3854 -566 3876
rect -546 3854 -542 3876
rect -522 3854 -518 3876
rect -498 3854 -494 3876
rect -474 3854 -470 3876
rect -450 3854 -446 3876
rect -426 3854 -422 3876
rect -402 3854 -398 3876
rect -378 3854 -374 3876
rect -354 3854 -350 3876
rect -330 3854 -326 3876
rect -306 3854 -302 3876
rect -282 3854 -278 3876
rect -258 3854 -254 3876
rect -234 3854 -230 3876
rect -210 3854 -206 3876
rect -186 3854 -182 3876
rect -162 3854 -158 3876
rect -138 3854 -134 3876
rect -114 3854 -110 3876
rect -90 3854 -86 3876
rect -66 3854 -62 3876
rect -42 3854 -38 3876
rect -18 3855 -14 3876
rect -29 3854 5 3855
rect -2393 3852 5 3854
rect -2371 3830 -2366 3852
rect -2348 3830 -2343 3852
rect -2325 3830 -2320 3852
rect -2000 3850 -1966 3852
rect -2309 3832 -2301 3840
rect -2062 3839 -2054 3846
rect -2092 3832 -2084 3839
rect -2062 3832 -2026 3834
rect -2317 3830 -2309 3832
rect -2062 3830 -2012 3832
rect -2000 3830 -1992 3850
rect -1982 3849 -1966 3850
rect -1846 3848 -1806 3852
rect -1846 3841 -1798 3846
rect -1806 3839 -1798 3841
rect -1854 3837 -1846 3839
rect -1854 3832 -1806 3837
rect -1655 3832 -1647 3840
rect -1864 3830 -1796 3831
rect -1663 3830 -1655 3832
rect -1642 3830 -1637 3852
rect -1619 3830 -1614 3852
rect -1530 3830 -1526 3852
rect -1506 3830 -1502 3852
rect -1482 3831 -1478 3852
rect -1493 3830 -1459 3831
rect -2393 3828 -1459 3830
rect -2371 3782 -2366 3828
rect -2348 3782 -2343 3828
rect -2325 3782 -2320 3828
rect -2317 3824 -2309 3828
rect -2062 3824 -2054 3828
rect -2154 3820 -2138 3822
rect -2057 3820 -2054 3824
rect -2292 3814 -2054 3820
rect -2052 3814 -2044 3824
rect -2092 3798 -2062 3800
rect -2094 3794 -2062 3798
rect -2000 3782 -1992 3828
rect -1846 3821 -1806 3828
rect -1663 3824 -1655 3828
rect -1846 3814 -1680 3820
rect -1854 3798 -1806 3800
rect -1854 3794 -1680 3798
rect -1642 3782 -1637 3828
rect -1619 3782 -1614 3828
rect -1530 3782 -1526 3828
rect -1506 3782 -1502 3828
rect -1493 3821 -1488 3828
rect -1482 3821 -1478 3828
rect -1483 3807 -1478 3821
rect -1493 3797 -1488 3807
rect -1483 3783 -1478 3797
rect -1482 3782 -1478 3783
rect -1458 3782 -1454 3852
rect -1434 3782 -1430 3852
rect -1410 3782 -1406 3852
rect -1386 3782 -1382 3852
rect -1362 3782 -1358 3852
rect -1338 3782 -1334 3852
rect -1314 3851 -1310 3852
rect -1314 3806 -1307 3851
rect -1290 3806 -1286 3852
rect -1266 3806 -1262 3852
rect -1242 3806 -1238 3852
rect -1218 3806 -1214 3852
rect -1194 3806 -1190 3852
rect -1170 3806 -1166 3852
rect -1146 3806 -1142 3852
rect -1122 3806 -1118 3852
rect -1098 3806 -1094 3852
rect -1074 3806 -1070 3852
rect -1050 3806 -1046 3852
rect -1026 3806 -1022 3852
rect -1002 3806 -998 3852
rect -978 3806 -974 3852
rect -954 3806 -950 3852
rect -930 3806 -926 3852
rect -906 3806 -902 3852
rect -882 3806 -878 3852
rect -858 3806 -854 3852
rect -834 3806 -830 3852
rect -810 3806 -806 3852
rect -786 3806 -782 3852
rect -762 3806 -758 3852
rect -738 3806 -734 3852
rect -714 3806 -710 3852
rect -690 3806 -686 3852
rect -666 3806 -662 3852
rect -642 3806 -638 3852
rect -618 3806 -614 3852
rect -594 3806 -590 3852
rect -570 3806 -566 3852
rect -546 3806 -542 3852
rect -522 3806 -518 3852
rect -498 3806 -494 3852
rect -474 3806 -470 3852
rect -450 3806 -446 3852
rect -426 3806 -422 3852
rect -402 3806 -398 3852
rect -378 3806 -374 3852
rect -354 3806 -350 3852
rect -330 3806 -326 3852
rect -306 3806 -302 3852
rect -282 3806 -278 3852
rect -258 3806 -254 3852
rect -234 3806 -230 3852
rect -210 3806 -206 3852
rect -186 3806 -182 3852
rect -162 3806 -158 3852
rect -138 3806 -134 3852
rect -114 3806 -110 3852
rect -90 3806 -86 3852
rect -66 3806 -62 3852
rect -42 3806 -38 3852
rect -29 3845 -24 3852
rect -18 3845 -14 3852
rect -19 3831 -14 3845
rect -29 3821 -24 3831
rect -19 3807 -14 3821
rect -18 3806 -14 3807
rect 6 3806 10 3876
rect 30 3806 34 3876
rect 54 3806 58 3876
rect 78 3806 82 3876
rect 102 3806 106 3876
rect 126 3806 130 3876
rect 150 3806 154 3876
rect 174 3806 178 3876
rect 198 3806 202 3876
rect 222 3806 226 3876
rect 246 3806 250 3876
rect 270 3806 274 3876
rect 294 3806 298 3876
rect 318 3806 322 3876
rect 342 3806 346 3876
rect 366 3806 370 3876
rect 390 3806 394 3876
rect 414 3806 418 3876
rect 438 3806 442 3876
rect 462 3806 466 3876
rect 486 3806 490 3876
rect 510 3806 514 3876
rect 534 3806 538 3876
rect 558 3875 562 3876
rect 558 3830 565 3875
rect 582 3830 586 3876
rect 606 3830 610 3876
rect 630 3830 634 3876
rect 654 3830 658 3876
rect 678 3830 682 3876
rect 702 3830 706 3876
rect 726 3830 730 3876
rect 750 3830 754 3876
rect 774 3830 778 3876
rect 798 3830 802 3876
rect 822 3830 826 3876
rect 846 3830 850 3876
rect 870 3830 874 3876
rect 894 3830 898 3876
rect 918 3830 922 3876
rect 942 3830 946 3876
rect 966 3830 970 3876
rect 990 3830 994 3876
rect 1014 3830 1018 3876
rect 1038 3830 1042 3876
rect 1062 3830 1066 3876
rect 1086 3830 1090 3876
rect 1110 3830 1114 3876
rect 1134 3830 1138 3876
rect 1158 3830 1162 3876
rect 1182 3830 1186 3876
rect 1206 3830 1210 3876
rect 1230 3830 1234 3876
rect 1254 3830 1258 3876
rect 1278 3830 1282 3876
rect 1302 3830 1306 3876
rect 1326 3830 1330 3876
rect 1350 3830 1354 3876
rect 1374 3830 1378 3876
rect 1398 3830 1402 3876
rect 1422 3830 1426 3876
rect 1446 3830 1450 3876
rect 1470 3830 1474 3876
rect 1494 3830 1498 3876
rect 1518 3830 1522 3876
rect 1542 3830 1546 3876
rect 1566 3830 1570 3876
rect 1590 3830 1594 3876
rect 1614 3830 1618 3876
rect 1638 3830 1642 3876
rect 1662 3830 1666 3876
rect 1686 3830 1690 3876
rect 1710 3830 1714 3876
rect 1734 3830 1738 3876
rect 1758 3830 1762 3876
rect 1782 3830 1786 3876
rect 1806 3830 1810 3876
rect 1830 3830 1834 3876
rect 1854 3830 1858 3876
rect 1878 3830 1882 3876
rect 1902 3830 1906 3876
rect 1926 3830 1930 3876
rect 1950 3830 1954 3876
rect 1974 3830 1978 3876
rect 1998 3830 2002 3876
rect 2022 3830 2026 3876
rect 2046 3830 2050 3876
rect 2070 3830 2074 3876
rect 2094 3830 2098 3876
rect 2118 3830 2122 3876
rect 2142 3830 2146 3876
rect 2166 3830 2170 3876
rect 2190 3830 2194 3876
rect 2214 3830 2218 3876
rect 2238 3830 2242 3876
rect 2262 3830 2266 3876
rect 2275 3869 2280 3876
rect 2285 3855 2290 3869
rect 2286 3831 2290 3855
rect 2275 3830 2309 3831
rect 541 3828 2309 3830
rect 541 3827 555 3828
rect 558 3827 565 3828
rect 558 3806 562 3827
rect 582 3806 586 3828
rect 606 3806 610 3828
rect 630 3806 634 3828
rect 654 3806 658 3828
rect 678 3806 682 3828
rect 702 3806 706 3828
rect 726 3806 730 3828
rect 750 3806 754 3828
rect 774 3806 778 3828
rect 798 3806 802 3828
rect 822 3806 826 3828
rect 846 3806 850 3828
rect 870 3806 874 3828
rect 894 3806 898 3828
rect 918 3806 922 3828
rect 942 3806 946 3828
rect 966 3806 970 3828
rect 990 3806 994 3828
rect 1014 3806 1018 3828
rect 1038 3806 1042 3828
rect 1062 3806 1066 3828
rect 1086 3806 1090 3828
rect 1110 3806 1114 3828
rect 1134 3806 1138 3828
rect 1158 3806 1162 3828
rect 1182 3806 1186 3828
rect 1206 3806 1210 3828
rect 1230 3806 1234 3828
rect 1254 3806 1258 3828
rect 1278 3806 1282 3828
rect 1302 3806 1306 3828
rect 1326 3806 1330 3828
rect 1350 3806 1354 3828
rect 1374 3806 1378 3828
rect 1398 3806 1402 3828
rect 1422 3806 1426 3828
rect 1446 3806 1450 3828
rect 1470 3806 1474 3828
rect 1494 3806 1498 3828
rect 1518 3806 1522 3828
rect 1542 3806 1546 3828
rect 1566 3806 1570 3828
rect 1590 3806 1594 3828
rect 1614 3806 1618 3828
rect 1638 3806 1642 3828
rect 1662 3806 1666 3828
rect 1686 3806 1690 3828
rect 1710 3806 1714 3828
rect 1734 3806 1738 3828
rect 1758 3806 1762 3828
rect 1782 3806 1786 3828
rect 1806 3806 1810 3828
rect 1830 3806 1834 3828
rect 1854 3806 1858 3828
rect 1878 3806 1882 3828
rect 1902 3806 1906 3828
rect 1926 3806 1930 3828
rect 1950 3806 1954 3828
rect 1974 3806 1978 3828
rect 1998 3806 2002 3828
rect 2022 3806 2026 3828
rect 2046 3806 2050 3828
rect 2070 3806 2074 3828
rect 2094 3806 2098 3828
rect 2118 3806 2122 3828
rect 2142 3806 2146 3828
rect 2166 3806 2170 3828
rect 2190 3806 2194 3828
rect 2214 3806 2218 3828
rect 2238 3806 2242 3828
rect 2262 3807 2266 3828
rect 2275 3821 2280 3828
rect 2286 3821 2290 3828
rect 2285 3807 2290 3821
rect 2299 3817 2307 3821
rect 2293 3807 2299 3817
rect 2251 3806 2285 3807
rect -1331 3804 2285 3806
rect -1331 3803 -1317 3804
rect -1314 3803 -1307 3804
rect -1314 3782 -1310 3803
rect -1290 3782 -1286 3804
rect -1266 3782 -1262 3804
rect -1242 3782 -1238 3804
rect -1218 3782 -1214 3804
rect -1194 3782 -1190 3804
rect -1170 3782 -1166 3804
rect -1146 3782 -1142 3804
rect -1122 3782 -1118 3804
rect -1098 3782 -1094 3804
rect -1074 3782 -1070 3804
rect -1050 3782 -1046 3804
rect -1026 3782 -1022 3804
rect -1002 3782 -998 3804
rect -978 3782 -974 3804
rect -954 3782 -950 3804
rect -930 3782 -926 3804
rect -906 3782 -902 3804
rect -882 3782 -878 3804
rect -858 3782 -854 3804
rect -834 3782 -830 3804
rect -810 3782 -806 3804
rect -786 3782 -782 3804
rect -762 3782 -758 3804
rect -738 3782 -734 3804
rect -714 3782 -710 3804
rect -690 3782 -686 3804
rect -666 3782 -662 3804
rect -642 3782 -638 3804
rect -618 3782 -614 3804
rect -594 3782 -590 3804
rect -570 3782 -566 3804
rect -546 3782 -542 3804
rect -522 3782 -518 3804
rect -498 3782 -494 3804
rect -474 3782 -470 3804
rect -450 3782 -446 3804
rect -426 3782 -422 3804
rect -402 3782 -398 3804
rect -378 3782 -374 3804
rect -354 3782 -350 3804
rect -330 3782 -326 3804
rect -306 3782 -302 3804
rect -282 3782 -278 3804
rect -258 3782 -254 3804
rect -234 3782 -230 3804
rect -210 3782 -206 3804
rect -186 3782 -182 3804
rect -162 3782 -158 3804
rect -138 3782 -134 3804
rect -114 3782 -110 3804
rect -90 3782 -86 3804
rect -66 3782 -62 3804
rect -42 3782 -38 3804
rect -18 3782 -14 3804
rect 6 3782 10 3804
rect 30 3782 34 3804
rect 54 3782 58 3804
rect 78 3782 82 3804
rect 102 3782 106 3804
rect 126 3782 130 3804
rect 150 3782 154 3804
rect 174 3782 178 3804
rect 198 3782 202 3804
rect 222 3782 226 3804
rect 246 3782 250 3804
rect 270 3782 274 3804
rect 294 3782 298 3804
rect 318 3782 322 3804
rect 342 3782 346 3804
rect 366 3782 370 3804
rect 390 3782 394 3804
rect 414 3782 418 3804
rect 438 3782 442 3804
rect 462 3782 466 3804
rect 486 3782 490 3804
rect 510 3782 514 3804
rect 534 3782 538 3804
rect 558 3782 562 3804
rect 582 3782 586 3804
rect 606 3782 610 3804
rect 630 3782 634 3804
rect 654 3782 658 3804
rect 678 3782 682 3804
rect 702 3782 706 3804
rect 726 3782 730 3804
rect 750 3782 754 3804
rect 774 3782 778 3804
rect 798 3782 802 3804
rect 822 3782 826 3804
rect 846 3782 850 3804
rect 870 3782 874 3804
rect 894 3782 898 3804
rect 918 3782 922 3804
rect 942 3782 946 3804
rect 966 3782 970 3804
rect 990 3782 994 3804
rect 1014 3782 1018 3804
rect 1038 3782 1042 3804
rect 1062 3782 1066 3804
rect 1086 3782 1090 3804
rect 1110 3782 1114 3804
rect 1134 3782 1138 3804
rect 1158 3782 1162 3804
rect 1182 3782 1186 3804
rect 1206 3782 1210 3804
rect 1230 3782 1234 3804
rect 1254 3782 1258 3804
rect 1278 3782 1282 3804
rect 1302 3782 1306 3804
rect 1326 3782 1330 3804
rect 1350 3782 1354 3804
rect 1374 3782 1378 3804
rect 1398 3782 1402 3804
rect 1422 3782 1426 3804
rect 1446 3782 1450 3804
rect 1470 3782 1474 3804
rect 1494 3782 1498 3804
rect 1518 3782 1522 3804
rect 1542 3782 1546 3804
rect 1566 3782 1570 3804
rect 1590 3782 1594 3804
rect 1614 3782 1618 3804
rect 1638 3782 1642 3804
rect 1662 3782 1666 3804
rect 1686 3782 1690 3804
rect 1710 3782 1714 3804
rect 1734 3782 1738 3804
rect 1758 3782 1762 3804
rect 1782 3782 1786 3804
rect 1806 3782 1810 3804
rect 1830 3782 1834 3804
rect 1854 3782 1858 3804
rect 1878 3782 1882 3804
rect 1902 3782 1906 3804
rect 1926 3782 1930 3804
rect 1950 3782 1954 3804
rect 1974 3782 1978 3804
rect 1998 3782 2002 3804
rect 2022 3782 2026 3804
rect 2046 3782 2050 3804
rect 2070 3782 2074 3804
rect 2094 3782 2098 3804
rect 2118 3782 2122 3804
rect 2142 3782 2146 3804
rect 2166 3782 2170 3804
rect 2190 3782 2194 3804
rect 2214 3782 2218 3804
rect 2238 3782 2242 3804
rect 2251 3797 2256 3804
rect 2262 3797 2266 3804
rect 2261 3783 2266 3797
rect 2251 3782 2285 3783
rect -2393 3780 2285 3782
rect -2371 3758 -2366 3780
rect -2348 3758 -2343 3780
rect -2325 3758 -2320 3780
rect -2072 3778 -2036 3779
rect -2072 3772 -2054 3778
rect -2309 3764 -2301 3772
rect -2317 3758 -2309 3764
rect -2092 3763 -2062 3768
rect -2000 3759 -1992 3780
rect -1938 3779 -1906 3780
rect -1920 3778 -1906 3779
rect -1806 3772 -1680 3778
rect -1854 3763 -1806 3768
rect -1655 3764 -1647 3772
rect -1982 3759 -1966 3760
rect -2000 3758 -1966 3759
rect -1846 3758 -1806 3761
rect -1663 3758 -1655 3764
rect -1642 3758 -1637 3780
rect -1619 3758 -1614 3780
rect -1530 3758 -1526 3780
rect -1506 3758 -1502 3780
rect -1482 3758 -1478 3780
rect -1458 3758 -1454 3780
rect -1434 3758 -1430 3780
rect -1410 3758 -1406 3780
rect -1386 3758 -1382 3780
rect -1362 3758 -1358 3780
rect -1338 3758 -1334 3780
rect -1314 3758 -1310 3780
rect -1290 3758 -1286 3780
rect -1266 3758 -1262 3780
rect -1242 3758 -1238 3780
rect -1218 3758 -1214 3780
rect -1194 3758 -1190 3780
rect -1170 3758 -1166 3780
rect -1146 3758 -1142 3780
rect -1122 3758 -1118 3780
rect -1098 3758 -1094 3780
rect -1074 3758 -1070 3780
rect -1050 3758 -1046 3780
rect -1026 3758 -1022 3780
rect -1002 3758 -998 3780
rect -978 3758 -974 3780
rect -954 3758 -950 3780
rect -930 3758 -926 3780
rect -906 3758 -902 3780
rect -882 3758 -878 3780
rect -858 3758 -854 3780
rect -834 3758 -830 3780
rect -810 3758 -806 3780
rect -786 3758 -782 3780
rect -762 3758 -758 3780
rect -738 3758 -734 3780
rect -714 3758 -710 3780
rect -690 3758 -686 3780
rect -666 3758 -662 3780
rect -642 3758 -638 3780
rect -618 3758 -614 3780
rect -594 3758 -590 3780
rect -570 3758 -566 3780
rect -546 3759 -542 3780
rect -557 3758 -523 3759
rect -2393 3756 -523 3758
rect -2371 3734 -2366 3756
rect -2348 3734 -2343 3756
rect -2325 3734 -2320 3756
rect -2000 3754 -1966 3756
rect -2309 3736 -2301 3744
rect -2062 3743 -2054 3750
rect -2092 3736 -2084 3743
rect -2062 3736 -2026 3738
rect -2317 3734 -2309 3736
rect -2062 3734 -2012 3736
rect -2000 3734 -1992 3754
rect -1982 3753 -1966 3754
rect -1846 3752 -1806 3756
rect -1846 3745 -1798 3750
rect -1806 3743 -1798 3745
rect -1854 3741 -1846 3743
rect -1854 3736 -1806 3741
rect -1655 3736 -1647 3744
rect -1864 3734 -1796 3735
rect -1663 3734 -1655 3736
rect -1642 3734 -1637 3756
rect -1619 3734 -1614 3756
rect -1530 3734 -1526 3756
rect -1506 3734 -1502 3756
rect -1482 3734 -1478 3756
rect -1458 3755 -1454 3756
rect -2393 3732 -1461 3734
rect -2371 3686 -2366 3732
rect -2348 3686 -2343 3732
rect -2325 3686 -2320 3732
rect -2317 3728 -2309 3732
rect -2062 3728 -2054 3732
rect -2154 3724 -2138 3726
rect -2057 3724 -2054 3728
rect -2292 3718 -2054 3724
rect -2052 3718 -2044 3728
rect -2092 3702 -2062 3704
rect -2094 3698 -2062 3702
rect -2000 3686 -1992 3732
rect -1846 3725 -1806 3732
rect -1663 3728 -1655 3732
rect -1846 3718 -1680 3724
rect -1854 3702 -1806 3704
rect -1854 3698 -1680 3702
rect -1642 3686 -1637 3732
rect -1619 3686 -1614 3732
rect -1530 3686 -1526 3732
rect -1506 3686 -1502 3732
rect -1482 3686 -1478 3732
rect -1475 3731 -1461 3732
rect -1458 3707 -1451 3755
rect -1458 3686 -1454 3707
rect -1434 3686 -1430 3756
rect -1410 3686 -1406 3756
rect -1386 3686 -1382 3756
rect -1362 3686 -1358 3756
rect -1338 3686 -1334 3756
rect -1314 3686 -1310 3756
rect -1290 3686 -1286 3756
rect -1266 3686 -1262 3756
rect -1242 3686 -1238 3756
rect -1218 3686 -1214 3756
rect -1194 3686 -1190 3756
rect -1170 3686 -1166 3756
rect -1146 3686 -1142 3756
rect -1122 3686 -1118 3756
rect -1098 3686 -1094 3756
rect -1074 3686 -1070 3756
rect -1050 3686 -1046 3756
rect -1026 3686 -1022 3756
rect -1002 3686 -998 3756
rect -978 3686 -974 3756
rect -954 3686 -950 3756
rect -930 3686 -926 3756
rect -906 3686 -902 3756
rect -893 3725 -888 3735
rect -882 3725 -878 3756
rect -883 3711 -878 3725
rect -893 3710 -859 3711
rect -858 3710 -854 3756
rect -834 3710 -830 3756
rect -810 3710 -806 3756
rect -786 3710 -782 3756
rect -762 3710 -758 3756
rect -738 3710 -734 3756
rect -714 3710 -710 3756
rect -690 3710 -686 3756
rect -666 3710 -662 3756
rect -642 3710 -638 3756
rect -618 3710 -614 3756
rect -594 3710 -590 3756
rect -570 3710 -566 3756
rect -557 3749 -552 3756
rect -546 3749 -542 3756
rect -547 3735 -542 3749
rect -557 3725 -552 3735
rect -547 3711 -542 3725
rect -546 3710 -542 3711
rect -522 3710 -518 3780
rect -498 3710 -494 3780
rect -474 3710 -470 3780
rect -450 3710 -446 3780
rect -426 3710 -422 3780
rect -402 3710 -398 3780
rect -378 3710 -374 3780
rect -354 3710 -350 3780
rect -330 3710 -326 3780
rect -306 3710 -302 3780
rect -282 3710 -278 3780
rect -258 3710 -254 3780
rect -234 3710 -230 3780
rect -210 3710 -206 3780
rect -186 3710 -182 3780
rect -162 3710 -158 3780
rect -138 3710 -134 3780
rect -114 3710 -110 3780
rect -90 3710 -86 3780
rect -66 3710 -62 3780
rect -42 3710 -38 3780
rect -18 3710 -14 3780
rect 6 3779 10 3780
rect 6 3734 13 3779
rect 30 3734 34 3780
rect 54 3734 58 3780
rect 78 3734 82 3780
rect 102 3734 106 3780
rect 126 3734 130 3780
rect 150 3734 154 3780
rect 174 3734 178 3780
rect 198 3734 202 3780
rect 222 3734 226 3780
rect 246 3734 250 3780
rect 270 3734 274 3780
rect 294 3734 298 3780
rect 318 3734 322 3780
rect 342 3734 346 3780
rect 366 3734 370 3780
rect 390 3734 394 3780
rect 414 3734 418 3780
rect 438 3734 442 3780
rect 462 3734 466 3780
rect 486 3734 490 3780
rect 510 3734 514 3780
rect 534 3734 538 3780
rect 558 3734 562 3780
rect 582 3734 586 3780
rect 606 3734 610 3780
rect 630 3734 634 3780
rect 654 3734 658 3780
rect 678 3734 682 3780
rect 702 3734 706 3780
rect 726 3734 730 3780
rect 750 3734 754 3780
rect 774 3734 778 3780
rect 798 3734 802 3780
rect 822 3734 826 3780
rect 846 3734 850 3780
rect 870 3734 874 3780
rect 894 3734 898 3780
rect 918 3734 922 3780
rect 942 3734 946 3780
rect 966 3734 970 3780
rect 990 3734 994 3780
rect 1014 3734 1018 3780
rect 1038 3734 1042 3780
rect 1062 3734 1066 3780
rect 1086 3734 1090 3780
rect 1110 3734 1114 3780
rect 1134 3734 1138 3780
rect 1158 3734 1162 3780
rect 1182 3734 1186 3780
rect 1206 3734 1210 3780
rect 1230 3734 1234 3780
rect 1254 3734 1258 3780
rect 1278 3734 1282 3780
rect 1302 3734 1306 3780
rect 1326 3734 1330 3780
rect 1350 3734 1354 3780
rect 1374 3734 1378 3780
rect 1398 3734 1402 3780
rect 1422 3734 1426 3780
rect 1446 3734 1450 3780
rect 1470 3734 1474 3780
rect 1494 3734 1498 3780
rect 1518 3734 1522 3780
rect 1542 3734 1546 3780
rect 1566 3734 1570 3780
rect 1590 3734 1594 3780
rect 1614 3734 1618 3780
rect 1638 3734 1642 3780
rect 1662 3734 1666 3780
rect 1686 3734 1690 3780
rect 1710 3734 1714 3780
rect 1734 3734 1738 3780
rect 1758 3734 1762 3780
rect 1782 3734 1786 3780
rect 1806 3734 1810 3780
rect 1830 3734 1834 3780
rect 1854 3734 1858 3780
rect 1878 3734 1882 3780
rect 1902 3734 1906 3780
rect 1926 3734 1930 3780
rect 1950 3734 1954 3780
rect 1974 3734 1978 3780
rect 1998 3734 2002 3780
rect 2022 3734 2026 3780
rect 2046 3734 2050 3780
rect 2070 3734 2074 3780
rect 2094 3734 2098 3780
rect 2118 3734 2122 3780
rect 2142 3734 2146 3780
rect 2166 3734 2170 3780
rect 2190 3734 2194 3780
rect 2214 3734 2218 3780
rect 2238 3734 2242 3780
rect 2251 3773 2256 3780
rect 2261 3759 2266 3773
rect 2262 3735 2266 3759
rect 2251 3734 2285 3735
rect -11 3732 2285 3734
rect -11 3731 3 3732
rect 6 3731 13 3732
rect 6 3710 10 3731
rect 30 3710 34 3732
rect 54 3710 58 3732
rect 78 3710 82 3732
rect 102 3710 106 3732
rect 126 3710 130 3732
rect 150 3710 154 3732
rect 174 3710 178 3732
rect 198 3710 202 3732
rect 222 3710 226 3732
rect 246 3710 250 3732
rect 270 3710 274 3732
rect 294 3710 298 3732
rect 318 3710 322 3732
rect 342 3710 346 3732
rect 366 3710 370 3732
rect 390 3710 394 3732
rect 414 3710 418 3732
rect 438 3710 442 3732
rect 462 3710 466 3732
rect 486 3710 490 3732
rect 510 3710 514 3732
rect 534 3710 538 3732
rect 558 3710 562 3732
rect 582 3710 586 3732
rect 606 3710 610 3732
rect 630 3710 634 3732
rect 654 3710 658 3732
rect 678 3710 682 3732
rect 702 3710 706 3732
rect 726 3710 730 3732
rect 750 3710 754 3732
rect 774 3710 778 3732
rect 798 3710 802 3732
rect 822 3710 826 3732
rect 846 3710 850 3732
rect 870 3710 874 3732
rect 894 3710 898 3732
rect 918 3710 922 3732
rect 942 3710 946 3732
rect 966 3710 970 3732
rect 990 3710 994 3732
rect 1014 3710 1018 3732
rect 1038 3710 1042 3732
rect 1062 3710 1066 3732
rect 1086 3710 1090 3732
rect 1110 3710 1114 3732
rect 1134 3710 1138 3732
rect 1158 3710 1162 3732
rect 1182 3710 1186 3732
rect 1206 3710 1210 3732
rect 1230 3710 1234 3732
rect 1254 3710 1258 3732
rect 1278 3710 1282 3732
rect 1302 3710 1306 3732
rect 1326 3710 1330 3732
rect 1350 3710 1354 3732
rect 1374 3710 1378 3732
rect 1398 3710 1402 3732
rect 1422 3710 1426 3732
rect 1446 3710 1450 3732
rect 1470 3710 1474 3732
rect 1494 3710 1498 3732
rect 1518 3710 1522 3732
rect 1542 3710 1546 3732
rect 1566 3710 1570 3732
rect 1590 3710 1594 3732
rect 1614 3710 1618 3732
rect 1638 3710 1642 3732
rect 1662 3710 1666 3732
rect 1686 3710 1690 3732
rect 1710 3710 1714 3732
rect 1734 3710 1738 3732
rect 1758 3710 1762 3732
rect 1782 3710 1786 3732
rect 1806 3710 1810 3732
rect 1830 3710 1834 3732
rect 1854 3710 1858 3732
rect 1878 3710 1882 3732
rect 1902 3710 1906 3732
rect 1926 3710 1930 3732
rect 1950 3710 1954 3732
rect 1974 3710 1978 3732
rect 1998 3710 2002 3732
rect 2022 3710 2026 3732
rect 2046 3710 2050 3732
rect 2070 3710 2074 3732
rect 2094 3710 2098 3732
rect 2118 3710 2122 3732
rect 2142 3710 2146 3732
rect 2166 3710 2170 3732
rect 2190 3710 2194 3732
rect 2214 3710 2218 3732
rect 2238 3711 2242 3732
rect 2251 3725 2256 3732
rect 2262 3725 2266 3732
rect 2261 3711 2266 3725
rect 2275 3721 2283 3725
rect 2269 3711 2275 3721
rect 2227 3710 2261 3711
rect -893 3708 2261 3710
rect -893 3701 -888 3708
rect -883 3687 -878 3701
rect -882 3686 -878 3687
rect -858 3686 -854 3708
rect -834 3686 -830 3708
rect -810 3686 -806 3708
rect -786 3686 -782 3708
rect -762 3686 -758 3708
rect -738 3686 -734 3708
rect -714 3686 -710 3708
rect -690 3686 -686 3708
rect -666 3686 -662 3708
rect -642 3686 -638 3708
rect -618 3686 -614 3708
rect -594 3686 -590 3708
rect -570 3686 -566 3708
rect -546 3686 -542 3708
rect -522 3686 -518 3708
rect -498 3686 -494 3708
rect -474 3686 -470 3708
rect -450 3686 -446 3708
rect -426 3686 -422 3708
rect -402 3686 -398 3708
rect -378 3686 -374 3708
rect -354 3686 -350 3708
rect -330 3686 -326 3708
rect -306 3686 -302 3708
rect -282 3686 -278 3708
rect -258 3686 -254 3708
rect -234 3686 -230 3708
rect -210 3686 -206 3708
rect -186 3686 -182 3708
rect -162 3686 -158 3708
rect -138 3686 -134 3708
rect -114 3686 -110 3708
rect -90 3686 -86 3708
rect -66 3686 -62 3708
rect -42 3686 -38 3708
rect -18 3686 -14 3708
rect 6 3686 10 3708
rect 30 3686 34 3708
rect 54 3686 58 3708
rect 78 3686 82 3708
rect 102 3686 106 3708
rect 126 3686 130 3708
rect 150 3686 154 3708
rect 174 3686 178 3708
rect 198 3686 202 3708
rect 222 3686 226 3708
rect 246 3686 250 3708
rect 270 3686 274 3708
rect 294 3686 298 3708
rect 318 3686 322 3708
rect 342 3686 346 3708
rect 366 3686 370 3708
rect 390 3686 394 3708
rect 414 3686 418 3708
rect 438 3686 442 3708
rect 462 3686 466 3708
rect 486 3686 490 3708
rect 510 3686 514 3708
rect 534 3686 538 3708
rect 558 3686 562 3708
rect 582 3686 586 3708
rect 606 3686 610 3708
rect 630 3686 634 3708
rect 654 3686 658 3708
rect 678 3686 682 3708
rect 702 3686 706 3708
rect 726 3686 730 3708
rect 750 3686 754 3708
rect 774 3686 778 3708
rect 798 3686 802 3708
rect 822 3686 826 3708
rect 846 3686 850 3708
rect 870 3686 874 3708
rect 894 3686 898 3708
rect 918 3686 922 3708
rect 942 3686 946 3708
rect 966 3686 970 3708
rect 990 3686 994 3708
rect 1014 3686 1018 3708
rect 1038 3686 1042 3708
rect 1062 3686 1066 3708
rect 1086 3686 1090 3708
rect 1110 3686 1114 3708
rect 1134 3686 1138 3708
rect 1158 3686 1162 3708
rect 1182 3686 1186 3708
rect 1206 3686 1210 3708
rect 1230 3686 1234 3708
rect 1254 3686 1258 3708
rect 1278 3686 1282 3708
rect 1302 3686 1306 3708
rect 1326 3686 1330 3708
rect 1350 3686 1354 3708
rect 1374 3686 1378 3708
rect 1398 3686 1402 3708
rect 1422 3686 1426 3708
rect 1446 3686 1450 3708
rect 1470 3686 1474 3708
rect 1494 3686 1498 3708
rect 1518 3686 1522 3708
rect 1542 3686 1546 3708
rect 1566 3686 1570 3708
rect 1590 3686 1594 3708
rect 1614 3686 1618 3708
rect 1638 3686 1642 3708
rect 1662 3686 1666 3708
rect 1686 3686 1690 3708
rect 1710 3686 1714 3708
rect 1734 3686 1738 3708
rect 1758 3686 1762 3708
rect 1782 3686 1786 3708
rect 1806 3686 1810 3708
rect 1830 3686 1834 3708
rect 1854 3686 1858 3708
rect 1878 3686 1882 3708
rect 1902 3686 1906 3708
rect 1926 3686 1930 3708
rect 1950 3686 1954 3708
rect 1974 3686 1978 3708
rect 1998 3686 2002 3708
rect 2022 3686 2026 3708
rect 2046 3686 2050 3708
rect 2070 3686 2074 3708
rect 2094 3686 2098 3708
rect 2118 3686 2122 3708
rect 2142 3686 2146 3708
rect 2166 3686 2170 3708
rect 2190 3686 2194 3708
rect 2214 3686 2218 3708
rect 2227 3701 2232 3708
rect 2238 3701 2242 3708
rect 2237 3687 2242 3701
rect 2227 3686 2261 3687
rect -2393 3684 2261 3686
rect -2371 3662 -2366 3684
rect -2348 3662 -2343 3684
rect -2325 3662 -2320 3684
rect -2072 3682 -2036 3683
rect -2072 3676 -2054 3682
rect -2309 3668 -2301 3676
rect -2317 3662 -2309 3668
rect -2092 3667 -2062 3672
rect -2000 3663 -1992 3684
rect -1938 3683 -1906 3684
rect -1920 3682 -1906 3683
rect -1806 3676 -1680 3682
rect -1854 3667 -1806 3672
rect -1655 3668 -1647 3676
rect -1982 3663 -1966 3664
rect -2000 3662 -1966 3663
rect -1846 3662 -1806 3665
rect -1663 3662 -1655 3668
rect -1642 3662 -1637 3684
rect -1619 3662 -1614 3684
rect -1530 3662 -1526 3684
rect -1506 3662 -1502 3684
rect -1482 3662 -1478 3684
rect -1458 3662 -1454 3684
rect -1434 3662 -1430 3684
rect -1410 3662 -1406 3684
rect -1386 3662 -1382 3684
rect -1362 3662 -1358 3684
rect -1338 3662 -1334 3684
rect -1314 3662 -1310 3684
rect -1290 3662 -1286 3684
rect -1266 3662 -1262 3684
rect -1242 3662 -1238 3684
rect -1218 3662 -1214 3684
rect -1194 3662 -1190 3684
rect -1170 3662 -1166 3684
rect -1146 3662 -1142 3684
rect -1122 3662 -1118 3684
rect -1098 3662 -1094 3684
rect -1074 3662 -1070 3684
rect -1050 3662 -1046 3684
rect -1026 3662 -1022 3684
rect -1002 3662 -998 3684
rect -978 3662 -974 3684
rect -954 3662 -950 3684
rect -930 3662 -926 3684
rect -906 3662 -902 3684
rect -882 3662 -878 3684
rect -858 3662 -854 3684
rect -834 3662 -830 3684
rect -810 3662 -806 3684
rect -786 3662 -782 3684
rect -762 3662 -758 3684
rect -738 3662 -734 3684
rect -714 3662 -710 3684
rect -690 3662 -686 3684
rect -666 3662 -662 3684
rect -642 3662 -638 3684
rect -618 3662 -614 3684
rect -594 3662 -590 3684
rect -570 3662 -566 3684
rect -546 3662 -542 3684
rect -522 3683 -518 3684
rect -2393 3660 -525 3662
rect -2371 3638 -2366 3660
rect -2348 3638 -2343 3660
rect -2325 3638 -2320 3660
rect -2000 3658 -1966 3660
rect -2309 3640 -2301 3648
rect -2062 3647 -2054 3654
rect -2092 3640 -2084 3647
rect -2062 3640 -2026 3642
rect -2317 3638 -2309 3640
rect -2062 3638 -2012 3640
rect -2000 3638 -1992 3658
rect -1982 3657 -1966 3658
rect -1846 3656 -1806 3660
rect -1846 3649 -1798 3654
rect -1806 3647 -1798 3649
rect -1854 3645 -1846 3647
rect -1854 3640 -1806 3645
rect -1655 3640 -1647 3648
rect -1864 3638 -1796 3639
rect -1663 3638 -1655 3640
rect -1642 3638 -1637 3660
rect -1619 3638 -1614 3660
rect -1530 3638 -1526 3660
rect -1506 3638 -1502 3660
rect -1482 3638 -1478 3660
rect -1458 3638 -1454 3660
rect -1434 3638 -1430 3660
rect -1410 3638 -1406 3660
rect -1386 3639 -1382 3660
rect -1397 3638 -1363 3639
rect -2393 3636 -1363 3638
rect -2371 3590 -2366 3636
rect -2348 3590 -2343 3636
rect -2325 3590 -2320 3636
rect -2317 3632 -2309 3636
rect -2062 3632 -2054 3636
rect -2154 3628 -2138 3630
rect -2057 3628 -2054 3632
rect -2292 3622 -2054 3628
rect -2052 3622 -2044 3632
rect -2092 3606 -2062 3608
rect -2094 3602 -2062 3606
rect -2000 3590 -1992 3636
rect -1846 3629 -1806 3636
rect -1663 3632 -1655 3636
rect -1846 3622 -1680 3628
rect -1854 3606 -1806 3608
rect -1854 3602 -1680 3606
rect -1979 3590 -1945 3592
rect -1642 3590 -1637 3636
rect -1619 3590 -1614 3636
rect -1530 3590 -1526 3636
rect -1506 3590 -1502 3636
rect -1482 3590 -1478 3636
rect -1458 3590 -1454 3636
rect -1434 3590 -1430 3636
rect -1410 3590 -1406 3636
rect -1397 3629 -1392 3636
rect -1386 3629 -1382 3636
rect -1387 3615 -1382 3629
rect -1386 3590 -1382 3615
rect -1362 3590 -1358 3660
rect -1338 3590 -1334 3660
rect -1314 3590 -1310 3660
rect -1290 3590 -1286 3660
rect -1266 3590 -1262 3660
rect -1242 3590 -1238 3660
rect -1218 3590 -1214 3660
rect -1194 3590 -1190 3660
rect -1170 3590 -1166 3660
rect -1146 3590 -1142 3660
rect -1122 3590 -1118 3660
rect -1098 3590 -1094 3660
rect -1074 3590 -1070 3660
rect -1050 3590 -1046 3660
rect -1026 3590 -1022 3660
rect -1002 3590 -998 3660
rect -978 3590 -974 3660
rect -954 3590 -950 3660
rect -930 3590 -926 3660
rect -906 3590 -902 3660
rect -882 3590 -878 3660
rect -858 3659 -854 3660
rect -858 3611 -851 3659
rect -858 3590 -854 3611
rect -834 3590 -830 3660
rect -810 3590 -806 3660
rect -786 3590 -782 3660
rect -762 3590 -758 3660
rect -738 3590 -734 3660
rect -714 3590 -710 3660
rect -690 3590 -686 3660
rect -666 3590 -662 3660
rect -642 3590 -638 3660
rect -618 3590 -614 3660
rect -594 3590 -590 3660
rect -570 3590 -566 3660
rect -546 3590 -542 3660
rect -539 3659 -525 3660
rect -522 3635 -515 3683
rect -522 3590 -518 3635
rect -498 3590 -494 3684
rect -474 3590 -470 3684
rect -450 3590 -446 3684
rect -426 3590 -422 3684
rect -402 3590 -398 3684
rect -378 3590 -374 3684
rect -354 3590 -350 3684
rect -330 3590 -326 3684
rect -306 3590 -302 3684
rect -282 3590 -278 3684
rect -258 3590 -254 3684
rect -234 3590 -230 3684
rect -210 3590 -206 3684
rect -186 3590 -182 3684
rect -162 3590 -158 3684
rect -138 3590 -134 3684
rect -125 3653 -120 3663
rect -114 3653 -110 3684
rect -115 3639 -110 3653
rect -125 3638 -91 3639
rect -90 3638 -86 3684
rect -66 3638 -62 3684
rect -42 3638 -38 3684
rect -18 3638 -14 3684
rect 6 3638 10 3684
rect 30 3638 34 3684
rect 54 3638 58 3684
rect 78 3638 82 3684
rect 102 3638 106 3684
rect 126 3638 130 3684
rect 150 3638 154 3684
rect 174 3638 178 3684
rect 198 3638 202 3684
rect 222 3638 226 3684
rect 246 3638 250 3684
rect 270 3638 274 3684
rect 294 3638 298 3684
rect 318 3638 322 3684
rect 342 3638 346 3684
rect 366 3638 370 3684
rect 390 3638 394 3684
rect 414 3638 418 3684
rect 438 3638 442 3684
rect 462 3638 466 3684
rect 486 3638 490 3684
rect 510 3638 514 3684
rect 534 3638 538 3684
rect 558 3638 562 3684
rect 582 3638 586 3684
rect 606 3638 610 3684
rect 630 3638 634 3684
rect 654 3638 658 3684
rect 678 3638 682 3684
rect 702 3638 706 3684
rect 726 3638 730 3684
rect 750 3638 754 3684
rect 774 3638 778 3684
rect 798 3638 802 3684
rect 822 3638 826 3684
rect 846 3638 850 3684
rect 870 3638 874 3684
rect 894 3638 898 3684
rect 918 3638 922 3684
rect 942 3638 946 3684
rect 966 3638 970 3684
rect 990 3638 994 3684
rect 1014 3638 1018 3684
rect 1038 3638 1042 3684
rect 1062 3638 1066 3684
rect 1086 3638 1090 3684
rect 1110 3638 1114 3684
rect 1134 3638 1138 3684
rect 1158 3638 1162 3684
rect 1182 3638 1186 3684
rect 1206 3638 1210 3684
rect 1230 3638 1234 3684
rect 1254 3638 1258 3684
rect 1278 3638 1282 3684
rect 1302 3638 1306 3684
rect 1326 3638 1330 3684
rect 1350 3638 1354 3684
rect 1374 3638 1378 3684
rect 1398 3638 1402 3684
rect 1422 3638 1426 3684
rect 1446 3638 1450 3684
rect 1470 3638 1474 3684
rect 1494 3638 1498 3684
rect 1518 3638 1522 3684
rect 1542 3638 1546 3684
rect 1566 3638 1570 3684
rect 1590 3638 1594 3684
rect 1614 3638 1618 3684
rect 1638 3638 1642 3684
rect 1662 3638 1666 3684
rect 1686 3638 1690 3684
rect 1710 3638 1714 3684
rect 1734 3638 1738 3684
rect 1758 3638 1762 3684
rect 1782 3638 1786 3684
rect 1806 3638 1810 3684
rect 1830 3638 1834 3684
rect 1854 3638 1858 3684
rect 1878 3638 1882 3684
rect 1902 3638 1906 3684
rect 1926 3638 1930 3684
rect 1950 3638 1954 3684
rect 1974 3638 1978 3684
rect 1998 3638 2002 3684
rect 2022 3638 2026 3684
rect 2046 3638 2050 3684
rect 2070 3638 2074 3684
rect 2094 3638 2098 3684
rect 2118 3638 2122 3684
rect 2142 3638 2146 3684
rect 2166 3638 2170 3684
rect 2190 3638 2194 3684
rect 2214 3638 2218 3684
rect 2227 3677 2232 3684
rect 2237 3663 2242 3677
rect 2238 3639 2242 3663
rect 2227 3638 2261 3639
rect -125 3636 2261 3638
rect -125 3629 -120 3636
rect -115 3615 -110 3629
rect -114 3590 -110 3615
rect -90 3590 -86 3636
rect -66 3590 -62 3636
rect -42 3590 -38 3636
rect -18 3590 -14 3636
rect 6 3590 10 3636
rect 30 3590 34 3636
rect 54 3590 58 3636
rect 78 3590 82 3636
rect 102 3590 106 3636
rect 126 3590 130 3636
rect 150 3590 154 3636
rect 174 3590 178 3636
rect 198 3590 202 3636
rect 222 3590 226 3636
rect 246 3590 250 3636
rect 270 3590 274 3636
rect 294 3590 298 3636
rect 318 3590 322 3636
rect 342 3590 346 3636
rect 366 3590 370 3636
rect 390 3590 394 3636
rect 414 3590 418 3636
rect 438 3590 442 3636
rect 462 3590 466 3636
rect 486 3590 490 3636
rect 510 3590 514 3636
rect 534 3590 538 3636
rect 558 3590 562 3636
rect 582 3590 586 3636
rect 606 3590 610 3636
rect 630 3590 634 3636
rect 654 3590 658 3636
rect 678 3590 682 3636
rect 702 3590 706 3636
rect 726 3590 730 3636
rect 750 3590 754 3636
rect 774 3590 778 3636
rect 798 3590 802 3636
rect 822 3590 826 3636
rect 846 3590 850 3636
rect 870 3590 874 3636
rect 894 3590 898 3636
rect 918 3590 922 3636
rect 942 3590 946 3636
rect 966 3590 970 3636
rect 990 3590 994 3636
rect 1014 3590 1018 3636
rect 1038 3590 1042 3636
rect 1062 3590 1066 3636
rect 1086 3590 1090 3636
rect 1110 3590 1114 3636
rect 1134 3590 1138 3636
rect 1158 3590 1162 3636
rect 1182 3590 1186 3636
rect 1206 3590 1210 3636
rect 1230 3590 1234 3636
rect 1254 3590 1258 3636
rect 1278 3590 1282 3636
rect 1302 3590 1306 3636
rect 1326 3590 1330 3636
rect 1350 3590 1354 3636
rect 1374 3590 1378 3636
rect 1398 3590 1402 3636
rect 1422 3590 1426 3636
rect 1446 3590 1450 3636
rect 1470 3590 1474 3636
rect 1494 3590 1498 3636
rect 1518 3590 1522 3636
rect 1542 3590 1546 3636
rect 1566 3590 1570 3636
rect 1590 3590 1594 3636
rect 1614 3590 1618 3636
rect 1638 3590 1642 3636
rect 1662 3590 1666 3636
rect 1686 3590 1690 3636
rect 1710 3590 1714 3636
rect 1734 3590 1738 3636
rect 1758 3590 1762 3636
rect 1782 3590 1786 3636
rect 1806 3590 1810 3636
rect 1830 3590 1834 3636
rect 1854 3590 1858 3636
rect 1878 3590 1882 3636
rect 1902 3590 1906 3636
rect 1926 3590 1930 3636
rect 1950 3590 1954 3636
rect 1974 3590 1978 3636
rect 1998 3590 2002 3636
rect 2022 3590 2026 3636
rect 2046 3590 2050 3636
rect 2070 3590 2074 3636
rect 2094 3590 2098 3636
rect 2118 3590 2122 3636
rect 2142 3590 2146 3636
rect 2166 3590 2170 3636
rect 2190 3590 2194 3636
rect 2214 3590 2218 3636
rect 2227 3629 2232 3636
rect 2238 3629 2242 3636
rect 2237 3615 2242 3629
rect 2251 3625 2259 3629
rect 2245 3615 2251 3625
rect 2227 3590 2259 3591
rect -2393 3588 2259 3590
rect -2371 3542 -2366 3588
rect -2348 3542 -2343 3588
rect -2325 3542 -2320 3588
rect -2080 3587 -1906 3588
rect -2080 3586 -2036 3587
rect -2080 3580 -2054 3586
rect -2309 3572 -2301 3578
rect -2317 3562 -2309 3572
rect -2070 3571 -2040 3578
rect -2054 3563 -2040 3566
rect -2000 3561 -1992 3587
rect -1920 3586 -1906 3587
rect -1850 3580 -1846 3588
rect -1840 3580 -1792 3588
rect -1969 3568 -1966 3577
rect -1850 3573 -1802 3578
rect -1906 3571 -1802 3573
rect -1655 3572 -1647 3578
rect -1906 3570 -1850 3571
rect -1846 3563 -1802 3569
rect -1663 3562 -1655 3572
rect -1860 3561 -1798 3562
rect -2078 3554 -2070 3561
rect -2309 3544 -2301 3550
rect -2317 3542 -2309 3544
rect -2154 3542 -2145 3552
rect -2044 3551 -2040 3556
rect -2028 3554 -1945 3561
rect -1929 3554 -1794 3561
rect -2070 3544 -2040 3551
rect -2044 3542 -2028 3544
rect -2000 3542 -1992 3554
rect -1860 3553 -1798 3554
rect -1850 3544 -1802 3551
rect -1655 3544 -1647 3550
rect -1978 3542 -1942 3543
rect -1663 3542 -1655 3544
rect -1642 3542 -1637 3588
rect -1619 3542 -1614 3588
rect -1530 3542 -1526 3588
rect -1506 3542 -1502 3588
rect -1482 3542 -1478 3588
rect -1458 3542 -1454 3588
rect -1434 3542 -1430 3588
rect -1410 3542 -1406 3588
rect -1386 3542 -1382 3588
rect -1362 3563 -1358 3588
rect -2393 3540 -1365 3542
rect -2371 3446 -2366 3540
rect -2348 3446 -2343 3540
rect -2325 3502 -2320 3540
rect -2317 3534 -2309 3540
rect -2145 3536 -2138 3540
rect -2070 3536 -2054 3540
rect -2078 3527 -2054 3534
rect -2062 3502 -2032 3503
rect -2000 3502 -1992 3540
rect -1846 3536 -1802 3540
rect -1846 3526 -1792 3535
rect -1663 3534 -1655 3540
rect -1942 3504 -1937 3516
rect -1850 3513 -1822 3514
rect -1850 3509 -1802 3513
rect -2325 3494 -2317 3502
rect -2062 3500 -1961 3502
rect -2325 3446 -2320 3494
rect -2317 3486 -2309 3494
rect -2062 3487 -2040 3498
rect -2032 3493 -1961 3500
rect -1947 3494 -1942 3502
rect -1842 3500 -1794 3503
rect -2070 3482 -2022 3486
rect -2000 3448 -1992 3493
rect -1942 3492 -1937 3494
rect -1932 3484 -1927 3492
rect -1912 3489 -1896 3495
rect -1842 3487 -1802 3498
rect -1671 3494 -1663 3502
rect -1663 3486 -1655 3494
rect -1850 3482 -1680 3486
rect -2000 3446 -1957 3448
rect -1642 3446 -1637 3540
rect -1619 3446 -1614 3540
rect -1530 3446 -1526 3540
rect -1506 3446 -1502 3540
rect -1482 3446 -1478 3540
rect -1458 3446 -1454 3540
rect -1434 3446 -1430 3540
rect -1410 3446 -1406 3540
rect -1397 3509 -1392 3519
rect -1386 3509 -1382 3540
rect -1379 3539 -1365 3540
rect -1362 3539 -1355 3563
rect -1387 3495 -1382 3509
rect -1397 3494 -1363 3495
rect -1362 3494 -1358 3539
rect -1338 3494 -1334 3588
rect -1314 3494 -1310 3588
rect -1290 3494 -1286 3588
rect -1266 3494 -1262 3588
rect -1242 3494 -1238 3588
rect -1218 3494 -1214 3588
rect -1194 3494 -1190 3588
rect -1170 3494 -1166 3588
rect -1146 3494 -1142 3588
rect -1122 3494 -1118 3588
rect -1098 3494 -1094 3588
rect -1074 3494 -1070 3588
rect -1050 3494 -1046 3588
rect -1026 3494 -1022 3588
rect -1002 3494 -998 3588
rect -978 3494 -974 3588
rect -954 3494 -950 3588
rect -930 3494 -926 3588
rect -906 3494 -902 3588
rect -882 3494 -878 3588
rect -858 3494 -854 3588
rect -834 3494 -830 3588
rect -810 3494 -806 3588
rect -786 3494 -782 3588
rect -762 3494 -758 3588
rect -738 3494 -734 3588
rect -714 3494 -710 3588
rect -690 3494 -686 3588
rect -666 3494 -662 3588
rect -642 3494 -638 3588
rect -618 3494 -614 3588
rect -594 3494 -590 3588
rect -570 3494 -566 3588
rect -546 3494 -542 3588
rect -522 3494 -518 3588
rect -498 3494 -494 3588
rect -474 3494 -470 3588
rect -450 3494 -446 3588
rect -437 3533 -432 3543
rect -426 3533 -422 3588
rect -427 3519 -422 3533
rect -437 3509 -432 3519
rect -427 3495 -422 3509
rect -426 3494 -422 3495
rect -402 3494 -398 3588
rect -378 3494 -374 3588
rect -354 3494 -350 3588
rect -330 3494 -326 3588
rect -306 3494 -302 3588
rect -282 3494 -278 3588
rect -258 3494 -254 3588
rect -234 3494 -230 3588
rect -210 3494 -206 3588
rect -186 3494 -182 3588
rect -162 3494 -158 3588
rect -138 3494 -134 3588
rect -114 3494 -110 3588
rect -90 3587 -86 3588
rect -90 3539 -83 3587
rect -90 3494 -86 3539
rect -66 3494 -62 3588
rect -42 3494 -38 3588
rect -18 3494 -14 3588
rect 6 3494 10 3588
rect 30 3494 34 3588
rect 54 3494 58 3588
rect 78 3494 82 3588
rect 102 3494 106 3588
rect 126 3494 130 3588
rect 150 3494 154 3588
rect 174 3494 178 3588
rect 198 3494 202 3588
rect 222 3494 226 3588
rect 246 3494 250 3588
rect 270 3494 274 3588
rect 294 3494 298 3588
rect 318 3494 322 3588
rect 342 3494 346 3588
rect 366 3494 370 3588
rect 390 3494 394 3588
rect 414 3494 418 3588
rect 438 3494 442 3588
rect 462 3494 466 3588
rect 486 3494 490 3588
rect 510 3494 514 3588
rect 534 3494 538 3588
rect 558 3494 562 3588
rect 582 3494 586 3588
rect 606 3494 610 3588
rect 630 3494 634 3588
rect 654 3494 658 3588
rect 678 3494 682 3588
rect 702 3494 706 3588
rect 726 3494 730 3588
rect 750 3494 754 3588
rect 774 3494 778 3588
rect 798 3494 802 3588
rect 822 3494 826 3588
rect 846 3494 850 3588
rect 870 3494 874 3588
rect 894 3494 898 3588
rect 918 3494 922 3588
rect 942 3494 946 3588
rect 966 3494 970 3588
rect 990 3494 994 3588
rect 1014 3494 1018 3588
rect 1038 3494 1042 3588
rect 1062 3494 1066 3588
rect 1086 3494 1090 3588
rect 1110 3494 1114 3588
rect 1134 3494 1138 3588
rect 1158 3494 1162 3588
rect 1182 3494 1186 3588
rect 1206 3494 1210 3588
rect 1230 3494 1234 3588
rect 1254 3494 1258 3588
rect 1278 3494 1282 3588
rect 1302 3494 1306 3588
rect 1326 3494 1330 3588
rect 1350 3494 1354 3588
rect 1374 3494 1378 3588
rect 1398 3494 1402 3588
rect 1422 3494 1426 3588
rect 1446 3494 1450 3588
rect 1470 3494 1474 3588
rect 1494 3494 1498 3588
rect 1518 3494 1522 3588
rect 1542 3494 1546 3588
rect 1566 3494 1570 3588
rect 1590 3494 1594 3588
rect 1614 3494 1618 3588
rect 1638 3494 1642 3588
rect 1662 3494 1666 3588
rect 1686 3494 1690 3588
rect 1710 3494 1714 3588
rect 1734 3494 1738 3588
rect 1758 3494 1762 3588
rect 1782 3494 1786 3588
rect 1806 3494 1810 3588
rect 1830 3494 1834 3588
rect 1854 3494 1858 3588
rect 1878 3494 1882 3588
rect 1902 3494 1906 3588
rect 1926 3494 1930 3588
rect 1950 3494 1954 3588
rect 1974 3494 1978 3588
rect 1998 3494 2002 3588
rect 2022 3494 2026 3588
rect 2046 3494 2050 3588
rect 2070 3494 2074 3588
rect 2094 3494 2098 3588
rect 2118 3494 2122 3588
rect 2142 3494 2146 3588
rect 2166 3494 2170 3588
rect 2190 3494 2194 3588
rect 2214 3495 2218 3588
rect 2227 3581 2232 3588
rect 2245 3587 2259 3588
rect 2237 3567 2242 3581
rect 2227 3509 2232 3519
rect 2238 3509 2242 3567
rect 2237 3495 2242 3509
rect 2251 3505 2259 3509
rect 2245 3495 2251 3505
rect 2203 3494 2237 3495
rect -1397 3492 2237 3494
rect -1397 3485 -1392 3492
rect -1387 3471 -1382 3485
rect -1386 3446 -1382 3471
rect -1362 3446 -1358 3492
rect -1338 3446 -1334 3492
rect -1314 3446 -1310 3492
rect -1290 3446 -1286 3492
rect -1266 3446 -1262 3492
rect -1242 3446 -1238 3492
rect -1218 3446 -1214 3492
rect -1194 3446 -1190 3492
rect -1170 3446 -1166 3492
rect -1146 3446 -1142 3492
rect -1122 3446 -1118 3492
rect -1098 3446 -1094 3492
rect -1074 3446 -1070 3492
rect -1050 3446 -1046 3492
rect -1026 3446 -1022 3492
rect -1002 3446 -998 3492
rect -978 3446 -974 3492
rect -954 3446 -950 3492
rect -930 3446 -926 3492
rect -906 3446 -902 3492
rect -882 3446 -878 3492
rect -858 3446 -854 3492
rect -834 3446 -830 3492
rect -810 3446 -806 3492
rect -786 3446 -782 3492
rect -762 3446 -758 3492
rect -738 3446 -734 3492
rect -714 3446 -710 3492
rect -690 3446 -686 3492
rect -666 3446 -662 3492
rect -642 3446 -638 3492
rect -618 3446 -614 3492
rect -594 3446 -590 3492
rect -570 3446 -566 3492
rect -546 3446 -542 3492
rect -522 3446 -518 3492
rect -498 3446 -494 3492
rect -474 3446 -470 3492
rect -450 3446 -446 3492
rect -426 3446 -422 3492
rect -402 3467 -398 3492
rect -2393 3444 -405 3446
rect -2371 2918 -2366 3444
rect -2348 2918 -2343 3444
rect -2325 3370 -2320 3444
rect -2317 3430 -2309 3444
rect -2317 3402 -2309 3418
rect -2062 3406 -2032 3410
rect -2325 3362 -2317 3370
rect -2325 3342 -2320 3362
rect -2317 3354 -2309 3362
rect -2325 3334 -2317 3342
rect -2325 3314 -2320 3334
rect -2317 3326 -2309 3334
rect -2127 3322 -2097 3323
rect -2325 3306 -2317 3314
rect -2325 3286 -2320 3306
rect -2317 3299 -2309 3306
rect -2127 3302 -2124 3311
rect -2119 3302 -2097 3315
rect -2092 3309 -2089 3315
rect -2087 3312 -2079 3325
rect -2127 3301 -2097 3302
rect -2317 3298 -2301 3299
rect -2309 3287 -2307 3298
rect -2145 3290 -2129 3297
rect -2066 3296 -2065 3297
rect -2325 3278 -2317 3286
rect -2325 3154 -2320 3278
rect -2317 3270 -2309 3278
rect -2297 3271 -2289 3287
rect -2150 3285 -2141 3287
rect -2129 3285 -2113 3287
rect -2119 3276 -2113 3285
rect -2125 3271 -2113 3276
rect -2101 3283 -2085 3287
rect -2101 3271 -2089 3283
rect -2317 3214 -2309 3230
rect -2317 3186 -2309 3202
rect -2193 3197 -2189 3207
rect -2199 3195 -2189 3197
rect -2177 3197 -2163 3207
rect -2177 3195 -2161 3197
rect -2325 3146 -2317 3154
rect -2325 3126 -2320 3146
rect -2317 3138 -2309 3146
rect -2325 3118 -2317 3126
rect -2325 3098 -2320 3118
rect -2317 3110 -2309 3118
rect -2127 3106 -2097 3107
rect -2325 3090 -2317 3098
rect -2325 3070 -2320 3090
rect -2317 3083 -2309 3090
rect -2127 3086 -2124 3095
rect -2119 3086 -2097 3099
rect -2092 3093 -2089 3099
rect -2087 3096 -2079 3109
rect -2127 3085 -2097 3086
rect -2317 3082 -2301 3083
rect -2309 3071 -2307 3082
rect -2145 3074 -2129 3081
rect -2066 3080 -2065 3081
rect -2325 3062 -2317 3070
rect -2325 3042 -2320 3062
rect -2317 3054 -2309 3062
rect -2297 3055 -2289 3071
rect -2150 3069 -2141 3071
rect -2129 3069 -2113 3071
rect -2119 3060 -2113 3069
rect -2125 3055 -2113 3060
rect -2101 3067 -2085 3071
rect -2101 3055 -2089 3067
rect -2325 3026 -2317 3042
rect -2325 3010 -2320 3026
rect -2309 3014 -2301 3026
rect -2317 3010 -2309 3014
rect -2325 2998 -2317 3010
rect -2103 3009 -2089 3012
rect -2036 3010 -2028 3014
rect -2079 3006 -2066 3010
rect -2061 3006 -2028 3010
rect -2325 2982 -2320 2998
rect -2309 2986 -2301 2998
rect -2066 2997 -2061 3000
rect -2093 2991 -2077 2995
rect -2317 2982 -2309 2986
rect -2121 2983 -2105 2985
rect -2093 2983 -2092 2985
rect -2091 2983 -2077 2991
rect -2058 2983 -2049 2997
rect -2018 2996 -2004 3004
rect -2018 2990 -2012 2996
rect -2292 2982 -2049 2983
rect -2036 2982 -2028 2990
rect -2325 2970 -2317 2982
rect -2292 2979 -2028 2982
rect -2020 2980 -2018 2990
rect -2026 2979 -2018 2980
rect -2325 2950 -2320 2970
rect -2325 2942 -2317 2950
rect -2325 2922 -2320 2942
rect -2317 2934 -2309 2942
rect -2325 2918 -2317 2922
rect -2000 2918 -1992 3444
rect -1974 3442 -1957 3444
rect -1960 3441 -1957 3442
rect -1832 3433 -1794 3434
rect -1663 3430 -1655 3444
rect -1824 3424 -1794 3426
rect -1954 3420 -1918 3424
rect -1904 3415 -1901 3424
rect -1794 3423 -1786 3424
rect -1904 3413 -1888 3415
rect -1822 3410 -1794 3422
rect -1857 3400 -1848 3410
rect -1842 3406 -1794 3410
rect -1663 3402 -1655 3418
rect -1847 3397 -1838 3400
rect -1671 3362 -1663 3370
rect -1663 3354 -1655 3362
rect -1946 3340 -1893 3348
rect -1927 3330 -1919 3338
rect -1901 3330 -1898 3340
rect -1671 3334 -1663 3342
rect -1927 3324 -1920 3330
rect -1936 3322 -1920 3324
rect -1919 3329 -1911 3330
rect -1919 3322 -1903 3329
rect -1901 3323 -1900 3330
rect -1663 3326 -1655 3334
rect -1901 3322 -1853 3323
rect -1893 3302 -1853 3315
rect -1671 3306 -1663 3314
rect -1901 3301 -1853 3302
rect -1663 3298 -1655 3306
rect -1915 3290 -1914 3297
rect -1767 3290 -1766 3297
rect -1671 3278 -1663 3286
rect -1663 3270 -1655 3278
rect -1977 3222 -1972 3232
rect -1663 3214 -1655 3230
rect -1972 3208 -1967 3211
rect -1944 3195 -1928 3198
rect -1927 3195 -1924 3198
rect -1663 3186 -1655 3202
rect -1671 3146 -1663 3154
rect -1663 3138 -1655 3146
rect -1946 3124 -1893 3132
rect -1927 3114 -1919 3122
rect -1901 3114 -1898 3124
rect -1671 3118 -1663 3126
rect -1927 3108 -1920 3114
rect -1936 3106 -1920 3108
rect -1919 3113 -1911 3114
rect -1919 3106 -1903 3113
rect -1901 3107 -1900 3114
rect -1663 3110 -1655 3118
rect -1901 3106 -1853 3107
rect -1893 3086 -1853 3099
rect -1671 3090 -1663 3098
rect -1901 3085 -1853 3086
rect -1663 3082 -1655 3090
rect -1915 3074 -1914 3081
rect -1767 3074 -1766 3081
rect -1671 3062 -1663 3070
rect -1663 3054 -1655 3062
rect -1671 3026 -1663 3042
rect -1655 3014 -1647 3026
rect -1663 3010 -1655 3014
rect -1980 2997 -1932 3000
rect -1671 2998 -1663 3010
rect -1972 2984 -1932 2995
rect -1655 2986 -1647 2998
rect -1972 2979 -1680 2983
rect -1663 2982 -1655 2986
rect -1671 2970 -1663 2982
rect -1671 2942 -1663 2950
rect -1663 2934 -1655 2942
rect -1671 2918 -1663 2922
rect -1642 2918 -1637 3444
rect -1619 2918 -1614 3444
rect -1530 2918 -1526 3444
rect -1506 2918 -1502 3444
rect -1482 2918 -1478 3444
rect -1458 2918 -1454 3444
rect -1434 2918 -1430 3444
rect -1410 2918 -1406 3444
rect -1386 2918 -1382 3444
rect -1362 3443 -1358 3444
rect -1362 3395 -1355 3443
rect -1362 2918 -1358 3395
rect -1338 2918 -1334 3444
rect -1314 2918 -1310 3444
rect -1290 2918 -1286 3444
rect -1266 2918 -1262 3444
rect -1242 2918 -1238 3444
rect -1218 2918 -1214 3444
rect -1194 2918 -1190 3444
rect -1170 2918 -1166 3444
rect -1146 2918 -1142 3444
rect -1122 2918 -1118 3444
rect -1098 2918 -1094 3444
rect -1074 2918 -1070 3444
rect -1050 2918 -1046 3444
rect -1037 3221 -1032 3231
rect -1026 3221 -1022 3444
rect -1027 3207 -1022 3221
rect -1026 2918 -1022 3207
rect -1002 3155 -998 3444
rect -1002 3131 -995 3155
rect -1002 2918 -998 3131
rect -978 2918 -974 3444
rect -954 2918 -950 3444
rect -930 2918 -926 3444
rect -906 2918 -902 3444
rect -882 2918 -878 3444
rect -858 2918 -854 3444
rect -834 2918 -830 3444
rect -810 2918 -806 3444
rect -786 2918 -782 3444
rect -762 2918 -758 3444
rect -738 2918 -734 3444
rect -714 2918 -710 3444
rect -690 2918 -686 3444
rect -666 2918 -662 3444
rect -642 2918 -638 3444
rect -618 2918 -614 3444
rect -594 2918 -590 3444
rect -570 2918 -566 3444
rect -546 2918 -542 3444
rect -522 2918 -518 3444
rect -498 2918 -494 3444
rect -474 2918 -470 3444
rect -450 2918 -446 3444
rect -426 2918 -422 3444
rect -419 3443 -405 3444
rect -402 3419 -395 3467
rect -402 2918 -398 3419
rect -378 2918 -374 3492
rect -354 2918 -350 3492
rect -330 2918 -326 3492
rect -306 2918 -302 3492
rect -282 2918 -278 3492
rect -258 2918 -254 3492
rect -234 2918 -230 3492
rect -210 2918 -206 3492
rect -186 2918 -182 3492
rect -162 2918 -158 3492
rect -138 2918 -134 3492
rect -114 2918 -110 3492
rect -90 2918 -86 3492
rect -66 2918 -62 3492
rect -42 2918 -38 3492
rect -18 2918 -14 3492
rect 6 2918 10 3492
rect 30 2918 34 3492
rect 54 2918 58 3492
rect 78 2918 82 3492
rect 102 2918 106 3492
rect 126 2918 130 3492
rect 150 2918 154 3492
rect 174 2918 178 3492
rect 198 2918 202 3492
rect 222 2918 226 3492
rect 246 2918 250 3492
rect 270 2918 274 3492
rect 294 2918 298 3492
rect 318 2918 322 3492
rect 331 3365 336 3375
rect 342 3365 346 3492
rect 341 3351 346 3365
rect 331 3149 336 3159
rect 342 3149 346 3351
rect 341 3135 346 3149
rect 366 3299 370 3492
rect 366 3275 373 3299
rect 331 3125 336 3135
rect 341 3111 346 3125
rect 342 2918 346 3111
rect 366 3083 370 3275
rect 366 3035 373 3083
rect 366 2918 370 3035
rect 390 2918 394 3492
rect 414 2918 418 3492
rect 438 2918 442 3492
rect 462 2918 466 3492
rect 486 2918 490 3492
rect 510 2918 514 3492
rect 534 2918 538 3492
rect 558 2918 562 3492
rect 582 2918 586 3492
rect 606 2918 610 3492
rect 630 2918 634 3492
rect 654 2918 658 3492
rect 667 3293 672 3303
rect 678 3293 682 3492
rect 677 3279 682 3293
rect 667 3269 672 3279
rect 677 3255 682 3269
rect 667 2957 672 2967
rect 678 2957 682 3255
rect 677 2943 682 2957
rect 702 3227 706 3492
rect 702 3179 709 3227
rect 667 2933 672 2943
rect 677 2919 682 2933
rect 678 2918 682 2919
rect 702 2918 706 3179
rect 715 3077 720 3087
rect 726 3077 730 3492
rect 725 3063 730 3077
rect 726 2918 730 3063
rect 750 3011 754 3492
rect 750 2987 757 3011
rect 750 2918 754 2987
rect 774 2918 778 3492
rect 798 2918 802 3492
rect 822 2918 826 3492
rect 846 2918 850 3492
rect 870 2918 874 3492
rect 894 2918 898 3492
rect 918 2918 922 3492
rect 942 2918 946 3492
rect 966 2918 970 3492
rect 990 2918 994 3492
rect 1014 2918 1018 3492
rect 1038 2918 1042 3492
rect 1062 2918 1066 3492
rect 1086 2918 1090 3492
rect 1110 2918 1114 3492
rect 1134 2918 1138 3492
rect 1158 2918 1162 3492
rect 1182 2918 1186 3492
rect 1206 2918 1210 3492
rect 1230 2918 1234 3492
rect 1254 2918 1258 3492
rect 1278 2918 1282 3492
rect 1302 2918 1306 3492
rect 1326 2918 1330 3492
rect 1350 2918 1354 3492
rect 1374 2918 1378 3492
rect 1398 2918 1402 3492
rect 1422 2918 1426 3492
rect 1446 2918 1450 3492
rect 1470 2918 1474 3492
rect 1494 2918 1498 3492
rect 1518 2918 1522 3492
rect 1542 2918 1546 3492
rect 1566 2918 1570 3492
rect 1590 2918 1594 3492
rect 1614 2918 1618 3492
rect 1638 2918 1642 3492
rect 1662 2918 1666 3492
rect 1686 2918 1690 3492
rect 1710 2918 1714 3492
rect 1734 2918 1738 3492
rect 1758 2918 1762 3492
rect 1782 2918 1786 3492
rect 1806 2918 1810 3492
rect 1830 2918 1834 3492
rect 1854 2918 1858 3492
rect 1878 2918 1882 3492
rect 1902 2918 1906 3492
rect 1926 2918 1930 3492
rect 1950 2918 1954 3492
rect 1974 2918 1978 3492
rect 1998 2918 2002 3492
rect 2022 2918 2026 3492
rect 2046 2918 2050 3492
rect 2070 2918 2074 3492
rect 2094 2918 2098 3492
rect 2118 2918 2122 3492
rect 2131 3437 2136 3447
rect 2142 3437 2146 3492
rect 2141 3423 2146 3437
rect 2131 3422 2165 3423
rect 2166 3422 2170 3492
rect 2190 3423 2194 3492
rect 2203 3485 2208 3492
rect 2214 3485 2218 3492
rect 2213 3471 2218 3485
rect 2179 3422 2213 3423
rect 2131 3420 2213 3422
rect 2131 3413 2136 3420
rect 2141 3399 2146 3413
rect 2131 3125 2136 3135
rect 2142 3125 2146 3399
rect 2166 3371 2170 3420
rect 2179 3413 2184 3420
rect 2190 3413 2194 3420
rect 2189 3399 2194 3413
rect 2166 3323 2173 3371
rect 2155 3269 2160 3279
rect 2166 3269 2170 3323
rect 2165 3255 2170 3269
rect 2141 3111 2146 3125
rect 2131 3005 2136 3015
rect 2141 2991 2146 3005
rect 2131 2933 2136 2943
rect 2142 2933 2146 2991
rect 2141 2919 2146 2933
rect 2155 2929 2163 2933
rect 2149 2919 2155 2929
rect 2131 2918 2163 2919
rect -2393 2916 -1969 2918
rect -1955 2916 2163 2918
rect -2371 2870 -2366 2916
rect -2348 2870 -2343 2916
rect -2325 2906 -2317 2916
rect -2080 2914 -1969 2916
rect -2080 2908 -2053 2914
rect -2325 2890 -2320 2906
rect -2309 2894 -2301 2906
rect -2070 2899 -2040 2906
rect -2000 2898 -1992 2914
rect -1972 2910 -1969 2914
rect -1972 2908 -1955 2910
rect -1955 2898 -1850 2907
rect -1671 2906 -1663 2916
rect -2317 2890 -2309 2894
rect -2070 2891 -2053 2897
rect -2027 2896 -1992 2898
rect -1969 2896 -1955 2897
rect -2325 2878 -2317 2890
rect -2292 2881 -2053 2890
rect -2325 2870 -2320 2878
rect -2309 2870 -2301 2878
rect -2000 2870 -1992 2896
rect -1655 2894 -1647 2906
rect -1663 2890 -1655 2894
rect -1972 2882 -1924 2889
rect -1945 2881 -1929 2882
rect -1860 2881 -1680 2890
rect -1671 2878 -1663 2890
rect -1978 2870 -1942 2871
rect -1655 2870 -1647 2878
rect -1642 2870 -1637 2916
rect -1619 2870 -1614 2916
rect -1530 2870 -1526 2916
rect -1506 2870 -1502 2916
rect -1482 2870 -1478 2916
rect -1458 2870 -1454 2916
rect -1434 2870 -1430 2916
rect -1410 2870 -1406 2916
rect -1386 2870 -1382 2916
rect -1362 2870 -1358 2916
rect -1338 2870 -1334 2916
rect -1314 2870 -1310 2916
rect -1290 2870 -1286 2916
rect -1266 2870 -1262 2916
rect -1242 2870 -1238 2916
rect -1218 2870 -1214 2916
rect -1194 2870 -1190 2916
rect -1170 2870 -1166 2916
rect -1146 2870 -1142 2916
rect -1122 2870 -1118 2916
rect -1098 2870 -1094 2916
rect -1074 2870 -1070 2916
rect -1050 2870 -1046 2916
rect -1026 2870 -1022 2916
rect -1002 2870 -998 2916
rect -978 2870 -974 2916
rect -954 2870 -950 2916
rect -930 2870 -926 2916
rect -906 2870 -902 2916
rect -882 2870 -878 2916
rect -858 2870 -854 2916
rect -834 2870 -830 2916
rect -810 2870 -806 2916
rect -786 2870 -782 2916
rect -762 2870 -758 2916
rect -738 2870 -734 2916
rect -714 2870 -710 2916
rect -690 2870 -686 2916
rect -666 2870 -662 2916
rect -642 2870 -638 2916
rect -618 2870 -614 2916
rect -594 2870 -590 2916
rect -570 2870 -566 2916
rect -546 2870 -542 2916
rect -522 2870 -518 2916
rect -498 2870 -494 2916
rect -474 2870 -470 2916
rect -450 2870 -446 2916
rect -426 2870 -422 2916
rect -402 2870 -398 2916
rect -378 2870 -374 2916
rect -354 2870 -350 2916
rect -330 2870 -326 2916
rect -306 2870 -302 2916
rect -282 2870 -278 2916
rect -258 2870 -254 2916
rect -234 2870 -230 2916
rect -210 2870 -206 2916
rect -186 2870 -182 2916
rect -162 2870 -158 2916
rect -138 2870 -134 2916
rect -114 2870 -110 2916
rect -90 2870 -86 2916
rect -66 2870 -62 2916
rect -42 2870 -38 2916
rect -18 2870 -14 2916
rect 6 2870 10 2916
rect 30 2870 34 2916
rect 54 2870 58 2916
rect 78 2870 82 2916
rect 102 2870 106 2916
rect 126 2870 130 2916
rect 150 2870 154 2916
rect 174 2870 178 2916
rect 198 2870 202 2916
rect 222 2870 226 2916
rect 246 2870 250 2916
rect 270 2870 274 2916
rect 294 2870 298 2916
rect 318 2870 322 2916
rect 342 2870 346 2916
rect 366 2870 370 2916
rect 390 2870 394 2916
rect 414 2870 418 2916
rect 438 2870 442 2916
rect 462 2870 466 2916
rect 486 2870 490 2916
rect 510 2870 514 2916
rect 534 2870 538 2916
rect 558 2870 562 2916
rect 582 2870 586 2916
rect 606 2870 610 2916
rect 630 2870 634 2916
rect 654 2870 658 2916
rect 678 2870 682 2916
rect 702 2891 706 2916
rect -2393 2868 699 2870
rect -2371 2774 -2366 2868
rect -2348 2774 -2343 2868
rect -2325 2862 -2320 2868
rect -2309 2866 -2301 2868
rect -2317 2862 -2309 2866
rect -2325 2850 -2317 2862
rect -2325 2830 -2320 2850
rect -2062 2830 -2032 2831
rect -2000 2830 -1992 2868
rect -1655 2866 -1647 2868
rect -1663 2862 -1655 2866
rect -1671 2850 -1663 2862
rect -1942 2832 -1937 2844
rect -1850 2841 -1822 2842
rect -1850 2837 -1802 2841
rect -2325 2822 -2317 2830
rect -2062 2828 -1961 2830
rect -2325 2802 -2320 2822
rect -2317 2814 -2309 2822
rect -2062 2815 -2040 2826
rect -2032 2821 -1961 2828
rect -1947 2822 -1942 2830
rect -1842 2828 -1794 2831
rect -2070 2810 -2022 2814
rect -2325 2790 -2317 2802
rect -2325 2774 -2320 2790
rect -2317 2786 -2309 2790
rect -2309 2774 -2301 2786
rect -2068 2779 -2038 2786
rect -2000 2776 -1992 2821
rect -1942 2820 -1937 2822
rect -1932 2812 -1927 2820
rect -1912 2817 -1896 2823
rect -1842 2815 -1802 2826
rect -1671 2822 -1663 2830
rect -1663 2814 -1655 2822
rect -1850 2810 -1680 2814
rect -1937 2796 -1934 2798
rect -1926 2796 -1921 2801
rect -1926 2791 -1924 2796
rect -1916 2788 -1914 2791
rect -1842 2788 -1794 2797
rect -1671 2790 -1663 2802
rect -1924 2778 -1916 2787
rect -1663 2786 -1655 2790
rect -1852 2779 -1804 2786
rect -1916 2777 -1914 2778
rect -2025 2775 -1991 2776
rect -2025 2774 -1975 2775
rect -1842 2774 -1804 2777
rect -1655 2774 -1647 2786
rect -1642 2774 -1637 2868
rect -1619 2774 -1614 2868
rect -1530 2774 -1526 2868
rect -1506 2774 -1502 2868
rect -1482 2774 -1478 2868
rect -1458 2774 -1454 2868
rect -1434 2774 -1430 2868
rect -1410 2774 -1406 2868
rect -1386 2774 -1382 2868
rect -1362 2774 -1358 2868
rect -1338 2774 -1334 2868
rect -1314 2774 -1310 2868
rect -1290 2774 -1286 2868
rect -1266 2774 -1262 2868
rect -1242 2774 -1238 2868
rect -1218 2774 -1214 2868
rect -1194 2774 -1190 2868
rect -1170 2774 -1166 2868
rect -1146 2774 -1142 2868
rect -1122 2774 -1118 2868
rect -1098 2774 -1094 2868
rect -1074 2774 -1070 2868
rect -1050 2774 -1046 2868
rect -1026 2774 -1022 2868
rect -1002 2774 -998 2868
rect -978 2774 -974 2868
rect -954 2774 -950 2868
rect -930 2774 -926 2868
rect -906 2774 -902 2868
rect -882 2774 -878 2868
rect -858 2774 -854 2868
rect -834 2774 -830 2868
rect -810 2774 -806 2868
rect -786 2774 -782 2868
rect -762 2774 -758 2868
rect -738 2774 -734 2868
rect -714 2774 -710 2868
rect -690 2774 -686 2868
rect -666 2774 -662 2868
rect -642 2774 -638 2868
rect -618 2774 -614 2868
rect -594 2774 -590 2868
rect -570 2774 -566 2868
rect -546 2774 -542 2868
rect -522 2774 -518 2868
rect -498 2774 -494 2868
rect -474 2774 -470 2868
rect -450 2774 -446 2868
rect -426 2774 -422 2868
rect -402 2774 -398 2868
rect -378 2774 -374 2868
rect -354 2774 -350 2868
rect -330 2774 -326 2868
rect -306 2774 -302 2868
rect -282 2774 -278 2868
rect -258 2774 -254 2868
rect -234 2774 -230 2868
rect -210 2774 -206 2868
rect -186 2774 -182 2868
rect -162 2774 -158 2868
rect -138 2774 -134 2868
rect -114 2774 -110 2868
rect -90 2774 -86 2868
rect -66 2774 -62 2868
rect -42 2774 -38 2868
rect -18 2774 -14 2868
rect 6 2774 10 2868
rect 30 2774 34 2868
rect 54 2774 58 2868
rect 78 2774 82 2868
rect 102 2774 106 2868
rect 126 2774 130 2868
rect 150 2774 154 2868
rect 174 2774 178 2868
rect 198 2774 202 2868
rect 222 2774 226 2868
rect 246 2774 250 2868
rect 270 2774 274 2868
rect 294 2774 298 2868
rect 318 2774 322 2868
rect 342 2774 346 2868
rect 366 2774 370 2868
rect 390 2774 394 2868
rect 414 2774 418 2868
rect 427 2837 432 2847
rect 438 2837 442 2868
rect 437 2823 442 2837
rect 427 2822 461 2823
rect 462 2822 466 2868
rect 486 2822 490 2868
rect 510 2822 514 2868
rect 534 2822 538 2868
rect 558 2822 562 2868
rect 582 2822 586 2868
rect 606 2822 610 2868
rect 630 2822 634 2868
rect 654 2822 658 2868
rect 678 2822 682 2868
rect 685 2867 699 2868
rect 702 2843 709 2891
rect 702 2822 706 2843
rect 726 2822 730 2916
rect 750 2822 754 2916
rect 774 2822 778 2916
rect 798 2822 802 2916
rect 822 2822 826 2916
rect 846 2822 850 2916
rect 870 2822 874 2916
rect 894 2822 898 2916
rect 918 2822 922 2916
rect 942 2822 946 2916
rect 966 2822 970 2916
rect 990 2822 994 2916
rect 1014 2822 1018 2916
rect 1038 2822 1042 2916
rect 1062 2822 1066 2916
rect 1086 2822 1090 2916
rect 1110 2822 1114 2916
rect 1134 2822 1138 2916
rect 1158 2822 1162 2916
rect 1182 2822 1186 2916
rect 1206 2822 1210 2916
rect 1230 2822 1234 2916
rect 1254 2822 1258 2916
rect 1278 2822 1282 2916
rect 1302 2822 1306 2916
rect 1326 2822 1330 2916
rect 1350 2822 1354 2916
rect 1374 2822 1378 2916
rect 1398 2822 1402 2916
rect 1422 2822 1426 2916
rect 1446 2822 1450 2916
rect 1470 2822 1474 2916
rect 1494 2822 1498 2916
rect 1518 2822 1522 2916
rect 1542 2822 1546 2916
rect 1566 2822 1570 2916
rect 1590 2822 1594 2916
rect 1614 2822 1618 2916
rect 1638 2822 1642 2916
rect 1662 2822 1666 2916
rect 1686 2822 1690 2916
rect 1710 2822 1714 2916
rect 1734 2822 1738 2916
rect 1758 2822 1762 2916
rect 1782 2822 1786 2916
rect 1806 2822 1810 2916
rect 1830 2822 1834 2916
rect 1854 2822 1858 2916
rect 1878 2822 1882 2916
rect 1902 2822 1906 2916
rect 1926 2822 1930 2916
rect 1939 2861 1944 2871
rect 1950 2861 1954 2916
rect 1949 2847 1954 2861
rect 1939 2846 1973 2847
rect 1974 2846 1978 2916
rect 1998 2846 2002 2916
rect 2022 2846 2026 2916
rect 2046 2846 2050 2916
rect 2070 2846 2074 2916
rect 2094 2846 2098 2916
rect 2118 2846 2122 2916
rect 2131 2909 2136 2916
rect 2149 2915 2163 2916
rect 2141 2895 2146 2909
rect 2142 2847 2146 2895
rect 2131 2846 2163 2847
rect 1939 2844 2163 2846
rect 1939 2837 1944 2844
rect 1949 2823 1954 2837
rect 1950 2822 1954 2823
rect 1974 2822 1978 2844
rect 1998 2822 2002 2844
rect 2022 2822 2026 2844
rect 2046 2822 2050 2844
rect 2070 2822 2074 2844
rect 2094 2822 2098 2844
rect 2118 2823 2122 2844
rect 2131 2837 2136 2844
rect 2142 2837 2146 2844
rect 2149 2843 2163 2844
rect 2141 2823 2146 2837
rect 2155 2833 2163 2837
rect 2149 2823 2155 2833
rect 2107 2822 2141 2823
rect 427 2820 2141 2822
rect 427 2813 432 2820
rect 437 2799 442 2813
rect 438 2774 442 2799
rect 462 2774 466 2820
rect 486 2774 490 2820
rect 510 2774 514 2820
rect 534 2774 538 2820
rect 558 2774 562 2820
rect 582 2774 586 2820
rect 606 2774 610 2820
rect 630 2774 634 2820
rect 654 2774 658 2820
rect 678 2774 682 2820
rect 702 2774 706 2820
rect 726 2774 730 2820
rect 750 2774 754 2820
rect 774 2774 778 2820
rect 798 2774 802 2820
rect 822 2774 826 2820
rect 846 2774 850 2820
rect 870 2774 874 2820
rect 894 2774 898 2820
rect 918 2774 922 2820
rect 942 2774 946 2820
rect 966 2774 970 2820
rect 990 2774 994 2820
rect 1014 2774 1018 2820
rect 1038 2774 1042 2820
rect 1062 2774 1066 2820
rect 1086 2774 1090 2820
rect 1110 2774 1114 2820
rect 1134 2774 1138 2820
rect 1158 2774 1162 2820
rect 1182 2774 1186 2820
rect 1206 2774 1210 2820
rect 1230 2774 1234 2820
rect 1254 2774 1258 2820
rect 1278 2774 1282 2820
rect 1302 2774 1306 2820
rect 1326 2774 1330 2820
rect 1350 2774 1354 2820
rect 1374 2774 1378 2820
rect 1398 2774 1402 2820
rect 1422 2774 1426 2820
rect 1446 2774 1450 2820
rect 1470 2774 1474 2820
rect 1494 2774 1498 2820
rect 1518 2774 1522 2820
rect 1542 2774 1546 2820
rect 1566 2774 1570 2820
rect 1590 2774 1594 2820
rect 1614 2774 1618 2820
rect 1638 2774 1642 2820
rect 1662 2774 1666 2820
rect 1686 2774 1690 2820
rect 1710 2774 1714 2820
rect 1734 2774 1738 2820
rect 1758 2774 1762 2820
rect 1782 2774 1786 2820
rect 1806 2774 1810 2820
rect 1830 2774 1834 2820
rect 1854 2774 1858 2820
rect 1878 2775 1882 2820
rect 1867 2774 1901 2775
rect -2393 2772 1901 2774
rect -2371 2750 -2366 2772
rect -2348 2750 -2343 2772
rect -2325 2762 -2317 2772
rect -2076 2762 -2068 2769
rect -2062 2762 -2001 2769
rect -2325 2750 -2320 2762
rect -2317 2758 -2309 2762
rect -2015 2761 -2001 2762
rect -2309 2750 -2301 2758
rect -2068 2752 -2062 2759
rect -2000 2754 -1992 2772
rect -1974 2770 -1960 2772
rect -1842 2771 -1804 2772
rect -1862 2769 -1794 2770
rect -1985 2767 -1794 2769
rect -1985 2762 -1852 2767
rect -1842 2761 -1794 2767
rect -1671 2762 -1663 2772
rect -2015 2752 -1985 2754
rect -1852 2752 -1804 2759
rect -1663 2758 -1655 2762
rect -2000 2750 -1992 2752
rect -1976 2750 -1940 2751
rect -1655 2750 -1647 2758
rect -1642 2750 -1637 2772
rect -1619 2750 -1614 2772
rect -1530 2750 -1526 2772
rect -1506 2750 -1502 2772
rect -1482 2750 -1478 2772
rect -1458 2750 -1454 2772
rect -1434 2750 -1430 2772
rect -1410 2750 -1406 2772
rect -1386 2750 -1382 2772
rect -1362 2750 -1358 2772
rect -1338 2750 -1334 2772
rect -1314 2750 -1310 2772
rect -1290 2750 -1286 2772
rect -1266 2750 -1262 2772
rect -1242 2750 -1238 2772
rect -1218 2750 -1214 2772
rect -1194 2750 -1190 2772
rect -1170 2750 -1166 2772
rect -1146 2750 -1142 2772
rect -1122 2750 -1118 2772
rect -1098 2750 -1094 2772
rect -1074 2750 -1070 2772
rect -1050 2750 -1046 2772
rect -1026 2750 -1022 2772
rect -1002 2750 -998 2772
rect -978 2750 -974 2772
rect -954 2750 -950 2772
rect -930 2750 -926 2772
rect -906 2750 -902 2772
rect -882 2750 -878 2772
rect -858 2750 -854 2772
rect -834 2750 -830 2772
rect -810 2750 -806 2772
rect -786 2750 -782 2772
rect -762 2750 -758 2772
rect -738 2750 -734 2772
rect -714 2750 -710 2772
rect -690 2750 -686 2772
rect -666 2750 -662 2772
rect -642 2750 -638 2772
rect -618 2750 -614 2772
rect -594 2750 -590 2772
rect -570 2750 -566 2772
rect -546 2750 -542 2772
rect -522 2750 -518 2772
rect -498 2750 -494 2772
rect -474 2750 -470 2772
rect -450 2750 -446 2772
rect -426 2750 -422 2772
rect -402 2750 -398 2772
rect -378 2750 -374 2772
rect -354 2750 -350 2772
rect -330 2750 -326 2772
rect -306 2750 -302 2772
rect -282 2750 -278 2772
rect -258 2750 -254 2772
rect -234 2750 -230 2772
rect -210 2750 -206 2772
rect -186 2750 -182 2772
rect -162 2750 -158 2772
rect -138 2750 -134 2772
rect -114 2750 -110 2772
rect -90 2750 -86 2772
rect -66 2750 -62 2772
rect -42 2750 -38 2772
rect -18 2750 -14 2772
rect 6 2750 10 2772
rect 30 2750 34 2772
rect 54 2751 58 2772
rect 43 2750 77 2751
rect -2393 2748 77 2750
rect -2371 2678 -2366 2748
rect -2348 2678 -2343 2748
rect -2325 2746 -2320 2748
rect -2309 2746 -2301 2748
rect -2325 2734 -2317 2746
rect -2062 2735 -2032 2742
rect -2325 2714 -2320 2734
rect -2317 2730 -2309 2734
rect -2325 2706 -2317 2714
rect -2060 2708 -2030 2711
rect -2325 2678 -2320 2706
rect -2317 2698 -2309 2706
rect -2060 2695 -2038 2706
rect -2033 2699 -2030 2708
rect -2028 2704 -2027 2708
rect -2068 2690 -2038 2693
rect -2000 2678 -1992 2748
rect -1888 2743 -1874 2748
rect -1842 2744 -1804 2748
rect -1655 2746 -1647 2748
rect -1902 2741 -1874 2743
rect -1842 2734 -1794 2743
rect -1671 2734 -1663 2746
rect -1663 2730 -1655 2734
rect -1912 2723 -1884 2725
rect -1852 2717 -1804 2721
rect -1844 2708 -1796 2711
rect -1671 2706 -1663 2714
rect -1844 2695 -1804 2706
rect -1663 2698 -1655 2706
rect -1852 2690 -1680 2694
rect -1642 2678 -1637 2748
rect -1619 2678 -1614 2748
rect -1530 2678 -1526 2748
rect -1506 2678 -1502 2748
rect -1482 2678 -1478 2748
rect -1458 2678 -1454 2748
rect -1434 2678 -1430 2748
rect -1410 2678 -1406 2748
rect -1386 2678 -1382 2748
rect -1362 2678 -1358 2748
rect -1338 2678 -1334 2748
rect -1314 2678 -1310 2748
rect -1290 2678 -1286 2748
rect -1277 2717 -1272 2727
rect -1266 2717 -1262 2748
rect -1267 2703 -1262 2717
rect -1277 2702 -1243 2703
rect -1242 2702 -1238 2748
rect -1218 2702 -1214 2748
rect -1194 2702 -1190 2748
rect -1170 2702 -1166 2748
rect -1146 2702 -1142 2748
rect -1122 2702 -1118 2748
rect -1098 2702 -1094 2748
rect -1074 2702 -1070 2748
rect -1050 2702 -1046 2748
rect -1026 2702 -1022 2748
rect -1002 2702 -998 2748
rect -978 2702 -974 2748
rect -954 2702 -950 2748
rect -930 2702 -926 2748
rect -906 2702 -902 2748
rect -882 2702 -878 2748
rect -858 2702 -854 2748
rect -834 2702 -830 2748
rect -810 2702 -806 2748
rect -786 2702 -782 2748
rect -762 2702 -758 2748
rect -738 2702 -734 2748
rect -714 2702 -710 2748
rect -690 2702 -686 2748
rect -666 2702 -662 2748
rect -642 2702 -638 2748
rect -618 2702 -614 2748
rect -594 2702 -590 2748
rect -570 2702 -566 2748
rect -546 2702 -542 2748
rect -522 2702 -518 2748
rect -498 2702 -494 2748
rect -474 2702 -470 2748
rect -450 2702 -446 2748
rect -426 2702 -422 2748
rect -402 2702 -398 2748
rect -378 2702 -374 2748
rect -354 2702 -350 2748
rect -330 2702 -326 2748
rect -306 2702 -302 2748
rect -282 2702 -278 2748
rect -258 2702 -254 2748
rect -234 2702 -230 2748
rect -210 2702 -206 2748
rect -186 2702 -182 2748
rect -162 2702 -158 2748
rect -138 2702 -134 2748
rect -114 2702 -110 2748
rect -90 2702 -86 2748
rect -66 2702 -62 2748
rect -42 2702 -38 2748
rect -18 2702 -14 2748
rect 6 2702 10 2748
rect 30 2702 34 2748
rect 43 2741 48 2748
rect 54 2741 58 2748
rect 53 2727 58 2741
rect 43 2717 48 2727
rect 53 2703 58 2717
rect 54 2702 58 2703
rect 78 2702 82 2772
rect 102 2702 106 2772
rect 126 2702 130 2772
rect 150 2702 154 2772
rect 174 2702 178 2772
rect 198 2702 202 2772
rect 222 2702 226 2772
rect 246 2702 250 2772
rect 270 2702 274 2772
rect 294 2702 298 2772
rect 318 2702 322 2772
rect 342 2702 346 2772
rect 366 2702 370 2772
rect 390 2702 394 2772
rect 414 2702 418 2772
rect 438 2702 442 2772
rect 462 2771 466 2772
rect 462 2726 469 2771
rect 486 2726 490 2772
rect 510 2726 514 2772
rect 534 2726 538 2772
rect 558 2726 562 2772
rect 582 2726 586 2772
rect 606 2726 610 2772
rect 630 2726 634 2772
rect 654 2726 658 2772
rect 678 2726 682 2772
rect 702 2726 706 2772
rect 726 2726 730 2772
rect 750 2726 754 2772
rect 774 2726 778 2772
rect 798 2726 802 2772
rect 822 2726 826 2772
rect 846 2726 850 2772
rect 870 2726 874 2772
rect 894 2726 898 2772
rect 918 2726 922 2772
rect 942 2726 946 2772
rect 966 2726 970 2772
rect 990 2726 994 2772
rect 1014 2726 1018 2772
rect 1038 2726 1042 2772
rect 1062 2726 1066 2772
rect 1086 2726 1090 2772
rect 1110 2726 1114 2772
rect 1134 2726 1138 2772
rect 1158 2726 1162 2772
rect 1182 2726 1186 2772
rect 1206 2726 1210 2772
rect 1230 2726 1234 2772
rect 1254 2726 1258 2772
rect 1278 2726 1282 2772
rect 1302 2726 1306 2772
rect 1326 2726 1330 2772
rect 1350 2726 1354 2772
rect 1374 2726 1378 2772
rect 1398 2726 1402 2772
rect 1422 2726 1426 2772
rect 1446 2726 1450 2772
rect 1470 2726 1474 2772
rect 1494 2726 1498 2772
rect 1518 2726 1522 2772
rect 1542 2726 1546 2772
rect 1566 2726 1570 2772
rect 1590 2726 1594 2772
rect 1614 2726 1618 2772
rect 1638 2726 1642 2772
rect 1662 2726 1666 2772
rect 1686 2726 1690 2772
rect 1710 2726 1714 2772
rect 1734 2726 1738 2772
rect 1758 2726 1762 2772
rect 1782 2726 1786 2772
rect 1806 2726 1810 2772
rect 1830 2726 1834 2772
rect 1854 2726 1858 2772
rect 1867 2765 1872 2772
rect 1878 2765 1882 2772
rect 1877 2751 1882 2765
rect 1867 2741 1872 2751
rect 1877 2727 1882 2741
rect 1878 2726 1882 2727
rect 1902 2726 1906 2820
rect 1926 2726 1930 2820
rect 1950 2726 1954 2820
rect 1974 2795 1978 2820
rect 1974 2750 1981 2795
rect 1998 2750 2002 2820
rect 2022 2750 2026 2820
rect 2046 2750 2050 2820
rect 2070 2750 2074 2820
rect 2094 2750 2098 2820
rect 2107 2813 2112 2820
rect 2118 2813 2122 2820
rect 2117 2799 2122 2813
rect 2107 2789 2112 2799
rect 2117 2775 2122 2789
rect 2118 2751 2122 2775
rect 2107 2750 2141 2751
rect 1957 2748 2141 2750
rect 1957 2747 1971 2748
rect 1974 2747 1981 2748
rect 1974 2726 1978 2747
rect 1998 2726 2002 2748
rect 2022 2726 2026 2748
rect 2046 2726 2050 2748
rect 2070 2726 2074 2748
rect 2094 2727 2098 2748
rect 2107 2741 2112 2748
rect 2118 2741 2122 2748
rect 2117 2727 2122 2741
rect 2131 2737 2139 2741
rect 2125 2727 2131 2737
rect 2083 2726 2117 2727
rect 445 2724 2117 2726
rect 445 2723 459 2724
rect 462 2723 469 2724
rect 462 2702 466 2723
rect 486 2702 490 2724
rect 510 2702 514 2724
rect 534 2702 538 2724
rect 558 2702 562 2724
rect 582 2702 586 2724
rect 606 2702 610 2724
rect 630 2702 634 2724
rect 654 2702 658 2724
rect 678 2702 682 2724
rect 702 2702 706 2724
rect 726 2702 730 2724
rect 750 2702 754 2724
rect 774 2702 778 2724
rect 798 2702 802 2724
rect 822 2702 826 2724
rect 846 2702 850 2724
rect 870 2702 874 2724
rect 894 2702 898 2724
rect 918 2702 922 2724
rect 942 2702 946 2724
rect 966 2702 970 2724
rect 990 2702 994 2724
rect 1014 2702 1018 2724
rect 1038 2702 1042 2724
rect 1062 2702 1066 2724
rect 1086 2702 1090 2724
rect 1110 2702 1114 2724
rect 1134 2702 1138 2724
rect 1158 2702 1162 2724
rect 1182 2702 1186 2724
rect 1206 2702 1210 2724
rect 1230 2702 1234 2724
rect 1254 2702 1258 2724
rect 1278 2702 1282 2724
rect 1302 2702 1306 2724
rect 1326 2702 1330 2724
rect 1350 2702 1354 2724
rect 1374 2702 1378 2724
rect 1398 2702 1402 2724
rect 1422 2702 1426 2724
rect 1446 2702 1450 2724
rect 1470 2702 1474 2724
rect 1494 2702 1498 2724
rect 1518 2702 1522 2724
rect 1542 2702 1546 2724
rect 1566 2702 1570 2724
rect 1590 2702 1594 2724
rect 1614 2702 1618 2724
rect 1638 2702 1642 2724
rect 1662 2702 1666 2724
rect 1686 2702 1690 2724
rect 1710 2702 1714 2724
rect 1734 2702 1738 2724
rect 1758 2702 1762 2724
rect 1782 2702 1786 2724
rect 1806 2702 1810 2724
rect 1830 2702 1834 2724
rect 1854 2702 1858 2724
rect 1878 2702 1882 2724
rect 1902 2702 1906 2724
rect 1926 2702 1930 2724
rect 1950 2702 1954 2724
rect 1974 2702 1978 2724
rect 1998 2702 2002 2724
rect 2022 2702 2026 2724
rect 2046 2702 2050 2724
rect 2070 2703 2074 2724
rect 2083 2717 2088 2724
rect 2094 2717 2098 2724
rect 2093 2703 2098 2717
rect 2059 2702 2093 2703
rect -1277 2700 2093 2702
rect -1277 2693 -1272 2700
rect -1267 2679 -1262 2693
rect -1266 2678 -1262 2679
rect -1242 2678 -1238 2700
rect -1218 2678 -1214 2700
rect -1194 2678 -1190 2700
rect -1170 2678 -1166 2700
rect -1146 2678 -1142 2700
rect -1122 2678 -1118 2700
rect -1098 2678 -1094 2700
rect -1074 2678 -1070 2700
rect -1050 2678 -1046 2700
rect -1026 2678 -1022 2700
rect -1002 2678 -998 2700
rect -978 2678 -974 2700
rect -954 2678 -950 2700
rect -930 2678 -926 2700
rect -906 2678 -902 2700
rect -882 2678 -878 2700
rect -858 2678 -854 2700
rect -834 2678 -830 2700
rect -810 2678 -806 2700
rect -786 2678 -782 2700
rect -762 2678 -758 2700
rect -738 2678 -734 2700
rect -714 2678 -710 2700
rect -690 2678 -686 2700
rect -666 2678 -662 2700
rect -642 2678 -638 2700
rect -618 2678 -614 2700
rect -594 2678 -590 2700
rect -570 2678 -566 2700
rect -546 2678 -542 2700
rect -522 2678 -518 2700
rect -498 2678 -494 2700
rect -474 2678 -470 2700
rect -450 2678 -446 2700
rect -426 2678 -422 2700
rect -402 2678 -398 2700
rect -378 2678 -374 2700
rect -354 2678 -350 2700
rect -330 2678 -326 2700
rect -306 2678 -302 2700
rect -282 2678 -278 2700
rect -258 2678 -254 2700
rect -234 2678 -230 2700
rect -210 2678 -206 2700
rect -186 2678 -182 2700
rect -162 2678 -158 2700
rect -138 2678 -134 2700
rect -114 2678 -110 2700
rect -90 2678 -86 2700
rect -66 2678 -62 2700
rect -42 2678 -38 2700
rect -18 2678 -14 2700
rect 6 2678 10 2700
rect 30 2678 34 2700
rect 54 2678 58 2700
rect 78 2678 82 2700
rect 102 2678 106 2700
rect 126 2678 130 2700
rect 150 2678 154 2700
rect 174 2678 178 2700
rect 198 2678 202 2700
rect 222 2678 226 2700
rect 246 2678 250 2700
rect 270 2678 274 2700
rect 294 2678 298 2700
rect 318 2678 322 2700
rect 342 2678 346 2700
rect 366 2678 370 2700
rect 390 2678 394 2700
rect 414 2678 418 2700
rect 438 2678 442 2700
rect 462 2678 466 2700
rect 486 2678 490 2700
rect 510 2678 514 2700
rect 534 2678 538 2700
rect 558 2678 562 2700
rect 582 2678 586 2700
rect 606 2678 610 2700
rect 630 2678 634 2700
rect 654 2678 658 2700
rect 678 2678 682 2700
rect 702 2678 706 2700
rect 726 2678 730 2700
rect 750 2678 754 2700
rect 774 2678 778 2700
rect 798 2678 802 2700
rect 822 2678 826 2700
rect 846 2678 850 2700
rect 870 2678 874 2700
rect 894 2678 898 2700
rect 918 2678 922 2700
rect 942 2678 946 2700
rect 966 2678 970 2700
rect 990 2678 994 2700
rect 1014 2678 1018 2700
rect 1038 2678 1042 2700
rect 1062 2678 1066 2700
rect 1086 2678 1090 2700
rect 1110 2678 1114 2700
rect 1134 2678 1138 2700
rect 1158 2678 1162 2700
rect 1182 2678 1186 2700
rect 1206 2678 1210 2700
rect 1230 2678 1234 2700
rect 1254 2678 1258 2700
rect 1278 2678 1282 2700
rect 1302 2678 1306 2700
rect 1326 2678 1330 2700
rect 1350 2678 1354 2700
rect 1374 2678 1378 2700
rect 1398 2678 1402 2700
rect 1422 2678 1426 2700
rect 1446 2678 1450 2700
rect 1470 2678 1474 2700
rect 1494 2678 1498 2700
rect 1518 2678 1522 2700
rect 1542 2678 1546 2700
rect 1566 2678 1570 2700
rect 1590 2679 1594 2700
rect 1579 2678 1613 2679
rect -2393 2676 1613 2678
rect -2371 2654 -2366 2676
rect -2348 2654 -2343 2676
rect -2325 2654 -2320 2676
rect -2309 2658 -2301 2668
rect -2068 2659 -2062 2664
rect -2317 2654 -2309 2658
rect -2060 2654 -2050 2659
rect -2000 2654 -1992 2676
rect -1806 2668 -1680 2674
rect -1854 2659 -1806 2664
rect -1655 2658 -1647 2668
rect -1972 2654 -1964 2655
rect -1958 2654 -1942 2656
rect -1844 2654 -1806 2657
rect -1663 2654 -1655 2658
rect -1642 2654 -1637 2676
rect -1619 2654 -1614 2676
rect -1530 2654 -1526 2676
rect -1506 2654 -1502 2676
rect -1482 2654 -1478 2676
rect -1458 2654 -1454 2676
rect -1434 2654 -1430 2676
rect -1410 2654 -1406 2676
rect -1386 2654 -1382 2676
rect -1362 2654 -1358 2676
rect -1338 2654 -1334 2676
rect -1314 2654 -1310 2676
rect -1290 2654 -1286 2676
rect -1266 2654 -1262 2676
rect -1242 2654 -1238 2676
rect -1218 2654 -1214 2676
rect -1194 2654 -1190 2676
rect -1170 2654 -1166 2676
rect -1146 2654 -1142 2676
rect -1122 2654 -1118 2676
rect -1098 2654 -1094 2676
rect -1074 2654 -1070 2676
rect -1050 2654 -1046 2676
rect -1026 2654 -1022 2676
rect -1002 2654 -998 2676
rect -978 2654 -974 2676
rect -954 2654 -950 2676
rect -930 2654 -926 2676
rect -906 2654 -902 2676
rect -882 2654 -878 2676
rect -858 2654 -854 2676
rect -834 2654 -830 2676
rect -810 2654 -806 2676
rect -786 2654 -782 2676
rect -762 2654 -758 2676
rect -738 2654 -734 2676
rect -714 2654 -710 2676
rect -690 2654 -686 2676
rect -666 2654 -662 2676
rect -642 2654 -638 2676
rect -618 2654 -614 2676
rect -594 2654 -590 2676
rect -570 2654 -566 2676
rect -546 2654 -542 2676
rect -522 2654 -518 2676
rect -498 2654 -494 2676
rect -474 2654 -470 2676
rect -450 2654 -446 2676
rect -426 2654 -422 2676
rect -402 2654 -398 2676
rect -378 2654 -374 2676
rect -354 2654 -350 2676
rect -330 2654 -326 2676
rect -306 2654 -302 2676
rect -282 2654 -278 2676
rect -258 2654 -254 2676
rect -234 2654 -230 2676
rect -210 2654 -206 2676
rect -186 2654 -182 2676
rect -162 2654 -158 2676
rect -138 2654 -134 2676
rect -114 2654 -110 2676
rect -90 2654 -86 2676
rect -66 2654 -62 2676
rect -42 2654 -38 2676
rect -18 2654 -14 2676
rect 6 2654 10 2676
rect 30 2654 34 2676
rect 54 2654 58 2676
rect 78 2675 82 2676
rect -2393 2652 75 2654
rect -2371 2630 -2366 2652
rect -2348 2630 -2343 2652
rect -2325 2630 -2320 2652
rect -2060 2646 -2050 2652
rect -2309 2630 -2301 2640
rect -2060 2639 -2030 2646
rect -2000 2642 -1992 2652
rect -1972 2650 -1942 2652
rect -1958 2649 -1942 2650
rect -1844 2648 -1806 2652
rect -2068 2632 -2062 2639
rect -2062 2630 -2036 2632
rect -2393 2628 -2036 2630
rect -2030 2630 -2012 2632
rect -2004 2630 -1990 2642
rect -1844 2641 -1798 2646
rect -1806 2639 -1798 2641
rect -1854 2637 -1844 2639
rect -1854 2632 -1806 2637
rect -1864 2630 -1796 2631
rect -1655 2630 -1647 2640
rect -1642 2630 -1637 2652
rect -1619 2630 -1614 2652
rect -1530 2630 -1526 2652
rect -1506 2630 -1502 2652
rect -1482 2630 -1478 2652
rect -1458 2630 -1454 2652
rect -1434 2630 -1430 2652
rect -1410 2630 -1406 2652
rect -1386 2630 -1382 2652
rect -1362 2630 -1358 2652
rect -1338 2631 -1334 2652
rect -1349 2630 -1315 2631
rect -2030 2628 -1315 2630
rect -2371 2558 -2366 2628
rect -2348 2558 -2343 2628
rect -2325 2558 -2320 2628
rect -2317 2624 -2309 2628
rect -2060 2624 -2050 2628
rect -2060 2622 -2036 2624
rect -2060 2620 -2030 2622
rect -2292 2614 -2030 2620
rect -2092 2598 -2062 2600
rect -2094 2594 -2062 2598
rect -2309 2564 -2301 2570
rect -2317 2558 -2309 2564
rect -2000 2558 -1992 2628
rect -1844 2621 -1806 2628
rect -1663 2624 -1655 2628
rect -1844 2614 -1680 2620
rect -1854 2598 -1806 2600
rect -1854 2594 -1680 2598
rect -1655 2564 -1647 2570
rect -1663 2558 -1655 2564
rect -1642 2558 -1637 2628
rect -1619 2558 -1614 2628
rect -1530 2558 -1526 2628
rect -1506 2558 -1502 2628
rect -1482 2558 -1478 2628
rect -1458 2558 -1454 2628
rect -1434 2558 -1430 2628
rect -1410 2558 -1406 2628
rect -1386 2558 -1382 2628
rect -1362 2558 -1358 2628
rect -1349 2621 -1344 2628
rect -1338 2621 -1334 2628
rect -1339 2607 -1334 2621
rect -1338 2558 -1334 2607
rect -1314 2558 -1310 2652
rect -1290 2558 -1286 2652
rect -1266 2558 -1262 2652
rect -1242 2651 -1238 2652
rect -1242 2603 -1235 2651
rect -1242 2558 -1238 2603
rect -1218 2558 -1214 2652
rect -1194 2558 -1190 2652
rect -1170 2558 -1166 2652
rect -1146 2558 -1142 2652
rect -1122 2558 -1118 2652
rect -1098 2558 -1094 2652
rect -1074 2558 -1070 2652
rect -1050 2558 -1046 2652
rect -1026 2558 -1022 2652
rect -1002 2558 -998 2652
rect -978 2558 -974 2652
rect -954 2558 -950 2652
rect -930 2558 -926 2652
rect -906 2558 -902 2652
rect -882 2558 -878 2652
rect -858 2558 -854 2652
rect -834 2558 -830 2652
rect -810 2558 -806 2652
rect -786 2558 -782 2652
rect -762 2558 -758 2652
rect -738 2558 -734 2652
rect -714 2558 -710 2652
rect -690 2558 -686 2652
rect -666 2558 -662 2652
rect -642 2558 -638 2652
rect -618 2558 -614 2652
rect -594 2558 -590 2652
rect -570 2558 -566 2652
rect -546 2558 -542 2652
rect -522 2558 -518 2652
rect -498 2558 -494 2652
rect -474 2558 -470 2652
rect -450 2558 -446 2652
rect -426 2558 -422 2652
rect -402 2558 -398 2652
rect -378 2558 -374 2652
rect -354 2558 -350 2652
rect -330 2558 -326 2652
rect -306 2558 -302 2652
rect -282 2558 -278 2652
rect -258 2558 -254 2652
rect -234 2558 -230 2652
rect -210 2558 -206 2652
rect -186 2558 -182 2652
rect -162 2558 -158 2652
rect -138 2559 -134 2652
rect -149 2558 -115 2559
rect -2393 2556 -115 2558
rect -2371 2462 -2366 2556
rect -2348 2462 -2343 2556
rect -2325 2494 -2320 2556
rect -2317 2554 -2309 2556
rect -2000 2555 -1966 2556
rect -2000 2554 -1982 2555
rect -1663 2554 -1655 2556
rect -2028 2546 -2018 2548
rect -2309 2536 -2301 2542
rect -2091 2536 -2061 2543
rect -2317 2526 -2309 2536
rect -2044 2534 -2028 2536
rect -2026 2534 -2014 2546
rect -2084 2528 -2061 2534
rect -2044 2532 -2014 2534
rect -2292 2518 -2054 2527
rect -2325 2486 -2317 2494
rect -2325 2466 -2320 2486
rect -2317 2478 -2309 2486
rect -2325 2462 -2317 2466
rect -2000 2462 -1992 2554
rect -1982 2553 -1966 2554
rect -1980 2536 -1932 2543
rect -1655 2536 -1647 2542
rect -1846 2518 -1680 2527
rect -1663 2526 -1655 2536
rect -1671 2486 -1663 2494
rect -1663 2478 -1655 2486
rect -1671 2462 -1663 2466
rect -1642 2462 -1637 2556
rect -1619 2462 -1614 2556
rect -1530 2462 -1526 2556
rect -1506 2462 -1502 2556
rect -1482 2462 -1478 2556
rect -1458 2462 -1454 2556
rect -1434 2462 -1430 2556
rect -1410 2462 -1406 2556
rect -1386 2462 -1382 2556
rect -1362 2462 -1358 2556
rect -1338 2462 -1334 2556
rect -1314 2555 -1310 2556
rect -1314 2531 -1307 2555
rect -1314 2462 -1310 2531
rect -1290 2462 -1286 2556
rect -1266 2462 -1262 2556
rect -1242 2462 -1238 2556
rect -1218 2462 -1214 2556
rect -1194 2462 -1190 2556
rect -1170 2462 -1166 2556
rect -1146 2462 -1142 2556
rect -1122 2462 -1118 2556
rect -1098 2462 -1094 2556
rect -1074 2462 -1070 2556
rect -1050 2462 -1046 2556
rect -1026 2462 -1022 2556
rect -1002 2462 -998 2556
rect -978 2462 -974 2556
rect -954 2462 -950 2556
rect -930 2462 -926 2556
rect -906 2462 -902 2556
rect -893 2501 -888 2511
rect -882 2501 -878 2556
rect -883 2487 -878 2501
rect -882 2462 -878 2487
rect -858 2462 -854 2556
rect -834 2462 -830 2556
rect -810 2462 -806 2556
rect -786 2462 -782 2556
rect -762 2462 -758 2556
rect -738 2462 -734 2556
rect -714 2462 -710 2556
rect -690 2462 -686 2556
rect -666 2462 -662 2556
rect -642 2462 -638 2556
rect -618 2462 -614 2556
rect -594 2462 -590 2556
rect -570 2462 -566 2556
rect -546 2462 -542 2556
rect -522 2462 -518 2556
rect -498 2462 -494 2556
rect -474 2462 -470 2556
rect -450 2462 -446 2556
rect -426 2462 -422 2556
rect -402 2462 -398 2556
rect -378 2462 -374 2556
rect -354 2462 -350 2556
rect -330 2462 -326 2556
rect -306 2462 -302 2556
rect -282 2462 -278 2556
rect -258 2462 -254 2556
rect -234 2462 -230 2556
rect -210 2462 -206 2556
rect -186 2462 -182 2556
rect -162 2462 -158 2556
rect -149 2549 -144 2556
rect -138 2549 -134 2556
rect -139 2535 -134 2549
rect -149 2525 -144 2535
rect -139 2511 -134 2525
rect -138 2462 -134 2511
rect -114 2483 -110 2652
rect -2393 2460 -117 2462
rect -2371 2414 -2366 2460
rect -2348 2414 -2343 2460
rect -2325 2452 -2317 2460
rect -2018 2459 -2004 2460
rect -2000 2459 -1992 2460
rect -2072 2458 -1928 2459
rect -2072 2452 -2053 2458
rect -2325 2436 -2320 2452
rect -2317 2450 -2309 2452
rect -2309 2438 -2301 2450
rect -2092 2443 -2062 2448
rect -2317 2436 -2309 2438
rect -2325 2424 -2317 2436
rect -2098 2430 -2096 2441
rect -2092 2430 -2084 2443
rect -2000 2442 -1992 2458
rect -1972 2452 -1928 2458
rect -1924 2452 -1918 2460
rect -1671 2452 -1663 2460
rect -1663 2450 -1655 2452
rect -2083 2432 -2062 2441
rect -2027 2440 -1992 2442
rect -2018 2432 -2002 2440
rect -2000 2432 -1992 2440
rect -2100 2425 -2096 2430
rect -2083 2425 -2053 2430
rect -2003 2428 -1990 2432
rect -1972 2430 -1964 2439
rect -1928 2438 -1924 2441
rect -1655 2438 -1647 2450
rect -1663 2436 -1655 2438
rect -2325 2414 -2320 2424
rect -2317 2422 -2309 2424
rect -2309 2414 -2301 2422
rect -2004 2418 -2003 2428
rect -2062 2414 -2012 2416
rect -2000 2414 -1992 2428
rect -1972 2425 -1924 2430
rect -1864 2425 -1796 2431
rect -1671 2424 -1663 2436
rect -1663 2422 -1655 2424
rect -1864 2414 -1796 2415
rect -1655 2414 -1647 2422
rect -1642 2414 -1637 2460
rect -1619 2414 -1614 2460
rect -1530 2414 -1526 2460
rect -1506 2414 -1502 2460
rect -1482 2414 -1478 2460
rect -1458 2414 -1454 2460
rect -1434 2414 -1430 2460
rect -1410 2414 -1406 2460
rect -1386 2414 -1382 2460
rect -1362 2414 -1358 2460
rect -1338 2414 -1334 2460
rect -1314 2414 -1310 2460
rect -1290 2414 -1286 2460
rect -1266 2414 -1262 2460
rect -1242 2414 -1238 2460
rect -1218 2414 -1214 2460
rect -1194 2414 -1190 2460
rect -1170 2414 -1166 2460
rect -1146 2414 -1142 2460
rect -1122 2414 -1118 2460
rect -1098 2414 -1094 2460
rect -1074 2414 -1070 2460
rect -1050 2414 -1046 2460
rect -1026 2414 -1022 2460
rect -1002 2414 -998 2460
rect -978 2414 -974 2460
rect -954 2414 -950 2460
rect -930 2414 -926 2460
rect -906 2414 -902 2460
rect -882 2414 -878 2460
rect -858 2435 -854 2460
rect -2393 2412 -861 2414
rect -2371 2366 -2366 2412
rect -2348 2366 -2343 2412
rect -2325 2408 -2320 2412
rect -2309 2410 -2301 2412
rect -2317 2408 -2309 2410
rect -2325 2396 -2317 2408
rect -2325 2366 -2320 2396
rect -2317 2394 -2309 2396
rect -2092 2382 -2062 2384
rect -2094 2378 -2062 2382
rect -2000 2366 -1992 2412
rect -1655 2410 -1647 2412
rect -1663 2408 -1655 2410
rect -1671 2396 -1663 2408
rect -1663 2394 -1655 2396
rect -1854 2382 -1806 2384
rect -1854 2378 -1680 2382
rect -1979 2366 -1945 2368
rect -1642 2366 -1637 2412
rect -1619 2366 -1614 2412
rect -1530 2366 -1526 2412
rect -1506 2366 -1502 2412
rect -1482 2366 -1478 2412
rect -1458 2366 -1454 2412
rect -1434 2366 -1430 2412
rect -1410 2366 -1406 2412
rect -1386 2366 -1382 2412
rect -1362 2366 -1358 2412
rect -1338 2366 -1334 2412
rect -1314 2366 -1310 2412
rect -1290 2366 -1286 2412
rect -1266 2366 -1262 2412
rect -1242 2366 -1238 2412
rect -1218 2366 -1214 2412
rect -1194 2366 -1190 2412
rect -1170 2366 -1166 2412
rect -1146 2366 -1142 2412
rect -1122 2366 -1118 2412
rect -1098 2366 -1094 2412
rect -1074 2366 -1070 2412
rect -1050 2366 -1046 2412
rect -1026 2366 -1022 2412
rect -1002 2366 -998 2412
rect -978 2366 -974 2412
rect -954 2366 -950 2412
rect -930 2366 -926 2412
rect -906 2366 -902 2412
rect -882 2366 -878 2412
rect -875 2411 -861 2412
rect -858 2411 -851 2435
rect -858 2366 -854 2411
rect -834 2366 -830 2460
rect -810 2366 -806 2460
rect -786 2366 -782 2460
rect -762 2366 -758 2460
rect -738 2366 -734 2460
rect -725 2429 -720 2439
rect -714 2429 -710 2460
rect -715 2415 -710 2429
rect -714 2366 -710 2415
rect -690 2366 -686 2460
rect -666 2366 -662 2460
rect -642 2366 -638 2460
rect -618 2366 -614 2460
rect -594 2366 -590 2460
rect -570 2366 -566 2460
rect -546 2366 -542 2460
rect -522 2366 -518 2460
rect -498 2366 -494 2460
rect -474 2366 -470 2460
rect -450 2366 -446 2460
rect -426 2366 -422 2460
rect -402 2366 -398 2460
rect -378 2366 -374 2460
rect -354 2366 -350 2460
rect -330 2366 -326 2460
rect -306 2366 -302 2460
rect -282 2366 -278 2460
rect -258 2366 -254 2460
rect -234 2366 -230 2460
rect -210 2366 -206 2460
rect -186 2366 -182 2460
rect -162 2366 -158 2460
rect -138 2366 -134 2460
rect -131 2459 -117 2460
rect -114 2435 -107 2483
rect -114 2366 -110 2435
rect -90 2366 -86 2652
rect -66 2366 -62 2652
rect -42 2366 -38 2652
rect -18 2366 -14 2652
rect 6 2366 10 2652
rect 30 2366 34 2652
rect 54 2366 58 2652
rect 61 2651 75 2652
rect 78 2627 85 2675
rect 78 2366 82 2627
rect 102 2366 106 2676
rect 126 2366 130 2676
rect 150 2366 154 2676
rect 174 2366 178 2676
rect 198 2366 202 2676
rect 222 2366 226 2676
rect 246 2366 250 2676
rect 270 2366 274 2676
rect 294 2366 298 2676
rect 318 2366 322 2676
rect 342 2366 346 2676
rect 366 2366 370 2676
rect 390 2366 394 2676
rect 414 2366 418 2676
rect 438 2366 442 2676
rect 462 2366 466 2676
rect 486 2366 490 2676
rect 510 2366 514 2676
rect 534 2366 538 2676
rect 558 2366 562 2676
rect 582 2366 586 2676
rect 606 2366 610 2676
rect 630 2366 634 2676
rect 654 2366 658 2676
rect 678 2366 682 2676
rect 702 2366 706 2676
rect 726 2366 730 2676
rect 750 2366 754 2676
rect 774 2366 778 2676
rect 798 2366 802 2676
rect 822 2366 826 2676
rect 846 2366 850 2676
rect 870 2366 874 2676
rect 894 2366 898 2676
rect 918 2366 922 2676
rect 942 2366 946 2676
rect 966 2366 970 2676
rect 990 2366 994 2676
rect 1014 2366 1018 2676
rect 1038 2366 1042 2676
rect 1051 2645 1056 2655
rect 1062 2645 1066 2676
rect 1061 2631 1066 2645
rect 1051 2630 1085 2631
rect 1086 2630 1090 2676
rect 1110 2630 1114 2676
rect 1134 2630 1138 2676
rect 1158 2630 1162 2676
rect 1182 2630 1186 2676
rect 1206 2630 1210 2676
rect 1230 2630 1234 2676
rect 1254 2630 1258 2676
rect 1278 2630 1282 2676
rect 1302 2630 1306 2676
rect 1326 2630 1330 2676
rect 1350 2630 1354 2676
rect 1374 2630 1378 2676
rect 1398 2630 1402 2676
rect 1422 2630 1426 2676
rect 1446 2630 1450 2676
rect 1470 2630 1474 2676
rect 1494 2630 1498 2676
rect 1518 2630 1522 2676
rect 1542 2630 1546 2676
rect 1566 2630 1570 2676
rect 1579 2669 1584 2676
rect 1590 2669 1594 2676
rect 1589 2655 1594 2669
rect 1579 2645 1584 2655
rect 1589 2631 1594 2645
rect 1590 2630 1594 2631
rect 1614 2630 1618 2700
rect 1638 2630 1642 2700
rect 1662 2630 1666 2700
rect 1686 2630 1690 2700
rect 1710 2630 1714 2700
rect 1734 2630 1738 2700
rect 1758 2630 1762 2700
rect 1782 2630 1786 2700
rect 1806 2630 1810 2700
rect 1830 2630 1834 2700
rect 1854 2630 1858 2700
rect 1878 2630 1882 2700
rect 1902 2699 1906 2700
rect 1902 2654 1909 2699
rect 1926 2654 1930 2700
rect 1950 2654 1954 2700
rect 1974 2654 1978 2700
rect 1998 2654 2002 2700
rect 2022 2654 2026 2700
rect 2046 2655 2050 2700
rect 2059 2693 2064 2700
rect 2070 2693 2074 2700
rect 2069 2679 2074 2693
rect 2035 2654 2069 2655
rect 1885 2652 2069 2654
rect 1885 2651 1899 2652
rect 1902 2651 1909 2652
rect 1902 2630 1906 2651
rect 1926 2630 1930 2652
rect 1950 2630 1954 2652
rect 1974 2630 1978 2652
rect 1998 2630 2002 2652
rect 2022 2631 2026 2652
rect 2035 2645 2040 2652
rect 2046 2645 2050 2652
rect 2045 2631 2050 2645
rect 2011 2630 2045 2631
rect 1051 2628 2045 2630
rect 1051 2621 1056 2628
rect 1061 2607 1066 2621
rect 1062 2366 1066 2607
rect 1086 2579 1090 2628
rect 1086 2534 1093 2579
rect 1110 2534 1114 2628
rect 1134 2534 1138 2628
rect 1158 2534 1162 2628
rect 1182 2534 1186 2628
rect 1206 2534 1210 2628
rect 1230 2534 1234 2628
rect 1254 2534 1258 2628
rect 1278 2534 1282 2628
rect 1302 2534 1306 2628
rect 1326 2534 1330 2628
rect 1350 2534 1354 2628
rect 1374 2534 1378 2628
rect 1398 2534 1402 2628
rect 1422 2534 1426 2628
rect 1446 2534 1450 2628
rect 1470 2534 1474 2628
rect 1494 2534 1498 2628
rect 1518 2534 1522 2628
rect 1542 2534 1546 2628
rect 1566 2534 1570 2628
rect 1590 2534 1594 2628
rect 1614 2603 1618 2628
rect 1614 2555 1621 2603
rect 1614 2534 1618 2555
rect 1638 2534 1642 2628
rect 1662 2534 1666 2628
rect 1686 2534 1690 2628
rect 1710 2534 1714 2628
rect 1734 2534 1738 2628
rect 1758 2534 1762 2628
rect 1782 2534 1786 2628
rect 1806 2534 1810 2628
rect 1830 2534 1834 2628
rect 1854 2534 1858 2628
rect 1878 2534 1882 2628
rect 1902 2534 1906 2628
rect 1926 2534 1930 2628
rect 1950 2534 1954 2628
rect 1974 2534 1978 2628
rect 1998 2535 2002 2628
rect 2011 2621 2016 2628
rect 2022 2621 2026 2628
rect 2021 2607 2026 2621
rect 1987 2534 2021 2535
rect 1069 2532 2021 2534
rect 1069 2531 1083 2532
rect 1086 2531 1093 2532
rect 1086 2366 1090 2531
rect 1110 2366 1114 2532
rect 1134 2366 1138 2532
rect 1158 2366 1162 2532
rect 1182 2366 1186 2532
rect 1206 2366 1210 2532
rect 1230 2366 1234 2532
rect 1254 2366 1258 2532
rect 1278 2366 1282 2532
rect 1302 2366 1306 2532
rect 1326 2366 1330 2532
rect 1350 2366 1354 2532
rect 1374 2366 1378 2532
rect 1398 2366 1402 2532
rect 1422 2366 1426 2532
rect 1446 2366 1450 2532
rect 1470 2366 1474 2532
rect 1494 2366 1498 2532
rect 1518 2366 1522 2532
rect 1542 2366 1546 2532
rect 1566 2366 1570 2532
rect 1590 2366 1594 2532
rect 1614 2366 1618 2532
rect 1638 2366 1642 2532
rect 1662 2366 1666 2532
rect 1686 2366 1690 2532
rect 1710 2366 1714 2532
rect 1734 2366 1738 2532
rect 1758 2366 1762 2532
rect 1782 2366 1786 2532
rect 1795 2405 1800 2415
rect 1806 2405 1810 2532
rect 1805 2391 1810 2405
rect 1795 2381 1800 2391
rect 1805 2367 1810 2381
rect 1806 2366 1810 2367
rect 1830 2366 1834 2532
rect 1854 2366 1858 2532
rect 1878 2366 1882 2532
rect 1902 2366 1906 2532
rect 1926 2366 1930 2532
rect 1950 2366 1954 2532
rect 1974 2366 1978 2532
rect 1987 2525 1992 2532
rect 1998 2525 2002 2532
rect 1997 2511 2002 2525
rect 1987 2453 1992 2463
rect 1997 2439 2002 2453
rect 2011 2449 2019 2453
rect 2005 2439 2011 2449
rect 1987 2381 1992 2391
rect 1998 2381 2002 2439
rect 1997 2367 2002 2381
rect 2011 2377 2019 2381
rect 2005 2367 2011 2377
rect 1987 2366 2019 2367
rect -2393 2364 2019 2366
rect -2371 2318 -2366 2364
rect -2348 2318 -2343 2364
rect -2325 2318 -2320 2364
rect -2080 2363 -1906 2364
rect -2080 2362 -2036 2363
rect -2080 2356 -2054 2362
rect -2309 2348 -2301 2354
rect -2317 2338 -2309 2348
rect -2070 2347 -2040 2354
rect -2054 2339 -2040 2342
rect -2000 2337 -1992 2363
rect -1920 2362 -1906 2363
rect -1850 2356 -1846 2364
rect -1840 2356 -1792 2364
rect -1969 2344 -1966 2353
rect -1850 2349 -1802 2354
rect -1906 2347 -1802 2349
rect -1655 2348 -1647 2354
rect -1906 2346 -1850 2347
rect -1846 2339 -1802 2345
rect -1663 2338 -1655 2348
rect -1860 2337 -1798 2338
rect -2078 2330 -2070 2337
rect -2309 2320 -2301 2326
rect -2317 2318 -2309 2320
rect -2154 2318 -2145 2328
rect -2044 2327 -2040 2332
rect -2028 2330 -1945 2337
rect -1929 2330 -1794 2337
rect -2070 2320 -2040 2327
rect -2044 2318 -2028 2320
rect -2000 2318 -1992 2330
rect -1860 2329 -1798 2330
rect -1850 2320 -1802 2327
rect -1655 2320 -1647 2326
rect -1978 2318 -1942 2319
rect -1663 2318 -1655 2320
rect -1642 2318 -1637 2364
rect -1619 2318 -1614 2364
rect -1530 2318 -1526 2364
rect -1506 2318 -1502 2364
rect -1482 2318 -1478 2364
rect -1458 2319 -1454 2364
rect -1469 2318 -1435 2319
rect -2393 2316 -1435 2318
rect -2371 2222 -2366 2316
rect -2348 2222 -2343 2316
rect -2325 2278 -2320 2316
rect -2317 2310 -2309 2316
rect -2145 2312 -2138 2316
rect -2070 2312 -2054 2316
rect -2078 2303 -2054 2310
rect -2062 2278 -2032 2279
rect -2000 2278 -1992 2316
rect -1846 2312 -1802 2316
rect -1846 2302 -1792 2311
rect -1663 2310 -1655 2316
rect -1942 2280 -1937 2292
rect -1850 2289 -1822 2290
rect -1850 2285 -1802 2289
rect -2325 2270 -2317 2278
rect -2062 2276 -1961 2278
rect -2325 2250 -2320 2270
rect -2317 2262 -2309 2270
rect -2062 2263 -2040 2274
rect -2032 2269 -1961 2276
rect -1947 2270 -1942 2278
rect -1842 2276 -1794 2279
rect -2070 2258 -2022 2262
rect -2325 2234 -2317 2250
rect -2325 2222 -2320 2234
rect -2309 2222 -2301 2234
rect -2000 2222 -1992 2269
rect -1942 2268 -1937 2270
rect -1932 2260 -1927 2268
rect -1912 2265 -1896 2271
rect -1842 2263 -1802 2274
rect -1671 2270 -1663 2278
rect -1663 2262 -1655 2270
rect -1850 2258 -1680 2262
rect -1671 2234 -1663 2250
rect -1655 2222 -1647 2234
rect -1642 2222 -1637 2316
rect -1619 2222 -1614 2316
rect -1530 2222 -1526 2316
rect -1506 2222 -1502 2316
rect -1482 2222 -1478 2316
rect -1469 2309 -1464 2316
rect -1458 2309 -1454 2316
rect -1459 2295 -1454 2309
rect -1469 2270 -1435 2271
rect -1434 2270 -1430 2364
rect -1410 2270 -1406 2364
rect -1386 2270 -1382 2364
rect -1362 2270 -1358 2364
rect -1338 2270 -1334 2364
rect -1314 2270 -1310 2364
rect -1290 2270 -1286 2364
rect -1266 2270 -1262 2364
rect -1242 2270 -1238 2364
rect -1218 2270 -1214 2364
rect -1194 2270 -1190 2364
rect -1170 2270 -1166 2364
rect -1146 2270 -1142 2364
rect -1122 2270 -1118 2364
rect -1098 2270 -1094 2364
rect -1074 2270 -1070 2364
rect -1050 2270 -1046 2364
rect -1026 2270 -1022 2364
rect -1013 2285 -1008 2295
rect -1002 2285 -998 2364
rect -1003 2271 -998 2285
rect -978 2270 -974 2364
rect -954 2270 -950 2364
rect -930 2270 -926 2364
rect -906 2270 -902 2364
rect -882 2270 -878 2364
rect -858 2270 -854 2364
rect -834 2270 -830 2364
rect -810 2270 -806 2364
rect -786 2270 -782 2364
rect -762 2270 -758 2364
rect -738 2270 -734 2364
rect -714 2270 -710 2364
rect -690 2363 -686 2364
rect -690 2339 -683 2363
rect -690 2270 -686 2339
rect -666 2270 -662 2364
rect -642 2270 -638 2364
rect -618 2270 -614 2364
rect -594 2270 -590 2364
rect -570 2270 -566 2364
rect -546 2270 -542 2364
rect -522 2270 -518 2364
rect -498 2270 -494 2364
rect -474 2270 -470 2364
rect -450 2270 -446 2364
rect -426 2270 -422 2364
rect -402 2270 -398 2364
rect -378 2270 -374 2364
rect -354 2270 -350 2364
rect -330 2270 -326 2364
rect -306 2270 -302 2364
rect -282 2270 -278 2364
rect -258 2270 -254 2364
rect -234 2270 -230 2364
rect -210 2270 -206 2364
rect -186 2270 -182 2364
rect -162 2270 -158 2364
rect -138 2270 -134 2364
rect -114 2270 -110 2364
rect -90 2270 -86 2364
rect -66 2270 -62 2364
rect -42 2270 -38 2364
rect -18 2270 -14 2364
rect 6 2270 10 2364
rect 30 2270 34 2364
rect 54 2270 58 2364
rect 78 2270 82 2364
rect 102 2270 106 2364
rect 126 2270 130 2364
rect 150 2270 154 2364
rect 174 2270 178 2364
rect 198 2270 202 2364
rect 222 2270 226 2364
rect 246 2270 250 2364
rect 270 2270 274 2364
rect 294 2270 298 2364
rect 318 2270 322 2364
rect 342 2270 346 2364
rect 366 2270 370 2364
rect 390 2270 394 2364
rect 414 2270 418 2364
rect 438 2270 442 2364
rect 462 2270 466 2364
rect 486 2270 490 2364
rect 510 2270 514 2364
rect 534 2270 538 2364
rect 558 2270 562 2364
rect 582 2270 586 2364
rect 606 2270 610 2364
rect 630 2270 634 2364
rect 654 2270 658 2364
rect 678 2270 682 2364
rect 702 2270 706 2364
rect 726 2270 730 2364
rect 750 2270 754 2364
rect 774 2270 778 2364
rect 798 2270 802 2364
rect 822 2270 826 2364
rect 846 2270 850 2364
rect 870 2270 874 2364
rect 894 2270 898 2364
rect 918 2270 922 2364
rect 942 2270 946 2364
rect 966 2270 970 2364
rect 990 2270 994 2364
rect 1014 2270 1018 2364
rect 1038 2270 1042 2364
rect 1062 2270 1066 2364
rect 1086 2270 1090 2364
rect 1110 2270 1114 2364
rect 1134 2270 1138 2364
rect 1158 2270 1162 2364
rect 1182 2270 1186 2364
rect 1206 2270 1210 2364
rect 1230 2270 1234 2364
rect 1254 2270 1258 2364
rect 1278 2270 1282 2364
rect 1302 2270 1306 2364
rect 1326 2270 1330 2364
rect 1350 2270 1354 2364
rect 1374 2270 1378 2364
rect 1398 2270 1402 2364
rect 1422 2270 1426 2364
rect 1446 2270 1450 2364
rect 1470 2270 1474 2364
rect 1494 2270 1498 2364
rect 1518 2270 1522 2364
rect 1542 2270 1546 2364
rect 1566 2270 1570 2364
rect 1590 2270 1594 2364
rect 1614 2270 1618 2364
rect 1638 2270 1642 2364
rect 1662 2270 1666 2364
rect 1686 2270 1690 2364
rect 1710 2270 1714 2364
rect 1734 2270 1738 2364
rect 1758 2270 1762 2364
rect 1782 2270 1786 2364
rect 1806 2270 1810 2364
rect 1830 2339 1834 2364
rect 1830 2291 1837 2339
rect 1830 2270 1834 2291
rect 1854 2270 1858 2364
rect 1878 2270 1882 2364
rect 1902 2270 1906 2364
rect 1926 2270 1930 2364
rect 1950 2270 1954 2364
rect 1974 2270 1978 2364
rect 1987 2357 1992 2364
rect 2005 2363 2019 2364
rect 1997 2343 2002 2357
rect 1998 2271 2002 2343
rect 1987 2270 2019 2271
rect -1469 2268 2019 2270
rect -1469 2261 -1464 2268
rect -1459 2247 -1454 2261
rect -1458 2222 -1454 2247
rect -1434 2243 -1430 2268
rect -2393 2220 -1437 2222
rect -2371 2126 -2366 2220
rect -2348 2126 -2343 2220
rect -2325 2218 -2320 2220
rect -2317 2218 -2309 2220
rect -2325 2206 -2317 2218
rect -2061 2207 -2046 2208
rect -2325 2190 -2320 2206
rect -2309 2194 -2301 2206
rect -2070 2200 -2046 2207
rect -2000 2202 -1992 2220
rect -1974 2218 -1960 2220
rect -1663 2218 -1655 2220
rect -1960 2217 -1944 2218
rect -1980 2202 -1932 2207
rect -1671 2206 -1663 2218
rect -2061 2198 -2046 2200
rect -2032 2200 -1932 2202
rect -2032 2198 -1980 2200
rect -2317 2190 -2309 2194
rect -2062 2192 -2061 2198
rect -2062 2190 -2051 2191
rect -2325 2178 -2317 2190
rect -2062 2183 -2032 2190
rect -2062 2182 -2051 2183
rect -2325 2158 -2320 2178
rect -2325 2150 -2317 2158
rect -2325 2130 -2320 2150
rect -2317 2142 -2309 2150
rect -2325 2126 -2317 2130
rect -2000 2126 -1992 2198
rect -1655 2194 -1647 2206
rect -1990 2182 -1924 2191
rect -1904 2189 -1874 2191
rect -1842 2182 -1680 2191
rect -1663 2190 -1655 2194
rect -1671 2178 -1663 2190
rect -1671 2150 -1663 2158
rect -1663 2142 -1655 2150
rect -1671 2126 -1663 2130
rect -1642 2126 -1637 2220
rect -1619 2126 -1614 2220
rect -1530 2126 -1526 2220
rect -1506 2126 -1502 2220
rect -1482 2126 -1478 2220
rect -1458 2126 -1454 2220
rect -1451 2219 -1437 2220
rect -1434 2219 -1427 2243
rect -1434 2174 -1427 2195
rect -1410 2174 -1406 2268
rect -1386 2174 -1382 2268
rect -1362 2174 -1358 2268
rect -1338 2174 -1334 2268
rect -1314 2174 -1310 2268
rect -1290 2174 -1286 2268
rect -1266 2174 -1262 2268
rect -1242 2174 -1238 2268
rect -1218 2174 -1214 2268
rect -1194 2174 -1190 2268
rect -1170 2174 -1166 2268
rect -1146 2174 -1142 2268
rect -1122 2174 -1118 2268
rect -1098 2174 -1094 2268
rect -1074 2174 -1070 2268
rect -1050 2174 -1046 2268
rect -1026 2174 -1022 2268
rect -1013 2237 -1008 2247
rect -1003 2223 -998 2237
rect -1002 2174 -998 2223
rect -978 2219 -974 2268
rect -978 2195 -971 2219
rect -954 2174 -950 2268
rect -930 2174 -926 2268
rect -906 2174 -902 2268
rect -882 2174 -878 2268
rect -858 2174 -854 2268
rect -834 2174 -830 2268
rect -810 2174 -806 2268
rect -786 2174 -782 2268
rect -762 2174 -758 2268
rect -738 2174 -734 2268
rect -714 2174 -710 2268
rect -690 2174 -686 2268
rect -666 2174 -662 2268
rect -642 2174 -638 2268
rect -618 2174 -614 2268
rect -594 2174 -590 2268
rect -570 2174 -566 2268
rect -546 2174 -542 2268
rect -522 2174 -518 2268
rect -498 2174 -494 2268
rect -474 2174 -470 2268
rect -450 2174 -446 2268
rect -426 2174 -422 2268
rect -402 2174 -398 2268
rect -378 2174 -374 2268
rect -354 2174 -350 2268
rect -330 2174 -326 2268
rect -306 2174 -302 2268
rect -282 2174 -278 2268
rect -258 2174 -254 2268
rect -234 2174 -230 2268
rect -210 2174 -206 2268
rect -186 2174 -182 2268
rect -162 2174 -158 2268
rect -138 2174 -134 2268
rect -114 2175 -110 2268
rect -125 2174 -91 2175
rect -1451 2172 -91 2174
rect -1451 2171 -1437 2172
rect -1434 2171 -1427 2172
rect -1434 2126 -1430 2171
rect -1410 2126 -1406 2172
rect -1386 2126 -1382 2172
rect -1362 2126 -1358 2172
rect -1338 2126 -1334 2172
rect -1314 2126 -1310 2172
rect -1290 2126 -1286 2172
rect -1266 2126 -1262 2172
rect -1242 2126 -1238 2172
rect -1218 2126 -1214 2172
rect -1194 2126 -1190 2172
rect -1170 2126 -1166 2172
rect -1146 2126 -1142 2172
rect -1122 2126 -1118 2172
rect -1098 2126 -1094 2172
rect -1074 2126 -1070 2172
rect -1050 2126 -1046 2172
rect -1026 2126 -1022 2172
rect -1002 2126 -998 2172
rect -978 2147 -971 2171
rect -978 2126 -974 2147
rect -954 2126 -950 2172
rect -930 2126 -926 2172
rect -906 2126 -902 2172
rect -882 2126 -878 2172
rect -858 2126 -854 2172
rect -834 2126 -830 2172
rect -810 2126 -806 2172
rect -786 2126 -782 2172
rect -762 2126 -758 2172
rect -738 2126 -734 2172
rect -714 2126 -710 2172
rect -690 2126 -686 2172
rect -666 2126 -662 2172
rect -642 2126 -638 2172
rect -618 2126 -614 2172
rect -594 2126 -590 2172
rect -570 2126 -566 2172
rect -546 2126 -542 2172
rect -522 2126 -518 2172
rect -498 2126 -494 2172
rect -474 2126 -470 2172
rect -450 2126 -446 2172
rect -426 2126 -422 2172
rect -402 2126 -398 2172
rect -378 2126 -374 2172
rect -354 2126 -350 2172
rect -330 2126 -326 2172
rect -306 2126 -302 2172
rect -282 2126 -278 2172
rect -258 2126 -254 2172
rect -234 2126 -230 2172
rect -210 2126 -206 2172
rect -186 2126 -182 2172
rect -162 2126 -158 2172
rect -138 2126 -134 2172
rect -125 2165 -120 2172
rect -114 2165 -110 2172
rect -115 2151 -110 2165
rect -114 2126 -110 2151
rect -90 2126 -86 2268
rect -66 2126 -62 2268
rect -42 2126 -38 2268
rect -18 2126 -14 2268
rect 6 2126 10 2268
rect 30 2126 34 2268
rect 54 2126 58 2268
rect 78 2126 82 2268
rect 102 2126 106 2268
rect 126 2126 130 2268
rect 150 2126 154 2268
rect 174 2126 178 2268
rect 198 2126 202 2268
rect 222 2126 226 2268
rect 246 2126 250 2268
rect 270 2126 274 2268
rect 294 2126 298 2268
rect 318 2126 322 2268
rect 342 2126 346 2268
rect 366 2126 370 2268
rect 390 2126 394 2268
rect 414 2126 418 2268
rect 438 2126 442 2268
rect 462 2126 466 2268
rect 486 2126 490 2268
rect 510 2126 514 2268
rect 534 2126 538 2268
rect 558 2126 562 2268
rect 582 2126 586 2268
rect 606 2126 610 2268
rect 630 2126 634 2268
rect 654 2126 658 2268
rect 678 2126 682 2268
rect 702 2126 706 2268
rect 726 2126 730 2268
rect 750 2126 754 2268
rect 774 2126 778 2268
rect 798 2126 802 2268
rect 822 2126 826 2268
rect 846 2126 850 2268
rect 870 2126 874 2268
rect 894 2126 898 2268
rect 918 2126 922 2268
rect 942 2126 946 2268
rect 966 2126 970 2268
rect 990 2126 994 2268
rect 1014 2126 1018 2268
rect 1038 2126 1042 2268
rect 1062 2126 1066 2268
rect 1086 2126 1090 2268
rect 1110 2126 1114 2268
rect 1134 2126 1138 2268
rect 1158 2126 1162 2268
rect 1182 2126 1186 2268
rect 1206 2126 1210 2268
rect 1230 2126 1234 2268
rect 1243 2213 1248 2223
rect 1254 2213 1258 2268
rect 1253 2199 1258 2213
rect 1243 2189 1248 2199
rect 1253 2175 1258 2189
rect 1254 2126 1258 2175
rect 1278 2147 1282 2268
rect -2393 2124 1275 2126
rect -2371 2078 -2366 2124
rect -2348 2078 -2343 2124
rect -2325 2116 -2317 2124
rect -2018 2123 -2004 2124
rect -2000 2123 -1992 2124
rect -2072 2122 -1928 2123
rect -2072 2116 -2053 2122
rect -2325 2100 -2320 2116
rect -2317 2114 -2309 2116
rect -2309 2102 -2301 2114
rect -2092 2107 -2062 2112
rect -2317 2100 -2309 2102
rect -2325 2088 -2317 2100
rect -2098 2094 -2096 2105
rect -2092 2094 -2084 2107
rect -2000 2106 -1992 2122
rect -1972 2116 -1928 2122
rect -1924 2116 -1918 2124
rect -1671 2116 -1663 2124
rect -1663 2114 -1655 2116
rect -2083 2096 -2062 2105
rect -2027 2104 -1992 2106
rect -2018 2096 -2002 2104
rect -2000 2096 -1992 2104
rect -2100 2089 -2096 2094
rect -2083 2089 -2053 2094
rect -2003 2092 -1990 2096
rect -1972 2094 -1964 2103
rect -1928 2102 -1924 2105
rect -1655 2102 -1647 2114
rect -1663 2100 -1655 2102
rect -2325 2078 -2320 2088
rect -2317 2086 -2309 2088
rect -2309 2078 -2301 2086
rect -2004 2082 -2003 2092
rect -2062 2078 -2012 2080
rect -2000 2078 -1992 2092
rect -1972 2089 -1924 2094
rect -1864 2089 -1796 2095
rect -1671 2088 -1663 2100
rect -1663 2086 -1655 2088
rect -1864 2078 -1796 2079
rect -1655 2078 -1647 2086
rect -1642 2078 -1637 2124
rect -1619 2078 -1614 2124
rect -1530 2078 -1526 2124
rect -1506 2078 -1502 2124
rect -1482 2078 -1478 2124
rect -1458 2078 -1454 2124
rect -1434 2078 -1430 2124
rect -1410 2078 -1406 2124
rect -1386 2078 -1382 2124
rect -1362 2078 -1358 2124
rect -1338 2078 -1334 2124
rect -1314 2078 -1310 2124
rect -1290 2078 -1286 2124
rect -1266 2078 -1262 2124
rect -1242 2078 -1238 2124
rect -1218 2078 -1214 2124
rect -1194 2078 -1190 2124
rect -1170 2078 -1166 2124
rect -1146 2078 -1142 2124
rect -1122 2078 -1118 2124
rect -1098 2078 -1094 2124
rect -1074 2078 -1070 2124
rect -1050 2079 -1046 2124
rect -1061 2078 -1027 2079
rect -2393 2076 -1027 2078
rect -2371 2030 -2366 2076
rect -2348 2030 -2343 2076
rect -2325 2072 -2320 2076
rect -2309 2074 -2301 2076
rect -2317 2072 -2309 2074
rect -2325 2060 -2317 2072
rect -2325 2030 -2320 2060
rect -2317 2058 -2309 2060
rect -2092 2046 -2062 2048
rect -2094 2042 -2062 2046
rect -2000 2030 -1992 2076
rect -1655 2074 -1647 2076
rect -1663 2072 -1655 2074
rect -1671 2060 -1663 2072
rect -1663 2058 -1655 2060
rect -1854 2046 -1806 2048
rect -1854 2042 -1680 2046
rect -1642 2030 -1637 2076
rect -1619 2030 -1614 2076
rect -1530 2030 -1526 2076
rect -1506 2030 -1502 2076
rect -1482 2030 -1478 2076
rect -1458 2030 -1454 2076
rect -1434 2030 -1430 2076
rect -1410 2030 -1406 2076
rect -1386 2030 -1382 2076
rect -1362 2030 -1358 2076
rect -1338 2030 -1334 2076
rect -1314 2030 -1310 2076
rect -1290 2030 -1286 2076
rect -1266 2030 -1262 2076
rect -1242 2030 -1238 2076
rect -1218 2030 -1214 2076
rect -1194 2030 -1190 2076
rect -1170 2030 -1166 2076
rect -1146 2030 -1142 2076
rect -1122 2030 -1118 2076
rect -1098 2030 -1094 2076
rect -1074 2030 -1070 2076
rect -1061 2069 -1056 2076
rect -1050 2069 -1046 2076
rect -1051 2055 -1046 2069
rect -1061 2045 -1056 2055
rect -1051 2031 -1046 2045
rect -1050 2030 -1046 2031
rect -1026 2030 -1022 2124
rect -1002 2030 -998 2124
rect -978 2030 -974 2124
rect -954 2030 -950 2124
rect -930 2030 -926 2124
rect -906 2030 -902 2124
rect -882 2030 -878 2124
rect -858 2030 -854 2124
rect -834 2030 -830 2124
rect -810 2030 -806 2124
rect -786 2030 -782 2124
rect -762 2030 -758 2124
rect -738 2030 -734 2124
rect -714 2030 -710 2124
rect -690 2030 -686 2124
rect -666 2030 -662 2124
rect -642 2030 -638 2124
rect -618 2030 -614 2124
rect -594 2030 -590 2124
rect -570 2030 -566 2124
rect -546 2030 -542 2124
rect -522 2030 -518 2124
rect -498 2030 -494 2124
rect -474 2030 -470 2124
rect -450 2030 -446 2124
rect -426 2030 -422 2124
rect -402 2030 -398 2124
rect -378 2030 -374 2124
rect -354 2030 -350 2124
rect -330 2030 -326 2124
rect -306 2030 -302 2124
rect -282 2030 -278 2124
rect -258 2030 -254 2124
rect -234 2030 -230 2124
rect -210 2030 -206 2124
rect -186 2030 -182 2124
rect -162 2030 -158 2124
rect -138 2030 -134 2124
rect -114 2030 -110 2124
rect -90 2099 -86 2124
rect -90 2075 -83 2099
rect -90 2030 -86 2075
rect -66 2030 -62 2124
rect -42 2030 -38 2124
rect -18 2030 -14 2124
rect 6 2030 10 2124
rect 30 2030 34 2124
rect 54 2030 58 2124
rect 78 2030 82 2124
rect 102 2030 106 2124
rect 126 2030 130 2124
rect 150 2030 154 2124
rect 174 2030 178 2124
rect 198 2030 202 2124
rect 222 2030 226 2124
rect 246 2030 250 2124
rect 270 2030 274 2124
rect 294 2030 298 2124
rect 318 2030 322 2124
rect 342 2030 346 2124
rect 366 2030 370 2124
rect 390 2030 394 2124
rect 414 2030 418 2124
rect 438 2030 442 2124
rect 462 2030 466 2124
rect 486 2030 490 2124
rect 510 2030 514 2124
rect 534 2030 538 2124
rect 558 2030 562 2124
rect 582 2030 586 2124
rect 606 2030 610 2124
rect 630 2030 634 2124
rect 654 2030 658 2124
rect 678 2030 682 2124
rect 702 2030 706 2124
rect 726 2030 730 2124
rect 750 2030 754 2124
rect 774 2030 778 2124
rect 798 2030 802 2124
rect 822 2030 826 2124
rect 846 2030 850 2124
rect 870 2030 874 2124
rect 894 2030 898 2124
rect 918 2030 922 2124
rect 942 2030 946 2124
rect 966 2030 970 2124
rect 990 2030 994 2124
rect 1014 2030 1018 2124
rect 1038 2030 1042 2124
rect 1051 2093 1056 2103
rect 1062 2093 1066 2124
rect 1061 2079 1066 2093
rect 1051 2069 1056 2079
rect 1061 2055 1066 2069
rect 1062 2030 1066 2055
rect 1086 2030 1090 2124
rect 1110 2030 1114 2124
rect 1134 2030 1138 2124
rect 1158 2030 1162 2124
rect 1182 2030 1186 2124
rect 1206 2030 1210 2124
rect 1230 2030 1234 2124
rect 1254 2030 1258 2124
rect 1261 2123 1275 2124
rect 1278 2099 1285 2147
rect 1278 2030 1282 2099
rect 1302 2030 1306 2268
rect 1326 2030 1330 2268
rect 1350 2030 1354 2268
rect 1374 2030 1378 2268
rect 1398 2030 1402 2268
rect 1422 2030 1426 2268
rect 1446 2030 1450 2268
rect 1470 2030 1474 2268
rect 1494 2030 1498 2268
rect 1518 2030 1522 2268
rect 1542 2030 1546 2268
rect 1566 2030 1570 2268
rect 1590 2030 1594 2268
rect 1614 2030 1618 2268
rect 1638 2030 1642 2268
rect 1662 2030 1666 2268
rect 1686 2030 1690 2268
rect 1710 2030 1714 2268
rect 1734 2030 1738 2268
rect 1758 2030 1762 2268
rect 1782 2030 1786 2268
rect 1806 2030 1810 2268
rect 1830 2030 1834 2268
rect 1854 2030 1858 2268
rect 1878 2030 1882 2268
rect 1902 2030 1906 2268
rect 1915 2045 1920 2055
rect 1926 2045 1930 2268
rect 1939 2189 1944 2199
rect 1950 2189 1954 2268
rect 1963 2237 1968 2247
rect 1974 2237 1978 2268
rect 1987 2261 1992 2268
rect 1998 2261 2002 2268
rect 2005 2267 2019 2268
rect 1997 2247 2002 2261
rect 1973 2223 1978 2237
rect 1949 2175 1954 2189
rect 1939 2117 1944 2127
rect 1949 2103 1954 2117
rect 1963 2113 1971 2117
rect 1957 2103 1963 2113
rect 1939 2069 1944 2079
rect 1950 2069 1954 2103
rect 1949 2055 1954 2069
rect 1925 2031 1930 2045
rect 1915 2030 1949 2031
rect -2393 2028 1949 2030
rect -2371 2006 -2366 2028
rect -2348 2006 -2343 2028
rect -2325 2006 -2320 2028
rect -2072 2026 -2036 2027
rect -2072 2020 -2054 2026
rect -2309 2012 -2301 2020
rect -2317 2006 -2309 2012
rect -2092 2011 -2062 2016
rect -2000 2007 -1992 2028
rect -1938 2027 -1906 2028
rect -1920 2026 -1906 2027
rect -1806 2020 -1680 2026
rect -1854 2011 -1806 2016
rect -1655 2012 -1647 2020
rect -1982 2007 -1966 2008
rect -2000 2006 -1966 2007
rect -1846 2006 -1806 2009
rect -1663 2006 -1655 2012
rect -1642 2006 -1637 2028
rect -1619 2006 -1614 2028
rect -1530 2006 -1526 2028
rect -1506 2006 -1502 2028
rect -1482 2006 -1478 2028
rect -1458 2006 -1454 2028
rect -1434 2006 -1430 2028
rect -1410 2006 -1406 2028
rect -1386 2006 -1382 2028
rect -1362 2006 -1358 2028
rect -1338 2006 -1334 2028
rect -1314 2006 -1310 2028
rect -1290 2006 -1286 2028
rect -1266 2006 -1262 2028
rect -1242 2006 -1238 2028
rect -1218 2006 -1214 2028
rect -1194 2006 -1190 2028
rect -1170 2006 -1166 2028
rect -1146 2006 -1142 2028
rect -1122 2006 -1118 2028
rect -1098 2006 -1094 2028
rect -1074 2006 -1070 2028
rect -1050 2006 -1046 2028
rect -1026 2006 -1022 2028
rect -1002 2006 -998 2028
rect -978 2006 -974 2028
rect -954 2006 -950 2028
rect -930 2006 -926 2028
rect -906 2006 -902 2028
rect -882 2006 -878 2028
rect -858 2006 -854 2028
rect -834 2006 -830 2028
rect -810 2006 -806 2028
rect -786 2006 -782 2028
rect -762 2006 -758 2028
rect -738 2006 -734 2028
rect -714 2007 -710 2028
rect -725 2006 -691 2007
rect -2393 2004 -691 2006
rect -2371 1982 -2366 2004
rect -2348 1982 -2343 2004
rect -2325 1982 -2320 2004
rect -2000 2002 -1966 2004
rect -2309 1984 -2301 1992
rect -2062 1991 -2054 1998
rect -2092 1984 -2084 1991
rect -2062 1984 -2026 1986
rect -2317 1982 -2309 1984
rect -2062 1982 -2012 1984
rect -2000 1982 -1992 2002
rect -1982 2001 -1966 2002
rect -1846 2000 -1806 2004
rect -1846 1993 -1798 1998
rect -1806 1991 -1798 1993
rect -1854 1989 -1846 1991
rect -1854 1984 -1806 1989
rect -1655 1984 -1647 1992
rect -1864 1982 -1796 1983
rect -1663 1982 -1655 1984
rect -1642 1982 -1637 2004
rect -1619 1982 -1614 2004
rect -1530 1982 -1526 2004
rect -1506 1982 -1502 2004
rect -1482 1982 -1478 2004
rect -1458 1982 -1454 2004
rect -1434 1982 -1430 2004
rect -1410 1982 -1406 2004
rect -1386 1982 -1382 2004
rect -1362 1982 -1358 2004
rect -1338 1982 -1334 2004
rect -1314 1982 -1310 2004
rect -1290 1982 -1286 2004
rect -1266 1982 -1262 2004
rect -1242 1982 -1238 2004
rect -1218 1982 -1214 2004
rect -1194 1982 -1190 2004
rect -1170 1982 -1166 2004
rect -1146 1982 -1142 2004
rect -1122 1982 -1118 2004
rect -1098 1982 -1094 2004
rect -1074 1982 -1070 2004
rect -1050 1982 -1046 2004
rect -1026 2003 -1022 2004
rect -2393 1980 -1029 1982
rect -2371 1934 -2366 1980
rect -2348 1934 -2343 1980
rect -2325 1944 -2320 1980
rect -2317 1976 -2309 1980
rect -2062 1976 -2054 1980
rect -2154 1972 -2138 1974
rect -2057 1972 -2054 1976
rect -2292 1966 -2054 1972
rect -2052 1966 -2044 1976
rect -2092 1950 -2062 1952
rect -2094 1946 -2062 1950
rect -2325 1934 -2317 1944
rect -2095 1936 -2084 1940
rect -2000 1937 -1992 1980
rect -1846 1973 -1806 1980
rect -1663 1976 -1655 1980
rect -1846 1966 -1680 1972
rect -1854 1950 -1806 1952
rect -1854 1946 -1680 1950
rect -2119 1934 -2069 1936
rect -2054 1934 -1892 1937
rect -1671 1934 -1663 1944
rect -1642 1934 -1637 1980
rect -1619 1934 -1614 1980
rect -1530 1934 -1526 1980
rect -1506 1934 -1502 1980
rect -1482 1934 -1478 1980
rect -1458 1934 -1454 1980
rect -1434 1934 -1430 1980
rect -1410 1934 -1406 1980
rect -1386 1934 -1382 1980
rect -1362 1934 -1358 1980
rect -1338 1934 -1334 1980
rect -1314 1934 -1310 1980
rect -1290 1934 -1286 1980
rect -1266 1934 -1262 1980
rect -1242 1934 -1238 1980
rect -1218 1934 -1214 1980
rect -1194 1934 -1190 1980
rect -1170 1934 -1166 1980
rect -1146 1934 -1142 1980
rect -1122 1934 -1118 1980
rect -1098 1934 -1094 1980
rect -1074 1934 -1070 1980
rect -1050 1934 -1046 1980
rect -1043 1979 -1029 1980
rect -1026 1955 -1019 2003
rect -1026 1934 -1022 1955
rect -1002 1934 -998 2004
rect -978 1934 -974 2004
rect -954 1934 -950 2004
rect -930 1934 -926 2004
rect -906 1934 -902 2004
rect -882 1934 -878 2004
rect -858 1934 -854 2004
rect -834 1934 -830 2004
rect -810 1934 -806 2004
rect -786 1934 -782 2004
rect -762 1934 -758 2004
rect -738 1934 -734 2004
rect -725 1997 -720 2004
rect -714 1997 -710 2004
rect -715 1983 -710 1997
rect -725 1958 -691 1959
rect -690 1958 -686 2028
rect -666 1958 -662 2028
rect -642 1958 -638 2028
rect -618 1958 -614 2028
rect -594 1958 -590 2028
rect -570 1958 -566 2028
rect -546 1958 -542 2028
rect -522 1958 -518 2028
rect -498 1958 -494 2028
rect -474 1958 -470 2028
rect -450 1958 -446 2028
rect -426 1958 -422 2028
rect -402 1958 -398 2028
rect -378 1958 -374 2028
rect -354 1958 -350 2028
rect -330 1958 -326 2028
rect -306 1958 -302 2028
rect -282 1958 -278 2028
rect -258 1958 -254 2028
rect -234 1958 -230 2028
rect -210 1958 -206 2028
rect -186 1958 -182 2028
rect -162 1958 -158 2028
rect -138 1958 -134 2028
rect -114 1958 -110 2028
rect -90 1958 -86 2028
rect -66 1958 -62 2028
rect -42 1958 -38 2028
rect -18 1958 -14 2028
rect 6 1958 10 2028
rect 30 1958 34 2028
rect 54 1958 58 2028
rect 78 1958 82 2028
rect 102 1958 106 2028
rect 126 1958 130 2028
rect 150 1958 154 2028
rect 174 1958 178 2028
rect 198 1958 202 2028
rect 222 1958 226 2028
rect 246 1958 250 2028
rect 270 1958 274 2028
rect 294 1958 298 2028
rect 318 1958 322 2028
rect 342 1958 346 2028
rect 366 1958 370 2028
rect 390 1958 394 2028
rect 414 1958 418 2028
rect 438 1958 442 2028
rect 462 1958 466 2028
rect 486 1958 490 2028
rect 510 1958 514 2028
rect 534 1958 538 2028
rect 558 1958 562 2028
rect 582 1958 586 2028
rect 606 1958 610 2028
rect 630 1958 634 2028
rect 654 1958 658 2028
rect 678 1958 682 2028
rect 702 1958 706 2028
rect 726 1958 730 2028
rect 750 1958 754 2028
rect 774 1958 778 2028
rect 798 1958 802 2028
rect 822 1958 826 2028
rect 846 1958 850 2028
rect 870 1958 874 2028
rect 894 1958 898 2028
rect 918 1958 922 2028
rect 942 1958 946 2028
rect 966 1958 970 2028
rect 990 1958 994 2028
rect 1014 1958 1018 2028
rect 1038 1958 1042 2028
rect 1062 1958 1066 2028
rect 1086 2027 1090 2028
rect 1086 1982 1093 2027
rect 1110 1982 1114 2028
rect 1134 1982 1138 2028
rect 1158 1982 1162 2028
rect 1182 1982 1186 2028
rect 1206 1982 1210 2028
rect 1230 1982 1234 2028
rect 1254 1982 1258 2028
rect 1278 1982 1282 2028
rect 1302 1982 1306 2028
rect 1326 1982 1330 2028
rect 1350 1982 1354 2028
rect 1374 1982 1378 2028
rect 1398 1982 1402 2028
rect 1422 1982 1426 2028
rect 1446 1982 1450 2028
rect 1470 1982 1474 2028
rect 1494 1982 1498 2028
rect 1518 1982 1522 2028
rect 1542 1983 1546 2028
rect 1531 1982 1565 1983
rect 1069 1980 1565 1982
rect 1069 1979 1083 1980
rect 1086 1979 1093 1980
rect 1086 1958 1090 1979
rect 1110 1958 1114 1980
rect 1134 1958 1138 1980
rect 1158 1958 1162 1980
rect 1182 1958 1186 1980
rect 1206 1958 1210 1980
rect 1230 1958 1234 1980
rect 1254 1958 1258 1980
rect 1278 1958 1282 1980
rect 1302 1958 1306 1980
rect 1326 1958 1330 1980
rect 1350 1958 1354 1980
rect 1374 1958 1378 1980
rect 1398 1958 1402 1980
rect 1422 1958 1426 1980
rect 1446 1958 1450 1980
rect 1470 1958 1474 1980
rect 1494 1958 1498 1980
rect 1518 1958 1522 1980
rect 1531 1973 1536 1980
rect 1542 1973 1546 1980
rect 1541 1959 1546 1973
rect 1566 1958 1570 2028
rect 1590 1958 1594 2028
rect 1614 1958 1618 2028
rect 1638 1958 1642 2028
rect 1662 1958 1666 2028
rect 1686 1958 1690 2028
rect 1710 1958 1714 2028
rect 1734 1958 1738 2028
rect 1758 1958 1762 2028
rect 1782 1958 1786 2028
rect 1806 1958 1810 2028
rect 1830 1958 1834 2028
rect 1854 1958 1858 2028
rect 1878 1958 1882 2028
rect 1902 1958 1906 2028
rect 1915 2021 1920 2028
rect 1925 2007 1930 2021
rect 1926 1959 1930 2007
rect 1915 1958 1947 1959
rect -725 1956 1947 1958
rect -725 1949 -720 1956
rect -715 1935 -710 1949
rect -714 1934 -710 1935
rect -690 1934 -686 1956
rect -666 1934 -662 1956
rect -642 1934 -638 1956
rect -618 1934 -614 1956
rect -594 1934 -590 1956
rect -570 1934 -566 1956
rect -546 1934 -542 1956
rect -522 1934 -518 1956
rect -498 1934 -494 1956
rect -474 1934 -470 1956
rect -450 1934 -446 1956
rect -426 1934 -422 1956
rect -402 1934 -398 1956
rect -378 1934 -374 1956
rect -354 1934 -350 1956
rect -330 1934 -326 1956
rect -306 1934 -302 1956
rect -282 1934 -278 1956
rect -258 1934 -254 1956
rect -234 1934 -230 1956
rect -210 1934 -206 1956
rect -186 1934 -182 1956
rect -162 1934 -158 1956
rect -138 1934 -134 1956
rect -114 1934 -110 1956
rect -90 1934 -86 1956
rect -66 1934 -62 1956
rect -42 1934 -38 1956
rect -18 1934 -14 1956
rect 6 1934 10 1956
rect 30 1934 34 1956
rect 54 1934 58 1956
rect 78 1934 82 1956
rect 102 1934 106 1956
rect 126 1934 130 1956
rect 150 1934 154 1956
rect 174 1934 178 1956
rect 198 1934 202 1956
rect 222 1934 226 1956
rect 246 1934 250 1956
rect 270 1934 274 1956
rect 294 1934 298 1956
rect 318 1934 322 1956
rect 342 1934 346 1956
rect 366 1934 370 1956
rect 390 1934 394 1956
rect 414 1934 418 1956
rect 438 1934 442 1956
rect 462 1934 466 1956
rect 486 1934 490 1956
rect 510 1934 514 1956
rect 534 1934 538 1956
rect 558 1934 562 1956
rect 582 1934 586 1956
rect 606 1934 610 1956
rect 630 1934 634 1956
rect 654 1934 658 1956
rect 678 1934 682 1956
rect 702 1934 706 1956
rect 726 1934 730 1956
rect 750 1934 754 1956
rect 774 1934 778 1956
rect 798 1934 802 1956
rect 822 1934 826 1956
rect 846 1934 850 1956
rect 870 1934 874 1956
rect 894 1934 898 1956
rect 918 1934 922 1956
rect 942 1934 946 1956
rect 966 1934 970 1956
rect 990 1934 994 1956
rect 1014 1934 1018 1956
rect 1038 1934 1042 1956
rect 1062 1934 1066 1956
rect 1086 1934 1090 1956
rect 1110 1934 1114 1956
rect 1134 1934 1138 1956
rect 1158 1934 1162 1956
rect 1182 1934 1186 1956
rect 1206 1934 1210 1956
rect 1230 1934 1234 1956
rect 1254 1934 1258 1956
rect 1278 1934 1282 1956
rect 1302 1934 1306 1956
rect 1326 1934 1330 1956
rect 1350 1934 1354 1956
rect 1374 1934 1378 1956
rect 1398 1934 1402 1956
rect 1422 1934 1426 1956
rect 1446 1934 1450 1956
rect 1470 1934 1474 1956
rect 1494 1934 1498 1956
rect 1518 1934 1522 1956
rect 1531 1934 1565 1935
rect -2393 1932 1565 1934
rect -2371 1910 -2366 1932
rect -2348 1910 -2343 1932
rect -2325 1928 -2317 1932
rect -2325 1912 -2320 1928
rect -2309 1916 -2301 1928
rect -2095 1926 -2084 1932
rect -2054 1931 -1906 1932
rect -2054 1930 -2036 1931
rect -2084 1924 -2079 1926
rect -2317 1912 -2309 1916
rect -2092 1915 -2079 1922
rect -2000 1918 -1992 1931
rect -1920 1930 -1906 1931
rect -1671 1928 -1663 1932
rect -1846 1924 -1806 1926
rect -1854 1918 -1806 1922
rect -2054 1915 -1982 1918
rect -1966 1915 -1806 1918
rect -1655 1916 -1647 1928
rect -2003 1912 -1992 1915
rect -1904 1913 -1902 1915
rect -1854 1913 -1846 1915
rect -2325 1910 -2317 1912
rect -2033 1910 -1992 1912
rect -1854 1911 -1806 1913
rect -1663 1912 -1655 1916
rect -1864 1910 -1796 1911
rect -1671 1910 -1663 1912
rect -1642 1910 -1637 1932
rect -1619 1910 -1614 1932
rect -1530 1910 -1526 1932
rect -1506 1910 -1502 1932
rect -1482 1910 -1478 1932
rect -1458 1910 -1454 1932
rect -1434 1910 -1430 1932
rect -1410 1910 -1406 1932
rect -1386 1910 -1382 1932
rect -1362 1910 -1358 1932
rect -1338 1910 -1334 1932
rect -1314 1910 -1310 1932
rect -1290 1910 -1286 1932
rect -1266 1910 -1262 1932
rect -1242 1910 -1238 1932
rect -1218 1910 -1214 1932
rect -1194 1910 -1190 1932
rect -1170 1910 -1166 1932
rect -1146 1910 -1142 1932
rect -1122 1910 -1118 1932
rect -1098 1910 -1094 1932
rect -1074 1910 -1070 1932
rect -1050 1910 -1046 1932
rect -1026 1910 -1022 1932
rect -1002 1910 -998 1932
rect -978 1910 -974 1932
rect -954 1910 -950 1932
rect -930 1910 -926 1932
rect -906 1910 -902 1932
rect -882 1910 -878 1932
rect -858 1910 -854 1932
rect -834 1910 -830 1932
rect -810 1910 -806 1932
rect -786 1910 -782 1932
rect -762 1910 -758 1932
rect -738 1910 -734 1932
rect -714 1910 -710 1932
rect -690 1931 -686 1932
rect -2393 1908 -693 1910
rect -2371 1886 -2366 1908
rect -2348 1886 -2343 1908
rect -2325 1900 -2317 1908
rect -2079 1905 -2018 1908
rect -2003 1907 -1966 1908
rect -2000 1906 -1982 1907
rect -2000 1905 -1992 1906
rect -2084 1901 -2009 1905
rect -2028 1900 -2009 1901
rect -2000 1901 -1854 1905
rect -1846 1901 -1798 1908
rect -2325 1886 -2320 1900
rect -2309 1888 -2301 1900
rect -2028 1898 -2018 1900
rect -2092 1888 -2084 1895
rect -2023 1891 -2014 1898
rect -2000 1891 -1992 1901
rect -1671 1900 -1663 1908
rect -1846 1897 -1806 1899
rect -1854 1891 -1806 1895
rect -2054 1888 -1806 1891
rect -1655 1888 -1647 1900
rect -2317 1886 -2309 1888
rect -2054 1886 -2024 1888
rect -2000 1886 -1992 1888
rect -1663 1886 -1655 1888
rect -1642 1886 -1637 1908
rect -1619 1886 -1614 1908
rect -1530 1886 -1526 1908
rect -1506 1886 -1502 1908
rect -1482 1886 -1478 1908
rect -1458 1886 -1454 1908
rect -1434 1886 -1430 1908
rect -1410 1886 -1406 1908
rect -1386 1886 -1382 1908
rect -1362 1886 -1358 1908
rect -1338 1886 -1334 1908
rect -1314 1886 -1310 1908
rect -1290 1886 -1286 1908
rect -1266 1886 -1262 1908
rect -1242 1886 -1238 1908
rect -1218 1886 -1214 1908
rect -1194 1886 -1190 1908
rect -1170 1886 -1166 1908
rect -1146 1886 -1142 1908
rect -1122 1886 -1118 1908
rect -1098 1886 -1094 1908
rect -1074 1886 -1070 1908
rect -1050 1886 -1046 1908
rect -1026 1886 -1022 1908
rect -1002 1886 -998 1908
rect -978 1886 -974 1908
rect -954 1886 -950 1908
rect -930 1886 -926 1908
rect -906 1886 -902 1908
rect -882 1886 -878 1908
rect -858 1886 -854 1908
rect -834 1886 -830 1908
rect -810 1886 -806 1908
rect -786 1886 -782 1908
rect -762 1886 -758 1908
rect -738 1886 -734 1908
rect -714 1886 -710 1908
rect -707 1907 -693 1908
rect -690 1907 -683 1931
rect -666 1886 -662 1932
rect -642 1886 -638 1932
rect -618 1886 -614 1932
rect -594 1886 -590 1932
rect -570 1886 -566 1932
rect -546 1886 -542 1932
rect -522 1886 -518 1932
rect -498 1886 -494 1932
rect -474 1886 -470 1932
rect -450 1886 -446 1932
rect -426 1886 -422 1932
rect -402 1886 -398 1932
rect -378 1886 -374 1932
rect -354 1886 -350 1932
rect -330 1886 -326 1932
rect -306 1886 -302 1932
rect -282 1886 -278 1932
rect -258 1886 -254 1932
rect -234 1886 -230 1932
rect -210 1886 -206 1932
rect -186 1886 -182 1932
rect -162 1886 -158 1932
rect -138 1886 -134 1932
rect -114 1886 -110 1932
rect -90 1886 -86 1932
rect -66 1886 -62 1932
rect -42 1886 -38 1932
rect -18 1886 -14 1932
rect 6 1886 10 1932
rect 30 1886 34 1932
rect 54 1886 58 1932
rect 78 1886 82 1932
rect 102 1886 106 1932
rect 126 1886 130 1932
rect 150 1886 154 1932
rect 174 1886 178 1932
rect 198 1886 202 1932
rect 222 1886 226 1932
rect 246 1886 250 1932
rect 270 1886 274 1932
rect 294 1886 298 1932
rect 318 1886 322 1932
rect 342 1886 346 1932
rect 366 1886 370 1932
rect 390 1886 394 1932
rect 414 1886 418 1932
rect 438 1886 442 1932
rect 462 1886 466 1932
rect 486 1886 490 1932
rect 510 1887 514 1932
rect 499 1886 533 1887
rect -2393 1884 -2064 1886
rect -2060 1884 533 1886
rect -2371 1838 -2366 1884
rect -2348 1838 -2343 1884
rect -2325 1872 -2317 1884
rect -2060 1881 -2054 1884
rect -2084 1874 -2054 1881
rect -2050 1878 -2044 1880
rect -2325 1852 -2320 1872
rect -2064 1870 -2054 1874
rect -2325 1844 -2317 1852
rect -2101 1847 -2071 1850
rect -2325 1838 -2320 1844
rect -2317 1838 -2309 1844
rect -2000 1842 -1992 1884
rect -1846 1883 -1806 1884
rect -1846 1874 -1798 1881
rect -1671 1872 -1663 1884
rect -1846 1870 -1806 1872
rect -1854 1856 -1680 1860
rect -1846 1847 -1798 1850
rect -2079 1841 -2043 1842
rect -2007 1841 -1991 1842
rect -2079 1840 -2071 1841
rect -2079 1838 -2029 1840
rect -2011 1838 -1991 1841
rect -1846 1839 -1806 1845
rect -1671 1844 -1663 1852
rect -1864 1838 -1796 1839
rect -1663 1838 -1655 1844
rect -1642 1838 -1637 1884
rect -1619 1838 -1614 1884
rect -1530 1838 -1526 1884
rect -1506 1838 -1502 1884
rect -1482 1838 -1478 1884
rect -1458 1838 -1454 1884
rect -1434 1838 -1430 1884
rect -1410 1838 -1406 1884
rect -1386 1838 -1382 1884
rect -1362 1838 -1358 1884
rect -1338 1838 -1334 1884
rect -1314 1838 -1310 1884
rect -1290 1838 -1286 1884
rect -1266 1838 -1262 1884
rect -1242 1838 -1238 1884
rect -1218 1838 -1214 1884
rect -1194 1838 -1190 1884
rect -1170 1838 -1166 1884
rect -1146 1838 -1142 1884
rect -1122 1838 -1118 1884
rect -1098 1838 -1094 1884
rect -1074 1838 -1070 1884
rect -1050 1838 -1046 1884
rect -1026 1838 -1022 1884
rect -1002 1838 -998 1884
rect -978 1838 -974 1884
rect -954 1838 -950 1884
rect -930 1838 -926 1884
rect -906 1838 -902 1884
rect -882 1838 -878 1884
rect -858 1838 -854 1884
rect -834 1838 -830 1884
rect -810 1838 -806 1884
rect -786 1838 -782 1884
rect -762 1838 -758 1884
rect -738 1838 -734 1884
rect -714 1838 -710 1884
rect -690 1862 -683 1883
rect -666 1862 -662 1884
rect -642 1862 -638 1884
rect -618 1862 -614 1884
rect -594 1862 -590 1884
rect -570 1862 -566 1884
rect -546 1862 -542 1884
rect -522 1862 -518 1884
rect -498 1862 -494 1884
rect -474 1862 -470 1884
rect -450 1862 -446 1884
rect -426 1862 -422 1884
rect -402 1862 -398 1884
rect -378 1862 -374 1884
rect -354 1862 -350 1884
rect -330 1862 -326 1884
rect -306 1862 -302 1884
rect -282 1862 -278 1884
rect -258 1862 -254 1884
rect -234 1862 -230 1884
rect -210 1862 -206 1884
rect -186 1862 -182 1884
rect -162 1862 -158 1884
rect -138 1862 -134 1884
rect -114 1862 -110 1884
rect -90 1862 -86 1884
rect -66 1862 -62 1884
rect -42 1862 -38 1884
rect -18 1862 -14 1884
rect 6 1862 10 1884
rect 30 1862 34 1884
rect 54 1862 58 1884
rect 78 1862 82 1884
rect 102 1862 106 1884
rect 126 1862 130 1884
rect 150 1862 154 1884
rect 174 1862 178 1884
rect 198 1862 202 1884
rect 222 1862 226 1884
rect 246 1862 250 1884
rect 270 1862 274 1884
rect 294 1862 298 1884
rect 318 1862 322 1884
rect 342 1862 346 1884
rect 366 1862 370 1884
rect 390 1862 394 1884
rect 414 1862 418 1884
rect 438 1862 442 1884
rect 462 1862 466 1884
rect 486 1862 490 1884
rect 499 1877 504 1884
rect 510 1877 514 1884
rect 509 1863 514 1877
rect 534 1862 538 1932
rect 558 1862 562 1932
rect 582 1862 586 1932
rect 606 1862 610 1932
rect 630 1862 634 1932
rect 654 1862 658 1932
rect 678 1862 682 1932
rect 702 1862 706 1932
rect 726 1862 730 1932
rect 750 1862 754 1932
rect 774 1862 778 1932
rect 798 1862 802 1932
rect 822 1862 826 1932
rect 846 1862 850 1932
rect 870 1862 874 1932
rect 894 1862 898 1932
rect 918 1862 922 1932
rect 942 1862 946 1932
rect 966 1863 970 1932
rect 955 1862 989 1863
rect -707 1860 989 1862
rect -707 1859 -693 1860
rect -690 1859 -683 1860
rect -690 1838 -686 1859
rect -666 1838 -662 1860
rect -642 1838 -638 1860
rect -618 1838 -614 1860
rect -594 1838 -590 1860
rect -570 1838 -566 1860
rect -546 1838 -542 1860
rect -522 1838 -518 1860
rect -498 1838 -494 1860
rect -474 1838 -470 1860
rect -450 1838 -446 1860
rect -426 1838 -422 1860
rect -402 1838 -398 1860
rect -378 1838 -374 1860
rect -354 1838 -350 1860
rect -330 1838 -326 1860
rect -306 1838 -302 1860
rect -282 1839 -278 1860
rect -293 1838 -259 1839
rect -2393 1836 -259 1838
rect -2371 1790 -2366 1836
rect -2348 1790 -2343 1836
rect -2325 1824 -2320 1836
rect -2079 1834 -2071 1836
rect -2072 1832 -2071 1834
rect -2109 1827 -2101 1832
rect -2101 1825 -2079 1827
rect -2069 1825 -2068 1832
rect -2325 1816 -2317 1824
rect -2079 1820 -2071 1825
rect -2325 1796 -2320 1816
rect -2317 1808 -2309 1816
rect -2074 1811 -2071 1820
rect -2069 1816 -2068 1820
rect -2109 1802 -2079 1805
rect -2325 1790 -2317 1796
rect -2000 1790 -1992 1836
rect -1846 1834 -1806 1836
rect -1854 1829 -1806 1833
rect -1854 1827 -1846 1829
rect -1846 1825 -1806 1827
rect -1806 1823 -1798 1825
rect -1846 1820 -1798 1823
rect -1846 1807 -1806 1818
rect -1671 1816 -1663 1824
rect -1663 1808 -1655 1816
rect -1854 1802 -1680 1806
rect -1671 1790 -1663 1796
rect -1642 1790 -1637 1836
rect -1619 1790 -1614 1836
rect -1530 1790 -1526 1836
rect -1506 1790 -1502 1836
rect -1482 1790 -1478 1836
rect -1458 1790 -1454 1836
rect -1434 1790 -1430 1836
rect -1410 1790 -1406 1836
rect -1386 1790 -1382 1836
rect -1362 1790 -1358 1836
rect -1338 1790 -1334 1836
rect -1314 1790 -1310 1836
rect -1290 1790 -1286 1836
rect -1266 1790 -1262 1836
rect -1242 1790 -1238 1836
rect -1218 1790 -1214 1836
rect -1194 1790 -1190 1836
rect -1170 1790 -1166 1836
rect -1146 1790 -1142 1836
rect -1122 1790 -1118 1836
rect -1098 1790 -1094 1836
rect -1074 1790 -1070 1836
rect -1050 1790 -1046 1836
rect -1026 1790 -1022 1836
rect -1002 1790 -998 1836
rect -978 1790 -974 1836
rect -954 1790 -950 1836
rect -930 1790 -926 1836
rect -906 1790 -902 1836
rect -882 1790 -878 1836
rect -858 1790 -854 1836
rect -834 1790 -830 1836
rect -810 1790 -806 1836
rect -786 1790 -782 1836
rect -762 1790 -758 1836
rect -738 1790 -734 1836
rect -714 1790 -710 1836
rect -690 1790 -686 1836
rect -666 1790 -662 1836
rect -642 1790 -638 1836
rect -618 1790 -614 1836
rect -594 1790 -590 1836
rect -570 1790 -566 1836
rect -546 1790 -542 1836
rect -522 1790 -518 1836
rect -498 1790 -494 1836
rect -474 1790 -470 1836
rect -450 1790 -446 1836
rect -426 1790 -422 1836
rect -402 1790 -398 1836
rect -378 1790 -374 1836
rect -354 1790 -350 1836
rect -330 1790 -326 1836
rect -306 1790 -302 1836
rect -293 1829 -288 1836
rect -282 1829 -278 1836
rect -283 1815 -278 1829
rect -293 1814 -259 1815
rect -258 1814 -254 1860
rect -234 1814 -230 1860
rect -210 1814 -206 1860
rect -186 1814 -182 1860
rect -162 1814 -158 1860
rect -138 1814 -134 1860
rect -114 1814 -110 1860
rect -90 1814 -86 1860
rect -66 1814 -62 1860
rect -42 1814 -38 1860
rect -18 1814 -14 1860
rect 6 1814 10 1860
rect 30 1814 34 1860
rect 54 1814 58 1860
rect 78 1814 82 1860
rect 102 1814 106 1860
rect 126 1814 130 1860
rect 150 1814 154 1860
rect 174 1814 178 1860
rect 198 1814 202 1860
rect 222 1814 226 1860
rect 246 1814 250 1860
rect 270 1814 274 1860
rect 294 1814 298 1860
rect 318 1814 322 1860
rect 342 1814 346 1860
rect 366 1814 370 1860
rect 390 1814 394 1860
rect 414 1814 418 1860
rect 438 1814 442 1860
rect 462 1814 466 1860
rect 486 1814 490 1860
rect 499 1838 533 1839
rect 534 1838 538 1860
rect 558 1838 562 1860
rect 582 1838 586 1860
rect 606 1838 610 1860
rect 630 1838 634 1860
rect 654 1838 658 1860
rect 678 1838 682 1860
rect 702 1838 706 1860
rect 726 1838 730 1860
rect 750 1838 754 1860
rect 774 1838 778 1860
rect 798 1838 802 1860
rect 822 1838 826 1860
rect 846 1838 850 1860
rect 870 1838 874 1860
rect 894 1838 898 1860
rect 918 1838 922 1860
rect 942 1838 946 1860
rect 955 1853 960 1860
rect 966 1853 970 1860
rect 965 1839 970 1853
rect 990 1838 994 1932
rect 1003 1901 1008 1911
rect 1014 1901 1018 1932
rect 1013 1887 1018 1901
rect 1003 1886 1037 1887
rect 1038 1886 1042 1932
rect 1062 1886 1066 1932
rect 1086 1886 1090 1932
rect 1110 1886 1114 1932
rect 1134 1886 1138 1932
rect 1158 1886 1162 1932
rect 1182 1886 1186 1932
rect 1206 1886 1210 1932
rect 1230 1886 1234 1932
rect 1254 1886 1258 1932
rect 1278 1886 1282 1932
rect 1302 1886 1306 1932
rect 1326 1886 1330 1932
rect 1350 1886 1354 1932
rect 1374 1886 1378 1932
rect 1398 1886 1402 1932
rect 1422 1886 1426 1932
rect 1446 1886 1450 1932
rect 1470 1886 1474 1932
rect 1494 1886 1498 1932
rect 1518 1886 1522 1932
rect 1531 1925 1536 1932
rect 1541 1911 1546 1925
rect 1542 1886 1546 1911
rect 1566 1907 1570 1956
rect 1003 1884 1563 1886
rect 1003 1877 1008 1884
rect 1013 1863 1018 1877
rect 1014 1838 1018 1863
rect 1038 1838 1042 1884
rect 1062 1838 1066 1884
rect 1086 1838 1090 1884
rect 1110 1838 1114 1884
rect 1134 1838 1138 1884
rect 1158 1838 1162 1884
rect 1182 1838 1186 1884
rect 1206 1838 1210 1884
rect 1230 1838 1234 1884
rect 1254 1838 1258 1884
rect 1278 1838 1282 1884
rect 1302 1838 1306 1884
rect 1326 1838 1330 1884
rect 1350 1838 1354 1884
rect 1374 1838 1378 1884
rect 1398 1838 1402 1884
rect 1422 1838 1426 1884
rect 1446 1838 1450 1884
rect 1470 1838 1474 1884
rect 1494 1838 1498 1884
rect 1518 1838 1522 1884
rect 1542 1838 1546 1884
rect 1549 1883 1563 1884
rect 1566 1883 1573 1907
rect 499 1836 1563 1838
rect 499 1829 504 1836
rect 509 1815 514 1829
rect 510 1814 514 1815
rect 534 1814 538 1836
rect 558 1814 562 1836
rect 582 1814 586 1836
rect 606 1814 610 1836
rect 630 1814 634 1836
rect 654 1814 658 1836
rect 678 1814 682 1836
rect 702 1814 706 1836
rect 726 1814 730 1836
rect 750 1814 754 1836
rect 774 1814 778 1836
rect 798 1814 802 1836
rect 822 1814 826 1836
rect 846 1814 850 1836
rect 870 1814 874 1836
rect 894 1814 898 1836
rect 918 1814 922 1836
rect 942 1814 946 1836
rect 990 1814 994 1836
rect 1014 1814 1018 1836
rect 1038 1835 1042 1836
rect -293 1812 1035 1814
rect -293 1805 -288 1812
rect -283 1791 -278 1805
rect -282 1790 -278 1791
rect -258 1790 -254 1812
rect -234 1790 -230 1812
rect -210 1790 -206 1812
rect -186 1790 -182 1812
rect -162 1790 -158 1812
rect -138 1790 -134 1812
rect -114 1790 -110 1812
rect -90 1790 -86 1812
rect -66 1790 -62 1812
rect -42 1790 -38 1812
rect -18 1790 -14 1812
rect 6 1790 10 1812
rect 30 1790 34 1812
rect 54 1790 58 1812
rect 78 1790 82 1812
rect 102 1790 106 1812
rect 126 1790 130 1812
rect 150 1790 154 1812
rect 174 1790 178 1812
rect 198 1790 202 1812
rect 222 1790 226 1812
rect 246 1790 250 1812
rect 270 1790 274 1812
rect 294 1790 298 1812
rect 318 1790 322 1812
rect 342 1790 346 1812
rect 366 1790 370 1812
rect 390 1790 394 1812
rect 414 1790 418 1812
rect 438 1790 442 1812
rect 462 1790 466 1812
rect 486 1790 490 1812
rect 510 1790 514 1812
rect 534 1811 538 1812
rect -2393 1788 531 1790
rect -2371 1766 -2366 1788
rect -2348 1766 -2343 1788
rect -2325 1780 -2317 1788
rect -2325 1766 -2320 1780
rect -2309 1768 -2301 1780
rect -2092 1771 -2062 1776
rect -2000 1768 -1992 1788
rect -2317 1766 -2309 1768
rect -2000 1766 -1983 1768
rect -1906 1766 -1904 1788
rect -1806 1780 -1680 1786
rect -1671 1780 -1663 1788
rect -1854 1771 -1806 1776
rect -1846 1766 -1806 1769
rect -1655 1768 -1647 1780
rect -1663 1766 -1655 1768
rect -1642 1766 -1637 1788
rect -1619 1766 -1614 1788
rect -1530 1766 -1526 1788
rect -1506 1766 -1502 1788
rect -1482 1766 -1478 1788
rect -1458 1766 -1454 1788
rect -1434 1766 -1430 1788
rect -1410 1766 -1406 1788
rect -1386 1766 -1382 1788
rect -1362 1766 -1358 1788
rect -1338 1766 -1334 1788
rect -1314 1766 -1310 1788
rect -1290 1766 -1286 1788
rect -1266 1766 -1262 1788
rect -1242 1766 -1238 1788
rect -1218 1766 -1214 1788
rect -1194 1766 -1190 1788
rect -1170 1766 -1166 1788
rect -1146 1766 -1142 1788
rect -1122 1766 -1118 1788
rect -1098 1766 -1094 1788
rect -1074 1766 -1070 1788
rect -1050 1766 -1046 1788
rect -1026 1766 -1022 1788
rect -1002 1766 -998 1788
rect -978 1766 -974 1788
rect -954 1766 -950 1788
rect -930 1766 -926 1788
rect -906 1767 -902 1788
rect -917 1766 -883 1767
rect -2393 1764 -883 1766
rect -2371 1742 -2366 1764
rect -2348 1742 -2343 1764
rect -2325 1752 -2317 1764
rect -2071 1760 -2062 1764
rect -2013 1762 -1983 1764
rect -2000 1761 -1983 1762
rect -2325 1742 -2320 1752
rect -2309 1742 -2301 1752
rect -2100 1751 -2092 1758
rect -2064 1756 -2062 1759
rect -2061 1751 -2059 1756
rect -2071 1746 -2062 1751
rect -2071 1744 -2026 1746
rect -2066 1742 -2012 1744
rect -2000 1742 -1992 1761
rect -1906 1759 -1904 1764
rect -1846 1760 -1806 1764
rect -1846 1753 -1798 1758
rect -1806 1751 -1798 1753
rect -1671 1752 -1663 1764
rect -1854 1749 -1846 1751
rect -1854 1744 -1806 1749
rect -1864 1742 -1796 1743
rect -1655 1742 -1647 1752
rect -1642 1742 -1637 1764
rect -1619 1742 -1614 1764
rect -1530 1742 -1526 1764
rect -1506 1742 -1502 1764
rect -1482 1742 -1478 1764
rect -1458 1742 -1454 1764
rect -1434 1742 -1430 1764
rect -1410 1742 -1406 1764
rect -1386 1742 -1382 1764
rect -1362 1742 -1358 1764
rect -1338 1742 -1334 1764
rect -1314 1742 -1310 1764
rect -1290 1742 -1286 1764
rect -1266 1742 -1262 1764
rect -1242 1742 -1238 1764
rect -1218 1742 -1214 1764
rect -1194 1742 -1190 1764
rect -1170 1742 -1166 1764
rect -1146 1742 -1142 1764
rect -1122 1742 -1118 1764
rect -1098 1742 -1094 1764
rect -1074 1742 -1070 1764
rect -1050 1742 -1046 1764
rect -1026 1742 -1022 1764
rect -1002 1742 -998 1764
rect -978 1742 -974 1764
rect -954 1742 -950 1764
rect -930 1742 -926 1764
rect -917 1757 -912 1764
rect -906 1757 -902 1764
rect -907 1743 -902 1757
rect -906 1742 -902 1743
rect -882 1742 -878 1788
rect -858 1742 -854 1788
rect -834 1742 -830 1788
rect -810 1742 -806 1788
rect -786 1742 -782 1788
rect -762 1742 -758 1788
rect -738 1742 -734 1788
rect -714 1742 -710 1788
rect -690 1742 -686 1788
rect -666 1742 -662 1788
rect -642 1742 -638 1788
rect -618 1742 -614 1788
rect -594 1742 -590 1788
rect -570 1742 -566 1788
rect -546 1742 -542 1788
rect -522 1742 -518 1788
rect -498 1742 -494 1788
rect -474 1742 -470 1788
rect -450 1742 -446 1788
rect -426 1743 -422 1788
rect -437 1742 -403 1743
rect -2393 1740 -403 1742
rect -2371 1694 -2366 1740
rect -2348 1694 -2343 1740
rect -2325 1736 -2320 1740
rect -2317 1736 -2309 1740
rect -2325 1724 -2317 1736
rect -2066 1735 -2062 1740
rect -2147 1732 -2134 1734
rect -2292 1726 -2071 1732
rect -2325 1694 -2320 1724
rect -2092 1710 -2062 1712
rect -2094 1706 -2062 1710
rect -2000 1694 -1992 1740
rect -1846 1733 -1806 1740
rect -1663 1736 -1655 1740
rect -1846 1726 -1680 1732
rect -1671 1724 -1663 1736
rect -1854 1710 -1806 1712
rect -1854 1706 -1680 1710
rect -1979 1694 -1945 1696
rect -1642 1694 -1637 1740
rect -1619 1694 -1614 1740
rect -1530 1694 -1526 1740
rect -1506 1694 -1502 1740
rect -1482 1694 -1478 1740
rect -1458 1694 -1454 1740
rect -1434 1694 -1430 1740
rect -1410 1694 -1406 1740
rect -1386 1694 -1382 1740
rect -1362 1694 -1358 1740
rect -1338 1694 -1334 1740
rect -1314 1694 -1310 1740
rect -1290 1694 -1286 1740
rect -1266 1694 -1262 1740
rect -1242 1694 -1238 1740
rect -1218 1694 -1214 1740
rect -1194 1694 -1190 1740
rect -1170 1694 -1166 1740
rect -1146 1694 -1142 1740
rect -1122 1694 -1118 1740
rect -1098 1694 -1094 1740
rect -1074 1694 -1070 1740
rect -1050 1694 -1046 1740
rect -1026 1694 -1022 1740
rect -1002 1694 -998 1740
rect -978 1694 -974 1740
rect -954 1694 -950 1740
rect -930 1694 -926 1740
rect -906 1694 -902 1740
rect -882 1694 -878 1740
rect -858 1694 -854 1740
rect -834 1694 -830 1740
rect -810 1694 -806 1740
rect -786 1694 -782 1740
rect -762 1694 -758 1740
rect -738 1694 -734 1740
rect -714 1694 -710 1740
rect -690 1694 -686 1740
rect -666 1694 -662 1740
rect -642 1694 -638 1740
rect -618 1694 -614 1740
rect -594 1694 -590 1740
rect -570 1694 -566 1740
rect -546 1694 -542 1740
rect -522 1694 -518 1740
rect -498 1694 -494 1740
rect -474 1694 -470 1740
rect -450 1694 -446 1740
rect -437 1733 -432 1740
rect -426 1733 -422 1740
rect -427 1719 -422 1733
rect -426 1694 -422 1719
rect -402 1694 -398 1788
rect -378 1694 -374 1788
rect -354 1694 -350 1788
rect -330 1694 -326 1788
rect -306 1694 -302 1788
rect -282 1694 -278 1788
rect -258 1763 -254 1788
rect -258 1715 -251 1763
rect -258 1694 -254 1715
rect -234 1694 -230 1788
rect -210 1694 -206 1788
rect -186 1694 -182 1788
rect -162 1694 -158 1788
rect -138 1694 -134 1788
rect -114 1694 -110 1788
rect -90 1694 -86 1788
rect -66 1694 -62 1788
rect -42 1694 -38 1788
rect -18 1694 -14 1788
rect 6 1694 10 1788
rect 30 1694 34 1788
rect 54 1694 58 1788
rect 78 1694 82 1788
rect 102 1694 106 1788
rect 126 1694 130 1788
rect 150 1694 154 1788
rect 174 1694 178 1788
rect 198 1694 202 1788
rect 222 1694 226 1788
rect 246 1694 250 1788
rect 270 1694 274 1788
rect 294 1694 298 1788
rect 318 1694 322 1788
rect 342 1694 346 1788
rect 366 1694 370 1788
rect 390 1694 394 1788
rect 414 1694 418 1788
rect 438 1694 442 1788
rect 462 1694 466 1788
rect 486 1694 490 1788
rect 510 1694 514 1788
rect 517 1787 531 1788
rect 534 1787 541 1811
rect 534 1739 541 1763
rect 534 1694 538 1739
rect 558 1694 562 1812
rect 582 1694 586 1812
rect 606 1694 610 1812
rect 630 1694 634 1812
rect 654 1694 658 1812
rect 678 1694 682 1812
rect 702 1694 706 1812
rect 726 1694 730 1812
rect 750 1694 754 1812
rect 774 1694 778 1812
rect 798 1694 802 1812
rect 822 1694 826 1812
rect 846 1694 850 1812
rect 870 1694 874 1812
rect 894 1694 898 1812
rect 918 1694 922 1812
rect 942 1694 946 1812
rect 955 1781 960 1791
rect 990 1787 994 1812
rect 965 1767 970 1781
rect 979 1777 987 1781
rect 973 1767 979 1777
rect 966 1694 970 1767
rect 990 1763 997 1787
rect -2393 1692 987 1694
rect -2371 1646 -2366 1692
rect -2348 1646 -2343 1692
rect -2325 1646 -2320 1692
rect -2080 1691 -1906 1692
rect -2080 1690 -2036 1691
rect -2080 1684 -2054 1690
rect -2309 1676 -2301 1682
rect -2317 1666 -2309 1676
rect -2070 1675 -2040 1682
rect -2054 1667 -2040 1670
rect -2000 1665 -1992 1691
rect -1920 1690 -1906 1691
rect -1850 1684 -1846 1692
rect -1840 1684 -1792 1692
rect -1969 1672 -1966 1681
rect -1850 1677 -1802 1682
rect -1906 1675 -1802 1677
rect -1655 1676 -1647 1682
rect -1906 1674 -1850 1675
rect -1846 1667 -1802 1673
rect -1663 1666 -1655 1676
rect -1860 1665 -1798 1666
rect -2078 1658 -2070 1665
rect -2309 1648 -2301 1654
rect -2317 1646 -2309 1648
rect -2154 1646 -2145 1656
rect -2044 1655 -2040 1660
rect -2028 1658 -1945 1665
rect -1929 1658 -1794 1665
rect -2070 1648 -2040 1655
rect -2044 1646 -2028 1648
rect -2000 1646 -1992 1658
rect -1860 1657 -1798 1658
rect -1850 1648 -1802 1655
rect -1655 1648 -1647 1654
rect -1978 1646 -1942 1647
rect -1663 1646 -1655 1648
rect -1642 1646 -1637 1692
rect -1619 1646 -1614 1692
rect -1530 1646 -1526 1692
rect -1506 1646 -1502 1692
rect -1482 1646 -1478 1692
rect -1458 1646 -1454 1692
rect -1434 1646 -1430 1692
rect -1410 1646 -1406 1692
rect -1386 1646 -1382 1692
rect -1362 1646 -1358 1692
rect -1338 1646 -1334 1692
rect -1314 1646 -1310 1692
rect -1290 1646 -1286 1692
rect -1266 1646 -1262 1692
rect -1242 1646 -1238 1692
rect -1218 1646 -1214 1692
rect -1194 1646 -1190 1692
rect -1170 1646 -1166 1692
rect -1146 1646 -1142 1692
rect -1122 1646 -1118 1692
rect -1098 1646 -1094 1692
rect -1074 1646 -1070 1692
rect -1050 1646 -1046 1692
rect -1026 1646 -1022 1692
rect -1002 1646 -998 1692
rect -978 1646 -974 1692
rect -954 1646 -950 1692
rect -930 1646 -926 1692
rect -906 1646 -902 1692
rect -882 1691 -878 1692
rect -882 1667 -875 1691
rect -882 1646 -878 1667
rect -858 1646 -854 1692
rect -834 1646 -830 1692
rect -810 1646 -806 1692
rect -786 1646 -782 1692
rect -762 1646 -758 1692
rect -738 1646 -734 1692
rect -714 1646 -710 1692
rect -690 1646 -686 1692
rect -666 1646 -662 1692
rect -642 1646 -638 1692
rect -618 1646 -614 1692
rect -594 1646 -590 1692
rect -570 1646 -566 1692
rect -546 1646 -542 1692
rect -522 1646 -518 1692
rect -498 1646 -494 1692
rect -474 1646 -470 1692
rect -450 1646 -446 1692
rect -426 1646 -422 1692
rect -402 1667 -398 1692
rect -2393 1644 -405 1646
rect -2371 1550 -2366 1644
rect -2348 1550 -2343 1644
rect -2325 1606 -2320 1644
rect -2317 1638 -2309 1644
rect -2145 1640 -2138 1644
rect -2070 1640 -2054 1644
rect -2078 1631 -2054 1638
rect -2062 1606 -2032 1607
rect -2000 1606 -1992 1644
rect -1846 1640 -1802 1644
rect -1846 1630 -1792 1639
rect -1663 1638 -1655 1644
rect -1942 1608 -1937 1620
rect -1850 1617 -1822 1618
rect -1850 1613 -1802 1617
rect -2325 1598 -2317 1606
rect -2062 1604 -1961 1606
rect -2325 1578 -2320 1598
rect -2317 1590 -2309 1598
rect -2062 1591 -2040 1602
rect -2032 1597 -1961 1604
rect -1947 1598 -1942 1606
rect -1842 1604 -1794 1607
rect -2070 1586 -2022 1590
rect -2325 1564 -2317 1578
rect -2072 1570 -2032 1571
rect -2102 1564 -2032 1570
rect -2325 1550 -2320 1564
rect -2317 1562 -2309 1564
rect -2309 1550 -2301 1562
rect -2070 1555 -2062 1560
rect -2000 1550 -1992 1597
rect -1942 1596 -1937 1598
rect -1932 1588 -1927 1596
rect -1912 1593 -1896 1599
rect -1842 1591 -1802 1602
rect -1671 1598 -1663 1606
rect -1663 1590 -1655 1598
rect -1850 1586 -1680 1590
rect -1924 1572 -1921 1574
rect -1806 1564 -1680 1570
rect -1671 1564 -1663 1578
rect -1663 1562 -1655 1564
rect -1854 1555 -1806 1560
rect -1974 1550 -1964 1551
rect -1960 1550 -1944 1552
rect -1842 1550 -1806 1553
rect -1655 1550 -1647 1562
rect -1642 1550 -1637 1644
rect -1619 1550 -1614 1644
rect -1530 1550 -1526 1644
rect -1506 1550 -1502 1644
rect -1482 1550 -1478 1644
rect -1458 1550 -1454 1644
rect -1434 1550 -1430 1644
rect -1410 1550 -1406 1644
rect -1386 1550 -1382 1644
rect -1362 1550 -1358 1644
rect -1338 1550 -1334 1644
rect -1314 1550 -1310 1644
rect -1290 1550 -1286 1644
rect -1266 1550 -1262 1644
rect -1242 1550 -1238 1644
rect -1218 1550 -1214 1644
rect -1194 1550 -1190 1644
rect -1170 1550 -1166 1644
rect -1146 1550 -1142 1644
rect -1122 1550 -1118 1644
rect -1098 1550 -1094 1644
rect -1074 1550 -1070 1644
rect -1050 1550 -1046 1644
rect -1026 1550 -1022 1644
rect -1002 1550 -998 1644
rect -978 1550 -974 1644
rect -954 1550 -950 1644
rect -930 1550 -926 1644
rect -906 1550 -902 1644
rect -882 1550 -878 1644
rect -858 1550 -854 1644
rect -834 1550 -830 1644
rect -810 1550 -806 1644
rect -786 1550 -782 1644
rect -762 1550 -758 1644
rect -738 1550 -734 1644
rect -714 1550 -710 1644
rect -690 1550 -686 1644
rect -666 1550 -662 1644
rect -642 1550 -638 1644
rect -618 1550 -614 1644
rect -594 1550 -590 1644
rect -570 1550 -566 1644
rect -557 1613 -552 1623
rect -546 1613 -542 1644
rect -547 1599 -542 1613
rect -557 1598 -523 1599
rect -522 1598 -518 1644
rect -498 1598 -494 1644
rect -474 1598 -470 1644
rect -450 1598 -446 1644
rect -426 1598 -422 1644
rect -419 1643 -405 1644
rect -402 1643 -395 1667
rect -402 1598 -398 1643
rect -378 1598 -374 1692
rect -354 1598 -350 1692
rect -330 1598 -326 1692
rect -306 1598 -302 1692
rect -282 1598 -278 1692
rect -258 1598 -254 1692
rect -234 1598 -230 1692
rect -210 1598 -206 1692
rect -186 1598 -182 1692
rect -162 1598 -158 1692
rect -138 1598 -134 1692
rect -114 1598 -110 1692
rect -90 1598 -86 1692
rect -66 1598 -62 1692
rect -42 1598 -38 1692
rect -18 1598 -14 1692
rect 6 1598 10 1692
rect 30 1598 34 1692
rect 54 1598 58 1692
rect 78 1598 82 1692
rect 102 1598 106 1692
rect 126 1598 130 1692
rect 150 1598 154 1692
rect 174 1598 178 1692
rect 198 1598 202 1692
rect 222 1598 226 1692
rect 246 1598 250 1692
rect 270 1598 274 1692
rect 294 1598 298 1692
rect 318 1598 322 1692
rect 342 1598 346 1692
rect 366 1598 370 1692
rect 390 1598 394 1692
rect 414 1598 418 1692
rect 438 1598 442 1692
rect 462 1598 466 1692
rect 486 1598 490 1692
rect 510 1598 514 1692
rect 534 1598 538 1692
rect 558 1598 562 1692
rect 582 1598 586 1692
rect 606 1598 610 1692
rect 630 1598 634 1692
rect 654 1598 658 1692
rect 678 1598 682 1692
rect 702 1598 706 1692
rect 726 1598 730 1692
rect 750 1598 754 1692
rect 774 1598 778 1692
rect 798 1598 802 1692
rect 822 1598 826 1692
rect 846 1598 850 1692
rect 870 1598 874 1692
rect 894 1598 898 1692
rect 918 1598 922 1692
rect 942 1598 946 1692
rect 966 1598 970 1692
rect 973 1691 987 1692
rect 990 1691 997 1715
rect 990 1598 994 1691
rect 1014 1598 1018 1812
rect 1021 1811 1035 1812
rect 1038 1787 1045 1835
rect 1038 1598 1042 1787
rect 1062 1598 1066 1836
rect 1086 1598 1090 1836
rect 1110 1598 1114 1836
rect 1134 1598 1138 1836
rect 1158 1598 1162 1836
rect 1182 1598 1186 1836
rect 1206 1598 1210 1836
rect 1230 1598 1234 1836
rect 1254 1598 1258 1836
rect 1278 1598 1282 1836
rect 1302 1598 1306 1836
rect 1326 1598 1330 1836
rect 1350 1598 1354 1836
rect 1374 1598 1378 1836
rect 1398 1598 1402 1836
rect 1422 1598 1426 1836
rect 1446 1598 1450 1836
rect 1470 1598 1474 1836
rect 1494 1598 1498 1836
rect 1518 1598 1522 1836
rect 1542 1598 1546 1836
rect 1549 1835 1563 1836
rect 1566 1835 1573 1859
rect 1566 1598 1570 1835
rect 1590 1598 1594 1956
rect 1603 1637 1608 1647
rect 1614 1637 1618 1956
rect 1613 1623 1618 1637
rect 1603 1613 1608 1623
rect 1613 1599 1618 1613
rect 1614 1598 1618 1599
rect 1638 1598 1642 1956
rect 1662 1598 1666 1956
rect 1686 1598 1690 1956
rect 1710 1598 1714 1956
rect 1734 1598 1738 1956
rect 1758 1598 1762 1956
rect 1782 1598 1786 1956
rect 1806 1598 1810 1956
rect 1830 1599 1834 1956
rect 1843 1805 1848 1815
rect 1854 1805 1858 1956
rect 1867 1829 1872 1839
rect 1878 1829 1882 1956
rect 1891 1877 1896 1887
rect 1902 1877 1906 1956
rect 1915 1949 1920 1956
rect 1926 1949 1930 1956
rect 1933 1955 1947 1956
rect 1925 1935 1930 1949
rect 1939 1945 1947 1949
rect 1933 1935 1939 1945
rect 1901 1863 1906 1877
rect 1877 1815 1882 1829
rect 1853 1791 1858 1805
rect 1843 1685 1848 1695
rect 1853 1671 1858 1685
rect 1843 1613 1848 1623
rect 1854 1613 1858 1671
rect 1853 1599 1858 1613
rect 1867 1609 1875 1613
rect 1861 1599 1867 1609
rect 1819 1598 1853 1599
rect -557 1596 1853 1598
rect -557 1589 -552 1596
rect -547 1575 -542 1589
rect -546 1550 -542 1575
rect -522 1550 -518 1596
rect -498 1550 -494 1596
rect -474 1550 -470 1596
rect -450 1550 -446 1596
rect -426 1550 -422 1596
rect -402 1550 -398 1596
rect -378 1550 -374 1596
rect -354 1550 -350 1596
rect -330 1550 -326 1596
rect -306 1550 -302 1596
rect -282 1550 -278 1596
rect -258 1550 -254 1596
rect -234 1550 -230 1596
rect -210 1550 -206 1596
rect -186 1550 -182 1596
rect -162 1550 -158 1596
rect -138 1550 -134 1596
rect -114 1550 -110 1596
rect -90 1550 -86 1596
rect -66 1550 -62 1596
rect -42 1550 -38 1596
rect -18 1550 -14 1596
rect 6 1550 10 1596
rect 30 1550 34 1596
rect 54 1550 58 1596
rect 78 1550 82 1596
rect 102 1550 106 1596
rect 126 1550 130 1596
rect 150 1550 154 1596
rect 174 1550 178 1596
rect 198 1550 202 1596
rect 222 1550 226 1596
rect 246 1550 250 1596
rect 270 1550 274 1596
rect 294 1550 298 1596
rect 318 1551 322 1596
rect 307 1550 341 1551
rect -2393 1548 341 1550
rect -2371 1526 -2366 1548
rect -2348 1526 -2343 1548
rect -2325 1536 -2317 1548
rect -2325 1526 -2320 1536
rect -2317 1534 -2309 1536
rect -2062 1535 -2032 1542
rect -2309 1526 -2301 1534
rect -2070 1528 -2062 1535
rect -2000 1530 -1992 1548
rect -1974 1546 -1944 1548
rect -1960 1545 -1944 1546
rect -1842 1544 -1806 1548
rect -1842 1537 -1798 1542
rect -1806 1535 -1798 1537
rect -1671 1536 -1663 1548
rect -1854 1533 -1842 1535
rect -1663 1534 -1655 1536
rect -2062 1526 -2036 1528
rect -2393 1524 -2036 1526
rect -2032 1526 -2012 1528
rect -2004 1526 -1974 1530
rect -1854 1528 -1806 1533
rect -1864 1526 -1796 1527
rect -1655 1526 -1647 1534
rect -1642 1526 -1637 1548
rect -1619 1526 -1614 1548
rect -1530 1526 -1526 1548
rect -1506 1526 -1502 1548
rect -1482 1526 -1478 1548
rect -1458 1526 -1454 1548
rect -1434 1526 -1430 1548
rect -1410 1526 -1406 1548
rect -1386 1526 -1382 1548
rect -1362 1526 -1358 1548
rect -1338 1526 -1334 1548
rect -1314 1526 -1310 1548
rect -1290 1526 -1286 1548
rect -1266 1526 -1262 1548
rect -1242 1526 -1238 1548
rect -1218 1526 -1214 1548
rect -1194 1526 -1190 1548
rect -1170 1526 -1166 1548
rect -1146 1526 -1142 1548
rect -1122 1526 -1118 1548
rect -1098 1526 -1094 1548
rect -1074 1526 -1070 1548
rect -1050 1526 -1046 1548
rect -1026 1526 -1022 1548
rect -1002 1526 -998 1548
rect -978 1526 -974 1548
rect -954 1526 -950 1548
rect -930 1526 -926 1548
rect -906 1526 -902 1548
rect -882 1526 -878 1548
rect -858 1526 -854 1548
rect -834 1526 -830 1548
rect -810 1526 -806 1548
rect -786 1526 -782 1548
rect -762 1526 -758 1548
rect -738 1526 -734 1548
rect -714 1526 -710 1548
rect -690 1526 -686 1548
rect -666 1526 -662 1548
rect -642 1526 -638 1548
rect -618 1526 -614 1548
rect -594 1526 -590 1548
rect -570 1526 -566 1548
rect -546 1526 -542 1548
rect -522 1547 -518 1548
rect -2032 1524 -525 1526
rect -2371 1478 -2366 1524
rect -2348 1478 -2343 1524
rect -2325 1520 -2320 1524
rect -2309 1522 -2301 1524
rect -2317 1520 -2309 1522
rect -2325 1508 -2317 1520
rect -2052 1518 -2036 1520
rect -2052 1516 -2032 1518
rect -2062 1510 -2032 1516
rect -2325 1488 -2320 1508
rect -2317 1506 -2309 1508
rect -2092 1494 -2062 1496
rect -2094 1490 -2062 1494
rect -2325 1478 -2317 1488
rect -2095 1480 -2084 1484
rect -2000 1481 -1992 1524
rect -1904 1517 -1874 1524
rect -1842 1517 -1806 1524
rect -1655 1522 -1647 1524
rect -1663 1520 -1655 1522
rect -1842 1510 -1680 1516
rect -1671 1508 -1663 1520
rect -1663 1506 -1655 1508
rect -1854 1494 -1806 1496
rect -1854 1490 -1680 1494
rect -2119 1478 -2069 1480
rect -2054 1478 -1892 1481
rect -1671 1478 -1663 1488
rect -1642 1478 -1637 1524
rect -1619 1478 -1614 1524
rect -1530 1478 -1526 1524
rect -1506 1478 -1502 1524
rect -1482 1478 -1478 1524
rect -1458 1478 -1454 1524
rect -1434 1478 -1430 1524
rect -1410 1478 -1406 1524
rect -1386 1478 -1382 1524
rect -1362 1478 -1358 1524
rect -1338 1478 -1334 1524
rect -1314 1478 -1310 1524
rect -1290 1478 -1286 1524
rect -1266 1478 -1262 1524
rect -1242 1478 -1238 1524
rect -1218 1478 -1214 1524
rect -1194 1478 -1190 1524
rect -1170 1478 -1166 1524
rect -1146 1478 -1142 1524
rect -1122 1478 -1118 1524
rect -1098 1478 -1094 1524
rect -1074 1478 -1070 1524
rect -1050 1478 -1046 1524
rect -1026 1478 -1022 1524
rect -1002 1478 -998 1524
rect -978 1478 -974 1524
rect -954 1478 -950 1524
rect -930 1478 -926 1524
rect -906 1478 -902 1524
rect -882 1478 -878 1524
rect -858 1478 -854 1524
rect -834 1478 -830 1524
rect -810 1478 -806 1524
rect -786 1478 -782 1524
rect -762 1478 -758 1524
rect -738 1478 -734 1524
rect -714 1478 -710 1524
rect -690 1478 -686 1524
rect -666 1478 -662 1524
rect -642 1478 -638 1524
rect -618 1478 -614 1524
rect -594 1478 -590 1524
rect -570 1478 -566 1524
rect -546 1478 -542 1524
rect -539 1523 -525 1524
rect -522 1499 -515 1547
rect -522 1478 -518 1499
rect -498 1478 -494 1548
rect -474 1478 -470 1548
rect -450 1478 -446 1548
rect -426 1478 -422 1548
rect -402 1478 -398 1548
rect -378 1478 -374 1548
rect -354 1478 -350 1548
rect -330 1478 -326 1548
rect -306 1478 -302 1548
rect -282 1478 -278 1548
rect -258 1478 -254 1548
rect -234 1478 -230 1548
rect -210 1478 -206 1548
rect -186 1478 -182 1548
rect -162 1478 -158 1548
rect -138 1478 -134 1548
rect -114 1478 -110 1548
rect -90 1478 -86 1548
rect -66 1478 -62 1548
rect -42 1478 -38 1548
rect -18 1478 -14 1548
rect 6 1478 10 1548
rect 30 1478 34 1548
rect 54 1478 58 1548
rect 78 1478 82 1548
rect 102 1478 106 1548
rect 126 1478 130 1548
rect 150 1478 154 1548
rect 163 1517 168 1527
rect 174 1517 178 1548
rect 173 1503 178 1517
rect 163 1502 197 1503
rect 198 1502 202 1548
rect 222 1502 226 1548
rect 246 1502 250 1548
rect 270 1502 274 1548
rect 294 1502 298 1548
rect 307 1541 312 1548
rect 318 1541 322 1548
rect 317 1527 322 1541
rect 307 1517 312 1527
rect 317 1503 322 1517
rect 318 1502 322 1503
rect 342 1502 346 1596
rect 366 1502 370 1596
rect 390 1502 394 1596
rect 414 1502 418 1596
rect 438 1502 442 1596
rect 462 1502 466 1596
rect 486 1502 490 1596
rect 510 1502 514 1596
rect 534 1502 538 1596
rect 558 1502 562 1596
rect 582 1502 586 1596
rect 606 1502 610 1596
rect 630 1502 634 1596
rect 654 1502 658 1596
rect 678 1502 682 1596
rect 702 1502 706 1596
rect 726 1502 730 1596
rect 750 1502 754 1596
rect 774 1502 778 1596
rect 798 1502 802 1596
rect 822 1502 826 1596
rect 846 1502 850 1596
rect 870 1502 874 1596
rect 894 1502 898 1596
rect 918 1502 922 1596
rect 942 1502 946 1596
rect 966 1502 970 1596
rect 990 1502 994 1596
rect 1014 1502 1018 1596
rect 1038 1502 1042 1596
rect 1062 1502 1066 1596
rect 1086 1502 1090 1596
rect 1110 1502 1114 1596
rect 1134 1502 1138 1596
rect 1158 1502 1162 1596
rect 1182 1502 1186 1596
rect 1206 1502 1210 1596
rect 1230 1502 1234 1596
rect 1254 1502 1258 1596
rect 1278 1502 1282 1596
rect 1302 1502 1306 1596
rect 1326 1502 1330 1596
rect 1350 1502 1354 1596
rect 1374 1502 1378 1596
rect 1398 1502 1402 1596
rect 1422 1502 1426 1596
rect 1446 1502 1450 1596
rect 1470 1502 1474 1596
rect 1494 1502 1498 1596
rect 1518 1502 1522 1596
rect 1542 1502 1546 1596
rect 1566 1502 1570 1596
rect 1590 1502 1594 1596
rect 1614 1502 1618 1596
rect 1638 1571 1642 1596
rect 1638 1526 1645 1571
rect 1662 1526 1666 1596
rect 1686 1526 1690 1596
rect 1710 1526 1714 1596
rect 1734 1526 1738 1596
rect 1758 1526 1762 1596
rect 1782 1526 1786 1596
rect 1806 1526 1810 1596
rect 1819 1589 1824 1596
rect 1830 1589 1834 1596
rect 1829 1575 1834 1589
rect 1819 1565 1824 1575
rect 1829 1551 1834 1565
rect 1830 1527 1834 1551
rect 1819 1526 1853 1527
rect 1621 1524 1853 1526
rect 1621 1523 1635 1524
rect 1638 1523 1645 1524
rect 1638 1502 1642 1523
rect 1662 1502 1666 1524
rect 1686 1502 1690 1524
rect 1710 1502 1714 1524
rect 1734 1502 1738 1524
rect 1758 1502 1762 1524
rect 1782 1502 1786 1524
rect 1806 1503 1810 1524
rect 1819 1517 1824 1524
rect 1830 1517 1834 1524
rect 1829 1503 1834 1517
rect 1843 1513 1851 1517
rect 1837 1503 1843 1513
rect 1795 1502 1829 1503
rect 163 1500 1829 1502
rect 163 1493 168 1500
rect 173 1479 178 1493
rect 174 1478 178 1479
rect 198 1478 202 1500
rect 222 1478 226 1500
rect 246 1478 250 1500
rect 270 1478 274 1500
rect 294 1478 298 1500
rect 318 1478 322 1500
rect 342 1478 346 1500
rect 366 1478 370 1500
rect 390 1478 394 1500
rect 414 1478 418 1500
rect 438 1478 442 1500
rect 462 1478 466 1500
rect 486 1478 490 1500
rect 510 1478 514 1500
rect 534 1478 538 1500
rect 558 1478 562 1500
rect 582 1478 586 1500
rect 606 1478 610 1500
rect 630 1478 634 1500
rect 654 1478 658 1500
rect 678 1478 682 1500
rect 702 1478 706 1500
rect 726 1478 730 1500
rect 750 1478 754 1500
rect 774 1478 778 1500
rect 798 1478 802 1500
rect 822 1478 826 1500
rect 846 1478 850 1500
rect 870 1478 874 1500
rect 894 1478 898 1500
rect 918 1478 922 1500
rect 942 1478 946 1500
rect 966 1478 970 1500
rect 990 1478 994 1500
rect 1014 1478 1018 1500
rect 1038 1478 1042 1500
rect 1062 1478 1066 1500
rect 1086 1478 1090 1500
rect 1110 1478 1114 1500
rect 1134 1478 1138 1500
rect 1158 1478 1162 1500
rect 1182 1478 1186 1500
rect 1206 1478 1210 1500
rect 1230 1478 1234 1500
rect 1254 1478 1258 1500
rect 1278 1478 1282 1500
rect 1302 1478 1306 1500
rect 1326 1478 1330 1500
rect 1350 1478 1354 1500
rect 1374 1478 1378 1500
rect 1398 1478 1402 1500
rect 1422 1478 1426 1500
rect 1446 1478 1450 1500
rect 1470 1478 1474 1500
rect 1494 1478 1498 1500
rect 1518 1478 1522 1500
rect 1542 1478 1546 1500
rect 1566 1478 1570 1500
rect 1590 1478 1594 1500
rect 1614 1478 1618 1500
rect 1638 1478 1642 1500
rect 1662 1478 1666 1500
rect 1686 1478 1690 1500
rect 1710 1478 1714 1500
rect 1734 1478 1738 1500
rect 1758 1478 1762 1500
rect 1782 1478 1786 1500
rect 1795 1493 1800 1500
rect 1806 1493 1810 1500
rect 1805 1479 1810 1493
rect 1795 1478 1829 1479
rect -2393 1476 1829 1478
rect -2371 1454 -2366 1476
rect -2348 1454 -2343 1476
rect -2325 1472 -2317 1476
rect -2325 1456 -2320 1472
rect -2309 1460 -2301 1472
rect -2095 1470 -2084 1476
rect -2054 1475 -1906 1476
rect -2054 1474 -2036 1475
rect -2084 1468 -2079 1470
rect -2317 1456 -2309 1460
rect -2092 1459 -2079 1466
rect -2000 1462 -1992 1475
rect -1920 1474 -1906 1475
rect -1671 1472 -1663 1476
rect -1846 1468 -1806 1470
rect -1854 1462 -1806 1466
rect -2054 1459 -1982 1462
rect -1966 1459 -1806 1462
rect -1655 1460 -1647 1472
rect -2003 1456 -1992 1459
rect -1904 1457 -1902 1459
rect -1854 1457 -1846 1459
rect -2325 1454 -2317 1456
rect -2033 1454 -1992 1456
rect -1854 1455 -1806 1457
rect -1663 1456 -1655 1460
rect -1864 1454 -1796 1455
rect -1671 1454 -1663 1456
rect -1642 1454 -1637 1476
rect -1619 1454 -1614 1476
rect -1530 1454 -1526 1476
rect -1506 1454 -1502 1476
rect -1482 1454 -1478 1476
rect -1458 1454 -1454 1476
rect -1434 1454 -1430 1476
rect -1410 1454 -1406 1476
rect -1386 1454 -1382 1476
rect -1362 1454 -1358 1476
rect -1338 1454 -1334 1476
rect -1314 1454 -1310 1476
rect -1290 1454 -1286 1476
rect -1266 1454 -1262 1476
rect -1242 1454 -1238 1476
rect -1218 1454 -1214 1476
rect -1194 1454 -1190 1476
rect -1170 1454 -1166 1476
rect -1146 1454 -1142 1476
rect -1122 1454 -1118 1476
rect -1098 1454 -1094 1476
rect -1074 1455 -1070 1476
rect -1085 1454 -1051 1455
rect -2393 1452 -1051 1454
rect -2371 1430 -2366 1452
rect -2348 1430 -2343 1452
rect -2325 1444 -2317 1452
rect -2079 1449 -2018 1452
rect -2003 1451 -1966 1452
rect -2000 1450 -1982 1451
rect -2000 1449 -1992 1450
rect -2084 1445 -2009 1449
rect -2028 1444 -2009 1445
rect -2000 1445 -1854 1449
rect -1846 1445 -1798 1452
rect -2325 1430 -2320 1444
rect -2309 1432 -2301 1444
rect -2028 1442 -2018 1444
rect -2092 1432 -2084 1439
rect -2023 1435 -2014 1442
rect -2000 1435 -1992 1445
rect -1671 1444 -1663 1452
rect -1846 1441 -1806 1443
rect -1854 1435 -1806 1439
rect -2054 1432 -1806 1435
rect -1655 1432 -1647 1444
rect -2317 1430 -2309 1432
rect -2054 1430 -2024 1432
rect -2000 1430 -1992 1432
rect -1663 1430 -1655 1432
rect -1642 1430 -1637 1452
rect -1619 1430 -1614 1452
rect -1589 1430 -1555 1431
rect -2393 1428 -2064 1430
rect -2060 1428 -1555 1430
rect -2371 1382 -2366 1428
rect -2348 1382 -2343 1428
rect -2325 1416 -2317 1428
rect -2060 1425 -2054 1428
rect -2084 1418 -2054 1425
rect -2050 1422 -2044 1424
rect -2325 1396 -2320 1416
rect -2064 1414 -2054 1418
rect -2325 1388 -2317 1396
rect -2101 1391 -2071 1394
rect -2325 1382 -2320 1388
rect -2317 1382 -2309 1388
rect -2000 1386 -1992 1428
rect -1846 1427 -1806 1428
rect -1846 1418 -1798 1425
rect -1671 1416 -1663 1428
rect -1846 1414 -1806 1416
rect -1854 1400 -1680 1404
rect -1846 1391 -1798 1394
rect -2079 1385 -2043 1386
rect -2007 1385 -1991 1386
rect -2079 1384 -2071 1385
rect -2079 1382 -2029 1384
rect -2011 1382 -1991 1385
rect -1846 1383 -1806 1389
rect -1671 1388 -1663 1396
rect -1864 1382 -1796 1383
rect -1663 1382 -1655 1388
rect -1642 1382 -1637 1428
rect -1619 1382 -1614 1428
rect -1589 1382 -1531 1383
rect -1530 1382 -1526 1452
rect -1506 1382 -1502 1452
rect -1482 1382 -1478 1452
rect -1458 1382 -1454 1452
rect -1434 1382 -1430 1452
rect -1410 1382 -1406 1452
rect -1386 1382 -1382 1452
rect -1362 1382 -1358 1452
rect -1338 1382 -1334 1452
rect -1314 1382 -1310 1452
rect -1290 1382 -1286 1452
rect -1266 1382 -1262 1452
rect -1242 1382 -1238 1452
rect -1218 1382 -1214 1452
rect -1194 1382 -1190 1452
rect -1170 1382 -1166 1452
rect -1146 1382 -1142 1452
rect -1122 1382 -1118 1452
rect -1098 1382 -1094 1452
rect -1085 1445 -1080 1452
rect -1074 1445 -1070 1452
rect -1075 1431 -1070 1445
rect -1085 1430 -1051 1431
rect -1050 1430 -1046 1476
rect -1026 1430 -1022 1476
rect -1002 1430 -998 1476
rect -978 1430 -974 1476
rect -954 1430 -950 1476
rect -930 1430 -926 1476
rect -906 1430 -902 1476
rect -882 1430 -878 1476
rect -858 1430 -854 1476
rect -834 1430 -830 1476
rect -810 1430 -806 1476
rect -786 1430 -782 1476
rect -762 1430 -758 1476
rect -738 1430 -734 1476
rect -714 1430 -710 1476
rect -690 1430 -686 1476
rect -666 1430 -662 1476
rect -642 1430 -638 1476
rect -618 1430 -614 1476
rect -594 1430 -590 1476
rect -570 1430 -566 1476
rect -546 1430 -542 1476
rect -522 1430 -518 1476
rect -498 1430 -494 1476
rect -474 1430 -470 1476
rect -450 1430 -446 1476
rect -426 1430 -422 1476
rect -402 1430 -398 1476
rect -378 1430 -374 1476
rect -354 1430 -350 1476
rect -330 1430 -326 1476
rect -306 1430 -302 1476
rect -282 1430 -278 1476
rect -258 1430 -254 1476
rect -234 1430 -230 1476
rect -210 1430 -206 1476
rect -186 1430 -182 1476
rect -162 1430 -158 1476
rect -138 1430 -134 1476
rect -114 1430 -110 1476
rect -90 1430 -86 1476
rect -66 1430 -62 1476
rect -42 1430 -38 1476
rect -18 1430 -14 1476
rect 6 1430 10 1476
rect 30 1430 34 1476
rect 54 1430 58 1476
rect 78 1430 82 1476
rect 102 1430 106 1476
rect 126 1430 130 1476
rect 150 1430 154 1476
rect 174 1430 178 1476
rect 198 1451 202 1476
rect -1085 1428 195 1430
rect -1085 1421 -1080 1428
rect -1075 1407 -1070 1421
rect -1074 1382 -1070 1407
rect -1050 1382 -1046 1428
rect -1026 1382 -1022 1428
rect -1002 1382 -998 1428
rect -978 1382 -974 1428
rect -954 1382 -950 1428
rect -930 1382 -926 1428
rect -906 1382 -902 1428
rect -882 1382 -878 1428
rect -858 1382 -854 1428
rect -834 1382 -830 1428
rect -810 1382 -806 1428
rect -786 1382 -782 1428
rect -762 1382 -758 1428
rect -738 1382 -734 1428
rect -714 1382 -710 1428
rect -690 1382 -686 1428
rect -666 1382 -662 1428
rect -642 1382 -638 1428
rect -618 1382 -614 1428
rect -594 1382 -590 1428
rect -570 1382 -566 1428
rect -546 1382 -542 1428
rect -522 1382 -518 1428
rect -498 1382 -494 1428
rect -474 1382 -470 1428
rect -450 1382 -446 1428
rect -426 1382 -422 1428
rect -402 1382 -398 1428
rect -378 1382 -374 1428
rect -354 1382 -350 1428
rect -330 1382 -326 1428
rect -306 1382 -302 1428
rect -282 1382 -278 1428
rect -258 1382 -254 1428
rect -245 1397 -240 1407
rect -234 1397 -230 1428
rect -235 1383 -230 1397
rect -210 1382 -206 1428
rect -186 1382 -182 1428
rect -162 1382 -158 1428
rect -138 1382 -134 1428
rect -114 1382 -110 1428
rect -90 1382 -86 1428
rect -66 1382 -62 1428
rect -42 1382 -38 1428
rect -18 1382 -14 1428
rect 6 1383 10 1428
rect -5 1382 29 1383
rect -2393 1380 29 1382
rect -2371 1334 -2366 1380
rect -2348 1334 -2343 1380
rect -2325 1368 -2320 1380
rect -2079 1378 -2071 1380
rect -2072 1376 -2071 1378
rect -2109 1371 -2101 1376
rect -2101 1369 -2079 1371
rect -2069 1369 -2068 1376
rect -2325 1360 -2317 1368
rect -2079 1364 -2071 1369
rect -2325 1340 -2320 1360
rect -2317 1352 -2309 1360
rect -2074 1355 -2071 1364
rect -2069 1360 -2068 1364
rect -2109 1346 -2079 1349
rect -2325 1334 -2317 1340
rect -2119 1334 -2069 1336
rect -2056 1334 -2026 1337
rect -2000 1334 -1992 1380
rect -1846 1378 -1806 1380
rect -1854 1373 -1806 1377
rect -1854 1371 -1846 1373
rect -1846 1369 -1806 1371
rect -1806 1367 -1798 1369
rect -1846 1364 -1798 1367
rect -1846 1351 -1806 1362
rect -1671 1360 -1663 1368
rect -1663 1352 -1655 1360
rect -1854 1346 -1680 1350
rect -1926 1334 -1892 1337
rect -1671 1334 -1663 1340
rect -1642 1334 -1637 1380
rect -1619 1334 -1614 1380
rect -1565 1358 -1531 1359
rect -1530 1358 -1526 1380
rect -1506 1358 -1502 1380
rect -1482 1358 -1478 1380
rect -1458 1358 -1454 1380
rect -1434 1358 -1430 1380
rect -1410 1358 -1406 1380
rect -1386 1358 -1382 1380
rect -1362 1358 -1358 1380
rect -1338 1358 -1334 1380
rect -1314 1358 -1310 1380
rect -1290 1358 -1286 1380
rect -1266 1358 -1262 1380
rect -1242 1358 -1238 1380
rect -1218 1358 -1214 1380
rect -1194 1358 -1190 1380
rect -1170 1358 -1166 1380
rect -1146 1358 -1142 1380
rect -1122 1358 -1118 1380
rect -1098 1358 -1094 1380
rect -1074 1358 -1070 1380
rect -1050 1379 -1046 1380
rect -1565 1356 -1053 1358
rect -1555 1335 -1547 1349
rect -2393 1332 -1557 1334
rect -1530 1332 -1526 1356
rect -2371 1310 -2366 1332
rect -2348 1310 -2343 1332
rect -2325 1328 -2317 1332
rect -2325 1312 -2320 1328
rect -2317 1324 -2309 1328
rect -2309 1312 -2301 1324
rect -2109 1315 -2079 1322
rect -2000 1321 -1992 1332
rect -1671 1328 -1663 1332
rect -1846 1324 -1806 1326
rect -1663 1324 -1655 1328
rect -2009 1318 -1992 1321
rect -1854 1318 -1806 1322
rect -2071 1315 -1992 1318
rect -1983 1315 -1806 1318
rect -2009 1312 -1992 1315
rect -2325 1310 -2317 1312
rect -2033 1310 -1992 1312
rect -1846 1311 -1806 1313
rect -1655 1312 -1647 1324
rect -1864 1310 -1796 1311
rect -1671 1310 -1663 1312
rect -1642 1310 -1637 1332
rect -1619 1310 -1614 1332
rect -1571 1331 -1557 1332
rect -1554 1318 -1547 1332
rect -1530 1310 -1523 1331
rect -1506 1310 -1502 1356
rect -1482 1310 -1478 1356
rect -1458 1310 -1454 1356
rect -1434 1310 -1430 1356
rect -1410 1310 -1406 1356
rect -1386 1310 -1382 1356
rect -1362 1310 -1358 1356
rect -1338 1310 -1334 1356
rect -1314 1310 -1310 1356
rect -1290 1310 -1286 1356
rect -1266 1310 -1262 1356
rect -1242 1310 -1238 1356
rect -1218 1310 -1214 1356
rect -1194 1310 -1190 1356
rect -1170 1311 -1166 1356
rect -1181 1310 -1147 1311
rect -2393 1308 -1557 1310
rect -1547 1308 -1147 1310
rect -2371 1286 -2366 1308
rect -2348 1286 -2343 1308
rect -2325 1300 -2317 1308
rect -2079 1305 -2035 1308
rect -2013 1306 -1992 1308
rect -2000 1305 -1992 1306
rect -1904 1305 -1798 1308
rect -2101 1301 -2009 1305
rect -2023 1300 -2009 1301
rect -2000 1303 -1798 1305
rect -2000 1301 -1854 1303
rect -1846 1301 -1798 1303
rect -2325 1286 -2320 1300
rect -2317 1296 -2309 1300
rect -2309 1286 -2301 1296
rect -2109 1288 -2101 1295
rect -2023 1291 -2021 1300
rect -2000 1291 -1992 1301
rect -1671 1300 -1663 1308
rect -1846 1297 -1806 1299
rect -1663 1296 -1655 1300
rect -1854 1291 -1806 1295
rect -2071 1288 -1806 1291
rect -2074 1286 -2031 1288
rect -2000 1286 -1992 1288
rect -1655 1286 -1647 1296
rect -1642 1286 -1637 1308
rect -1619 1286 -1614 1308
rect -1571 1307 -1557 1308
rect -1554 1307 -1533 1308
rect -1554 1294 -1547 1307
rect -1530 1286 -1523 1308
rect -1506 1286 -1502 1308
rect -1482 1286 -1478 1308
rect -1458 1286 -1454 1308
rect -1434 1286 -1430 1308
rect -1410 1286 -1406 1308
rect -1386 1286 -1382 1308
rect -1362 1286 -1358 1308
rect -1338 1286 -1334 1308
rect -1314 1286 -1310 1308
rect -1290 1286 -1286 1308
rect -1266 1286 -1262 1308
rect -1242 1286 -1238 1308
rect -1218 1286 -1214 1308
rect -1194 1286 -1190 1308
rect -1181 1301 -1176 1308
rect -1170 1301 -1166 1308
rect -1171 1287 -1166 1301
rect -1170 1286 -1166 1287
rect -1146 1286 -1142 1356
rect -1122 1286 -1118 1356
rect -1098 1286 -1094 1356
rect -1074 1286 -1070 1356
rect -1067 1355 -1053 1356
rect -1050 1334 -1043 1379
rect -1026 1334 -1022 1380
rect -1002 1334 -998 1380
rect -978 1334 -974 1380
rect -954 1334 -950 1380
rect -930 1334 -926 1380
rect -906 1334 -902 1380
rect -882 1334 -878 1380
rect -858 1334 -854 1380
rect -834 1334 -830 1380
rect -810 1334 -806 1380
rect -786 1334 -782 1380
rect -762 1334 -758 1380
rect -738 1334 -734 1380
rect -714 1334 -710 1380
rect -690 1334 -686 1380
rect -666 1334 -662 1380
rect -642 1334 -638 1380
rect -618 1334 -614 1380
rect -594 1334 -590 1380
rect -570 1334 -566 1380
rect -546 1334 -542 1380
rect -522 1334 -518 1380
rect -498 1334 -494 1380
rect -474 1334 -470 1380
rect -450 1334 -446 1380
rect -426 1334 -422 1380
rect -402 1334 -398 1380
rect -378 1334 -374 1380
rect -354 1334 -350 1380
rect -330 1334 -326 1380
rect -306 1334 -302 1380
rect -282 1334 -278 1380
rect -258 1334 -254 1380
rect -210 1334 -206 1380
rect -186 1334 -182 1380
rect -162 1334 -158 1380
rect -138 1334 -134 1380
rect -114 1334 -110 1380
rect -90 1334 -86 1380
rect -66 1334 -62 1380
rect -42 1334 -38 1380
rect -18 1334 -14 1380
rect -5 1373 0 1380
rect 6 1373 10 1380
rect 5 1359 10 1373
rect 30 1334 34 1428
rect 54 1334 58 1428
rect 78 1334 82 1428
rect 102 1334 106 1428
rect 126 1335 130 1428
rect 115 1334 149 1335
rect -1067 1332 149 1334
rect -1067 1331 -1053 1332
rect -1050 1331 -1043 1332
rect -1050 1286 -1046 1331
rect -1026 1286 -1022 1332
rect -1002 1286 -998 1332
rect -978 1286 -974 1332
rect -954 1286 -950 1332
rect -930 1286 -926 1332
rect -906 1286 -902 1332
rect -882 1286 -878 1332
rect -858 1286 -854 1332
rect -834 1286 -830 1332
rect -810 1286 -806 1332
rect -786 1286 -782 1332
rect -762 1286 -758 1332
rect -738 1286 -734 1332
rect -714 1286 -710 1332
rect -690 1286 -686 1332
rect -666 1286 -662 1332
rect -642 1286 -638 1332
rect -618 1286 -614 1332
rect -594 1286 -590 1332
rect -570 1286 -566 1332
rect -546 1286 -542 1332
rect -522 1286 -518 1332
rect -498 1286 -494 1332
rect -474 1286 -470 1332
rect -450 1286 -446 1332
rect -426 1286 -422 1332
rect -402 1286 -398 1332
rect -378 1286 -374 1332
rect -354 1286 -350 1332
rect -330 1286 -326 1332
rect -306 1286 -302 1332
rect -282 1286 -278 1332
rect -258 1286 -254 1332
rect -210 1331 -206 1332
rect -245 1308 -213 1311
rect -245 1301 -240 1308
rect -227 1307 -213 1308
rect -210 1307 -203 1331
rect -235 1287 -230 1301
rect -234 1286 -230 1287
rect -186 1286 -182 1332
rect -162 1286 -158 1332
rect -138 1286 -134 1332
rect -114 1286 -110 1332
rect -90 1286 -86 1332
rect -66 1286 -62 1332
rect -42 1286 -38 1332
rect -18 1286 -14 1332
rect 30 1307 34 1332
rect -2393 1284 -1557 1286
rect -1547 1284 27 1286
rect -2371 1238 -2366 1284
rect -2348 1238 -2343 1284
rect -2325 1272 -2317 1284
rect -2074 1281 -2071 1284
rect -2101 1274 -2071 1281
rect -2325 1252 -2320 1272
rect -2317 1268 -2309 1272
rect -2064 1270 -2061 1278
rect -2325 1244 -2317 1252
rect -2101 1247 -2071 1250
rect -2325 1238 -2320 1244
rect -2317 1238 -2309 1244
rect -2000 1242 -1992 1284
rect -1846 1283 -1806 1284
rect -1846 1274 -1798 1281
rect -1671 1272 -1663 1284
rect -1846 1270 -1806 1272
rect -1663 1268 -1655 1272
rect -1854 1256 -1680 1260
rect -1846 1247 -1798 1250
rect -2079 1241 -2043 1242
rect -2007 1241 -1991 1242
rect -2079 1240 -2071 1241
rect -2079 1238 -2029 1240
rect -2011 1238 -1991 1241
rect -1846 1239 -1806 1245
rect -1671 1244 -1663 1252
rect -1864 1238 -1796 1239
rect -1663 1238 -1655 1244
rect -1642 1238 -1637 1284
rect -1619 1238 -1614 1284
rect -1571 1283 -1557 1284
rect -1554 1283 -1533 1284
rect -1530 1262 -1523 1284
rect -1506 1262 -1502 1284
rect -1482 1262 -1478 1284
rect -1458 1262 -1454 1284
rect -1434 1262 -1430 1284
rect -1410 1262 -1406 1284
rect -1386 1262 -1382 1284
rect -1362 1262 -1358 1284
rect -1338 1262 -1334 1284
rect -1314 1262 -1310 1284
rect -1290 1262 -1286 1284
rect -1266 1262 -1262 1284
rect -1242 1262 -1238 1284
rect -1218 1262 -1214 1284
rect -1194 1262 -1190 1284
rect -1170 1262 -1166 1284
rect -1146 1262 -1142 1284
rect -1122 1262 -1118 1284
rect -1098 1262 -1094 1284
rect -1074 1262 -1070 1284
rect -1050 1262 -1046 1284
rect -1026 1262 -1022 1284
rect -1002 1262 -998 1284
rect -978 1262 -974 1284
rect -954 1262 -950 1284
rect -930 1262 -926 1284
rect -906 1262 -902 1284
rect -882 1262 -878 1284
rect -858 1262 -854 1284
rect -834 1262 -830 1284
rect -810 1262 -806 1284
rect -786 1262 -782 1284
rect -762 1262 -758 1284
rect -738 1263 -734 1284
rect -749 1262 -715 1263
rect -1547 1260 -715 1262
rect -1547 1259 -1533 1260
rect -1530 1259 -1523 1260
rect -1530 1238 -1526 1259
rect -1506 1238 -1502 1260
rect -1482 1238 -1478 1260
rect -1458 1238 -1454 1260
rect -1434 1238 -1430 1260
rect -1410 1238 -1406 1260
rect -1386 1238 -1382 1260
rect -1362 1238 -1358 1260
rect -1338 1238 -1334 1260
rect -1314 1238 -1310 1260
rect -1290 1238 -1286 1260
rect -1266 1238 -1262 1260
rect -1242 1238 -1238 1260
rect -1218 1238 -1214 1260
rect -1194 1238 -1190 1260
rect -1170 1238 -1166 1260
rect -1146 1238 -1142 1260
rect -1122 1238 -1118 1260
rect -1098 1238 -1094 1260
rect -1074 1238 -1070 1260
rect -1050 1238 -1046 1260
rect -1026 1238 -1022 1260
rect -1002 1238 -998 1260
rect -978 1238 -974 1260
rect -954 1238 -950 1260
rect -930 1238 -926 1260
rect -906 1238 -902 1260
rect -882 1238 -878 1260
rect -858 1238 -854 1260
rect -834 1238 -830 1260
rect -810 1238 -806 1260
rect -786 1238 -782 1260
rect -762 1238 -758 1260
rect -749 1253 -744 1260
rect -738 1253 -734 1260
rect -739 1239 -734 1253
rect -714 1238 -710 1284
rect -690 1238 -686 1284
rect -666 1238 -662 1284
rect -642 1238 -638 1284
rect -618 1238 -614 1284
rect -594 1238 -590 1284
rect -570 1238 -566 1284
rect -546 1238 -542 1284
rect -522 1238 -518 1284
rect -498 1238 -494 1284
rect -474 1238 -470 1284
rect -450 1238 -446 1284
rect -426 1238 -422 1284
rect -402 1238 -398 1284
rect -378 1238 -374 1284
rect -354 1238 -350 1284
rect -330 1238 -326 1284
rect -306 1238 -302 1284
rect -282 1238 -278 1284
rect -258 1238 -254 1284
rect -234 1238 -230 1284
rect -186 1238 -182 1284
rect -162 1238 -158 1284
rect -138 1238 -134 1284
rect -114 1238 -110 1284
rect -90 1238 -86 1284
rect -66 1238 -62 1284
rect -42 1238 -38 1284
rect -18 1238 -14 1284
rect 13 1283 27 1284
rect 30 1283 37 1307
rect -5 1262 29 1263
rect 54 1262 58 1332
rect 78 1262 82 1332
rect 102 1262 106 1332
rect 115 1325 120 1332
rect 126 1325 130 1332
rect 125 1311 130 1325
rect 150 1262 154 1428
rect 174 1262 178 1428
rect 181 1427 195 1428
rect 198 1403 205 1451
rect 198 1262 202 1403
rect 222 1262 226 1476
rect 246 1262 250 1476
rect 270 1262 274 1476
rect 294 1262 298 1476
rect 318 1262 322 1476
rect 342 1475 346 1476
rect 342 1430 349 1475
rect 366 1430 370 1476
rect 390 1430 394 1476
rect 414 1430 418 1476
rect 438 1430 442 1476
rect 462 1430 466 1476
rect 486 1430 490 1476
rect 510 1430 514 1476
rect 534 1430 538 1476
rect 558 1430 562 1476
rect 582 1430 586 1476
rect 606 1430 610 1476
rect 630 1430 634 1476
rect 654 1430 658 1476
rect 678 1430 682 1476
rect 702 1430 706 1476
rect 726 1430 730 1476
rect 750 1430 754 1476
rect 774 1430 778 1476
rect 798 1430 802 1476
rect 822 1430 826 1476
rect 846 1430 850 1476
rect 870 1430 874 1476
rect 894 1430 898 1476
rect 918 1430 922 1476
rect 942 1430 946 1476
rect 966 1430 970 1476
rect 990 1430 994 1476
rect 1014 1430 1018 1476
rect 1038 1430 1042 1476
rect 1062 1430 1066 1476
rect 1086 1430 1090 1476
rect 1110 1430 1114 1476
rect 1134 1430 1138 1476
rect 1158 1430 1162 1476
rect 1182 1430 1186 1476
rect 1206 1430 1210 1476
rect 1230 1430 1234 1476
rect 1254 1430 1258 1476
rect 1278 1430 1282 1476
rect 1302 1430 1306 1476
rect 1326 1430 1330 1476
rect 1350 1430 1354 1476
rect 1374 1430 1378 1476
rect 1398 1430 1402 1476
rect 1422 1430 1426 1476
rect 1446 1430 1450 1476
rect 1470 1430 1474 1476
rect 1494 1430 1498 1476
rect 1518 1430 1522 1476
rect 1542 1430 1546 1476
rect 1566 1430 1570 1476
rect 1590 1430 1594 1476
rect 1614 1430 1618 1476
rect 1638 1430 1642 1476
rect 1662 1430 1666 1476
rect 1686 1430 1690 1476
rect 1710 1430 1714 1476
rect 1734 1430 1738 1476
rect 1758 1430 1762 1476
rect 1782 1430 1786 1476
rect 1795 1469 1800 1476
rect 1805 1455 1810 1469
rect 1806 1431 1810 1455
rect 1795 1430 1829 1431
rect 325 1428 1829 1430
rect 325 1427 339 1428
rect 342 1427 349 1428
rect 342 1262 346 1427
rect 366 1262 370 1428
rect 390 1262 394 1428
rect 414 1262 418 1428
rect 438 1262 442 1428
rect 462 1262 466 1428
rect 486 1262 490 1428
rect 510 1262 514 1428
rect 534 1262 538 1428
rect 558 1262 562 1428
rect 582 1262 586 1428
rect 606 1262 610 1428
rect 630 1262 634 1428
rect 654 1262 658 1428
rect 678 1262 682 1428
rect 702 1262 706 1428
rect 726 1262 730 1428
rect 750 1262 754 1428
rect 774 1262 778 1428
rect 798 1262 802 1428
rect 822 1262 826 1428
rect 846 1262 850 1428
rect 870 1262 874 1428
rect 894 1262 898 1428
rect 918 1262 922 1428
rect 931 1277 936 1287
rect 942 1277 946 1428
rect 941 1263 946 1277
rect 966 1262 970 1428
rect 990 1262 994 1428
rect 1014 1262 1018 1428
rect 1038 1262 1042 1428
rect 1062 1262 1066 1428
rect 1086 1262 1090 1428
rect 1110 1262 1114 1428
rect 1134 1262 1138 1428
rect 1158 1262 1162 1428
rect 1182 1262 1186 1428
rect 1206 1262 1210 1428
rect 1230 1262 1234 1428
rect 1254 1262 1258 1428
rect 1278 1262 1282 1428
rect 1302 1262 1306 1428
rect 1326 1262 1330 1428
rect 1350 1262 1354 1428
rect 1374 1262 1378 1428
rect 1398 1262 1402 1428
rect 1422 1262 1426 1428
rect 1446 1262 1450 1428
rect 1470 1262 1474 1428
rect 1494 1262 1498 1428
rect 1518 1262 1522 1428
rect 1542 1262 1546 1428
rect 1566 1262 1570 1428
rect 1590 1262 1594 1428
rect 1614 1262 1618 1428
rect 1638 1262 1642 1428
rect 1662 1262 1666 1428
rect 1686 1262 1690 1428
rect 1710 1262 1714 1428
rect 1734 1263 1738 1428
rect 1747 1301 1752 1311
rect 1758 1301 1762 1428
rect 1771 1349 1776 1359
rect 1782 1349 1786 1428
rect 1795 1421 1800 1428
rect 1806 1421 1810 1428
rect 1805 1407 1810 1421
rect 1819 1417 1827 1421
rect 1813 1407 1819 1417
rect 1781 1335 1786 1349
rect 1757 1287 1762 1301
rect 1723 1262 1757 1263
rect -5 1260 1757 1262
rect -5 1253 0 1260
rect 5 1239 10 1253
rect 6 1238 10 1239
rect 54 1238 58 1260
rect 78 1238 82 1260
rect 102 1238 106 1260
rect 150 1259 154 1260
rect -2393 1236 147 1238
rect -2371 1190 -2366 1236
rect -2348 1190 -2343 1236
rect -2325 1224 -2320 1236
rect -2079 1234 -2071 1236
rect -2072 1232 -2071 1234
rect -2109 1227 -2101 1232
rect -2101 1225 -2079 1227
rect -2069 1225 -2068 1232
rect -2325 1216 -2317 1224
rect -2079 1220 -2071 1225
rect -2325 1196 -2320 1216
rect -2317 1208 -2309 1216
rect -2074 1211 -2071 1220
rect -2069 1216 -2068 1220
rect -2109 1202 -2079 1205
rect -2325 1190 -2317 1196
rect -2119 1190 -2069 1192
rect -2056 1190 -2026 1193
rect -2000 1190 -1992 1236
rect -1846 1234 -1806 1236
rect -1854 1229 -1806 1233
rect -1854 1227 -1846 1229
rect -1846 1225 -1806 1227
rect -1806 1223 -1798 1225
rect -1846 1220 -1798 1223
rect -1846 1207 -1806 1218
rect -1671 1216 -1663 1224
rect -1663 1208 -1655 1216
rect -1854 1202 -1680 1206
rect -1926 1190 -1892 1193
rect -1671 1190 -1663 1196
rect -1642 1190 -1637 1236
rect -1619 1190 -1614 1236
rect -1530 1190 -1526 1236
rect -1506 1190 -1502 1236
rect -1482 1190 -1478 1236
rect -1458 1190 -1454 1236
rect -1434 1190 -1430 1236
rect -1410 1190 -1406 1236
rect -1386 1190 -1382 1236
rect -1362 1190 -1358 1236
rect -1338 1190 -1334 1236
rect -1314 1190 -1310 1236
rect -1290 1190 -1286 1236
rect -1266 1190 -1262 1236
rect -1242 1190 -1238 1236
rect -1218 1190 -1214 1236
rect -1194 1190 -1190 1236
rect -1170 1190 -1166 1236
rect -1146 1235 -1142 1236
rect -1146 1211 -1139 1235
rect -1146 1190 -1142 1211
rect -1122 1190 -1118 1236
rect -1098 1190 -1094 1236
rect -1074 1190 -1070 1236
rect -1050 1190 -1046 1236
rect -1026 1190 -1022 1236
rect -1002 1190 -998 1236
rect -978 1190 -974 1236
rect -954 1190 -950 1236
rect -930 1190 -926 1236
rect -906 1190 -902 1236
rect -882 1190 -878 1236
rect -858 1190 -854 1236
rect -834 1190 -830 1236
rect -810 1190 -806 1236
rect -786 1190 -782 1236
rect -762 1190 -758 1236
rect -749 1205 -744 1215
rect -739 1191 -734 1205
rect -738 1190 -734 1191
rect -714 1190 -710 1236
rect -690 1190 -686 1236
rect -666 1190 -662 1236
rect -642 1190 -638 1236
rect -618 1190 -614 1236
rect -594 1190 -590 1236
rect -570 1191 -566 1236
rect -581 1190 -547 1191
rect -2393 1188 -547 1190
rect -2371 1166 -2366 1188
rect -2348 1166 -2343 1188
rect -2325 1184 -2317 1188
rect -2325 1168 -2320 1184
rect -2317 1180 -2309 1184
rect -2309 1168 -2301 1180
rect -2109 1171 -2079 1178
rect -2000 1177 -1992 1188
rect -1671 1184 -1663 1188
rect -1846 1180 -1806 1182
rect -1663 1180 -1655 1184
rect -2009 1174 -1992 1177
rect -1854 1174 -1806 1178
rect -2071 1171 -1992 1174
rect -1983 1171 -1806 1174
rect -2009 1168 -1992 1171
rect -2325 1166 -2317 1168
rect -2033 1166 -1992 1168
rect -1846 1167 -1806 1169
rect -1655 1168 -1647 1180
rect -1864 1166 -1796 1167
rect -1671 1166 -1663 1168
rect -1642 1166 -1637 1188
rect -1619 1166 -1614 1188
rect -1530 1166 -1526 1188
rect -1506 1166 -1502 1188
rect -1482 1166 -1478 1188
rect -1458 1166 -1454 1188
rect -1434 1166 -1430 1188
rect -1410 1166 -1406 1188
rect -1386 1166 -1382 1188
rect -1362 1166 -1358 1188
rect -1338 1166 -1334 1188
rect -1314 1166 -1310 1188
rect -1290 1166 -1286 1188
rect -1266 1166 -1262 1188
rect -1242 1166 -1238 1188
rect -1218 1166 -1214 1188
rect -1194 1166 -1190 1188
rect -1170 1166 -1166 1188
rect -1146 1166 -1142 1188
rect -1122 1166 -1118 1188
rect -1098 1166 -1094 1188
rect -1074 1166 -1070 1188
rect -1050 1166 -1046 1188
rect -1026 1166 -1022 1188
rect -1002 1166 -998 1188
rect -978 1166 -974 1188
rect -954 1166 -950 1188
rect -930 1166 -926 1188
rect -906 1166 -902 1188
rect -882 1166 -878 1188
rect -858 1166 -854 1188
rect -834 1166 -830 1188
rect -810 1166 -806 1188
rect -786 1166 -782 1188
rect -762 1166 -758 1188
rect -738 1166 -734 1188
rect -714 1187 -710 1188
rect -2393 1164 -717 1166
rect -2371 1142 -2366 1164
rect -2348 1142 -2343 1164
rect -2325 1156 -2317 1164
rect -2079 1161 -2035 1164
rect -2013 1162 -1992 1164
rect -2000 1161 -1992 1162
rect -1904 1161 -1798 1164
rect -2101 1157 -2009 1161
rect -2023 1156 -2009 1157
rect -2000 1159 -1798 1161
rect -2000 1157 -1854 1159
rect -1846 1157 -1798 1159
rect -2325 1142 -2320 1156
rect -2317 1152 -2309 1156
rect -2309 1142 -2301 1152
rect -2109 1144 -2101 1151
rect -2023 1147 -2021 1156
rect -2000 1147 -1992 1157
rect -1671 1156 -1663 1164
rect -1846 1153 -1806 1155
rect -1663 1152 -1655 1156
rect -1854 1147 -1806 1151
rect -2071 1144 -1806 1147
rect -2074 1142 -2031 1144
rect -2000 1142 -1992 1144
rect -1655 1142 -1647 1152
rect -1642 1142 -1637 1164
rect -1619 1142 -1614 1164
rect -1530 1142 -1526 1164
rect -1506 1142 -1502 1164
rect -1482 1142 -1478 1164
rect -1458 1142 -1454 1164
rect -1434 1142 -1430 1164
rect -1410 1142 -1406 1164
rect -1386 1142 -1382 1164
rect -1362 1142 -1358 1164
rect -1338 1142 -1334 1164
rect -1314 1142 -1310 1164
rect -1290 1142 -1286 1164
rect -1266 1142 -1262 1164
rect -1242 1142 -1238 1164
rect -1218 1142 -1214 1164
rect -1194 1142 -1190 1164
rect -1170 1142 -1166 1164
rect -1146 1142 -1142 1164
rect -1122 1142 -1118 1164
rect -1098 1142 -1094 1164
rect -1074 1142 -1070 1164
rect -1050 1142 -1046 1164
rect -1026 1142 -1022 1164
rect -1002 1142 -998 1164
rect -978 1142 -974 1164
rect -954 1142 -950 1164
rect -930 1142 -926 1164
rect -906 1142 -902 1164
rect -882 1142 -878 1164
rect -858 1142 -854 1164
rect -834 1142 -830 1164
rect -810 1142 -806 1164
rect -786 1142 -782 1164
rect -762 1142 -758 1164
rect -738 1142 -734 1164
rect -731 1163 -717 1164
rect -714 1163 -707 1187
rect -690 1142 -686 1188
rect -666 1142 -662 1188
rect -642 1142 -638 1188
rect -618 1142 -614 1188
rect -594 1142 -590 1188
rect -581 1181 -576 1188
rect -570 1181 -566 1188
rect -571 1167 -566 1181
rect -581 1157 -576 1167
rect -571 1143 -566 1157
rect -570 1142 -566 1143
rect -546 1142 -542 1236
rect -522 1142 -518 1236
rect -498 1142 -494 1236
rect -474 1142 -470 1236
rect -450 1142 -446 1236
rect -426 1142 -422 1236
rect -402 1142 -398 1236
rect -378 1142 -374 1236
rect -354 1142 -350 1236
rect -330 1142 -326 1236
rect -306 1142 -302 1236
rect -282 1142 -278 1236
rect -258 1142 -254 1236
rect -234 1142 -230 1236
rect -210 1214 -203 1235
rect -186 1214 -182 1236
rect -162 1214 -158 1236
rect -138 1214 -134 1236
rect -114 1214 -110 1236
rect -90 1214 -86 1236
rect -66 1214 -62 1236
rect -42 1214 -38 1236
rect -18 1214 -14 1236
rect 6 1214 10 1236
rect 54 1214 58 1236
rect 78 1214 82 1236
rect 102 1214 106 1236
rect 133 1235 147 1236
rect 150 1235 157 1259
rect 174 1214 178 1260
rect 198 1214 202 1260
rect 222 1214 226 1260
rect 246 1214 250 1260
rect 270 1214 274 1260
rect 294 1214 298 1260
rect 318 1214 322 1260
rect 342 1214 346 1260
rect 366 1214 370 1260
rect 390 1214 394 1260
rect 414 1214 418 1260
rect 438 1214 442 1260
rect 462 1214 466 1260
rect 486 1214 490 1260
rect 510 1214 514 1260
rect 534 1214 538 1260
rect 558 1214 562 1260
rect 582 1214 586 1260
rect 606 1214 610 1260
rect 630 1214 634 1260
rect 654 1214 658 1260
rect 678 1214 682 1260
rect 702 1214 706 1260
rect 726 1214 730 1260
rect 750 1214 754 1260
rect 774 1214 778 1260
rect 798 1214 802 1260
rect 822 1214 826 1260
rect 846 1214 850 1260
rect 870 1214 874 1260
rect 894 1214 898 1260
rect 918 1214 922 1260
rect 966 1214 970 1260
rect 990 1214 994 1260
rect 1014 1214 1018 1260
rect 1038 1214 1042 1260
rect 1062 1214 1066 1260
rect 1086 1214 1090 1260
rect 1110 1214 1114 1260
rect 1123 1229 1128 1239
rect 1134 1229 1138 1260
rect 1133 1215 1138 1229
rect 1158 1214 1162 1260
rect 1182 1214 1186 1260
rect 1206 1214 1210 1260
rect 1230 1214 1234 1260
rect 1254 1214 1258 1260
rect 1278 1214 1282 1260
rect 1302 1214 1306 1260
rect 1326 1214 1330 1260
rect 1350 1214 1354 1260
rect 1374 1214 1378 1260
rect 1398 1214 1402 1260
rect 1422 1214 1426 1260
rect 1446 1214 1450 1260
rect 1470 1214 1474 1260
rect 1494 1214 1498 1260
rect 1518 1214 1522 1260
rect 1542 1214 1546 1260
rect 1566 1214 1570 1260
rect 1590 1214 1594 1260
rect 1614 1214 1618 1260
rect 1638 1214 1642 1260
rect 1662 1214 1666 1260
rect 1686 1214 1690 1260
rect 1710 1215 1714 1260
rect 1723 1253 1728 1260
rect 1734 1253 1738 1260
rect 1733 1239 1738 1253
rect 1699 1214 1733 1215
rect -227 1212 1733 1214
rect -227 1211 -213 1212
rect -210 1211 -203 1212
rect -210 1142 -206 1211
rect -186 1142 -182 1212
rect -162 1142 -158 1212
rect -138 1142 -134 1212
rect -114 1142 -110 1212
rect -90 1142 -86 1212
rect -66 1142 -62 1212
rect -42 1142 -38 1212
rect -18 1142 -14 1212
rect 6 1142 10 1212
rect 30 1166 37 1187
rect 54 1167 58 1212
rect 43 1166 77 1167
rect 13 1164 77 1166
rect 13 1163 27 1164
rect 30 1163 37 1164
rect 30 1142 34 1163
rect 43 1157 48 1164
rect 54 1157 58 1164
rect 53 1143 58 1157
rect 78 1142 82 1212
rect 102 1142 106 1212
rect 115 1190 149 1191
rect 174 1190 178 1212
rect 198 1190 202 1212
rect 222 1190 226 1212
rect 246 1190 250 1212
rect 270 1190 274 1212
rect 294 1190 298 1212
rect 318 1190 322 1212
rect 342 1190 346 1212
rect 366 1190 370 1212
rect 390 1190 394 1212
rect 414 1190 418 1212
rect 438 1190 442 1212
rect 462 1190 466 1212
rect 486 1190 490 1212
rect 510 1190 514 1212
rect 534 1190 538 1212
rect 558 1190 562 1212
rect 582 1190 586 1212
rect 606 1190 610 1212
rect 630 1190 634 1212
rect 654 1190 658 1212
rect 678 1190 682 1212
rect 702 1190 706 1212
rect 726 1190 730 1212
rect 750 1190 754 1212
rect 774 1190 778 1212
rect 798 1190 802 1212
rect 822 1190 826 1212
rect 846 1190 850 1212
rect 870 1190 874 1212
rect 894 1190 898 1212
rect 918 1190 922 1212
rect 966 1211 970 1212
rect 115 1188 963 1190
rect 115 1181 120 1188
rect 125 1167 130 1181
rect 126 1142 130 1167
rect 174 1142 178 1188
rect 198 1142 202 1188
rect 222 1142 226 1188
rect 246 1142 250 1188
rect 270 1142 274 1188
rect 294 1142 298 1188
rect 318 1142 322 1188
rect 342 1142 346 1188
rect 366 1142 370 1188
rect 390 1142 394 1188
rect 414 1142 418 1188
rect 438 1142 442 1188
rect 462 1142 466 1188
rect 486 1142 490 1188
rect 510 1142 514 1188
rect 534 1142 538 1188
rect 558 1142 562 1188
rect 582 1142 586 1188
rect 606 1142 610 1188
rect 630 1142 634 1188
rect 654 1142 658 1188
rect 678 1142 682 1188
rect 702 1142 706 1188
rect 726 1142 730 1188
rect 750 1142 754 1188
rect 774 1142 778 1188
rect 798 1142 802 1188
rect 822 1142 826 1188
rect 846 1143 850 1188
rect 835 1142 869 1143
rect -2393 1140 869 1142
rect -2371 1094 -2366 1140
rect -2348 1094 -2343 1140
rect -2325 1128 -2317 1140
rect -2074 1137 -2071 1140
rect -2101 1130 -2071 1137
rect -2325 1108 -2320 1128
rect -2317 1124 -2309 1128
rect -2064 1126 -2061 1134
rect -2325 1100 -2317 1108
rect -2101 1103 -2071 1106
rect -2325 1094 -2320 1100
rect -2317 1094 -2309 1100
rect -2000 1098 -1992 1140
rect -1846 1139 -1806 1140
rect -1846 1130 -1798 1137
rect -1671 1128 -1663 1140
rect -1846 1126 -1806 1128
rect -1663 1124 -1655 1128
rect -1854 1112 -1680 1116
rect -1846 1103 -1798 1106
rect -2079 1097 -2043 1098
rect -2007 1097 -1991 1098
rect -2079 1096 -2071 1097
rect -2079 1094 -2029 1096
rect -2011 1094 -1991 1097
rect -1846 1095 -1806 1101
rect -1671 1100 -1663 1108
rect -1864 1094 -1796 1095
rect -1663 1094 -1655 1100
rect -1642 1094 -1637 1140
rect -1619 1094 -1614 1140
rect -1530 1094 -1526 1140
rect -1506 1094 -1502 1140
rect -1482 1094 -1478 1140
rect -1458 1094 -1454 1140
rect -1434 1094 -1430 1140
rect -1410 1094 -1406 1140
rect -1386 1094 -1382 1140
rect -1362 1094 -1358 1140
rect -1338 1094 -1334 1140
rect -1314 1094 -1310 1140
rect -1290 1094 -1286 1140
rect -1266 1094 -1262 1140
rect -1242 1094 -1238 1140
rect -1218 1094 -1214 1140
rect -1194 1094 -1190 1140
rect -1170 1094 -1166 1140
rect -1146 1094 -1142 1140
rect -1122 1094 -1118 1140
rect -1098 1094 -1094 1140
rect -1074 1094 -1070 1140
rect -1050 1094 -1046 1140
rect -1026 1094 -1022 1140
rect -1002 1094 -998 1140
rect -978 1094 -974 1140
rect -954 1094 -950 1140
rect -930 1094 -926 1140
rect -906 1094 -902 1140
rect -882 1094 -878 1140
rect -858 1094 -854 1140
rect -834 1094 -830 1140
rect -810 1094 -806 1140
rect -786 1094 -782 1140
rect -762 1094 -758 1140
rect -738 1094 -734 1140
rect -714 1118 -707 1139
rect -690 1118 -686 1140
rect -666 1118 -662 1140
rect -642 1118 -638 1140
rect -618 1118 -614 1140
rect -594 1118 -590 1140
rect -570 1118 -566 1140
rect -546 1118 -542 1140
rect -522 1118 -518 1140
rect -498 1118 -494 1140
rect -474 1118 -470 1140
rect -450 1118 -446 1140
rect -426 1118 -422 1140
rect -402 1118 -398 1140
rect -378 1118 -374 1140
rect -354 1118 -350 1140
rect -330 1118 -326 1140
rect -306 1118 -302 1140
rect -282 1118 -278 1140
rect -258 1118 -254 1140
rect -234 1118 -230 1140
rect -210 1118 -206 1140
rect -186 1118 -182 1140
rect -162 1118 -158 1140
rect -138 1118 -134 1140
rect -114 1118 -110 1140
rect -90 1118 -86 1140
rect -66 1118 -62 1140
rect -42 1118 -38 1140
rect -18 1118 -14 1140
rect 6 1118 10 1140
rect 30 1118 34 1140
rect 43 1118 77 1119
rect 78 1118 82 1140
rect 102 1118 106 1140
rect 126 1119 130 1140
rect 115 1118 149 1119
rect -731 1116 149 1118
rect -731 1115 -717 1116
rect -714 1115 -707 1116
rect -714 1094 -710 1115
rect -690 1094 -686 1116
rect -666 1094 -662 1116
rect -642 1094 -638 1116
rect -618 1094 -614 1116
rect -594 1094 -590 1116
rect -570 1094 -566 1116
rect -546 1115 -542 1116
rect -2393 1092 -549 1094
rect -2371 1046 -2366 1092
rect -2348 1046 -2343 1092
rect -2325 1080 -2320 1092
rect -2079 1090 -2071 1092
rect -2072 1088 -2071 1090
rect -2109 1083 -2101 1088
rect -2101 1081 -2079 1083
rect -2069 1081 -2068 1088
rect -2325 1072 -2317 1080
rect -2079 1076 -2071 1081
rect -2325 1052 -2320 1072
rect -2317 1064 -2309 1072
rect -2074 1067 -2071 1076
rect -2069 1072 -2068 1076
rect -2109 1058 -2079 1061
rect -2325 1046 -2317 1052
rect -2119 1046 -2069 1048
rect -2056 1046 -2026 1049
rect -2000 1046 -1992 1092
rect -1846 1090 -1806 1092
rect -1854 1085 -1806 1089
rect -1854 1083 -1846 1085
rect -1846 1081 -1806 1083
rect -1806 1079 -1798 1081
rect -1846 1076 -1798 1079
rect -1846 1063 -1806 1074
rect -1671 1072 -1663 1080
rect -1663 1064 -1655 1072
rect -1854 1058 -1680 1062
rect -1926 1046 -1892 1049
rect -1671 1046 -1663 1052
rect -1642 1046 -1637 1092
rect -1619 1046 -1614 1092
rect -1530 1046 -1526 1092
rect -1506 1046 -1502 1092
rect -1482 1046 -1478 1092
rect -1458 1046 -1454 1092
rect -1434 1046 -1430 1092
rect -1410 1046 -1406 1092
rect -1386 1046 -1382 1092
rect -1362 1046 -1358 1092
rect -1338 1046 -1334 1092
rect -1314 1046 -1310 1092
rect -1290 1046 -1286 1092
rect -1266 1046 -1262 1092
rect -1242 1046 -1238 1092
rect -1218 1046 -1214 1092
rect -1194 1046 -1190 1092
rect -1170 1046 -1166 1092
rect -1146 1046 -1142 1092
rect -1122 1046 -1118 1092
rect -1098 1046 -1094 1092
rect -1074 1046 -1070 1092
rect -1050 1046 -1046 1092
rect -1026 1046 -1022 1092
rect -1002 1046 -998 1092
rect -978 1046 -974 1092
rect -954 1046 -950 1092
rect -930 1046 -926 1092
rect -906 1046 -902 1092
rect -882 1046 -878 1092
rect -858 1046 -854 1092
rect -834 1046 -830 1092
rect -810 1046 -806 1092
rect -786 1047 -782 1092
rect -797 1046 -763 1047
rect -2393 1044 -763 1046
rect -2371 1022 -2366 1044
rect -2348 1022 -2343 1044
rect -2325 1040 -2317 1044
rect -2325 1024 -2320 1040
rect -2317 1036 -2309 1040
rect -2309 1024 -2301 1036
rect -2109 1027 -2079 1034
rect -2000 1033 -1992 1044
rect -1671 1040 -1663 1044
rect -1846 1036 -1806 1038
rect -1663 1036 -1655 1040
rect -2009 1030 -1992 1033
rect -1854 1030 -1806 1034
rect -2071 1027 -1992 1030
rect -1983 1027 -1806 1030
rect -2009 1024 -1992 1027
rect -2325 1022 -2317 1024
rect -2033 1022 -1992 1024
rect -1846 1023 -1806 1025
rect -1655 1024 -1647 1036
rect -1864 1022 -1796 1023
rect -1671 1022 -1663 1024
rect -1642 1022 -1637 1044
rect -1619 1022 -1614 1044
rect -1530 1022 -1526 1044
rect -1506 1022 -1502 1044
rect -1482 1022 -1478 1044
rect -1458 1022 -1454 1044
rect -1434 1022 -1430 1044
rect -1410 1022 -1406 1044
rect -1386 1022 -1382 1044
rect -1362 1022 -1358 1044
rect -1338 1022 -1334 1044
rect -1314 1022 -1310 1044
rect -1290 1022 -1286 1044
rect -1266 1022 -1262 1044
rect -1242 1022 -1238 1044
rect -1218 1022 -1214 1044
rect -1194 1022 -1190 1044
rect -1170 1022 -1166 1044
rect -1146 1022 -1142 1044
rect -1122 1022 -1118 1044
rect -1098 1022 -1094 1044
rect -1074 1022 -1070 1044
rect -1050 1022 -1046 1044
rect -1026 1022 -1022 1044
rect -1002 1022 -998 1044
rect -978 1022 -974 1044
rect -954 1022 -950 1044
rect -930 1022 -926 1044
rect -906 1022 -902 1044
rect -882 1022 -878 1044
rect -858 1022 -854 1044
rect -834 1022 -830 1044
rect -810 1022 -806 1044
rect -797 1037 -792 1044
rect -786 1037 -782 1044
rect -787 1023 -782 1037
rect -797 1022 -763 1023
rect -762 1022 -758 1092
rect -738 1022 -734 1092
rect -714 1022 -710 1092
rect -690 1022 -686 1092
rect -666 1022 -662 1092
rect -642 1022 -638 1092
rect -618 1022 -614 1092
rect -594 1022 -590 1092
rect -570 1022 -566 1092
rect -563 1091 -549 1092
rect -546 1067 -539 1115
rect -546 1022 -542 1067
rect -522 1022 -518 1116
rect -498 1023 -494 1116
rect -509 1022 -475 1023
rect -2393 1020 -475 1022
rect -2371 998 -2366 1020
rect -2348 998 -2343 1020
rect -2325 1012 -2317 1020
rect -2079 1017 -2035 1020
rect -2013 1018 -1992 1020
rect -2000 1017 -1992 1018
rect -1904 1017 -1798 1020
rect -2101 1013 -2009 1017
rect -2023 1012 -2009 1013
rect -2000 1015 -1798 1017
rect -2000 1013 -1854 1015
rect -1846 1013 -1798 1015
rect -2325 998 -2320 1012
rect -2317 1008 -2309 1012
rect -2309 998 -2301 1008
rect -2109 1000 -2101 1007
rect -2023 1003 -2021 1012
rect -2000 1003 -1992 1013
rect -1671 1012 -1663 1020
rect -1846 1009 -1806 1011
rect -1663 1008 -1655 1012
rect -1854 1003 -1806 1007
rect -2071 1000 -1806 1003
rect -2074 998 -2031 1000
rect -2000 998 -1992 1000
rect -1655 998 -1647 1008
rect -1642 998 -1637 1020
rect -1619 998 -1614 1020
rect -1530 998 -1526 1020
rect -1506 998 -1502 1020
rect -1482 998 -1478 1020
rect -1458 998 -1454 1020
rect -1434 998 -1430 1020
rect -1410 998 -1406 1020
rect -1386 998 -1382 1020
rect -1362 998 -1358 1020
rect -1338 998 -1334 1020
rect -1314 998 -1310 1020
rect -1290 998 -1286 1020
rect -1266 998 -1262 1020
rect -1242 998 -1238 1020
rect -1218 998 -1214 1020
rect -1194 998 -1190 1020
rect -1170 998 -1166 1020
rect -1146 998 -1142 1020
rect -1122 998 -1118 1020
rect -1098 998 -1094 1020
rect -1074 998 -1070 1020
rect -1050 998 -1046 1020
rect -1026 998 -1022 1020
rect -1002 998 -998 1020
rect -978 998 -974 1020
rect -954 998 -950 1020
rect -930 998 -926 1020
rect -906 998 -902 1020
rect -882 998 -878 1020
rect -858 998 -854 1020
rect -834 998 -830 1020
rect -810 998 -806 1020
rect -797 1013 -792 1020
rect -787 999 -782 1013
rect -786 998 -782 999
rect -762 998 -758 1020
rect -738 998 -734 1020
rect -714 998 -710 1020
rect -690 998 -686 1020
rect -666 998 -662 1020
rect -642 998 -638 1020
rect -618 998 -614 1020
rect -594 998 -590 1020
rect -570 998 -566 1020
rect -546 998 -542 1020
rect -522 998 -518 1020
rect -509 1013 -504 1020
rect -498 1013 -494 1020
rect -499 999 -494 1013
rect -509 998 -475 999
rect -474 998 -470 1116
rect -450 998 -446 1116
rect -426 998 -422 1116
rect -402 998 -398 1116
rect -378 998 -374 1116
rect -354 998 -350 1116
rect -330 998 -326 1116
rect -306 998 -302 1116
rect -282 998 -278 1116
rect -258 998 -254 1116
rect -234 998 -230 1116
rect -210 998 -206 1116
rect -186 998 -182 1116
rect -162 998 -158 1116
rect -138 998 -134 1116
rect -114 998 -110 1116
rect -90 998 -86 1116
rect -66 998 -62 1116
rect -42 998 -38 1116
rect -18 998 -14 1116
rect 6 998 10 1116
rect 30 998 34 1116
rect 43 1109 48 1116
rect 53 1095 58 1109
rect 54 998 58 1095
rect 78 1091 82 1116
rect 78 1067 85 1091
rect 78 1019 85 1043
rect 78 998 82 1019
rect 102 998 106 1116
rect 115 1109 120 1116
rect 126 1109 130 1116
rect 125 1095 130 1109
rect 139 1105 147 1109
rect 133 1095 139 1105
rect 150 1094 157 1115
rect 174 1094 178 1140
rect 198 1094 202 1140
rect 222 1094 226 1140
rect 246 1094 250 1140
rect 270 1094 274 1140
rect 294 1094 298 1140
rect 318 1094 322 1140
rect 342 1094 346 1140
rect 366 1094 370 1140
rect 390 1094 394 1140
rect 414 1094 418 1140
rect 438 1094 442 1140
rect 462 1094 466 1140
rect 486 1094 490 1140
rect 510 1094 514 1140
rect 534 1094 538 1140
rect 558 1094 562 1140
rect 582 1094 586 1140
rect 606 1094 610 1140
rect 630 1094 634 1140
rect 654 1094 658 1140
rect 678 1094 682 1140
rect 702 1094 706 1140
rect 726 1094 730 1140
rect 750 1094 754 1140
rect 774 1094 778 1140
rect 798 1094 802 1140
rect 822 1094 826 1140
rect 835 1133 840 1140
rect 846 1133 850 1140
rect 845 1119 850 1133
rect 835 1118 869 1119
rect 870 1118 874 1188
rect 894 1118 898 1188
rect 918 1118 922 1188
rect 949 1187 963 1188
rect 966 1187 973 1211
rect 931 1166 965 1167
rect 990 1166 994 1212
rect 1014 1166 1018 1212
rect 1038 1166 1042 1212
rect 1062 1166 1066 1212
rect 1086 1166 1090 1212
rect 1110 1166 1114 1212
rect 1158 1166 1162 1212
rect 1182 1166 1186 1212
rect 1206 1166 1210 1212
rect 1230 1166 1234 1212
rect 1254 1166 1258 1212
rect 1278 1166 1282 1212
rect 1302 1166 1306 1212
rect 1326 1166 1330 1212
rect 1350 1166 1354 1212
rect 1374 1166 1378 1212
rect 1398 1166 1402 1212
rect 1422 1166 1426 1212
rect 1446 1166 1450 1212
rect 1470 1166 1474 1212
rect 1494 1166 1498 1212
rect 1518 1166 1522 1212
rect 1542 1166 1546 1212
rect 1566 1166 1570 1212
rect 1590 1166 1594 1212
rect 1614 1166 1618 1212
rect 1638 1166 1642 1212
rect 1662 1167 1666 1212
rect 1675 1181 1680 1191
rect 1686 1181 1690 1212
rect 1699 1205 1704 1212
rect 1710 1205 1714 1212
rect 1709 1191 1714 1205
rect 1685 1167 1690 1181
rect 1651 1166 1685 1167
rect 931 1164 1685 1166
rect 931 1157 936 1164
rect 941 1143 946 1157
rect 942 1118 946 1143
rect 990 1118 994 1164
rect 1014 1118 1018 1164
rect 1038 1118 1042 1164
rect 1062 1118 1066 1164
rect 1086 1118 1090 1164
rect 1110 1118 1114 1164
rect 1158 1163 1162 1164
rect 1123 1140 1155 1143
rect 1123 1133 1128 1140
rect 1141 1139 1155 1140
rect 1158 1139 1165 1163
rect 1133 1119 1138 1133
rect 1134 1118 1138 1119
rect 1182 1118 1186 1164
rect 1206 1118 1210 1164
rect 1230 1118 1234 1164
rect 1254 1118 1258 1164
rect 1278 1118 1282 1164
rect 1302 1118 1306 1164
rect 1326 1118 1330 1164
rect 1350 1118 1354 1164
rect 1374 1118 1378 1164
rect 1398 1118 1402 1164
rect 1422 1118 1426 1164
rect 1446 1118 1450 1164
rect 1470 1118 1474 1164
rect 1494 1118 1498 1164
rect 1518 1118 1522 1164
rect 1542 1118 1546 1164
rect 1566 1118 1570 1164
rect 1590 1118 1594 1164
rect 1614 1119 1618 1164
rect 1627 1133 1632 1143
rect 1638 1133 1642 1164
rect 1651 1157 1656 1164
rect 1662 1157 1666 1164
rect 1661 1143 1666 1157
rect 1637 1119 1642 1133
rect 1603 1118 1637 1119
rect 835 1116 1637 1118
rect 835 1109 840 1116
rect 845 1095 850 1109
rect 846 1094 850 1095
rect 870 1094 874 1116
rect 894 1095 898 1116
rect 883 1094 917 1095
rect 133 1092 917 1094
rect 133 1091 147 1092
rect 150 1091 157 1092
rect 115 1061 120 1071
rect 125 1047 130 1061
rect 126 998 130 1047
rect 150 1043 154 1091
rect 150 1019 157 1043
rect 174 998 178 1092
rect 198 998 202 1092
rect 222 998 226 1092
rect 246 998 250 1092
rect 270 998 274 1092
rect 294 998 298 1092
rect 318 998 322 1092
rect 342 998 346 1092
rect 366 998 370 1092
rect 390 998 394 1092
rect 414 998 418 1092
rect 438 998 442 1092
rect 462 998 466 1092
rect 486 998 490 1092
rect 510 998 514 1092
rect 534 998 538 1092
rect 558 998 562 1092
rect 582 998 586 1092
rect 606 998 610 1092
rect 630 998 634 1092
rect 654 998 658 1092
rect 678 998 682 1092
rect 702 998 706 1092
rect 726 998 730 1092
rect 750 998 754 1092
rect 774 998 778 1092
rect 798 998 802 1092
rect 822 998 826 1092
rect 846 998 850 1092
rect 870 1067 874 1092
rect 883 1085 888 1092
rect 894 1085 898 1092
rect 893 1071 898 1085
rect 870 1019 877 1067
rect 883 1037 888 1047
rect 893 1023 898 1037
rect 870 998 874 1019
rect 894 998 898 1023
rect 918 1019 922 1116
rect -2393 996 915 998
rect -2371 950 -2366 996
rect -2348 950 -2343 996
rect -2325 984 -2317 996
rect -2074 993 -2071 996
rect -2101 986 -2071 993
rect -2325 964 -2320 984
rect -2317 980 -2309 984
rect -2064 982 -2061 990
rect -2325 956 -2317 964
rect -2101 959 -2071 962
rect -2325 950 -2320 956
rect -2317 950 -2309 956
rect -2000 954 -1992 996
rect -1846 995 -1806 996
rect -1846 986 -1798 993
rect -1671 984 -1663 996
rect -1846 982 -1806 984
rect -1663 980 -1655 984
rect -1854 968 -1680 972
rect -1846 959 -1798 962
rect -2079 953 -2043 954
rect -2007 953 -1991 954
rect -2079 952 -2071 953
rect -2079 950 -2029 952
rect -2011 950 -1991 953
rect -1846 951 -1806 957
rect -1671 956 -1663 964
rect -1864 950 -1796 951
rect -1663 950 -1655 956
rect -1642 950 -1637 996
rect -1619 950 -1614 996
rect -1530 950 -1526 996
rect -1506 950 -1502 996
rect -1482 950 -1478 996
rect -1458 950 -1454 996
rect -1434 950 -1430 996
rect -1410 950 -1406 996
rect -1386 950 -1382 996
rect -1362 950 -1358 996
rect -1338 950 -1334 996
rect -1314 950 -1310 996
rect -1290 950 -1286 996
rect -1266 950 -1262 996
rect -1242 950 -1238 996
rect -1218 950 -1214 996
rect -1194 950 -1190 996
rect -1170 950 -1166 996
rect -1146 950 -1142 996
rect -1122 950 -1118 996
rect -1098 950 -1094 996
rect -1074 950 -1070 996
rect -1050 950 -1046 996
rect -1026 950 -1022 996
rect -1002 950 -998 996
rect -978 950 -974 996
rect -954 950 -950 996
rect -930 950 -926 996
rect -906 950 -902 996
rect -882 950 -878 996
rect -858 950 -854 996
rect -834 950 -830 996
rect -810 950 -806 996
rect -786 950 -782 996
rect -762 971 -758 996
rect -2393 948 -765 950
rect -2371 902 -2366 948
rect -2348 902 -2343 948
rect -2325 936 -2320 948
rect -2079 946 -2071 948
rect -2072 944 -2071 946
rect -2109 939 -2101 944
rect -2101 937 -2079 939
rect -2069 937 -2068 944
rect -2325 928 -2317 936
rect -2079 932 -2071 937
rect -2325 908 -2320 928
rect -2317 920 -2309 928
rect -2074 923 -2071 932
rect -2069 928 -2068 932
rect -2109 914 -2079 917
rect -2325 902 -2317 908
rect -2119 902 -2069 904
rect -2056 902 -2026 905
rect -2000 902 -1992 948
rect -1846 946 -1806 948
rect -1854 941 -1806 945
rect -1854 939 -1846 941
rect -1846 937 -1806 939
rect -1806 935 -1798 937
rect -1846 932 -1798 935
rect -1846 919 -1806 930
rect -1671 928 -1663 936
rect -1663 920 -1655 928
rect -1854 914 -1680 918
rect -1926 902 -1892 905
rect -1671 902 -1663 908
rect -1642 902 -1637 948
rect -1619 902 -1614 948
rect -1530 902 -1526 948
rect -1506 902 -1502 948
rect -1482 902 -1478 948
rect -1458 902 -1454 948
rect -1434 902 -1430 948
rect -1410 902 -1406 948
rect -1386 902 -1382 948
rect -1362 902 -1358 948
rect -1338 902 -1334 948
rect -1314 902 -1310 948
rect -1290 902 -1286 948
rect -1266 902 -1262 948
rect -1242 902 -1238 948
rect -1218 902 -1214 948
rect -1194 902 -1190 948
rect -1170 902 -1166 948
rect -1146 902 -1142 948
rect -1122 902 -1118 948
rect -1098 902 -1094 948
rect -1074 902 -1070 948
rect -1050 902 -1046 948
rect -1026 902 -1022 948
rect -1002 902 -998 948
rect -978 902 -974 948
rect -954 902 -950 948
rect -930 902 -926 948
rect -906 902 -902 948
rect -882 902 -878 948
rect -858 902 -854 948
rect -834 902 -830 948
rect -810 902 -806 948
rect -786 902 -782 948
rect -779 947 -765 948
rect -762 923 -755 971
rect -762 902 -758 923
rect -738 902 -734 996
rect -714 902 -710 996
rect -690 902 -686 996
rect -666 902 -662 996
rect -642 902 -638 996
rect -618 902 -614 996
rect -594 902 -590 996
rect -570 902 -566 996
rect -546 902 -542 996
rect -522 902 -518 996
rect -509 989 -504 996
rect -499 975 -494 989
rect -498 902 -494 975
rect -474 947 -470 996
rect -474 902 -467 947
rect -450 902 -446 996
rect -426 902 -422 996
rect -402 902 -398 996
rect -378 902 -374 996
rect -354 902 -350 996
rect -330 902 -326 996
rect -306 902 -302 996
rect -282 902 -278 996
rect -258 902 -254 996
rect -234 902 -230 996
rect -210 902 -206 996
rect -186 902 -182 996
rect -162 902 -158 996
rect -138 902 -134 996
rect -114 902 -110 996
rect -90 902 -86 996
rect -66 902 -62 996
rect -42 902 -38 996
rect -18 902 -14 996
rect 6 902 10 996
rect 30 902 34 996
rect 54 902 58 996
rect 78 902 82 996
rect 102 902 106 996
rect 115 941 120 951
rect 126 941 130 996
rect 150 974 157 995
rect 174 974 178 996
rect 198 974 202 996
rect 222 974 226 996
rect 246 974 250 996
rect 270 975 274 996
rect 259 974 293 975
rect 133 972 293 974
rect 133 971 147 972
rect 150 971 157 972
rect 125 927 130 941
rect 115 917 120 927
rect 125 903 130 917
rect 126 902 130 903
rect 150 902 154 971
rect 174 902 178 972
rect 198 902 202 972
rect 222 903 226 972
rect 211 902 245 903
rect -2393 900 245 902
rect -2371 878 -2366 900
rect -2348 878 -2343 900
rect -2325 896 -2317 900
rect -2325 880 -2320 896
rect -2317 892 -2309 896
rect -2309 880 -2301 892
rect -2109 883 -2079 890
rect -2000 889 -1992 900
rect -1671 896 -1663 900
rect -1846 892 -1806 894
rect -1663 892 -1655 896
rect -2009 886 -1992 889
rect -1854 886 -1806 890
rect -2071 883 -1992 886
rect -1983 883 -1806 886
rect -2009 880 -1992 883
rect -2325 878 -2317 880
rect -2033 878 -1992 880
rect -1846 879 -1806 881
rect -1655 880 -1647 892
rect -1864 878 -1796 879
rect -1671 878 -1663 880
rect -1642 878 -1637 900
rect -1619 878 -1614 900
rect -1530 878 -1526 900
rect -1506 878 -1502 900
rect -1482 878 -1478 900
rect -1458 878 -1454 900
rect -1434 878 -1430 900
rect -1410 878 -1406 900
rect -1386 878 -1382 900
rect -1362 878 -1358 900
rect -1338 878 -1334 900
rect -1314 878 -1310 900
rect -1290 878 -1286 900
rect -1266 878 -1262 900
rect -1242 878 -1238 900
rect -1218 878 -1214 900
rect -1194 878 -1190 900
rect -1170 878 -1166 900
rect -1146 878 -1142 900
rect -1122 878 -1118 900
rect -1098 878 -1094 900
rect -1074 878 -1070 900
rect -1050 878 -1046 900
rect -1026 878 -1022 900
rect -1002 878 -998 900
rect -978 878 -974 900
rect -954 878 -950 900
rect -930 878 -926 900
rect -906 878 -902 900
rect -882 878 -878 900
rect -858 878 -854 900
rect -834 878 -830 900
rect -810 878 -806 900
rect -786 878 -782 900
rect -762 878 -758 900
rect -738 878 -734 900
rect -714 878 -710 900
rect -690 878 -686 900
rect -666 878 -662 900
rect -642 878 -638 900
rect -618 878 -614 900
rect -594 878 -590 900
rect -570 878 -566 900
rect -546 878 -542 900
rect -522 878 -518 900
rect -498 878 -494 900
rect -491 899 -477 900
rect -474 899 -467 900
rect -474 878 -470 899
rect -450 878 -446 900
rect -426 878 -422 900
rect -402 878 -398 900
rect -378 878 -374 900
rect -354 878 -350 900
rect -330 878 -326 900
rect -306 878 -302 900
rect -282 878 -278 900
rect -258 878 -254 900
rect -234 878 -230 900
rect -210 878 -206 900
rect -186 878 -182 900
rect -162 878 -158 900
rect -138 878 -134 900
rect -114 878 -110 900
rect -90 878 -86 900
rect -66 878 -62 900
rect -42 879 -38 900
rect -53 878 -19 879
rect -2393 876 -19 878
rect -2371 854 -2366 876
rect -2348 854 -2343 876
rect -2325 868 -2317 876
rect -2079 873 -2035 876
rect -2013 874 -1992 876
rect -2000 873 -1992 874
rect -1904 873 -1798 876
rect -2101 869 -2009 873
rect -2023 868 -2009 869
rect -2000 871 -1798 873
rect -2000 869 -1854 871
rect -1846 869 -1798 871
rect -2325 854 -2320 868
rect -2317 864 -2309 868
rect -2309 854 -2301 864
rect -2109 856 -2101 863
rect -2023 859 -2021 868
rect -2000 859 -1992 869
rect -1671 868 -1663 876
rect -1846 865 -1806 867
rect -1663 864 -1655 868
rect -1854 859 -1806 863
rect -2071 856 -1806 859
rect -2074 854 -2031 856
rect -2000 854 -1992 856
rect -1655 854 -1647 864
rect -1642 854 -1637 876
rect -1619 854 -1614 876
rect -1530 854 -1526 876
rect -1506 854 -1502 876
rect -1482 854 -1478 876
rect -1458 854 -1454 876
rect -1434 854 -1430 876
rect -1410 854 -1406 876
rect -1386 854 -1382 876
rect -1362 854 -1358 876
rect -1338 854 -1334 876
rect -1314 854 -1310 876
rect -1290 854 -1286 876
rect -1266 854 -1262 876
rect -1242 854 -1238 876
rect -1218 854 -1214 876
rect -1194 854 -1190 876
rect -1170 854 -1166 876
rect -1146 854 -1142 876
rect -1122 854 -1118 876
rect -1098 854 -1094 876
rect -1074 854 -1070 876
rect -1050 854 -1046 876
rect -1026 854 -1022 876
rect -1002 854 -998 876
rect -978 854 -974 876
rect -954 854 -950 876
rect -930 854 -926 876
rect -906 854 -902 876
rect -882 854 -878 876
rect -858 854 -854 876
rect -834 854 -830 876
rect -810 854 -806 876
rect -786 854 -782 876
rect -762 854 -758 876
rect -738 854 -734 876
rect -714 854 -710 876
rect -690 854 -686 876
rect -666 854 -662 876
rect -642 854 -638 876
rect -618 854 -614 876
rect -594 854 -590 876
rect -570 854 -566 876
rect -546 854 -542 876
rect -522 854 -518 876
rect -498 854 -494 876
rect -474 854 -470 876
rect -450 854 -446 876
rect -426 854 -422 876
rect -402 854 -398 876
rect -378 854 -374 876
rect -354 854 -350 876
rect -330 854 -326 876
rect -306 854 -302 876
rect -282 855 -278 876
rect -293 854 -259 855
rect -2393 852 -259 854
rect -2371 806 -2366 852
rect -2348 806 -2343 852
rect -2325 840 -2317 852
rect -2074 849 -2071 852
rect -2101 842 -2071 849
rect -2325 820 -2320 840
rect -2317 836 -2309 840
rect -2064 838 -2061 846
rect -2325 812 -2317 820
rect -2101 815 -2071 818
rect -2325 806 -2320 812
rect -2317 806 -2309 812
rect -2000 810 -1992 852
rect -1846 851 -1806 852
rect -1846 842 -1798 849
rect -1671 840 -1663 852
rect -1846 838 -1806 840
rect -1663 836 -1655 840
rect -1854 824 -1680 828
rect -1846 815 -1798 818
rect -2079 809 -2043 810
rect -2007 809 -1991 810
rect -2079 808 -2071 809
rect -2079 806 -2029 808
rect -2011 806 -1991 809
rect -1846 807 -1806 813
rect -1671 812 -1663 820
rect -1864 806 -1796 807
rect -1663 806 -1655 812
rect -1642 806 -1637 852
rect -1619 806 -1614 852
rect -1530 806 -1526 852
rect -1506 806 -1502 852
rect -1482 806 -1478 852
rect -1458 806 -1454 852
rect -1434 806 -1430 852
rect -1410 806 -1406 852
rect -1386 806 -1382 852
rect -1362 806 -1358 852
rect -1338 806 -1334 852
rect -1325 821 -1320 831
rect -1314 821 -1310 852
rect -1315 807 -1310 821
rect -1325 806 -1291 807
rect -1290 806 -1286 852
rect -1266 806 -1262 852
rect -1242 806 -1238 852
rect -1218 807 -1214 852
rect -1229 806 -1195 807
rect -2393 804 -1195 806
rect -2371 758 -2366 804
rect -2348 758 -2343 804
rect -2325 792 -2320 804
rect -2079 802 -2071 804
rect -2072 800 -2071 802
rect -2109 795 -2101 800
rect -2101 793 -2079 795
rect -2069 793 -2068 800
rect -2325 784 -2317 792
rect -2079 788 -2071 793
rect -2325 764 -2320 784
rect -2317 776 -2309 784
rect -2074 779 -2071 788
rect -2069 784 -2068 788
rect -2109 770 -2079 773
rect -2325 758 -2317 764
rect -2000 758 -1992 804
rect -1846 802 -1806 804
rect -1854 797 -1806 801
rect -1854 795 -1846 797
rect -1846 793 -1806 795
rect -1806 791 -1798 793
rect -1846 788 -1798 791
rect -1846 775 -1806 786
rect -1671 784 -1663 792
rect -1663 776 -1655 784
rect -1854 770 -1680 774
rect -1671 758 -1663 764
rect -1642 758 -1637 804
rect -1619 758 -1614 804
rect -1530 758 -1526 804
rect -1506 758 -1502 804
rect -1482 758 -1478 804
rect -1458 758 -1454 804
rect -1434 758 -1430 804
rect -1410 759 -1406 804
rect -1421 758 -1387 759
rect -2393 756 -1387 758
rect -2371 734 -2366 756
rect -2348 734 -2343 756
rect -2325 748 -2317 756
rect -2325 734 -2320 748
rect -2309 736 -2301 748
rect -2092 739 -2062 744
rect -2000 736 -1992 756
rect -2317 734 -2309 736
rect -2000 734 -1983 736
rect -1906 734 -1904 756
rect -1806 748 -1680 754
rect -1671 748 -1663 756
rect -1854 739 -1806 744
rect -1846 734 -1806 737
rect -1655 736 -1647 748
rect -1663 734 -1655 736
rect -1642 734 -1637 756
rect -1619 734 -1614 756
rect -1530 734 -1526 756
rect -1506 734 -1502 756
rect -1482 734 -1478 756
rect -1458 734 -1454 756
rect -1434 734 -1430 756
rect -1421 749 -1416 756
rect -1410 749 -1406 756
rect -1411 735 -1406 749
rect -1386 734 -1382 804
rect -1362 734 -1358 804
rect -1338 734 -1334 804
rect -1325 797 -1320 804
rect -1315 783 -1310 797
rect -1314 734 -1310 783
rect -1290 755 -1286 804
rect -2393 732 -1293 734
rect -2371 710 -2366 732
rect -2348 710 -2343 732
rect -2325 720 -2317 732
rect -2071 728 -2062 732
rect -2013 730 -1983 732
rect -2000 729 -1983 730
rect -2325 710 -2320 720
rect -2309 710 -2301 720
rect -2100 719 -2092 726
rect -2064 724 -2062 727
rect -2061 719 -2059 724
rect -2071 714 -2062 719
rect -2071 712 -2026 714
rect -2066 710 -2012 712
rect -2000 710 -1992 729
rect -1906 727 -1904 732
rect -1846 728 -1806 732
rect -1846 721 -1798 726
rect -1806 719 -1798 721
rect -1671 720 -1663 732
rect -1854 717 -1846 719
rect -1854 712 -1806 717
rect -1864 710 -1796 711
rect -1655 710 -1647 720
rect -1642 710 -1637 732
rect -1619 710 -1614 732
rect -1530 710 -1526 732
rect -1506 710 -1502 732
rect -1482 710 -1478 732
rect -1458 710 -1454 732
rect -1434 710 -1430 732
rect -1386 710 -1382 732
rect -1362 710 -1358 732
rect -1338 710 -1334 732
rect -1314 710 -1310 732
rect -1307 731 -1293 732
rect -1290 710 -1283 755
rect -1266 710 -1262 804
rect -1242 710 -1238 804
rect -1229 797 -1224 804
rect -1218 797 -1214 804
rect -1219 783 -1214 797
rect -1229 782 -1195 783
rect -1194 782 -1190 852
rect -1170 782 -1166 852
rect -1146 782 -1142 852
rect -1122 782 -1118 852
rect -1098 782 -1094 852
rect -1074 782 -1070 852
rect -1050 782 -1046 852
rect -1026 782 -1022 852
rect -1002 782 -998 852
rect -978 782 -974 852
rect -954 782 -950 852
rect -930 782 -926 852
rect -906 782 -902 852
rect -882 782 -878 852
rect -858 782 -854 852
rect -834 782 -830 852
rect -810 782 -806 852
rect -786 782 -782 852
rect -762 782 -758 852
rect -738 782 -734 852
rect -714 782 -710 852
rect -690 782 -686 852
rect -666 782 -662 852
rect -642 782 -638 852
rect -618 782 -614 852
rect -594 782 -590 852
rect -570 782 -566 852
rect -546 782 -542 852
rect -522 782 -518 852
rect -498 782 -494 852
rect -474 782 -470 852
rect -450 782 -446 852
rect -426 782 -422 852
rect -402 782 -398 852
rect -378 782 -374 852
rect -354 782 -350 852
rect -330 782 -326 852
rect -306 782 -302 852
rect -293 845 -288 852
rect -282 845 -278 852
rect -283 831 -278 845
rect -293 821 -288 831
rect -283 807 -278 821
rect -282 782 -278 807
rect -258 782 -254 876
rect -234 782 -230 876
rect -210 782 -206 876
rect -186 782 -182 876
rect -162 782 -158 876
rect -138 782 -134 876
rect -114 782 -110 876
rect -90 782 -86 876
rect -66 782 -62 876
rect -53 869 -48 876
rect -42 869 -38 876
rect -43 855 -38 869
rect -53 854 -19 855
rect -18 854 -14 900
rect 6 854 10 900
rect 30 854 34 900
rect 54 854 58 900
rect 78 854 82 900
rect 102 854 106 900
rect 126 854 130 900
rect 150 875 154 900
rect -53 852 147 854
rect -53 845 -48 852
rect -43 831 -38 845
rect -42 782 -38 831
rect -18 803 -14 852
rect -1229 780 -21 782
rect -1229 773 -1224 780
rect -1219 759 -1214 773
rect -1218 710 -1214 759
rect -1194 731 -1190 780
rect -2393 708 -1197 710
rect -2371 662 -2366 708
rect -2348 662 -2343 708
rect -2325 704 -2320 708
rect -2317 704 -2309 708
rect -2325 692 -2317 704
rect -2066 703 -2062 708
rect -2147 700 -2134 702
rect -2292 694 -2071 700
rect -2325 672 -2320 692
rect -2092 678 -2062 680
rect -2094 674 -2062 678
rect -2325 662 -2317 672
rect -2095 664 -2084 668
rect -2000 665 -1992 708
rect -1846 701 -1806 708
rect -1663 704 -1655 708
rect -1846 694 -1680 700
rect -1671 692 -1663 704
rect -1854 678 -1806 680
rect -1854 674 -1680 678
rect -2119 662 -2069 664
rect -2054 662 -1892 665
rect -1671 662 -1663 672
rect -1642 662 -1637 708
rect -1619 662 -1614 708
rect -1530 662 -1526 708
rect -1506 662 -1502 708
rect -1482 662 -1478 708
rect -1458 662 -1454 708
rect -1434 662 -1430 708
rect -1421 677 -1416 687
rect -1386 683 -1382 708
rect -1411 663 -1406 677
rect -1397 673 -1389 677
rect -1403 663 -1397 673
rect -1421 662 -1389 663
rect -2393 660 -1389 662
rect -2371 638 -2366 660
rect -2348 638 -2343 660
rect -2325 656 -2317 660
rect -2325 640 -2320 656
rect -2309 644 -2301 656
rect -2095 654 -2084 660
rect -2054 659 -1906 660
rect -2054 658 -2036 659
rect -2084 652 -2079 654
rect -2317 640 -2309 644
rect -2092 643 -2079 650
rect -2000 646 -1992 659
rect -1920 658 -1906 659
rect -1671 656 -1663 660
rect -1846 652 -1806 654
rect -1854 646 -1806 650
rect -2054 643 -1982 646
rect -1966 643 -1806 646
rect -1655 644 -1647 656
rect -2003 640 -1992 643
rect -1904 641 -1902 643
rect -1854 641 -1846 643
rect -2325 638 -2317 640
rect -2033 638 -1992 640
rect -1854 639 -1806 641
rect -1663 640 -1655 644
rect -1864 638 -1796 639
rect -1671 638 -1663 640
rect -1642 638 -1637 660
rect -1619 638 -1614 660
rect -1530 638 -1526 660
rect -1506 638 -1502 660
rect -1482 638 -1478 660
rect -1458 638 -1454 660
rect -1434 638 -1430 660
rect -1421 653 -1416 660
rect -1410 653 -1406 660
rect -1403 659 -1389 660
rect -1386 659 -1379 683
rect -1411 639 -1406 653
rect -1362 638 -1358 708
rect -1338 638 -1334 708
rect -1314 638 -1310 708
rect -1307 707 -1293 708
rect -1290 707 -1283 708
rect -1290 638 -1286 707
rect -1266 638 -1262 708
rect -1242 638 -1238 708
rect -1218 638 -1214 708
rect -1211 707 -1197 708
rect -1194 686 -1187 731
rect -1170 686 -1166 780
rect -1146 686 -1142 780
rect -1122 686 -1118 780
rect -1098 686 -1094 780
rect -1074 686 -1070 780
rect -1050 686 -1046 780
rect -1026 686 -1022 780
rect -1002 686 -998 780
rect -978 686 -974 780
rect -954 686 -950 780
rect -930 686 -926 780
rect -906 686 -902 780
rect -893 701 -888 711
rect -882 701 -878 780
rect -883 687 -878 701
rect -858 686 -854 780
rect -834 686 -830 780
rect -810 686 -806 780
rect -786 686 -782 780
rect -773 725 -768 735
rect -762 725 -758 780
rect -763 711 -758 725
rect -773 701 -768 711
rect -763 687 -758 701
rect -762 686 -758 687
rect -738 686 -734 780
rect -714 686 -710 780
rect -690 686 -686 780
rect -666 686 -662 780
rect -642 686 -638 780
rect -618 686 -614 780
rect -594 686 -590 780
rect -570 686 -566 780
rect -546 686 -542 780
rect -522 686 -518 780
rect -498 686 -494 780
rect -474 686 -470 780
rect -450 686 -446 780
rect -426 686 -422 780
rect -402 686 -398 780
rect -378 686 -374 780
rect -354 686 -350 780
rect -330 686 -326 780
rect -306 686 -302 780
rect -282 686 -278 780
rect -258 779 -254 780
rect -258 731 -251 779
rect -258 686 -254 731
rect -234 686 -230 780
rect -210 686 -206 780
rect -186 686 -182 780
rect -162 686 -158 780
rect -138 686 -134 780
rect -114 686 -110 780
rect -90 686 -86 780
rect -66 686 -62 780
rect -42 686 -38 780
rect -35 779 -21 780
rect -18 755 -11 803
rect -18 686 -14 755
rect 6 686 10 852
rect 30 686 34 852
rect 54 686 58 852
rect 78 686 82 852
rect 102 686 106 852
rect 126 686 130 852
rect 133 851 147 852
rect 150 830 157 875
rect 174 830 178 900
rect 198 830 202 900
rect 211 893 216 900
rect 222 893 226 900
rect 221 879 226 893
rect 211 878 245 879
rect 246 878 250 972
rect 259 965 264 972
rect 270 965 274 972
rect 269 951 274 965
rect 259 941 264 951
rect 269 927 274 941
rect 270 878 274 927
rect 294 899 298 996
rect 211 876 291 878
rect 211 869 216 876
rect 221 855 226 869
rect 222 830 226 855
rect 246 830 250 876
rect 270 830 274 876
rect 277 875 291 876
rect 294 854 301 899
rect 318 854 322 996
rect 342 854 346 996
rect 366 854 370 996
rect 390 854 394 996
rect 414 854 418 996
rect 438 854 442 996
rect 462 854 466 996
rect 486 854 490 996
rect 510 854 514 996
rect 534 854 538 996
rect 558 854 562 996
rect 582 854 586 996
rect 606 854 610 996
rect 630 854 634 996
rect 654 854 658 996
rect 678 854 682 996
rect 702 854 706 996
rect 726 854 730 996
rect 750 854 754 996
rect 774 854 778 996
rect 798 854 802 996
rect 822 854 826 996
rect 846 854 850 996
rect 870 854 874 996
rect 894 854 898 996
rect 901 995 915 996
rect 918 995 925 1019
rect 918 950 925 971
rect 942 950 946 1116
rect 966 1070 973 1091
rect 990 1070 994 1116
rect 1014 1070 1018 1116
rect 1038 1070 1042 1116
rect 1062 1070 1066 1116
rect 1086 1070 1090 1116
rect 1110 1070 1114 1116
rect 1134 1070 1138 1116
rect 1182 1070 1186 1116
rect 1206 1070 1210 1116
rect 1230 1070 1234 1116
rect 1254 1070 1258 1116
rect 1278 1070 1282 1116
rect 1302 1070 1306 1116
rect 1326 1070 1330 1116
rect 1350 1070 1354 1116
rect 1374 1070 1378 1116
rect 1398 1070 1402 1116
rect 1422 1070 1426 1116
rect 1446 1070 1450 1116
rect 1470 1070 1474 1116
rect 1494 1070 1498 1116
rect 1518 1070 1522 1116
rect 1542 1070 1546 1116
rect 1566 1070 1570 1116
rect 1590 1071 1594 1116
rect 1603 1109 1608 1116
rect 1614 1109 1618 1116
rect 1613 1095 1618 1109
rect 1579 1070 1613 1071
rect 949 1068 1613 1070
rect 949 1067 963 1068
rect 966 1067 973 1068
rect 966 950 970 1067
rect 990 950 994 1068
rect 1014 950 1018 1068
rect 1038 950 1042 1068
rect 1062 950 1066 1068
rect 1086 950 1090 1068
rect 1110 950 1114 1068
rect 1134 950 1138 1068
rect 1158 1046 1165 1067
rect 1182 1046 1186 1068
rect 1206 1046 1210 1068
rect 1230 1046 1234 1068
rect 1254 1046 1258 1068
rect 1278 1046 1282 1068
rect 1302 1046 1306 1068
rect 1326 1046 1330 1068
rect 1350 1046 1354 1068
rect 1374 1046 1378 1068
rect 1398 1046 1402 1068
rect 1422 1046 1426 1068
rect 1446 1046 1450 1068
rect 1470 1046 1474 1068
rect 1494 1046 1498 1068
rect 1518 1046 1522 1068
rect 1542 1046 1546 1068
rect 1566 1047 1570 1068
rect 1579 1061 1584 1068
rect 1590 1061 1594 1068
rect 1589 1047 1594 1061
rect 1555 1046 1589 1047
rect 1141 1044 1589 1046
rect 1141 1043 1155 1044
rect 1158 1043 1165 1044
rect 1158 950 1162 1043
rect 1182 950 1186 1044
rect 1206 950 1210 1044
rect 1230 950 1234 1044
rect 1254 950 1258 1044
rect 1278 950 1282 1044
rect 1302 950 1306 1044
rect 1326 950 1330 1044
rect 1350 950 1354 1044
rect 1374 950 1378 1044
rect 1398 950 1402 1044
rect 1422 950 1426 1044
rect 1446 950 1450 1044
rect 1470 950 1474 1044
rect 1483 989 1488 999
rect 1494 989 1498 1044
rect 1493 975 1498 989
rect 1483 974 1517 975
rect 1518 974 1522 1044
rect 1542 975 1546 1044
rect 1555 1037 1560 1044
rect 1566 1037 1570 1044
rect 1565 1023 1570 1037
rect 1531 974 1565 975
rect 1483 972 1565 974
rect 1483 965 1488 972
rect 1493 951 1498 965
rect 1518 951 1522 972
rect 1531 965 1536 972
rect 1542 965 1546 972
rect 1541 951 1546 965
rect 1494 950 1498 951
rect 1507 950 1541 951
rect 901 948 1541 950
rect 901 947 915 948
rect 918 947 925 948
rect 918 854 922 947
rect 942 854 946 948
rect 966 854 970 948
rect 990 854 994 948
rect 1014 854 1018 948
rect 1038 854 1042 948
rect 1062 854 1066 948
rect 1086 854 1090 948
rect 1110 854 1114 948
rect 1134 854 1138 948
rect 1158 854 1162 948
rect 1182 854 1186 948
rect 1206 854 1210 948
rect 1230 854 1234 948
rect 1254 854 1258 948
rect 1278 854 1282 948
rect 1302 854 1306 948
rect 1326 854 1330 948
rect 1350 854 1354 948
rect 1374 854 1378 948
rect 1398 854 1402 948
rect 1422 854 1426 948
rect 1446 855 1450 948
rect 1459 869 1464 879
rect 1470 869 1474 948
rect 1483 917 1488 927
rect 1494 917 1498 948
rect 1507 941 1512 948
rect 1518 941 1522 948
rect 1517 927 1522 941
rect 1493 903 1498 917
rect 1507 913 1515 917
rect 1501 903 1507 913
rect 1469 855 1474 869
rect 1435 854 1469 855
rect 277 852 1469 854
rect 277 851 291 852
rect 294 851 301 852
rect 294 830 298 851
rect 318 830 322 852
rect 342 830 346 852
rect 366 830 370 852
rect 390 830 394 852
rect 414 830 418 852
rect 438 830 442 852
rect 462 830 466 852
rect 486 830 490 852
rect 510 830 514 852
rect 534 830 538 852
rect 558 830 562 852
rect 582 830 586 852
rect 606 830 610 852
rect 630 830 634 852
rect 654 830 658 852
rect 678 830 682 852
rect 702 830 706 852
rect 726 830 730 852
rect 750 830 754 852
rect 774 830 778 852
rect 798 830 802 852
rect 822 830 826 852
rect 846 830 850 852
rect 870 830 874 852
rect 894 830 898 852
rect 918 830 922 852
rect 942 830 946 852
rect 966 830 970 852
rect 990 830 994 852
rect 1014 830 1018 852
rect 1038 830 1042 852
rect 1062 830 1066 852
rect 1086 830 1090 852
rect 1110 830 1114 852
rect 1134 830 1138 852
rect 1158 830 1162 852
rect 1182 830 1186 852
rect 1206 830 1210 852
rect 1230 830 1234 852
rect 1254 830 1258 852
rect 1278 830 1282 852
rect 1302 830 1306 852
rect 1326 830 1330 852
rect 1350 830 1354 852
rect 1374 830 1378 852
rect 1398 830 1402 852
rect 1422 831 1426 852
rect 1435 845 1440 852
rect 1446 845 1450 852
rect 1445 831 1450 845
rect 1411 830 1445 831
rect 133 828 1445 830
rect 133 827 147 828
rect 150 827 157 828
rect 150 686 154 827
rect 174 686 178 828
rect 198 686 202 828
rect 222 686 226 828
rect 246 827 250 828
rect 246 782 253 827
rect 270 782 274 828
rect 294 782 298 828
rect 318 782 322 828
rect 342 782 346 828
rect 366 782 370 828
rect 390 782 394 828
rect 414 782 418 828
rect 438 782 442 828
rect 462 782 466 828
rect 486 782 490 828
rect 510 782 514 828
rect 534 782 538 828
rect 558 782 562 828
rect 582 782 586 828
rect 606 782 610 828
rect 630 782 634 828
rect 654 782 658 828
rect 678 782 682 828
rect 702 782 706 828
rect 726 782 730 828
rect 750 782 754 828
rect 774 782 778 828
rect 798 782 802 828
rect 822 782 826 828
rect 846 782 850 828
rect 870 782 874 828
rect 894 782 898 828
rect 918 782 922 828
rect 942 782 946 828
rect 966 782 970 828
rect 990 782 994 828
rect 1014 782 1018 828
rect 1038 782 1042 828
rect 1062 782 1066 828
rect 1086 782 1090 828
rect 1110 782 1114 828
rect 1134 782 1138 828
rect 1158 782 1162 828
rect 1182 782 1186 828
rect 1206 782 1210 828
rect 1230 782 1234 828
rect 1254 782 1258 828
rect 1278 782 1282 828
rect 1302 782 1306 828
rect 1326 782 1330 828
rect 1350 782 1354 828
rect 1374 782 1378 828
rect 1398 783 1402 828
rect 1411 821 1416 828
rect 1422 821 1426 828
rect 1421 807 1426 821
rect 1387 782 1421 783
rect 229 780 1421 782
rect 229 779 243 780
rect 246 779 253 780
rect 246 686 250 779
rect 270 686 274 780
rect 294 686 298 780
rect 318 686 322 780
rect 342 686 346 780
rect 366 686 370 780
rect 390 686 394 780
rect 414 686 418 780
rect 438 686 442 780
rect 462 686 466 780
rect 486 686 490 780
rect 510 686 514 780
rect 534 686 538 780
rect 558 686 562 780
rect 582 686 586 780
rect 606 686 610 780
rect 630 686 634 780
rect 654 686 658 780
rect 678 686 682 780
rect 702 686 706 780
rect 726 686 730 780
rect 750 686 754 780
rect 774 686 778 780
rect 798 686 802 780
rect 822 686 826 780
rect 846 686 850 780
rect 870 686 874 780
rect 894 686 898 780
rect 918 686 922 780
rect 942 686 946 780
rect 966 686 970 780
rect 990 686 994 780
rect 1014 686 1018 780
rect 1038 686 1042 780
rect 1062 686 1066 780
rect 1086 686 1090 780
rect 1110 686 1114 780
rect 1134 686 1138 780
rect 1158 686 1162 780
rect 1182 686 1186 780
rect 1206 686 1210 780
rect 1230 686 1234 780
rect 1254 686 1258 780
rect 1278 686 1282 780
rect 1302 686 1306 780
rect 1326 686 1330 780
rect 1350 687 1354 780
rect 1363 701 1368 711
rect 1374 701 1378 780
rect 1387 773 1392 780
rect 1398 773 1402 780
rect 1397 759 1402 773
rect 1373 687 1378 701
rect 1339 686 1373 687
rect -1211 684 1373 686
rect -1211 683 -1197 684
rect -1194 683 -1187 684
rect -1194 638 -1190 683
rect -1170 638 -1166 684
rect -1146 638 -1142 684
rect -1122 638 -1118 684
rect -1098 638 -1094 684
rect -1074 638 -1070 684
rect -1050 638 -1046 684
rect -1026 638 -1022 684
rect -1002 638 -998 684
rect -978 638 -974 684
rect -954 638 -950 684
rect -930 638 -926 684
rect -906 638 -902 684
rect -893 653 -888 663
rect -883 639 -878 653
rect -882 638 -878 639
rect -858 638 -854 684
rect -834 638 -830 684
rect -810 638 -806 684
rect -786 638 -782 684
rect -762 638 -758 684
rect -738 659 -734 684
rect -2393 636 -741 638
rect -2371 614 -2366 636
rect -2348 614 -2343 636
rect -2325 628 -2317 636
rect -2079 633 -2018 636
rect -2003 635 -1966 636
rect -2000 634 -1982 635
rect -2000 633 -1992 634
rect -2084 629 -2009 633
rect -2028 628 -2009 629
rect -2000 629 -1854 633
rect -1846 629 -1798 636
rect -2325 614 -2320 628
rect -2309 616 -2301 628
rect -2028 626 -2018 628
rect -2092 616 -2084 623
rect -2023 619 -2014 626
rect -2000 619 -1992 629
rect -1671 628 -1663 636
rect -1846 625 -1806 627
rect -1854 619 -1806 623
rect -2054 616 -1806 619
rect -1655 616 -1647 628
rect -2317 614 -2309 616
rect -2054 614 -2024 616
rect -2000 614 -1992 616
rect -1663 614 -1655 616
rect -1642 614 -1637 636
rect -1619 614 -1614 636
rect -1530 614 -1526 636
rect -1506 614 -1502 636
rect -1482 614 -1478 636
rect -1458 614 -1454 636
rect -1434 614 -1430 636
rect -1362 614 -1358 636
rect -1338 614 -1334 636
rect -1314 614 -1310 636
rect -1290 614 -1286 636
rect -1266 614 -1262 636
rect -1242 614 -1238 636
rect -1218 614 -1214 636
rect -1194 614 -1190 636
rect -1170 614 -1166 636
rect -1146 614 -1142 636
rect -1122 614 -1118 636
rect -1098 614 -1094 636
rect -1074 614 -1070 636
rect -1050 614 -1046 636
rect -1026 614 -1022 636
rect -1002 614 -998 636
rect -978 614 -974 636
rect -954 614 -950 636
rect -930 615 -926 636
rect -941 614 -907 615
rect -2393 612 -2064 614
rect -2060 612 -907 614
rect -2371 566 -2366 612
rect -2348 566 -2343 612
rect -2325 600 -2317 612
rect -2060 609 -2054 612
rect -2084 602 -2054 609
rect -2050 606 -2044 608
rect -2325 580 -2320 600
rect -2064 598 -2054 602
rect -2325 572 -2317 580
rect -2101 575 -2071 578
rect -2325 566 -2320 572
rect -2317 566 -2309 572
rect -2000 570 -1992 612
rect -1846 611 -1806 612
rect -1846 602 -1798 609
rect -1671 600 -1663 612
rect -1846 598 -1806 600
rect -1854 584 -1680 588
rect -1846 575 -1798 578
rect -2079 569 -2043 570
rect -2007 569 -1991 570
rect -2079 568 -2071 569
rect -2079 566 -2029 568
rect -2011 566 -1991 569
rect -1846 567 -1806 573
rect -1671 572 -1663 580
rect -1864 566 -1796 567
rect -1663 566 -1655 572
rect -1642 566 -1637 612
rect -1619 566 -1614 612
rect -1530 566 -1526 612
rect -1506 566 -1502 612
rect -1482 566 -1478 612
rect -1458 566 -1454 612
rect -1434 566 -1430 612
rect -1386 590 -1379 611
rect -1362 590 -1358 612
rect -1338 590 -1334 612
rect -1314 590 -1310 612
rect -1290 590 -1286 612
rect -1266 590 -1262 612
rect -1242 590 -1238 612
rect -1218 590 -1214 612
rect -1194 590 -1190 612
rect -1170 590 -1166 612
rect -1146 590 -1142 612
rect -1122 590 -1118 612
rect -1098 590 -1094 612
rect -1074 590 -1070 612
rect -1050 590 -1046 612
rect -1026 590 -1022 612
rect -1002 590 -998 612
rect -978 590 -974 612
rect -954 590 -950 612
rect -941 605 -936 612
rect -930 605 -926 612
rect -931 591 -926 605
rect -906 590 -902 636
rect -882 590 -878 636
rect -858 635 -854 636
rect -858 611 -851 635
rect -834 590 -830 636
rect -810 590 -806 636
rect -786 590 -782 636
rect -762 590 -758 636
rect -755 635 -741 636
rect -738 611 -731 659
rect -738 590 -734 611
rect -714 590 -710 684
rect -690 590 -686 684
rect -666 590 -662 684
rect -642 590 -638 684
rect -618 590 -614 684
rect -594 590 -590 684
rect -570 590 -566 684
rect -546 590 -542 684
rect -522 590 -518 684
rect -498 590 -494 684
rect -474 590 -470 684
rect -450 590 -446 684
rect -426 590 -422 684
rect -402 590 -398 684
rect -378 590 -374 684
rect -354 590 -350 684
rect -330 590 -326 684
rect -306 590 -302 684
rect -282 590 -278 684
rect -258 590 -254 684
rect -234 590 -230 684
rect -210 590 -206 684
rect -186 590 -182 684
rect -162 590 -158 684
rect -138 590 -134 684
rect -114 590 -110 684
rect -90 590 -86 684
rect -66 590 -62 684
rect -53 629 -48 639
rect -42 629 -38 684
rect -43 615 -38 629
rect -53 614 -19 615
rect -18 614 -14 684
rect 6 614 10 684
rect 30 614 34 684
rect 54 614 58 684
rect 78 614 82 684
rect 102 614 106 684
rect 126 614 130 684
rect 150 614 154 684
rect 174 614 178 684
rect 198 614 202 684
rect 222 614 226 684
rect 246 614 250 684
rect 270 614 274 684
rect 294 614 298 684
rect 318 614 322 684
rect 342 614 346 684
rect 366 614 370 684
rect 390 614 394 684
rect 414 614 418 684
rect 438 614 442 684
rect 462 614 466 684
rect 486 614 490 684
rect 510 614 514 684
rect 534 614 538 684
rect 558 614 562 684
rect 582 614 586 684
rect 606 614 610 684
rect 630 614 634 684
rect 654 614 658 684
rect 678 614 682 684
rect 702 614 706 684
rect 726 614 730 684
rect 750 614 754 684
rect 774 614 778 684
rect 798 614 802 684
rect 822 614 826 684
rect 846 614 850 684
rect 870 614 874 684
rect 894 614 898 684
rect 918 614 922 684
rect 942 614 946 684
rect 966 614 970 684
rect 990 614 994 684
rect 1014 614 1018 684
rect 1038 614 1042 684
rect 1062 614 1066 684
rect 1086 614 1090 684
rect 1110 614 1114 684
rect 1134 614 1138 684
rect 1158 614 1162 684
rect 1182 614 1186 684
rect 1206 614 1210 684
rect 1230 614 1234 684
rect 1254 614 1258 684
rect 1278 614 1282 684
rect 1302 615 1306 684
rect 1315 653 1320 663
rect 1326 653 1330 684
rect 1339 677 1344 684
rect 1350 677 1354 684
rect 1349 663 1354 677
rect 1325 639 1330 653
rect 1291 614 1325 615
rect -53 612 1325 614
rect -53 605 -48 612
rect -43 591 -38 605
rect -42 590 -38 591
rect -18 590 -14 612
rect 6 590 10 612
rect 30 590 34 612
rect 54 590 58 612
rect 78 590 82 612
rect 102 590 106 612
rect 126 590 130 612
rect 150 590 154 612
rect 174 590 178 612
rect 198 590 202 612
rect 222 590 226 612
rect 246 590 250 612
rect 270 591 274 612
rect 259 590 293 591
rect -1403 588 293 590
rect -1403 587 -1389 588
rect -2393 564 -1389 566
rect -2371 518 -2366 564
rect -2348 518 -2343 564
rect -2325 552 -2320 564
rect -2079 562 -2071 564
rect -2072 560 -2071 562
rect -2109 555 -2101 560
rect -2101 553 -2079 555
rect -2069 553 -2068 560
rect -2325 544 -2317 552
rect -2079 548 -2071 553
rect -2325 524 -2320 544
rect -2317 536 -2309 544
rect -2074 539 -2071 548
rect -2069 544 -2068 548
rect -2109 530 -2079 533
rect -2325 518 -2317 524
rect -2000 518 -1992 564
rect -1846 562 -1806 564
rect -1854 557 -1806 561
rect -1854 555 -1846 557
rect -1846 553 -1806 555
rect -1806 551 -1798 553
rect -1846 548 -1798 551
rect -1846 535 -1806 546
rect -1671 544 -1663 552
rect -1663 536 -1655 544
rect -1854 530 -1680 534
rect -1671 518 -1663 524
rect -1642 518 -1637 564
rect -1619 518 -1614 564
rect -1530 518 -1526 564
rect -1506 518 -1502 564
rect -1482 518 -1478 564
rect -1458 518 -1454 564
rect -1434 518 -1430 564
rect -1403 563 -1389 564
rect -1386 563 -1379 588
rect -1421 542 -1387 543
rect -1362 542 -1358 588
rect -1338 542 -1334 588
rect -1314 542 -1310 588
rect -1290 542 -1286 588
rect -1266 542 -1262 588
rect -1242 542 -1238 588
rect -1218 542 -1214 588
rect -1194 542 -1190 588
rect -1170 542 -1166 588
rect -1146 542 -1142 588
rect -1122 542 -1118 588
rect -1098 542 -1094 588
rect -1074 542 -1070 588
rect -1050 542 -1046 588
rect -1026 542 -1022 588
rect -1002 542 -998 588
rect -978 542 -974 588
rect -954 542 -950 588
rect -906 542 -902 588
rect -882 542 -878 588
rect -858 566 -851 587
rect -834 566 -830 588
rect -810 566 -806 588
rect -786 566 -782 588
rect -762 566 -758 588
rect -738 566 -734 588
rect -714 566 -710 588
rect -690 566 -686 588
rect -666 566 -662 588
rect -642 566 -638 588
rect -618 566 -614 588
rect -594 566 -590 588
rect -570 566 -566 588
rect -546 566 -542 588
rect -522 566 -518 588
rect -498 566 -494 588
rect -474 566 -470 588
rect -450 566 -446 588
rect -426 566 -422 588
rect -402 566 -398 588
rect -378 566 -374 588
rect -354 566 -350 588
rect -330 566 -326 588
rect -306 566 -302 588
rect -282 566 -278 588
rect -258 566 -254 588
rect -234 566 -230 588
rect -210 566 -206 588
rect -186 566 -182 588
rect -162 566 -158 588
rect -138 566 -134 588
rect -114 566 -110 588
rect -90 566 -86 588
rect -66 566 -62 588
rect -42 566 -38 588
rect -18 566 -14 588
rect 6 566 10 588
rect 30 566 34 588
rect 54 566 58 588
rect 78 566 82 588
rect 102 566 106 588
rect 126 566 130 588
rect 150 566 154 588
rect 174 566 178 588
rect 198 566 202 588
rect 222 566 226 588
rect 246 566 250 588
rect 259 581 264 588
rect 270 581 274 588
rect 269 567 274 581
rect 294 566 298 612
rect 318 566 322 612
rect 342 566 346 612
rect 366 566 370 612
rect 390 566 394 612
rect 414 566 418 612
rect 438 566 442 612
rect 462 566 466 612
rect 486 566 490 612
rect 510 566 514 612
rect 534 566 538 612
rect 558 566 562 612
rect 582 566 586 612
rect 606 566 610 612
rect 630 566 634 612
rect 654 566 658 612
rect 678 566 682 612
rect 702 566 706 612
rect 726 566 730 612
rect 750 566 754 612
rect 774 566 778 612
rect 798 566 802 612
rect 822 566 826 612
rect 846 566 850 612
rect 870 566 874 612
rect 894 566 898 612
rect 918 566 922 612
rect 942 566 946 612
rect 966 566 970 612
rect 990 566 994 612
rect 1014 566 1018 612
rect 1038 566 1042 612
rect 1062 566 1066 612
rect 1086 566 1090 612
rect 1110 566 1114 612
rect 1134 566 1138 612
rect 1158 567 1162 612
rect 1147 566 1181 567
rect -875 564 1181 566
rect -875 563 -861 564
rect -858 563 -851 564
rect -858 542 -854 563
rect -834 542 -830 564
rect -810 542 -806 564
rect -786 542 -782 564
rect -762 542 -758 564
rect -738 542 -734 564
rect -714 542 -710 564
rect -690 542 -686 564
rect -666 542 -662 564
rect -642 542 -638 564
rect -618 542 -614 564
rect -594 542 -590 564
rect -570 542 -566 564
rect -546 542 -542 564
rect -522 542 -518 564
rect -498 542 -494 564
rect -474 542 -470 564
rect -450 542 -446 564
rect -426 542 -422 564
rect -402 542 -398 564
rect -378 542 -374 564
rect -354 542 -350 564
rect -330 542 -326 564
rect -306 542 -302 564
rect -282 542 -278 564
rect -258 542 -254 564
rect -234 542 -230 564
rect -210 542 -206 564
rect -186 542 -182 564
rect -162 542 -158 564
rect -138 542 -134 564
rect -114 542 -110 564
rect -90 542 -86 564
rect -66 542 -62 564
rect -42 542 -38 564
rect -18 563 -14 564
rect -1421 540 -21 542
rect -1421 533 -1416 540
rect -1411 519 -1406 533
rect -1410 518 -1406 519
rect -1362 518 -1358 540
rect -1338 518 -1334 540
rect -1314 518 -1310 540
rect -1290 518 -1286 540
rect -1266 518 -1262 540
rect -1242 518 -1238 540
rect -1218 518 -1214 540
rect -1194 518 -1190 540
rect -1170 518 -1166 540
rect -1146 518 -1142 540
rect -1122 518 -1118 540
rect -1098 518 -1094 540
rect -1074 518 -1070 540
rect -1050 518 -1046 540
rect -1026 518 -1022 540
rect -1002 518 -998 540
rect -978 518 -974 540
rect -954 518 -950 540
rect -906 539 -902 540
rect -941 518 -909 519
rect -2393 516 -909 518
rect -2371 494 -2366 516
rect -2348 494 -2343 516
rect -2325 508 -2317 516
rect -2325 494 -2320 508
rect -2309 496 -2301 508
rect -2092 499 -2062 504
rect -2000 496 -1992 516
rect -2317 494 -2309 496
rect -2000 494 -1983 496
rect -1906 494 -1904 516
rect -1806 508 -1680 514
rect -1671 508 -1663 516
rect -1854 499 -1806 504
rect -1846 494 -1806 497
rect -1655 496 -1647 508
rect -1663 494 -1655 496
rect -1642 494 -1637 516
rect -1619 494 -1614 516
rect -1530 494 -1526 516
rect -1506 494 -1502 516
rect -1482 494 -1478 516
rect -1458 494 -1454 516
rect -1434 494 -1430 516
rect -1410 494 -1406 516
rect -1362 494 -1358 516
rect -1338 494 -1334 516
rect -1314 494 -1310 516
rect -1290 494 -1286 516
rect -1266 494 -1262 516
rect -1242 494 -1238 516
rect -1218 494 -1214 516
rect -1194 494 -1190 516
rect -1170 494 -1166 516
rect -1146 494 -1142 516
rect -1122 494 -1118 516
rect -1098 494 -1094 516
rect -1074 494 -1070 516
rect -1050 494 -1046 516
rect -1026 494 -1022 516
rect -1002 494 -998 516
rect -978 494 -974 516
rect -954 494 -950 516
rect -941 509 -936 516
rect -923 515 -909 516
rect -906 515 -899 539
rect -931 495 -926 509
rect -930 494 -926 495
rect -882 494 -878 540
rect -858 494 -854 540
rect -834 494 -830 540
rect -810 494 -806 540
rect -786 494 -782 540
rect -762 495 -758 540
rect -773 494 -739 495
rect -2393 492 -739 494
rect -2371 470 -2366 492
rect -2348 470 -2343 492
rect -2325 480 -2317 492
rect -2071 488 -2062 492
rect -2013 490 -1983 492
rect -2000 489 -1983 490
rect -2325 470 -2320 480
rect -2309 470 -2301 480
rect -2100 479 -2092 486
rect -2064 484 -2062 487
rect -2061 479 -2059 484
rect -2071 474 -2062 479
rect -2071 472 -2026 474
rect -2066 470 -2012 472
rect -2000 470 -1992 489
rect -1906 487 -1904 492
rect -1846 488 -1806 492
rect -1846 481 -1798 486
rect -1806 479 -1798 481
rect -1671 480 -1663 492
rect -1854 477 -1846 479
rect -1854 472 -1806 477
rect -1864 470 -1796 471
rect -1655 470 -1647 480
rect -1642 470 -1637 492
rect -1619 470 -1614 492
rect -1530 470 -1526 492
rect -1506 470 -1502 492
rect -1482 470 -1478 492
rect -1458 470 -1454 492
rect -1434 470 -1430 492
rect -1410 470 -1406 492
rect -1362 470 -1358 492
rect -1338 470 -1334 492
rect -1314 470 -1310 492
rect -1290 470 -1286 492
rect -1266 470 -1262 492
rect -1242 470 -1238 492
rect -1218 470 -1214 492
rect -1194 470 -1190 492
rect -1170 470 -1166 492
rect -1146 470 -1142 492
rect -1122 470 -1118 492
rect -1098 470 -1094 492
rect -1074 470 -1070 492
rect -1050 470 -1046 492
rect -1026 470 -1022 492
rect -1002 470 -998 492
rect -978 470 -974 492
rect -954 470 -950 492
rect -930 470 -926 492
rect -882 470 -878 492
rect -858 470 -854 492
rect -834 470 -830 492
rect -810 470 -806 492
rect -786 470 -782 492
rect -773 485 -768 492
rect -762 485 -758 492
rect -763 471 -758 485
rect -738 470 -734 540
rect -714 470 -710 540
rect -690 470 -686 540
rect -666 470 -662 540
rect -642 470 -638 540
rect -618 470 -614 540
rect -594 470 -590 540
rect -570 470 -566 540
rect -546 470 -542 540
rect -522 470 -518 540
rect -498 470 -494 540
rect -474 470 -470 540
rect -450 470 -446 540
rect -426 470 -422 540
rect -402 470 -398 540
rect -378 470 -374 540
rect -354 470 -350 540
rect -330 470 -326 540
rect -306 470 -302 540
rect -282 470 -278 540
rect -258 470 -254 540
rect -234 470 -230 540
rect -210 470 -206 540
rect -186 470 -182 540
rect -162 470 -158 540
rect -138 470 -134 540
rect -114 470 -110 540
rect -90 470 -86 540
rect -66 470 -62 540
rect -42 470 -38 540
rect -35 539 -21 540
rect -18 515 -11 563
rect -18 470 -14 515
rect 6 470 10 564
rect 30 470 34 564
rect 54 470 58 564
rect 78 470 82 564
rect 102 470 106 564
rect 126 470 130 564
rect 150 470 154 564
rect 174 470 178 564
rect 198 470 202 564
rect 222 470 226 564
rect 246 470 250 564
rect 259 518 293 519
rect 294 518 298 564
rect 318 518 322 564
rect 342 518 346 564
rect 366 518 370 564
rect 390 518 394 564
rect 414 518 418 564
rect 438 518 442 564
rect 462 518 466 564
rect 486 518 490 564
rect 510 518 514 564
rect 534 518 538 564
rect 558 518 562 564
rect 582 518 586 564
rect 606 518 610 564
rect 630 518 634 564
rect 654 518 658 564
rect 678 518 682 564
rect 702 518 706 564
rect 726 518 730 564
rect 750 518 754 564
rect 774 518 778 564
rect 798 518 802 564
rect 822 518 826 564
rect 846 518 850 564
rect 870 518 874 564
rect 894 518 898 564
rect 918 518 922 564
rect 942 518 946 564
rect 966 518 970 564
rect 990 518 994 564
rect 1014 518 1018 564
rect 1038 518 1042 564
rect 1062 518 1066 564
rect 1086 518 1090 564
rect 1110 518 1114 564
rect 1134 518 1138 564
rect 1147 557 1152 564
rect 1158 557 1162 564
rect 1157 543 1162 557
rect 1182 518 1186 612
rect 1206 518 1210 612
rect 1230 518 1234 612
rect 1254 519 1258 612
rect 1267 533 1272 543
rect 1278 533 1282 612
rect 1291 605 1296 612
rect 1302 605 1306 612
rect 1301 591 1306 605
rect 1277 519 1282 533
rect 1243 518 1277 519
rect 259 516 1277 518
rect 259 509 264 516
rect 294 515 298 516
rect 269 495 274 509
rect 283 505 291 509
rect 277 495 283 505
rect 270 470 274 495
rect 294 491 301 515
rect 318 470 322 516
rect 342 470 346 516
rect 366 470 370 516
rect 390 470 394 516
rect 414 470 418 516
rect 438 470 442 516
rect 462 470 466 516
rect 486 470 490 516
rect 510 470 514 516
rect 534 470 538 516
rect 558 470 562 516
rect 582 471 586 516
rect 571 470 605 471
rect -2393 468 605 470
rect -2371 422 -2366 468
rect -2348 422 -2343 468
rect -2325 464 -2320 468
rect -2317 464 -2309 468
rect -2325 452 -2317 464
rect -2066 463 -2062 468
rect -2147 460 -2134 462
rect -2292 454 -2071 460
rect -2325 432 -2320 452
rect -2092 438 -2062 440
rect -2094 434 -2062 438
rect -2325 422 -2317 432
rect -2095 424 -2084 428
rect -2000 425 -1992 468
rect -1846 461 -1806 468
rect -1663 464 -1655 468
rect -1846 454 -1680 460
rect -1671 452 -1663 464
rect -1854 438 -1806 440
rect -1854 434 -1680 438
rect -2119 422 -2069 424
rect -2054 422 -1892 425
rect -1671 422 -1663 432
rect -1642 422 -1637 468
rect -1619 422 -1614 468
rect -1530 422 -1526 468
rect -1506 422 -1502 468
rect -1482 422 -1478 468
rect -1458 422 -1454 468
rect -1434 422 -1430 468
rect -1410 422 -1406 468
rect -1386 443 -1379 467
rect -1386 422 -1382 443
rect -1362 422 -1358 468
rect -1338 422 -1334 468
rect -1314 422 -1310 468
rect -1290 422 -1286 468
rect -1266 422 -1262 468
rect -1242 422 -1238 468
rect -1218 422 -1214 468
rect -1194 422 -1190 468
rect -1170 422 -1166 468
rect -1146 422 -1142 468
rect -1122 422 -1118 468
rect -1098 422 -1094 468
rect -1074 422 -1070 468
rect -1050 422 -1046 468
rect -1026 422 -1022 468
rect -1002 422 -998 468
rect -978 422 -974 468
rect -954 422 -950 468
rect -930 422 -926 468
rect -2393 420 -909 422
rect -2371 398 -2366 420
rect -2348 398 -2343 420
rect -2325 416 -2317 420
rect -2325 400 -2320 416
rect -2309 404 -2301 416
rect -2095 414 -2084 420
rect -2054 419 -1906 420
rect -2054 418 -2036 419
rect -2084 412 -2079 414
rect -2317 400 -2309 404
rect -2092 403 -2079 410
rect -2000 406 -1992 419
rect -1920 418 -1906 419
rect -1671 416 -1663 420
rect -1846 412 -1806 414
rect -1854 406 -1806 410
rect -2054 403 -1982 406
rect -1966 403 -1806 406
rect -1655 404 -1647 416
rect -2003 400 -1992 403
rect -1904 401 -1902 403
rect -1854 401 -1846 403
rect -2325 398 -2317 400
rect -2033 398 -1992 400
rect -1854 399 -1806 401
rect -1663 400 -1655 404
rect -1864 398 -1796 399
rect -1671 398 -1663 400
rect -1642 398 -1637 420
rect -1619 398 -1614 420
rect -1530 398 -1526 420
rect -1506 398 -1502 420
rect -1482 398 -1478 420
rect -1458 398 -1454 420
rect -1434 398 -1430 420
rect -1410 398 -1406 420
rect -1386 398 -1382 420
rect -1362 398 -1358 420
rect -1338 398 -1334 420
rect -1314 398 -1310 420
rect -1290 398 -1286 420
rect -1266 398 -1262 420
rect -1242 398 -1238 420
rect -1218 398 -1214 420
rect -1194 398 -1190 420
rect -1170 398 -1166 420
rect -1146 398 -1142 420
rect -1122 398 -1118 420
rect -1098 398 -1094 420
rect -1074 398 -1070 420
rect -1050 398 -1046 420
rect -1026 398 -1022 420
rect -1002 398 -998 420
rect -978 398 -974 420
rect -954 398 -950 420
rect -930 398 -926 420
rect -923 419 -909 420
rect -906 419 -899 443
rect -906 398 -902 419
rect -882 398 -878 468
rect -858 398 -854 468
rect -834 398 -830 468
rect -810 398 -806 468
rect -786 398 -782 468
rect -773 446 -739 447
rect -738 446 -734 468
rect -714 446 -710 468
rect -690 446 -686 468
rect -666 446 -662 468
rect -642 446 -638 468
rect -618 446 -614 468
rect -594 446 -590 468
rect -570 446 -566 468
rect -546 446 -542 468
rect -522 446 -518 468
rect -498 446 -494 468
rect -474 446 -470 468
rect -450 446 -446 468
rect -426 446 -422 468
rect -402 446 -398 468
rect -378 446 -374 468
rect -354 446 -350 468
rect -330 446 -326 468
rect -306 446 -302 468
rect -282 446 -278 468
rect -258 446 -254 468
rect -234 446 -230 468
rect -210 446 -206 468
rect -186 446 -182 468
rect -162 446 -158 468
rect -138 446 -134 468
rect -114 446 -110 468
rect -90 446 -86 468
rect -66 446 -62 468
rect -42 446 -38 468
rect -18 446 -14 468
rect 6 446 10 468
rect 30 446 34 468
rect 54 446 58 468
rect 78 446 82 468
rect 102 446 106 468
rect 126 446 130 468
rect 150 446 154 468
rect 174 446 178 468
rect 198 446 202 468
rect 222 446 226 468
rect 246 446 250 468
rect 270 446 274 468
rect 318 446 322 468
rect 342 446 346 468
rect 366 446 370 468
rect 390 446 394 468
rect 414 446 418 468
rect 438 446 442 468
rect 462 446 466 468
rect 486 446 490 468
rect 510 446 514 468
rect 534 446 538 468
rect 558 446 562 468
rect 571 461 576 468
rect 582 461 586 468
rect 581 447 586 461
rect 606 446 610 516
rect 630 446 634 516
rect 654 446 658 516
rect 678 446 682 516
rect 702 446 706 516
rect 726 446 730 516
rect 750 446 754 516
rect 774 446 778 516
rect 798 446 802 516
rect 822 446 826 516
rect 846 446 850 516
rect 870 446 874 516
rect 894 446 898 516
rect 918 446 922 516
rect 942 446 946 516
rect 966 446 970 516
rect 990 446 994 516
rect 1014 446 1018 516
rect 1038 446 1042 516
rect 1062 446 1066 516
rect 1086 446 1090 516
rect 1110 446 1114 516
rect 1134 446 1138 516
rect 1147 485 1152 495
rect 1182 491 1186 516
rect 1157 471 1162 485
rect 1171 481 1179 485
rect 1165 471 1171 481
rect 1158 446 1162 471
rect 1182 467 1189 491
rect 1206 447 1210 516
rect 1219 485 1224 495
rect 1230 485 1234 516
rect 1243 509 1248 516
rect 1254 509 1258 516
rect 1253 495 1258 509
rect 1229 471 1234 485
rect 1195 446 1229 447
rect -773 444 1229 446
rect -773 437 -768 444
rect -763 423 -758 437
rect -762 398 -758 423
rect -738 419 -734 444
rect -2393 396 -741 398
rect -2371 374 -2366 396
rect -2348 374 -2343 396
rect -2325 388 -2317 396
rect -2079 393 -2018 396
rect -2003 395 -1966 396
rect -2000 394 -1982 395
rect -2000 393 -1992 394
rect -2084 389 -2009 393
rect -2028 388 -2009 389
rect -2000 389 -1854 393
rect -1846 389 -1798 396
rect -2325 374 -2320 388
rect -2309 376 -2301 388
rect -2028 386 -2018 388
rect -2092 376 -2084 383
rect -2023 379 -2014 386
rect -2000 379 -1992 389
rect -1671 388 -1663 396
rect -1846 385 -1806 387
rect -1854 379 -1806 383
rect -2054 376 -1806 379
rect -1655 376 -1647 388
rect -2317 374 -2309 376
rect -2054 374 -2024 376
rect -2000 374 -1992 376
rect -1663 374 -1655 376
rect -1642 374 -1637 396
rect -1619 374 -1614 396
rect -1530 374 -1526 396
rect -1506 374 -1502 396
rect -1482 374 -1478 396
rect -1458 374 -1454 396
rect -1434 374 -1430 396
rect -1410 374 -1406 396
rect -1386 374 -1382 396
rect -1362 374 -1358 396
rect -1338 374 -1334 396
rect -1314 374 -1310 396
rect -1290 374 -1286 396
rect -1266 374 -1262 396
rect -1242 374 -1238 396
rect -1218 374 -1214 396
rect -1194 374 -1190 396
rect -1170 374 -1166 396
rect -1146 374 -1142 396
rect -1122 374 -1118 396
rect -1098 374 -1094 396
rect -1074 374 -1070 396
rect -1050 374 -1046 396
rect -1026 374 -1022 396
rect -1002 374 -998 396
rect -978 374 -974 396
rect -954 374 -950 396
rect -930 374 -926 396
rect -906 374 -902 396
rect -882 374 -878 396
rect -858 374 -854 396
rect -834 374 -830 396
rect -810 374 -806 396
rect -786 374 -782 396
rect -762 374 -758 396
rect -755 395 -741 396
rect -738 395 -731 419
rect -714 374 -710 444
rect -690 374 -686 444
rect -666 374 -662 444
rect -642 374 -638 444
rect -618 374 -614 444
rect -594 374 -590 444
rect -570 374 -566 444
rect -546 374 -542 444
rect -522 374 -518 444
rect -498 374 -494 444
rect -474 374 -470 444
rect -450 374 -446 444
rect -426 374 -422 444
rect -402 374 -398 444
rect -378 374 -374 444
rect -354 374 -350 444
rect -330 374 -326 444
rect -306 374 -302 444
rect -282 374 -278 444
rect -258 374 -254 444
rect -234 374 -230 444
rect -210 374 -206 444
rect -186 374 -182 444
rect -162 374 -158 444
rect -138 374 -134 444
rect -114 374 -110 444
rect -90 374 -86 444
rect -66 374 -62 444
rect -42 374 -38 444
rect -18 374 -14 444
rect 6 375 10 444
rect -5 374 29 375
rect -2393 372 -2064 374
rect -2060 372 29 374
rect -2371 326 -2366 372
rect -2348 326 -2343 372
rect -2325 360 -2317 372
rect -2060 369 -2054 372
rect -2084 362 -2054 369
rect -2050 366 -2044 368
rect -2325 340 -2320 360
rect -2064 358 -2054 362
rect -2325 332 -2317 340
rect -2101 335 -2071 338
rect -2325 326 -2320 332
rect -2317 326 -2309 332
rect -2000 330 -1992 372
rect -1846 371 -1806 372
rect -1846 362 -1798 369
rect -1671 360 -1663 372
rect -1846 358 -1806 360
rect -1854 344 -1680 348
rect -1846 335 -1798 338
rect -2079 329 -2043 330
rect -2007 329 -1991 330
rect -2079 328 -2071 329
rect -2079 326 -2029 328
rect -2011 326 -1991 329
rect -1846 327 -1806 333
rect -1671 332 -1663 340
rect -1864 326 -1796 327
rect -1663 326 -1655 332
rect -1642 326 -1637 372
rect -1619 326 -1614 372
rect -1530 326 -1526 372
rect -1506 326 -1502 372
rect -1482 326 -1478 372
rect -1458 326 -1454 372
rect -1434 326 -1430 372
rect -1410 326 -1406 372
rect -1386 326 -1382 372
rect -1362 326 -1358 372
rect -1338 326 -1334 372
rect -1314 326 -1310 372
rect -1290 326 -1286 372
rect -1266 326 -1262 372
rect -1242 326 -1238 372
rect -1218 326 -1214 372
rect -1194 326 -1190 372
rect -1170 326 -1166 372
rect -1146 326 -1142 372
rect -1122 326 -1118 372
rect -1098 326 -1094 372
rect -1074 326 -1070 372
rect -1050 326 -1046 372
rect -1026 326 -1022 372
rect -1002 326 -998 372
rect -978 326 -974 372
rect -954 326 -950 372
rect -930 326 -926 372
rect -906 326 -902 372
rect -882 326 -878 372
rect -858 326 -854 372
rect -834 326 -830 372
rect -810 326 -806 372
rect -786 326 -782 372
rect -762 326 -758 372
rect -738 350 -731 371
rect -714 350 -710 372
rect -690 350 -686 372
rect -666 350 -662 372
rect -642 350 -638 372
rect -618 350 -614 372
rect -594 350 -590 372
rect -570 350 -566 372
rect -546 350 -542 372
rect -522 350 -518 372
rect -498 350 -494 372
rect -474 350 -470 372
rect -450 350 -446 372
rect -426 350 -422 372
rect -402 350 -398 372
rect -378 350 -374 372
rect -354 350 -350 372
rect -330 350 -326 372
rect -306 350 -302 372
rect -282 350 -278 372
rect -258 350 -254 372
rect -234 350 -230 372
rect -210 350 -206 372
rect -186 350 -182 372
rect -162 350 -158 372
rect -138 350 -134 372
rect -114 350 -110 372
rect -90 350 -86 372
rect -66 350 -62 372
rect -42 350 -38 372
rect -18 350 -14 372
rect -5 365 0 372
rect 6 365 10 372
rect 5 351 10 365
rect 6 350 10 351
rect 30 350 34 444
rect 54 350 58 444
rect 78 350 82 444
rect 102 350 106 444
rect 126 350 130 444
rect 150 350 154 444
rect 174 350 178 444
rect 198 350 202 444
rect 222 350 226 444
rect 246 350 250 444
rect 270 350 274 444
rect 294 422 301 443
rect 318 422 322 444
rect 342 422 346 444
rect 366 422 370 444
rect 390 422 394 444
rect 414 422 418 444
rect 438 422 442 444
rect 462 422 466 444
rect 486 422 490 444
rect 510 422 514 444
rect 534 422 538 444
rect 558 422 562 444
rect 571 422 605 423
rect 277 420 605 422
rect 277 419 291 420
rect 294 419 301 420
rect 294 350 298 419
rect 318 350 322 420
rect 342 351 346 420
rect 331 350 365 351
rect -755 348 365 350
rect -755 347 -741 348
rect -738 347 -731 348
rect -738 326 -734 347
rect -714 326 -710 348
rect -690 326 -686 348
rect -666 326 -662 348
rect -642 326 -638 348
rect -618 326 -614 348
rect -594 326 -590 348
rect -570 326 -566 348
rect -546 326 -542 348
rect -522 326 -518 348
rect -498 326 -494 348
rect -474 326 -470 348
rect -450 326 -446 348
rect -426 326 -422 348
rect -402 326 -398 348
rect -378 326 -374 348
rect -354 326 -350 348
rect -330 326 -326 348
rect -306 326 -302 348
rect -282 326 -278 348
rect -258 326 -254 348
rect -234 326 -230 348
rect -210 326 -206 348
rect -186 326 -182 348
rect -162 326 -158 348
rect -138 326 -134 348
rect -114 326 -110 348
rect -90 326 -86 348
rect -66 326 -62 348
rect -42 326 -38 348
rect -18 326 -14 348
rect 6 326 10 348
rect 30 326 34 348
rect 54 326 58 348
rect 78 326 82 348
rect 102 326 106 348
rect 126 326 130 348
rect 150 326 154 348
rect 174 326 178 348
rect 198 326 202 348
rect 222 326 226 348
rect 246 326 250 348
rect 270 326 274 348
rect 294 326 298 348
rect 318 326 322 348
rect 331 341 336 348
rect 342 341 346 348
rect 341 327 346 341
rect 366 326 370 420
rect 390 326 394 420
rect 414 326 418 420
rect 438 326 442 420
rect 462 326 466 420
rect 486 326 490 420
rect 510 326 514 420
rect 534 326 538 420
rect 558 326 562 420
rect 571 413 576 420
rect 581 399 586 413
rect 582 326 586 399
rect 606 395 610 444
rect 606 371 613 395
rect -2393 324 603 326
rect -2371 278 -2366 324
rect -2348 278 -2343 324
rect -2325 312 -2320 324
rect -2079 322 -2071 324
rect -2072 320 -2071 322
rect -2109 315 -2101 320
rect -2101 313 -2079 315
rect -2069 313 -2068 320
rect -2325 304 -2317 312
rect -2079 308 -2071 313
rect -2325 284 -2320 304
rect -2317 296 -2309 304
rect -2074 299 -2071 308
rect -2069 304 -2068 308
rect -2109 290 -2079 293
rect -2325 278 -2317 284
rect -2080 278 -2071 279
rect -2000 278 -1992 324
rect -1846 322 -1806 324
rect -1854 317 -1806 321
rect -1854 315 -1846 317
rect -1846 313 -1806 315
rect -1806 311 -1798 313
rect -1846 308 -1798 311
rect -1846 295 -1806 306
rect -1671 304 -1663 312
rect -1663 296 -1655 304
rect -1854 290 -1680 294
rect -1926 278 -1892 281
rect -1671 278 -1663 284
rect -1642 278 -1637 324
rect -1619 278 -1614 324
rect -1530 278 -1526 324
rect -1506 278 -1502 324
rect -1482 278 -1478 324
rect -1458 278 -1454 324
rect -1434 278 -1430 324
rect -1410 278 -1406 324
rect -1386 278 -1382 324
rect -1362 278 -1358 324
rect -1338 278 -1334 324
rect -1314 278 -1310 324
rect -1290 278 -1286 324
rect -1266 278 -1262 324
rect -1242 278 -1238 324
rect -1218 278 -1214 324
rect -1194 278 -1190 324
rect -1170 278 -1166 324
rect -1146 278 -1142 324
rect -1122 278 -1118 324
rect -1098 278 -1094 324
rect -1074 278 -1070 324
rect -1050 278 -1046 324
rect -1026 278 -1022 324
rect -1002 278 -998 324
rect -978 278 -974 324
rect -954 278 -950 324
rect -930 278 -926 324
rect -906 278 -902 324
rect -882 278 -878 324
rect -858 278 -854 324
rect -834 278 -830 324
rect -810 278 -806 324
rect -786 278 -782 324
rect -762 278 -758 324
rect -738 278 -734 324
rect -714 278 -710 324
rect -690 278 -686 324
rect -666 278 -662 324
rect -642 278 -638 324
rect -618 278 -614 324
rect -594 278 -590 324
rect -570 278 -566 324
rect -546 279 -542 324
rect -557 278 -523 279
rect -2393 276 -523 278
rect -2371 254 -2366 276
rect -2348 254 -2343 276
rect -2325 270 -2317 276
rect -2325 254 -2320 270
rect -2317 268 -2309 270
rect -2309 256 -2301 268
rect -2080 267 -2071 276
rect -2068 266 -2059 267
rect -2068 259 -2038 266
rect -2317 254 -2309 256
rect -2068 254 -2059 259
rect -2000 258 -1992 276
rect -1846 268 -1794 276
rect -1671 270 -1663 276
rect -1663 268 -1655 270
rect -1852 259 -1804 266
rect -2011 256 -1983 258
rect -2025 255 -1983 256
rect -2025 254 -1975 255
rect -1846 254 -1804 257
rect -1655 256 -1647 268
rect -1663 254 -1655 256
rect -1642 254 -1637 276
rect -1619 254 -1614 276
rect -1530 254 -1526 276
rect -1506 254 -1502 276
rect -1482 254 -1478 276
rect -1458 254 -1454 276
rect -1434 254 -1430 276
rect -1410 254 -1406 276
rect -1386 254 -1382 276
rect -1362 254 -1358 276
rect -1338 254 -1334 276
rect -1314 254 -1310 276
rect -1290 254 -1286 276
rect -1266 254 -1262 276
rect -1242 254 -1238 276
rect -1218 254 -1214 276
rect -1194 254 -1190 276
rect -1170 254 -1166 276
rect -1146 254 -1142 276
rect -1122 254 -1118 276
rect -1098 254 -1094 276
rect -1074 254 -1070 276
rect -1050 254 -1046 276
rect -1026 254 -1022 276
rect -1002 254 -998 276
rect -978 254 -974 276
rect -954 254 -950 276
rect -930 254 -926 276
rect -906 254 -902 276
rect -882 254 -878 276
rect -858 254 -854 276
rect -834 254 -830 276
rect -810 254 -806 276
rect -786 255 -782 276
rect -797 254 -763 255
rect -2393 252 -763 254
rect -2371 230 -2366 252
rect -2348 230 -2343 252
rect -2325 242 -2317 252
rect -2068 251 -2038 252
rect -2068 249 -2059 251
rect -2013 250 -1983 252
rect -1846 251 -1804 252
rect -2000 249 -1983 250
rect -1862 249 -1798 250
rect -2076 242 -2068 249
rect -2061 242 -2045 244
rect -2038 242 -2001 249
rect -2325 230 -2320 242
rect -2317 240 -2309 242
rect -2309 230 -2301 240
rect -2068 239 -2045 242
rect -2015 241 -2001 242
rect -2068 232 -2038 239
rect -2068 230 -2045 232
rect -2000 230 -1992 249
rect -1985 247 -1796 249
rect -1985 242 -1852 247
rect -1846 242 -1796 247
rect -1671 242 -1663 252
rect -1846 241 -1798 242
rect -1663 240 -1655 242
rect -1852 232 -1804 239
rect -1976 230 -1940 231
rect -1655 230 -1647 240
rect -1642 230 -1637 252
rect -1619 230 -1614 252
rect -1530 230 -1526 252
rect -1506 230 -1502 252
rect -1482 230 -1478 252
rect -1458 230 -1454 252
rect -1434 230 -1430 252
rect -1410 230 -1406 252
rect -1386 230 -1382 252
rect -1362 230 -1358 252
rect -1338 230 -1334 252
rect -1314 230 -1310 252
rect -1290 230 -1286 252
rect -1266 230 -1262 252
rect -1242 230 -1238 252
rect -1218 230 -1214 252
rect -1194 230 -1190 252
rect -1170 230 -1166 252
rect -1146 230 -1142 252
rect -1122 230 -1118 252
rect -1098 230 -1094 252
rect -1074 230 -1070 252
rect -1050 230 -1046 252
rect -1026 230 -1022 252
rect -1002 230 -998 252
rect -978 230 -974 252
rect -954 230 -950 252
rect -930 230 -926 252
rect -906 230 -902 252
rect -882 230 -878 252
rect -858 230 -854 252
rect -834 230 -830 252
rect -810 230 -806 252
rect -797 245 -792 252
rect -786 245 -782 252
rect -787 231 -782 245
rect -786 230 -782 231
rect -762 230 -758 276
rect -738 230 -734 276
rect -714 230 -710 276
rect -690 230 -686 276
rect -666 230 -662 276
rect -642 230 -638 276
rect -618 230 -614 276
rect -594 230 -590 276
rect -570 230 -566 276
rect -557 269 -552 276
rect -546 269 -542 276
rect -547 255 -542 269
rect -546 230 -542 255
rect -522 230 -518 324
rect -498 230 -494 324
rect -474 230 -470 324
rect -450 230 -446 324
rect -426 230 -422 324
rect -402 230 -398 324
rect -378 230 -374 324
rect -354 230 -350 324
rect -330 230 -326 324
rect -306 230 -302 324
rect -282 230 -278 324
rect -258 230 -254 324
rect -234 230 -230 324
rect -210 230 -206 324
rect -186 231 -182 324
rect -197 230 -163 231
rect -2393 228 -163 230
rect -2371 158 -2366 228
rect -2348 158 -2343 228
rect -2325 226 -2320 228
rect -2317 226 -2309 228
rect -2325 214 -2317 226
rect -2068 222 -2059 228
rect -2076 215 -2071 222
rect -2068 214 -2059 215
rect -2325 194 -2320 214
rect -2317 212 -2309 214
rect -2325 186 -2317 194
rect -2060 188 -2030 191
rect -2325 166 -2320 186
rect -2317 178 -2309 186
rect -2060 175 -2038 186
rect -2033 179 -2030 188
rect -2028 184 -2027 188
rect -2068 170 -2038 173
rect -2325 158 -2317 166
rect -2000 161 -1992 228
rect -1846 224 -1804 228
rect -1663 226 -1655 228
rect -1846 214 -1794 223
rect -1671 214 -1663 226
rect -1663 212 -1655 214
rect -1912 203 -1884 205
rect -1852 197 -1804 201
rect -1844 188 -1796 191
rect -1671 186 -1663 194
rect -1844 175 -1804 186
rect -1663 178 -1655 186
rect -1852 170 -1680 174
rect -2119 158 -2069 160
rect -2007 158 -1977 161
rect -1926 158 -1892 161
rect -1671 158 -1663 166
rect -1642 158 -1637 228
rect -1619 158 -1614 228
rect -1530 158 -1526 228
rect -1506 158 -1502 228
rect -1482 158 -1478 228
rect -1458 158 -1454 228
rect -1434 158 -1430 228
rect -1410 158 -1406 228
rect -1386 158 -1382 228
rect -1362 158 -1358 228
rect -1338 158 -1334 228
rect -1314 158 -1310 228
rect -1290 158 -1286 228
rect -1266 158 -1262 228
rect -1242 158 -1238 228
rect -1218 158 -1214 228
rect -1194 158 -1190 228
rect -1170 158 -1166 228
rect -1146 158 -1142 228
rect -1122 158 -1118 228
rect -1098 158 -1094 228
rect -1074 158 -1070 228
rect -1050 158 -1046 228
rect -1026 158 -1022 228
rect -1002 158 -998 228
rect -978 158 -974 228
rect -954 158 -950 228
rect -930 158 -926 228
rect -906 158 -902 228
rect -882 158 -878 228
rect -858 158 -854 228
rect -834 158 -830 228
rect -810 158 -806 228
rect -786 158 -782 228
rect -762 179 -758 228
rect -2393 156 -765 158
rect -2371 134 -2366 156
rect -2348 134 -2343 156
rect -2325 152 -2317 156
rect -2325 136 -2320 152
rect -2317 150 -2309 152
rect -2309 138 -2301 150
rect -2000 142 -1992 156
rect -1671 152 -1663 156
rect -1663 150 -1655 152
rect -1844 148 -1806 150
rect -1854 142 -1806 146
rect -2068 139 -2060 142
rect -2030 139 -1958 142
rect -1942 139 -1806 142
rect -2317 136 -2309 138
rect -2000 136 -1992 139
rect -1655 138 -1647 150
rect -2325 134 -2317 136
rect -2033 134 -1992 136
rect -1844 135 -1806 137
rect -1663 136 -1655 138
rect -1864 134 -1796 135
rect -1671 134 -1663 136
rect -1642 134 -1637 156
rect -1619 134 -1614 156
rect -1530 134 -1526 156
rect -1506 134 -1502 156
rect -1482 134 -1478 156
rect -1458 134 -1454 156
rect -1434 134 -1430 156
rect -1410 134 -1406 156
rect -1386 134 -1382 156
rect -1362 134 -1358 156
rect -1338 134 -1334 156
rect -1314 134 -1310 156
rect -1290 134 -1286 156
rect -1266 134 -1262 156
rect -1242 134 -1238 156
rect -1218 134 -1214 156
rect -1194 134 -1190 156
rect -1170 134 -1166 156
rect -1146 134 -1142 156
rect -1122 134 -1118 156
rect -1098 134 -1094 156
rect -1074 134 -1070 156
rect -1050 134 -1046 156
rect -1026 134 -1022 156
rect -1002 134 -998 156
rect -978 134 -974 156
rect -954 134 -950 156
rect -930 134 -926 156
rect -906 134 -902 156
rect -882 134 -878 156
rect -858 134 -854 156
rect -834 134 -830 156
rect -810 134 -806 156
rect -786 134 -782 156
rect -779 155 -765 156
rect -762 155 -755 179
rect -762 134 -758 155
rect -738 134 -734 228
rect -714 134 -710 228
rect -690 134 -686 228
rect -666 134 -662 228
rect -653 197 -648 207
rect -642 197 -638 228
rect -643 183 -638 197
rect -653 182 -619 183
rect -618 182 -614 228
rect -594 182 -590 228
rect -570 182 -566 228
rect -546 182 -542 228
rect -522 203 -518 228
rect -653 180 -525 182
rect -653 173 -648 180
rect -643 159 -638 173
rect -642 134 -638 159
rect -618 134 -614 180
rect -594 134 -590 180
rect -570 134 -566 180
rect -546 134 -542 180
rect -539 179 -525 180
rect -522 179 -515 203
rect -522 134 -518 179
rect -498 134 -494 228
rect -474 134 -470 228
rect -450 134 -446 228
rect -426 134 -422 228
rect -402 134 -398 228
rect -378 134 -374 228
rect -354 134 -350 228
rect -330 134 -326 228
rect -306 134 -302 228
rect -282 134 -278 228
rect -258 134 -254 228
rect -234 134 -230 228
rect -210 134 -206 228
rect -197 221 -192 228
rect -186 221 -182 228
rect -187 207 -182 221
rect -197 197 -192 207
rect -187 183 -182 197
rect -186 134 -182 183
rect -162 155 -158 324
rect -2393 132 -165 134
rect -2371 110 -2366 132
rect -2348 110 -2343 132
rect -2325 124 -2317 132
rect -2060 129 -2030 132
rect -2000 129 -1992 132
rect -1972 130 -1958 132
rect -1904 129 -1798 132
rect -2078 125 -2020 129
rect -2023 124 -2020 125
rect -2000 127 -1798 129
rect -2000 125 -1854 127
rect -1844 125 -1798 127
rect -2325 110 -2320 124
rect -2317 122 -2309 124
rect -2020 122 -2004 124
rect -2000 122 -1992 125
rect -1671 124 -1663 132
rect -2309 110 -2301 122
rect -2020 120 -1992 122
rect -1844 121 -1806 123
rect -1663 122 -1655 124
rect -2023 115 -1992 120
rect -1854 115 -1806 119
rect -2068 112 -2060 115
rect -2030 112 -1806 115
rect -2074 110 -2060 112
rect -2020 110 -2004 112
rect -2000 110 -1992 112
rect -1655 110 -1647 122
rect -1642 110 -1637 132
rect -1619 110 -1614 132
rect -1530 110 -1526 132
rect -1506 110 -1502 132
rect -1482 110 -1478 132
rect -1458 110 -1454 132
rect -1434 110 -1430 132
rect -1410 110 -1406 132
rect -1386 110 -1382 132
rect -1362 110 -1358 132
rect -1338 110 -1334 132
rect -1314 110 -1310 132
rect -1290 110 -1286 132
rect -1266 110 -1262 132
rect -1242 110 -1238 132
rect -1218 110 -1214 132
rect -1194 110 -1190 132
rect -1170 110 -1166 132
rect -1146 110 -1142 132
rect -1122 110 -1118 132
rect -1098 110 -1094 132
rect -1074 110 -1070 132
rect -1050 110 -1046 132
rect -1026 110 -1022 132
rect -1002 110 -998 132
rect -978 110 -974 132
rect -954 110 -950 132
rect -930 110 -926 132
rect -906 110 -902 132
rect -882 110 -878 132
rect -858 110 -854 132
rect -834 110 -830 132
rect -810 110 -806 132
rect -786 110 -782 132
rect -762 110 -758 132
rect -738 110 -734 132
rect -714 110 -710 132
rect -690 110 -686 132
rect -666 110 -662 132
rect -642 110 -638 132
rect -618 131 -614 132
rect -2393 108 -2060 110
rect -2050 108 -621 110
rect -2371 62 -2366 108
rect -2348 62 -2343 108
rect -2325 96 -2317 108
rect -2109 105 -2108 108
rect -2117 98 -2108 105
rect -2325 76 -2320 96
rect -2317 94 -2309 96
rect -2109 94 -2108 98
rect -2060 98 -2030 105
rect -2060 94 -2034 98
rect -2325 68 -2317 76
rect -2101 71 -2071 74
rect -2325 62 -2320 68
rect -2317 62 -2309 68
rect -2000 66 -1992 108
rect -1844 107 -1806 108
rect -1844 98 -1798 105
rect -1671 96 -1663 108
rect -1844 94 -1806 96
rect -1663 94 -1655 96
rect -1854 80 -1680 84
rect -1846 71 -1798 74
rect -2079 65 -2043 66
rect -2007 65 -1991 66
rect -2079 64 -2071 65
rect -2079 62 -2029 64
rect -2011 62 -1991 65
rect -1846 63 -1806 69
rect -1671 68 -1663 76
rect -1864 62 -1796 63
rect -1663 62 -1655 68
rect -1642 62 -1637 108
rect -1619 62 -1614 108
rect -1530 62 -1526 108
rect -1506 62 -1502 108
rect -1482 62 -1478 108
rect -1458 62 -1454 108
rect -1434 62 -1430 108
rect -1410 62 -1406 108
rect -1386 62 -1382 108
rect -1362 62 -1358 108
rect -1338 62 -1334 108
rect -1314 62 -1310 108
rect -1290 62 -1286 108
rect -1266 62 -1262 108
rect -1242 62 -1238 108
rect -1218 62 -1214 108
rect -1194 62 -1190 108
rect -1170 62 -1166 108
rect -1146 62 -1142 108
rect -1122 62 -1118 108
rect -1098 62 -1094 108
rect -1074 62 -1070 108
rect -1050 62 -1046 108
rect -1026 62 -1022 108
rect -1002 62 -998 108
rect -978 62 -974 108
rect -954 62 -950 108
rect -930 62 -926 108
rect -906 62 -902 108
rect -882 62 -878 108
rect -858 62 -854 108
rect -834 62 -830 108
rect -810 62 -806 108
rect -786 62 -782 108
rect -762 62 -758 108
rect -738 62 -734 108
rect -714 62 -710 108
rect -690 62 -686 108
rect -666 62 -662 108
rect -642 62 -638 108
rect -635 107 -621 108
rect -618 86 -611 131
rect -594 86 -590 132
rect -570 86 -566 132
rect -546 86 -542 132
rect -522 86 -518 132
rect -498 86 -494 132
rect -474 86 -470 132
rect -450 86 -446 132
rect -426 86 -422 132
rect -402 86 -398 132
rect -378 86 -374 132
rect -354 86 -350 132
rect -330 86 -326 132
rect -306 86 -302 132
rect -282 86 -278 132
rect -258 86 -254 132
rect -234 86 -230 132
rect -210 86 -206 132
rect -186 86 -182 132
rect -179 131 -165 132
rect -162 110 -155 155
rect -138 110 -134 324
rect -114 110 -110 324
rect -90 110 -86 324
rect -66 110 -62 324
rect -42 110 -38 324
rect -18 110 -14 324
rect 6 110 10 324
rect 30 299 34 324
rect 30 275 37 299
rect 30 110 34 275
rect 54 110 58 324
rect 78 110 82 324
rect 102 110 106 324
rect 126 110 130 324
rect 150 110 154 324
rect 174 110 178 324
rect 198 110 202 324
rect 222 110 226 324
rect 246 110 250 324
rect 270 110 274 324
rect 294 110 298 324
rect 318 110 322 324
rect 331 302 365 303
rect 366 302 370 324
rect 390 302 394 324
rect 414 302 418 324
rect 438 302 442 324
rect 462 302 466 324
rect 486 302 490 324
rect 510 302 514 324
rect 534 302 538 324
rect 558 302 562 324
rect 582 302 586 324
rect 589 323 603 324
rect 606 323 613 347
rect 606 302 610 323
rect 630 302 634 444
rect 643 317 648 327
rect 654 317 658 444
rect 653 303 658 317
rect 678 302 682 444
rect 702 302 706 444
rect 726 302 730 444
rect 750 302 754 444
rect 774 302 778 444
rect 798 302 802 444
rect 822 302 826 444
rect 846 302 850 444
rect 870 302 874 444
rect 894 302 898 444
rect 918 302 922 444
rect 942 302 946 444
rect 966 302 970 444
rect 990 302 994 444
rect 1014 302 1018 444
rect 1038 302 1042 444
rect 1062 302 1066 444
rect 1086 302 1090 444
rect 1110 302 1114 444
rect 1134 302 1138 444
rect 1158 303 1162 444
rect 1195 437 1200 444
rect 1206 437 1210 444
rect 1205 423 1210 437
rect 1182 399 1189 419
rect 1171 398 1205 399
rect 1165 396 1205 398
rect 1165 395 1179 396
rect 1182 395 1189 396
rect 1171 389 1176 395
rect 1182 389 1186 395
rect 1181 375 1186 389
rect 1147 302 1181 303
rect 331 300 1181 302
rect 331 293 336 300
rect 341 279 346 293
rect 342 110 346 279
rect 366 275 370 300
rect 366 251 373 275
rect 366 206 373 227
rect 390 206 394 300
rect 414 206 418 300
rect 438 206 442 300
rect 462 206 466 300
rect 486 206 490 300
rect 510 206 514 300
rect 534 206 538 300
rect 558 206 562 300
rect 582 206 586 300
rect 606 206 610 300
rect 630 206 634 300
rect 643 269 648 279
rect 653 255 658 269
rect 654 206 658 255
rect 678 251 682 300
rect 678 227 685 251
rect 702 206 706 300
rect 726 206 730 300
rect 750 206 754 300
rect 774 206 778 300
rect 798 206 802 300
rect 822 206 826 300
rect 846 206 850 300
rect 870 206 874 300
rect 894 206 898 300
rect 918 206 922 300
rect 942 206 946 300
rect 966 206 970 300
rect 990 206 994 300
rect 1014 206 1018 300
rect 1038 206 1042 300
rect 1062 206 1066 300
rect 1086 206 1090 300
rect 1110 207 1114 300
rect 1123 269 1128 279
rect 1134 269 1138 300
rect 1147 293 1152 300
rect 1158 293 1162 300
rect 1157 279 1162 293
rect 1133 255 1138 269
rect 1099 206 1133 207
rect 349 204 1133 206
rect 349 203 363 204
rect 366 203 373 204
rect 366 110 370 203
rect 390 110 394 204
rect 414 110 418 204
rect 438 110 442 204
rect 462 110 466 204
rect 486 111 490 204
rect 475 110 509 111
rect -179 108 509 110
rect -179 107 -165 108
rect -162 107 -155 108
rect -162 87 -158 107
rect -173 86 -139 87
rect -635 84 -139 86
rect -635 83 -621 84
rect -618 83 -611 84
rect -618 62 -614 83
rect -594 62 -590 84
rect -570 62 -566 84
rect -546 62 -542 84
rect -522 62 -518 84
rect -498 62 -494 84
rect -474 62 -470 84
rect -450 62 -446 84
rect -426 62 -422 84
rect -402 62 -398 84
rect -378 62 -374 84
rect -354 62 -350 84
rect -330 62 -326 84
rect -306 62 -302 84
rect -282 62 -278 84
rect -258 62 -254 84
rect -234 62 -230 84
rect -210 62 -206 84
rect -186 62 -182 84
rect -173 77 -168 84
rect -162 77 -158 84
rect -163 63 -158 77
rect -138 62 -134 108
rect -114 62 -110 108
rect -90 62 -86 108
rect -66 62 -62 108
rect -42 62 -38 108
rect -18 62 -14 108
rect 6 62 10 108
rect 30 62 34 108
rect 54 62 58 108
rect 78 62 82 108
rect 102 62 106 108
rect 126 62 130 108
rect 150 62 154 108
rect 174 62 178 108
rect 198 62 202 108
rect 222 62 226 108
rect 246 62 250 108
rect 270 62 274 108
rect 294 63 298 108
rect 283 62 317 63
rect -2393 60 317 62
rect -2371 14 -2366 60
rect -2348 14 -2343 60
rect -2325 48 -2320 60
rect -2079 58 -2071 60
rect -2072 56 -2071 58
rect -2109 51 -2101 56
rect -2101 49 -2079 51
rect -2069 49 -2068 56
rect -2325 40 -2317 48
rect -2079 44 -2071 49
rect -2325 20 -2320 40
rect -2317 32 -2309 40
rect -2074 35 -2071 44
rect -2069 40 -2068 44
rect -2109 26 -2079 29
rect -2325 14 -2317 20
rect -2119 14 -2069 16
rect -2056 14 -2026 17
rect -2000 14 -1992 60
rect -1846 58 -1806 60
rect -1854 53 -1806 57
rect -1854 51 -1846 53
rect -1846 49 -1806 51
rect -1806 47 -1798 49
rect -1846 44 -1798 47
rect -1846 31 -1806 42
rect -1671 40 -1663 48
rect -1663 32 -1655 40
rect -1854 26 -1680 30
rect -1926 14 -1892 17
rect -1671 14 -1663 20
rect -1642 14 -1637 60
rect -1619 14 -1614 60
rect -1530 14 -1526 60
rect -1506 14 -1502 60
rect -1482 14 -1478 60
rect -1458 14 -1454 60
rect -1434 14 -1430 60
rect -1410 14 -1406 60
rect -1386 14 -1382 60
rect -1362 14 -1358 60
rect -1338 14 -1334 60
rect -1314 14 -1310 60
rect -1290 14 -1286 60
rect -1266 14 -1262 60
rect -1242 14 -1238 60
rect -1218 14 -1214 60
rect -1194 14 -1190 60
rect -1170 14 -1166 60
rect -1146 14 -1142 60
rect -1122 14 -1118 60
rect -1098 14 -1094 60
rect -1074 14 -1070 60
rect -1050 14 -1046 60
rect -1026 14 -1022 60
rect -1002 14 -998 60
rect -978 14 -974 60
rect -954 14 -950 60
rect -930 14 -926 60
rect -906 14 -902 60
rect -882 14 -878 60
rect -858 14 -854 60
rect -834 14 -830 60
rect -810 14 -806 60
rect -786 14 -782 60
rect -762 14 -758 60
rect -738 14 -734 60
rect -714 14 -710 60
rect -690 14 -686 60
rect -666 14 -662 60
rect -642 14 -638 60
rect -618 14 -614 60
rect -594 14 -590 60
rect -570 14 -566 60
rect -546 14 -542 60
rect -522 14 -518 60
rect -498 14 -494 60
rect -474 14 -470 60
rect -450 14 -446 60
rect -426 14 -422 60
rect -402 14 -398 60
rect -378 14 -374 60
rect -354 14 -350 60
rect -330 14 -326 60
rect -306 14 -302 60
rect -282 14 -278 60
rect -258 14 -254 60
rect -234 14 -230 60
rect -210 14 -206 60
rect -186 14 -182 60
rect -173 38 -139 39
rect -138 38 -134 60
rect -114 38 -110 60
rect -90 38 -86 60
rect -66 38 -62 60
rect -42 38 -38 60
rect -18 38 -14 60
rect 6 38 10 60
rect 30 38 34 60
rect 54 38 58 60
rect 78 38 82 60
rect 102 38 106 60
rect 126 38 130 60
rect 150 38 154 60
rect 174 38 178 60
rect 198 38 202 60
rect 222 38 226 60
rect 246 38 250 60
rect 270 38 274 60
rect 283 53 288 60
rect 294 53 298 60
rect 293 39 298 53
rect 318 38 322 108
rect 342 38 346 108
rect 366 38 370 108
rect 390 38 394 108
rect 414 38 418 108
rect 438 38 442 108
rect 462 38 466 108
rect 475 101 480 108
rect 486 101 490 108
rect 485 87 490 101
rect 475 86 509 87
rect 510 86 514 204
rect 534 86 538 204
rect 558 86 562 204
rect 582 86 586 204
rect 606 86 610 204
rect 630 86 634 204
rect 654 86 658 204
rect 678 182 685 203
rect 702 182 706 204
rect 726 182 730 204
rect 750 182 754 204
rect 774 182 778 204
rect 798 182 802 204
rect 822 182 826 204
rect 846 182 850 204
rect 870 182 874 204
rect 894 182 898 204
rect 918 182 922 204
rect 942 182 946 204
rect 966 182 970 204
rect 990 182 994 204
rect 1014 182 1018 204
rect 1038 182 1042 204
rect 1062 182 1066 204
rect 1086 183 1090 204
rect 1099 197 1104 204
rect 1110 197 1114 204
rect 1109 183 1114 197
rect 1075 182 1109 183
rect 661 180 1109 182
rect 661 179 675 180
rect 678 179 685 180
rect 678 86 682 179
rect 702 86 706 180
rect 726 86 730 180
rect 750 86 754 180
rect 774 86 778 180
rect 787 125 792 135
rect 798 125 802 180
rect 797 111 802 125
rect 787 110 821 111
rect 822 110 826 180
rect 846 110 850 180
rect 870 110 874 180
rect 894 110 898 180
rect 918 110 922 180
rect 942 110 946 180
rect 966 110 970 180
rect 990 110 994 180
rect 1014 110 1018 180
rect 1038 110 1042 180
rect 1062 110 1066 180
rect 1075 173 1080 180
rect 1086 173 1090 180
rect 1085 159 1090 173
rect 1075 149 1080 159
rect 1085 135 1090 149
rect 1086 111 1090 135
rect 1075 110 1109 111
rect 787 108 1109 110
rect 787 101 792 108
rect 797 87 802 101
rect 798 86 802 87
rect 822 86 826 108
rect 846 86 850 108
rect 870 86 874 108
rect 894 86 898 108
rect 918 86 922 108
rect 942 86 946 108
rect 966 86 970 108
rect 990 86 994 108
rect 1014 86 1018 108
rect 1038 86 1042 108
rect 1062 87 1066 108
rect 1075 101 1080 108
rect 1086 101 1090 108
rect 1085 87 1090 101
rect 1099 97 1107 101
rect 1093 87 1099 97
rect 1051 86 1085 87
rect 475 84 1085 86
rect 475 77 480 84
rect 485 63 490 77
rect 486 38 490 63
rect 510 38 514 84
rect 534 38 538 84
rect 558 38 562 84
rect 582 38 586 84
rect 606 38 610 84
rect 630 38 634 84
rect 654 38 658 84
rect 678 38 682 84
rect 702 38 706 84
rect 726 38 730 84
rect 750 38 754 84
rect 774 38 778 84
rect 798 38 802 84
rect 822 59 826 84
rect -173 36 819 38
rect -173 29 -168 36
rect -163 15 -158 29
rect -162 14 -158 15
rect -138 14 -134 36
rect -114 14 -110 36
rect -90 14 -86 36
rect -66 14 -62 36
rect -42 14 -38 36
rect -18 14 -14 36
rect 6 14 10 36
rect 30 14 34 36
rect 54 14 58 36
rect 78 14 82 36
rect 102 14 106 36
rect 126 14 130 36
rect 150 14 154 36
rect 174 14 178 36
rect 198 14 202 36
rect 222 14 226 36
rect 246 14 250 36
rect 270 14 274 36
rect 283 14 317 15
rect -2393 12 317 14
rect -2371 -10 -2366 12
rect -2348 -10 -2343 12
rect -2325 8 -2317 12
rect -2325 -8 -2320 8
rect -2317 4 -2309 8
rect -2309 -8 -2301 4
rect -2109 -5 -2079 2
rect -2000 1 -1992 12
rect -1671 8 -1663 12
rect -1846 4 -1806 6
rect -1663 4 -1655 8
rect -2009 -2 -1992 1
rect -1854 -2 -1806 2
rect -2071 -5 -1992 -2
rect -1983 -5 -1806 -2
rect -2009 -8 -1992 -5
rect -2325 -10 -2317 -8
rect -2033 -10 -1992 -8
rect -1846 -9 -1806 -7
rect -1655 -8 -1647 4
rect -1864 -10 -1796 -9
rect -1671 -10 -1663 -8
rect -1642 -10 -1637 12
rect -1619 -10 -1614 12
rect -1530 -10 -1526 12
rect -1506 -10 -1502 12
rect -1482 -10 -1478 12
rect -1458 -10 -1454 12
rect -1434 -10 -1430 12
rect -1410 -10 -1406 12
rect -1386 -10 -1382 12
rect -1362 -10 -1358 12
rect -1338 -10 -1334 12
rect -1314 -9 -1310 12
rect -1325 -10 -1291 -9
rect -2393 -12 -1291 -10
rect -2371 -34 -2366 -12
rect -2348 -34 -2343 -12
rect -2325 -20 -2317 -12
rect -2079 -15 -2035 -12
rect -2013 -14 -1992 -12
rect -2000 -15 -1992 -14
rect -1904 -15 -1798 -12
rect -2101 -19 -2009 -15
rect -2023 -20 -2009 -19
rect -2000 -17 -1798 -15
rect -2000 -19 -1854 -17
rect -1846 -19 -1798 -17
rect -2325 -34 -2320 -20
rect -2317 -24 -2309 -20
rect -2309 -34 -2301 -24
rect -2109 -32 -2101 -25
rect -2023 -29 -2021 -20
rect -2000 -29 -1992 -19
rect -1671 -20 -1663 -12
rect -1846 -23 -1806 -21
rect -1663 -24 -1655 -20
rect -1854 -29 -1806 -25
rect -2071 -32 -1806 -29
rect -2074 -34 -2031 -32
rect -2000 -34 -1992 -32
rect -1655 -34 -1647 -24
rect -1642 -34 -1637 -12
rect -1619 -34 -1614 -12
rect -1530 -34 -1526 -12
rect -1506 -34 -1502 -12
rect -1482 -34 -1478 -12
rect -1458 -34 -1454 -12
rect -1434 -34 -1430 -12
rect -1410 -34 -1406 -12
rect -1386 -34 -1382 -12
rect -1362 -34 -1358 -12
rect -1338 -34 -1334 -12
rect -1325 -19 -1320 -12
rect -1314 -19 -1310 -12
rect -1315 -33 -1310 -19
rect -1290 -34 -1286 12
rect -1266 -34 -1262 12
rect -1242 -34 -1238 12
rect -1218 -34 -1214 12
rect -1194 -34 -1190 12
rect -1170 -34 -1166 12
rect -1146 -34 -1142 12
rect -1122 -34 -1118 12
rect -1098 -34 -1094 12
rect -1074 -34 -1070 12
rect -1050 -34 -1046 12
rect -1026 -34 -1022 12
rect -1002 -34 -998 12
rect -978 -34 -974 12
rect -954 -34 -950 12
rect -930 -34 -926 12
rect -906 -34 -902 12
rect -882 -34 -878 12
rect -858 -34 -854 12
rect -834 -34 -830 12
rect -810 -34 -806 12
rect -786 -34 -782 12
rect -762 -34 -758 12
rect -738 -34 -734 12
rect -714 -34 -710 12
rect -690 -34 -686 12
rect -666 -34 -662 12
rect -642 -34 -638 12
rect -618 -34 -614 12
rect -594 -34 -590 12
rect -570 -34 -566 12
rect -546 -34 -542 12
rect -522 -34 -518 12
rect -498 -34 -494 12
rect -474 -34 -470 12
rect -450 -34 -446 12
rect -426 -34 -422 12
rect -402 -34 -398 12
rect -378 -34 -374 12
rect -354 -34 -350 12
rect -330 -34 -326 12
rect -306 -34 -302 12
rect -282 -34 -278 12
rect -258 -34 -254 12
rect -234 -34 -230 12
rect -210 -34 -206 12
rect -186 -34 -182 12
rect -162 -34 -158 12
rect -138 11 -134 12
rect -138 -13 -131 11
rect -114 -34 -110 12
rect -90 -34 -86 12
rect -66 -34 -62 12
rect -42 -34 -38 12
rect -18 -34 -14 12
rect 6 -34 10 12
rect 30 -34 34 12
rect 54 -34 58 12
rect 78 -34 82 12
rect 102 -34 106 12
rect 126 -34 130 12
rect 150 -34 154 12
rect 174 -34 178 12
rect 198 -34 202 12
rect 222 -34 226 12
rect 246 -34 250 12
rect 270 -34 274 12
rect 283 5 288 12
rect 293 -9 298 5
rect 294 -34 298 -9
rect 318 -13 322 36
rect -2393 -36 315 -34
rect -2371 -82 -2366 -36
rect -2348 -82 -2343 -36
rect -2325 -48 -2317 -36
rect -2074 -39 -2071 -36
rect -2101 -46 -2071 -39
rect -2325 -68 -2320 -48
rect -2317 -52 -2309 -48
rect -2064 -50 -2061 -42
rect -2325 -76 -2317 -68
rect -2101 -73 -2071 -70
rect -2325 -82 -2320 -76
rect -2317 -82 -2309 -76
rect -2000 -78 -1992 -36
rect -1846 -37 -1806 -36
rect -1846 -46 -1798 -39
rect -1671 -48 -1663 -36
rect -1846 -50 -1806 -48
rect -1663 -52 -1655 -48
rect -1854 -64 -1680 -60
rect -1846 -73 -1798 -70
rect -2079 -79 -2043 -78
rect -2007 -79 -1991 -78
rect -2079 -80 -2071 -79
rect -2079 -82 -2029 -80
rect -2011 -82 -1991 -79
rect -1846 -81 -1806 -75
rect -1671 -76 -1663 -68
rect -1864 -82 -1796 -81
rect -1663 -82 -1655 -76
rect -1642 -82 -1637 -36
rect -1619 -82 -1614 -36
rect -1530 -82 -1526 -36
rect -1506 -82 -1502 -36
rect -1482 -82 -1478 -36
rect -1458 -82 -1454 -36
rect -1434 -82 -1430 -36
rect -1410 -82 -1406 -36
rect -1386 -82 -1382 -36
rect -1362 -82 -1358 -36
rect -1338 -82 -1334 -36
rect -1290 -82 -1286 -36
rect -1266 -82 -1262 -36
rect -1242 -82 -1238 -36
rect -1218 -82 -1214 -36
rect -1194 -82 -1190 -36
rect -1170 -82 -1166 -36
rect -1146 -82 -1142 -36
rect -1122 -82 -1118 -36
rect -1098 -82 -1094 -36
rect -1074 -82 -1070 -36
rect -1050 -82 -1046 -36
rect -1026 -82 -1022 -36
rect -1002 -82 -998 -36
rect -989 -67 -984 -57
rect -978 -67 -974 -36
rect -979 -81 -974 -67
rect -954 -82 -950 -36
rect -930 -82 -926 -36
rect -906 -82 -902 -36
rect -882 -82 -878 -36
rect -858 -82 -854 -36
rect -834 -82 -830 -36
rect -810 -82 -806 -36
rect -786 -82 -782 -36
rect -762 -82 -758 -36
rect -738 -82 -734 -36
rect -714 -82 -710 -36
rect -690 -82 -686 -36
rect -666 -82 -662 -36
rect -642 -82 -638 -36
rect -618 -82 -614 -36
rect -594 -82 -590 -36
rect -570 -82 -566 -36
rect -546 -82 -542 -36
rect -522 -82 -518 -36
rect -498 -82 -494 -36
rect -474 -82 -470 -36
rect -450 -82 -446 -36
rect -426 -82 -422 -36
rect -402 -82 -398 -36
rect -378 -82 -374 -36
rect -354 -82 -350 -36
rect -330 -82 -326 -36
rect -306 -82 -302 -36
rect -282 -82 -278 -36
rect -258 -82 -254 -36
rect -234 -82 -230 -36
rect -210 -82 -206 -36
rect -186 -82 -182 -36
rect -162 -82 -158 -36
rect -138 -61 -131 -37
rect -138 -82 -134 -61
rect -114 -82 -110 -36
rect -90 -82 -86 -36
rect -66 -82 -62 -36
rect -42 -82 -38 -36
rect -18 -82 -14 -36
rect 6 -82 10 -36
rect 30 -82 34 -36
rect 54 -82 58 -36
rect 78 -82 82 -36
rect 102 -82 106 -36
rect 126 -82 130 -36
rect 150 -82 154 -36
rect 174 -82 178 -36
rect 198 -82 202 -36
rect 222 -82 226 -36
rect 246 -82 250 -36
rect 270 -82 274 -36
rect 294 -82 298 -36
rect 301 -37 315 -36
rect 318 -37 325 -13
rect -2393 -84 315 -82
rect -2371 -154 -2366 -84
rect -2348 -154 -2343 -84
rect -2325 -96 -2320 -84
rect -2079 -86 -2071 -84
rect -2072 -88 -2071 -86
rect -2109 -93 -2101 -88
rect -2101 -95 -2079 -93
rect -2069 -95 -2068 -88
rect -2325 -104 -2317 -96
rect -2079 -100 -2071 -95
rect -2325 -154 -2320 -104
rect -2317 -112 -2309 -104
rect -2074 -109 -2071 -100
rect -2069 -104 -2068 -100
rect -2109 -118 -2079 -115
rect -2309 -152 -2301 -142
rect -2317 -154 -2309 -152
rect -2000 -154 -1992 -84
rect -1846 -86 -1806 -84
rect -1854 -91 -1806 -87
rect -1854 -93 -1846 -91
rect -1846 -95 -1806 -93
rect -1806 -97 -1798 -95
rect -1846 -100 -1798 -97
rect -1846 -113 -1806 -102
rect -1671 -104 -1663 -96
rect -1663 -112 -1655 -104
rect -1854 -118 -1680 -114
rect -1655 -152 -1647 -142
rect -1663 -154 -1655 -152
rect -1642 -154 -1637 -84
rect -1619 -154 -1614 -84
rect -1530 -154 -1526 -84
rect -1506 -154 -1502 -84
rect -1482 -154 -1478 -84
rect -1458 -154 -1454 -84
rect -1434 -154 -1430 -84
rect -1410 -154 -1406 -84
rect -1386 -154 -1382 -84
rect -1362 -154 -1358 -84
rect -1338 -154 -1334 -84
rect -1290 -85 -1286 -84
rect -1325 -108 -1293 -105
rect -1325 -115 -1320 -108
rect -1307 -109 -1293 -108
rect -1290 -109 -1283 -85
rect -1315 -129 -1310 -115
rect -1314 -154 -1310 -129
rect -1266 -154 -1262 -84
rect -1242 -154 -1238 -84
rect -1218 -154 -1214 -84
rect -1194 -154 -1190 -84
rect -1170 -154 -1166 -84
rect -1146 -154 -1142 -84
rect -1122 -154 -1118 -84
rect -1098 -154 -1094 -84
rect -1074 -154 -1070 -84
rect -1050 -154 -1046 -84
rect -1026 -154 -1022 -84
rect -1002 -154 -998 -84
rect -989 -130 -955 -129
rect -954 -130 -950 -84
rect -930 -130 -926 -84
rect -906 -130 -902 -84
rect -882 -130 -878 -84
rect -858 -130 -854 -84
rect -834 -130 -830 -84
rect -810 -130 -806 -84
rect -786 -130 -782 -84
rect -762 -130 -758 -84
rect -738 -130 -734 -84
rect -714 -130 -710 -84
rect -690 -130 -686 -84
rect -666 -130 -662 -84
rect -642 -130 -638 -84
rect -618 -130 -614 -84
rect -594 -130 -590 -84
rect -570 -130 -566 -84
rect -546 -130 -542 -84
rect -522 -130 -518 -84
rect -498 -130 -494 -84
rect -474 -130 -470 -84
rect -450 -130 -446 -84
rect -426 -130 -422 -84
rect -402 -130 -398 -84
rect -378 -130 -374 -84
rect -354 -130 -350 -84
rect -330 -130 -326 -84
rect -306 -130 -302 -84
rect -282 -130 -278 -84
rect -258 -130 -254 -84
rect -234 -130 -230 -84
rect -210 -130 -206 -84
rect -186 -130 -182 -84
rect -162 -130 -158 -84
rect -138 -130 -134 -84
rect -114 -130 -110 -84
rect -90 -130 -86 -84
rect -66 -130 -62 -84
rect -42 -130 -38 -84
rect -18 -130 -14 -84
rect 6 -130 10 -84
rect 30 -130 34 -84
rect 54 -130 58 -84
rect 78 -130 82 -84
rect 102 -130 106 -84
rect 126 -130 130 -84
rect 150 -130 154 -84
rect 174 -130 178 -84
rect 198 -130 202 -84
rect 222 -130 226 -84
rect 246 -130 250 -84
rect 270 -130 274 -84
rect 294 -130 298 -84
rect 301 -85 315 -84
rect 318 -85 325 -61
rect 318 -130 322 -85
rect 342 -130 346 36
rect 355 -43 360 -33
rect 366 -43 370 36
rect 365 -57 370 -43
rect 355 -58 389 -57
rect 390 -58 394 36
rect 414 -58 418 36
rect 438 -58 442 36
rect 462 -58 466 36
rect 486 -58 490 36
rect 510 35 514 36
rect 510 -13 517 35
rect 510 -58 514 -13
rect 534 -58 538 36
rect 558 -58 562 36
rect 582 -58 586 36
rect 606 -58 610 36
rect 630 -58 634 36
rect 654 -58 658 36
rect 678 -58 682 36
rect 702 -58 706 36
rect 726 -58 730 36
rect 750 -58 754 36
rect 774 -58 778 36
rect 798 -58 802 36
rect 805 35 819 36
rect 822 11 829 59
rect 822 -58 826 11
rect 846 -58 850 84
rect 870 -58 874 84
rect 894 -58 898 84
rect 918 -58 922 84
rect 942 -58 946 84
rect 966 -58 970 84
rect 990 -58 994 84
rect 1014 -57 1018 84
rect 1027 29 1032 39
rect 1038 29 1042 84
rect 1051 77 1056 84
rect 1062 77 1066 84
rect 1061 63 1066 77
rect 1037 15 1042 29
rect 1003 -58 1037 -57
rect 355 -60 1037 -58
rect 355 -67 360 -60
rect 365 -81 370 -67
rect 366 -130 370 -81
rect 390 -109 394 -60
rect -989 -132 387 -130
rect -989 -139 -984 -132
rect -954 -133 -950 -132
rect -979 -153 -974 -139
rect -965 -143 -957 -139
rect -971 -153 -965 -143
rect -978 -154 -974 -153
rect -2393 -156 -957 -154
rect -2371 -250 -2366 -156
rect -2348 -250 -2343 -156
rect -2325 -218 -2320 -156
rect -2317 -158 -2309 -156
rect -2013 -158 -1992 -156
rect -1663 -158 -1655 -156
rect -2000 -159 -1983 -158
rect -2026 -168 -2021 -164
rect -2062 -169 -2061 -168
rect -2309 -180 -2301 -170
rect -2091 -176 -2061 -169
rect -2317 -186 -2309 -180
rect -2132 -185 -2131 -183
rect -2101 -185 -2092 -183
rect -2091 -184 -2071 -178
rect -2062 -180 -2045 -176
rect -2036 -180 -2031 -178
rect -2292 -194 -2071 -185
rect -2107 -199 -2104 -195
rect -2325 -226 -2317 -218
rect -2325 -246 -2320 -226
rect -2317 -234 -2309 -226
rect -2325 -250 -2317 -246
rect -2000 -250 -1992 -159
rect -1980 -176 -1932 -169
rect -1655 -180 -1647 -170
rect -1846 -194 -1680 -185
rect -1663 -186 -1655 -180
rect -1671 -226 -1663 -218
rect -1663 -234 -1655 -226
rect -1671 -250 -1663 -246
rect -1642 -250 -1637 -156
rect -1619 -250 -1614 -156
rect -1530 -250 -1526 -156
rect -1506 -250 -1502 -156
rect -1482 -250 -1478 -156
rect -1458 -250 -1454 -156
rect -1434 -250 -1430 -156
rect -1410 -250 -1406 -156
rect -1386 -250 -1382 -156
rect -1362 -250 -1358 -156
rect -1338 -250 -1334 -156
rect -1314 -250 -1310 -156
rect -1290 -202 -1283 -181
rect -1266 -202 -1262 -156
rect -1242 -202 -1238 -156
rect -1218 -202 -1214 -156
rect -1194 -202 -1190 -156
rect -1170 -202 -1166 -156
rect -1146 -202 -1142 -156
rect -1122 -202 -1118 -156
rect -1098 -202 -1094 -156
rect -1074 -202 -1070 -156
rect -1050 -202 -1046 -156
rect -1026 -202 -1022 -156
rect -1002 -202 -998 -156
rect -978 -202 -974 -156
rect -971 -157 -957 -156
rect -954 -157 -947 -133
rect -930 -202 -926 -132
rect -906 -202 -902 -132
rect -882 -202 -878 -132
rect -858 -202 -854 -132
rect -834 -202 -830 -132
rect -810 -202 -806 -132
rect -786 -202 -782 -132
rect -762 -202 -758 -132
rect -738 -202 -734 -132
rect -714 -202 -710 -132
rect -690 -202 -686 -132
rect -666 -202 -662 -132
rect -642 -202 -638 -132
rect -618 -202 -614 -132
rect -594 -202 -590 -132
rect -570 -202 -566 -132
rect -546 -202 -542 -132
rect -522 -202 -518 -132
rect -498 -202 -494 -132
rect -474 -202 -470 -132
rect -450 -202 -446 -132
rect -426 -202 -422 -132
rect -402 -202 -398 -132
rect -378 -202 -374 -132
rect -354 -202 -350 -132
rect -330 -202 -326 -132
rect -306 -202 -302 -132
rect -282 -202 -278 -132
rect -258 -202 -254 -132
rect -234 -202 -230 -132
rect -210 -202 -206 -132
rect -186 -202 -182 -132
rect -162 -202 -158 -132
rect -138 -202 -134 -132
rect -114 -202 -110 -132
rect -90 -202 -86 -132
rect -66 -202 -62 -132
rect -42 -202 -38 -132
rect -18 -202 -14 -132
rect 6 -202 10 -132
rect 30 -202 34 -132
rect 54 -202 58 -132
rect 78 -202 82 -132
rect 102 -202 106 -132
rect 126 -201 130 -132
rect 115 -202 149 -201
rect -1307 -204 149 -202
rect -1307 -205 -1293 -204
rect -1290 -205 -1283 -204
rect -1290 -250 -1286 -205
rect -1266 -250 -1262 -204
rect -1242 -250 -1238 -204
rect -1218 -250 -1214 -204
rect -1194 -250 -1190 -204
rect -1170 -250 -1166 -204
rect -1146 -250 -1142 -204
rect -1122 -250 -1118 -204
rect -1098 -250 -1094 -204
rect -1074 -250 -1070 -204
rect -1050 -250 -1046 -204
rect -1026 -250 -1022 -204
rect -1002 -250 -998 -204
rect -978 -250 -974 -204
rect -954 -229 -947 -205
rect -954 -250 -950 -229
rect -930 -250 -926 -204
rect -906 -250 -902 -204
rect -882 -250 -878 -204
rect -858 -250 -854 -204
rect -834 -250 -830 -204
rect -810 -250 -806 -204
rect -786 -250 -782 -204
rect -762 -250 -758 -204
rect -738 -250 -734 -204
rect -714 -250 -710 -204
rect -690 -250 -686 -204
rect -666 -250 -662 -204
rect -642 -250 -638 -204
rect -618 -250 -614 -204
rect -594 -250 -590 -204
rect -570 -250 -566 -204
rect -546 -250 -542 -204
rect -522 -250 -518 -204
rect -498 -250 -494 -204
rect -474 -250 -470 -204
rect -450 -250 -446 -204
rect -426 -250 -422 -204
rect -402 -250 -398 -204
rect -378 -250 -374 -204
rect -354 -250 -350 -204
rect -330 -250 -326 -204
rect -306 -250 -302 -204
rect -282 -250 -278 -204
rect -258 -250 -254 -204
rect -234 -250 -230 -204
rect -210 -250 -206 -204
rect -186 -250 -182 -204
rect -162 -250 -158 -204
rect -138 -250 -134 -204
rect -114 -250 -110 -204
rect -90 -250 -86 -204
rect -66 -250 -62 -204
rect -42 -250 -38 -204
rect -18 -250 -14 -204
rect 6 -250 10 -204
rect 30 -250 34 -204
rect 54 -250 58 -204
rect 78 -250 82 -204
rect 102 -250 106 -204
rect 115 -211 120 -204
rect 126 -211 130 -204
rect 125 -225 130 -211
rect 115 -226 149 -225
rect 150 -226 154 -132
rect 174 -226 178 -132
rect 198 -226 202 -132
rect 222 -226 226 -132
rect 246 -226 250 -132
rect 270 -226 274 -132
rect 294 -226 298 -132
rect 318 -226 322 -132
rect 342 -226 346 -132
rect 366 -226 370 -132
rect 373 -133 387 -132
rect 390 -154 397 -109
rect 414 -154 418 -60
rect 438 -154 442 -60
rect 462 -154 466 -60
rect 486 -154 490 -60
rect 510 -154 514 -60
rect 534 -154 538 -60
rect 558 -154 562 -60
rect 582 -154 586 -60
rect 606 -154 610 -60
rect 630 -154 634 -60
rect 654 -154 658 -60
rect 678 -154 682 -60
rect 702 -154 706 -60
rect 726 -154 730 -60
rect 739 -91 744 -81
rect 750 -91 754 -60
rect 749 -105 754 -91
rect 739 -154 773 -153
rect 373 -156 773 -154
rect 373 -157 387 -156
rect 390 -157 397 -156
rect 390 -226 394 -157
rect 414 -226 418 -156
rect 438 -226 442 -156
rect 462 -226 466 -156
rect 486 -226 490 -156
rect 510 -226 514 -156
rect 534 -226 538 -156
rect 558 -226 562 -156
rect 582 -226 586 -156
rect 606 -226 610 -156
rect 630 -226 634 -156
rect 654 -226 658 -156
rect 678 -226 682 -156
rect 702 -226 706 -156
rect 726 -226 730 -156
rect 739 -163 744 -156
rect 774 -157 778 -60
rect 749 -177 754 -163
rect 763 -167 771 -163
rect 757 -177 763 -167
rect 750 -226 754 -177
rect 774 -181 781 -157
rect 798 -226 802 -60
rect 822 -226 826 -60
rect 846 -226 850 -60
rect 870 -226 874 -60
rect 894 -226 898 -60
rect 918 -226 922 -60
rect 942 -225 946 -60
rect 955 -139 960 -129
rect 966 -139 970 -60
rect 979 -115 984 -105
rect 990 -115 994 -60
rect 1003 -67 1008 -60
rect 1014 -67 1018 -60
rect 1013 -81 1018 -67
rect 989 -129 994 -115
rect 965 -153 970 -139
rect 931 -226 965 -225
rect 115 -228 965 -226
rect 115 -235 120 -228
rect 125 -249 130 -235
rect 126 -250 130 -249
rect 150 -250 154 -228
rect 174 -250 178 -228
rect 198 -250 202 -228
rect 222 -250 226 -228
rect 246 -250 250 -228
rect 270 -250 274 -228
rect 294 -250 298 -228
rect 318 -250 322 -228
rect 342 -250 346 -228
rect 366 -250 370 -228
rect 390 -250 394 -228
rect 414 -250 418 -228
rect 438 -250 442 -228
rect 462 -250 466 -228
rect 486 -250 490 -228
rect 510 -250 514 -228
rect 534 -250 538 -228
rect 558 -250 562 -228
rect 582 -250 586 -228
rect 606 -250 610 -228
rect 630 -250 634 -228
rect 654 -250 658 -228
rect 678 -250 682 -228
rect 702 -250 706 -228
rect 726 -250 730 -228
rect 750 -250 754 -228
rect -2393 -252 771 -250
rect -2371 -298 -2366 -252
rect -2348 -298 -2343 -252
rect -2325 -260 -2317 -252
rect -2018 -253 -2004 -252
rect -2000 -253 -1992 -252
rect -2072 -254 -1928 -253
rect -2072 -260 -2053 -254
rect -2325 -276 -2320 -260
rect -2317 -262 -2309 -260
rect -2309 -274 -2301 -262
rect -2092 -269 -2062 -264
rect -2317 -276 -2309 -274
rect -2325 -288 -2317 -276
rect -2098 -282 -2096 -271
rect -2092 -282 -2084 -269
rect -2000 -270 -1992 -254
rect -1972 -260 -1928 -254
rect -1924 -260 -1918 -252
rect -1671 -260 -1663 -252
rect -1663 -262 -1655 -260
rect -2083 -280 -2062 -271
rect -2027 -272 -1992 -270
rect -2018 -280 -2002 -272
rect -2000 -280 -1992 -272
rect -2100 -287 -2096 -282
rect -2083 -287 -2053 -282
rect -2003 -284 -1990 -280
rect -1972 -282 -1964 -273
rect -1928 -274 -1924 -271
rect -1655 -274 -1647 -262
rect -1663 -276 -1655 -274
rect -2325 -298 -2320 -288
rect -2317 -290 -2309 -288
rect -2309 -298 -2301 -290
rect -2004 -294 -2003 -284
rect -2062 -298 -2012 -296
rect -2000 -298 -1992 -284
rect -1972 -287 -1924 -282
rect -1864 -287 -1796 -281
rect -1671 -288 -1663 -276
rect -1663 -290 -1655 -288
rect -1864 -298 -1796 -297
rect -1655 -298 -1647 -290
rect -1642 -298 -1637 -252
rect -1619 -298 -1614 -252
rect -1530 -298 -1526 -252
rect -1506 -298 -1502 -252
rect -1482 -298 -1478 -252
rect -1458 -298 -1454 -252
rect -1434 -298 -1430 -252
rect -1410 -298 -1406 -252
rect -1386 -298 -1382 -252
rect -1362 -298 -1358 -252
rect -1338 -298 -1334 -252
rect -1325 -283 -1320 -273
rect -1314 -283 -1310 -252
rect -1315 -297 -1310 -283
rect -1325 -298 -1291 -297
rect -2393 -300 -1291 -298
rect -2371 -346 -2366 -300
rect -2348 -346 -2343 -300
rect -2325 -304 -2320 -300
rect -2309 -302 -2301 -300
rect -2317 -304 -2309 -302
rect -2325 -316 -2317 -304
rect -2325 -346 -2320 -316
rect -2317 -318 -2309 -316
rect -2092 -330 -2062 -328
rect -2094 -334 -2062 -330
rect -2000 -346 -1992 -300
rect -1655 -302 -1647 -300
rect -1663 -304 -1655 -302
rect -1671 -316 -1663 -304
rect -1663 -318 -1655 -316
rect -1854 -330 -1806 -328
rect -1854 -334 -1680 -330
rect -1642 -346 -1637 -300
rect -1619 -346 -1614 -300
rect -1530 -346 -1526 -300
rect -1506 -346 -1502 -300
rect -1482 -346 -1478 -300
rect -1458 -346 -1454 -300
rect -1434 -346 -1430 -300
rect -1410 -346 -1406 -300
rect -1386 -346 -1382 -300
rect -1362 -346 -1358 -300
rect -1338 -346 -1334 -300
rect -1325 -307 -1320 -300
rect -1315 -321 -1310 -307
rect -1314 -346 -1310 -321
rect -1290 -346 -1286 -252
rect -1266 -346 -1262 -252
rect -1242 -346 -1238 -252
rect -1218 -346 -1214 -252
rect -1194 -346 -1190 -252
rect -1170 -346 -1166 -252
rect -1146 -346 -1142 -252
rect -1122 -346 -1118 -252
rect -1098 -346 -1094 -252
rect -1074 -346 -1070 -252
rect -1050 -346 -1046 -252
rect -1026 -346 -1022 -252
rect -1002 -346 -998 -252
rect -978 -346 -974 -252
rect -954 -346 -950 -252
rect -930 -346 -926 -252
rect -906 -346 -902 -252
rect -882 -346 -878 -252
rect -858 -346 -854 -252
rect -834 -346 -830 -252
rect -810 -346 -806 -252
rect -786 -346 -782 -252
rect -762 -346 -758 -252
rect -738 -346 -734 -252
rect -714 -346 -710 -252
rect -690 -346 -686 -252
rect -666 -346 -662 -252
rect -642 -346 -638 -252
rect -618 -346 -614 -252
rect -594 -346 -590 -252
rect -570 -346 -566 -252
rect -546 -346 -542 -252
rect -522 -346 -518 -252
rect -498 -346 -494 -252
rect -474 -346 -470 -252
rect -450 -346 -446 -252
rect -426 -346 -422 -252
rect -402 -346 -398 -252
rect -378 -346 -374 -252
rect -354 -346 -350 -252
rect -330 -346 -326 -252
rect -306 -346 -302 -252
rect -282 -346 -278 -252
rect -258 -346 -254 -252
rect -234 -346 -230 -252
rect -210 -346 -206 -252
rect -186 -346 -182 -252
rect -162 -346 -158 -252
rect -138 -346 -134 -252
rect -114 -346 -110 -252
rect -90 -346 -86 -252
rect -66 -346 -62 -252
rect -42 -346 -38 -252
rect -18 -346 -14 -252
rect 6 -346 10 -252
rect 30 -346 34 -252
rect 54 -346 58 -252
rect 78 -346 82 -252
rect 102 -346 106 -252
rect 126 -346 130 -252
rect 150 -277 154 -252
rect 150 -325 157 -277
rect 150 -346 154 -325
rect 174 -346 178 -252
rect 198 -346 202 -252
rect 222 -346 226 -252
rect 246 -346 250 -252
rect 270 -346 274 -252
rect 294 -346 298 -252
rect 318 -346 322 -252
rect 342 -346 346 -252
rect 366 -346 370 -252
rect 390 -346 394 -252
rect 414 -346 418 -252
rect 438 -346 442 -252
rect 462 -346 466 -252
rect 486 -346 490 -252
rect 510 -346 514 -252
rect 534 -346 538 -252
rect 558 -346 562 -252
rect 582 -346 586 -252
rect 606 -346 610 -252
rect 630 -346 634 -252
rect 654 -346 658 -252
rect 678 -346 682 -252
rect 702 -346 706 -252
rect 726 -346 730 -252
rect 750 -346 754 -252
rect 757 -253 771 -252
rect 774 -253 781 -229
rect 774 -346 778 -253
rect 798 -346 802 -228
rect 822 -346 826 -228
rect 846 -346 850 -228
rect 870 -346 874 -228
rect 894 -346 898 -228
rect 918 -346 922 -228
rect 931 -235 936 -228
rect 942 -235 946 -228
rect 941 -249 946 -235
rect 931 -259 936 -249
rect 941 -273 946 -259
rect 942 -346 946 -273
rect 955 -346 963 -345
rect -2393 -348 963 -346
rect -2371 -394 -2366 -348
rect -2348 -394 -2343 -348
rect -2325 -394 -2320 -348
rect -2309 -364 -2301 -354
rect -2317 -370 -2309 -364
rect -2097 -370 -2095 -361
rect -2309 -392 -2301 -382
rect -2097 -384 -2095 -380
rect -2292 -385 -2095 -384
rect -2097 -387 -2095 -385
rect -2084 -392 -2083 -349
rect -2069 -356 -2054 -354
rect -2054 -372 -2018 -370
rect -2054 -374 -2004 -372
rect -2059 -378 -2045 -374
rect -2054 -380 -2049 -378
rect -2317 -394 -2309 -392
rect -2084 -394 -2054 -392
rect -2044 -394 -2039 -380
rect -2025 -390 -2014 -384
rect -2000 -390 -1992 -348
rect -1920 -350 -1906 -348
rect -1977 -365 -1929 -359
rect -1655 -364 -1647 -354
rect -1977 -375 -1966 -365
rect -1663 -370 -1655 -364
rect -1977 -387 -1929 -385
rect -2033 -394 -1992 -390
rect -1655 -392 -1647 -382
rect -1663 -394 -1655 -392
rect -1642 -394 -1637 -348
rect -1619 -394 -1614 -348
rect -1530 -394 -1526 -348
rect -1506 -394 -1502 -348
rect -1482 -394 -1478 -348
rect -1458 -393 -1454 -348
rect -1469 -394 -1435 -393
rect -2393 -396 -1435 -394
rect -2371 -490 -2366 -396
rect -2348 -490 -2343 -396
rect -2325 -430 -2320 -396
rect -2317 -398 -2309 -396
rect -2084 -409 -2083 -396
rect -2084 -410 -2054 -409
rect -2325 -438 -2317 -430
rect -2325 -490 -2320 -438
rect -2317 -446 -2309 -438
rect -2117 -447 -2095 -437
rect -2045 -440 -2037 -426
rect -2309 -486 -2301 -478
rect -2317 -490 -2309 -486
rect -2000 -490 -1992 -396
rect -1663 -398 -1655 -396
rect -1969 -447 -1929 -435
rect -1671 -438 -1663 -430
rect -1663 -446 -1655 -438
rect -1655 -486 -1647 -478
rect -1663 -490 -1655 -486
rect -1642 -490 -1637 -396
rect -1619 -490 -1614 -396
rect -1530 -490 -1526 -396
rect -1506 -490 -1502 -396
rect -1482 -490 -1478 -396
rect -1469 -403 -1464 -396
rect -1458 -403 -1454 -396
rect -1459 -417 -1454 -403
rect -1469 -442 -1435 -441
rect -1434 -442 -1430 -348
rect -1410 -442 -1406 -348
rect -1386 -442 -1382 -348
rect -1362 -442 -1358 -348
rect -1338 -442 -1334 -348
rect -1314 -442 -1310 -348
rect -1290 -349 -1286 -348
rect -1290 -397 -1283 -349
rect -1290 -442 -1286 -397
rect -1266 -442 -1262 -348
rect -1242 -442 -1238 -348
rect -1218 -442 -1214 -348
rect -1194 -442 -1190 -348
rect -1170 -442 -1166 -348
rect -1146 -442 -1142 -348
rect -1122 -442 -1118 -348
rect -1098 -442 -1094 -348
rect -1074 -442 -1070 -348
rect -1050 -442 -1046 -348
rect -1026 -442 -1022 -348
rect -1013 -427 -1008 -417
rect -1002 -427 -998 -348
rect -1003 -441 -998 -427
rect -978 -442 -974 -348
rect -954 -442 -950 -348
rect -930 -442 -926 -348
rect -906 -442 -902 -348
rect -882 -442 -878 -348
rect -858 -442 -854 -348
rect -834 -442 -830 -348
rect -810 -442 -806 -348
rect -786 -442 -782 -348
rect -762 -442 -758 -348
rect -738 -442 -734 -348
rect -714 -442 -710 -348
rect -690 -442 -686 -348
rect -666 -442 -662 -348
rect -642 -442 -638 -348
rect -618 -442 -614 -348
rect -594 -442 -590 -348
rect -570 -442 -566 -348
rect -546 -442 -542 -348
rect -522 -442 -518 -348
rect -498 -442 -494 -348
rect -474 -442 -470 -348
rect -450 -442 -446 -348
rect -426 -442 -422 -348
rect -402 -442 -398 -348
rect -378 -442 -374 -348
rect -354 -442 -350 -348
rect -330 -442 -326 -348
rect -306 -442 -302 -348
rect -282 -442 -278 -348
rect -258 -442 -254 -348
rect -234 -442 -230 -348
rect -210 -442 -206 -348
rect -186 -442 -182 -348
rect -162 -442 -158 -348
rect -138 -442 -134 -348
rect -114 -442 -110 -348
rect -90 -442 -86 -348
rect -66 -442 -62 -348
rect -42 -442 -38 -348
rect -18 -442 -14 -348
rect 6 -442 10 -348
rect 30 -442 34 -348
rect 54 -442 58 -348
rect 78 -442 82 -348
rect 102 -442 106 -348
rect 126 -442 130 -348
rect 150 -442 154 -348
rect 174 -442 178 -348
rect 198 -442 202 -348
rect 222 -442 226 -348
rect 246 -442 250 -348
rect 270 -442 274 -348
rect 294 -442 298 -348
rect 318 -442 322 -348
rect 342 -442 346 -348
rect 366 -442 370 -348
rect 390 -442 394 -348
rect 414 -442 418 -348
rect 438 -442 442 -348
rect 462 -442 466 -348
rect 486 -442 490 -348
rect 510 -442 514 -348
rect 534 -442 538 -348
rect 558 -442 562 -348
rect 582 -442 586 -348
rect 606 -442 610 -348
rect 630 -442 634 -348
rect 654 -442 658 -348
rect 678 -442 682 -348
rect 702 -442 706 -348
rect 726 -442 730 -348
rect 750 -442 754 -348
rect 774 -442 778 -348
rect 798 -442 802 -348
rect 822 -442 826 -348
rect 846 -442 850 -348
rect 870 -442 874 -348
rect 894 -442 898 -348
rect 918 -442 922 -348
rect 942 -442 946 -348
rect 949 -349 963 -348
rect 955 -355 960 -349
rect 965 -369 970 -355
rect 966 -441 970 -369
rect 955 -442 987 -441
rect -1469 -444 987 -442
rect -1469 -451 -1464 -444
rect -1459 -465 -1454 -451
rect -1458 -490 -1454 -465
rect -1434 -469 -1430 -444
rect -2393 -492 -2026 -490
rect -2021 -492 -1437 -490
rect -2371 -586 -2366 -492
rect -2348 -586 -2343 -492
rect -2325 -554 -2320 -492
rect -2317 -494 -2309 -492
rect -2309 -514 -2301 -506
rect -2317 -522 -2309 -514
rect -2123 -519 -2116 -514
rect -2123 -521 -2092 -519
rect -2091 -520 -2087 -504
rect -2026 -512 -2021 -500
rect -2037 -516 -2021 -512
rect -2292 -523 -2087 -521
rect -2123 -525 -2116 -523
rect -2325 -562 -2317 -554
rect -2325 -582 -2320 -562
rect -2317 -570 -2309 -562
rect -2325 -586 -2317 -582
rect -2000 -586 -1992 -492
rect -1663 -494 -1655 -492
rect -1969 -520 -1932 -504
rect -1655 -514 -1647 -506
rect -1969 -523 -1680 -521
rect -1663 -522 -1655 -514
rect -1671 -562 -1663 -554
rect -1663 -570 -1655 -562
rect -1671 -586 -1663 -582
rect -1642 -586 -1637 -492
rect -1619 -586 -1614 -492
rect -1530 -586 -1526 -492
rect -1506 -586 -1502 -492
rect -1482 -586 -1478 -492
rect -1458 -586 -1454 -492
rect -1451 -493 -1437 -492
rect -1434 -493 -1427 -469
rect -1434 -538 -1427 -517
rect -1410 -538 -1406 -444
rect -1386 -538 -1382 -444
rect -1362 -538 -1358 -444
rect -1338 -538 -1334 -444
rect -1314 -538 -1310 -444
rect -1290 -538 -1286 -444
rect -1266 -538 -1262 -444
rect -1242 -538 -1238 -444
rect -1218 -538 -1214 -444
rect -1194 -538 -1190 -444
rect -1170 -538 -1166 -444
rect -1146 -538 -1142 -444
rect -1122 -538 -1118 -444
rect -1098 -538 -1094 -444
rect -1074 -537 -1070 -444
rect -1085 -538 -1051 -537
rect -1451 -540 -1051 -538
rect -1451 -541 -1437 -540
rect -1434 -541 -1427 -540
rect -1434 -586 -1430 -541
rect -1410 -586 -1406 -540
rect -1386 -586 -1382 -540
rect -1362 -586 -1358 -540
rect -1338 -586 -1334 -540
rect -1314 -586 -1310 -540
rect -1290 -586 -1286 -540
rect -1266 -586 -1262 -540
rect -1242 -586 -1238 -540
rect -1218 -586 -1214 -540
rect -1194 -586 -1190 -540
rect -1170 -586 -1166 -540
rect -1146 -586 -1142 -540
rect -1122 -586 -1118 -540
rect -1098 -586 -1094 -540
rect -1085 -547 -1080 -540
rect -1074 -547 -1070 -540
rect -1075 -561 -1070 -547
rect -1085 -571 -1080 -561
rect -1075 -585 -1070 -571
rect -1074 -586 -1070 -585
rect -1050 -586 -1046 -444
rect -1026 -586 -1022 -444
rect -1013 -475 -1008 -465
rect -1003 -489 -998 -475
rect -1002 -586 -998 -489
rect -978 -493 -974 -444
rect -978 -517 -971 -493
rect -978 -562 -971 -541
rect -954 -562 -950 -444
rect -930 -562 -926 -444
rect -906 -562 -902 -444
rect -882 -562 -878 -444
rect -858 -562 -854 -444
rect -834 -562 -830 -444
rect -810 -562 -806 -444
rect -786 -562 -782 -444
rect -762 -562 -758 -444
rect -738 -562 -734 -444
rect -714 -562 -710 -444
rect -690 -562 -686 -444
rect -666 -562 -662 -444
rect -642 -562 -638 -444
rect -618 -562 -614 -444
rect -594 -562 -590 -444
rect -570 -562 -566 -444
rect -546 -562 -542 -444
rect -522 -562 -518 -444
rect -498 -562 -494 -444
rect -474 -562 -470 -444
rect -450 -562 -446 -444
rect -426 -562 -422 -444
rect -402 -562 -398 -444
rect -378 -562 -374 -444
rect -354 -562 -350 -444
rect -330 -562 -326 -444
rect -306 -562 -302 -444
rect -282 -562 -278 -444
rect -258 -562 -254 -444
rect -234 -562 -230 -444
rect -210 -562 -206 -444
rect -186 -562 -182 -444
rect -162 -562 -158 -444
rect -138 -562 -134 -444
rect -114 -562 -110 -444
rect -90 -562 -86 -444
rect -66 -562 -62 -444
rect -42 -562 -38 -444
rect -18 -562 -14 -444
rect 6 -562 10 -444
rect 30 -562 34 -444
rect 54 -562 58 -444
rect 78 -562 82 -444
rect 102 -562 106 -444
rect 126 -562 130 -444
rect 150 -562 154 -444
rect 174 -562 178 -444
rect 198 -562 202 -444
rect 222 -562 226 -444
rect 246 -562 250 -444
rect 270 -562 274 -444
rect 294 -562 298 -444
rect 318 -562 322 -444
rect 342 -562 346 -444
rect 366 -562 370 -444
rect 390 -562 394 -444
rect 414 -562 418 -444
rect 438 -562 442 -444
rect 462 -562 466 -444
rect 486 -562 490 -444
rect 510 -562 514 -444
rect 534 -562 538 -444
rect 558 -562 562 -444
rect 582 -562 586 -444
rect 606 -562 610 -444
rect 630 -562 634 -444
rect 654 -562 658 -444
rect 678 -562 682 -444
rect 702 -562 706 -444
rect 726 -562 730 -444
rect 750 -562 754 -444
rect 774 -562 778 -444
rect 798 -562 802 -444
rect 822 -562 826 -444
rect 846 -562 850 -444
rect 870 -562 874 -444
rect 894 -562 898 -444
rect 918 -562 922 -444
rect 931 -475 936 -465
rect 942 -475 946 -444
rect 955 -451 960 -444
rect 966 -451 970 -444
rect 973 -445 987 -444
rect 965 -465 970 -451
rect 941 -489 946 -475
rect 931 -499 936 -489
rect 941 -513 946 -499
rect 942 -561 946 -513
rect 931 -562 963 -561
rect -995 -564 963 -562
rect -995 -565 -981 -564
rect -978 -565 -971 -564
rect -978 -586 -974 -565
rect -954 -586 -950 -564
rect -930 -586 -926 -564
rect -906 -586 -902 -564
rect -882 -586 -878 -564
rect -858 -586 -854 -564
rect -834 -586 -830 -564
rect -810 -586 -806 -564
rect -786 -586 -782 -564
rect -762 -586 -758 -564
rect -738 -586 -734 -564
rect -714 -586 -710 -564
rect -690 -586 -686 -564
rect -666 -586 -662 -564
rect -642 -586 -638 -564
rect -618 -586 -614 -564
rect -594 -586 -590 -564
rect -570 -586 -566 -564
rect -546 -586 -542 -564
rect -522 -586 -518 -564
rect -498 -586 -494 -564
rect -474 -586 -470 -564
rect -450 -586 -446 -564
rect -426 -586 -422 -564
rect -402 -586 -398 -564
rect -378 -586 -374 -564
rect -354 -586 -350 -564
rect -330 -586 -326 -564
rect -306 -586 -302 -564
rect -282 -586 -278 -564
rect -258 -586 -254 -564
rect -234 -586 -230 -564
rect -210 -586 -206 -564
rect -186 -586 -182 -564
rect -162 -586 -158 -564
rect -138 -586 -134 -564
rect -114 -586 -110 -564
rect -90 -586 -86 -564
rect -66 -586 -62 -564
rect -42 -586 -38 -564
rect -18 -586 -14 -564
rect 6 -586 10 -564
rect 30 -586 34 -564
rect 54 -586 58 -564
rect 78 -586 82 -564
rect 102 -586 106 -564
rect 126 -586 130 -564
rect 150 -586 154 -564
rect 174 -586 178 -564
rect 198 -586 202 -564
rect 222 -586 226 -564
rect 246 -586 250 -564
rect 270 -586 274 -564
rect 294 -586 298 -564
rect 318 -586 322 -564
rect 342 -586 346 -564
rect 366 -586 370 -564
rect 390 -586 394 -564
rect 414 -586 418 -564
rect 438 -586 442 -564
rect 462 -586 466 -564
rect 486 -586 490 -564
rect 510 -586 514 -564
rect 534 -586 538 -564
rect 558 -586 562 -564
rect 582 -586 586 -564
rect 606 -586 610 -564
rect 630 -586 634 -564
rect 654 -586 658 -564
rect 678 -586 682 -564
rect 702 -585 706 -564
rect 691 -586 725 -585
rect -2393 -588 725 -586
rect -2371 -634 -2366 -588
rect -2348 -634 -2343 -588
rect -2325 -596 -2317 -588
rect -2018 -589 -2004 -588
rect -2000 -589 -1992 -588
rect -2072 -590 -1928 -589
rect -2072 -596 -2053 -590
rect -2325 -612 -2320 -596
rect -2317 -598 -2309 -596
rect -2309 -610 -2301 -598
rect -2092 -605 -2062 -600
rect -2317 -612 -2309 -610
rect -2325 -624 -2317 -612
rect -2098 -618 -2096 -607
rect -2092 -618 -2084 -605
rect -2000 -606 -1992 -590
rect -1972 -596 -1928 -590
rect -1924 -596 -1918 -588
rect -1671 -596 -1663 -588
rect -1663 -598 -1655 -596
rect -2083 -616 -2062 -607
rect -2027 -608 -1992 -606
rect -2018 -616 -2002 -608
rect -2000 -616 -1992 -608
rect -2100 -623 -2096 -618
rect -2083 -623 -2053 -618
rect -2003 -620 -1990 -616
rect -1972 -618 -1964 -609
rect -1928 -610 -1924 -607
rect -1655 -610 -1647 -598
rect -1663 -612 -1655 -610
rect -2325 -634 -2320 -624
rect -2317 -626 -2309 -624
rect -2309 -634 -2301 -626
rect -2004 -630 -2003 -620
rect -2062 -634 -2012 -632
rect -2000 -634 -1992 -620
rect -1972 -623 -1924 -618
rect -1864 -623 -1796 -617
rect -1671 -624 -1663 -612
rect -1663 -626 -1655 -624
rect -1864 -634 -1796 -633
rect -1655 -634 -1647 -626
rect -1642 -634 -1637 -588
rect -1619 -634 -1614 -588
rect -1530 -634 -1526 -588
rect -1506 -634 -1502 -588
rect -1482 -634 -1478 -588
rect -1458 -634 -1454 -588
rect -1434 -634 -1430 -588
rect -1410 -634 -1406 -588
rect -1386 -634 -1382 -588
rect -1362 -634 -1358 -588
rect -1338 -634 -1334 -588
rect -1314 -634 -1310 -588
rect -1290 -634 -1286 -588
rect -1266 -634 -1262 -588
rect -1242 -634 -1238 -588
rect -1229 -619 -1224 -609
rect -1218 -619 -1214 -588
rect -1219 -633 -1214 -619
rect -1194 -634 -1190 -588
rect -1170 -634 -1166 -588
rect -1146 -634 -1142 -588
rect -1122 -634 -1118 -588
rect -1098 -634 -1094 -588
rect -1074 -634 -1070 -588
rect -1050 -613 -1046 -588
rect -2393 -636 -1053 -634
rect -2371 -682 -2366 -636
rect -2348 -682 -2343 -636
rect -2325 -640 -2320 -636
rect -2309 -638 -2301 -636
rect -2317 -640 -2309 -638
rect -2325 -652 -2317 -640
rect -2325 -672 -2320 -652
rect -2317 -654 -2309 -652
rect -2092 -666 -2062 -664
rect -2094 -670 -2062 -666
rect -2325 -682 -2317 -672
rect -2095 -680 -2084 -676
rect -2000 -679 -1992 -636
rect -1655 -638 -1647 -636
rect -1663 -640 -1655 -638
rect -1671 -652 -1663 -640
rect -1663 -654 -1655 -652
rect -1854 -666 -1806 -664
rect -1854 -670 -1680 -666
rect -2119 -682 -2069 -680
rect -2054 -682 -1892 -679
rect -1671 -682 -1663 -672
rect -1642 -682 -1637 -636
rect -1619 -682 -1614 -636
rect -1530 -682 -1526 -636
rect -1506 -682 -1502 -636
rect -1482 -682 -1478 -636
rect -1458 -682 -1454 -636
rect -1434 -682 -1430 -636
rect -1410 -682 -1406 -636
rect -1386 -682 -1382 -636
rect -1362 -682 -1358 -636
rect -1338 -682 -1334 -636
rect -1314 -682 -1310 -636
rect -1290 -682 -1286 -636
rect -1266 -682 -1262 -636
rect -1242 -682 -1238 -636
rect -1229 -667 -1224 -657
rect -1219 -681 -1214 -667
rect -1194 -681 -1190 -636
rect -1218 -682 -1214 -681
rect -1205 -682 -1171 -681
rect -2393 -684 -1171 -682
rect -2371 -706 -2366 -684
rect -2348 -706 -2343 -684
rect -2325 -688 -2317 -684
rect -2325 -704 -2320 -688
rect -2309 -700 -2301 -688
rect -2095 -690 -2084 -684
rect -2054 -685 -1906 -684
rect -2054 -686 -2036 -685
rect -2084 -692 -2079 -690
rect -2317 -704 -2309 -700
rect -2092 -701 -2079 -694
rect -2000 -698 -1992 -685
rect -1920 -686 -1906 -685
rect -1671 -688 -1663 -684
rect -1846 -692 -1806 -690
rect -1854 -698 -1806 -694
rect -2054 -701 -1982 -698
rect -1966 -701 -1806 -698
rect -1655 -700 -1647 -688
rect -2003 -704 -1992 -701
rect -1904 -703 -1902 -701
rect -1854 -703 -1846 -701
rect -2325 -706 -2317 -704
rect -2033 -706 -1992 -704
rect -1854 -705 -1806 -703
rect -1663 -704 -1655 -700
rect -1864 -706 -1796 -705
rect -1671 -706 -1663 -704
rect -1642 -706 -1637 -684
rect -1619 -706 -1614 -684
rect -1530 -706 -1526 -684
rect -1506 -706 -1502 -684
rect -1482 -706 -1478 -684
rect -1458 -706 -1454 -684
rect -1434 -706 -1430 -684
rect -1410 -706 -1406 -684
rect -1386 -706 -1382 -684
rect -1362 -706 -1358 -684
rect -1338 -706 -1334 -684
rect -1314 -706 -1310 -684
rect -1290 -706 -1286 -684
rect -1266 -706 -1262 -684
rect -1242 -706 -1238 -684
rect -1218 -706 -1214 -684
rect -1205 -691 -1200 -684
rect -1194 -685 -1190 -684
rect -1194 -691 -1187 -685
rect -1195 -705 -1187 -691
rect -2393 -708 -1197 -706
rect -2371 -730 -2366 -708
rect -2348 -730 -2343 -708
rect -2325 -716 -2317 -708
rect -2079 -711 -2018 -708
rect -2003 -709 -1966 -708
rect -2000 -710 -1982 -709
rect -2000 -711 -1992 -710
rect -2084 -715 -2009 -711
rect -2028 -716 -2009 -715
rect -2000 -715 -1854 -711
rect -1846 -715 -1798 -708
rect -2325 -730 -2320 -716
rect -2309 -728 -2301 -716
rect -2028 -718 -2018 -716
rect -2092 -728 -2084 -721
rect -2023 -725 -2014 -718
rect -2000 -725 -1992 -715
rect -1671 -716 -1663 -708
rect -1846 -719 -1806 -717
rect -1854 -725 -1806 -721
rect -2054 -728 -1806 -725
rect -1655 -728 -1647 -716
rect -2317 -730 -2309 -728
rect -2054 -730 -2024 -728
rect -2000 -730 -1992 -728
rect -1663 -730 -1655 -728
rect -1642 -730 -1637 -708
rect -1619 -730 -1614 -708
rect -1530 -730 -1526 -708
rect -1506 -730 -1502 -708
rect -1482 -730 -1478 -708
rect -1458 -730 -1454 -708
rect -1434 -730 -1430 -708
rect -1410 -730 -1406 -708
rect -1386 -730 -1382 -708
rect -1362 -730 -1358 -708
rect -1338 -730 -1334 -708
rect -1314 -730 -1310 -708
rect -1290 -730 -1286 -708
rect -1266 -730 -1262 -708
rect -1242 -730 -1238 -708
rect -1218 -730 -1214 -708
rect -1211 -709 -1197 -708
rect -1205 -730 -1171 -729
rect -1170 -730 -1166 -636
rect -1146 -730 -1142 -636
rect -1122 -730 -1118 -636
rect -1098 -730 -1094 -636
rect -1074 -730 -1070 -636
rect -1067 -637 -1053 -636
rect -1050 -658 -1043 -613
rect -1026 -658 -1022 -588
rect -1002 -658 -998 -588
rect -978 -658 -974 -588
rect -954 -658 -950 -588
rect -930 -658 -926 -588
rect -906 -658 -902 -588
rect -882 -658 -878 -588
rect -858 -658 -854 -588
rect -834 -658 -830 -588
rect -810 -658 -806 -588
rect -786 -658 -782 -588
rect -762 -658 -758 -588
rect -738 -658 -734 -588
rect -725 -643 -720 -633
rect -714 -643 -710 -588
rect -715 -657 -710 -643
rect -690 -658 -686 -588
rect -666 -658 -662 -588
rect -642 -658 -638 -588
rect -618 -658 -614 -588
rect -594 -658 -590 -588
rect -570 -658 -566 -588
rect -546 -658 -542 -588
rect -522 -658 -518 -588
rect -498 -658 -494 -588
rect -474 -658 -470 -588
rect -450 -658 -446 -588
rect -426 -658 -422 -588
rect -402 -658 -398 -588
rect -378 -658 -374 -588
rect -354 -658 -350 -588
rect -330 -658 -326 -588
rect -306 -658 -302 -588
rect -282 -658 -278 -588
rect -258 -658 -254 -588
rect -234 -658 -230 -588
rect -210 -658 -206 -588
rect -186 -658 -182 -588
rect -162 -658 -158 -588
rect -138 -658 -134 -588
rect -114 -658 -110 -588
rect -90 -658 -86 -588
rect -66 -658 -62 -588
rect -42 -658 -38 -588
rect -18 -658 -14 -588
rect 6 -658 10 -588
rect 30 -658 34 -588
rect 54 -658 58 -588
rect 78 -658 82 -588
rect 102 -658 106 -588
rect 126 -658 130 -588
rect 150 -658 154 -588
rect 174 -658 178 -588
rect 198 -658 202 -588
rect 222 -658 226 -588
rect 246 -658 250 -588
rect 270 -658 274 -588
rect 294 -658 298 -588
rect 318 -658 322 -588
rect 342 -658 346 -588
rect 366 -658 370 -588
rect 390 -658 394 -588
rect 414 -658 418 -588
rect 438 -658 442 -588
rect 462 -658 466 -588
rect 486 -658 490 -588
rect 510 -658 514 -588
rect 534 -658 538 -588
rect 558 -658 562 -588
rect 582 -658 586 -588
rect 606 -658 610 -588
rect 630 -658 634 -588
rect 654 -658 658 -588
rect 678 -658 682 -588
rect 691 -595 696 -588
rect 702 -595 706 -588
rect 701 -609 706 -595
rect 691 -619 696 -609
rect 701 -633 706 -619
rect 702 -658 706 -633
rect 726 -658 730 -564
rect 750 -658 754 -564
rect 774 -658 778 -564
rect 798 -658 802 -564
rect 822 -658 826 -564
rect 846 -658 850 -564
rect 870 -658 874 -564
rect 894 -657 898 -564
rect 907 -619 912 -609
rect 918 -619 922 -564
rect 931 -571 936 -564
rect 942 -571 946 -564
rect 949 -565 963 -564
rect 941 -585 946 -571
rect 955 -575 963 -571
rect 949 -585 955 -575
rect 917 -633 922 -619
rect 883 -658 917 -657
rect -1067 -660 917 -658
rect -1067 -661 -1053 -660
rect -1050 -661 -1043 -660
rect -1050 -730 -1046 -661
rect -1026 -730 -1022 -660
rect -1002 -730 -998 -660
rect -978 -730 -974 -660
rect -954 -730 -950 -660
rect -930 -730 -926 -660
rect -906 -730 -902 -660
rect -882 -730 -878 -660
rect -858 -730 -854 -660
rect -834 -730 -830 -660
rect -810 -730 -806 -660
rect -786 -730 -782 -660
rect -762 -730 -758 -660
rect -738 -730 -734 -660
rect -725 -682 -691 -681
rect -690 -682 -686 -660
rect -666 -682 -662 -660
rect -642 -682 -638 -660
rect -618 -682 -614 -660
rect -594 -682 -590 -660
rect -570 -682 -566 -660
rect -546 -682 -542 -660
rect -522 -682 -518 -660
rect -498 -682 -494 -660
rect -474 -682 -470 -660
rect -450 -682 -446 -660
rect -426 -682 -422 -660
rect -402 -682 -398 -660
rect -378 -682 -374 -660
rect -354 -682 -350 -660
rect -330 -682 -326 -660
rect -306 -682 -302 -660
rect -282 -682 -278 -660
rect -258 -682 -254 -660
rect -234 -682 -230 -660
rect -210 -682 -206 -660
rect -186 -682 -182 -660
rect -162 -682 -158 -660
rect -138 -682 -134 -660
rect -114 -682 -110 -660
rect -90 -682 -86 -660
rect -66 -682 -62 -660
rect -42 -682 -38 -660
rect -18 -682 -14 -660
rect 6 -682 10 -660
rect 30 -682 34 -660
rect 54 -682 58 -660
rect 78 -682 82 -660
rect 102 -682 106 -660
rect 126 -682 130 -660
rect 150 -682 154 -660
rect 174 -682 178 -660
rect 198 -682 202 -660
rect 222 -682 226 -660
rect 246 -682 250 -660
rect 270 -682 274 -660
rect 294 -682 298 -660
rect 318 -682 322 -660
rect 342 -682 346 -660
rect 366 -682 370 -660
rect 390 -682 394 -660
rect 414 -682 418 -660
rect 438 -682 442 -660
rect 462 -682 466 -660
rect 486 -682 490 -660
rect 510 -682 514 -660
rect 534 -682 538 -660
rect 558 -682 562 -660
rect 582 -682 586 -660
rect 606 -682 610 -660
rect 630 -682 634 -660
rect 654 -682 658 -660
rect 678 -682 682 -660
rect 702 -682 706 -660
rect 726 -661 730 -660
rect -725 -684 723 -682
rect -725 -691 -720 -684
rect -715 -705 -710 -691
rect -714 -730 -710 -705
rect -690 -709 -686 -684
rect -2393 -732 -2064 -730
rect -2060 -732 -693 -730
rect -2371 -778 -2366 -732
rect -2348 -778 -2343 -732
rect -2325 -744 -2317 -732
rect -2060 -735 -2054 -732
rect -2084 -742 -2054 -735
rect -2050 -738 -2044 -736
rect -2325 -764 -2320 -744
rect -2064 -746 -2054 -742
rect -2325 -772 -2317 -764
rect -2101 -769 -2071 -766
rect -2325 -778 -2320 -772
rect -2317 -778 -2309 -772
rect -2000 -774 -1992 -732
rect -1846 -733 -1806 -732
rect -1846 -742 -1798 -735
rect -1671 -744 -1663 -732
rect -1846 -746 -1806 -744
rect -1854 -760 -1680 -756
rect -1846 -769 -1798 -766
rect -2079 -775 -2043 -774
rect -2007 -775 -1991 -774
rect -2079 -776 -2071 -775
rect -2079 -778 -2029 -776
rect -2011 -778 -1991 -775
rect -1846 -777 -1806 -771
rect -1671 -772 -1663 -764
rect -1864 -778 -1796 -777
rect -1663 -778 -1655 -772
rect -1642 -778 -1637 -732
rect -1619 -778 -1614 -732
rect -1530 -778 -1526 -732
rect -1506 -778 -1502 -732
rect -1482 -778 -1478 -732
rect -1458 -778 -1454 -732
rect -1434 -778 -1430 -732
rect -1410 -778 -1406 -732
rect -1386 -778 -1382 -732
rect -1362 -778 -1358 -732
rect -1338 -778 -1334 -732
rect -1314 -778 -1310 -732
rect -1290 -778 -1286 -732
rect -1266 -778 -1262 -732
rect -1242 -778 -1238 -732
rect -1218 -778 -1214 -732
rect -1195 -753 -1187 -739
rect -1194 -754 -1187 -753
rect -1170 -754 -1166 -732
rect -1146 -754 -1142 -732
rect -1122 -754 -1118 -732
rect -1098 -754 -1094 -732
rect -1074 -754 -1070 -732
rect -1050 -754 -1046 -732
rect -1026 -754 -1022 -732
rect -1002 -754 -998 -732
rect -978 -754 -974 -732
rect -954 -754 -950 -732
rect -930 -754 -926 -732
rect -906 -754 -902 -732
rect -882 -754 -878 -732
rect -858 -754 -854 -732
rect -834 -754 -830 -732
rect -810 -754 -806 -732
rect -786 -754 -782 -732
rect -762 -754 -758 -732
rect -738 -754 -734 -732
rect -714 -754 -710 -732
rect -707 -733 -693 -732
rect -690 -733 -683 -709
rect -666 -754 -662 -684
rect -642 -754 -638 -684
rect -629 -715 -624 -705
rect -618 -715 -614 -684
rect -619 -729 -614 -715
rect -594 -754 -590 -684
rect -570 -754 -566 -684
rect -546 -754 -542 -684
rect -522 -754 -518 -684
rect -498 -754 -494 -684
rect -474 -754 -470 -684
rect -450 -754 -446 -684
rect -426 -754 -422 -684
rect -402 -754 -398 -684
rect -378 -754 -374 -684
rect -354 -754 -350 -684
rect -341 -739 -336 -729
rect -330 -739 -326 -684
rect -331 -753 -326 -739
rect -306 -754 -302 -684
rect -282 -754 -278 -684
rect -258 -754 -254 -684
rect -234 -754 -230 -684
rect -210 -754 -206 -684
rect -186 -754 -182 -684
rect -162 -754 -158 -684
rect -138 -754 -134 -684
rect -114 -754 -110 -684
rect -90 -754 -86 -684
rect -66 -754 -62 -684
rect -42 -754 -38 -684
rect -18 -754 -14 -684
rect 6 -754 10 -684
rect 30 -754 34 -684
rect 54 -754 58 -684
rect 78 -754 82 -684
rect 102 -754 106 -684
rect 126 -754 130 -684
rect 150 -754 154 -684
rect 174 -754 178 -684
rect 198 -754 202 -684
rect 222 -754 226 -684
rect 246 -753 250 -684
rect 235 -754 269 -753
rect -1211 -756 269 -754
rect -1211 -757 -1197 -756
rect -1194 -757 -1187 -756
rect -1170 -757 -1166 -756
rect -1194 -778 -1190 -757
rect -2393 -780 -1173 -778
rect -2371 -826 -2366 -780
rect -2348 -826 -2343 -780
rect -2325 -792 -2320 -780
rect -2079 -782 -2071 -780
rect -2072 -784 -2071 -782
rect -2109 -789 -2101 -784
rect -2101 -791 -2079 -789
rect -2069 -791 -2068 -784
rect -2325 -800 -2317 -792
rect -2079 -796 -2071 -791
rect -2325 -820 -2320 -800
rect -2317 -808 -2309 -800
rect -2074 -805 -2071 -796
rect -2069 -800 -2068 -796
rect -2109 -814 -2079 -811
rect -2325 -826 -2317 -820
rect -2080 -826 -2071 -825
rect -2000 -826 -1992 -780
rect -1846 -782 -1806 -780
rect -1854 -787 -1806 -783
rect -1854 -789 -1846 -787
rect -1846 -791 -1806 -789
rect -1806 -793 -1798 -791
rect -1846 -796 -1798 -793
rect -1846 -809 -1806 -798
rect -1671 -800 -1663 -792
rect -1663 -808 -1655 -800
rect -1854 -814 -1680 -810
rect -1926 -826 -1892 -823
rect -1671 -826 -1663 -820
rect -1642 -826 -1637 -780
rect -1619 -826 -1614 -780
rect -1530 -826 -1526 -780
rect -1506 -826 -1502 -780
rect -1482 -826 -1478 -780
rect -1458 -826 -1454 -780
rect -1434 -826 -1430 -780
rect -1410 -826 -1406 -780
rect -1386 -826 -1382 -780
rect -1362 -826 -1358 -780
rect -1338 -826 -1334 -780
rect -1314 -826 -1310 -780
rect -1290 -826 -1286 -780
rect -1266 -826 -1262 -780
rect -1242 -825 -1238 -780
rect -1253 -826 -1219 -825
rect -2393 -828 -1219 -826
rect -2371 -850 -2366 -828
rect -2348 -850 -2343 -828
rect -2325 -834 -2317 -828
rect -2325 -850 -2320 -834
rect -2317 -836 -2309 -834
rect -2309 -848 -2301 -836
rect -2080 -837 -2071 -828
rect -2068 -838 -2059 -837
rect -2068 -845 -2038 -838
rect -2317 -850 -2309 -848
rect -2068 -850 -2059 -845
rect -2000 -846 -1992 -828
rect -1846 -836 -1794 -828
rect -1671 -834 -1663 -828
rect -1663 -836 -1655 -834
rect -1852 -845 -1804 -838
rect -2011 -848 -1983 -846
rect -2025 -849 -1983 -848
rect -2025 -850 -1975 -849
rect -1846 -850 -1804 -847
rect -1655 -848 -1647 -836
rect -1663 -850 -1655 -848
rect -1642 -850 -1637 -828
rect -1619 -850 -1614 -828
rect -1530 -850 -1526 -828
rect -1506 -850 -1502 -828
rect -1482 -850 -1478 -828
rect -1458 -850 -1454 -828
rect -1434 -850 -1430 -828
rect -1410 -850 -1406 -828
rect -1386 -850 -1382 -828
rect -1362 -850 -1358 -828
rect -1338 -850 -1334 -828
rect -1314 -850 -1310 -828
rect -1290 -850 -1286 -828
rect -1266 -850 -1262 -828
rect -1253 -835 -1248 -828
rect -1242 -835 -1238 -828
rect -1243 -849 -1238 -835
rect -1218 -850 -1214 -780
rect -1194 -850 -1190 -780
rect -1187 -781 -1173 -780
rect -1170 -781 -1163 -757
rect -1170 -829 -1163 -805
rect -1170 -850 -1166 -829
rect -1146 -850 -1142 -756
rect -1122 -850 -1118 -756
rect -1098 -850 -1094 -756
rect -1074 -850 -1070 -756
rect -1050 -850 -1046 -756
rect -1026 -850 -1022 -756
rect -1002 -850 -998 -756
rect -978 -850 -974 -756
rect -954 -850 -950 -756
rect -930 -850 -926 -756
rect -906 -850 -902 -756
rect -882 -850 -878 -756
rect -858 -850 -854 -756
rect -834 -850 -830 -756
rect -810 -850 -806 -756
rect -786 -850 -782 -756
rect -762 -850 -758 -756
rect -738 -850 -734 -756
rect -714 -850 -710 -756
rect -690 -778 -683 -757
rect -666 -778 -662 -756
rect -642 -778 -638 -756
rect -594 -778 -590 -756
rect -570 -778 -566 -756
rect -546 -778 -542 -756
rect -522 -778 -518 -756
rect -498 -778 -494 -756
rect -474 -778 -470 -756
rect -450 -778 -446 -756
rect -426 -778 -422 -756
rect -402 -778 -398 -756
rect -378 -778 -374 -756
rect -354 -778 -350 -756
rect -306 -778 -302 -756
rect -282 -778 -278 -756
rect -258 -778 -254 -756
rect -234 -778 -230 -756
rect -210 -778 -206 -756
rect -186 -778 -182 -756
rect -162 -778 -158 -756
rect -138 -778 -134 -756
rect -114 -778 -110 -756
rect -90 -778 -86 -756
rect -66 -778 -62 -756
rect -42 -778 -38 -756
rect -18 -777 -14 -756
rect -29 -778 5 -777
rect -707 -780 5 -778
rect -707 -781 -693 -780
rect -690 -781 -683 -780
rect -690 -850 -686 -781
rect -666 -850 -662 -780
rect -642 -850 -638 -780
rect -594 -781 -590 -780
rect -629 -804 -597 -801
rect -629 -811 -624 -804
rect -611 -805 -597 -804
rect -594 -805 -587 -781
rect -619 -825 -614 -811
rect -618 -850 -614 -825
rect -570 -850 -566 -780
rect -546 -850 -542 -780
rect -522 -850 -518 -780
rect -498 -850 -494 -780
rect -474 -850 -470 -780
rect -450 -850 -446 -780
rect -426 -850 -422 -780
rect -402 -850 -398 -780
rect -378 -850 -374 -780
rect -354 -850 -350 -780
rect -306 -805 -302 -780
rect -341 -828 -309 -825
rect -341 -835 -336 -828
rect -323 -829 -309 -828
rect -306 -829 -299 -805
rect -331 -849 -326 -835
rect -330 -850 -326 -849
rect -282 -850 -278 -780
rect -258 -850 -254 -780
rect -234 -850 -230 -780
rect -210 -850 -206 -780
rect -186 -850 -182 -780
rect -162 -850 -158 -780
rect -138 -850 -134 -780
rect -114 -850 -110 -780
rect -90 -850 -86 -780
rect -66 -850 -62 -780
rect -42 -850 -38 -780
rect -29 -787 -24 -780
rect -18 -787 -14 -780
rect -19 -801 -14 -787
rect 6 -850 10 -756
rect 30 -850 34 -756
rect 54 -850 58 -756
rect 78 -850 82 -756
rect 102 -850 106 -756
rect 126 -850 130 -756
rect 150 -850 154 -756
rect 174 -850 178 -756
rect 198 -850 202 -756
rect 222 -850 226 -756
rect 235 -763 240 -756
rect 246 -763 250 -756
rect 245 -777 250 -763
rect 235 -778 269 -777
rect 270 -778 274 -684
rect 294 -778 298 -684
rect 318 -778 322 -684
rect 342 -778 346 -684
rect 366 -778 370 -684
rect 390 -778 394 -684
rect 414 -778 418 -684
rect 438 -778 442 -684
rect 462 -778 466 -684
rect 486 -778 490 -684
rect 510 -778 514 -684
rect 534 -778 538 -684
rect 558 -778 562 -684
rect 582 -778 586 -684
rect 606 -778 610 -684
rect 630 -778 634 -684
rect 654 -778 658 -684
rect 678 -778 682 -684
rect 702 -778 706 -684
rect 709 -685 723 -684
rect 726 -709 733 -661
rect 726 -778 730 -709
rect 750 -778 754 -660
rect 774 -778 778 -660
rect 798 -778 802 -660
rect 822 -778 826 -660
rect 846 -777 850 -660
rect 859 -691 864 -681
rect 870 -691 874 -660
rect 883 -667 888 -660
rect 894 -667 898 -660
rect 893 -681 898 -667
rect 869 -705 874 -691
rect 835 -778 869 -777
rect 235 -780 869 -778
rect 235 -787 240 -780
rect 245 -801 250 -787
rect 246 -850 250 -801
rect 270 -829 274 -780
rect -2393 -852 267 -850
rect -2371 -874 -2366 -852
rect -2348 -874 -2343 -852
rect -2325 -862 -2317 -852
rect -2068 -853 -2038 -852
rect -2068 -855 -2059 -853
rect -2013 -854 -1983 -852
rect -1846 -853 -1804 -852
rect -2000 -855 -1983 -854
rect -1862 -855 -1798 -854
rect -2076 -862 -2068 -855
rect -2061 -862 -2045 -860
rect -2038 -862 -2001 -855
rect -2325 -874 -2320 -862
rect -2317 -864 -2309 -862
rect -2309 -874 -2301 -864
rect -2068 -865 -2045 -862
rect -2015 -863 -2001 -862
rect -2068 -872 -2038 -865
rect -2068 -874 -2045 -872
rect -2000 -874 -1992 -855
rect -1985 -857 -1796 -855
rect -1985 -862 -1852 -857
rect -1846 -862 -1796 -857
rect -1671 -862 -1663 -852
rect -1846 -863 -1798 -862
rect -1663 -864 -1655 -862
rect -1852 -872 -1804 -865
rect -1976 -874 -1940 -873
rect -1655 -874 -1647 -864
rect -1642 -874 -1637 -852
rect -1619 -874 -1614 -852
rect -1530 -874 -1526 -852
rect -1506 -874 -1502 -852
rect -1482 -874 -1478 -852
rect -1458 -874 -1454 -852
rect -1434 -874 -1430 -852
rect -1410 -874 -1406 -852
rect -1386 -874 -1382 -852
rect -1362 -874 -1358 -852
rect -1338 -874 -1334 -852
rect -1314 -874 -1310 -852
rect -1290 -874 -1286 -852
rect -1266 -874 -1262 -852
rect -1253 -874 -1219 -873
rect -1218 -874 -1214 -852
rect -1194 -873 -1190 -852
rect -1205 -874 -1171 -873
rect -2393 -876 -1171 -874
rect -2371 -946 -2366 -876
rect -2348 -946 -2343 -876
rect -2325 -878 -2320 -876
rect -2317 -878 -2309 -876
rect -2325 -890 -2317 -878
rect -2068 -882 -2059 -876
rect -2076 -889 -2071 -882
rect -2068 -890 -2059 -889
rect -2325 -910 -2320 -890
rect -2317 -892 -2309 -890
rect -2325 -918 -2317 -910
rect -2060 -916 -2030 -913
rect -2325 -938 -2320 -918
rect -2317 -926 -2309 -918
rect -2060 -929 -2038 -918
rect -2033 -925 -2030 -916
rect -2028 -920 -2027 -916
rect -2068 -934 -2038 -931
rect -2325 -946 -2317 -938
rect -2000 -943 -1992 -876
rect -1846 -880 -1804 -876
rect -1663 -878 -1655 -876
rect -1846 -890 -1794 -881
rect -1671 -890 -1663 -878
rect -1663 -892 -1655 -890
rect -1912 -901 -1884 -899
rect -1852 -907 -1804 -903
rect -1844 -916 -1796 -913
rect -1671 -918 -1663 -910
rect -1844 -929 -1804 -918
rect -1663 -926 -1655 -918
rect -1852 -934 -1680 -930
rect -2119 -946 -2069 -944
rect -2007 -946 -1977 -943
rect -1926 -946 -1892 -943
rect -1671 -946 -1663 -938
rect -1642 -946 -1637 -876
rect -1619 -946 -1614 -876
rect -1530 -946 -1526 -876
rect -1506 -946 -1502 -876
rect -1482 -946 -1478 -876
rect -1458 -946 -1454 -876
rect -1434 -946 -1430 -876
rect -1410 -946 -1406 -876
rect -1386 -946 -1382 -876
rect -1362 -946 -1358 -876
rect -1338 -946 -1334 -876
rect -1314 -946 -1310 -876
rect -1290 -946 -1286 -876
rect -1266 -946 -1262 -876
rect -1253 -883 -1248 -876
rect -1243 -897 -1238 -883
rect -1242 -946 -1238 -897
rect -1218 -901 -1214 -876
rect -1205 -883 -1200 -876
rect -1194 -883 -1190 -876
rect -1195 -897 -1190 -883
rect -1218 -925 -1211 -901
rect -1205 -931 -1200 -921
rect -1195 -945 -1190 -931
rect -1194 -946 -1190 -945
rect -1170 -946 -1166 -852
rect -1146 -946 -1142 -852
rect -1122 -946 -1118 -852
rect -1098 -946 -1094 -852
rect -1074 -946 -1070 -852
rect -1050 -946 -1046 -852
rect -1026 -946 -1022 -852
rect -1002 -946 -998 -852
rect -978 -946 -974 -852
rect -954 -946 -950 -852
rect -930 -946 -926 -852
rect -906 -946 -902 -852
rect -882 -946 -878 -852
rect -858 -946 -854 -852
rect -834 -946 -830 -852
rect -810 -946 -806 -852
rect -786 -946 -782 -852
rect -762 -946 -758 -852
rect -738 -946 -734 -852
rect -714 -946 -710 -852
rect -690 -946 -686 -852
rect -666 -946 -662 -852
rect -642 -946 -638 -852
rect -618 -946 -614 -852
rect -594 -898 -587 -877
rect -570 -898 -566 -852
rect -546 -898 -542 -852
rect -522 -898 -518 -852
rect -498 -898 -494 -852
rect -474 -898 -470 -852
rect -450 -898 -446 -852
rect -426 -898 -422 -852
rect -402 -897 -398 -852
rect -413 -898 -379 -897
rect -611 -900 -379 -898
rect -611 -901 -597 -900
rect -594 -901 -587 -900
rect -594 -946 -590 -901
rect -570 -946 -566 -900
rect -546 -946 -542 -900
rect -522 -946 -518 -900
rect -498 -946 -494 -900
rect -474 -946 -470 -900
rect -450 -946 -446 -900
rect -426 -946 -422 -900
rect -413 -907 -408 -900
rect -402 -907 -398 -900
rect -403 -921 -398 -907
rect -413 -946 -379 -945
rect -2393 -948 -379 -946
rect -2371 -970 -2366 -948
rect -2348 -970 -2343 -948
rect -2325 -952 -2317 -948
rect -2325 -968 -2320 -952
rect -2317 -954 -2309 -952
rect -2309 -966 -2301 -954
rect -2000 -962 -1992 -948
rect -1671 -952 -1663 -948
rect -1663 -954 -1655 -952
rect -1844 -956 -1806 -954
rect -1854 -962 -1806 -958
rect -2068 -965 -2060 -962
rect -2030 -965 -1958 -962
rect -1942 -965 -1806 -962
rect -2317 -968 -2309 -966
rect -2000 -968 -1992 -965
rect -1655 -966 -1647 -954
rect -2325 -970 -2317 -968
rect -2033 -970 -1992 -968
rect -1844 -969 -1806 -967
rect -1663 -968 -1655 -966
rect -1864 -970 -1796 -969
rect -1671 -970 -1663 -968
rect -1642 -970 -1637 -948
rect -1619 -970 -1614 -948
rect -1530 -970 -1526 -948
rect -1506 -970 -1502 -948
rect -1482 -970 -1478 -948
rect -1458 -970 -1454 -948
rect -1434 -970 -1430 -948
rect -1410 -970 -1406 -948
rect -1386 -970 -1382 -948
rect -1362 -970 -1358 -948
rect -1338 -970 -1334 -948
rect -1314 -970 -1310 -948
rect -1290 -970 -1286 -948
rect -1266 -970 -1262 -948
rect -1242 -970 -1238 -948
rect -1218 -970 -1211 -949
rect -1194 -970 -1190 -948
rect -1170 -949 -1166 -948
rect -2393 -972 -1173 -970
rect -2371 -994 -2366 -972
rect -2348 -994 -2343 -972
rect -2325 -980 -2317 -972
rect -2060 -975 -2030 -972
rect -2000 -975 -1992 -972
rect -1972 -974 -1958 -972
rect -1904 -975 -1798 -972
rect -2078 -979 -2020 -975
rect -2023 -980 -2020 -979
rect -2000 -977 -1798 -975
rect -2000 -979 -1854 -977
rect -1844 -979 -1798 -977
rect -2325 -994 -2320 -980
rect -2317 -982 -2309 -980
rect -2020 -982 -2004 -980
rect -2000 -982 -1992 -979
rect -1671 -980 -1663 -972
rect -2309 -994 -2301 -982
rect -2020 -984 -1992 -982
rect -1844 -983 -1806 -981
rect -1663 -982 -1655 -980
rect -2023 -989 -1992 -984
rect -1854 -989 -1806 -985
rect -2068 -992 -2060 -989
rect -2030 -992 -1806 -989
rect -2074 -994 -2060 -992
rect -2020 -994 -2004 -992
rect -2000 -994 -1992 -992
rect -1655 -994 -1647 -982
rect -1642 -994 -1637 -972
rect -1619 -994 -1614 -972
rect -1530 -994 -1526 -972
rect -1506 -994 -1502 -972
rect -1482 -994 -1478 -972
rect -1458 -994 -1454 -972
rect -1434 -994 -1430 -972
rect -1410 -994 -1406 -972
rect -1386 -994 -1382 -972
rect -1362 -994 -1358 -972
rect -1338 -994 -1334 -972
rect -1314 -994 -1310 -972
rect -1290 -994 -1286 -972
rect -1266 -994 -1262 -972
rect -1242 -994 -1238 -972
rect -1235 -973 -1221 -972
rect -1218 -973 -1211 -972
rect -1218 -994 -1214 -973
rect -1194 -994 -1190 -972
rect -1187 -973 -1173 -972
rect -1170 -973 -1163 -949
rect -1146 -994 -1142 -948
rect -1122 -994 -1118 -948
rect -1098 -994 -1094 -948
rect -1074 -994 -1070 -948
rect -1050 -994 -1046 -948
rect -1026 -994 -1022 -948
rect -1002 -994 -998 -948
rect -978 -994 -974 -948
rect -954 -994 -950 -948
rect -930 -994 -926 -948
rect -906 -994 -902 -948
rect -882 -994 -878 -948
rect -858 -994 -854 -948
rect -834 -994 -830 -948
rect -821 -979 -816 -969
rect -810 -979 -806 -948
rect -811 -993 -806 -979
rect -786 -994 -782 -948
rect -762 -994 -758 -948
rect -738 -994 -734 -948
rect -714 -994 -710 -948
rect -690 -994 -686 -948
rect -666 -994 -662 -948
rect -642 -994 -638 -948
rect -618 -994 -614 -948
rect -594 -994 -590 -948
rect -570 -994 -566 -948
rect -546 -994 -542 -948
rect -522 -994 -518 -948
rect -498 -994 -494 -948
rect -474 -994 -470 -948
rect -450 -994 -446 -948
rect -426 -994 -422 -948
rect -413 -955 -408 -948
rect -403 -969 -398 -955
rect -378 -958 -374 -852
rect -412 -982 -408 -972
rect -389 -979 -384 -969
rect -402 -994 -398 -982
rect -379 -993 -371 -979
rect -2393 -996 -2060 -994
rect -2050 -996 -381 -994
rect -2371 -1042 -2366 -996
rect -2348 -1042 -2343 -996
rect -2325 -1008 -2317 -996
rect -2109 -999 -2108 -996
rect -2117 -1006 -2108 -999
rect -2325 -1028 -2320 -1008
rect -2317 -1010 -2309 -1008
rect -2109 -1010 -2108 -1006
rect -2060 -1006 -2030 -999
rect -2060 -1010 -2034 -1006
rect -2325 -1036 -2317 -1028
rect -2101 -1033 -2071 -1030
rect -2325 -1042 -2320 -1036
rect -2317 -1042 -2309 -1036
rect -2000 -1038 -1992 -996
rect -1844 -997 -1806 -996
rect -1844 -1006 -1798 -999
rect -1671 -1008 -1663 -996
rect -1844 -1010 -1806 -1008
rect -1663 -1010 -1655 -1008
rect -1854 -1024 -1680 -1020
rect -1846 -1033 -1798 -1030
rect -2079 -1039 -2043 -1038
rect -2007 -1039 -1991 -1038
rect -2079 -1040 -2071 -1039
rect -2079 -1042 -2029 -1040
rect -2011 -1042 -1991 -1039
rect -1846 -1041 -1806 -1035
rect -1671 -1036 -1663 -1028
rect -1864 -1042 -1796 -1041
rect -1663 -1042 -1655 -1036
rect -1642 -1042 -1637 -996
rect -1619 -1042 -1614 -996
rect -1530 -1042 -1526 -996
rect -1506 -1042 -1502 -996
rect -1482 -1042 -1478 -996
rect -1458 -1042 -1454 -996
rect -1434 -1042 -1430 -996
rect -1410 -1042 -1406 -996
rect -1386 -1042 -1382 -996
rect -1362 -1042 -1358 -996
rect -1338 -1042 -1334 -996
rect -1314 -1042 -1310 -996
rect -1290 -1042 -1286 -996
rect -1266 -1041 -1262 -996
rect -1277 -1042 -1243 -1041
rect -2393 -1044 -1243 -1042
rect -2371 -1114 -2366 -1044
rect -2348 -1114 -2343 -1044
rect -2325 -1056 -2320 -1044
rect -2079 -1046 -2071 -1044
rect -2072 -1048 -2071 -1046
rect -2109 -1053 -2101 -1048
rect -2101 -1055 -2079 -1053
rect -2069 -1055 -2068 -1048
rect -2325 -1064 -2317 -1056
rect -2079 -1060 -2071 -1055
rect -2325 -1114 -2320 -1064
rect -2317 -1072 -2309 -1064
rect -2074 -1069 -2071 -1060
rect -2069 -1064 -2068 -1060
rect -2109 -1078 -2079 -1075
rect -2309 -1112 -2301 -1102
rect -2317 -1114 -2309 -1112
rect -2000 -1114 -1992 -1044
rect -1846 -1046 -1806 -1044
rect -1854 -1051 -1806 -1047
rect -1854 -1053 -1846 -1051
rect -1846 -1055 -1806 -1053
rect -1806 -1057 -1798 -1055
rect -1846 -1060 -1798 -1057
rect -1846 -1073 -1806 -1062
rect -1671 -1064 -1663 -1056
rect -1663 -1072 -1655 -1064
rect -1854 -1078 -1680 -1074
rect -1655 -1112 -1647 -1102
rect -1663 -1114 -1655 -1112
rect -1642 -1114 -1637 -1044
rect -1619 -1114 -1614 -1044
rect -1530 -1114 -1526 -1044
rect -1506 -1114 -1502 -1044
rect -1482 -1114 -1478 -1044
rect -1458 -1114 -1454 -1044
rect -1434 -1114 -1430 -1044
rect -1410 -1114 -1406 -1044
rect -1386 -1114 -1382 -1044
rect -1362 -1114 -1358 -1044
rect -1338 -1114 -1334 -1044
rect -1314 -1114 -1310 -1044
rect -1290 -1114 -1286 -1044
rect -1277 -1051 -1272 -1044
rect -1266 -1051 -1262 -1044
rect -1267 -1065 -1262 -1051
rect -1277 -1066 -1243 -1065
rect -1242 -1066 -1238 -996
rect -1218 -1066 -1214 -996
rect -1194 -1066 -1190 -996
rect -1170 -1018 -1163 -997
rect -1146 -1018 -1142 -996
rect -1122 -1018 -1118 -996
rect -1098 -1018 -1094 -996
rect -1074 -1018 -1070 -996
rect -1050 -1018 -1046 -996
rect -1026 -1018 -1022 -996
rect -1002 -1018 -998 -996
rect -978 -1018 -974 -996
rect -954 -1018 -950 -996
rect -930 -1018 -926 -996
rect -906 -1018 -902 -996
rect -882 -1018 -878 -996
rect -858 -1018 -854 -996
rect -834 -1018 -830 -996
rect -821 -1018 -787 -1017
rect -786 -1018 -782 -996
rect -762 -1018 -758 -996
rect -738 -1018 -734 -996
rect -714 -1018 -710 -996
rect -690 -1018 -686 -996
rect -666 -1018 -662 -996
rect -642 -1018 -638 -996
rect -618 -1018 -614 -996
rect -594 -1018 -590 -996
rect -570 -1018 -566 -996
rect -546 -1018 -542 -996
rect -522 -1018 -518 -996
rect -498 -1018 -494 -996
rect -474 -1018 -470 -996
rect -450 -1018 -446 -996
rect -426 -1018 -422 -996
rect -402 -1018 -398 -996
rect -395 -997 -381 -996
rect -354 -1018 -350 -852
rect -330 -1018 -326 -852
rect -306 -922 -299 -901
rect -282 -922 -278 -852
rect -258 -922 -254 -852
rect -234 -922 -230 -852
rect -210 -922 -206 -852
rect -186 -922 -182 -852
rect -162 -922 -158 -852
rect -138 -922 -134 -852
rect -114 -922 -110 -852
rect -90 -922 -86 -852
rect -66 -922 -62 -852
rect -42 -922 -38 -852
rect 6 -853 10 -852
rect -29 -876 3 -873
rect -29 -883 -24 -876
rect -11 -877 3 -876
rect 6 -877 13 -853
rect -19 -897 -14 -883
rect -18 -922 -14 -897
rect 30 -922 34 -852
rect 54 -922 58 -852
rect 78 -922 82 -852
rect 102 -922 106 -852
rect 126 -922 130 -852
rect 150 -922 154 -852
rect 174 -922 178 -852
rect 198 -922 202 -852
rect 222 -922 226 -852
rect 246 -922 250 -852
rect 253 -853 267 -852
rect 270 -874 277 -829
rect 294 -874 298 -780
rect 318 -874 322 -780
rect 342 -874 346 -780
rect 366 -874 370 -780
rect 390 -874 394 -780
rect 414 -874 418 -780
rect 438 -874 442 -780
rect 462 -874 466 -780
rect 486 -874 490 -780
rect 510 -874 514 -780
rect 534 -874 538 -780
rect 558 -874 562 -780
rect 582 -874 586 -780
rect 595 -859 600 -849
rect 606 -859 610 -780
rect 605 -873 610 -859
rect 630 -874 634 -780
rect 654 -874 658 -780
rect 678 -874 682 -780
rect 702 -874 706 -780
rect 726 -874 730 -780
rect 750 -874 754 -780
rect 774 -873 778 -780
rect 787 -835 792 -825
rect 798 -835 802 -780
rect 811 -811 816 -801
rect 822 -811 826 -780
rect 835 -787 840 -780
rect 846 -787 850 -780
rect 845 -801 850 -787
rect 821 -825 826 -811
rect 797 -849 802 -835
rect 763 -874 797 -873
rect 253 -876 797 -874
rect 253 -877 267 -876
rect 270 -877 277 -876
rect 270 -922 274 -877
rect 294 -922 298 -876
rect 318 -922 322 -876
rect 342 -922 346 -876
rect 366 -922 370 -876
rect 390 -922 394 -876
rect 414 -922 418 -876
rect 438 -922 442 -876
rect 462 -922 466 -876
rect 486 -922 490 -876
rect 510 -922 514 -876
rect 534 -922 538 -876
rect 558 -922 562 -876
rect 582 -922 586 -876
rect 595 -898 629 -897
rect 630 -898 634 -876
rect 654 -898 658 -876
rect 678 -898 682 -876
rect 702 -898 706 -876
rect 726 -898 730 -876
rect 750 -897 754 -876
rect 763 -883 768 -876
rect 774 -883 778 -876
rect 773 -897 778 -883
rect 739 -898 773 -897
rect 595 -900 773 -898
rect 595 -907 600 -900
rect 605 -921 610 -907
rect 606 -922 610 -921
rect 630 -922 634 -900
rect 654 -922 658 -900
rect 678 -922 682 -900
rect 702 -922 706 -900
rect 726 -921 730 -900
rect 739 -907 744 -900
rect 750 -907 754 -900
rect 749 -921 754 -907
rect 715 -922 749 -921
rect -323 -924 749 -922
rect -323 -925 -309 -924
rect -306 -925 -299 -924
rect -306 -1018 -302 -925
rect -282 -1018 -278 -924
rect -258 -1018 -254 -924
rect -234 -1018 -230 -924
rect -210 -1018 -206 -924
rect -186 -1018 -182 -924
rect -162 -1018 -158 -924
rect -138 -1018 -134 -924
rect -125 -1003 -120 -993
rect -114 -1003 -110 -924
rect -115 -1017 -110 -1003
rect -90 -1018 -86 -924
rect -66 -1018 -62 -924
rect -42 -1018 -38 -924
rect -18 -1018 -14 -924
rect 6 -970 13 -949
rect 30 -970 34 -924
rect 54 -970 58 -924
rect 78 -970 82 -924
rect 102 -970 106 -924
rect 126 -970 130 -924
rect 150 -970 154 -924
rect 174 -970 178 -924
rect 198 -970 202 -924
rect 222 -970 226 -924
rect 246 -970 250 -924
rect 270 -970 274 -924
rect 294 -970 298 -924
rect 318 -970 322 -924
rect 342 -970 346 -924
rect 366 -970 370 -924
rect 390 -970 394 -924
rect 414 -970 418 -924
rect 438 -970 442 -924
rect 462 -970 466 -924
rect 486 -970 490 -924
rect 510 -970 514 -924
rect 534 -970 538 -924
rect 558 -970 562 -924
rect 582 -970 586 -924
rect 606 -970 610 -924
rect 630 -925 634 -924
rect 630 -949 637 -925
rect 654 -970 658 -924
rect 678 -970 682 -924
rect 702 -969 706 -924
rect 715 -931 720 -924
rect 726 -931 730 -924
rect 725 -945 730 -931
rect 691 -970 725 -969
rect -11 -972 725 -970
rect -11 -973 3 -972
rect 6 -973 13 -972
rect 6 -1018 10 -973
rect 30 -1018 34 -972
rect 54 -1018 58 -972
rect 78 -1018 82 -972
rect 102 -1017 106 -972
rect 91 -1018 125 -1017
rect -1187 -1020 125 -1018
rect -1187 -1021 -1173 -1020
rect -1170 -1021 -1163 -1020
rect -1170 -1066 -1166 -1021
rect -1146 -1066 -1142 -1020
rect -1122 -1066 -1118 -1020
rect -1098 -1066 -1094 -1020
rect -1074 -1066 -1070 -1020
rect -1050 -1066 -1046 -1020
rect -1026 -1066 -1022 -1020
rect -1002 -1066 -998 -1020
rect -978 -1066 -974 -1020
rect -954 -1066 -950 -1020
rect -930 -1066 -926 -1020
rect -906 -1066 -902 -1020
rect -882 -1066 -878 -1020
rect -858 -1066 -854 -1020
rect -834 -1066 -830 -1020
rect -821 -1027 -816 -1020
rect -811 -1041 -806 -1027
rect -810 -1066 -806 -1041
rect -786 -1045 -782 -1020
rect -1277 -1068 -789 -1066
rect -1277 -1075 -1272 -1068
rect -1267 -1089 -1262 -1075
rect -1266 -1114 -1262 -1089
rect -1242 -1114 -1238 -1068
rect -1218 -1114 -1214 -1068
rect -1194 -1114 -1190 -1068
rect -1170 -1114 -1166 -1068
rect -1146 -1114 -1142 -1068
rect -1122 -1114 -1118 -1068
rect -1098 -1114 -1094 -1068
rect -1074 -1114 -1070 -1068
rect -1050 -1114 -1046 -1068
rect -1026 -1114 -1022 -1068
rect -1002 -1114 -998 -1068
rect -978 -1114 -974 -1068
rect -954 -1114 -950 -1068
rect -930 -1114 -926 -1068
rect -906 -1114 -902 -1068
rect -882 -1114 -878 -1068
rect -858 -1114 -854 -1068
rect -834 -1114 -830 -1068
rect -810 -1114 -806 -1068
rect -803 -1069 -789 -1068
rect -786 -1069 -779 -1045
rect -786 -1114 -779 -1093
rect -762 -1114 -758 -1020
rect -738 -1114 -734 -1020
rect -714 -1114 -710 -1020
rect -690 -1114 -686 -1020
rect -666 -1114 -662 -1020
rect -642 -1114 -638 -1020
rect -618 -1114 -614 -1020
rect -594 -1114 -590 -1020
rect -570 -1114 -566 -1020
rect -546 -1114 -542 -1020
rect -522 -1114 -518 -1020
rect -498 -1114 -494 -1020
rect -474 -1114 -470 -1020
rect -450 -1114 -446 -1020
rect -426 -1114 -422 -1020
rect -402 -1114 -398 -1020
rect -389 -1044 -360 -1041
rect -354 -1044 -350 -1020
rect -389 -1045 -381 -1044
rect -365 -1055 -357 -1051
rect -371 -1065 -365 -1055
rect -354 -1066 -347 -1045
rect -330 -1066 -326 -1020
rect -306 -1066 -302 -1020
rect -282 -1066 -278 -1020
rect -258 -1066 -254 -1020
rect -234 -1066 -230 -1020
rect -210 -1066 -206 -1020
rect -186 -1066 -182 -1020
rect -162 -1066 -158 -1020
rect -138 -1066 -134 -1020
rect -90 -1066 -86 -1020
rect -66 -1066 -62 -1020
rect -42 -1066 -38 -1020
rect -18 -1066 -14 -1020
rect 6 -1066 10 -1020
rect 30 -1066 34 -1020
rect 54 -1066 58 -1020
rect 78 -1066 82 -1020
rect 91 -1027 96 -1020
rect 102 -1027 106 -1020
rect 101 -1041 106 -1027
rect 126 -1066 130 -972
rect 150 -1066 154 -972
rect 174 -1066 178 -972
rect 198 -1066 202 -972
rect 222 -1066 226 -972
rect 246 -1066 250 -972
rect 270 -1066 274 -972
rect 294 -1066 298 -972
rect 318 -1066 322 -972
rect 342 -1066 346 -972
rect 366 -1066 370 -972
rect 390 -1066 394 -972
rect 414 -1066 418 -972
rect 438 -1066 442 -972
rect 462 -1066 466 -972
rect 486 -1066 490 -972
rect 510 -1066 514 -972
rect 534 -1066 538 -972
rect 558 -1066 562 -972
rect 582 -1066 586 -972
rect 606 -1066 610 -972
rect 630 -997 637 -973
rect 630 -1066 634 -997
rect 654 -1065 658 -972
rect 667 -1051 672 -1041
rect 678 -1051 682 -972
rect 691 -979 696 -972
rect 702 -979 706 -972
rect 701 -993 706 -979
rect 677 -1065 682 -1051
rect 643 -1066 677 -1065
rect -371 -1068 677 -1066
rect -378 -1114 -374 -1068
rect -371 -1069 -357 -1068
rect -354 -1069 -347 -1068
rect -330 -1114 -326 -1068
rect -306 -1114 -302 -1068
rect -282 -1114 -278 -1068
rect -258 -1114 -254 -1068
rect -234 -1114 -230 -1068
rect -210 -1114 -206 -1068
rect -186 -1114 -182 -1068
rect -162 -1114 -158 -1068
rect -138 -1114 -134 -1068
rect -90 -1069 -86 -1068
rect -125 -1092 -93 -1089
rect -125 -1099 -120 -1092
rect -107 -1093 -93 -1092
rect -90 -1093 -83 -1069
rect -115 -1113 -110 -1099
rect -114 -1114 -110 -1113
rect -66 -1114 -62 -1068
rect -42 -1114 -38 -1068
rect -18 -1114 -14 -1068
rect 6 -1114 10 -1068
rect 30 -1114 34 -1068
rect 54 -1114 58 -1068
rect 78 -1114 82 -1068
rect 126 -1093 130 -1068
rect 91 -1114 123 -1113
rect -2393 -1116 123 -1114
rect -2371 -1210 -2366 -1116
rect -2348 -1210 -2343 -1116
rect -2325 -1178 -2320 -1116
rect -2317 -1118 -2309 -1116
rect -2013 -1118 -1992 -1116
rect -1663 -1118 -1655 -1116
rect -2000 -1119 -1983 -1118
rect -2026 -1128 -2021 -1124
rect -2062 -1129 -2061 -1128
rect -2309 -1140 -2301 -1130
rect -2091 -1136 -2061 -1129
rect -2317 -1146 -2309 -1140
rect -2132 -1145 -2131 -1143
rect -2101 -1145 -2092 -1143
rect -2091 -1144 -2071 -1138
rect -2062 -1140 -2045 -1136
rect -2036 -1140 -2031 -1138
rect -2292 -1154 -2071 -1145
rect -2107 -1159 -2104 -1155
rect -2325 -1186 -2317 -1178
rect -2325 -1206 -2320 -1186
rect -2317 -1194 -2309 -1186
rect -2325 -1210 -2317 -1206
rect -2000 -1210 -1992 -1119
rect -1980 -1136 -1932 -1129
rect -1655 -1140 -1647 -1130
rect -1846 -1154 -1680 -1145
rect -1663 -1146 -1655 -1140
rect -1671 -1186 -1663 -1178
rect -1663 -1194 -1655 -1186
rect -1926 -1210 -1892 -1207
rect -1671 -1210 -1663 -1206
rect -1642 -1210 -1637 -1116
rect -1619 -1210 -1614 -1116
rect -1530 -1210 -1526 -1116
rect -1506 -1210 -1502 -1116
rect -1482 -1210 -1478 -1116
rect -1458 -1210 -1454 -1116
rect -1434 -1210 -1430 -1116
rect -1410 -1210 -1406 -1116
rect -1386 -1210 -1382 -1116
rect -1362 -1210 -1358 -1116
rect -1338 -1210 -1334 -1116
rect -1314 -1210 -1310 -1116
rect -1290 -1210 -1286 -1116
rect -1266 -1210 -1262 -1116
rect -1242 -1117 -1238 -1116
rect -1242 -1162 -1235 -1117
rect -1218 -1162 -1214 -1116
rect -1194 -1162 -1190 -1116
rect -1170 -1162 -1166 -1116
rect -1146 -1162 -1142 -1116
rect -1122 -1162 -1118 -1116
rect -1098 -1162 -1094 -1116
rect -1074 -1162 -1070 -1116
rect -1050 -1162 -1046 -1116
rect -1026 -1162 -1022 -1116
rect -1002 -1162 -998 -1116
rect -978 -1162 -974 -1116
rect -954 -1162 -950 -1116
rect -930 -1162 -926 -1116
rect -906 -1162 -902 -1116
rect -882 -1162 -878 -1116
rect -858 -1162 -854 -1116
rect -834 -1162 -830 -1116
rect -810 -1162 -806 -1116
rect -803 -1117 -789 -1116
rect -786 -1117 -779 -1116
rect -786 -1162 -782 -1117
rect -762 -1162 -758 -1116
rect -738 -1162 -734 -1116
rect -714 -1162 -710 -1116
rect -690 -1162 -686 -1116
rect -666 -1162 -662 -1116
rect -642 -1162 -638 -1116
rect -618 -1162 -614 -1116
rect -594 -1162 -590 -1116
rect -570 -1162 -566 -1116
rect -546 -1161 -542 -1116
rect -557 -1162 -523 -1161
rect -1259 -1164 -523 -1162
rect -1259 -1165 -1245 -1164
rect -1242 -1165 -1235 -1164
rect -1242 -1210 -1238 -1165
rect -1218 -1210 -1214 -1164
rect -1194 -1210 -1190 -1164
rect -1170 -1210 -1166 -1164
rect -1146 -1210 -1142 -1164
rect -1122 -1210 -1118 -1164
rect -1098 -1210 -1094 -1164
rect -1074 -1210 -1070 -1164
rect -1050 -1210 -1046 -1164
rect -1026 -1210 -1022 -1164
rect -1002 -1210 -998 -1164
rect -978 -1210 -974 -1164
rect -954 -1210 -950 -1164
rect -930 -1210 -926 -1164
rect -906 -1210 -902 -1164
rect -882 -1210 -878 -1164
rect -858 -1210 -854 -1164
rect -834 -1210 -830 -1164
rect -810 -1210 -806 -1164
rect -786 -1210 -782 -1164
rect -762 -1210 -758 -1164
rect -738 -1210 -734 -1164
rect -714 -1210 -710 -1164
rect -690 -1210 -686 -1164
rect -666 -1210 -662 -1164
rect -642 -1210 -638 -1164
rect -618 -1210 -614 -1164
rect -594 -1210 -590 -1164
rect -570 -1210 -566 -1164
rect -557 -1171 -552 -1164
rect -546 -1171 -542 -1164
rect -547 -1185 -542 -1171
rect -557 -1195 -552 -1185
rect -547 -1209 -542 -1195
rect -546 -1210 -542 -1209
rect -522 -1210 -518 -1116
rect -498 -1210 -494 -1116
rect -474 -1210 -470 -1116
rect -450 -1210 -446 -1116
rect -426 -1210 -422 -1116
rect -402 -1210 -398 -1116
rect -378 -1210 -374 -1116
rect -354 -1141 -347 -1117
rect -354 -1210 -350 -1141
rect -330 -1210 -326 -1116
rect -306 -1210 -302 -1116
rect -282 -1210 -278 -1116
rect -258 -1210 -254 -1116
rect -234 -1210 -230 -1116
rect -210 -1210 -206 -1116
rect -186 -1210 -182 -1116
rect -162 -1210 -158 -1116
rect -138 -1210 -134 -1116
rect -114 -1210 -110 -1116
rect -90 -1186 -83 -1165
rect -66 -1186 -62 -1116
rect -42 -1186 -38 -1116
rect -18 -1186 -14 -1116
rect 6 -1186 10 -1116
rect 30 -1186 34 -1116
rect 54 -1186 58 -1116
rect 78 -1186 82 -1116
rect 91 -1123 96 -1116
rect 109 -1117 123 -1116
rect 126 -1117 133 -1093
rect 101 -1137 106 -1123
rect 102 -1186 106 -1137
rect 150 -1186 154 -1068
rect 174 -1186 178 -1068
rect 198 -1186 202 -1068
rect 222 -1186 226 -1068
rect 246 -1186 250 -1068
rect 270 -1186 274 -1068
rect 294 -1186 298 -1068
rect 318 -1186 322 -1068
rect 342 -1186 346 -1068
rect 366 -1186 370 -1068
rect 390 -1186 394 -1068
rect 414 -1186 418 -1068
rect 438 -1186 442 -1068
rect 462 -1186 466 -1068
rect 486 -1186 490 -1068
rect 510 -1186 514 -1068
rect 534 -1186 538 -1068
rect 558 -1186 562 -1068
rect 582 -1186 586 -1068
rect 606 -1185 610 -1068
rect 619 -1099 624 -1089
rect 630 -1099 634 -1068
rect 643 -1075 648 -1068
rect 654 -1075 658 -1068
rect 653 -1089 658 -1075
rect 629 -1113 634 -1099
rect 595 -1186 629 -1185
rect -107 -1188 629 -1186
rect -107 -1189 -93 -1188
rect -90 -1189 -83 -1188
rect -90 -1210 -86 -1189
rect -66 -1210 -62 -1188
rect -42 -1210 -38 -1188
rect -18 -1210 -14 -1188
rect 6 -1210 10 -1188
rect 30 -1210 34 -1188
rect 54 -1210 58 -1188
rect 78 -1210 82 -1188
rect 102 -1210 106 -1188
rect -2393 -1212 123 -1210
rect -2371 -1258 -2366 -1212
rect -2348 -1258 -2343 -1212
rect -2325 -1218 -2317 -1212
rect -2053 -1214 -1972 -1212
rect -2325 -1234 -2320 -1218
rect -2317 -1222 -2309 -1218
rect -2069 -1222 -2068 -1221
rect -2309 -1234 -2301 -1222
rect -2069 -1229 -2038 -1222
rect -2069 -1231 -2068 -1229
rect -2000 -1230 -1992 -1214
rect -1926 -1217 -1924 -1212
rect -1916 -1220 -1914 -1217
rect -1671 -1218 -1663 -1212
rect -1982 -1230 -1916 -1221
rect -1663 -1222 -1655 -1218
rect -2325 -1246 -2317 -1234
rect -2068 -1237 -2053 -1231
rect -2027 -1232 -1992 -1230
rect -2076 -1246 -2053 -1239
rect -2011 -1240 -2002 -1232
rect -2000 -1240 -1992 -1232
rect -1655 -1234 -1647 -1222
rect -2003 -1242 -1992 -1240
rect -2325 -1258 -2320 -1246
rect -2317 -1250 -2309 -1246
rect -2309 -1258 -2301 -1250
rect -2015 -1254 -2003 -1242
rect -2000 -1258 -1992 -1242
rect -1972 -1246 -1924 -1239
rect -1862 -1247 -1680 -1238
rect -1671 -1246 -1663 -1234
rect -1663 -1250 -1655 -1246
rect -1976 -1258 -1940 -1257
rect -1655 -1258 -1647 -1250
rect -1642 -1258 -1637 -1212
rect -1619 -1258 -1614 -1212
rect -1530 -1258 -1526 -1212
rect -1506 -1258 -1502 -1212
rect -1482 -1258 -1478 -1212
rect -1458 -1258 -1454 -1212
rect -1434 -1258 -1430 -1212
rect -1410 -1258 -1406 -1212
rect -1386 -1258 -1382 -1212
rect -1362 -1258 -1358 -1212
rect -1338 -1258 -1334 -1212
rect -1314 -1258 -1310 -1212
rect -1290 -1258 -1286 -1212
rect -1266 -1258 -1262 -1212
rect -1242 -1258 -1238 -1212
rect -1218 -1258 -1214 -1212
rect -1194 -1258 -1190 -1212
rect -1170 -1258 -1166 -1212
rect -1146 -1258 -1142 -1212
rect -1122 -1258 -1118 -1212
rect -1098 -1258 -1094 -1212
rect -1074 -1258 -1070 -1212
rect -1050 -1258 -1046 -1212
rect -1026 -1258 -1022 -1212
rect -1002 -1258 -998 -1212
rect -978 -1258 -974 -1212
rect -954 -1258 -950 -1212
rect -930 -1258 -926 -1212
rect -917 -1243 -912 -1233
rect -906 -1243 -902 -1212
rect -907 -1257 -902 -1243
rect -882 -1258 -878 -1212
rect -858 -1258 -854 -1212
rect -834 -1258 -830 -1212
rect -810 -1258 -806 -1212
rect -786 -1258 -782 -1212
rect -762 -1258 -758 -1212
rect -738 -1258 -734 -1212
rect -714 -1258 -710 -1212
rect -690 -1258 -686 -1212
rect -666 -1258 -662 -1212
rect -642 -1258 -638 -1212
rect -618 -1258 -614 -1212
rect -594 -1258 -590 -1212
rect -570 -1258 -566 -1212
rect -546 -1258 -542 -1212
rect -522 -1237 -518 -1212
rect -2393 -1260 -525 -1258
rect -2371 -1330 -2366 -1260
rect -2348 -1330 -2343 -1260
rect -2325 -1262 -2320 -1260
rect -2309 -1262 -2301 -1260
rect -2325 -1274 -2317 -1262
rect -2325 -1294 -2320 -1274
rect -2317 -1278 -2309 -1274
rect -2325 -1302 -2317 -1294
rect -2060 -1300 -2030 -1297
rect -2325 -1330 -2320 -1302
rect -2317 -1310 -2309 -1302
rect -2060 -1313 -2038 -1302
rect -2033 -1309 -2030 -1300
rect -2028 -1304 -2027 -1300
rect -2068 -1318 -2038 -1315
rect -2000 -1330 -1992 -1260
rect -1655 -1262 -1647 -1260
rect -1671 -1274 -1663 -1262
rect -1663 -1278 -1655 -1274
rect -1912 -1285 -1884 -1283
rect -1852 -1291 -1804 -1287
rect -1844 -1300 -1796 -1297
rect -1671 -1302 -1663 -1294
rect -1844 -1313 -1804 -1302
rect -1663 -1310 -1655 -1302
rect -1852 -1318 -1680 -1314
rect -1642 -1330 -1637 -1260
rect -1619 -1330 -1614 -1260
rect -1530 -1330 -1526 -1260
rect -1506 -1330 -1502 -1260
rect -1482 -1330 -1478 -1260
rect -1458 -1330 -1454 -1260
rect -1434 -1330 -1430 -1260
rect -1410 -1330 -1406 -1260
rect -1386 -1330 -1382 -1260
rect -1362 -1330 -1358 -1260
rect -1338 -1330 -1334 -1260
rect -1314 -1330 -1310 -1260
rect -1290 -1330 -1286 -1260
rect -1266 -1330 -1262 -1260
rect -1242 -1330 -1238 -1260
rect -1218 -1330 -1214 -1260
rect -1194 -1330 -1190 -1260
rect -1170 -1330 -1166 -1260
rect -1146 -1330 -1142 -1260
rect -1122 -1330 -1118 -1260
rect -1098 -1330 -1094 -1260
rect -1074 -1330 -1070 -1260
rect -1050 -1330 -1046 -1260
rect -1026 -1330 -1022 -1260
rect -1002 -1330 -998 -1260
rect -978 -1330 -974 -1260
rect -954 -1330 -950 -1260
rect -930 -1330 -926 -1260
rect -917 -1291 -912 -1281
rect -907 -1305 -902 -1291
rect -906 -1330 -902 -1305
rect -882 -1309 -878 -1260
rect -2393 -1332 -885 -1330
rect -2371 -1354 -2366 -1332
rect -2348 -1354 -2343 -1332
rect -2325 -1354 -2320 -1332
rect -2309 -1350 -2301 -1340
rect -2068 -1349 -2062 -1344
rect -2317 -1354 -2309 -1350
rect -2060 -1354 -2050 -1349
rect -2000 -1354 -1992 -1332
rect -1806 -1340 -1680 -1334
rect -1854 -1349 -1806 -1344
rect -1655 -1350 -1647 -1340
rect -1972 -1354 -1964 -1353
rect -1958 -1354 -1942 -1352
rect -1844 -1354 -1806 -1351
rect -1663 -1354 -1655 -1350
rect -1642 -1354 -1637 -1332
rect -1619 -1354 -1614 -1332
rect -1530 -1354 -1526 -1332
rect -1506 -1354 -1502 -1332
rect -1482 -1354 -1478 -1332
rect -1458 -1354 -1454 -1332
rect -1434 -1354 -1430 -1332
rect -1410 -1354 -1406 -1332
rect -1386 -1354 -1382 -1332
rect -1362 -1354 -1358 -1332
rect -1338 -1354 -1334 -1332
rect -1314 -1354 -1310 -1332
rect -1290 -1354 -1286 -1332
rect -1266 -1354 -1262 -1332
rect -1242 -1354 -1238 -1332
rect -1218 -1354 -1214 -1332
rect -1194 -1354 -1190 -1332
rect -1170 -1354 -1166 -1332
rect -1146 -1354 -1142 -1332
rect -1122 -1354 -1118 -1332
rect -1098 -1354 -1094 -1332
rect -1074 -1354 -1070 -1332
rect -1050 -1354 -1046 -1332
rect -1026 -1354 -1022 -1332
rect -1002 -1354 -998 -1332
rect -978 -1354 -974 -1332
rect -954 -1354 -950 -1332
rect -930 -1354 -926 -1332
rect -906 -1354 -902 -1332
rect -899 -1333 -885 -1332
rect -882 -1333 -875 -1309
rect -858 -1354 -854 -1260
rect -834 -1354 -830 -1260
rect -810 -1354 -806 -1260
rect -786 -1354 -782 -1260
rect -762 -1354 -758 -1260
rect -738 -1354 -734 -1260
rect -714 -1354 -710 -1260
rect -690 -1354 -686 -1260
rect -666 -1354 -662 -1260
rect -642 -1354 -638 -1260
rect -618 -1354 -614 -1260
rect -594 -1353 -590 -1260
rect -605 -1354 -571 -1353
rect -2393 -1356 -571 -1354
rect -2371 -1378 -2366 -1356
rect -2348 -1378 -2343 -1356
rect -2325 -1378 -2320 -1356
rect -2060 -1362 -2050 -1356
rect -2309 -1378 -2301 -1368
rect -2060 -1369 -2030 -1362
rect -2000 -1366 -1992 -1356
rect -1972 -1358 -1942 -1356
rect -1958 -1359 -1942 -1358
rect -1844 -1360 -1806 -1356
rect -2068 -1376 -2062 -1369
rect -2062 -1378 -2036 -1376
rect -2393 -1380 -2036 -1378
rect -2030 -1378 -2012 -1376
rect -2004 -1378 -1990 -1366
rect -1844 -1367 -1798 -1362
rect -1806 -1369 -1798 -1367
rect -1854 -1371 -1844 -1369
rect -1854 -1376 -1806 -1371
rect -1864 -1378 -1796 -1377
rect -1655 -1378 -1647 -1368
rect -1642 -1378 -1637 -1356
rect -1619 -1378 -1614 -1356
rect -1530 -1378 -1526 -1356
rect -1506 -1378 -1502 -1356
rect -1482 -1378 -1478 -1356
rect -1458 -1378 -1454 -1356
rect -1434 -1378 -1430 -1356
rect -1410 -1378 -1406 -1356
rect -1386 -1378 -1382 -1356
rect -1362 -1378 -1358 -1356
rect -1338 -1378 -1334 -1356
rect -1314 -1378 -1310 -1356
rect -1290 -1378 -1286 -1356
rect -1266 -1378 -1262 -1356
rect -1242 -1378 -1238 -1356
rect -1218 -1378 -1214 -1356
rect -1194 -1378 -1190 -1356
rect -1170 -1378 -1166 -1356
rect -1146 -1378 -1142 -1356
rect -1122 -1378 -1118 -1356
rect -1098 -1378 -1094 -1356
rect -1074 -1378 -1070 -1356
rect -1050 -1378 -1046 -1356
rect -1026 -1378 -1022 -1356
rect -1002 -1378 -998 -1356
rect -978 -1378 -974 -1356
rect -954 -1378 -950 -1356
rect -930 -1378 -926 -1356
rect -906 -1378 -902 -1356
rect -882 -1378 -875 -1357
rect -858 -1378 -854 -1356
rect -834 -1378 -830 -1356
rect -810 -1378 -806 -1356
rect -786 -1378 -782 -1356
rect -762 -1378 -758 -1356
rect -738 -1378 -734 -1356
rect -714 -1378 -710 -1356
rect -690 -1378 -686 -1356
rect -666 -1378 -662 -1356
rect -642 -1378 -638 -1356
rect -618 -1378 -614 -1356
rect -605 -1363 -600 -1356
rect -594 -1363 -590 -1356
rect -595 -1377 -590 -1363
rect -605 -1378 -571 -1377
rect -570 -1378 -566 -1260
rect -546 -1378 -542 -1260
rect -539 -1261 -525 -1260
rect -522 -1282 -515 -1237
rect -498 -1282 -494 -1212
rect -474 -1282 -470 -1212
rect -450 -1282 -446 -1212
rect -437 -1267 -432 -1257
rect -426 -1267 -422 -1212
rect -427 -1281 -422 -1267
rect -402 -1282 -398 -1212
rect -378 -1282 -374 -1212
rect -354 -1282 -350 -1212
rect -330 -1282 -326 -1212
rect -306 -1282 -302 -1212
rect -282 -1282 -278 -1212
rect -258 -1282 -254 -1212
rect -234 -1282 -230 -1212
rect -210 -1282 -206 -1212
rect -186 -1282 -182 -1212
rect -162 -1282 -158 -1212
rect -138 -1282 -134 -1212
rect -114 -1282 -110 -1212
rect -90 -1281 -86 -1212
rect -101 -1282 -67 -1281
rect -539 -1284 -67 -1282
rect -539 -1285 -525 -1284
rect -522 -1285 -515 -1284
rect -522 -1378 -518 -1285
rect -498 -1378 -494 -1284
rect -474 -1378 -470 -1284
rect -450 -1378 -446 -1284
rect -437 -1306 -403 -1305
rect -402 -1306 -398 -1284
rect -378 -1306 -374 -1284
rect -354 -1306 -350 -1284
rect -330 -1306 -326 -1284
rect -306 -1306 -302 -1284
rect -282 -1306 -278 -1284
rect -258 -1306 -254 -1284
rect -234 -1306 -230 -1284
rect -210 -1306 -206 -1284
rect -186 -1306 -182 -1284
rect -162 -1306 -158 -1284
rect -138 -1306 -134 -1284
rect -114 -1306 -110 -1284
rect -101 -1291 -96 -1284
rect -90 -1291 -86 -1284
rect -91 -1305 -86 -1291
rect -66 -1306 -62 -1212
rect -42 -1306 -38 -1212
rect -18 -1306 -14 -1212
rect 6 -1306 10 -1212
rect 30 -1306 34 -1212
rect 54 -1306 58 -1212
rect 78 -1306 82 -1212
rect 102 -1306 106 -1212
rect 109 -1213 123 -1212
rect 126 -1213 133 -1189
rect 126 -1306 130 -1213
rect 150 -1306 154 -1188
rect 174 -1306 178 -1188
rect 198 -1306 202 -1188
rect 222 -1306 226 -1188
rect 246 -1306 250 -1188
rect 270 -1306 274 -1188
rect 294 -1306 298 -1188
rect 318 -1306 322 -1188
rect 342 -1306 346 -1188
rect 366 -1306 370 -1188
rect 390 -1306 394 -1188
rect 414 -1306 418 -1188
rect 438 -1306 442 -1188
rect 462 -1306 466 -1188
rect 486 -1306 490 -1188
rect 510 -1306 514 -1188
rect 534 -1306 538 -1188
rect 558 -1306 562 -1188
rect 582 -1306 586 -1188
rect 595 -1195 600 -1188
rect 606 -1195 610 -1188
rect 605 -1209 610 -1195
rect 595 -1219 600 -1209
rect 605 -1233 610 -1219
rect 606 -1305 610 -1233
rect 595 -1306 627 -1305
rect -437 -1308 627 -1306
rect -437 -1315 -432 -1308
rect -427 -1329 -422 -1315
rect -426 -1378 -422 -1329
rect -402 -1333 -398 -1308
rect -402 -1357 -395 -1333
rect -378 -1378 -374 -1308
rect -354 -1378 -350 -1308
rect -330 -1378 -326 -1308
rect -306 -1378 -302 -1308
rect -282 -1378 -278 -1308
rect -258 -1378 -254 -1308
rect -234 -1378 -230 -1308
rect -210 -1378 -206 -1308
rect -186 -1378 -182 -1308
rect -162 -1378 -158 -1308
rect -138 -1378 -134 -1308
rect -114 -1378 -110 -1308
rect -101 -1339 -96 -1329
rect -91 -1353 -86 -1339
rect -90 -1378 -86 -1353
rect -66 -1357 -62 -1308
rect -2030 -1380 -69 -1378
rect -2371 -1426 -2366 -1380
rect -2348 -1426 -2343 -1380
rect -2325 -1426 -2320 -1380
rect -2317 -1384 -2309 -1380
rect -2060 -1384 -2050 -1380
rect -2060 -1386 -2036 -1384
rect -2060 -1388 -2030 -1386
rect -2292 -1394 -2030 -1388
rect -2092 -1410 -2062 -1408
rect -2094 -1414 -2062 -1410
rect -2000 -1426 -1992 -1380
rect -1844 -1387 -1806 -1380
rect -1663 -1384 -1655 -1380
rect -1844 -1394 -1680 -1388
rect -1854 -1410 -1806 -1408
rect -1854 -1414 -1680 -1410
rect -1642 -1426 -1637 -1380
rect -1619 -1426 -1614 -1380
rect -1530 -1426 -1526 -1380
rect -1506 -1426 -1502 -1380
rect -1482 -1426 -1478 -1380
rect -1458 -1426 -1454 -1380
rect -1434 -1426 -1430 -1380
rect -1410 -1426 -1406 -1380
rect -1386 -1426 -1382 -1380
rect -1362 -1426 -1358 -1380
rect -1338 -1426 -1334 -1380
rect -1314 -1426 -1310 -1380
rect -1290 -1426 -1286 -1380
rect -1266 -1426 -1262 -1380
rect -1242 -1426 -1238 -1380
rect -1218 -1426 -1214 -1380
rect -1194 -1426 -1190 -1380
rect -1170 -1426 -1166 -1380
rect -1146 -1426 -1142 -1380
rect -1122 -1426 -1118 -1380
rect -1098 -1426 -1094 -1380
rect -1074 -1426 -1070 -1380
rect -1050 -1426 -1046 -1380
rect -1026 -1426 -1022 -1380
rect -1002 -1426 -998 -1380
rect -978 -1426 -974 -1380
rect -954 -1426 -950 -1380
rect -930 -1426 -926 -1380
rect -906 -1426 -902 -1380
rect -899 -1381 -885 -1380
rect -882 -1381 -875 -1380
rect -882 -1426 -878 -1381
rect -858 -1426 -854 -1380
rect -834 -1426 -830 -1380
rect -810 -1426 -806 -1380
rect -786 -1426 -782 -1380
rect -762 -1426 -758 -1380
rect -738 -1426 -734 -1380
rect -714 -1426 -710 -1380
rect -690 -1426 -686 -1380
rect -666 -1426 -662 -1380
rect -642 -1426 -638 -1380
rect -618 -1426 -614 -1380
rect -605 -1387 -600 -1380
rect -595 -1401 -590 -1387
rect -594 -1426 -590 -1401
rect -570 -1426 -566 -1380
rect -546 -1426 -542 -1380
rect -522 -1426 -518 -1380
rect -498 -1426 -494 -1380
rect -474 -1426 -470 -1380
rect -450 -1426 -446 -1380
rect -426 -1426 -422 -1380
rect -402 -1405 -395 -1381
rect -402 -1426 -398 -1405
rect -378 -1426 -374 -1380
rect -354 -1426 -350 -1380
rect -330 -1426 -326 -1380
rect -306 -1426 -302 -1380
rect -282 -1426 -278 -1380
rect -258 -1426 -254 -1380
rect -234 -1426 -230 -1380
rect -210 -1426 -206 -1380
rect -186 -1426 -182 -1380
rect -162 -1426 -158 -1380
rect -138 -1426 -134 -1380
rect -114 -1426 -110 -1380
rect -90 -1426 -86 -1380
rect -83 -1381 -69 -1380
rect -66 -1381 -59 -1357
rect -2393 -1428 -69 -1426
rect -2371 -1450 -2366 -1428
rect -2348 -1450 -2343 -1428
rect -2325 -1450 -2320 -1428
rect -2072 -1430 -2036 -1429
rect -2072 -1436 -2054 -1430
rect -2309 -1444 -2301 -1436
rect -2317 -1450 -2309 -1444
rect -2092 -1445 -2062 -1440
rect -2000 -1449 -1992 -1428
rect -1938 -1429 -1906 -1428
rect -1920 -1430 -1906 -1429
rect -1806 -1436 -1680 -1430
rect -1854 -1445 -1806 -1440
rect -1655 -1444 -1647 -1436
rect -1982 -1449 -1966 -1448
rect -2000 -1450 -1966 -1449
rect -1846 -1450 -1806 -1447
rect -1663 -1450 -1655 -1444
rect -1642 -1450 -1637 -1428
rect -1619 -1450 -1614 -1428
rect -1530 -1450 -1526 -1428
rect -1506 -1450 -1502 -1428
rect -1482 -1450 -1478 -1428
rect -1458 -1450 -1454 -1428
rect -1434 -1450 -1430 -1428
rect -1410 -1450 -1406 -1428
rect -1386 -1450 -1382 -1428
rect -1362 -1450 -1358 -1428
rect -1338 -1450 -1334 -1428
rect -1314 -1450 -1310 -1428
rect -1290 -1450 -1286 -1428
rect -1266 -1450 -1262 -1428
rect -1242 -1450 -1238 -1428
rect -1218 -1450 -1214 -1428
rect -1194 -1450 -1190 -1428
rect -1170 -1450 -1166 -1428
rect -1146 -1450 -1142 -1428
rect -1122 -1450 -1118 -1428
rect -1098 -1450 -1094 -1428
rect -1074 -1450 -1070 -1428
rect -1050 -1450 -1046 -1428
rect -1026 -1450 -1022 -1428
rect -1002 -1450 -998 -1428
rect -978 -1450 -974 -1428
rect -954 -1450 -950 -1428
rect -930 -1450 -926 -1428
rect -906 -1450 -902 -1428
rect -882 -1450 -878 -1428
rect -858 -1450 -854 -1428
rect -834 -1450 -830 -1428
rect -810 -1450 -806 -1428
rect -786 -1450 -782 -1428
rect -762 -1450 -758 -1428
rect -738 -1450 -734 -1428
rect -714 -1450 -710 -1428
rect -690 -1450 -686 -1428
rect -666 -1450 -662 -1428
rect -642 -1450 -638 -1428
rect -618 -1450 -614 -1428
rect -594 -1450 -590 -1428
rect -570 -1429 -566 -1428
rect -2393 -1452 -573 -1450
rect -2371 -1474 -2366 -1452
rect -2348 -1474 -2343 -1452
rect -2325 -1474 -2320 -1452
rect -2000 -1454 -1966 -1452
rect -2309 -1472 -2301 -1464
rect -2062 -1465 -2054 -1458
rect -2092 -1472 -2084 -1465
rect -2062 -1472 -2026 -1470
rect -2317 -1474 -2309 -1472
rect -2062 -1474 -2012 -1472
rect -2000 -1474 -1992 -1454
rect -1982 -1455 -1966 -1454
rect -1846 -1456 -1806 -1452
rect -1846 -1463 -1798 -1458
rect -1806 -1465 -1798 -1463
rect -1854 -1467 -1846 -1465
rect -1854 -1472 -1806 -1467
rect -1655 -1472 -1647 -1464
rect -1864 -1474 -1796 -1473
rect -1663 -1474 -1655 -1472
rect -1642 -1474 -1637 -1452
rect -1619 -1474 -1614 -1452
rect -1530 -1474 -1526 -1452
rect -1506 -1474 -1502 -1452
rect -1482 -1474 -1478 -1452
rect -1458 -1474 -1454 -1452
rect -1434 -1474 -1430 -1452
rect -1410 -1474 -1406 -1452
rect -1386 -1474 -1382 -1452
rect -1362 -1474 -1358 -1452
rect -1338 -1474 -1334 -1452
rect -1314 -1474 -1310 -1452
rect -1290 -1474 -1286 -1452
rect -1266 -1474 -1262 -1452
rect -1242 -1474 -1238 -1452
rect -1218 -1474 -1214 -1452
rect -1194 -1474 -1190 -1452
rect -1170 -1474 -1166 -1452
rect -1146 -1474 -1142 -1452
rect -1122 -1474 -1118 -1452
rect -1098 -1474 -1094 -1452
rect -1074 -1474 -1070 -1452
rect -1050 -1474 -1046 -1452
rect -1026 -1474 -1022 -1452
rect -1002 -1474 -998 -1452
rect -978 -1474 -974 -1452
rect -954 -1474 -950 -1452
rect -930 -1474 -926 -1452
rect -906 -1474 -902 -1452
rect -882 -1474 -878 -1452
rect -858 -1474 -854 -1452
rect -834 -1474 -830 -1452
rect -810 -1474 -806 -1452
rect -786 -1474 -782 -1452
rect -762 -1474 -758 -1452
rect -738 -1474 -734 -1452
rect -714 -1474 -710 -1452
rect -690 -1474 -686 -1452
rect -666 -1474 -662 -1452
rect -642 -1474 -638 -1452
rect -618 -1474 -614 -1452
rect -594 -1474 -590 -1452
rect -587 -1453 -573 -1452
rect -570 -1474 -563 -1429
rect -546 -1474 -542 -1428
rect -522 -1474 -518 -1428
rect -498 -1474 -494 -1428
rect -474 -1474 -470 -1428
rect -450 -1474 -446 -1428
rect -426 -1474 -422 -1428
rect -402 -1474 -398 -1428
rect -378 -1474 -374 -1428
rect -354 -1474 -350 -1428
rect -330 -1474 -326 -1428
rect -306 -1474 -302 -1428
rect -282 -1474 -278 -1428
rect -258 -1474 -254 -1428
rect -234 -1474 -230 -1428
rect -210 -1474 -206 -1428
rect -186 -1474 -182 -1428
rect -162 -1474 -158 -1428
rect -138 -1474 -134 -1428
rect -114 -1474 -110 -1428
rect -90 -1474 -86 -1428
rect -83 -1429 -69 -1428
rect -66 -1429 -59 -1405
rect -66 -1474 -62 -1429
rect -42 -1474 -38 -1308
rect -18 -1474 -14 -1308
rect 6 -1474 10 -1308
rect 30 -1474 34 -1308
rect 54 -1474 58 -1308
rect 78 -1474 82 -1308
rect 102 -1474 106 -1308
rect 126 -1474 130 -1308
rect 150 -1474 154 -1308
rect 174 -1474 178 -1308
rect 198 -1474 202 -1308
rect 222 -1474 226 -1308
rect 246 -1474 250 -1308
rect 270 -1474 274 -1308
rect 294 -1474 298 -1308
rect 318 -1474 322 -1308
rect 342 -1474 346 -1308
rect 366 -1474 370 -1308
rect 379 -1459 384 -1449
rect 390 -1459 394 -1308
rect 389 -1473 394 -1459
rect 390 -1474 394 -1473
rect 414 -1474 418 -1308
rect 438 -1474 442 -1308
rect 462 -1474 466 -1308
rect 475 -1387 480 -1377
rect 486 -1387 490 -1308
rect 485 -1401 490 -1387
rect 475 -1402 509 -1401
rect 510 -1402 514 -1308
rect 534 -1402 538 -1308
rect 558 -1402 562 -1308
rect 582 -1401 586 -1308
rect 595 -1315 600 -1308
rect 606 -1315 610 -1308
rect 613 -1309 627 -1308
rect 605 -1329 610 -1315
rect 571 -1402 605 -1401
rect 475 -1404 605 -1402
rect 475 -1411 480 -1404
rect 485 -1425 490 -1411
rect 486 -1474 490 -1425
rect 510 -1453 514 -1404
rect 499 -1474 507 -1473
rect -2393 -1476 507 -1474
rect -2371 -1522 -2366 -1476
rect -2348 -1522 -2343 -1476
rect -2325 -1522 -2320 -1476
rect -2317 -1480 -2309 -1476
rect -2062 -1480 -2054 -1476
rect -2154 -1484 -2138 -1482
rect -2057 -1484 -2054 -1480
rect -2292 -1490 -2054 -1484
rect -2052 -1490 -2044 -1480
rect -2092 -1506 -2062 -1504
rect -2094 -1510 -2062 -1506
rect -2000 -1522 -1992 -1476
rect -1846 -1483 -1806 -1476
rect -1663 -1480 -1655 -1476
rect -1846 -1490 -1680 -1484
rect -1854 -1506 -1806 -1504
rect -1854 -1510 -1680 -1506
rect -1642 -1522 -1637 -1476
rect -1619 -1522 -1614 -1476
rect -1530 -1522 -1526 -1476
rect -1506 -1522 -1502 -1476
rect -1482 -1522 -1478 -1476
rect -1458 -1522 -1454 -1476
rect -1434 -1522 -1430 -1476
rect -1410 -1522 -1406 -1476
rect -1386 -1522 -1382 -1476
rect -1362 -1522 -1358 -1476
rect -1338 -1522 -1334 -1476
rect -1314 -1522 -1310 -1476
rect -1290 -1522 -1286 -1476
rect -1266 -1522 -1262 -1476
rect -1242 -1522 -1238 -1476
rect -1218 -1522 -1214 -1476
rect -1194 -1522 -1190 -1476
rect -1170 -1522 -1166 -1476
rect -1146 -1522 -1142 -1476
rect -1122 -1522 -1118 -1476
rect -1098 -1522 -1094 -1476
rect -1074 -1522 -1070 -1476
rect -1050 -1522 -1046 -1476
rect -1026 -1522 -1022 -1476
rect -1002 -1522 -998 -1476
rect -978 -1522 -974 -1476
rect -954 -1522 -950 -1476
rect -930 -1522 -926 -1476
rect -906 -1522 -902 -1476
rect -882 -1522 -878 -1476
rect -858 -1522 -854 -1476
rect -834 -1522 -830 -1476
rect -810 -1522 -806 -1476
rect -786 -1522 -782 -1476
rect -762 -1522 -758 -1476
rect -738 -1522 -734 -1476
rect -714 -1522 -710 -1476
rect -690 -1522 -686 -1476
rect -666 -1522 -662 -1476
rect -642 -1522 -638 -1476
rect -618 -1522 -614 -1476
rect -594 -1522 -590 -1476
rect -587 -1477 -573 -1476
rect -570 -1477 -563 -1476
rect -570 -1522 -566 -1477
rect -546 -1522 -542 -1476
rect -522 -1522 -518 -1476
rect -498 -1522 -494 -1476
rect -474 -1522 -470 -1476
rect -450 -1522 -446 -1476
rect -426 -1522 -422 -1476
rect -402 -1522 -398 -1476
rect -378 -1522 -374 -1476
rect -354 -1522 -350 -1476
rect -330 -1522 -326 -1476
rect -306 -1522 -302 -1476
rect -282 -1522 -278 -1476
rect -258 -1522 -254 -1476
rect -234 -1522 -230 -1476
rect -210 -1522 -206 -1476
rect -186 -1522 -182 -1476
rect -162 -1522 -158 -1476
rect -138 -1522 -134 -1476
rect -114 -1522 -110 -1476
rect -90 -1522 -86 -1476
rect -66 -1522 -62 -1476
rect -42 -1522 -38 -1476
rect -18 -1522 -14 -1476
rect 6 -1522 10 -1476
rect 30 -1522 34 -1476
rect 54 -1522 58 -1476
rect 78 -1522 82 -1476
rect 102 -1522 106 -1476
rect 126 -1522 130 -1476
rect 150 -1522 154 -1476
rect 174 -1522 178 -1476
rect 198 -1522 202 -1476
rect 222 -1522 226 -1476
rect 246 -1522 250 -1476
rect 270 -1522 274 -1476
rect 294 -1522 298 -1476
rect 318 -1522 322 -1476
rect 342 -1522 346 -1476
rect 366 -1522 370 -1476
rect 390 -1522 394 -1476
rect 414 -1522 418 -1476
rect 438 -1522 442 -1476
rect 462 -1522 466 -1476
rect 486 -1522 490 -1476
rect 493 -1477 507 -1476
rect 510 -1483 517 -1453
rect 509 -1497 517 -1483
rect 510 -1501 517 -1497
rect 510 -1522 514 -1501
rect 534 -1522 538 -1404
rect 558 -1522 562 -1404
rect 571 -1411 576 -1404
rect 582 -1411 586 -1404
rect 581 -1425 586 -1411
rect 571 -1435 576 -1425
rect 581 -1449 586 -1435
rect 582 -1522 586 -1449
rect 595 -1522 603 -1521
rect -2393 -1524 603 -1522
rect -2371 -1546 -2366 -1524
rect -2348 -1546 -2343 -1524
rect -2325 -1546 -2320 -1524
rect -2072 -1526 -2036 -1525
rect -2072 -1532 -2054 -1526
rect -2309 -1540 -2301 -1532
rect -2317 -1546 -2309 -1540
rect -2092 -1541 -2062 -1536
rect -2000 -1545 -1992 -1524
rect -1938 -1525 -1906 -1524
rect -1920 -1526 -1906 -1525
rect -1806 -1532 -1680 -1526
rect -1854 -1541 -1806 -1536
rect -1655 -1540 -1647 -1532
rect -1982 -1545 -1966 -1544
rect -2000 -1546 -1966 -1545
rect -1846 -1546 -1806 -1543
rect -1663 -1546 -1655 -1540
rect -1642 -1546 -1637 -1524
rect -1619 -1546 -1614 -1524
rect -1530 -1546 -1526 -1524
rect -1506 -1546 -1502 -1524
rect -1482 -1546 -1478 -1524
rect -1458 -1546 -1454 -1524
rect -1434 -1546 -1430 -1524
rect -1410 -1546 -1406 -1524
rect -1386 -1546 -1382 -1524
rect -1362 -1546 -1358 -1524
rect -1338 -1546 -1334 -1524
rect -1314 -1546 -1310 -1524
rect -1290 -1546 -1286 -1524
rect -1266 -1546 -1262 -1524
rect -1242 -1546 -1238 -1524
rect -1218 -1546 -1214 -1524
rect -1194 -1546 -1190 -1524
rect -1170 -1546 -1166 -1524
rect -1146 -1546 -1142 -1524
rect -1122 -1546 -1118 -1524
rect -1098 -1546 -1094 -1524
rect -1074 -1546 -1070 -1524
rect -1050 -1546 -1046 -1524
rect -1026 -1546 -1022 -1524
rect -1002 -1546 -998 -1524
rect -978 -1546 -974 -1524
rect -954 -1546 -950 -1524
rect -930 -1546 -926 -1524
rect -906 -1546 -902 -1524
rect -882 -1546 -878 -1524
rect -858 -1546 -854 -1524
rect -834 -1546 -830 -1524
rect -810 -1546 -806 -1524
rect -786 -1546 -782 -1524
rect -762 -1546 -758 -1524
rect -738 -1546 -734 -1524
rect -714 -1546 -710 -1524
rect -690 -1546 -686 -1524
rect -666 -1546 -662 -1524
rect -642 -1546 -638 -1524
rect -618 -1546 -614 -1524
rect -594 -1546 -590 -1524
rect -570 -1546 -566 -1524
rect -546 -1546 -542 -1524
rect -522 -1546 -518 -1524
rect -498 -1546 -494 -1524
rect -474 -1546 -470 -1524
rect -450 -1546 -446 -1524
rect -426 -1546 -422 -1524
rect -402 -1546 -398 -1524
rect -378 -1546 -374 -1524
rect -354 -1546 -350 -1524
rect -330 -1546 -326 -1524
rect -306 -1546 -302 -1524
rect -282 -1546 -278 -1524
rect -258 -1546 -254 -1524
rect -234 -1546 -230 -1524
rect -210 -1546 -206 -1524
rect -186 -1546 -182 -1524
rect -162 -1546 -158 -1524
rect -138 -1546 -134 -1524
rect -114 -1546 -110 -1524
rect -90 -1546 -86 -1524
rect -66 -1545 -62 -1524
rect -77 -1546 -43 -1545
rect -2393 -1548 -43 -1546
rect -2371 -1570 -2366 -1548
rect -2348 -1570 -2343 -1548
rect -2325 -1570 -2320 -1548
rect -2000 -1550 -1966 -1548
rect -2309 -1568 -2301 -1560
rect -2062 -1561 -2054 -1554
rect -2092 -1568 -2084 -1561
rect -2062 -1568 -2026 -1566
rect -2317 -1570 -2309 -1568
rect -2062 -1570 -2012 -1568
rect -2000 -1570 -1992 -1550
rect -1982 -1551 -1966 -1550
rect -1846 -1552 -1806 -1548
rect -1846 -1559 -1798 -1554
rect -1806 -1561 -1798 -1559
rect -1854 -1563 -1846 -1561
rect -1854 -1568 -1806 -1563
rect -1655 -1568 -1647 -1560
rect -1864 -1570 -1796 -1569
rect -1663 -1570 -1655 -1568
rect -1642 -1570 -1637 -1548
rect -1619 -1570 -1614 -1548
rect -1530 -1570 -1526 -1548
rect -1506 -1570 -1502 -1548
rect -1482 -1570 -1478 -1548
rect -1458 -1570 -1454 -1548
rect -1434 -1570 -1430 -1548
rect -1410 -1570 -1406 -1548
rect -1386 -1570 -1382 -1548
rect -1362 -1570 -1358 -1548
rect -1338 -1570 -1334 -1548
rect -1314 -1570 -1310 -1548
rect -1290 -1570 -1286 -1548
rect -1266 -1570 -1262 -1548
rect -1242 -1570 -1238 -1548
rect -1218 -1570 -1214 -1548
rect -1194 -1570 -1190 -1548
rect -1170 -1570 -1166 -1548
rect -1146 -1570 -1142 -1548
rect -1122 -1570 -1118 -1548
rect -1098 -1570 -1094 -1548
rect -1074 -1570 -1070 -1548
rect -1050 -1570 -1046 -1548
rect -1026 -1570 -1022 -1548
rect -1002 -1570 -998 -1548
rect -978 -1570 -974 -1548
rect -954 -1570 -950 -1548
rect -930 -1570 -926 -1548
rect -906 -1570 -902 -1548
rect -882 -1570 -878 -1548
rect -858 -1570 -854 -1548
rect -834 -1570 -830 -1548
rect -810 -1570 -806 -1548
rect -786 -1570 -782 -1548
rect -762 -1570 -758 -1548
rect -738 -1570 -734 -1548
rect -714 -1570 -710 -1548
rect -690 -1570 -686 -1548
rect -666 -1570 -662 -1548
rect -642 -1570 -638 -1548
rect -618 -1570 -614 -1548
rect -594 -1569 -590 -1548
rect -605 -1570 -571 -1569
rect -2393 -1572 -571 -1570
rect -2371 -1618 -2366 -1572
rect -2348 -1618 -2343 -1572
rect -2325 -1618 -2320 -1572
rect -2317 -1576 -2309 -1572
rect -2062 -1576 -2054 -1572
rect -2154 -1580 -2138 -1578
rect -2057 -1580 -2054 -1576
rect -2292 -1586 -2054 -1580
rect -2052 -1586 -2044 -1576
rect -2092 -1602 -2062 -1600
rect -2094 -1606 -2062 -1602
rect -2000 -1618 -1992 -1572
rect -1846 -1579 -1806 -1572
rect -1663 -1576 -1655 -1572
rect -1846 -1586 -1680 -1580
rect -1854 -1602 -1806 -1600
rect -1854 -1606 -1680 -1602
rect -1642 -1618 -1637 -1572
rect -1619 -1618 -1614 -1572
rect -1530 -1618 -1526 -1572
rect -1506 -1618 -1502 -1572
rect -1482 -1618 -1478 -1572
rect -1458 -1618 -1454 -1572
rect -1434 -1618 -1430 -1572
rect -1410 -1618 -1406 -1572
rect -1386 -1618 -1382 -1572
rect -1362 -1618 -1358 -1572
rect -1338 -1618 -1334 -1572
rect -1314 -1618 -1310 -1572
rect -1290 -1618 -1286 -1572
rect -1266 -1618 -1262 -1572
rect -1242 -1618 -1238 -1572
rect -1218 -1618 -1214 -1572
rect -1194 -1618 -1190 -1572
rect -1170 -1618 -1166 -1572
rect -1146 -1618 -1142 -1572
rect -1122 -1618 -1118 -1572
rect -1098 -1618 -1094 -1572
rect -1074 -1618 -1070 -1572
rect -1050 -1618 -1046 -1572
rect -1026 -1618 -1022 -1572
rect -1002 -1618 -998 -1572
rect -978 -1618 -974 -1572
rect -954 -1618 -950 -1572
rect -930 -1618 -926 -1572
rect -906 -1618 -902 -1572
rect -882 -1618 -878 -1572
rect -858 -1618 -854 -1572
rect -834 -1618 -830 -1572
rect -810 -1618 -806 -1572
rect -786 -1618 -782 -1572
rect -762 -1618 -758 -1572
rect -738 -1618 -734 -1572
rect -714 -1618 -710 -1572
rect -690 -1618 -686 -1572
rect -666 -1618 -662 -1572
rect -642 -1618 -638 -1572
rect -618 -1618 -614 -1572
rect -605 -1579 -600 -1572
rect -594 -1579 -590 -1572
rect -595 -1593 -590 -1579
rect -594 -1618 -590 -1593
rect -570 -1618 -566 -1548
rect -546 -1618 -542 -1548
rect -522 -1618 -518 -1548
rect -498 -1618 -494 -1548
rect -474 -1618 -470 -1548
rect -450 -1618 -446 -1548
rect -426 -1618 -422 -1548
rect -402 -1618 -398 -1548
rect -378 -1618 -374 -1548
rect -354 -1618 -350 -1548
rect -330 -1618 -326 -1548
rect -306 -1618 -302 -1548
rect -282 -1618 -278 -1548
rect -258 -1618 -254 -1548
rect -234 -1618 -230 -1548
rect -210 -1618 -206 -1548
rect -186 -1618 -182 -1548
rect -162 -1618 -158 -1548
rect -138 -1618 -134 -1548
rect -114 -1618 -110 -1548
rect -90 -1618 -86 -1548
rect -77 -1555 -72 -1548
rect -66 -1555 -62 -1548
rect -67 -1569 -62 -1555
rect -77 -1570 -43 -1569
rect -42 -1570 -38 -1524
rect -18 -1570 -14 -1524
rect 6 -1570 10 -1524
rect 30 -1570 34 -1524
rect 54 -1570 58 -1524
rect 78 -1570 82 -1524
rect 102 -1570 106 -1524
rect 126 -1570 130 -1524
rect 150 -1570 154 -1524
rect 174 -1570 178 -1524
rect 198 -1570 202 -1524
rect 222 -1570 226 -1524
rect 246 -1570 250 -1524
rect 270 -1570 274 -1524
rect 294 -1570 298 -1524
rect 318 -1570 322 -1524
rect 342 -1570 346 -1524
rect 366 -1570 370 -1524
rect 390 -1570 394 -1524
rect 414 -1525 418 -1524
rect 414 -1549 421 -1525
rect 414 -1570 418 -1549
rect 438 -1570 442 -1524
rect 462 -1570 466 -1524
rect 486 -1570 490 -1524
rect 510 -1570 514 -1524
rect 534 -1549 538 -1524
rect -77 -1572 531 -1570
rect -77 -1579 -72 -1572
rect -67 -1593 -62 -1579
rect -66 -1618 -62 -1593
rect -42 -1618 -38 -1572
rect -18 -1618 -14 -1572
rect 6 -1618 10 -1572
rect 30 -1618 34 -1572
rect 54 -1618 58 -1572
rect 78 -1618 82 -1572
rect 102 -1618 106 -1572
rect 126 -1618 130 -1572
rect 150 -1618 154 -1572
rect 174 -1618 178 -1572
rect 198 -1618 202 -1572
rect 222 -1618 226 -1572
rect 246 -1618 250 -1572
rect 270 -1618 274 -1572
rect 294 -1618 298 -1572
rect 318 -1618 322 -1572
rect 342 -1618 346 -1572
rect 366 -1618 370 -1572
rect 390 -1618 394 -1572
rect 414 -1618 418 -1572
rect 438 -1618 442 -1572
rect 462 -1618 466 -1572
rect 486 -1618 490 -1572
rect 510 -1618 514 -1572
rect 517 -1573 531 -1572
rect 534 -1573 541 -1549
rect 534 -1618 538 -1573
rect 558 -1618 562 -1524
rect 582 -1618 586 -1524
rect 589 -1525 603 -1524
rect 595 -1531 600 -1525
rect 605 -1545 610 -1531
rect 595 -1579 600 -1569
rect 606 -1579 610 -1545
rect 605 -1593 610 -1579
rect 595 -1618 627 -1617
rect -2393 -1620 627 -1618
rect -2371 -1642 -2366 -1620
rect -2348 -1642 -2343 -1620
rect -2325 -1642 -2320 -1620
rect -2072 -1622 -2036 -1621
rect -2072 -1628 -2054 -1622
rect -2309 -1636 -2301 -1628
rect -2317 -1642 -2309 -1636
rect -2092 -1637 -2062 -1632
rect -2000 -1641 -1992 -1620
rect -1938 -1621 -1906 -1620
rect -1920 -1622 -1906 -1621
rect -1806 -1628 -1680 -1622
rect -1854 -1637 -1806 -1632
rect -1655 -1636 -1647 -1628
rect -1982 -1641 -1966 -1640
rect -2000 -1642 -1966 -1641
rect -1846 -1642 -1806 -1639
rect -1663 -1642 -1655 -1636
rect -1642 -1642 -1637 -1620
rect -1619 -1642 -1614 -1620
rect -1530 -1642 -1526 -1620
rect -1506 -1642 -1502 -1620
rect -1482 -1642 -1478 -1620
rect -1458 -1642 -1454 -1620
rect -1434 -1642 -1430 -1620
rect -1410 -1642 -1406 -1620
rect -1386 -1642 -1382 -1620
rect -1362 -1642 -1358 -1620
rect -1338 -1642 -1334 -1620
rect -1314 -1642 -1310 -1620
rect -1290 -1642 -1286 -1620
rect -1266 -1642 -1262 -1620
rect -1242 -1642 -1238 -1620
rect -1218 -1642 -1214 -1620
rect -1194 -1641 -1190 -1620
rect -1205 -1642 -1171 -1641
rect -2393 -1644 -1171 -1642
rect -2371 -1666 -2366 -1644
rect -2348 -1666 -2343 -1644
rect -2325 -1666 -2320 -1644
rect -2000 -1646 -1966 -1644
rect -2309 -1664 -2301 -1656
rect -2062 -1657 -2054 -1650
rect -2092 -1664 -2084 -1657
rect -2062 -1664 -2026 -1662
rect -2317 -1666 -2309 -1664
rect -2062 -1666 -2012 -1664
rect -2000 -1666 -1992 -1646
rect -1982 -1647 -1966 -1646
rect -1846 -1648 -1806 -1644
rect -1846 -1655 -1798 -1650
rect -1806 -1657 -1798 -1655
rect -1854 -1659 -1846 -1657
rect -1854 -1664 -1806 -1659
rect -1655 -1664 -1647 -1656
rect -1864 -1666 -1796 -1665
rect -1663 -1666 -1655 -1664
rect -1642 -1666 -1637 -1644
rect -1619 -1666 -1614 -1644
rect -1530 -1666 -1526 -1644
rect -1506 -1666 -1502 -1644
rect -1482 -1666 -1478 -1644
rect -1458 -1666 -1454 -1644
rect -1434 -1666 -1430 -1644
rect -1410 -1666 -1406 -1644
rect -1386 -1666 -1382 -1644
rect -1362 -1666 -1358 -1644
rect -1338 -1666 -1334 -1644
rect -1314 -1666 -1310 -1644
rect -1290 -1666 -1286 -1644
rect -1266 -1666 -1262 -1644
rect -1242 -1666 -1238 -1644
rect -1218 -1666 -1214 -1644
rect -1205 -1651 -1200 -1644
rect -1194 -1651 -1190 -1644
rect -1195 -1665 -1190 -1651
rect -1194 -1666 -1190 -1665
rect -1170 -1666 -1166 -1620
rect -1146 -1666 -1142 -1620
rect -1122 -1666 -1118 -1620
rect -1098 -1666 -1094 -1620
rect -1074 -1666 -1070 -1620
rect -1050 -1666 -1046 -1620
rect -1026 -1666 -1022 -1620
rect -1002 -1666 -998 -1620
rect -978 -1666 -974 -1620
rect -954 -1666 -950 -1620
rect -930 -1666 -926 -1620
rect -906 -1666 -902 -1620
rect -882 -1666 -878 -1620
rect -858 -1666 -854 -1620
rect -834 -1666 -830 -1620
rect -810 -1666 -806 -1620
rect -786 -1666 -782 -1620
rect -762 -1666 -758 -1620
rect -738 -1666 -734 -1620
rect -714 -1666 -710 -1620
rect -690 -1666 -686 -1620
rect -666 -1666 -662 -1620
rect -642 -1666 -638 -1620
rect -618 -1666 -614 -1620
rect -594 -1666 -590 -1620
rect -570 -1645 -566 -1620
rect -2393 -1668 -573 -1666
rect -2371 -1714 -2366 -1668
rect -2348 -1714 -2343 -1668
rect -2325 -1714 -2320 -1668
rect -2317 -1672 -2309 -1668
rect -2062 -1672 -2054 -1668
rect -2154 -1676 -2138 -1674
rect -2057 -1676 -2054 -1672
rect -2292 -1682 -2054 -1676
rect -2052 -1682 -2044 -1672
rect -2092 -1698 -2062 -1696
rect -2094 -1702 -2062 -1698
rect -2000 -1714 -1992 -1668
rect -1846 -1675 -1806 -1668
rect -1663 -1672 -1655 -1668
rect -1846 -1682 -1680 -1676
rect -1854 -1698 -1806 -1696
rect -1854 -1702 -1680 -1698
rect -1642 -1714 -1637 -1668
rect -1619 -1714 -1614 -1668
rect -1530 -1714 -1526 -1668
rect -1506 -1714 -1502 -1668
rect -1482 -1714 -1478 -1668
rect -1458 -1714 -1454 -1668
rect -1434 -1714 -1430 -1668
rect -1410 -1714 -1406 -1668
rect -1386 -1714 -1382 -1668
rect -1362 -1714 -1358 -1668
rect -1338 -1714 -1334 -1668
rect -1314 -1714 -1310 -1668
rect -1290 -1714 -1286 -1668
rect -1266 -1714 -1262 -1668
rect -1242 -1714 -1238 -1668
rect -1218 -1714 -1214 -1668
rect -1194 -1714 -1190 -1668
rect -1170 -1714 -1166 -1668
rect -1146 -1714 -1142 -1668
rect -1122 -1714 -1118 -1668
rect -1098 -1714 -1094 -1668
rect -1074 -1714 -1070 -1668
rect -1050 -1714 -1046 -1668
rect -1026 -1714 -1022 -1668
rect -1002 -1714 -998 -1668
rect -978 -1714 -974 -1668
rect -954 -1714 -950 -1668
rect -930 -1714 -926 -1668
rect -906 -1714 -902 -1668
rect -882 -1714 -878 -1668
rect -858 -1714 -854 -1668
rect -834 -1714 -830 -1668
rect -810 -1714 -806 -1668
rect -786 -1714 -782 -1668
rect -762 -1714 -758 -1668
rect -738 -1714 -734 -1668
rect -714 -1714 -710 -1668
rect -690 -1714 -686 -1668
rect -666 -1714 -662 -1668
rect -642 -1714 -638 -1668
rect -618 -1714 -614 -1668
rect -594 -1714 -590 -1668
rect -587 -1669 -573 -1668
rect -570 -1669 -563 -1645
rect -570 -1714 -566 -1669
rect -546 -1714 -542 -1620
rect -522 -1714 -518 -1620
rect -498 -1714 -494 -1620
rect -474 -1714 -470 -1620
rect -450 -1714 -446 -1620
rect -426 -1714 -422 -1620
rect -402 -1714 -398 -1620
rect -378 -1714 -374 -1620
rect -354 -1714 -350 -1620
rect -330 -1714 -326 -1620
rect -306 -1714 -302 -1620
rect -282 -1714 -278 -1620
rect -258 -1714 -254 -1620
rect -234 -1714 -230 -1620
rect -210 -1714 -206 -1620
rect -186 -1714 -182 -1620
rect -162 -1714 -158 -1620
rect -138 -1714 -134 -1620
rect -114 -1714 -110 -1620
rect -90 -1714 -86 -1620
rect -66 -1714 -62 -1620
rect -42 -1621 -38 -1620
rect -42 -1666 -35 -1621
rect -18 -1666 -14 -1620
rect 6 -1666 10 -1620
rect 30 -1666 34 -1620
rect 54 -1666 58 -1620
rect 78 -1666 82 -1620
rect 102 -1666 106 -1620
rect 126 -1666 130 -1620
rect 150 -1666 154 -1620
rect 174 -1666 178 -1620
rect 198 -1666 202 -1620
rect 222 -1666 226 -1620
rect 246 -1666 250 -1620
rect 270 -1666 274 -1620
rect 294 -1666 298 -1620
rect 318 -1666 322 -1620
rect 342 -1666 346 -1620
rect 366 -1666 370 -1620
rect 390 -1666 394 -1620
rect 414 -1666 418 -1620
rect 438 -1666 442 -1620
rect 462 -1666 466 -1620
rect 486 -1666 490 -1620
rect 510 -1665 514 -1620
rect 499 -1666 533 -1665
rect -59 -1668 533 -1666
rect -59 -1669 -45 -1668
rect -42 -1669 -35 -1668
rect -42 -1714 -38 -1669
rect -18 -1714 -14 -1668
rect 6 -1714 10 -1668
rect 30 -1714 34 -1668
rect 54 -1714 58 -1668
rect 78 -1714 82 -1668
rect 102 -1714 106 -1668
rect 126 -1714 130 -1668
rect 150 -1714 154 -1668
rect 174 -1714 178 -1668
rect 198 -1714 202 -1668
rect 222 -1714 226 -1668
rect 246 -1714 250 -1668
rect 270 -1714 274 -1668
rect 294 -1714 298 -1668
rect 318 -1714 322 -1668
rect 342 -1714 346 -1668
rect 366 -1714 370 -1668
rect 390 -1714 394 -1668
rect 414 -1714 418 -1668
rect 438 -1714 442 -1668
rect 462 -1714 466 -1668
rect 486 -1714 490 -1668
rect 499 -1675 504 -1668
rect 510 -1675 514 -1668
rect 509 -1689 514 -1675
rect 510 -1714 514 -1689
rect 534 -1714 538 -1620
rect 558 -1714 562 -1620
rect 582 -1714 586 -1620
rect 595 -1627 600 -1620
rect 613 -1621 627 -1620
rect 605 -1641 610 -1627
rect 606 -1714 610 -1641
rect 619 -1714 627 -1713
rect -2393 -1716 627 -1714
rect -2371 -1738 -2366 -1716
rect -2348 -1738 -2343 -1716
rect -2325 -1738 -2320 -1716
rect -2072 -1718 -2036 -1717
rect -2072 -1724 -2054 -1718
rect -2309 -1732 -2301 -1724
rect -2317 -1738 -2309 -1732
rect -2092 -1733 -2062 -1728
rect -2000 -1737 -1992 -1716
rect -1938 -1717 -1906 -1716
rect -1920 -1718 -1906 -1717
rect -1806 -1724 -1680 -1718
rect -1854 -1733 -1806 -1728
rect -1655 -1732 -1647 -1724
rect -1982 -1737 -1966 -1736
rect -2000 -1738 -1966 -1737
rect -1846 -1738 -1806 -1735
rect -1663 -1738 -1655 -1732
rect -1642 -1738 -1637 -1716
rect -1619 -1738 -1614 -1716
rect -1530 -1738 -1526 -1716
rect -1506 -1738 -1502 -1716
rect -1482 -1738 -1478 -1716
rect -1458 -1738 -1454 -1716
rect -1434 -1738 -1430 -1716
rect -1410 -1737 -1406 -1716
rect -1421 -1738 -1387 -1737
rect -2393 -1740 -1387 -1738
rect -2371 -1762 -2366 -1740
rect -2348 -1762 -2343 -1740
rect -2325 -1762 -2320 -1740
rect -2000 -1742 -1966 -1740
rect -2309 -1760 -2301 -1752
rect -2062 -1753 -2054 -1746
rect -2092 -1760 -2084 -1753
rect -2062 -1760 -2026 -1758
rect -2317 -1762 -2309 -1760
rect -2062 -1762 -2012 -1760
rect -2000 -1762 -1992 -1742
rect -1982 -1743 -1966 -1742
rect -1846 -1744 -1806 -1740
rect -1846 -1751 -1798 -1746
rect -1806 -1753 -1798 -1751
rect -1854 -1755 -1846 -1753
rect -1854 -1760 -1806 -1755
rect -1655 -1760 -1647 -1752
rect -1864 -1762 -1796 -1761
rect -1663 -1762 -1655 -1760
rect -1642 -1762 -1637 -1740
rect -1619 -1762 -1614 -1740
rect -1530 -1762 -1526 -1740
rect -1506 -1762 -1502 -1740
rect -1482 -1762 -1478 -1740
rect -1458 -1762 -1454 -1740
rect -1434 -1762 -1430 -1740
rect -1421 -1747 -1416 -1740
rect -1410 -1747 -1406 -1740
rect -1411 -1761 -1406 -1747
rect -1421 -1762 -1387 -1761
rect -1386 -1762 -1382 -1716
rect -1362 -1762 -1358 -1716
rect -1338 -1762 -1334 -1716
rect -1314 -1762 -1310 -1716
rect -1290 -1762 -1286 -1716
rect -1266 -1762 -1262 -1716
rect -1242 -1762 -1238 -1716
rect -1218 -1762 -1214 -1716
rect -1194 -1762 -1190 -1716
rect -1170 -1717 -1166 -1716
rect -1170 -1741 -1163 -1717
rect -1170 -1762 -1166 -1741
rect -1146 -1762 -1142 -1716
rect -1122 -1762 -1118 -1716
rect -1098 -1762 -1094 -1716
rect -1074 -1762 -1070 -1716
rect -1050 -1762 -1046 -1716
rect -1026 -1762 -1022 -1716
rect -1002 -1762 -998 -1716
rect -978 -1762 -974 -1716
rect -954 -1762 -950 -1716
rect -930 -1762 -926 -1716
rect -906 -1762 -902 -1716
rect -882 -1762 -878 -1716
rect -858 -1762 -854 -1716
rect -834 -1762 -830 -1716
rect -810 -1762 -806 -1716
rect -786 -1762 -782 -1716
rect -762 -1762 -758 -1716
rect -738 -1762 -734 -1716
rect -714 -1762 -710 -1716
rect -690 -1762 -686 -1716
rect -666 -1762 -662 -1716
rect -642 -1762 -638 -1716
rect -618 -1762 -614 -1716
rect -594 -1761 -590 -1716
rect -605 -1762 -571 -1761
rect -2393 -1764 -571 -1762
rect -2371 -1810 -2366 -1764
rect -2348 -1810 -2343 -1764
rect -2325 -1810 -2320 -1764
rect -2317 -1768 -2309 -1764
rect -2062 -1768 -2054 -1764
rect -2154 -1772 -2138 -1770
rect -2057 -1772 -2054 -1768
rect -2292 -1778 -2054 -1772
rect -2052 -1778 -2044 -1768
rect -2092 -1794 -2062 -1792
rect -2094 -1798 -2062 -1794
rect -2000 -1810 -1992 -1764
rect -1846 -1771 -1806 -1764
rect -1663 -1768 -1655 -1764
rect -1846 -1778 -1680 -1772
rect -1854 -1794 -1806 -1792
rect -1854 -1798 -1680 -1794
rect -1642 -1810 -1637 -1764
rect -1619 -1810 -1614 -1764
rect -1530 -1810 -1526 -1764
rect -1506 -1810 -1502 -1764
rect -1482 -1810 -1478 -1764
rect -1458 -1810 -1454 -1764
rect -1434 -1810 -1430 -1764
rect -1421 -1771 -1416 -1764
rect -1411 -1785 -1406 -1771
rect -1410 -1810 -1406 -1785
rect -1386 -1810 -1382 -1764
rect -1362 -1810 -1358 -1764
rect -1338 -1810 -1334 -1764
rect -1314 -1810 -1310 -1764
rect -1290 -1810 -1286 -1764
rect -1266 -1810 -1262 -1764
rect -1242 -1810 -1238 -1764
rect -1218 -1810 -1214 -1764
rect -1194 -1810 -1190 -1764
rect -1170 -1810 -1166 -1764
rect -1146 -1810 -1142 -1764
rect -1122 -1810 -1118 -1764
rect -1098 -1810 -1094 -1764
rect -1074 -1810 -1070 -1764
rect -1050 -1810 -1046 -1764
rect -1026 -1810 -1022 -1764
rect -1002 -1810 -998 -1764
rect -978 -1810 -974 -1764
rect -954 -1810 -950 -1764
rect -930 -1810 -926 -1764
rect -906 -1810 -902 -1764
rect -882 -1810 -878 -1764
rect -858 -1810 -854 -1764
rect -834 -1810 -830 -1764
rect -810 -1810 -806 -1764
rect -786 -1810 -782 -1764
rect -762 -1810 -758 -1764
rect -738 -1810 -734 -1764
rect -714 -1810 -710 -1764
rect -690 -1810 -686 -1764
rect -666 -1810 -662 -1764
rect -642 -1810 -638 -1764
rect -618 -1810 -614 -1764
rect -605 -1771 -600 -1764
rect -594 -1771 -590 -1764
rect -595 -1785 -590 -1771
rect -605 -1795 -600 -1785
rect -595 -1809 -590 -1795
rect -594 -1810 -590 -1809
rect -570 -1810 -566 -1716
rect -546 -1810 -542 -1716
rect -522 -1810 -518 -1716
rect -498 -1810 -494 -1716
rect -474 -1810 -470 -1716
rect -450 -1810 -446 -1716
rect -426 -1810 -422 -1716
rect -402 -1810 -398 -1716
rect -378 -1810 -374 -1716
rect -354 -1810 -350 -1716
rect -330 -1810 -326 -1716
rect -306 -1810 -302 -1716
rect -282 -1810 -278 -1716
rect -258 -1810 -254 -1716
rect -234 -1810 -230 -1716
rect -210 -1810 -206 -1716
rect -186 -1810 -182 -1716
rect -162 -1810 -158 -1716
rect -138 -1810 -134 -1716
rect -114 -1810 -110 -1716
rect -90 -1810 -86 -1716
rect -66 -1810 -62 -1716
rect -42 -1810 -38 -1716
rect -18 -1810 -14 -1716
rect 6 -1810 10 -1716
rect 30 -1810 34 -1716
rect 54 -1810 58 -1716
rect 78 -1810 82 -1716
rect 102 -1810 106 -1716
rect 126 -1810 130 -1716
rect 150 -1810 154 -1716
rect 174 -1810 178 -1716
rect 198 -1810 202 -1716
rect 222 -1810 226 -1716
rect 246 -1810 250 -1716
rect 270 -1810 274 -1716
rect 294 -1810 298 -1716
rect 318 -1810 322 -1716
rect 342 -1810 346 -1716
rect 366 -1810 370 -1716
rect 390 -1810 394 -1716
rect 414 -1810 418 -1716
rect 438 -1810 442 -1716
rect 462 -1810 466 -1716
rect 486 -1810 490 -1716
rect 510 -1810 514 -1716
rect 534 -1741 538 -1716
rect 534 -1765 541 -1741
rect 534 -1810 538 -1765
rect 558 -1810 562 -1716
rect 582 -1810 586 -1716
rect 606 -1810 610 -1716
rect 613 -1717 627 -1716
rect 619 -1723 624 -1717
rect 629 -1737 634 -1723
rect 619 -1795 624 -1785
rect 630 -1795 634 -1737
rect 629 -1809 634 -1795
rect 643 -1799 651 -1795
rect 637 -1809 643 -1799
rect 619 -1810 651 -1809
rect -2393 -1812 651 -1810
rect -2371 -1834 -2366 -1812
rect -2348 -1834 -2343 -1812
rect -2325 -1834 -2320 -1812
rect -2072 -1814 -2036 -1813
rect -2072 -1820 -2054 -1814
rect -2309 -1828 -2301 -1820
rect -2317 -1834 -2309 -1828
rect -2092 -1829 -2062 -1824
rect -2000 -1833 -1992 -1812
rect -1938 -1813 -1906 -1812
rect -1920 -1814 -1906 -1813
rect -1806 -1820 -1680 -1814
rect -1854 -1829 -1806 -1824
rect -1655 -1828 -1647 -1820
rect -1982 -1833 -1966 -1832
rect -2000 -1834 -1966 -1833
rect -1846 -1834 -1806 -1831
rect -1663 -1834 -1655 -1828
rect -1642 -1834 -1637 -1812
rect -1619 -1834 -1614 -1812
rect -1530 -1834 -1526 -1812
rect -1506 -1834 -1502 -1812
rect -1482 -1834 -1478 -1812
rect -1458 -1834 -1454 -1812
rect -1434 -1834 -1430 -1812
rect -1410 -1834 -1406 -1812
rect -1386 -1813 -1382 -1812
rect -2393 -1836 -1389 -1834
rect -2371 -1858 -2366 -1836
rect -2348 -1858 -2343 -1836
rect -2325 -1858 -2320 -1836
rect -2000 -1838 -1966 -1836
rect -2309 -1856 -2301 -1848
rect -2062 -1849 -2054 -1842
rect -2092 -1856 -2084 -1849
rect -2062 -1856 -2026 -1854
rect -2317 -1858 -2309 -1856
rect -2062 -1858 -2012 -1856
rect -2000 -1858 -1992 -1838
rect -1982 -1839 -1966 -1838
rect -1846 -1840 -1806 -1836
rect -1846 -1847 -1798 -1842
rect -1806 -1849 -1798 -1847
rect -1854 -1851 -1846 -1849
rect -1854 -1856 -1806 -1851
rect -1655 -1856 -1647 -1848
rect -1864 -1858 -1796 -1857
rect -1663 -1858 -1655 -1856
rect -1642 -1858 -1637 -1836
rect -1619 -1858 -1614 -1836
rect -1530 -1858 -1526 -1836
rect -1506 -1858 -1502 -1836
rect -1482 -1858 -1478 -1836
rect -1458 -1858 -1454 -1836
rect -1434 -1858 -1430 -1836
rect -1410 -1858 -1406 -1836
rect -1403 -1837 -1389 -1836
rect -1386 -1858 -1379 -1813
rect -1362 -1858 -1358 -1812
rect -1338 -1858 -1334 -1812
rect -1314 -1858 -1310 -1812
rect -1290 -1858 -1286 -1812
rect -1266 -1858 -1262 -1812
rect -1242 -1858 -1238 -1812
rect -1218 -1858 -1214 -1812
rect -1194 -1858 -1190 -1812
rect -1170 -1858 -1166 -1812
rect -1146 -1858 -1142 -1812
rect -1122 -1858 -1118 -1812
rect -1098 -1858 -1094 -1812
rect -1074 -1858 -1070 -1812
rect -1050 -1858 -1046 -1812
rect -1026 -1858 -1022 -1812
rect -1002 -1858 -998 -1812
rect -978 -1858 -974 -1812
rect -954 -1858 -950 -1812
rect -930 -1858 -926 -1812
rect -906 -1858 -902 -1812
rect -882 -1858 -878 -1812
rect -858 -1858 -854 -1812
rect -834 -1858 -830 -1812
rect -810 -1858 -806 -1812
rect -786 -1858 -782 -1812
rect -762 -1858 -758 -1812
rect -738 -1858 -734 -1812
rect -714 -1858 -710 -1812
rect -690 -1858 -686 -1812
rect -666 -1858 -662 -1812
rect -642 -1858 -638 -1812
rect -618 -1858 -614 -1812
rect -594 -1858 -590 -1812
rect -570 -1837 -566 -1812
rect -2393 -1860 -573 -1858
rect -2371 -1906 -2366 -1860
rect -2348 -1906 -2343 -1860
rect -2325 -1906 -2320 -1860
rect -2317 -1864 -2309 -1860
rect -2062 -1864 -2054 -1860
rect -2154 -1868 -2138 -1866
rect -2057 -1868 -2054 -1864
rect -2292 -1874 -2054 -1868
rect -2052 -1874 -2044 -1864
rect -2092 -1890 -2062 -1888
rect -2094 -1894 -2062 -1890
rect -2000 -1906 -1992 -1860
rect -1846 -1867 -1806 -1860
rect -1663 -1864 -1655 -1860
rect -1846 -1874 -1680 -1868
rect -1854 -1890 -1806 -1888
rect -1854 -1894 -1680 -1890
rect -1642 -1906 -1637 -1860
rect -1619 -1906 -1614 -1860
rect -1530 -1906 -1526 -1860
rect -1506 -1906 -1502 -1860
rect -1482 -1906 -1478 -1860
rect -1458 -1906 -1454 -1860
rect -1434 -1906 -1430 -1860
rect -1410 -1906 -1406 -1860
rect -1403 -1861 -1389 -1860
rect -1386 -1861 -1379 -1860
rect -1386 -1906 -1382 -1861
rect -1362 -1906 -1358 -1860
rect -1338 -1906 -1334 -1860
rect -1314 -1906 -1310 -1860
rect -1290 -1906 -1286 -1860
rect -1266 -1906 -1262 -1860
rect -1242 -1906 -1238 -1860
rect -1218 -1906 -1214 -1860
rect -1194 -1906 -1190 -1860
rect -1170 -1906 -1166 -1860
rect -1146 -1906 -1142 -1860
rect -1122 -1906 -1118 -1860
rect -1098 -1906 -1094 -1860
rect -1074 -1906 -1070 -1860
rect -1050 -1906 -1046 -1860
rect -1026 -1906 -1022 -1860
rect -1002 -1906 -998 -1860
rect -978 -1906 -974 -1860
rect -954 -1906 -950 -1860
rect -930 -1906 -926 -1860
rect -906 -1906 -902 -1860
rect -882 -1906 -878 -1860
rect -858 -1906 -854 -1860
rect -834 -1906 -830 -1860
rect -810 -1906 -806 -1860
rect -786 -1906 -782 -1860
rect -762 -1906 -758 -1860
rect -738 -1906 -734 -1860
rect -714 -1906 -710 -1860
rect -690 -1906 -686 -1860
rect -666 -1906 -662 -1860
rect -642 -1906 -638 -1860
rect -618 -1906 -614 -1860
rect -594 -1906 -590 -1860
rect -587 -1861 -573 -1860
rect -570 -1885 -563 -1837
rect -570 -1906 -566 -1885
rect -546 -1906 -542 -1812
rect -522 -1906 -518 -1812
rect -498 -1906 -494 -1812
rect -474 -1906 -470 -1812
rect -450 -1906 -446 -1812
rect -426 -1906 -422 -1812
rect -402 -1906 -398 -1812
rect -378 -1906 -374 -1812
rect -354 -1906 -350 -1812
rect -330 -1906 -326 -1812
rect -306 -1906 -302 -1812
rect -282 -1906 -278 -1812
rect -258 -1906 -254 -1812
rect -234 -1906 -230 -1812
rect -210 -1906 -206 -1812
rect -186 -1906 -182 -1812
rect -162 -1906 -158 -1812
rect -138 -1906 -134 -1812
rect -114 -1906 -110 -1812
rect -90 -1906 -86 -1812
rect -66 -1906 -62 -1812
rect -42 -1906 -38 -1812
rect -18 -1906 -14 -1812
rect 6 -1906 10 -1812
rect 30 -1906 34 -1812
rect 54 -1906 58 -1812
rect 78 -1906 82 -1812
rect 102 -1906 106 -1812
rect 126 -1906 130 -1812
rect 150 -1906 154 -1812
rect 174 -1906 178 -1812
rect 198 -1906 202 -1812
rect 222 -1906 226 -1812
rect 246 -1906 250 -1812
rect 270 -1906 274 -1812
rect 294 -1906 298 -1812
rect 318 -1906 322 -1812
rect 342 -1906 346 -1812
rect 366 -1906 370 -1812
rect 390 -1906 394 -1812
rect 403 -1843 408 -1833
rect 414 -1843 418 -1812
rect 413 -1857 418 -1843
rect 414 -1906 418 -1857
rect 438 -1906 442 -1812
rect 462 -1906 466 -1812
rect 486 -1906 490 -1812
rect 499 -1867 504 -1857
rect 510 -1867 514 -1812
rect 509 -1881 514 -1867
rect 510 -1906 514 -1881
rect 534 -1906 538 -1812
rect 558 -1906 562 -1812
rect 582 -1906 586 -1812
rect 606 -1906 610 -1812
rect 619 -1819 624 -1812
rect 637 -1813 651 -1812
rect 629 -1833 634 -1819
rect 630 -1906 634 -1833
rect 643 -1906 651 -1905
rect -2393 -1908 651 -1906
rect -2371 -1930 -2366 -1908
rect -2348 -1930 -2343 -1908
rect -2325 -1930 -2320 -1908
rect -2072 -1910 -2036 -1909
rect -2072 -1916 -2054 -1910
rect -2309 -1924 -2301 -1916
rect -2317 -1930 -2309 -1924
rect -2092 -1925 -2062 -1920
rect -2000 -1929 -1992 -1908
rect -1938 -1909 -1906 -1908
rect -1920 -1910 -1906 -1909
rect -1806 -1916 -1680 -1910
rect -1854 -1925 -1806 -1920
rect -1655 -1924 -1647 -1916
rect -1982 -1929 -1966 -1928
rect -2000 -1930 -1966 -1929
rect -1846 -1930 -1806 -1927
rect -1663 -1930 -1655 -1924
rect -1642 -1930 -1637 -1908
rect -1619 -1930 -1614 -1908
rect -1530 -1930 -1526 -1908
rect -1506 -1930 -1502 -1908
rect -1482 -1930 -1478 -1908
rect -1458 -1930 -1454 -1908
rect -1434 -1930 -1430 -1908
rect -1410 -1930 -1406 -1908
rect -1386 -1930 -1382 -1908
rect -1362 -1930 -1358 -1908
rect -1338 -1930 -1334 -1908
rect -1314 -1930 -1310 -1908
rect -1290 -1930 -1286 -1908
rect -1266 -1930 -1262 -1908
rect -1242 -1930 -1238 -1908
rect -1218 -1930 -1214 -1908
rect -1194 -1930 -1190 -1908
rect -1170 -1930 -1166 -1908
rect -1146 -1930 -1142 -1908
rect -1122 -1930 -1118 -1908
rect -1098 -1930 -1094 -1908
rect -1074 -1930 -1070 -1908
rect -1050 -1930 -1046 -1908
rect -1026 -1930 -1022 -1908
rect -1002 -1930 -998 -1908
rect -978 -1930 -974 -1908
rect -954 -1930 -950 -1908
rect -930 -1930 -926 -1908
rect -906 -1930 -902 -1908
rect -882 -1930 -878 -1908
rect -858 -1930 -854 -1908
rect -834 -1930 -830 -1908
rect -810 -1930 -806 -1908
rect -786 -1930 -782 -1908
rect -762 -1930 -758 -1908
rect -738 -1929 -734 -1908
rect -749 -1930 -715 -1929
rect -2393 -1932 -715 -1930
rect -2371 -1954 -2366 -1932
rect -2348 -1954 -2343 -1932
rect -2325 -1954 -2320 -1932
rect -2000 -1934 -1966 -1932
rect -2309 -1952 -2301 -1944
rect -2062 -1945 -2054 -1938
rect -2092 -1952 -2084 -1945
rect -2062 -1952 -2026 -1950
rect -2317 -1954 -2309 -1952
rect -2062 -1954 -2012 -1952
rect -2000 -1954 -1992 -1934
rect -1982 -1935 -1966 -1934
rect -1846 -1936 -1806 -1932
rect -1846 -1943 -1798 -1938
rect -1806 -1945 -1798 -1943
rect -1854 -1947 -1846 -1945
rect -1854 -1952 -1806 -1947
rect -1655 -1952 -1647 -1944
rect -1864 -1954 -1796 -1953
rect -1663 -1954 -1655 -1952
rect -1642 -1954 -1637 -1932
rect -1619 -1954 -1614 -1932
rect -1530 -1954 -1526 -1932
rect -1506 -1954 -1502 -1932
rect -1482 -1954 -1478 -1932
rect -1458 -1954 -1454 -1932
rect -1434 -1954 -1430 -1932
rect -1410 -1954 -1406 -1932
rect -1386 -1954 -1382 -1932
rect -1362 -1954 -1358 -1932
rect -1338 -1954 -1334 -1932
rect -1314 -1954 -1310 -1932
rect -1290 -1954 -1286 -1932
rect -1266 -1954 -1262 -1932
rect -1242 -1954 -1238 -1932
rect -1218 -1954 -1214 -1932
rect -1194 -1954 -1190 -1932
rect -1170 -1954 -1166 -1932
rect -1146 -1954 -1142 -1932
rect -1122 -1954 -1118 -1932
rect -1098 -1954 -1094 -1932
rect -1074 -1954 -1070 -1932
rect -1050 -1954 -1046 -1932
rect -1026 -1954 -1022 -1932
rect -1002 -1954 -998 -1932
rect -978 -1954 -974 -1932
rect -954 -1954 -950 -1932
rect -930 -1954 -926 -1932
rect -906 -1954 -902 -1932
rect -882 -1954 -878 -1932
rect -858 -1954 -854 -1932
rect -834 -1954 -830 -1932
rect -810 -1954 -806 -1932
rect -786 -1954 -782 -1932
rect -762 -1954 -758 -1932
rect -749 -1939 -744 -1932
rect -738 -1939 -734 -1932
rect -739 -1953 -734 -1939
rect -738 -1954 -734 -1953
rect -714 -1954 -710 -1908
rect -690 -1954 -686 -1908
rect -666 -1954 -662 -1908
rect -642 -1954 -638 -1908
rect -618 -1954 -614 -1908
rect -594 -1954 -590 -1908
rect -570 -1954 -566 -1908
rect -546 -1954 -542 -1908
rect -522 -1954 -518 -1908
rect -498 -1954 -494 -1908
rect -474 -1954 -470 -1908
rect -450 -1954 -446 -1908
rect -426 -1954 -422 -1908
rect -402 -1954 -398 -1908
rect -378 -1954 -374 -1908
rect -354 -1954 -350 -1908
rect -330 -1954 -326 -1908
rect -306 -1954 -302 -1908
rect -282 -1954 -278 -1908
rect -258 -1954 -254 -1908
rect -234 -1954 -230 -1908
rect -210 -1954 -206 -1908
rect -186 -1954 -182 -1908
rect -162 -1954 -158 -1908
rect -138 -1954 -134 -1908
rect -114 -1954 -110 -1908
rect -90 -1954 -86 -1908
rect -66 -1954 -62 -1908
rect -42 -1954 -38 -1908
rect -18 -1954 -14 -1908
rect 6 -1954 10 -1908
rect 30 -1954 34 -1908
rect 54 -1954 58 -1908
rect 78 -1954 82 -1908
rect 102 -1954 106 -1908
rect 126 -1954 130 -1908
rect 150 -1954 154 -1908
rect 174 -1954 178 -1908
rect 198 -1954 202 -1908
rect 222 -1954 226 -1908
rect 246 -1954 250 -1908
rect 270 -1954 274 -1908
rect 294 -1954 298 -1908
rect 318 -1954 322 -1908
rect 342 -1954 346 -1908
rect 366 -1954 370 -1908
rect 390 -1954 394 -1908
rect 414 -1954 418 -1908
rect 438 -1909 442 -1908
rect 438 -1933 445 -1909
rect 438 -1954 442 -1933
rect 462 -1954 466 -1908
rect 486 -1954 490 -1908
rect 510 -1953 514 -1908
rect 534 -1933 538 -1908
rect 499 -1954 531 -1953
rect -2393 -1956 531 -1954
rect -2371 -2002 -2366 -1956
rect -2348 -2002 -2343 -1956
rect -2325 -2002 -2320 -1956
rect -2317 -1960 -2309 -1956
rect -2062 -1960 -2054 -1956
rect -2154 -1964 -2138 -1962
rect -2057 -1964 -2054 -1960
rect -2292 -1970 -2054 -1964
rect -2052 -1970 -2044 -1960
rect -2092 -1986 -2062 -1984
rect -2094 -1990 -2062 -1986
rect -2000 -2002 -1992 -1956
rect -1846 -1963 -1806 -1956
rect -1663 -1960 -1655 -1956
rect -1846 -1970 -1680 -1964
rect -1854 -1986 -1806 -1984
rect -1854 -1990 -1680 -1986
rect -1642 -2002 -1637 -1956
rect -1619 -2002 -1614 -1956
rect -1530 -2002 -1526 -1956
rect -1506 -2002 -1502 -1956
rect -1482 -2002 -1478 -1956
rect -1458 -2002 -1454 -1956
rect -1434 -2002 -1430 -1956
rect -1410 -2002 -1406 -1956
rect -1386 -2002 -1382 -1956
rect -1362 -2002 -1358 -1956
rect -1338 -2002 -1334 -1956
rect -1314 -2002 -1310 -1956
rect -1290 -2002 -1286 -1956
rect -1266 -2002 -1262 -1956
rect -1242 -2002 -1238 -1956
rect -1218 -2002 -1214 -1956
rect -1194 -2002 -1190 -1956
rect -1170 -2002 -1166 -1956
rect -1146 -2002 -1142 -1956
rect -1122 -2002 -1118 -1956
rect -1098 -2002 -1094 -1956
rect -1074 -2002 -1070 -1956
rect -1050 -2002 -1046 -1956
rect -1026 -2002 -1022 -1956
rect -1002 -2002 -998 -1956
rect -978 -2002 -974 -1956
rect -954 -2002 -950 -1956
rect -930 -2002 -926 -1956
rect -906 -2002 -902 -1956
rect -882 -2002 -878 -1956
rect -858 -2002 -854 -1956
rect -834 -2002 -830 -1956
rect -810 -2002 -806 -1956
rect -786 -2002 -782 -1956
rect -762 -2002 -758 -1956
rect -738 -2002 -734 -1956
rect -714 -2002 -710 -1956
rect -690 -2002 -686 -1956
rect -666 -2002 -662 -1956
rect -642 -2002 -638 -1956
rect -618 -2002 -614 -1956
rect -594 -2002 -590 -1956
rect -570 -2002 -566 -1956
rect -546 -2002 -542 -1956
rect -522 -2002 -518 -1956
rect -498 -2002 -494 -1956
rect -474 -2002 -470 -1956
rect -450 -2002 -446 -1956
rect -426 -2002 -422 -1956
rect -402 -2002 -398 -1956
rect -378 -2002 -374 -1956
rect -354 -2002 -350 -1956
rect -330 -2002 -326 -1956
rect -306 -2002 -302 -1956
rect -282 -2002 -278 -1956
rect -258 -2002 -254 -1956
rect -234 -2002 -230 -1956
rect -210 -2002 -206 -1956
rect -186 -2002 -182 -1956
rect -162 -2002 -158 -1956
rect -138 -2002 -134 -1956
rect -114 -2002 -110 -1956
rect -90 -2002 -86 -1956
rect -66 -2002 -62 -1956
rect -42 -2002 -38 -1956
rect -18 -2002 -14 -1956
rect 6 -2002 10 -1956
rect 30 -2002 34 -1956
rect 54 -2002 58 -1956
rect 78 -2002 82 -1956
rect 102 -2002 106 -1956
rect 126 -2002 130 -1956
rect 150 -2002 154 -1956
rect 174 -2002 178 -1956
rect 198 -2002 202 -1956
rect 222 -2002 226 -1956
rect 246 -2002 250 -1956
rect 270 -2002 274 -1956
rect 294 -2002 298 -1956
rect 318 -2002 322 -1956
rect 342 -2002 346 -1956
rect 366 -2002 370 -1956
rect 390 -2002 394 -1956
rect 414 -2002 418 -1956
rect 438 -2002 442 -1956
rect 462 -2002 466 -1956
rect 486 -2002 490 -1956
rect 499 -1963 504 -1956
rect 510 -1963 514 -1956
rect 517 -1957 531 -1956
rect 534 -1957 541 -1933
rect 509 -1977 514 -1963
rect 499 -1987 504 -1977
rect 509 -2001 514 -1987
rect 510 -2002 514 -2001
rect 534 -2002 538 -1957
rect 558 -2002 562 -1908
rect 582 -2002 586 -1908
rect 606 -2002 610 -1908
rect 630 -2002 634 -1908
rect 637 -1909 651 -1908
rect 643 -1915 648 -1909
rect 653 -1929 658 -1915
rect 643 -1987 648 -1977
rect 654 -1987 658 -1929
rect 653 -2001 658 -1987
rect 667 -1991 675 -1987
rect 661 -2001 667 -1991
rect 643 -2002 675 -2001
rect -2393 -2004 675 -2002
rect -2371 -2026 -2366 -2004
rect -2348 -2026 -2343 -2004
rect -2325 -2026 -2320 -2004
rect -2072 -2006 -2036 -2005
rect -2072 -2012 -2054 -2006
rect -2309 -2020 -2301 -2012
rect -2317 -2026 -2309 -2020
rect -2092 -2021 -2062 -2016
rect -2000 -2025 -1992 -2004
rect -1938 -2005 -1906 -2004
rect -1920 -2006 -1906 -2005
rect -1806 -2012 -1680 -2006
rect -1854 -2021 -1806 -2016
rect -1655 -2020 -1647 -2012
rect -1982 -2025 -1966 -2024
rect -2000 -2026 -1966 -2025
rect -1846 -2026 -1806 -2023
rect -1663 -2026 -1655 -2020
rect -1642 -2026 -1637 -2004
rect -1619 -2026 -1614 -2004
rect -1530 -2026 -1526 -2004
rect -1506 -2026 -1502 -2004
rect -1482 -2026 -1478 -2004
rect -1458 -2026 -1454 -2004
rect -1434 -2026 -1430 -2004
rect -1410 -2026 -1406 -2004
rect -1386 -2026 -1382 -2004
rect -1362 -2026 -1358 -2004
rect -1338 -2026 -1334 -2004
rect -1314 -2026 -1310 -2004
rect -1290 -2026 -1286 -2004
rect -1266 -2025 -1262 -2004
rect -1277 -2026 -1243 -2025
rect -2393 -2028 -1243 -2026
rect -2371 -2050 -2366 -2028
rect -2348 -2050 -2343 -2028
rect -2325 -2050 -2320 -2028
rect -2000 -2030 -1966 -2028
rect -2309 -2048 -2301 -2040
rect -2062 -2041 -2054 -2034
rect -2092 -2048 -2084 -2041
rect -2062 -2048 -2026 -2046
rect -2317 -2050 -2309 -2048
rect -2062 -2050 -2012 -2048
rect -2000 -2050 -1992 -2030
rect -1982 -2031 -1966 -2030
rect -1846 -2032 -1806 -2028
rect -1846 -2039 -1798 -2034
rect -1806 -2041 -1798 -2039
rect -1854 -2043 -1846 -2041
rect -1854 -2048 -1806 -2043
rect -1655 -2048 -1647 -2040
rect -1864 -2050 -1796 -2049
rect -1663 -2050 -1655 -2048
rect -1642 -2050 -1637 -2028
rect -1619 -2050 -1614 -2028
rect -1530 -2050 -1526 -2028
rect -1506 -2050 -1502 -2028
rect -1482 -2050 -1478 -2028
rect -1458 -2050 -1454 -2028
rect -1434 -2050 -1430 -2028
rect -1410 -2049 -1406 -2028
rect -1421 -2050 -1387 -2049
rect -2393 -2052 -1387 -2050
rect -2371 -2098 -2366 -2052
rect -2348 -2098 -2343 -2052
rect -2325 -2088 -2320 -2052
rect -2317 -2056 -2309 -2052
rect -2062 -2056 -2054 -2052
rect -2154 -2060 -2138 -2058
rect -2057 -2060 -2054 -2056
rect -2292 -2066 -2054 -2060
rect -2052 -2066 -2044 -2056
rect -2092 -2082 -2062 -2080
rect -2094 -2086 -2062 -2082
rect -2325 -2098 -2317 -2088
rect -2095 -2096 -2084 -2092
rect -2000 -2095 -1992 -2052
rect -1846 -2059 -1806 -2052
rect -1663 -2056 -1655 -2052
rect -1846 -2066 -1680 -2060
rect -1854 -2082 -1806 -2080
rect -1854 -2086 -1680 -2082
rect -2119 -2098 -2069 -2096
rect -2054 -2098 -1892 -2095
rect -1671 -2098 -1663 -2088
rect -1642 -2098 -1637 -2052
rect -1619 -2098 -1614 -2052
rect -1530 -2098 -1526 -2052
rect -1506 -2098 -1502 -2052
rect -1482 -2098 -1478 -2052
rect -1458 -2098 -1454 -2052
rect -1434 -2098 -1430 -2052
rect -1421 -2059 -1416 -2052
rect -1410 -2059 -1406 -2052
rect -1411 -2073 -1406 -2059
rect -1421 -2083 -1416 -2073
rect -1411 -2097 -1406 -2083
rect -1410 -2098 -1406 -2097
rect -1386 -2098 -1382 -2028
rect -1362 -2098 -1358 -2028
rect -1338 -2098 -1334 -2028
rect -1314 -2098 -1310 -2028
rect -1290 -2098 -1286 -2028
rect -1277 -2035 -1272 -2028
rect -1266 -2035 -1262 -2028
rect -1267 -2049 -1262 -2035
rect -1277 -2050 -1243 -2049
rect -1242 -2050 -1238 -2004
rect -1218 -2050 -1214 -2004
rect -1194 -2050 -1190 -2004
rect -1170 -2050 -1166 -2004
rect -1146 -2050 -1142 -2004
rect -1122 -2050 -1118 -2004
rect -1098 -2050 -1094 -2004
rect -1074 -2050 -1070 -2004
rect -1050 -2050 -1046 -2004
rect -1026 -2050 -1022 -2004
rect -1002 -2050 -998 -2004
rect -978 -2050 -974 -2004
rect -954 -2050 -950 -2004
rect -930 -2050 -926 -2004
rect -906 -2050 -902 -2004
rect -882 -2050 -878 -2004
rect -858 -2050 -854 -2004
rect -834 -2050 -830 -2004
rect -810 -2050 -806 -2004
rect -786 -2050 -782 -2004
rect -762 -2050 -758 -2004
rect -738 -2050 -734 -2004
rect -714 -2005 -710 -2004
rect -714 -2029 -707 -2005
rect -714 -2050 -710 -2029
rect -690 -2050 -686 -2004
rect -666 -2050 -662 -2004
rect -642 -2050 -638 -2004
rect -618 -2050 -614 -2004
rect -594 -2050 -590 -2004
rect -570 -2050 -566 -2004
rect -546 -2050 -542 -2004
rect -522 -2050 -518 -2004
rect -498 -2050 -494 -2004
rect -474 -2050 -470 -2004
rect -450 -2050 -446 -2004
rect -426 -2050 -422 -2004
rect -402 -2050 -398 -2004
rect -378 -2050 -374 -2004
rect -354 -2050 -350 -2004
rect -330 -2050 -326 -2004
rect -306 -2050 -302 -2004
rect -282 -2050 -278 -2004
rect -258 -2050 -254 -2004
rect -234 -2050 -230 -2004
rect -210 -2050 -206 -2004
rect -186 -2050 -182 -2004
rect -162 -2050 -158 -2004
rect -138 -2050 -134 -2004
rect -114 -2050 -110 -2004
rect -90 -2050 -86 -2004
rect -66 -2050 -62 -2004
rect -42 -2050 -38 -2004
rect -18 -2050 -14 -2004
rect 6 -2050 10 -2004
rect 30 -2050 34 -2004
rect 54 -2050 58 -2004
rect 78 -2050 82 -2004
rect 102 -2050 106 -2004
rect 126 -2050 130 -2004
rect 150 -2050 154 -2004
rect 174 -2050 178 -2004
rect 198 -2050 202 -2004
rect 222 -2050 226 -2004
rect 246 -2050 250 -2004
rect 270 -2050 274 -2004
rect 294 -2050 298 -2004
rect 318 -2050 322 -2004
rect 342 -2050 346 -2004
rect 366 -2050 370 -2004
rect 390 -2050 394 -2004
rect 414 -2050 418 -2004
rect 438 -2050 442 -2004
rect 462 -2050 466 -2004
rect 486 -2050 490 -2004
rect 510 -2050 514 -2004
rect 534 -2029 538 -2004
rect -1277 -2052 531 -2050
rect -1277 -2059 -1272 -2052
rect -1267 -2073 -1262 -2059
rect -1266 -2098 -1262 -2073
rect -1242 -2098 -1238 -2052
rect -1218 -2098 -1214 -2052
rect -1194 -2098 -1190 -2052
rect -1170 -2098 -1166 -2052
rect -1146 -2098 -1142 -2052
rect -1122 -2098 -1118 -2052
rect -1098 -2098 -1094 -2052
rect -1074 -2098 -1070 -2052
rect -1050 -2098 -1046 -2052
rect -1026 -2098 -1022 -2052
rect -1002 -2098 -998 -2052
rect -978 -2098 -974 -2052
rect -954 -2098 -950 -2052
rect -930 -2098 -926 -2052
rect -906 -2098 -902 -2052
rect -882 -2098 -878 -2052
rect -858 -2098 -854 -2052
rect -834 -2098 -830 -2052
rect -810 -2098 -806 -2052
rect -786 -2098 -782 -2052
rect -762 -2098 -758 -2052
rect -738 -2098 -734 -2052
rect -714 -2098 -710 -2052
rect -690 -2098 -686 -2052
rect -666 -2098 -662 -2052
rect -642 -2098 -638 -2052
rect -618 -2098 -614 -2052
rect -594 -2098 -590 -2052
rect -570 -2098 -566 -2052
rect -546 -2098 -542 -2052
rect -522 -2098 -518 -2052
rect -498 -2098 -494 -2052
rect -474 -2098 -470 -2052
rect -450 -2098 -446 -2052
rect -426 -2098 -422 -2052
rect -402 -2098 -398 -2052
rect -378 -2098 -374 -2052
rect -354 -2098 -350 -2052
rect -330 -2098 -326 -2052
rect -306 -2098 -302 -2052
rect -282 -2098 -278 -2052
rect -258 -2098 -254 -2052
rect -234 -2098 -230 -2052
rect -210 -2098 -206 -2052
rect -186 -2098 -182 -2052
rect -162 -2098 -158 -2052
rect -138 -2098 -134 -2052
rect -114 -2098 -110 -2052
rect -90 -2098 -86 -2052
rect -66 -2098 -62 -2052
rect -42 -2098 -38 -2052
rect -18 -2098 -14 -2052
rect 6 -2098 10 -2052
rect 30 -2098 34 -2052
rect 54 -2098 58 -2052
rect 78 -2098 82 -2052
rect 102 -2098 106 -2052
rect 126 -2098 130 -2052
rect 150 -2098 154 -2052
rect 174 -2098 178 -2052
rect 198 -2098 202 -2052
rect 222 -2098 226 -2052
rect 246 -2098 250 -2052
rect 270 -2098 274 -2052
rect 294 -2098 298 -2052
rect 318 -2098 322 -2052
rect 342 -2098 346 -2052
rect 366 -2098 370 -2052
rect 390 -2098 394 -2052
rect 414 -2098 418 -2052
rect 438 -2098 442 -2052
rect 462 -2098 466 -2052
rect 486 -2098 490 -2052
rect 510 -2098 514 -2052
rect 517 -2053 531 -2052
rect 534 -2074 541 -2029
rect 558 -2074 562 -2004
rect 582 -2074 586 -2004
rect 606 -2074 610 -2004
rect 630 -2073 634 -2004
rect 643 -2011 648 -2004
rect 661 -2005 675 -2004
rect 653 -2025 658 -2011
rect 643 -2059 648 -2049
rect 654 -2059 658 -2025
rect 653 -2073 658 -2059
rect 667 -2063 675 -2059
rect 661 -2073 667 -2063
rect 619 -2074 653 -2073
rect 517 -2076 653 -2074
rect 517 -2077 531 -2076
rect 534 -2077 541 -2076
rect 534 -2098 538 -2077
rect 558 -2098 562 -2076
rect 582 -2098 586 -2076
rect 606 -2098 610 -2076
rect 619 -2083 624 -2076
rect 630 -2083 634 -2076
rect 629 -2097 634 -2083
rect 619 -2098 653 -2097
rect -2393 -2100 653 -2098
rect -2371 -2122 -2366 -2100
rect -2348 -2122 -2343 -2100
rect -2325 -2104 -2317 -2100
rect -2325 -2120 -2320 -2104
rect -2309 -2116 -2301 -2104
rect -2095 -2106 -2084 -2100
rect -2054 -2101 -1906 -2100
rect -2054 -2102 -2036 -2101
rect -2084 -2108 -2079 -2106
rect -2317 -2120 -2309 -2116
rect -2092 -2117 -2079 -2110
rect -2000 -2114 -1992 -2101
rect -1920 -2102 -1906 -2101
rect -1671 -2104 -1663 -2100
rect -1846 -2108 -1806 -2106
rect -1854 -2114 -1806 -2110
rect -2054 -2117 -1982 -2114
rect -1966 -2117 -1806 -2114
rect -1655 -2116 -1647 -2104
rect -2003 -2120 -1992 -2117
rect -1904 -2119 -1902 -2117
rect -1854 -2119 -1846 -2117
rect -2325 -2122 -2317 -2120
rect -2033 -2122 -1992 -2120
rect -1854 -2121 -1806 -2119
rect -1663 -2120 -1655 -2116
rect -1864 -2122 -1796 -2121
rect -1671 -2122 -1663 -2120
rect -1642 -2122 -1637 -2100
rect -1619 -2122 -1614 -2100
rect -1530 -2122 -1526 -2100
rect -1506 -2122 -1502 -2100
rect -1482 -2122 -1478 -2100
rect -1458 -2122 -1454 -2100
rect -1434 -2122 -1430 -2100
rect -1410 -2122 -1406 -2100
rect -1386 -2122 -1382 -2100
rect -1362 -2122 -1358 -2100
rect -1338 -2122 -1334 -2100
rect -1314 -2122 -1310 -2100
rect -1290 -2122 -1286 -2100
rect -1266 -2122 -1262 -2100
rect -1242 -2101 -1238 -2100
rect -2393 -2124 -1245 -2122
rect -2371 -2146 -2366 -2124
rect -2348 -2146 -2343 -2124
rect -2325 -2132 -2317 -2124
rect -2079 -2127 -2018 -2124
rect -2003 -2125 -1966 -2124
rect -2000 -2126 -1982 -2125
rect -2000 -2127 -1992 -2126
rect -2084 -2131 -2009 -2127
rect -2028 -2132 -2009 -2131
rect -2000 -2131 -1854 -2127
rect -1846 -2131 -1798 -2124
rect -2325 -2146 -2320 -2132
rect -2309 -2144 -2301 -2132
rect -2028 -2134 -2018 -2132
rect -2092 -2144 -2084 -2137
rect -2023 -2141 -2014 -2134
rect -2000 -2141 -1992 -2131
rect -1671 -2132 -1663 -2124
rect -1846 -2135 -1806 -2133
rect -1854 -2141 -1806 -2137
rect -2054 -2144 -1806 -2141
rect -1655 -2144 -1647 -2132
rect -2317 -2146 -2309 -2144
rect -2054 -2146 -2024 -2144
rect -2000 -2146 -1992 -2144
rect -1663 -2146 -1655 -2144
rect -1642 -2146 -1637 -2124
rect -1619 -2146 -1614 -2124
rect -1530 -2146 -1526 -2124
rect -1506 -2146 -1502 -2124
rect -1482 -2146 -1478 -2124
rect -1458 -2146 -1454 -2124
rect -1434 -2146 -1430 -2124
rect -1410 -2146 -1406 -2124
rect -1386 -2125 -1382 -2124
rect -2393 -2148 -2064 -2146
rect -2060 -2148 -1389 -2146
rect -2371 -2194 -2366 -2148
rect -2348 -2194 -2343 -2148
rect -2325 -2160 -2317 -2148
rect -2060 -2151 -2054 -2148
rect -2084 -2158 -2054 -2151
rect -2050 -2154 -2044 -2152
rect -2325 -2180 -2320 -2160
rect -2064 -2162 -2054 -2158
rect -2325 -2188 -2317 -2180
rect -2101 -2185 -2071 -2182
rect -2325 -2194 -2320 -2188
rect -2317 -2194 -2309 -2188
rect -2000 -2190 -1992 -2148
rect -1846 -2149 -1806 -2148
rect -1846 -2158 -1798 -2151
rect -1671 -2160 -1663 -2148
rect -1846 -2162 -1806 -2160
rect -1854 -2176 -1680 -2172
rect -1846 -2185 -1798 -2182
rect -2079 -2191 -2043 -2190
rect -2007 -2191 -1991 -2190
rect -2079 -2192 -2071 -2191
rect -2079 -2194 -2029 -2192
rect -2011 -2194 -1991 -2191
rect -1846 -2193 -1806 -2187
rect -1671 -2188 -1663 -2180
rect -1864 -2194 -1796 -2193
rect -1663 -2194 -1655 -2188
rect -1642 -2194 -1637 -2148
rect -1619 -2194 -1614 -2148
rect -1530 -2194 -1526 -2148
rect -1506 -2194 -1502 -2148
rect -1482 -2194 -1478 -2148
rect -1458 -2194 -1454 -2148
rect -1434 -2194 -1430 -2148
rect -1410 -2194 -1406 -2148
rect -1403 -2149 -1389 -2148
rect -1386 -2170 -1379 -2125
rect -1362 -2170 -1358 -2124
rect -1338 -2170 -1334 -2124
rect -1314 -2170 -1310 -2124
rect -1290 -2170 -1286 -2124
rect -1266 -2170 -1262 -2124
rect -1259 -2125 -1245 -2124
rect -1242 -2146 -1235 -2101
rect -1218 -2146 -1214 -2100
rect -1194 -2146 -1190 -2100
rect -1170 -2146 -1166 -2100
rect -1146 -2146 -1142 -2100
rect -1122 -2146 -1118 -2100
rect -1098 -2146 -1094 -2100
rect -1074 -2146 -1070 -2100
rect -1050 -2146 -1046 -2100
rect -1026 -2146 -1022 -2100
rect -1002 -2146 -998 -2100
rect -978 -2146 -974 -2100
rect -954 -2146 -950 -2100
rect -930 -2146 -926 -2100
rect -906 -2146 -902 -2100
rect -882 -2146 -878 -2100
rect -869 -2131 -864 -2121
rect -858 -2131 -854 -2100
rect -859 -2145 -854 -2131
rect -834 -2146 -830 -2100
rect -810 -2146 -806 -2100
rect -786 -2146 -782 -2100
rect -762 -2146 -758 -2100
rect -738 -2146 -734 -2100
rect -714 -2146 -710 -2100
rect -690 -2146 -686 -2100
rect -666 -2146 -662 -2100
rect -642 -2146 -638 -2100
rect -618 -2146 -614 -2100
rect -594 -2146 -590 -2100
rect -570 -2146 -566 -2100
rect -546 -2146 -542 -2100
rect -522 -2146 -518 -2100
rect -498 -2146 -494 -2100
rect -474 -2146 -470 -2100
rect -450 -2146 -446 -2100
rect -426 -2146 -422 -2100
rect -402 -2146 -398 -2100
rect -378 -2146 -374 -2100
rect -354 -2146 -350 -2100
rect -330 -2146 -326 -2100
rect -306 -2146 -302 -2100
rect -282 -2146 -278 -2100
rect -258 -2146 -254 -2100
rect -234 -2146 -230 -2100
rect -210 -2146 -206 -2100
rect -186 -2146 -182 -2100
rect -162 -2146 -158 -2100
rect -138 -2146 -134 -2100
rect -114 -2146 -110 -2100
rect -90 -2146 -86 -2100
rect -66 -2146 -62 -2100
rect -42 -2146 -38 -2100
rect -18 -2146 -14 -2100
rect 6 -2146 10 -2100
rect 30 -2146 34 -2100
rect 54 -2146 58 -2100
rect 78 -2146 82 -2100
rect 102 -2146 106 -2100
rect 126 -2146 130 -2100
rect 150 -2146 154 -2100
rect 174 -2146 178 -2100
rect 198 -2146 202 -2100
rect 222 -2146 226 -2100
rect 246 -2146 250 -2100
rect 270 -2146 274 -2100
rect 294 -2146 298 -2100
rect 318 -2146 322 -2100
rect 342 -2146 346 -2100
rect 366 -2146 370 -2100
rect 390 -2146 394 -2100
rect 414 -2146 418 -2100
rect 438 -2145 442 -2100
rect 427 -2146 461 -2145
rect -1259 -2148 461 -2146
rect -1259 -2149 -1245 -2148
rect -1242 -2149 -1235 -2148
rect -1242 -2170 -1238 -2149
rect -1218 -2170 -1214 -2148
rect -1194 -2170 -1190 -2148
rect -1170 -2170 -1166 -2148
rect -1146 -2170 -1142 -2148
rect -1122 -2170 -1118 -2148
rect -1098 -2170 -1094 -2148
rect -1074 -2170 -1070 -2148
rect -1050 -2170 -1046 -2148
rect -1026 -2170 -1022 -2148
rect -1002 -2170 -998 -2148
rect -978 -2170 -974 -2148
rect -954 -2170 -950 -2148
rect -930 -2170 -926 -2148
rect -906 -2170 -902 -2148
rect -882 -2170 -878 -2148
rect -834 -2170 -830 -2148
rect -810 -2170 -806 -2148
rect -786 -2170 -782 -2148
rect -762 -2170 -758 -2148
rect -738 -2170 -734 -2148
rect -714 -2170 -710 -2148
rect -690 -2170 -686 -2148
rect -666 -2170 -662 -2148
rect -642 -2170 -638 -2148
rect -618 -2170 -614 -2148
rect -594 -2170 -590 -2148
rect -570 -2170 -566 -2148
rect -546 -2170 -542 -2148
rect -522 -2170 -518 -2148
rect -498 -2170 -494 -2148
rect -474 -2170 -470 -2148
rect -450 -2170 -446 -2148
rect -426 -2170 -422 -2148
rect -402 -2170 -398 -2148
rect -378 -2170 -374 -2148
rect -354 -2170 -350 -2148
rect -330 -2170 -326 -2148
rect -306 -2170 -302 -2148
rect -282 -2170 -278 -2148
rect -258 -2170 -254 -2148
rect -234 -2170 -230 -2148
rect -210 -2170 -206 -2148
rect -186 -2170 -182 -2148
rect -162 -2170 -158 -2148
rect -138 -2170 -134 -2148
rect -114 -2170 -110 -2148
rect -90 -2170 -86 -2148
rect -66 -2170 -62 -2148
rect -42 -2170 -38 -2148
rect -18 -2170 -14 -2148
rect 6 -2170 10 -2148
rect 30 -2170 34 -2148
rect 54 -2170 58 -2148
rect 78 -2170 82 -2148
rect 102 -2170 106 -2148
rect 126 -2170 130 -2148
rect 150 -2170 154 -2148
rect 174 -2170 178 -2148
rect 198 -2170 202 -2148
rect 222 -2170 226 -2148
rect 246 -2170 250 -2148
rect 270 -2169 274 -2148
rect 259 -2170 293 -2169
rect -1403 -2172 293 -2170
rect -1403 -2173 -1389 -2172
rect -1386 -2173 -1379 -2172
rect -1386 -2194 -1382 -2173
rect -1362 -2194 -1358 -2172
rect -1338 -2194 -1334 -2172
rect -1314 -2194 -1310 -2172
rect -1290 -2194 -1286 -2172
rect -1266 -2194 -1262 -2172
rect -1242 -2194 -1238 -2172
rect -1218 -2194 -1214 -2172
rect -1194 -2194 -1190 -2172
rect -1170 -2194 -1166 -2172
rect -1146 -2194 -1142 -2172
rect -1122 -2194 -1118 -2172
rect -1098 -2194 -1094 -2172
rect -1074 -2194 -1070 -2172
rect -1050 -2194 -1046 -2172
rect -1026 -2194 -1022 -2172
rect -1002 -2194 -998 -2172
rect -978 -2194 -974 -2172
rect -954 -2194 -950 -2172
rect -930 -2194 -926 -2172
rect -906 -2194 -902 -2172
rect -882 -2194 -878 -2172
rect -834 -2194 -830 -2172
rect -810 -2194 -806 -2172
rect -786 -2194 -782 -2172
rect -762 -2194 -758 -2172
rect -738 -2194 -734 -2172
rect -714 -2193 -710 -2172
rect -725 -2194 -691 -2193
rect -2393 -2196 -691 -2194
rect -2371 -2242 -2366 -2196
rect -2348 -2242 -2343 -2196
rect -2325 -2208 -2320 -2196
rect -2079 -2198 -2071 -2196
rect -2072 -2200 -2071 -2198
rect -2109 -2205 -2101 -2200
rect -2101 -2207 -2079 -2205
rect -2069 -2207 -2068 -2200
rect -2325 -2216 -2317 -2208
rect -2079 -2212 -2071 -2207
rect -2325 -2236 -2320 -2216
rect -2317 -2224 -2309 -2216
rect -2074 -2221 -2071 -2212
rect -2069 -2216 -2068 -2212
rect -2109 -2230 -2079 -2227
rect -2325 -2242 -2317 -2236
rect -2000 -2242 -1992 -2196
rect -1846 -2198 -1806 -2196
rect -1854 -2203 -1806 -2199
rect -1854 -2205 -1846 -2203
rect -1846 -2207 -1806 -2205
rect -1806 -2209 -1798 -2207
rect -1846 -2212 -1798 -2209
rect -1846 -2225 -1806 -2214
rect -1671 -2216 -1663 -2208
rect -1663 -2224 -1655 -2216
rect -1854 -2230 -1680 -2226
rect -1671 -2242 -1663 -2236
rect -1642 -2242 -1637 -2196
rect -1619 -2242 -1614 -2196
rect -1530 -2242 -1526 -2196
rect -1506 -2242 -1502 -2196
rect -1482 -2242 -1478 -2196
rect -1458 -2242 -1454 -2196
rect -1434 -2242 -1430 -2196
rect -1410 -2242 -1406 -2196
rect -1386 -2242 -1382 -2196
rect -1362 -2242 -1358 -2196
rect -1338 -2242 -1334 -2196
rect -1314 -2242 -1310 -2196
rect -1290 -2242 -1286 -2196
rect -1266 -2242 -1262 -2196
rect -1242 -2242 -1238 -2196
rect -1218 -2242 -1214 -2196
rect -1194 -2242 -1190 -2196
rect -1170 -2242 -1166 -2196
rect -1146 -2242 -1142 -2196
rect -1122 -2242 -1118 -2196
rect -1098 -2242 -1094 -2196
rect -1074 -2242 -1070 -2196
rect -1050 -2242 -1046 -2196
rect -1026 -2242 -1022 -2196
rect -1002 -2242 -998 -2196
rect -978 -2242 -974 -2196
rect -954 -2242 -950 -2196
rect -930 -2242 -926 -2196
rect -906 -2242 -902 -2196
rect -882 -2242 -878 -2196
rect -834 -2197 -830 -2196
rect -869 -2220 -837 -2217
rect -869 -2227 -864 -2220
rect -851 -2221 -837 -2220
rect -834 -2221 -827 -2197
rect -859 -2241 -854 -2227
rect -858 -2242 -854 -2241
rect -810 -2242 -806 -2196
rect -786 -2242 -782 -2196
rect -762 -2242 -758 -2196
rect -738 -2242 -734 -2196
rect -725 -2203 -720 -2196
rect -714 -2203 -710 -2196
rect -715 -2217 -710 -2203
rect -725 -2242 -691 -2241
rect -2393 -2244 -691 -2242
rect -2371 -2266 -2366 -2244
rect -2348 -2266 -2343 -2244
rect -2325 -2252 -2317 -2244
rect -2325 -2266 -2320 -2252
rect -2309 -2264 -2301 -2252
rect -2092 -2261 -2062 -2256
rect -2000 -2264 -1992 -2244
rect -2317 -2266 -2309 -2264
rect -2000 -2266 -1983 -2264
rect -1906 -2266 -1904 -2244
rect -1806 -2252 -1680 -2246
rect -1671 -2252 -1663 -2244
rect -1854 -2261 -1806 -2256
rect -1846 -2266 -1806 -2263
rect -1655 -2264 -1647 -2252
rect -1663 -2266 -1655 -2264
rect -1642 -2266 -1637 -2244
rect -1619 -2266 -1614 -2244
rect -1530 -2266 -1526 -2244
rect -1506 -2266 -1502 -2244
rect -1482 -2266 -1478 -2244
rect -1458 -2266 -1454 -2244
rect -1434 -2266 -1430 -2244
rect -1410 -2266 -1406 -2244
rect -1386 -2266 -1382 -2244
rect -1362 -2266 -1358 -2244
rect -1338 -2266 -1334 -2244
rect -1314 -2266 -1310 -2244
rect -1290 -2266 -1286 -2244
rect -1266 -2266 -1262 -2244
rect -1242 -2266 -1238 -2244
rect -1218 -2266 -1214 -2244
rect -1194 -2266 -1190 -2244
rect -1170 -2266 -1166 -2244
rect -1146 -2266 -1142 -2244
rect -1122 -2266 -1118 -2244
rect -1098 -2266 -1094 -2244
rect -1074 -2266 -1070 -2244
rect -1050 -2266 -1046 -2244
rect -1026 -2266 -1022 -2244
rect -1002 -2266 -998 -2244
rect -978 -2266 -974 -2244
rect -954 -2266 -950 -2244
rect -930 -2266 -926 -2244
rect -906 -2266 -902 -2244
rect -882 -2266 -878 -2244
rect -858 -2266 -854 -2244
rect -810 -2266 -806 -2244
rect -786 -2265 -782 -2244
rect -797 -2266 -763 -2265
rect -2393 -2268 -763 -2266
rect -2371 -2290 -2366 -2268
rect -2348 -2290 -2343 -2268
rect -2325 -2280 -2317 -2268
rect -2071 -2272 -2062 -2268
rect -2013 -2270 -1983 -2268
rect -2000 -2271 -1983 -2270
rect -2325 -2290 -2320 -2280
rect -2309 -2290 -2301 -2280
rect -2100 -2281 -2092 -2274
rect -2064 -2276 -2062 -2273
rect -2061 -2281 -2059 -2276
rect -2071 -2286 -2062 -2281
rect -2071 -2288 -2026 -2286
rect -2066 -2290 -2012 -2288
rect -2000 -2290 -1992 -2271
rect -1906 -2273 -1904 -2268
rect -1846 -2272 -1806 -2268
rect -1846 -2279 -1798 -2274
rect -1806 -2281 -1798 -2279
rect -1671 -2280 -1663 -2268
rect -1854 -2283 -1846 -2281
rect -1854 -2288 -1806 -2283
rect -1864 -2290 -1796 -2289
rect -1655 -2290 -1647 -2280
rect -1642 -2290 -1637 -2268
rect -1619 -2290 -1614 -2268
rect -1530 -2290 -1526 -2268
rect -1506 -2290 -1502 -2268
rect -1482 -2290 -1478 -2268
rect -1458 -2290 -1454 -2268
rect -1434 -2290 -1430 -2268
rect -1410 -2290 -1406 -2268
rect -1386 -2290 -1382 -2268
rect -1362 -2290 -1358 -2268
rect -1338 -2290 -1334 -2268
rect -1314 -2290 -1310 -2268
rect -1290 -2290 -1286 -2268
rect -1266 -2290 -1262 -2268
rect -1242 -2290 -1238 -2268
rect -1218 -2290 -1214 -2268
rect -1194 -2290 -1190 -2268
rect -1170 -2290 -1166 -2268
rect -1146 -2290 -1142 -2268
rect -1122 -2290 -1118 -2268
rect -1098 -2290 -1094 -2268
rect -1074 -2290 -1070 -2268
rect -1050 -2290 -1046 -2268
rect -1026 -2290 -1022 -2268
rect -1002 -2290 -998 -2268
rect -978 -2289 -974 -2268
rect -989 -2290 -955 -2289
rect -2393 -2292 -955 -2290
rect -2371 -2338 -2366 -2292
rect -2348 -2338 -2343 -2292
rect -2325 -2296 -2320 -2292
rect -2317 -2296 -2309 -2292
rect -2325 -2308 -2317 -2296
rect -2066 -2297 -2062 -2292
rect -2147 -2300 -2134 -2298
rect -2292 -2306 -2071 -2300
rect -2325 -2338 -2320 -2308
rect -2092 -2322 -2062 -2320
rect -2094 -2326 -2062 -2322
rect -2000 -2338 -1992 -2292
rect -1846 -2299 -1806 -2292
rect -1663 -2296 -1655 -2292
rect -1846 -2306 -1680 -2300
rect -1671 -2308 -1663 -2296
rect -1854 -2322 -1806 -2320
rect -1854 -2326 -1680 -2322
rect -1642 -2338 -1637 -2292
rect -1619 -2338 -1614 -2292
rect -1530 -2338 -1526 -2292
rect -1506 -2338 -1502 -2292
rect -1482 -2338 -1478 -2292
rect -1458 -2338 -1454 -2292
rect -1434 -2338 -1430 -2292
rect -1410 -2338 -1406 -2292
rect -1386 -2338 -1382 -2292
rect -1362 -2338 -1358 -2292
rect -1338 -2338 -1334 -2292
rect -1314 -2338 -1310 -2292
rect -1290 -2338 -1286 -2292
rect -1266 -2338 -1262 -2292
rect -1242 -2338 -1238 -2292
rect -1218 -2338 -1214 -2292
rect -1194 -2338 -1190 -2292
rect -1170 -2338 -1166 -2292
rect -1146 -2338 -1142 -2292
rect -1122 -2338 -1118 -2292
rect -1098 -2338 -1094 -2292
rect -1074 -2338 -1070 -2292
rect -1050 -2338 -1046 -2292
rect -1026 -2338 -1022 -2292
rect -1002 -2338 -998 -2292
rect -989 -2299 -984 -2292
rect -978 -2299 -974 -2292
rect -979 -2313 -974 -2299
rect -978 -2338 -974 -2313
rect -954 -2338 -950 -2268
rect -930 -2338 -926 -2268
rect -906 -2338 -902 -2268
rect -882 -2338 -878 -2268
rect -858 -2338 -854 -2268
rect -834 -2317 -827 -2293
rect -834 -2338 -830 -2317
rect -810 -2338 -806 -2268
rect -797 -2275 -792 -2268
rect -786 -2275 -782 -2268
rect -787 -2289 -782 -2275
rect -786 -2338 -782 -2289
rect -762 -2338 -758 -2244
rect -738 -2338 -734 -2244
rect -725 -2251 -720 -2244
rect -715 -2265 -710 -2251
rect -714 -2338 -710 -2265
rect -690 -2269 -686 -2172
rect -690 -2293 -683 -2269
rect -2393 -2340 -693 -2338
rect -2371 -2386 -2366 -2340
rect -2348 -2386 -2343 -2340
rect -2325 -2386 -2320 -2340
rect -2309 -2356 -2301 -2346
rect -2317 -2362 -2309 -2356
rect -2097 -2362 -2095 -2353
rect -2309 -2384 -2301 -2374
rect -2097 -2376 -2095 -2372
rect -2292 -2377 -2095 -2376
rect -2097 -2379 -2095 -2377
rect -2084 -2384 -2083 -2341
rect -2069 -2348 -2054 -2346
rect -2054 -2364 -2018 -2362
rect -2054 -2366 -2004 -2364
rect -2059 -2370 -2045 -2366
rect -2054 -2372 -2049 -2370
rect -2317 -2386 -2309 -2384
rect -2084 -2386 -2054 -2384
rect -2044 -2386 -2039 -2372
rect -2025 -2382 -2014 -2376
rect -2000 -2382 -1992 -2340
rect -1920 -2342 -1906 -2340
rect -1977 -2357 -1929 -2351
rect -1655 -2356 -1647 -2346
rect -1977 -2367 -1966 -2357
rect -1663 -2362 -1655 -2356
rect -1977 -2379 -1929 -2377
rect -2033 -2386 -1992 -2382
rect -1655 -2384 -1647 -2374
rect -1663 -2386 -1655 -2384
rect -1642 -2386 -1637 -2340
rect -1619 -2386 -1614 -2340
rect -1530 -2386 -1526 -2340
rect -1506 -2386 -1502 -2340
rect -1482 -2386 -1478 -2340
rect -1458 -2386 -1454 -2340
rect -1434 -2386 -1430 -2340
rect -1410 -2386 -1406 -2340
rect -1386 -2386 -1382 -2340
rect -1362 -2386 -1358 -2340
rect -1338 -2386 -1334 -2340
rect -1314 -2386 -1310 -2340
rect -1290 -2386 -1286 -2340
rect -1266 -2386 -1262 -2340
rect -1242 -2386 -1238 -2340
rect -1218 -2386 -1214 -2340
rect -1194 -2386 -1190 -2340
rect -1170 -2386 -1166 -2340
rect -1146 -2386 -1142 -2340
rect -1122 -2386 -1118 -2340
rect -1098 -2386 -1094 -2340
rect -1074 -2386 -1070 -2340
rect -1050 -2386 -1046 -2340
rect -1026 -2386 -1022 -2340
rect -1002 -2386 -998 -2340
rect -978 -2386 -974 -2340
rect -954 -2365 -950 -2340
rect -2393 -2388 -957 -2386
rect -2371 -2482 -2366 -2388
rect -2348 -2482 -2343 -2388
rect -2325 -2422 -2320 -2388
rect -2317 -2390 -2309 -2388
rect -2084 -2401 -2083 -2388
rect -2084 -2402 -2054 -2401
rect -2325 -2430 -2317 -2422
rect -2325 -2482 -2320 -2430
rect -2317 -2438 -2309 -2430
rect -2117 -2439 -2095 -2429
rect -2045 -2432 -2037 -2418
rect -2309 -2478 -2301 -2468
rect -2087 -2472 -2076 -2464
rect -2017 -2468 -2015 -2461
rect -2317 -2482 -2309 -2478
rect -2092 -2480 -2087 -2472
rect -2092 -2482 -2077 -2481
rect -2000 -2482 -1992 -2388
rect -1663 -2390 -1655 -2388
rect -1969 -2439 -1929 -2427
rect -1671 -2430 -1663 -2422
rect -1663 -2438 -1655 -2430
rect -1655 -2478 -1647 -2468
rect -1928 -2482 -1924 -2481
rect -1854 -2482 -1680 -2481
rect -1663 -2482 -1655 -2478
rect -1642 -2482 -1637 -2388
rect -1619 -2482 -1614 -2388
rect -1530 -2482 -1526 -2388
rect -1506 -2482 -1502 -2388
rect -1482 -2482 -1478 -2388
rect -1458 -2482 -1454 -2388
rect -1434 -2482 -1430 -2388
rect -1410 -2482 -1406 -2388
rect -1386 -2482 -1382 -2388
rect -1362 -2482 -1358 -2388
rect -1338 -2482 -1334 -2388
rect -1314 -2482 -1310 -2388
rect -1290 -2482 -1286 -2388
rect -1266 -2482 -1262 -2388
rect -1242 -2482 -1238 -2388
rect -1218 -2482 -1214 -2388
rect -1194 -2482 -1190 -2388
rect -1170 -2481 -1166 -2388
rect -1181 -2482 -1147 -2481
rect -2393 -2484 -1147 -2482
rect -2371 -2506 -2366 -2484
rect -2348 -2506 -2343 -2484
rect -2325 -2506 -2320 -2484
rect -2092 -2489 -2037 -2484
rect -2021 -2489 -1969 -2484
rect -1921 -2489 -1913 -2484
rect -1854 -2488 -1680 -2484
rect -2100 -2491 -2092 -2490
rect -2309 -2506 -2301 -2496
rect -2100 -2497 -2087 -2491
rect -2051 -2504 -2026 -2502
rect -2062 -2506 -2012 -2504
rect -2000 -2506 -1992 -2489
rect -1969 -2497 -1921 -2490
rect -1969 -2506 -1964 -2497
rect -1864 -2506 -1796 -2505
rect -1655 -2506 -1647 -2496
rect -1642 -2506 -1637 -2484
rect -1619 -2506 -1614 -2484
rect -1530 -2506 -1526 -2484
rect -1506 -2506 -1502 -2484
rect -1482 -2506 -1478 -2484
rect -1458 -2506 -1454 -2484
rect -1434 -2506 -1430 -2484
rect -1410 -2506 -1406 -2484
rect -1386 -2506 -1382 -2484
rect -1362 -2506 -1358 -2484
rect -1338 -2506 -1334 -2484
rect -1314 -2506 -1310 -2484
rect -1290 -2506 -1286 -2484
rect -1266 -2506 -1262 -2484
rect -1242 -2506 -1238 -2484
rect -1218 -2506 -1214 -2484
rect -1194 -2506 -1190 -2484
rect -1181 -2491 -1176 -2484
rect -1170 -2491 -1166 -2484
rect -1171 -2505 -1166 -2491
rect -1146 -2506 -1142 -2388
rect -1122 -2506 -1118 -2388
rect -1098 -2506 -1094 -2388
rect -1074 -2506 -1070 -2388
rect -1050 -2506 -1046 -2388
rect -1026 -2506 -1022 -2388
rect -1002 -2505 -998 -2388
rect -1013 -2506 -979 -2505
rect -2393 -2508 -979 -2506
rect -2371 -2554 -2366 -2508
rect -2348 -2554 -2343 -2508
rect -2325 -2554 -2320 -2508
rect -2317 -2512 -2309 -2508
rect -2105 -2515 -2092 -2512
rect -2092 -2538 -2062 -2536
rect -2094 -2542 -2062 -2538
rect -2000 -2554 -1992 -2508
rect -1663 -2512 -1655 -2508
rect -1969 -2515 -1921 -2512
rect -1854 -2538 -1806 -2536
rect -1854 -2542 -1680 -2538
rect -1926 -2554 -1892 -2551
rect -1642 -2554 -1637 -2508
rect -1619 -2554 -1614 -2508
rect -1530 -2554 -1526 -2508
rect -1506 -2554 -1502 -2508
rect -1482 -2554 -1478 -2508
rect -1458 -2554 -1454 -2508
rect -1434 -2554 -1430 -2508
rect -1410 -2554 -1406 -2508
rect -1386 -2554 -1382 -2508
rect -1362 -2554 -1358 -2508
rect -1338 -2554 -1334 -2508
rect -1314 -2554 -1310 -2508
rect -1290 -2554 -1286 -2508
rect -1266 -2554 -1262 -2508
rect -1242 -2554 -1238 -2508
rect -1218 -2553 -1214 -2508
rect -1229 -2554 -1195 -2553
rect -2393 -2556 -1195 -2554
rect -2371 -2578 -2366 -2556
rect -2348 -2578 -2343 -2556
rect -2325 -2578 -2320 -2556
rect -2054 -2557 -1906 -2556
rect -2054 -2558 -2036 -2557
rect -2309 -2572 -2301 -2562
rect -2317 -2578 -2309 -2572
rect -2068 -2573 -2038 -2566
rect -2000 -2574 -1992 -2557
rect -1920 -2558 -1906 -2557
rect -1846 -2564 -1794 -2556
rect -1852 -2571 -1804 -2566
rect -1902 -2573 -1804 -2571
rect -1655 -2572 -1647 -2562
rect -2000 -2576 -1975 -2574
rect -1902 -2575 -1852 -2573
rect -2025 -2578 -1975 -2576
rect -1846 -2578 -1804 -2575
rect -1663 -2578 -1655 -2572
rect -1642 -2578 -1637 -2556
rect -1619 -2578 -1614 -2556
rect -1530 -2578 -1526 -2556
rect -1506 -2578 -1502 -2556
rect -1482 -2578 -1478 -2556
rect -1458 -2578 -1454 -2556
rect -1434 -2578 -1430 -2556
rect -1410 -2578 -1406 -2556
rect -1386 -2578 -1382 -2556
rect -1362 -2578 -1358 -2556
rect -1338 -2578 -1334 -2556
rect -1314 -2578 -1310 -2556
rect -1290 -2578 -1286 -2556
rect -1266 -2578 -1262 -2556
rect -1242 -2578 -1238 -2556
rect -1229 -2563 -1224 -2556
rect -1218 -2563 -1214 -2556
rect -1219 -2577 -1214 -2563
rect -1194 -2578 -1190 -2508
rect -1181 -2539 -1176 -2529
rect -1171 -2553 -1166 -2539
rect -1170 -2578 -1166 -2553
rect -1146 -2557 -1142 -2508
rect -2393 -2580 -1149 -2578
rect -2371 -2602 -2366 -2580
rect -2348 -2602 -2343 -2580
rect -2325 -2602 -2320 -2580
rect -2054 -2581 -2038 -2580
rect -2000 -2581 -1966 -2580
rect -1846 -2581 -1804 -2580
rect -2000 -2582 -1975 -2581
rect -2076 -2590 -2054 -2583
rect -2309 -2600 -2301 -2590
rect -2044 -2593 -2038 -2588
rect -2028 -2590 -2001 -2583
rect -2054 -2600 -2038 -2593
rect -2015 -2591 -2001 -2590
rect -2015 -2600 -2014 -2591
rect -2317 -2602 -2309 -2600
rect -2044 -2602 -2028 -2600
rect -2000 -2602 -1992 -2582
rect -1982 -2583 -1975 -2582
rect -1862 -2583 -1798 -2582
rect -1985 -2590 -1796 -2583
rect -1862 -2591 -1798 -2590
rect -1852 -2600 -1804 -2593
rect -1655 -2600 -1647 -2590
rect -1976 -2602 -1940 -2601
rect -1663 -2602 -1655 -2600
rect -1642 -2602 -1637 -2580
rect -1619 -2602 -1614 -2580
rect -1530 -2602 -1526 -2580
rect -1506 -2602 -1502 -2580
rect -1482 -2602 -1478 -2580
rect -1458 -2602 -1454 -2580
rect -1434 -2602 -1430 -2580
rect -1410 -2602 -1406 -2580
rect -1386 -2602 -1382 -2580
rect -1362 -2602 -1358 -2580
rect -1338 -2602 -1334 -2580
rect -1314 -2602 -1310 -2580
rect -1290 -2602 -1286 -2580
rect -1266 -2602 -1262 -2580
rect -1242 -2602 -1238 -2580
rect -1229 -2602 -1195 -2601
rect -1194 -2602 -1190 -2580
rect -1170 -2602 -1166 -2580
rect -1163 -2581 -1149 -2580
rect -1146 -2581 -1139 -2557
rect -1122 -2602 -1118 -2508
rect -1098 -2602 -1094 -2508
rect -1074 -2602 -1070 -2508
rect -1050 -2602 -1046 -2508
rect -1026 -2602 -1022 -2508
rect -1013 -2515 -1008 -2508
rect -1002 -2515 -998 -2508
rect -1003 -2529 -998 -2515
rect -1013 -2554 -979 -2553
rect -978 -2554 -974 -2388
rect -971 -2389 -957 -2388
rect -954 -2389 -947 -2365
rect -954 -2554 -950 -2389
rect -930 -2554 -926 -2340
rect -906 -2554 -902 -2340
rect -882 -2554 -878 -2340
rect -858 -2554 -854 -2340
rect -834 -2554 -830 -2340
rect -810 -2554 -806 -2340
rect -786 -2554 -782 -2340
rect -762 -2341 -758 -2340
rect -762 -2365 -755 -2341
rect -762 -2554 -758 -2365
rect -738 -2554 -734 -2340
rect -714 -2554 -710 -2340
rect -707 -2341 -693 -2340
rect -690 -2341 -683 -2317
rect -690 -2554 -686 -2341
rect -666 -2554 -662 -2172
rect -642 -2554 -638 -2172
rect -618 -2554 -614 -2172
rect -594 -2554 -590 -2172
rect -570 -2554 -566 -2172
rect -546 -2554 -542 -2172
rect -522 -2554 -518 -2172
rect -498 -2554 -494 -2172
rect -474 -2554 -470 -2172
rect -450 -2554 -446 -2172
rect -426 -2554 -422 -2172
rect -413 -2395 -408 -2385
rect -402 -2395 -398 -2172
rect -403 -2409 -398 -2395
rect -413 -2434 -379 -2433
rect -378 -2434 -374 -2172
rect -354 -2434 -350 -2172
rect -341 -2419 -336 -2409
rect -330 -2419 -326 -2172
rect -331 -2433 -326 -2419
rect -306 -2434 -302 -2172
rect -282 -2434 -278 -2172
rect -258 -2434 -254 -2172
rect -234 -2434 -230 -2172
rect -210 -2434 -206 -2172
rect -186 -2434 -182 -2172
rect -162 -2434 -158 -2172
rect -138 -2434 -134 -2172
rect -114 -2434 -110 -2172
rect -90 -2434 -86 -2172
rect -66 -2434 -62 -2172
rect -42 -2434 -38 -2172
rect -18 -2434 -14 -2172
rect 6 -2434 10 -2172
rect 30 -2434 34 -2172
rect 54 -2434 58 -2172
rect 78 -2434 82 -2172
rect 102 -2434 106 -2172
rect 126 -2434 130 -2172
rect 150 -2434 154 -2172
rect 174 -2434 178 -2172
rect 198 -2434 202 -2172
rect 222 -2434 226 -2172
rect 246 -2434 250 -2172
rect 259 -2179 264 -2172
rect 270 -2179 274 -2172
rect 269 -2193 274 -2179
rect 259 -2194 293 -2193
rect 294 -2194 298 -2148
rect 318 -2194 322 -2148
rect 342 -2194 346 -2148
rect 366 -2194 370 -2148
rect 390 -2194 394 -2148
rect 414 -2194 418 -2148
rect 427 -2155 432 -2148
rect 438 -2155 442 -2148
rect 437 -2169 442 -2155
rect 427 -2170 461 -2169
rect 462 -2170 466 -2100
rect 486 -2170 490 -2100
rect 510 -2170 514 -2100
rect 534 -2170 538 -2100
rect 558 -2170 562 -2100
rect 582 -2170 586 -2100
rect 606 -2170 610 -2100
rect 619 -2107 624 -2100
rect 629 -2121 634 -2107
rect 630 -2169 634 -2121
rect 619 -2170 651 -2169
rect 427 -2172 651 -2170
rect 427 -2179 432 -2172
rect 437 -2193 442 -2179
rect 438 -2194 442 -2193
rect 462 -2194 466 -2172
rect 486 -2194 490 -2172
rect 510 -2194 514 -2172
rect 534 -2194 538 -2172
rect 558 -2194 562 -2172
rect 582 -2194 586 -2172
rect 606 -2193 610 -2172
rect 619 -2179 624 -2172
rect 630 -2179 634 -2172
rect 637 -2173 651 -2172
rect 629 -2193 634 -2179
rect 643 -2183 651 -2179
rect 637 -2193 643 -2183
rect 595 -2194 629 -2193
rect 259 -2196 629 -2194
rect 259 -2203 264 -2196
rect 269 -2217 274 -2203
rect 270 -2434 274 -2217
rect 294 -2245 298 -2196
rect 294 -2293 301 -2245
rect 294 -2434 298 -2293
rect 318 -2434 322 -2196
rect 342 -2434 346 -2196
rect 366 -2434 370 -2196
rect 390 -2434 394 -2196
rect 414 -2434 418 -2196
rect 438 -2434 442 -2196
rect 462 -2221 466 -2196
rect 462 -2269 469 -2221
rect 462 -2434 466 -2269
rect 486 -2434 490 -2196
rect 510 -2434 514 -2196
rect 534 -2434 538 -2196
rect 558 -2434 562 -2196
rect 571 -2227 576 -2217
rect 582 -2227 586 -2196
rect 595 -2203 600 -2196
rect 606 -2203 610 -2196
rect 605 -2217 610 -2203
rect 581 -2241 586 -2227
rect 571 -2347 576 -2337
rect 581 -2361 586 -2347
rect 582 -2433 586 -2361
rect 571 -2434 603 -2433
rect -413 -2436 603 -2434
rect -413 -2443 -408 -2436
rect -403 -2457 -398 -2443
rect -402 -2554 -398 -2457
rect -378 -2461 -374 -2436
rect -378 -2485 -371 -2461
rect -378 -2530 -371 -2509
rect -354 -2530 -350 -2436
rect -341 -2467 -336 -2457
rect -331 -2481 -326 -2467
rect -330 -2530 -326 -2481
rect -306 -2485 -302 -2436
rect -306 -2509 -299 -2485
rect -282 -2530 -278 -2436
rect -258 -2530 -254 -2436
rect -234 -2530 -230 -2436
rect -210 -2530 -206 -2436
rect -186 -2530 -182 -2436
rect -162 -2530 -158 -2436
rect -138 -2530 -134 -2436
rect -114 -2530 -110 -2436
rect -90 -2530 -86 -2436
rect -66 -2530 -62 -2436
rect -42 -2530 -38 -2436
rect -18 -2530 -14 -2436
rect 6 -2530 10 -2436
rect 30 -2530 34 -2436
rect 54 -2530 58 -2436
rect 78 -2530 82 -2436
rect 102 -2530 106 -2436
rect 126 -2530 130 -2436
rect 150 -2530 154 -2436
rect 174 -2530 178 -2436
rect 198 -2530 202 -2436
rect 222 -2530 226 -2436
rect 246 -2530 250 -2436
rect 270 -2530 274 -2436
rect 294 -2530 298 -2436
rect 318 -2530 322 -2436
rect 342 -2530 346 -2436
rect 366 -2530 370 -2436
rect 390 -2530 394 -2436
rect 414 -2530 418 -2436
rect 438 -2530 442 -2436
rect 462 -2530 466 -2436
rect 486 -2530 490 -2436
rect 510 -2530 514 -2436
rect 534 -2530 538 -2436
rect 558 -2529 562 -2436
rect 571 -2443 576 -2436
rect 582 -2443 586 -2436
rect 589 -2437 603 -2436
rect 581 -2457 586 -2443
rect 547 -2530 581 -2529
rect -395 -2532 581 -2530
rect -395 -2533 -381 -2532
rect -378 -2533 -371 -2532
rect -378 -2554 -374 -2533
rect -354 -2554 -350 -2532
rect -330 -2554 -326 -2532
rect -1013 -2556 -309 -2554
rect -1013 -2563 -1008 -2556
rect -1003 -2577 -998 -2563
rect -1002 -2602 -998 -2577
rect -978 -2581 -974 -2556
rect -2393 -2604 -981 -2602
rect -2371 -2674 -2366 -2604
rect -2348 -2674 -2343 -2604
rect -2325 -2638 -2320 -2604
rect -2317 -2606 -2309 -2604
rect -2076 -2617 -2054 -2610
rect -2325 -2646 -2317 -2638
rect -2060 -2644 -2030 -2641
rect -2325 -2666 -2320 -2646
rect -2317 -2654 -2309 -2646
rect -2060 -2657 -2038 -2646
rect -2033 -2653 -2030 -2644
rect -2028 -2648 -2027 -2644
rect -2068 -2662 -2038 -2659
rect -2325 -2674 -2317 -2666
rect -2000 -2674 -1992 -2604
rect -1846 -2608 -1804 -2604
rect -1663 -2606 -1655 -2604
rect -1846 -2618 -1794 -2609
rect -1912 -2629 -1884 -2627
rect -1852 -2635 -1804 -2631
rect -1844 -2644 -1796 -2641
rect -1671 -2646 -1663 -2638
rect -1844 -2657 -1804 -2646
rect -1663 -2654 -1655 -2646
rect -1852 -2662 -1680 -2658
rect -1926 -2674 -1892 -2671
rect -1671 -2674 -1663 -2666
rect -1642 -2674 -1637 -2604
rect -1619 -2674 -1614 -2604
rect -1530 -2674 -1526 -2604
rect -1506 -2674 -1502 -2604
rect -1482 -2674 -1478 -2604
rect -1458 -2674 -1454 -2604
rect -1434 -2674 -1430 -2604
rect -1410 -2674 -1406 -2604
rect -1386 -2674 -1382 -2604
rect -1362 -2674 -1358 -2604
rect -1338 -2674 -1334 -2604
rect -1314 -2674 -1310 -2604
rect -1290 -2674 -1286 -2604
rect -1266 -2674 -1262 -2604
rect -1242 -2674 -1238 -2604
rect -1229 -2611 -1224 -2604
rect -1219 -2625 -1214 -2611
rect -1218 -2674 -1214 -2625
rect -1194 -2629 -1190 -2604
rect -1194 -2653 -1187 -2629
rect -1170 -2674 -1166 -2604
rect -1146 -2626 -1139 -2605
rect -1122 -2626 -1118 -2604
rect -1098 -2626 -1094 -2604
rect -1074 -2626 -1070 -2604
rect -1050 -2626 -1046 -2604
rect -1026 -2626 -1022 -2604
rect -1002 -2625 -998 -2604
rect -995 -2605 -981 -2604
rect -978 -2605 -971 -2581
rect -1013 -2626 -979 -2625
rect -1163 -2628 -979 -2626
rect -1163 -2629 -1149 -2628
rect -1146 -2629 -1139 -2628
rect -1146 -2674 -1142 -2629
rect -1122 -2674 -1118 -2628
rect -1098 -2674 -1094 -2628
rect -1074 -2674 -1070 -2628
rect -1050 -2674 -1046 -2628
rect -1026 -2674 -1022 -2628
rect -1013 -2635 -1008 -2628
rect -1002 -2635 -998 -2628
rect -1003 -2649 -998 -2635
rect -989 -2639 -981 -2635
rect -995 -2649 -989 -2639
rect -1013 -2659 -1008 -2649
rect -995 -2650 -979 -2649
rect -978 -2650 -971 -2629
rect -954 -2650 -950 -2556
rect -930 -2650 -926 -2556
rect -906 -2650 -902 -2556
rect -882 -2650 -878 -2556
rect -858 -2650 -854 -2556
rect -834 -2650 -830 -2556
rect -810 -2650 -806 -2556
rect -786 -2650 -782 -2556
rect -762 -2650 -758 -2556
rect -738 -2650 -734 -2556
rect -714 -2650 -710 -2556
rect -690 -2650 -686 -2556
rect -666 -2650 -662 -2556
rect -642 -2650 -638 -2556
rect -629 -2587 -624 -2577
rect -618 -2587 -614 -2556
rect -619 -2601 -614 -2587
rect -629 -2626 -595 -2625
rect -594 -2626 -590 -2556
rect -570 -2626 -566 -2556
rect -546 -2626 -542 -2556
rect -522 -2626 -518 -2556
rect -498 -2626 -494 -2556
rect -474 -2626 -470 -2556
rect -450 -2626 -446 -2556
rect -426 -2626 -422 -2556
rect -402 -2626 -398 -2556
rect -378 -2626 -374 -2556
rect -354 -2626 -350 -2556
rect -330 -2626 -326 -2556
rect -323 -2557 -309 -2556
rect -306 -2557 -299 -2533
rect -306 -2626 -302 -2557
rect -282 -2626 -278 -2532
rect -258 -2626 -254 -2532
rect -234 -2626 -230 -2532
rect -210 -2626 -206 -2532
rect -186 -2626 -182 -2532
rect -162 -2626 -158 -2532
rect -138 -2626 -134 -2532
rect -114 -2626 -110 -2532
rect -90 -2626 -86 -2532
rect -66 -2626 -62 -2532
rect -42 -2626 -38 -2532
rect -18 -2626 -14 -2532
rect 6 -2626 10 -2532
rect 30 -2626 34 -2532
rect 54 -2626 58 -2532
rect 78 -2626 82 -2532
rect 102 -2626 106 -2532
rect 126 -2626 130 -2532
rect 150 -2626 154 -2532
rect 163 -2611 168 -2601
rect 174 -2611 178 -2532
rect 173 -2625 178 -2611
rect 198 -2626 202 -2532
rect 222 -2626 226 -2532
rect 246 -2626 250 -2532
rect 270 -2626 274 -2532
rect 294 -2626 298 -2532
rect 318 -2626 322 -2532
rect 342 -2626 346 -2532
rect 366 -2626 370 -2532
rect 390 -2626 394 -2532
rect 414 -2626 418 -2532
rect 438 -2626 442 -2532
rect 462 -2626 466 -2532
rect 486 -2626 490 -2532
rect 510 -2625 514 -2532
rect 523 -2563 528 -2553
rect 534 -2563 538 -2532
rect 547 -2539 552 -2532
rect 558 -2539 562 -2532
rect 557 -2553 562 -2539
rect 533 -2577 538 -2563
rect 499 -2626 533 -2625
rect -629 -2628 533 -2626
rect -629 -2635 -624 -2628
rect -619 -2649 -614 -2635
rect -618 -2650 -614 -2649
rect -594 -2650 -590 -2628
rect -570 -2650 -566 -2628
rect -546 -2650 -542 -2628
rect -522 -2650 -518 -2628
rect -498 -2650 -494 -2628
rect -474 -2650 -470 -2628
rect -450 -2650 -446 -2628
rect -426 -2650 -422 -2628
rect -402 -2650 -398 -2628
rect -378 -2650 -374 -2628
rect -354 -2650 -350 -2628
rect -330 -2650 -326 -2628
rect -306 -2650 -302 -2628
rect -282 -2650 -278 -2628
rect -258 -2650 -254 -2628
rect -234 -2650 -230 -2628
rect -210 -2650 -206 -2628
rect -186 -2650 -182 -2628
rect -162 -2650 -158 -2628
rect -138 -2650 -134 -2628
rect -114 -2650 -110 -2628
rect -90 -2650 -86 -2628
rect -66 -2650 -62 -2628
rect -42 -2650 -38 -2628
rect -18 -2650 -14 -2628
rect 6 -2650 10 -2628
rect 30 -2650 34 -2628
rect 54 -2650 58 -2628
rect 78 -2650 82 -2628
rect 102 -2650 106 -2628
rect 126 -2650 130 -2628
rect 150 -2650 154 -2628
rect 198 -2650 202 -2628
rect 222 -2650 226 -2628
rect 246 -2650 250 -2628
rect 270 -2650 274 -2628
rect 294 -2650 298 -2628
rect 318 -2650 322 -2628
rect 342 -2650 346 -2628
rect 366 -2650 370 -2628
rect 390 -2650 394 -2628
rect 414 -2650 418 -2628
rect 438 -2650 442 -2628
rect 462 -2650 466 -2628
rect 486 -2649 490 -2628
rect 499 -2635 504 -2628
rect 510 -2635 514 -2628
rect 509 -2649 514 -2635
rect 475 -2650 509 -2649
rect -995 -2652 509 -2650
rect -995 -2653 -981 -2652
rect -978 -2653 -971 -2652
rect -1003 -2673 -998 -2659
rect -1002 -2674 -998 -2673
rect -978 -2674 -974 -2653
rect -954 -2674 -950 -2652
rect -930 -2674 -926 -2652
rect -906 -2674 -902 -2652
rect -882 -2674 -878 -2652
rect -858 -2674 -854 -2652
rect -834 -2674 -830 -2652
rect -810 -2674 -806 -2652
rect -786 -2674 -782 -2652
rect -762 -2674 -758 -2652
rect -738 -2674 -734 -2652
rect -714 -2674 -710 -2652
rect -690 -2674 -686 -2652
rect -666 -2674 -662 -2652
rect -642 -2674 -638 -2652
rect -618 -2674 -614 -2652
rect -594 -2653 -590 -2652
rect -2393 -2676 -597 -2674
rect -2371 -2698 -2366 -2676
rect -2348 -2698 -2343 -2676
rect -2325 -2682 -2317 -2676
rect -2325 -2698 -2320 -2682
rect -2309 -2694 -2301 -2682
rect -2068 -2693 -2038 -2686
rect -2317 -2698 -2309 -2694
rect -2000 -2696 -1992 -2676
rect -1844 -2684 -1794 -2676
rect -1671 -2682 -1663 -2676
rect -1852 -2693 -1804 -2686
rect -1655 -2694 -1647 -2682
rect -2025 -2697 -1991 -2696
rect -2025 -2698 -1975 -2697
rect -1844 -2698 -1804 -2695
rect -1663 -2698 -1655 -2694
rect -1642 -2698 -1637 -2676
rect -1619 -2698 -1614 -2676
rect -1530 -2698 -1526 -2676
rect -1506 -2698 -1502 -2676
rect -1482 -2698 -1478 -2676
rect -1458 -2698 -1454 -2676
rect -1434 -2698 -1430 -2676
rect -1410 -2698 -1406 -2676
rect -1386 -2698 -1382 -2676
rect -1362 -2698 -1358 -2676
rect -1338 -2698 -1334 -2676
rect -1314 -2698 -1310 -2676
rect -1290 -2698 -1286 -2676
rect -1266 -2698 -1262 -2676
rect -1242 -2698 -1238 -2676
rect -1218 -2698 -1214 -2676
rect -1194 -2698 -1187 -2677
rect -1170 -2698 -1166 -2676
rect -1146 -2698 -1142 -2676
rect -1122 -2697 -1118 -2676
rect -1133 -2698 -1099 -2697
rect -2393 -2700 -1099 -2698
rect -2371 -2722 -2366 -2700
rect -2348 -2722 -2343 -2700
rect -2325 -2710 -2317 -2700
rect -2060 -2710 -2020 -2703
rect -2004 -2708 -2001 -2703
rect -2015 -2710 -2001 -2708
rect -2000 -2710 -1992 -2700
rect -1972 -2702 -1958 -2700
rect -1844 -2701 -1804 -2700
rect -1862 -2703 -1796 -2702
rect -1985 -2705 -1796 -2703
rect -1985 -2710 -1852 -2705
rect -2325 -2722 -2320 -2710
rect -2309 -2722 -2301 -2710
rect -2068 -2720 -2060 -2713
rect -2015 -2720 -1990 -2710
rect -1844 -2711 -1796 -2705
rect -1671 -2710 -1663 -2700
rect -1852 -2720 -1804 -2713
rect -2020 -2722 -2004 -2720
rect -2000 -2722 -1992 -2720
rect -1976 -2722 -1940 -2721
rect -1655 -2722 -1647 -2710
rect -1642 -2722 -1637 -2700
rect -1619 -2722 -1614 -2700
rect -1530 -2722 -1526 -2700
rect -1506 -2722 -1502 -2700
rect -1482 -2722 -1478 -2700
rect -1458 -2722 -1454 -2700
rect -1434 -2722 -1430 -2700
rect -1410 -2722 -1406 -2700
rect -1386 -2722 -1382 -2700
rect -1362 -2722 -1358 -2700
rect -1338 -2722 -1334 -2700
rect -1314 -2722 -1310 -2700
rect -1290 -2722 -1286 -2700
rect -1266 -2722 -1262 -2700
rect -1242 -2722 -1238 -2700
rect -1218 -2721 -1214 -2700
rect -1211 -2701 -1197 -2700
rect -1194 -2701 -1187 -2700
rect -1229 -2722 -1195 -2721
rect -2393 -2724 -1195 -2722
rect -2371 -2794 -2366 -2724
rect -2348 -2794 -2343 -2724
rect -2325 -2726 -2320 -2724
rect -2317 -2726 -2309 -2724
rect -2325 -2738 -2317 -2726
rect -2060 -2737 -2030 -2730
rect -2325 -2758 -2320 -2738
rect -2325 -2766 -2317 -2758
rect -2060 -2764 -2030 -2761
rect -2325 -2786 -2320 -2766
rect -2317 -2774 -2309 -2766
rect -2060 -2777 -2038 -2766
rect -2033 -2773 -2030 -2764
rect -2028 -2768 -2027 -2764
rect -2068 -2782 -2038 -2779
rect -2325 -2794 -2317 -2786
rect -2000 -2791 -1992 -2724
rect -1844 -2728 -1804 -2724
rect -1663 -2726 -1655 -2724
rect -1844 -2738 -1794 -2729
rect -1671 -2738 -1663 -2726
rect -1912 -2749 -1884 -2747
rect -1852 -2755 -1804 -2751
rect -1844 -2764 -1796 -2761
rect -1671 -2766 -1663 -2758
rect -1844 -2777 -1804 -2766
rect -1663 -2774 -1655 -2766
rect -1852 -2782 -1680 -2778
rect -2119 -2794 -2069 -2792
rect -2007 -2794 -1977 -2791
rect -1926 -2794 -1892 -2791
rect -1671 -2794 -1663 -2786
rect -1642 -2794 -1637 -2724
rect -1619 -2794 -1614 -2724
rect -1530 -2794 -1526 -2724
rect -1506 -2794 -1502 -2724
rect -1482 -2794 -1478 -2724
rect -1458 -2794 -1454 -2724
rect -1434 -2794 -1430 -2724
rect -1410 -2794 -1406 -2724
rect -1386 -2794 -1382 -2724
rect -1362 -2794 -1358 -2724
rect -1338 -2794 -1334 -2724
rect -1314 -2794 -1310 -2724
rect -1290 -2794 -1286 -2724
rect -1266 -2794 -1262 -2724
rect -1242 -2794 -1238 -2724
rect -1229 -2731 -1224 -2724
rect -1218 -2731 -1214 -2724
rect -1219 -2745 -1214 -2731
rect -1229 -2770 -1195 -2769
rect -1194 -2770 -1190 -2701
rect -1170 -2770 -1166 -2700
rect -1146 -2770 -1142 -2700
rect -1133 -2707 -1128 -2700
rect -1122 -2707 -1118 -2700
rect -1123 -2721 -1118 -2707
rect -1133 -2722 -1099 -2721
rect -1098 -2722 -1094 -2676
rect -1074 -2722 -1070 -2676
rect -1050 -2722 -1046 -2676
rect -1026 -2722 -1022 -2676
rect -1002 -2722 -998 -2676
rect -978 -2701 -974 -2676
rect -1133 -2724 -981 -2722
rect -1133 -2731 -1128 -2724
rect -1123 -2745 -1118 -2731
rect -1122 -2770 -1118 -2745
rect -1098 -2770 -1094 -2724
rect -1074 -2770 -1070 -2724
rect -1050 -2770 -1046 -2724
rect -1026 -2770 -1022 -2724
rect -1002 -2770 -998 -2724
rect -995 -2725 -981 -2724
rect -978 -2746 -971 -2701
rect -954 -2746 -950 -2676
rect -930 -2746 -926 -2676
rect -906 -2746 -902 -2676
rect -882 -2746 -878 -2676
rect -858 -2746 -854 -2676
rect -834 -2746 -830 -2676
rect -810 -2746 -806 -2676
rect -786 -2746 -782 -2676
rect -762 -2746 -758 -2676
rect -738 -2746 -734 -2676
rect -714 -2746 -710 -2676
rect -690 -2746 -686 -2676
rect -666 -2746 -662 -2676
rect -642 -2746 -638 -2676
rect -618 -2746 -614 -2676
rect -611 -2677 -597 -2676
rect -594 -2677 -587 -2653
rect -594 -2722 -587 -2701
rect -570 -2722 -566 -2652
rect -546 -2722 -542 -2652
rect -522 -2722 -518 -2652
rect -498 -2722 -494 -2652
rect -474 -2722 -470 -2652
rect -450 -2722 -446 -2652
rect -426 -2722 -422 -2652
rect -402 -2722 -398 -2652
rect -378 -2722 -374 -2652
rect -354 -2722 -350 -2652
rect -330 -2722 -326 -2652
rect -306 -2722 -302 -2652
rect -282 -2722 -278 -2652
rect -258 -2722 -254 -2652
rect -234 -2722 -230 -2652
rect -210 -2722 -206 -2652
rect -186 -2722 -182 -2652
rect -162 -2722 -158 -2652
rect -138 -2722 -134 -2652
rect -114 -2722 -110 -2652
rect -90 -2722 -86 -2652
rect -66 -2722 -62 -2652
rect -53 -2683 -48 -2673
rect -42 -2683 -38 -2652
rect -43 -2697 -38 -2683
rect -53 -2698 -19 -2697
rect -18 -2698 -14 -2652
rect 6 -2698 10 -2652
rect 30 -2698 34 -2652
rect 54 -2698 58 -2652
rect 78 -2698 82 -2652
rect 102 -2698 106 -2652
rect 126 -2698 130 -2652
rect 150 -2698 154 -2652
rect 163 -2683 168 -2673
rect 198 -2677 202 -2652
rect 173 -2697 178 -2683
rect 187 -2687 195 -2683
rect 181 -2697 187 -2687
rect 174 -2698 178 -2697
rect -53 -2700 195 -2698
rect -53 -2707 -48 -2700
rect -43 -2721 -38 -2707
rect -42 -2722 -38 -2721
rect -18 -2722 -14 -2700
rect 6 -2722 10 -2700
rect 30 -2722 34 -2700
rect 54 -2722 58 -2700
rect 78 -2722 82 -2700
rect 102 -2722 106 -2700
rect 126 -2722 130 -2700
rect 150 -2722 154 -2700
rect 174 -2722 178 -2700
rect 181 -2701 195 -2700
rect 198 -2701 205 -2677
rect 222 -2722 226 -2652
rect 246 -2722 250 -2652
rect 270 -2722 274 -2652
rect 294 -2722 298 -2652
rect 318 -2722 322 -2652
rect 342 -2722 346 -2652
rect 366 -2722 370 -2652
rect 390 -2722 394 -2652
rect 414 -2721 418 -2652
rect 427 -2707 432 -2697
rect 438 -2707 442 -2652
rect 451 -2683 456 -2673
rect 462 -2683 466 -2652
rect 475 -2659 480 -2652
rect 486 -2659 490 -2652
rect 485 -2673 490 -2659
rect 461 -2697 466 -2683
rect 437 -2721 442 -2707
rect 403 -2722 437 -2721
rect -611 -2724 437 -2722
rect -611 -2725 -597 -2724
rect -594 -2725 -587 -2724
rect -594 -2746 -590 -2725
rect -570 -2746 -566 -2724
rect -546 -2746 -542 -2724
rect -522 -2746 -518 -2724
rect -498 -2746 -494 -2724
rect -474 -2746 -470 -2724
rect -450 -2746 -446 -2724
rect -426 -2746 -422 -2724
rect -402 -2746 -398 -2724
rect -378 -2746 -374 -2724
rect -354 -2746 -350 -2724
rect -330 -2746 -326 -2724
rect -306 -2746 -302 -2724
rect -282 -2746 -278 -2724
rect -258 -2746 -254 -2724
rect -234 -2746 -230 -2724
rect -210 -2746 -206 -2724
rect -186 -2746 -182 -2724
rect -162 -2745 -158 -2724
rect -173 -2746 -139 -2745
rect -995 -2748 -139 -2746
rect -995 -2749 -981 -2748
rect -978 -2749 -971 -2748
rect -978 -2770 -974 -2749
rect -954 -2770 -950 -2748
rect -930 -2770 -926 -2748
rect -906 -2770 -902 -2748
rect -882 -2770 -878 -2748
rect -858 -2770 -854 -2748
rect -834 -2770 -830 -2748
rect -810 -2770 -806 -2748
rect -786 -2770 -782 -2748
rect -762 -2770 -758 -2748
rect -738 -2770 -734 -2748
rect -714 -2770 -710 -2748
rect -690 -2770 -686 -2748
rect -666 -2770 -662 -2748
rect -642 -2770 -638 -2748
rect -618 -2770 -614 -2748
rect -594 -2770 -590 -2748
rect -570 -2770 -566 -2748
rect -546 -2770 -542 -2748
rect -522 -2770 -518 -2748
rect -498 -2770 -494 -2748
rect -474 -2770 -470 -2748
rect -450 -2770 -446 -2748
rect -426 -2770 -422 -2748
rect -402 -2770 -398 -2748
rect -378 -2770 -374 -2748
rect -354 -2770 -350 -2748
rect -330 -2770 -326 -2748
rect -306 -2770 -302 -2748
rect -282 -2770 -278 -2748
rect -258 -2770 -254 -2748
rect -234 -2770 -230 -2748
rect -210 -2770 -206 -2748
rect -186 -2770 -182 -2748
rect -173 -2755 -168 -2748
rect -162 -2755 -158 -2748
rect -163 -2769 -158 -2755
rect -138 -2770 -134 -2724
rect -114 -2770 -110 -2724
rect -90 -2770 -86 -2724
rect -66 -2770 -62 -2724
rect -42 -2770 -38 -2724
rect -18 -2749 -14 -2724
rect -1229 -2772 -21 -2770
rect -1229 -2779 -1224 -2772
rect -1219 -2793 -1214 -2779
rect -1218 -2794 -1214 -2793
rect -1194 -2794 -1190 -2772
rect -1170 -2794 -1166 -2772
rect -1146 -2794 -1142 -2772
rect -1122 -2794 -1118 -2772
rect -1098 -2773 -1094 -2772
rect -2393 -2796 -1101 -2794
rect -2371 -2818 -2366 -2796
rect -2348 -2818 -2343 -2796
rect -2325 -2800 -2317 -2796
rect -2325 -2816 -2320 -2800
rect -2317 -2802 -2309 -2800
rect -2309 -2814 -2301 -2802
rect -2000 -2810 -1992 -2796
rect -1671 -2800 -1663 -2796
rect -1663 -2802 -1655 -2800
rect -1844 -2804 -1806 -2802
rect -1854 -2810 -1806 -2806
rect -2068 -2813 -2060 -2810
rect -2030 -2813 -1958 -2810
rect -1942 -2813 -1806 -2810
rect -2317 -2816 -2309 -2814
rect -2000 -2816 -1992 -2813
rect -1655 -2814 -1647 -2802
rect -2325 -2818 -2317 -2816
rect -2033 -2818 -1992 -2816
rect -1844 -2817 -1806 -2815
rect -1663 -2816 -1655 -2814
rect -1864 -2818 -1796 -2817
rect -1671 -2818 -1663 -2816
rect -1642 -2818 -1637 -2796
rect -1619 -2818 -1614 -2796
rect -1530 -2818 -1526 -2796
rect -1506 -2818 -1502 -2796
rect -1482 -2818 -1478 -2796
rect -1458 -2818 -1454 -2796
rect -1434 -2818 -1430 -2796
rect -1410 -2818 -1406 -2796
rect -1386 -2818 -1382 -2796
rect -1362 -2818 -1358 -2796
rect -1338 -2818 -1334 -2796
rect -1314 -2818 -1310 -2796
rect -1290 -2818 -1286 -2796
rect -1266 -2818 -1262 -2796
rect -1242 -2818 -1238 -2796
rect -1218 -2818 -1214 -2796
rect -1194 -2797 -1190 -2796
rect -2393 -2820 -1197 -2818
rect -2371 -2842 -2366 -2820
rect -2348 -2842 -2343 -2820
rect -2325 -2828 -2317 -2820
rect -2060 -2823 -2030 -2820
rect -2000 -2823 -1992 -2820
rect -1972 -2822 -1958 -2820
rect -1904 -2823 -1798 -2820
rect -2078 -2827 -2020 -2823
rect -2023 -2828 -2020 -2827
rect -2000 -2825 -1798 -2823
rect -2000 -2827 -1854 -2825
rect -1844 -2827 -1798 -2825
rect -2325 -2842 -2320 -2828
rect -2317 -2830 -2309 -2828
rect -2020 -2830 -2004 -2828
rect -2000 -2830 -1992 -2827
rect -1671 -2828 -1663 -2820
rect -2309 -2842 -2301 -2830
rect -2020 -2832 -1992 -2830
rect -1844 -2831 -1806 -2829
rect -1663 -2830 -1655 -2828
rect -2023 -2837 -1992 -2832
rect -1854 -2837 -1806 -2833
rect -2068 -2840 -2060 -2837
rect -2030 -2840 -1806 -2837
rect -2074 -2842 -2060 -2840
rect -2020 -2842 -2004 -2840
rect -2000 -2842 -1992 -2840
rect -1655 -2842 -1647 -2830
rect -1642 -2842 -1637 -2820
rect -1619 -2842 -1614 -2820
rect -1530 -2842 -1526 -2820
rect -1506 -2842 -1502 -2820
rect -1482 -2842 -1478 -2820
rect -1458 -2842 -1454 -2820
rect -1434 -2842 -1430 -2820
rect -1410 -2842 -1406 -2820
rect -1386 -2842 -1382 -2820
rect -1362 -2842 -1358 -2820
rect -1338 -2842 -1334 -2820
rect -1314 -2842 -1310 -2820
rect -1290 -2842 -1286 -2820
rect -1266 -2842 -1262 -2820
rect -1242 -2842 -1238 -2820
rect -1218 -2842 -1214 -2820
rect -1211 -2821 -1197 -2820
rect -1194 -2821 -1187 -2797
rect -1170 -2842 -1166 -2796
rect -1146 -2842 -1142 -2796
rect -1122 -2842 -1118 -2796
rect -1115 -2797 -1101 -2796
rect -1098 -2818 -1091 -2773
rect -1074 -2818 -1070 -2772
rect -1050 -2818 -1046 -2772
rect -1026 -2818 -1022 -2772
rect -1002 -2818 -998 -2772
rect -978 -2818 -974 -2772
rect -954 -2818 -950 -2772
rect -930 -2818 -926 -2772
rect -906 -2818 -902 -2772
rect -893 -2803 -888 -2793
rect -882 -2803 -878 -2772
rect -883 -2817 -878 -2803
rect -858 -2818 -854 -2772
rect -834 -2818 -830 -2772
rect -810 -2818 -806 -2772
rect -786 -2818 -782 -2772
rect -762 -2818 -758 -2772
rect -738 -2818 -734 -2772
rect -714 -2818 -710 -2772
rect -690 -2818 -686 -2772
rect -666 -2818 -662 -2772
rect -642 -2818 -638 -2772
rect -618 -2818 -614 -2772
rect -594 -2818 -590 -2772
rect -570 -2818 -566 -2772
rect -546 -2818 -542 -2772
rect -522 -2818 -518 -2772
rect -498 -2818 -494 -2772
rect -474 -2818 -470 -2772
rect -450 -2818 -446 -2772
rect -426 -2818 -422 -2772
rect -402 -2818 -398 -2772
rect -378 -2818 -374 -2772
rect -354 -2817 -350 -2772
rect -365 -2818 -331 -2817
rect -1115 -2820 -331 -2818
rect -1115 -2821 -1101 -2820
rect -1098 -2821 -1091 -2820
rect -1098 -2842 -1094 -2821
rect -1074 -2842 -1070 -2820
rect -1050 -2842 -1046 -2820
rect -1026 -2842 -1022 -2820
rect -1002 -2842 -998 -2820
rect -978 -2842 -974 -2820
rect -954 -2842 -950 -2820
rect -930 -2842 -926 -2820
rect -906 -2842 -902 -2820
rect -858 -2842 -854 -2820
rect -834 -2842 -830 -2820
rect -810 -2842 -806 -2820
rect -786 -2842 -782 -2820
rect -762 -2842 -758 -2820
rect -738 -2842 -734 -2820
rect -714 -2842 -710 -2820
rect -690 -2842 -686 -2820
rect -666 -2842 -662 -2820
rect -642 -2842 -638 -2820
rect -618 -2842 -614 -2820
rect -594 -2842 -590 -2820
rect -570 -2842 -566 -2820
rect -546 -2842 -542 -2820
rect -522 -2842 -518 -2820
rect -498 -2842 -494 -2820
rect -474 -2842 -470 -2820
rect -450 -2842 -446 -2820
rect -426 -2842 -422 -2820
rect -402 -2842 -398 -2820
rect -378 -2841 -374 -2820
rect -365 -2827 -360 -2820
rect -354 -2827 -350 -2820
rect -355 -2841 -350 -2827
rect -389 -2842 -331 -2841
rect -330 -2842 -326 -2772
rect -306 -2842 -302 -2772
rect -282 -2842 -278 -2772
rect -258 -2842 -254 -2772
rect -234 -2842 -230 -2772
rect -210 -2842 -206 -2772
rect -186 -2842 -182 -2772
rect -173 -2803 -168 -2793
rect -163 -2817 -158 -2803
rect -162 -2842 -158 -2817
rect -138 -2821 -134 -2772
rect -2393 -2844 -2060 -2842
rect -2050 -2844 -141 -2842
rect -2371 -2890 -2366 -2844
rect -2348 -2890 -2343 -2844
rect -2325 -2856 -2317 -2844
rect -2109 -2847 -2108 -2844
rect -2117 -2854 -2108 -2847
rect -2325 -2876 -2320 -2856
rect -2317 -2858 -2309 -2856
rect -2109 -2858 -2108 -2854
rect -2060 -2854 -2030 -2847
rect -2060 -2858 -2034 -2854
rect -2325 -2884 -2317 -2876
rect -2101 -2881 -2071 -2878
rect -2325 -2890 -2320 -2884
rect -2317 -2890 -2309 -2884
rect -2000 -2886 -1992 -2844
rect -1844 -2845 -1806 -2844
rect -1844 -2854 -1798 -2847
rect -1671 -2856 -1663 -2844
rect -1844 -2858 -1806 -2856
rect -1663 -2858 -1655 -2856
rect -1854 -2872 -1680 -2868
rect -1846 -2881 -1798 -2878
rect -2079 -2887 -2043 -2886
rect -2007 -2887 -1991 -2886
rect -2079 -2888 -2071 -2887
rect -2079 -2890 -2029 -2888
rect -2011 -2890 -1991 -2887
rect -1846 -2889 -1806 -2883
rect -1671 -2884 -1663 -2876
rect -1864 -2890 -1796 -2889
rect -1663 -2890 -1655 -2884
rect -1642 -2890 -1637 -2844
rect -1619 -2890 -1614 -2844
rect -1530 -2890 -1526 -2844
rect -1506 -2890 -1502 -2844
rect -1482 -2890 -1478 -2844
rect -1458 -2890 -1454 -2844
rect -1434 -2890 -1430 -2844
rect -1410 -2890 -1406 -2844
rect -1386 -2890 -1382 -2844
rect -1362 -2890 -1358 -2844
rect -1338 -2890 -1334 -2844
rect -1314 -2890 -1310 -2844
rect -1290 -2890 -1286 -2844
rect -1266 -2890 -1262 -2844
rect -1242 -2890 -1238 -2844
rect -1218 -2890 -1214 -2844
rect -1194 -2866 -1187 -2845
rect -1170 -2866 -1166 -2844
rect -1146 -2866 -1142 -2844
rect -1122 -2866 -1118 -2844
rect -1098 -2866 -1094 -2844
rect -1074 -2866 -1070 -2844
rect -1050 -2866 -1046 -2844
rect -1026 -2866 -1022 -2844
rect -1002 -2866 -998 -2844
rect -978 -2866 -974 -2844
rect -954 -2866 -950 -2844
rect -930 -2866 -926 -2844
rect -906 -2866 -902 -2844
rect -893 -2866 -859 -2865
rect -858 -2866 -854 -2844
rect -834 -2866 -830 -2844
rect -810 -2866 -806 -2844
rect -786 -2866 -782 -2844
rect -762 -2866 -758 -2844
rect -738 -2866 -734 -2844
rect -714 -2866 -710 -2844
rect -690 -2866 -686 -2844
rect -666 -2866 -662 -2844
rect -642 -2866 -638 -2844
rect -618 -2866 -614 -2844
rect -594 -2866 -590 -2844
rect -570 -2866 -566 -2844
rect -546 -2866 -542 -2844
rect -522 -2866 -518 -2844
rect -498 -2866 -494 -2844
rect -474 -2866 -470 -2844
rect -450 -2865 -446 -2844
rect -461 -2866 -427 -2865
rect -1211 -2868 -427 -2866
rect -1211 -2869 -1197 -2868
rect -1194 -2869 -1187 -2868
rect -1194 -2890 -1190 -2869
rect -1170 -2890 -1166 -2868
rect -1146 -2890 -1142 -2868
rect -1122 -2890 -1118 -2868
rect -1098 -2890 -1094 -2868
rect -1074 -2890 -1070 -2868
rect -1050 -2890 -1046 -2868
rect -1026 -2890 -1022 -2868
rect -1002 -2890 -998 -2868
rect -978 -2890 -974 -2868
rect -954 -2890 -950 -2868
rect -930 -2890 -926 -2868
rect -906 -2890 -902 -2868
rect -893 -2875 -888 -2868
rect -858 -2869 -854 -2868
rect -883 -2889 -878 -2875
rect -869 -2879 -861 -2875
rect -875 -2889 -869 -2879
rect -882 -2890 -878 -2889
rect -2393 -2892 -861 -2890
rect -2371 -2938 -2366 -2892
rect -2348 -2938 -2343 -2892
rect -2325 -2904 -2320 -2892
rect -2079 -2894 -2071 -2892
rect -2072 -2896 -2071 -2894
rect -2109 -2901 -2101 -2896
rect -2101 -2903 -2079 -2901
rect -2069 -2903 -2068 -2896
rect -2325 -2912 -2317 -2904
rect -2079 -2908 -2071 -2903
rect -2325 -2932 -2320 -2912
rect -2317 -2920 -2309 -2912
rect -2074 -2917 -2071 -2908
rect -2069 -2912 -2068 -2908
rect -2109 -2926 -2079 -2923
rect -2325 -2938 -2317 -2932
rect -2000 -2938 -1992 -2892
rect -1846 -2894 -1806 -2892
rect -1854 -2899 -1806 -2895
rect -1854 -2901 -1846 -2899
rect -1846 -2903 -1806 -2901
rect -1806 -2905 -1798 -2903
rect -1846 -2908 -1798 -2905
rect -1846 -2921 -1806 -2910
rect -1671 -2912 -1663 -2904
rect -1663 -2920 -1655 -2912
rect -1854 -2926 -1680 -2922
rect -1671 -2938 -1663 -2932
rect -1642 -2938 -1637 -2892
rect -1619 -2938 -1614 -2892
rect -1530 -2938 -1526 -2892
rect -1506 -2938 -1502 -2892
rect -1482 -2938 -1478 -2892
rect -1458 -2938 -1454 -2892
rect -1434 -2938 -1430 -2892
rect -1410 -2938 -1406 -2892
rect -1386 -2938 -1382 -2892
rect -1362 -2938 -1358 -2892
rect -1338 -2938 -1334 -2892
rect -1314 -2938 -1310 -2892
rect -1290 -2938 -1286 -2892
rect -1266 -2938 -1262 -2892
rect -1242 -2938 -1238 -2892
rect -1218 -2938 -1214 -2892
rect -1194 -2938 -1190 -2892
rect -1170 -2938 -1166 -2892
rect -1146 -2938 -1142 -2892
rect -1122 -2938 -1118 -2892
rect -1098 -2938 -1094 -2892
rect -1074 -2938 -1070 -2892
rect -1050 -2938 -1046 -2892
rect -1026 -2938 -1022 -2892
rect -1002 -2938 -998 -2892
rect -978 -2938 -974 -2892
rect -954 -2938 -950 -2892
rect -930 -2938 -926 -2892
rect -906 -2938 -902 -2892
rect -882 -2938 -878 -2892
rect -875 -2893 -861 -2892
rect -858 -2893 -851 -2869
rect -834 -2938 -830 -2868
rect -810 -2938 -806 -2868
rect -786 -2938 -782 -2868
rect -762 -2938 -758 -2868
rect -738 -2938 -734 -2868
rect -714 -2938 -710 -2868
rect -690 -2938 -686 -2868
rect -666 -2938 -662 -2868
rect -642 -2938 -638 -2868
rect -618 -2938 -614 -2868
rect -594 -2938 -590 -2868
rect -570 -2938 -566 -2868
rect -546 -2938 -542 -2868
rect -522 -2938 -518 -2868
rect -498 -2938 -494 -2868
rect -474 -2938 -470 -2868
rect -461 -2875 -456 -2868
rect -450 -2875 -446 -2868
rect -451 -2889 -446 -2875
rect -461 -2914 -427 -2913
rect -426 -2914 -422 -2844
rect -402 -2914 -398 -2844
rect -389 -2851 -384 -2844
rect -378 -2851 -374 -2844
rect -365 -2851 -360 -2844
rect -379 -2865 -374 -2851
rect -355 -2865 -350 -2851
rect -389 -2866 -355 -2865
rect -354 -2866 -350 -2865
rect -330 -2866 -326 -2844
rect -306 -2866 -302 -2844
rect -282 -2866 -278 -2844
rect -258 -2866 -254 -2844
rect -234 -2866 -230 -2844
rect -210 -2866 -206 -2844
rect -186 -2866 -182 -2844
rect -162 -2866 -158 -2844
rect -155 -2845 -141 -2844
rect -138 -2845 -131 -2821
rect -114 -2866 -110 -2772
rect -90 -2866 -86 -2772
rect -66 -2866 -62 -2772
rect -42 -2866 -38 -2772
rect -35 -2773 -21 -2772
rect -18 -2794 -11 -2749
rect 6 -2794 10 -2724
rect 30 -2794 34 -2724
rect 54 -2794 58 -2724
rect 78 -2794 82 -2724
rect 102 -2794 106 -2724
rect 126 -2794 130 -2724
rect 150 -2794 154 -2724
rect 174 -2794 178 -2724
rect 198 -2770 205 -2749
rect 222 -2770 226 -2724
rect 246 -2770 250 -2724
rect 270 -2770 274 -2724
rect 294 -2770 298 -2724
rect 318 -2770 322 -2724
rect 342 -2770 346 -2724
rect 366 -2770 370 -2724
rect 390 -2769 394 -2724
rect 403 -2731 408 -2724
rect 414 -2731 418 -2724
rect 413 -2745 418 -2731
rect 379 -2770 413 -2769
rect 181 -2772 413 -2770
rect 181 -2773 195 -2772
rect 198 -2773 205 -2772
rect 198 -2794 202 -2773
rect 222 -2794 226 -2772
rect 246 -2794 250 -2772
rect 270 -2794 274 -2772
rect 294 -2794 298 -2772
rect 318 -2794 322 -2772
rect 342 -2794 346 -2772
rect 366 -2793 370 -2772
rect 379 -2779 384 -2772
rect 390 -2779 394 -2772
rect 389 -2793 394 -2779
rect 355 -2794 389 -2793
rect -35 -2796 389 -2794
rect -35 -2797 -21 -2796
rect -18 -2797 -11 -2796
rect -18 -2866 -14 -2797
rect 6 -2866 10 -2796
rect 30 -2866 34 -2796
rect 54 -2866 58 -2796
rect 78 -2866 82 -2796
rect 102 -2866 106 -2796
rect 126 -2866 130 -2796
rect 150 -2866 154 -2796
rect 174 -2866 178 -2796
rect 198 -2866 202 -2796
rect 222 -2866 226 -2796
rect 246 -2866 250 -2796
rect 270 -2866 274 -2796
rect 294 -2866 298 -2796
rect 318 -2865 322 -2796
rect 331 -2851 336 -2841
rect 342 -2851 346 -2796
rect 355 -2803 360 -2796
rect 366 -2803 370 -2796
rect 365 -2817 370 -2803
rect 341 -2865 346 -2851
rect 307 -2866 341 -2865
rect -389 -2868 341 -2866
rect -389 -2875 -384 -2868
rect -379 -2889 -374 -2875
rect -378 -2914 -374 -2889
rect -354 -2914 -350 -2868
rect -330 -2893 -326 -2868
rect -461 -2916 -333 -2914
rect -461 -2923 -456 -2916
rect -451 -2937 -446 -2923
rect -450 -2938 -446 -2937
rect -426 -2938 -422 -2916
rect -402 -2938 -398 -2916
rect -378 -2938 -374 -2916
rect -354 -2917 -350 -2916
rect -347 -2917 -333 -2916
rect -354 -2938 -347 -2917
rect -330 -2938 -323 -2893
rect -317 -2899 -312 -2889
rect -306 -2899 -302 -2868
rect -307 -2913 -302 -2899
rect -317 -2938 -283 -2937
rect -2393 -2940 -357 -2938
rect -2371 -2962 -2366 -2940
rect -2348 -2962 -2343 -2940
rect -2325 -2948 -2317 -2940
rect -2325 -2962 -2320 -2948
rect -2309 -2960 -2301 -2948
rect -2092 -2957 -2062 -2952
rect -2000 -2960 -1992 -2940
rect -2317 -2962 -2309 -2960
rect -2000 -2962 -1983 -2960
rect -1906 -2962 -1904 -2940
rect -1806 -2948 -1680 -2942
rect -1671 -2948 -1663 -2940
rect -1854 -2957 -1806 -2952
rect -1846 -2962 -1806 -2959
rect -1655 -2960 -1647 -2948
rect -1663 -2962 -1655 -2960
rect -1642 -2962 -1637 -2940
rect -1619 -2962 -1614 -2940
rect -1530 -2962 -1526 -2940
rect -1506 -2962 -1502 -2940
rect -1482 -2962 -1478 -2940
rect -1458 -2962 -1454 -2940
rect -1434 -2962 -1430 -2940
rect -1410 -2962 -1406 -2940
rect -1386 -2962 -1382 -2940
rect -1362 -2962 -1358 -2940
rect -1338 -2962 -1334 -2940
rect -1314 -2962 -1310 -2940
rect -1290 -2962 -1286 -2940
rect -1266 -2962 -1262 -2940
rect -1242 -2962 -1238 -2940
rect -1218 -2962 -1214 -2940
rect -1194 -2962 -1190 -2940
rect -1170 -2961 -1166 -2940
rect -1181 -2962 -1147 -2961
rect -2393 -2964 -1147 -2962
rect -2371 -2986 -2366 -2964
rect -2348 -2986 -2343 -2964
rect -2325 -2976 -2317 -2964
rect -2071 -2968 -2062 -2964
rect -2013 -2966 -1983 -2964
rect -2000 -2967 -1983 -2966
rect -2325 -2986 -2320 -2976
rect -2309 -2986 -2301 -2976
rect -2100 -2977 -2092 -2970
rect -2064 -2972 -2062 -2969
rect -2061 -2977 -2059 -2972
rect -2071 -2982 -2062 -2977
rect -2071 -2984 -2026 -2982
rect -2066 -2986 -2012 -2984
rect -2000 -2986 -1992 -2967
rect -1906 -2969 -1904 -2964
rect -1846 -2968 -1806 -2964
rect -1846 -2975 -1798 -2970
rect -1806 -2977 -1798 -2975
rect -1671 -2976 -1663 -2964
rect -1854 -2979 -1846 -2977
rect -1854 -2984 -1806 -2979
rect -1864 -2986 -1796 -2985
rect -1655 -2986 -1647 -2976
rect -1642 -2986 -1637 -2964
rect -1619 -2986 -1614 -2964
rect -1530 -2986 -1526 -2964
rect -1506 -2986 -1502 -2964
rect -1482 -2986 -1478 -2964
rect -1458 -2986 -1454 -2964
rect -1434 -2986 -1430 -2964
rect -1410 -2986 -1406 -2964
rect -1386 -2986 -1382 -2964
rect -1362 -2986 -1358 -2964
rect -1338 -2986 -1334 -2964
rect -1314 -2986 -1310 -2964
rect -1290 -2986 -1286 -2964
rect -1266 -2986 -1262 -2964
rect -1242 -2986 -1238 -2964
rect -1218 -2986 -1214 -2964
rect -1194 -2986 -1190 -2964
rect -1181 -2971 -1176 -2964
rect -1170 -2971 -1166 -2964
rect -1171 -2985 -1166 -2971
rect -1170 -2986 -1166 -2985
rect -1146 -2986 -1142 -2940
rect -1122 -2986 -1118 -2940
rect -1098 -2986 -1094 -2940
rect -1074 -2986 -1070 -2940
rect -1050 -2986 -1046 -2940
rect -1026 -2986 -1022 -2940
rect -1002 -2986 -998 -2940
rect -978 -2986 -974 -2940
rect -954 -2986 -950 -2940
rect -930 -2986 -926 -2940
rect -906 -2986 -902 -2940
rect -882 -2986 -878 -2940
rect -858 -2965 -851 -2941
rect -858 -2986 -854 -2965
rect -834 -2985 -830 -2940
rect -845 -2986 -811 -2985
rect -2393 -2988 -811 -2986
rect -2371 -3405 -2366 -2988
rect -2361 -3385 -2353 -3375
rect -2348 -3385 -2343 -2988
rect -2351 -3401 -2343 -3385
rect -2371 -3431 -2363 -3405
rect -2383 -3603 -2376 -3593
rect -2371 -3603 -2366 -3431
rect -2373 -3614 -2366 -3603
rect -2348 -3614 -2343 -3401
rect -2325 -2992 -2320 -2988
rect -2317 -2992 -2309 -2988
rect -2325 -3004 -2317 -2992
rect -2066 -2993 -2062 -2988
rect -2147 -2996 -2134 -2994
rect -2292 -3002 -2071 -2996
rect -2325 -3119 -2320 -3004
rect -2092 -3018 -2062 -3016
rect -2094 -3022 -2062 -3018
rect -2309 -3052 -2301 -3043
rect -2317 -3059 -2309 -3052
rect -2309 -3080 -2301 -3072
rect -2251 -3078 -2093 -3072
rect -2317 -3088 -2309 -3080
rect -2154 -3085 -2138 -3082
rect -2084 -3085 -2054 -3080
rect -2143 -3098 -2138 -3092
rect -2325 -3129 -2317 -3119
rect -2325 -3148 -2320 -3129
rect -2317 -3135 -2309 -3129
rect -2243 -3146 -2221 -3138
rect -2211 -3146 -2201 -3126
rect -2073 -3146 -2065 -3128
rect -2000 -3146 -1992 -2988
rect -1846 -2995 -1806 -2988
rect -1663 -2992 -1655 -2988
rect -1846 -3002 -1680 -2996
rect -1671 -3004 -1663 -2992
rect -1854 -3018 -1806 -3016
rect -1854 -3022 -1680 -3018
rect -1915 -3052 -1906 -3042
rect -1846 -3044 -1837 -3042
rect -1790 -3044 -1680 -3042
rect -1655 -3052 -1647 -3046
rect -1905 -3061 -1896 -3052
rect -1837 -3053 -1790 -3052
rect -1837 -3068 -1798 -3055
rect -1663 -3062 -1655 -3052
rect -1798 -3078 -1790 -3073
rect -1837 -3080 -1798 -3078
rect -1655 -3080 -1647 -3074
rect -1846 -3082 -1837 -3080
rect -1846 -3085 -1798 -3082
rect -1837 -3098 -1798 -3088
rect -1663 -3090 -1655 -3080
rect -1671 -3130 -1663 -3122
rect -1655 -3130 -1647 -3128
rect -1663 -3138 -1647 -3130
rect -1642 -3138 -1637 -2988
rect -1885 -3146 -1877 -3144
rect -1708 -3146 -1672 -3144
rect -2243 -3147 -2213 -3146
rect -2325 -3157 -2317 -3148
rect -2259 -3153 -2211 -3147
rect -2183 -3153 -1877 -3146
rect -1869 -3153 -1758 -3146
rect -1710 -3152 -1672 -3146
rect -1710 -3153 -1692 -3152
rect -2211 -3157 -2201 -3153
rect -2325 -3177 -2320 -3157
rect -2317 -3164 -2309 -3157
rect -2211 -3164 -2198 -3157
rect -2325 -3185 -2317 -3177
rect -2300 -3184 -2292 -3174
rect -2243 -3183 -2228 -3172
rect -2211 -3180 -2181 -3164
rect -2211 -3183 -2201 -3180
rect -2325 -3205 -2320 -3185
rect -2317 -3193 -2309 -3185
rect -2325 -3213 -2317 -3205
rect -2325 -3233 -2320 -3213
rect -2317 -3221 -2309 -3213
rect -2325 -3242 -2317 -3233
rect -2325 -3261 -2320 -3242
rect -2317 -3249 -2309 -3242
rect -2325 -3270 -2317 -3261
rect -2325 -3290 -2320 -3270
rect -2317 -3277 -2309 -3270
rect -2325 -3298 -2317 -3290
rect -2290 -3297 -2282 -3184
rect -2251 -3194 -2240 -3190
rect -2211 -3194 -2181 -3190
rect -2251 -3197 -2181 -3194
rect -2176 -3204 -2173 -3202
rect -2240 -3211 -2173 -3204
rect -2169 -3209 -2163 -3154
rect -2073 -3190 -2065 -3153
rect -2073 -3194 -2043 -3190
rect -2000 -3194 -1992 -3153
rect -1915 -3184 -1907 -3175
rect -1963 -3190 -1955 -3184
rect -1963 -3194 -1915 -3190
rect -1885 -3194 -1877 -3153
rect -1875 -3158 -1869 -3154
rect -1829 -3176 -1781 -3174
rect -1847 -3180 -1781 -3176
rect -1778 -3180 -1771 -3154
rect -1758 -3161 -1710 -3154
rect -1718 -3168 -1710 -3161
rect -1768 -3178 -1760 -3168
rect -1718 -3170 -1700 -3168
rect -2146 -3197 -2135 -3194
rect -2105 -3197 -2043 -3194
rect -2035 -3197 -1989 -3194
rect -1973 -3197 -1915 -3194
rect -1907 -3197 -1854 -3194
rect -2073 -3199 -2043 -3197
rect -2135 -3211 -2105 -3204
rect -2065 -3206 -2043 -3199
rect -2243 -3222 -2240 -3213
rect -2221 -3219 -2213 -3211
rect -2211 -3219 -2208 -3211
rect -2203 -3218 -2173 -3211
rect -2251 -3229 -2240 -3222
rect -2211 -3222 -2203 -3219
rect -2211 -3229 -2181 -3222
rect -2073 -3229 -2043 -3222
rect -2203 -3252 -2173 -3245
rect -2262 -3270 -2240 -3260
rect -2203 -3261 -2176 -3252
rect -2083 -3263 -2075 -3253
rect -2040 -3263 -2035 -3259
rect -2073 -3275 -2043 -3263
rect -2028 -3275 -2023 -3263
rect -2000 -3270 -1992 -3197
rect -1963 -3200 -1955 -3197
rect -1963 -3201 -1915 -3200
rect -1955 -3211 -1907 -3204
rect -1885 -3208 -1877 -3197
rect -1837 -3202 -1828 -3186
rect -1758 -3193 -1750 -3178
rect -1758 -3194 -1692 -3193
rect -1837 -3204 -1833 -3202
rect -1837 -3206 -1835 -3204
rect -1887 -3211 -1851 -3208
rect -1750 -3211 -1702 -3204
rect -1885 -3216 -1877 -3211
rect -1963 -3229 -1915 -3222
rect -1905 -3261 -1897 -3216
rect -1857 -3234 -1851 -3211
rect -1760 -3219 -1758 -3218
rect -1837 -3229 -1789 -3222
rect -1758 -3228 -1750 -3222
rect -1758 -3229 -1710 -3228
rect -1955 -3264 -1915 -3261
rect -1963 -3270 -1962 -3268
rect -2000 -3273 -1981 -3270
rect -1965 -3273 -1962 -3270
rect -1955 -3270 -1907 -3266
rect -1885 -3270 -1877 -3251
rect -1857 -3264 -1851 -3252
rect -1750 -3256 -1702 -3249
rect -1829 -3264 -1789 -3262
rect -1766 -3266 -1760 -3256
rect -1829 -3270 -1781 -3266
rect -1756 -3270 -1740 -3266
rect -1680 -3270 -1672 -3152
rect -1671 -3158 -1663 -3150
rect -1645 -3154 -1637 -3138
rect -1663 -3166 -1655 -3158
rect -1671 -3186 -1663 -3178
rect -1663 -3194 -1655 -3186
rect -1671 -3214 -1663 -3206
rect -1671 -3230 -1669 -3217
rect -1663 -3222 -1655 -3214
rect -1671 -3242 -1663 -3234
rect -1663 -3250 -1655 -3242
rect -1671 -3270 -1663 -3262
rect -1955 -3273 -1837 -3270
rect -1829 -3273 -1740 -3270
rect -2206 -3283 -2176 -3280
rect -2206 -3286 -2203 -3283
rect -2161 -3285 -2145 -3276
rect -2073 -3278 -2065 -3275
rect -2073 -3279 -2043 -3278
rect -2028 -3279 -2012 -3275
rect -2073 -3286 -2065 -3280
rect -2203 -3287 -2176 -3286
rect -2065 -3287 -2043 -3286
rect -2262 -3293 -2232 -3287
rect -2176 -3293 -2173 -3287
rect -2043 -3293 -2035 -3287
rect -2325 -3318 -2320 -3298
rect -2317 -3306 -2309 -3298
rect -2153 -3299 -2146 -3295
rect -2325 -3326 -2317 -3318
rect -2300 -3322 -2292 -3312
rect -2325 -3346 -2320 -3326
rect -2317 -3334 -2309 -3326
rect -2325 -3354 -2317 -3346
rect -2325 -3374 -2320 -3354
rect -2317 -3362 -2309 -3354
rect -2290 -3355 -2282 -3322
rect -2273 -3326 -2264 -3321
rect -2206 -3326 -2176 -3321
rect -2262 -3333 -2232 -3328
rect -2198 -3337 -2176 -3326
rect -2198 -3351 -2176 -3343
rect -2166 -3359 -2158 -3311
rect -2143 -3315 -2136 -3299
rect -2143 -3326 -2113 -3321
rect -2073 -3326 -2065 -3321
rect -2065 -3328 -2043 -3326
rect -2043 -3333 -2035 -3328
rect -2065 -3354 -2043 -3339
rect -2006 -3355 -2004 -3339
rect -2265 -3369 -2260 -3363
rect -2143 -3369 -2113 -3362
rect -2270 -3370 -2240 -3369
rect -2270 -3373 -2265 -3370
rect -2325 -3382 -2317 -3374
rect -2325 -3402 -2320 -3382
rect -2317 -3390 -2309 -3382
rect -2113 -3385 -2105 -3375
rect -2291 -3397 -2270 -3390
rect -2198 -3392 -2168 -3390
rect -2135 -3391 -2105 -3390
rect -2103 -3391 -2095 -3385
rect -2113 -3392 -2105 -3391
rect -2065 -3392 -2035 -3390
rect -2000 -3392 -1992 -3273
rect -1963 -3280 -1960 -3273
rect -1915 -3277 -1905 -3273
rect -1963 -3281 -1955 -3280
rect -1963 -3287 -1915 -3281
rect -1989 -3314 -1973 -3311
rect -1915 -3314 -1907 -3307
rect -1990 -3349 -1989 -3328
rect -1983 -3392 -1981 -3329
rect -1885 -3338 -1877 -3273
rect -1789 -3278 -1778 -3273
rect -1837 -3281 -1829 -3280
rect -1837 -3287 -1789 -3281
rect -1756 -3282 -1740 -3273
rect -1837 -3297 -1829 -3287
rect -1872 -3316 -1867 -3306
rect -1789 -3314 -1781 -3307
rect -1776 -3314 -1769 -3297
rect -1756 -3304 -1750 -3282
rect -1671 -3286 -1669 -3275
rect -1663 -3278 -1655 -3270
rect -1671 -3298 -1663 -3290
rect -1663 -3306 -1655 -3298
rect -1702 -3316 -1696 -3310
rect -1955 -3340 -1915 -3338
rect -1963 -3342 -1955 -3340
rect -1963 -3349 -1915 -3342
rect -1963 -3357 -1955 -3349
rect -1963 -3358 -1915 -3357
rect -1973 -3364 -1965 -3361
rect -1955 -3364 -1907 -3360
rect -1974 -3367 -1907 -3364
rect -1973 -3371 -1965 -3367
rect -1963 -3371 -1960 -3369
rect -1963 -3375 -1915 -3371
rect -1963 -3383 -1955 -3375
rect -1963 -3387 -1915 -3383
rect -1963 -3390 -1955 -3387
rect -2240 -3397 -2206 -3392
rect -2198 -3397 -2143 -3392
rect -2113 -3397 -1981 -3392
rect -1915 -3397 -1907 -3390
rect -2270 -3402 -2266 -3398
rect -2086 -3401 -2070 -3397
rect -2325 -3410 -2317 -3402
rect -2270 -3409 -2240 -3402
rect -2206 -3409 -2176 -3402
rect -2325 -3430 -2320 -3410
rect -2317 -3418 -2309 -3410
rect -2270 -3414 -2266 -3409
rect -2270 -3418 -2266 -3415
rect -2198 -3418 -2176 -3411
rect -2166 -3418 -2158 -3401
rect -2143 -3409 -2113 -3402
rect -2198 -3427 -2168 -3423
rect -2325 -3438 -2317 -3430
rect -2143 -3432 -2136 -3418
rect -2085 -3423 -2060 -3422
rect -2039 -3423 -2035 -3414
rect -2135 -3430 -2105 -3423
rect -2085 -3430 -2035 -3423
rect -2029 -3430 -2025 -3423
rect -2325 -3451 -2320 -3438
rect -2317 -3446 -2309 -3438
rect -2235 -3448 -2232 -3445
rect -2325 -3477 -2317 -3451
rect -2325 -3486 -2320 -3477
rect -2325 -3494 -2317 -3486
rect -2135 -3494 -2119 -3481
rect -2000 -3489 -1992 -3397
rect -1983 -3415 -1981 -3397
rect -1955 -3415 -1915 -3414
rect -1862 -3418 -1857 -3316
rect -1706 -3320 -1702 -3316
rect -1829 -3332 -1789 -3324
rect -1671 -3326 -1663 -3318
rect -1849 -3340 -1842 -3332
rect -1790 -3340 -1781 -3332
rect -1663 -3334 -1655 -3326
rect -1837 -3349 -1829 -3342
rect -1758 -3349 -1732 -3342
rect -1748 -3358 -1732 -3349
rect -1671 -3354 -1663 -3346
rect -1829 -3367 -1781 -3360
rect -1663 -3362 -1655 -3354
rect -1829 -3373 -1789 -3369
rect -1768 -3372 -1760 -3362
rect -1758 -3373 -1750 -3372
rect -1671 -3382 -1663 -3374
rect -1837 -3385 -1780 -3382
rect -1758 -3388 -1748 -3382
rect -1708 -3388 -1690 -3382
rect -1829 -3397 -1781 -3390
rect -1680 -3399 -1672 -3382
rect -1663 -3390 -1655 -3382
rect -1829 -3408 -1791 -3402
rect -1758 -3408 -1710 -3406
rect -1758 -3415 -1692 -3408
rect -1671 -3410 -1663 -3402
rect -1955 -3426 -1907 -3423
rect -1791 -3426 -1781 -3423
rect -1991 -3430 -1839 -3426
rect -1791 -3430 -1780 -3426
rect -1680 -3433 -1672 -3415
rect -1663 -3418 -1655 -3410
rect -1839 -3443 -1791 -3436
rect -1671 -3438 -1663 -3430
rect -1829 -3449 -1791 -3445
rect -1671 -3448 -1669 -3438
rect -1663 -3446 -1655 -3438
rect -1680 -3464 -1672 -3449
rect -1642 -3464 -1637 -3154
rect -1619 -3204 -1614 -2988
rect -1619 -3230 -1611 -3204
rect -1768 -3480 -1760 -3470
rect -1758 -3487 -1710 -3480
rect -2325 -3514 -2320 -3494
rect -2317 -3502 -2306 -3494
rect -2031 -3497 -1992 -3489
rect -1750 -3491 -1710 -3487
rect -1674 -3492 -1663 -3486
rect -2307 -3510 -2306 -3502
rect -2149 -3499 -2135 -3498
rect -2149 -3503 -2119 -3499
rect -2024 -3508 -2021 -3499
rect -2325 -3522 -2317 -3514
rect -2325 -3570 -2320 -3522
rect -2317 -3530 -2306 -3522
rect -2185 -3524 -2169 -3512
rect -2056 -3515 -2040 -3511
rect -2021 -3515 -2008 -3508
rect -2056 -3526 -2054 -3516
rect -2056 -3527 -2048 -3526
rect -2307 -3566 -2306 -3558
rect -2111 -3559 -2054 -3553
rect -2325 -3578 -2314 -3570
rect -2104 -3577 -2101 -3573
rect -2325 -3598 -2320 -3578
rect -2314 -3586 -2306 -3578
rect -2104 -3580 -2101 -3578
rect -2084 -3580 -2054 -3579
rect -2000 -3580 -1992 -3497
rect -1758 -3498 -1750 -3497
rect -1758 -3499 -1749 -3498
rect -1758 -3500 -1710 -3499
rect -1663 -3502 -1658 -3492
rect -1831 -3510 -1783 -3506
rect -1784 -3523 -1783 -3510
rect -1674 -3520 -1663 -3514
rect -1826 -3525 -1796 -3524
rect -1663 -3530 -1658 -3520
rect -1654 -3524 -1647 -3514
rect -1644 -3538 -1637 -3524
rect -1758 -3556 -1750 -3553
rect -1758 -3559 -1710 -3556
rect -1844 -3571 -1828 -3569
rect -1844 -3572 -1792 -3571
rect -1828 -3573 -1792 -3572
rect -1772 -3573 -1758 -3565
rect -1750 -3568 -1702 -3561
rect -1750 -3576 -1710 -3572
rect -1700 -3576 -1692 -3556
rect -1674 -3564 -1665 -3556
rect -1674 -3576 -1666 -3568
rect -1758 -3580 -1710 -3579
rect -2307 -3594 -2306 -3586
rect -2139 -3590 -2123 -3581
rect -2111 -3586 -2016 -3580
rect -2139 -3597 -2111 -3590
rect -2325 -3606 -2314 -3598
rect -2177 -3604 -2161 -3603
rect -2141 -3604 -2119 -3602
rect -2104 -3604 -2101 -3586
rect -2076 -3597 -2046 -3592
rect -2325 -3614 -2320 -3606
rect -2314 -3614 -2306 -3606
rect -2076 -3608 -2054 -3602
rect -2021 -3605 -2016 -3586
rect -2000 -3586 -1818 -3580
rect -1802 -3586 -1776 -3580
rect -1760 -3586 -1710 -3580
rect -1666 -3584 -1658 -3576
rect -2189 -3614 -2175 -3609
rect -2373 -3616 -2175 -3614
rect -2373 -3617 -2359 -3616
rect -2371 -4029 -2366 -3617
rect -2348 -3669 -2343 -3616
rect -2325 -3626 -2320 -3616
rect -2307 -3622 -2306 -3616
rect -2189 -3617 -2175 -3616
rect -2149 -3618 -2119 -3609
rect -2084 -3610 -2036 -3609
rect -2000 -3610 -1992 -3586
rect -1758 -3588 -1710 -3586
rect -1758 -3590 -1755 -3588
rect -1828 -3597 -1792 -3590
rect -1768 -3599 -1760 -3592
rect -1758 -3597 -1757 -3590
rect -1710 -3591 -1702 -3590
rect -1750 -3597 -1702 -3591
rect -1674 -3592 -1665 -3584
rect -1768 -3602 -1764 -3599
rect -1758 -3602 -1755 -3597
rect -1818 -3610 -1789 -3602
rect -1758 -3609 -1754 -3602
rect -1750 -3607 -1710 -3602
rect -1674 -3604 -1666 -3596
rect -1758 -3610 -1692 -3609
rect -2084 -3612 -1692 -3610
rect -1666 -3612 -1658 -3604
rect -2084 -3615 -1690 -3612
rect -2084 -3618 -2054 -3615
rect -2046 -3617 -1710 -3615
rect -2325 -3634 -2314 -3626
rect -2076 -3627 -2046 -3620
rect -2325 -3654 -2320 -3634
rect -2314 -3642 -2306 -3634
rect -2076 -3635 -2054 -3629
rect -2084 -3639 -2054 -3637
rect -2104 -3642 -2054 -3639
rect -2307 -3650 -2306 -3642
rect -2084 -3645 -2054 -3642
rect -2325 -3666 -2314 -3654
rect -2348 -3693 -2341 -3669
rect -2325 -3683 -2320 -3666
rect -2314 -3670 -2309 -3666
rect -2309 -3682 -2298 -3670
rect -2314 -3683 -2309 -3682
rect -2361 -4009 -2353 -3999
rect -2348 -4009 -2343 -3693
rect -2351 -4025 -2343 -4009
rect -2371 -4055 -2363 -4029
rect -2383 -4227 -2376 -4217
rect -2371 -4227 -2366 -4055
rect -2373 -4238 -2366 -4227
rect -2348 -4238 -2343 -4025
rect -2325 -3695 -2314 -3683
rect -2076 -3694 -2073 -3678
rect -2325 -3712 -2320 -3695
rect -2314 -3698 -2309 -3695
rect -2309 -3710 -2298 -3698
rect -2251 -3702 -2101 -3695
rect -2141 -3709 -2111 -3703
rect -2086 -3705 -2083 -3695
rect -2076 -3709 -2046 -3703
rect -2314 -3712 -2309 -3710
rect -2325 -3724 -2314 -3712
rect -2141 -3721 -2113 -3716
rect -2076 -3721 -2073 -3718
rect -2325 -3743 -2320 -3724
rect -2314 -3726 -2309 -3724
rect -2325 -3753 -2317 -3743
rect -2325 -3772 -2320 -3753
rect -2317 -3759 -2309 -3753
rect -2243 -3770 -2221 -3762
rect -2211 -3770 -2201 -3750
rect -2073 -3770 -2065 -3752
rect -2000 -3770 -1992 -3617
rect -1758 -3618 -1710 -3617
rect -1680 -3620 -1665 -3612
rect -1750 -3627 -1702 -3620
rect -1680 -3624 -1672 -3620
rect -1680 -3629 -1666 -3624
rect -1836 -3633 -1820 -3632
rect -1837 -3637 -1820 -3633
rect -1750 -3635 -1710 -3629
rect -1674 -3632 -1666 -3629
rect -1837 -3644 -1789 -3637
rect -1758 -3638 -1710 -3637
rect -1760 -3641 -1692 -3638
rect -1666 -3640 -1658 -3632
rect -1837 -3645 -1820 -3644
rect -1764 -3645 -1692 -3641
rect -1674 -3645 -1665 -3640
rect -1680 -3648 -1665 -3645
rect -1680 -3676 -1672 -3648
rect -1666 -3668 -1665 -3658
rect -1837 -3678 -1789 -3676
rect -1829 -3692 -1789 -3678
rect -1655 -3680 -1650 -3670
rect -1666 -3686 -1655 -3680
rect -1778 -3694 -1771 -3692
rect -1710 -3694 -1702 -3692
rect -1666 -3696 -1665 -3686
rect -1837 -3702 -1829 -3696
rect -1829 -3703 -1789 -3702
rect -1726 -3703 -1710 -3702
rect -1789 -3705 -1781 -3703
rect -1829 -3709 -1781 -3705
rect -1750 -3709 -1710 -3703
rect -1829 -3721 -1789 -3712
rect -1726 -3718 -1710 -3709
rect -1706 -3718 -1702 -3705
rect -1655 -3708 -1650 -3698
rect -1666 -3714 -1655 -3708
rect -1666 -3724 -1665 -3714
rect -1671 -3754 -1663 -3746
rect -1655 -3754 -1647 -3752
rect -1663 -3762 -1647 -3754
rect -1642 -3762 -1637 -3538
rect -1619 -3540 -1614 -3230
rect -1885 -3770 -1877 -3768
rect -1708 -3770 -1672 -3768
rect -2243 -3771 -2213 -3770
rect -2325 -3781 -2317 -3772
rect -2259 -3777 -2211 -3771
rect -2183 -3777 -1877 -3770
rect -1869 -3777 -1758 -3770
rect -1710 -3776 -1672 -3770
rect -1710 -3777 -1692 -3776
rect -2211 -3781 -2201 -3777
rect -2325 -3801 -2320 -3781
rect -2317 -3788 -2309 -3781
rect -2211 -3788 -2198 -3781
rect -2325 -3809 -2317 -3801
rect -2300 -3808 -2292 -3798
rect -2243 -3807 -2228 -3796
rect -2211 -3804 -2181 -3788
rect -2211 -3807 -2201 -3804
rect -2325 -3829 -2320 -3809
rect -2317 -3817 -2309 -3809
rect -2325 -3837 -2317 -3829
rect -2325 -3857 -2320 -3837
rect -2317 -3845 -2309 -3837
rect -2325 -3866 -2317 -3857
rect -2325 -3885 -2320 -3866
rect -2317 -3873 -2309 -3866
rect -2325 -3894 -2317 -3885
rect -2325 -3914 -2320 -3894
rect -2317 -3901 -2309 -3894
rect -2325 -3922 -2317 -3914
rect -2290 -3921 -2282 -3808
rect -2251 -3818 -2240 -3814
rect -2211 -3818 -2181 -3814
rect -2251 -3821 -2181 -3818
rect -2176 -3828 -2173 -3826
rect -2240 -3835 -2173 -3828
rect -2169 -3833 -2163 -3778
rect -2073 -3814 -2065 -3777
rect -2073 -3818 -2043 -3814
rect -2000 -3818 -1992 -3777
rect -1915 -3808 -1907 -3799
rect -1963 -3814 -1955 -3808
rect -1963 -3818 -1915 -3814
rect -1885 -3818 -1877 -3777
rect -1875 -3782 -1869 -3778
rect -1829 -3800 -1781 -3798
rect -1847 -3804 -1781 -3800
rect -1778 -3804 -1771 -3778
rect -1758 -3785 -1710 -3778
rect -1718 -3792 -1710 -3785
rect -1768 -3802 -1760 -3792
rect -1718 -3794 -1700 -3792
rect -2146 -3821 -2135 -3818
rect -2105 -3821 -2043 -3818
rect -2035 -3821 -1989 -3818
rect -1973 -3821 -1915 -3818
rect -1907 -3821 -1854 -3818
rect -2073 -3823 -2043 -3821
rect -2135 -3835 -2105 -3828
rect -2065 -3830 -2043 -3823
rect -2243 -3846 -2240 -3837
rect -2221 -3843 -2213 -3835
rect -2211 -3843 -2208 -3835
rect -2203 -3842 -2173 -3835
rect -2251 -3853 -2240 -3846
rect -2211 -3846 -2203 -3843
rect -2211 -3853 -2181 -3846
rect -2073 -3853 -2043 -3846
rect -2203 -3876 -2173 -3869
rect -2262 -3894 -2240 -3884
rect -2203 -3885 -2176 -3876
rect -2083 -3887 -2075 -3877
rect -2040 -3887 -2035 -3883
rect -2073 -3899 -2043 -3887
rect -2028 -3899 -2023 -3887
rect -2000 -3894 -1992 -3821
rect -1963 -3824 -1955 -3821
rect -1963 -3825 -1915 -3824
rect -1955 -3835 -1907 -3828
rect -1885 -3832 -1877 -3821
rect -1837 -3826 -1828 -3810
rect -1758 -3817 -1750 -3802
rect -1758 -3818 -1692 -3817
rect -1837 -3828 -1833 -3826
rect -1837 -3830 -1835 -3828
rect -1887 -3835 -1851 -3832
rect -1750 -3835 -1702 -3828
rect -1885 -3840 -1877 -3835
rect -1963 -3853 -1915 -3846
rect -1905 -3885 -1897 -3840
rect -1857 -3858 -1851 -3835
rect -1760 -3843 -1758 -3842
rect -1837 -3853 -1789 -3846
rect -1758 -3852 -1750 -3846
rect -1758 -3853 -1710 -3852
rect -1955 -3888 -1915 -3885
rect -1963 -3894 -1962 -3892
rect -2000 -3897 -1981 -3894
rect -1965 -3897 -1962 -3894
rect -1955 -3894 -1907 -3890
rect -1885 -3894 -1877 -3875
rect -1857 -3888 -1851 -3876
rect -1750 -3880 -1702 -3873
rect -1829 -3888 -1789 -3886
rect -1766 -3890 -1760 -3880
rect -1829 -3894 -1781 -3890
rect -1756 -3894 -1740 -3890
rect -1680 -3894 -1672 -3776
rect -1671 -3782 -1663 -3774
rect -1645 -3778 -1637 -3762
rect -1663 -3790 -1655 -3782
rect -1671 -3810 -1663 -3802
rect -1663 -3818 -1655 -3810
rect -1671 -3838 -1663 -3830
rect -1671 -3854 -1669 -3841
rect -1663 -3846 -1655 -3838
rect -1671 -3866 -1663 -3858
rect -1663 -3874 -1655 -3866
rect -1671 -3894 -1663 -3886
rect -1955 -3897 -1837 -3894
rect -1829 -3897 -1740 -3894
rect -2206 -3907 -2176 -3904
rect -2206 -3910 -2203 -3907
rect -2161 -3909 -2145 -3900
rect -2073 -3902 -2065 -3899
rect -2073 -3903 -2043 -3902
rect -2028 -3903 -2012 -3899
rect -2073 -3910 -2065 -3904
rect -2203 -3911 -2176 -3910
rect -2065 -3911 -2043 -3910
rect -2262 -3917 -2232 -3911
rect -2176 -3917 -2173 -3911
rect -2043 -3917 -2035 -3911
rect -2325 -3942 -2320 -3922
rect -2317 -3930 -2309 -3922
rect -2153 -3923 -2146 -3919
rect -2325 -3950 -2317 -3942
rect -2300 -3946 -2292 -3936
rect -2325 -3970 -2320 -3950
rect -2317 -3958 -2309 -3950
rect -2325 -3978 -2317 -3970
rect -2325 -3998 -2320 -3978
rect -2317 -3986 -2309 -3978
rect -2290 -3979 -2282 -3946
rect -2273 -3950 -2264 -3945
rect -2206 -3950 -2176 -3945
rect -2262 -3957 -2232 -3952
rect -2198 -3961 -2176 -3950
rect -2198 -3975 -2176 -3967
rect -2166 -3983 -2158 -3935
rect -2143 -3939 -2136 -3923
rect -2143 -3950 -2113 -3945
rect -2073 -3950 -2065 -3945
rect -2065 -3952 -2043 -3950
rect -2043 -3957 -2035 -3952
rect -2065 -3978 -2043 -3963
rect -2006 -3979 -2004 -3963
rect -2265 -3993 -2260 -3987
rect -2143 -3993 -2113 -3986
rect -2270 -3994 -2240 -3993
rect -2270 -3997 -2265 -3994
rect -2325 -4006 -2317 -3998
rect -2325 -4026 -2320 -4006
rect -2317 -4014 -2309 -4006
rect -2113 -4009 -2105 -3999
rect -2291 -4021 -2270 -4014
rect -2198 -4016 -2168 -4014
rect -2135 -4015 -2105 -4014
rect -2103 -4015 -2095 -4009
rect -2113 -4016 -2105 -4015
rect -2065 -4016 -2035 -4014
rect -2000 -4016 -1992 -3897
rect -1963 -3904 -1960 -3897
rect -1915 -3901 -1905 -3897
rect -1963 -3905 -1955 -3904
rect -1963 -3911 -1915 -3905
rect -1989 -3938 -1973 -3935
rect -1915 -3938 -1907 -3931
rect -1990 -3973 -1989 -3952
rect -1983 -4016 -1981 -3953
rect -1885 -3962 -1877 -3897
rect -1789 -3902 -1778 -3897
rect -1837 -3905 -1829 -3904
rect -1837 -3911 -1789 -3905
rect -1756 -3906 -1740 -3897
rect -1837 -3921 -1829 -3911
rect -1872 -3940 -1867 -3930
rect -1789 -3938 -1781 -3931
rect -1776 -3938 -1769 -3921
rect -1756 -3928 -1750 -3906
rect -1671 -3910 -1669 -3899
rect -1663 -3902 -1655 -3894
rect -1671 -3922 -1663 -3914
rect -1663 -3930 -1655 -3922
rect -1702 -3940 -1696 -3934
rect -1955 -3964 -1915 -3962
rect -1963 -3966 -1955 -3964
rect -1963 -3973 -1915 -3966
rect -1963 -3981 -1955 -3973
rect -1963 -3982 -1915 -3981
rect -1973 -3988 -1965 -3985
rect -1955 -3988 -1907 -3984
rect -1974 -3991 -1907 -3988
rect -1973 -3995 -1965 -3991
rect -1963 -3995 -1960 -3993
rect -1963 -3999 -1915 -3995
rect -1963 -4007 -1955 -3999
rect -1963 -4011 -1915 -4007
rect -1963 -4014 -1955 -4011
rect -2240 -4021 -2206 -4016
rect -2198 -4021 -2143 -4016
rect -2113 -4021 -1981 -4016
rect -1915 -4021 -1907 -4014
rect -2270 -4026 -2266 -4022
rect -2086 -4025 -2070 -4021
rect -2325 -4034 -2317 -4026
rect -2270 -4033 -2240 -4026
rect -2206 -4033 -2176 -4026
rect -2325 -4054 -2320 -4034
rect -2317 -4042 -2309 -4034
rect -2270 -4038 -2266 -4033
rect -2270 -4042 -2266 -4039
rect -2198 -4042 -2176 -4035
rect -2166 -4042 -2158 -4025
rect -2143 -4033 -2113 -4026
rect -2198 -4051 -2168 -4047
rect -2325 -4062 -2317 -4054
rect -2143 -4056 -2136 -4042
rect -2085 -4047 -2060 -4046
rect -2039 -4047 -2035 -4038
rect -2135 -4054 -2105 -4047
rect -2085 -4054 -2035 -4047
rect -2029 -4054 -2025 -4047
rect -2325 -4075 -2320 -4062
rect -2317 -4070 -2309 -4062
rect -2235 -4072 -2232 -4069
rect -2325 -4101 -2317 -4075
rect -2325 -4110 -2320 -4101
rect -2325 -4118 -2317 -4110
rect -2135 -4118 -2119 -4105
rect -2000 -4113 -1992 -4021
rect -1983 -4039 -1981 -4021
rect -1955 -4039 -1915 -4038
rect -1862 -4042 -1857 -3940
rect -1706 -3944 -1702 -3940
rect -1829 -3956 -1789 -3948
rect -1671 -3950 -1663 -3942
rect -1849 -3964 -1842 -3956
rect -1790 -3964 -1781 -3956
rect -1663 -3958 -1655 -3950
rect -1837 -3973 -1829 -3966
rect -1758 -3973 -1732 -3966
rect -1748 -3982 -1732 -3973
rect -1671 -3978 -1663 -3970
rect -1829 -3991 -1781 -3984
rect -1663 -3986 -1655 -3978
rect -1829 -3997 -1789 -3993
rect -1768 -3996 -1760 -3986
rect -1758 -3997 -1750 -3996
rect -1671 -4006 -1663 -3998
rect -1837 -4009 -1780 -4006
rect -1758 -4012 -1748 -4006
rect -1708 -4012 -1690 -4006
rect -1829 -4021 -1781 -4014
rect -1680 -4023 -1672 -4006
rect -1663 -4014 -1655 -4006
rect -1829 -4032 -1791 -4026
rect -1758 -4032 -1710 -4030
rect -1758 -4039 -1692 -4032
rect -1671 -4034 -1663 -4026
rect -1955 -4050 -1907 -4047
rect -1791 -4050 -1781 -4047
rect -1991 -4054 -1839 -4050
rect -1791 -4054 -1780 -4050
rect -1680 -4057 -1672 -4039
rect -1663 -4042 -1655 -4034
rect -1839 -4067 -1791 -4060
rect -1671 -4062 -1663 -4054
rect -1829 -4073 -1791 -4069
rect -1671 -4072 -1669 -4062
rect -1663 -4070 -1655 -4062
rect -1680 -4088 -1672 -4073
rect -1642 -4088 -1637 -3778
rect -1619 -3614 -1612 -3590
rect -1619 -3828 -1614 -3614
rect -1619 -3854 -1611 -3828
rect -1768 -4104 -1760 -4094
rect -1758 -4111 -1710 -4104
rect -2325 -4138 -2320 -4118
rect -2317 -4126 -2306 -4118
rect -2031 -4121 -1992 -4113
rect -1750 -4115 -1710 -4111
rect -1674 -4116 -1663 -4110
rect -2307 -4134 -2306 -4126
rect -2149 -4123 -2135 -4122
rect -2149 -4127 -2119 -4123
rect -2024 -4132 -2021 -4123
rect -2325 -4146 -2317 -4138
rect -2325 -4194 -2320 -4146
rect -2317 -4154 -2306 -4146
rect -2185 -4148 -2169 -4136
rect -2056 -4139 -2040 -4135
rect -2021 -4139 -2008 -4132
rect -2056 -4150 -2054 -4140
rect -2056 -4151 -2048 -4150
rect -2307 -4190 -2306 -4182
rect -2111 -4183 -2054 -4177
rect -2325 -4202 -2314 -4194
rect -2104 -4201 -2101 -4197
rect -2325 -4222 -2320 -4202
rect -2314 -4210 -2306 -4202
rect -2104 -4204 -2101 -4202
rect -2084 -4204 -2054 -4203
rect -2000 -4204 -1992 -4121
rect -1758 -4122 -1750 -4121
rect -1758 -4123 -1749 -4122
rect -1758 -4124 -1710 -4123
rect -1663 -4126 -1658 -4116
rect -1831 -4134 -1783 -4130
rect -1784 -4147 -1783 -4134
rect -1674 -4144 -1663 -4138
rect -1826 -4149 -1796 -4148
rect -1663 -4154 -1658 -4144
rect -1654 -4148 -1647 -4138
rect -1644 -4162 -1637 -4148
rect -1758 -4180 -1750 -4177
rect -1758 -4183 -1710 -4180
rect -1844 -4195 -1828 -4193
rect -1844 -4196 -1792 -4195
rect -1828 -4197 -1792 -4196
rect -1772 -4197 -1758 -4189
rect -1750 -4192 -1702 -4185
rect -1750 -4200 -1710 -4196
rect -1700 -4200 -1692 -4180
rect -1674 -4188 -1665 -4180
rect -1674 -4200 -1666 -4192
rect -1758 -4204 -1710 -4203
rect -2307 -4218 -2306 -4210
rect -2139 -4214 -2123 -4205
rect -2111 -4210 -2016 -4204
rect -2139 -4221 -2111 -4214
rect -2325 -4230 -2314 -4222
rect -2177 -4228 -2161 -4227
rect -2141 -4228 -2119 -4226
rect -2104 -4228 -2101 -4210
rect -2076 -4221 -2046 -4216
rect -2325 -4238 -2320 -4230
rect -2314 -4238 -2306 -4230
rect -2076 -4232 -2054 -4226
rect -2021 -4229 -2016 -4210
rect -2000 -4210 -1818 -4204
rect -1802 -4210 -1776 -4204
rect -1760 -4210 -1710 -4204
rect -1666 -4208 -1658 -4200
rect -2189 -4238 -2175 -4233
rect -2373 -4240 -2175 -4238
rect -2373 -4241 -2359 -4240
rect -2371 -4378 -2366 -4241
rect -2348 -4293 -2343 -4240
rect -2325 -4250 -2320 -4240
rect -2307 -4246 -2306 -4240
rect -2189 -4241 -2175 -4240
rect -2149 -4242 -2119 -4233
rect -2084 -4234 -2036 -4233
rect -2000 -4234 -1992 -4210
rect -1758 -4212 -1710 -4210
rect -1758 -4214 -1755 -4212
rect -1828 -4221 -1792 -4214
rect -1768 -4223 -1760 -4216
rect -1758 -4221 -1757 -4214
rect -1710 -4215 -1702 -4214
rect -1750 -4221 -1702 -4215
rect -1674 -4216 -1665 -4208
rect -1768 -4226 -1764 -4223
rect -1758 -4226 -1755 -4221
rect -1818 -4234 -1789 -4226
rect -1758 -4233 -1754 -4226
rect -1750 -4231 -1710 -4226
rect -1674 -4228 -1666 -4220
rect -1758 -4234 -1692 -4233
rect -2084 -4236 -1692 -4234
rect -1666 -4236 -1658 -4228
rect -2084 -4239 -1690 -4236
rect -2084 -4242 -2054 -4239
rect -2046 -4241 -1710 -4239
rect -2325 -4258 -2314 -4250
rect -2076 -4251 -2046 -4244
rect -2325 -4278 -2320 -4258
rect -2314 -4266 -2306 -4258
rect -2076 -4259 -2054 -4253
rect -2084 -4263 -2054 -4261
rect -2104 -4266 -2054 -4263
rect -2307 -4274 -2306 -4266
rect -2084 -4269 -2054 -4266
rect -2325 -4292 -2314 -4278
rect -2348 -4317 -2341 -4293
rect -2325 -4308 -2320 -4292
rect -2314 -4294 -2309 -4292
rect -2309 -4306 -2298 -4294
rect -2092 -4297 -2060 -4296
rect -2062 -4302 -2060 -4297
rect -2314 -4308 -2309 -4306
rect -2348 -4378 -2343 -4317
rect -2325 -4320 -2314 -4308
rect -2076 -4312 -2062 -4302
rect -2076 -4318 -2046 -4314
rect -2014 -4315 -2003 -4306
rect -2062 -4320 -2046 -4318
rect -2325 -4336 -2320 -4320
rect -2314 -4322 -2309 -4320
rect -2076 -4321 -2062 -4320
rect -2309 -4334 -2298 -4322
rect -2092 -4327 -2076 -4321
rect -2046 -4327 -2026 -4326
rect -2314 -4336 -2309 -4334
rect -2046 -4336 -2042 -4335
rect -2325 -4348 -2314 -4336
rect -2141 -4340 -2134 -4338
rect -2052 -4340 -2046 -4336
rect -2292 -4345 -2111 -4340
rect -2096 -4342 -2046 -4340
rect -2076 -4345 -2046 -4342
rect -2325 -4378 -2320 -4348
rect -2314 -4350 -2309 -4348
rect -2092 -4362 -2062 -4360
rect -2094 -4366 -2062 -4362
rect -2000 -4378 -1992 -4241
rect -1758 -4242 -1710 -4241
rect -1680 -4244 -1665 -4236
rect -1750 -4251 -1702 -4244
rect -1680 -4248 -1672 -4244
rect -1680 -4253 -1666 -4248
rect -1836 -4257 -1820 -4256
rect -1837 -4261 -1820 -4257
rect -1750 -4259 -1710 -4253
rect -1674 -4256 -1666 -4253
rect -1837 -4268 -1789 -4261
rect -1758 -4262 -1710 -4261
rect -1760 -4265 -1692 -4262
rect -1666 -4264 -1658 -4256
rect -1837 -4269 -1820 -4268
rect -1764 -4269 -1692 -4265
rect -1674 -4269 -1665 -4264
rect -1680 -4272 -1665 -4269
rect -1750 -4288 -1702 -4286
rect -1680 -4296 -1672 -4272
rect -1671 -4292 -1666 -4276
rect -1854 -4297 -1806 -4296
rect -1829 -4312 -1806 -4302
rect -1655 -4304 -1650 -4292
rect -1666 -4308 -1655 -4304
rect -1829 -4318 -1798 -4314
rect -1680 -4315 -1672 -4312
rect -1806 -4320 -1798 -4318
rect -1671 -4320 -1666 -4308
rect -1829 -4321 -1806 -4320
rect -1854 -4323 -1829 -4321
rect -1854 -4327 -1806 -4323
rect -1829 -4339 -1806 -4329
rect -1655 -4332 -1650 -4320
rect -1666 -4336 -1655 -4332
rect -1829 -4345 -1680 -4340
rect -1671 -4348 -1666 -4336
rect -1854 -4362 -1806 -4360
rect -1854 -4366 -1680 -4362
rect -1979 -4378 -1945 -4376
rect -1642 -4378 -1637 -4162
rect -1619 -4164 -1614 -3854
rect -1619 -4238 -1612 -4214
rect -1619 -4378 -1614 -4238
rect -1530 -4378 -1526 -2988
rect -1506 -4378 -1502 -2988
rect -1482 -4378 -1478 -2988
rect -1458 -4378 -1454 -2988
rect -1445 -3811 -1440 -3801
rect -1434 -3811 -1430 -2988
rect -1435 -3825 -1430 -3811
rect -1445 -3835 -1440 -3825
rect -1435 -3849 -1430 -3835
rect -1434 -4378 -1430 -3849
rect -1410 -3877 -1406 -2988
rect -1410 -3925 -1403 -3877
rect -1410 -4378 -1406 -3925
rect -1386 -4378 -1382 -2988
rect -1373 -3139 -1368 -3129
rect -1362 -3139 -1358 -2988
rect -1363 -3153 -1358 -3139
rect -1373 -3163 -1368 -3153
rect -1363 -3177 -1358 -3163
rect -1362 -4378 -1358 -3177
rect -1338 -3205 -1334 -2988
rect -1338 -3253 -1331 -3205
rect -1338 -4378 -1334 -3253
rect -1314 -4378 -1310 -2988
rect -1290 -4378 -1286 -2988
rect -1266 -4378 -1262 -2988
rect -1242 -4378 -1238 -2988
rect -1218 -4378 -1214 -2988
rect -1194 -4378 -1190 -2988
rect -1181 -4315 -1176 -4305
rect -1170 -4315 -1166 -2988
rect -1171 -4329 -1166 -4315
rect -1170 -4378 -1166 -4329
rect -1146 -3037 -1142 -2988
rect -1146 -3061 -1139 -3037
rect -1146 -4378 -1142 -3061
rect -1122 -4378 -1118 -2988
rect -1098 -4378 -1094 -2988
rect -1074 -4378 -1070 -2988
rect -1050 -4378 -1046 -2988
rect -1037 -4339 -1032 -4329
rect -1026 -4339 -1022 -2988
rect -1027 -4353 -1022 -4339
rect -1037 -4363 -1032 -4353
rect -1027 -4377 -1022 -4363
rect -1026 -4378 -1022 -4377
rect -1002 -4378 -998 -2988
rect -978 -4378 -974 -2988
rect -954 -4378 -950 -2988
rect -941 -3547 -936 -3537
rect -930 -3547 -926 -2988
rect -931 -3561 -926 -3547
rect -941 -3571 -936 -3561
rect -931 -3585 -926 -3571
rect -930 -4378 -926 -3585
rect -906 -3613 -902 -2988
rect -906 -3661 -899 -3613
rect -906 -4378 -902 -3661
rect -882 -4378 -878 -2988
rect -858 -4378 -854 -2988
rect -845 -2995 -840 -2988
rect -834 -2995 -830 -2988
rect -835 -3009 -830 -2995
rect -845 -3019 -840 -3009
rect -835 -3033 -830 -3019
rect -834 -4378 -830 -3033
rect -810 -3061 -806 -2940
rect -810 -3109 -803 -3061
rect -810 -4378 -806 -3109
rect -786 -4378 -782 -2940
rect -762 -4378 -758 -2940
rect -738 -4378 -734 -2940
rect -714 -4378 -710 -2940
rect -690 -4378 -686 -2940
rect -666 -4378 -662 -2940
rect -642 -4378 -638 -2940
rect -618 -4378 -614 -2940
rect -594 -4378 -590 -2940
rect -570 -4378 -566 -2940
rect -546 -4378 -542 -2940
rect -522 -4378 -518 -2940
rect -498 -4378 -494 -2940
rect -474 -4378 -470 -2940
rect -461 -4171 -456 -4161
rect -450 -4171 -446 -2940
rect -426 -2941 -422 -2940
rect -426 -2965 -419 -2941
rect -426 -3010 -419 -2989
rect -402 -3010 -398 -2940
rect -378 -3010 -374 -2940
rect -371 -2941 -357 -2940
rect -354 -2940 -283 -2938
rect -354 -2941 -333 -2940
rect -330 -2941 -323 -2940
rect -354 -2965 -347 -2941
rect -354 -3010 -350 -2965
rect -330 -3010 -326 -2941
rect -317 -2947 -312 -2940
rect -307 -2961 -302 -2947
rect -306 -3010 -302 -2961
rect -282 -2965 -278 -2868
rect -282 -2989 -275 -2965
rect -258 -3010 -254 -2868
rect -234 -3010 -230 -2868
rect -210 -3010 -206 -2868
rect -186 -3010 -182 -2868
rect -162 -3010 -158 -2868
rect -138 -2893 -131 -2869
rect -138 -3010 -134 -2893
rect -114 -3010 -110 -2868
rect -90 -3010 -86 -2868
rect -66 -3010 -62 -2868
rect -42 -3010 -38 -2868
rect -18 -3010 -14 -2868
rect 6 -3010 10 -2868
rect 30 -3010 34 -2868
rect 54 -3010 58 -2868
rect 78 -3010 82 -2868
rect 102 -3010 106 -2868
rect 126 -3010 130 -2868
rect 150 -3010 154 -2868
rect 174 -3010 178 -2868
rect 198 -3010 202 -2868
rect 222 -3010 226 -2868
rect 246 -3010 250 -2868
rect 270 -3009 274 -2868
rect 283 -2923 288 -2913
rect 294 -2923 298 -2868
rect 307 -2875 312 -2868
rect 318 -2875 322 -2868
rect 317 -2889 322 -2875
rect 293 -2937 298 -2923
rect 259 -3010 293 -3009
rect -443 -3012 293 -3010
rect -443 -3013 -429 -3012
rect -426 -3013 -419 -3012
rect -451 -4185 -446 -4171
rect -461 -4195 -456 -4185
rect -451 -4209 -446 -4195
rect -450 -4378 -446 -4209
rect -426 -4237 -422 -3013
rect -426 -4282 -419 -4237
rect -402 -4282 -398 -3012
rect -378 -4282 -374 -3012
rect -354 -4282 -350 -3012
rect -330 -4282 -326 -3012
rect -306 -4282 -302 -3012
rect -282 -3037 -275 -3013
rect -282 -4282 -278 -3037
rect -258 -4282 -254 -3012
rect -234 -4282 -230 -3012
rect -210 -4282 -206 -3012
rect -186 -4282 -182 -3012
rect -162 -4282 -158 -3012
rect -138 -4282 -134 -3012
rect -125 -3763 -120 -3753
rect -114 -3763 -110 -3012
rect -115 -3777 -110 -3763
rect -125 -3787 -120 -3777
rect -115 -3801 -110 -3787
rect -114 -4282 -110 -3801
rect -90 -3829 -86 -3012
rect -90 -3877 -83 -3829
rect -90 -4282 -86 -3877
rect -66 -4282 -62 -3012
rect -42 -4282 -38 -3012
rect -18 -4282 -14 -3012
rect 6 -4282 10 -3012
rect 30 -4282 34 -3012
rect 54 -4282 58 -3012
rect 78 -4282 82 -3012
rect 102 -4282 106 -3012
rect 126 -4282 130 -3012
rect 139 -4195 144 -4185
rect 150 -4195 154 -3012
rect 163 -3835 168 -3825
rect 174 -3835 178 -3012
rect 187 -3787 192 -3777
rect 198 -3787 202 -3012
rect 211 -3571 216 -3561
rect 222 -3571 226 -3012
rect 235 -3163 240 -3153
rect 246 -3163 250 -3012
rect 259 -3019 264 -3012
rect 270 -3019 274 -3012
rect 269 -3033 274 -3019
rect 245 -3177 250 -3163
rect 221 -3585 226 -3571
rect 197 -3801 202 -3787
rect 173 -3849 178 -3835
rect 149 -4209 154 -4195
rect 139 -4282 171 -4281
rect -443 -4284 171 -4282
rect -443 -4285 -429 -4284
rect -426 -4285 -419 -4284
rect -426 -4378 -422 -4285
rect -402 -4378 -398 -4284
rect -378 -4378 -374 -4284
rect -354 -4378 -350 -4284
rect -330 -4378 -326 -4284
rect -306 -4378 -302 -4284
rect -282 -4378 -278 -4284
rect -258 -4378 -254 -4284
rect -234 -4378 -230 -4284
rect -210 -4378 -206 -4284
rect -186 -4378 -182 -4284
rect -162 -4378 -158 -4284
rect -138 -4378 -134 -4284
rect -114 -4378 -110 -4284
rect -90 -4378 -86 -4284
rect -66 -4378 -62 -4284
rect -42 -4378 -38 -4284
rect -18 -4378 -14 -4284
rect 6 -4378 10 -4284
rect 30 -4378 34 -4284
rect 54 -4378 58 -4284
rect 78 -4378 82 -4284
rect 102 -4378 106 -4284
rect 126 -4378 130 -4284
rect 139 -4291 144 -4284
rect 157 -4285 171 -4284
rect 149 -4305 154 -4291
rect 139 -4363 144 -4353
rect 150 -4363 154 -4305
rect 149 -4377 154 -4363
rect 163 -4367 171 -4363
rect 157 -4377 163 -4367
rect 139 -4378 171 -4377
rect -2393 -4380 171 -4378
rect -2371 -4426 -2366 -4380
rect -2348 -4426 -2343 -4380
rect -2325 -4426 -2320 -4380
rect -2080 -4381 -1906 -4380
rect -2080 -4382 -2036 -4381
rect -2080 -4388 -2054 -4382
rect -2309 -4396 -2301 -4390
rect -2317 -4406 -2309 -4396
rect -2070 -4397 -2040 -4390
rect -2054 -4405 -2040 -4402
rect -2000 -4407 -1992 -4381
rect -1920 -4382 -1906 -4381
rect -1850 -4388 -1846 -4380
rect -1840 -4388 -1792 -4380
rect -1969 -4400 -1966 -4391
rect -1850 -4395 -1802 -4390
rect -1906 -4397 -1802 -4395
rect -1655 -4396 -1647 -4390
rect -1906 -4398 -1850 -4397
rect -1846 -4405 -1802 -4399
rect -1663 -4406 -1655 -4396
rect -1860 -4407 -1798 -4406
rect -2078 -4414 -2070 -4407
rect -2309 -4424 -2301 -4418
rect -2317 -4426 -2309 -4424
rect -2154 -4426 -2145 -4416
rect -2044 -4417 -2040 -4412
rect -2028 -4414 -1945 -4407
rect -1929 -4414 -1794 -4407
rect -2070 -4424 -2040 -4417
rect -2044 -4426 -2028 -4424
rect -2000 -4426 -1992 -4414
rect -1860 -4415 -1798 -4414
rect -1850 -4424 -1802 -4417
rect -1655 -4424 -1647 -4418
rect -1978 -4426 -1942 -4425
rect -1663 -4426 -1655 -4424
rect -1642 -4426 -1637 -4380
rect -1619 -4426 -1614 -4380
rect -1530 -4426 -1526 -4380
rect -1506 -4426 -1502 -4380
rect -1482 -4426 -1478 -4380
rect -1458 -4426 -1454 -4380
rect -1434 -4426 -1430 -4380
rect -1410 -4426 -1406 -4380
rect -1386 -4426 -1382 -4380
rect -1362 -4426 -1358 -4380
rect -1338 -4426 -1334 -4380
rect -1314 -4426 -1310 -4380
rect -1290 -4426 -1286 -4380
rect -1266 -4426 -1262 -4380
rect -1242 -4426 -1238 -4380
rect -1218 -4426 -1214 -4380
rect -1194 -4426 -1190 -4380
rect -1170 -4426 -1166 -4380
rect -1146 -4381 -1142 -4380
rect -1146 -4405 -1139 -4381
rect -1146 -4426 -1142 -4405
rect -1122 -4426 -1118 -4380
rect -1098 -4426 -1094 -4380
rect -1074 -4426 -1070 -4380
rect -1050 -4426 -1046 -4380
rect -1026 -4426 -1022 -4380
rect -1002 -4405 -998 -4380
rect -2393 -4428 -1005 -4426
rect -2371 -4522 -2366 -4428
rect -2348 -4522 -2343 -4428
rect -2325 -4466 -2320 -4428
rect -2317 -4434 -2309 -4428
rect -2145 -4432 -2138 -4428
rect -2070 -4432 -2054 -4428
rect -2078 -4441 -2054 -4434
rect -2062 -4466 -2032 -4465
rect -2000 -4466 -1992 -4428
rect -1846 -4432 -1802 -4428
rect -1846 -4442 -1792 -4433
rect -1663 -4434 -1655 -4428
rect -1942 -4464 -1937 -4452
rect -1850 -4455 -1822 -4454
rect -1850 -4459 -1802 -4455
rect -2325 -4474 -2317 -4466
rect -2062 -4468 -1961 -4466
rect -2325 -4494 -2320 -4474
rect -2317 -4482 -2309 -4474
rect -2062 -4481 -2040 -4470
rect -2032 -4475 -1961 -4468
rect -1947 -4474 -1942 -4466
rect -1842 -4468 -1794 -4465
rect -2070 -4486 -2022 -4482
rect -2325 -4508 -2317 -4494
rect -2072 -4502 -2032 -4501
rect -2102 -4508 -2032 -4502
rect -2325 -4522 -2320 -4508
rect -2317 -4510 -2309 -4508
rect -2309 -4522 -2301 -4510
rect -2070 -4517 -2062 -4512
rect -2000 -4522 -1992 -4475
rect -1942 -4476 -1937 -4474
rect -1932 -4484 -1927 -4476
rect -1912 -4479 -1896 -4473
rect -1842 -4481 -1802 -4470
rect -1671 -4474 -1663 -4466
rect -1663 -4482 -1655 -4474
rect -1850 -4486 -1680 -4482
rect -1924 -4500 -1921 -4498
rect -1806 -4508 -1680 -4502
rect -1671 -4508 -1663 -4494
rect -1663 -4510 -1655 -4508
rect -1854 -4517 -1806 -4512
rect -1974 -4522 -1964 -4521
rect -1960 -4522 -1944 -4520
rect -1842 -4522 -1806 -4519
rect -1655 -4522 -1647 -4510
rect -1642 -4522 -1637 -4428
rect -1619 -4522 -1614 -4428
rect -1530 -4522 -1526 -4428
rect -1506 -4522 -1502 -4428
rect -1482 -4522 -1478 -4428
rect -1458 -4522 -1454 -4428
rect -1434 -4522 -1430 -4428
rect -1410 -4522 -1406 -4428
rect -1386 -4522 -1382 -4428
rect -1362 -4522 -1358 -4428
rect -1338 -4522 -1334 -4428
rect -1314 -4522 -1310 -4428
rect -1290 -4522 -1286 -4428
rect -1266 -4522 -1262 -4428
rect -1242 -4522 -1238 -4428
rect -1218 -4522 -1214 -4428
rect -1194 -4522 -1190 -4428
rect -1170 -4521 -1166 -4428
rect -1181 -4522 -1147 -4521
rect -2393 -4524 -1147 -4522
rect -2371 -4546 -2366 -4524
rect -2348 -4546 -2343 -4524
rect -2325 -4536 -2317 -4524
rect -2325 -4546 -2320 -4536
rect -2317 -4538 -2309 -4536
rect -2062 -4537 -2032 -4530
rect -2309 -4546 -2301 -4538
rect -2070 -4544 -2062 -4537
rect -2000 -4542 -1992 -4524
rect -1974 -4526 -1944 -4524
rect -1960 -4527 -1944 -4526
rect -1842 -4528 -1806 -4524
rect -1842 -4535 -1798 -4530
rect -1806 -4537 -1798 -4535
rect -1671 -4536 -1663 -4524
rect -1854 -4539 -1842 -4537
rect -1663 -4538 -1655 -4536
rect -2062 -4546 -2036 -4544
rect -2393 -4548 -2036 -4546
rect -2032 -4546 -2012 -4544
rect -2004 -4546 -1974 -4542
rect -1854 -4544 -1806 -4539
rect -1864 -4546 -1796 -4545
rect -1655 -4546 -1647 -4538
rect -1642 -4546 -1637 -4524
rect -1619 -4546 -1614 -4524
rect -1530 -4546 -1526 -4524
rect -1506 -4546 -1502 -4524
rect -1482 -4545 -1478 -4524
rect -1493 -4546 -1459 -4545
rect -2032 -4548 -1459 -4546
rect -2371 -4594 -2366 -4548
rect -2348 -4594 -2343 -4548
rect -2325 -4552 -2320 -4548
rect -2309 -4550 -2301 -4548
rect -2317 -4552 -2309 -4550
rect -2325 -4564 -2317 -4552
rect -2052 -4554 -2036 -4552
rect -2052 -4556 -2032 -4554
rect -2062 -4562 -2032 -4556
rect -2325 -4594 -2320 -4564
rect -2317 -4566 -2309 -4564
rect -2092 -4578 -2062 -4576
rect -2094 -4582 -2062 -4578
rect -2000 -4594 -1992 -4548
rect -1904 -4555 -1874 -4548
rect -1842 -4555 -1806 -4548
rect -1655 -4550 -1647 -4548
rect -1663 -4552 -1655 -4550
rect -1842 -4562 -1680 -4556
rect -1671 -4564 -1663 -4552
rect -1663 -4566 -1655 -4564
rect -1854 -4578 -1806 -4576
rect -1854 -4582 -1680 -4578
rect -1642 -4594 -1637 -4548
rect -1619 -4594 -1614 -4548
rect -1530 -4594 -1526 -4548
rect -1506 -4594 -1502 -4548
rect -1493 -4555 -1488 -4548
rect -1482 -4555 -1478 -4548
rect -1483 -4569 -1478 -4555
rect -1493 -4579 -1488 -4569
rect -1483 -4593 -1478 -4579
rect -1482 -4594 -1478 -4593
rect -1458 -4594 -1454 -4524
rect -1434 -4594 -1430 -4524
rect -1410 -4594 -1406 -4524
rect -1386 -4594 -1382 -4524
rect -1362 -4594 -1358 -4524
rect -1338 -4594 -1334 -4524
rect -1314 -4594 -1310 -4524
rect -1290 -4594 -1286 -4524
rect -1266 -4594 -1262 -4524
rect -1242 -4594 -1238 -4524
rect -1218 -4594 -1214 -4524
rect -1194 -4594 -1190 -4524
rect -1181 -4531 -1176 -4524
rect -1170 -4531 -1166 -4524
rect -1171 -4545 -1166 -4531
rect -1170 -4594 -1166 -4545
rect -1146 -4594 -1142 -4428
rect -1122 -4594 -1118 -4428
rect -1098 -4594 -1094 -4428
rect -1074 -4594 -1070 -4428
rect -1050 -4594 -1046 -4428
rect -1026 -4594 -1022 -4428
rect -1019 -4429 -1005 -4428
rect -1002 -4450 -995 -4405
rect -978 -4450 -974 -4380
rect -954 -4450 -950 -4380
rect -930 -4450 -926 -4380
rect -906 -4450 -902 -4380
rect -882 -4450 -878 -4380
rect -858 -4450 -854 -4380
rect -834 -4450 -830 -4380
rect -810 -4450 -806 -4380
rect -786 -4450 -782 -4380
rect -762 -4450 -758 -4380
rect -738 -4450 -734 -4380
rect -714 -4450 -710 -4380
rect -690 -4450 -686 -4380
rect -666 -4450 -662 -4380
rect -642 -4450 -638 -4380
rect -618 -4450 -614 -4380
rect -594 -4450 -590 -4380
rect -570 -4450 -566 -4380
rect -546 -4450 -542 -4380
rect -522 -4450 -518 -4380
rect -498 -4450 -494 -4380
rect -485 -4435 -480 -4425
rect -474 -4435 -470 -4380
rect -475 -4449 -470 -4435
rect -450 -4450 -446 -4380
rect -426 -4450 -422 -4380
rect -402 -4450 -398 -4380
rect -378 -4449 -374 -4380
rect -389 -4450 -355 -4449
rect -1019 -4452 -355 -4450
rect -1019 -4453 -1005 -4452
rect -1002 -4453 -995 -4452
rect -1002 -4594 -998 -4453
rect -978 -4594 -974 -4452
rect -954 -4594 -950 -4452
rect -930 -4594 -926 -4452
rect -906 -4594 -902 -4452
rect -882 -4594 -878 -4452
rect -858 -4594 -854 -4452
rect -834 -4594 -830 -4452
rect -810 -4594 -806 -4452
rect -786 -4594 -782 -4452
rect -762 -4594 -758 -4452
rect -738 -4594 -734 -4452
rect -714 -4594 -710 -4452
rect -690 -4594 -686 -4452
rect -666 -4594 -662 -4452
rect -642 -4594 -638 -4452
rect -618 -4594 -614 -4452
rect -594 -4594 -590 -4452
rect -570 -4594 -566 -4452
rect -546 -4594 -542 -4452
rect -522 -4594 -518 -4452
rect -498 -4594 -494 -4452
rect -485 -4474 -451 -4473
rect -450 -4474 -446 -4452
rect -426 -4474 -422 -4452
rect -402 -4474 -398 -4452
rect -389 -4459 -384 -4452
rect -378 -4459 -374 -4452
rect -379 -4473 -374 -4459
rect -354 -4474 -350 -4380
rect -330 -4474 -326 -4380
rect -306 -4474 -302 -4380
rect -282 -4474 -278 -4380
rect -258 -4474 -254 -4380
rect -234 -4474 -230 -4380
rect -210 -4474 -206 -4380
rect -186 -4474 -182 -4380
rect -162 -4474 -158 -4380
rect -138 -4474 -134 -4380
rect -114 -4474 -110 -4380
rect -90 -4474 -86 -4380
rect -66 -4474 -62 -4380
rect -42 -4474 -38 -4380
rect -18 -4474 -14 -4380
rect 6 -4474 10 -4380
rect 30 -4474 34 -4380
rect 54 -4474 58 -4380
rect 78 -4474 82 -4380
rect 102 -4474 106 -4380
rect 126 -4474 130 -4380
rect 139 -4387 144 -4380
rect 157 -4381 171 -4380
rect 149 -4401 154 -4387
rect 150 -4473 154 -4401
rect 139 -4474 171 -4473
rect -485 -4476 171 -4474
rect -485 -4483 -480 -4476
rect -475 -4497 -470 -4483
rect -474 -4594 -470 -4497
rect -450 -4501 -446 -4476
rect -450 -4525 -443 -4501
rect -450 -4570 -443 -4549
rect -426 -4570 -422 -4476
rect -402 -4570 -398 -4476
rect -389 -4507 -384 -4497
rect -379 -4521 -374 -4507
rect -378 -4570 -374 -4521
rect -354 -4525 -350 -4476
rect -354 -4549 -347 -4525
rect -330 -4570 -326 -4476
rect -306 -4570 -302 -4476
rect -282 -4570 -278 -4476
rect -258 -4570 -254 -4476
rect -234 -4570 -230 -4476
rect -210 -4570 -206 -4476
rect -186 -4570 -182 -4476
rect -162 -4570 -158 -4476
rect -138 -4570 -134 -4476
rect -114 -4570 -110 -4476
rect -90 -4570 -86 -4476
rect -66 -4570 -62 -4476
rect -42 -4570 -38 -4476
rect -18 -4570 -14 -4476
rect 6 -4570 10 -4476
rect 30 -4570 34 -4476
rect 54 -4570 58 -4476
rect 78 -4570 82 -4476
rect 102 -4570 106 -4476
rect 126 -4569 130 -4476
rect 139 -4483 144 -4476
rect 150 -4483 154 -4476
rect 157 -4477 171 -4476
rect 149 -4497 154 -4483
rect 115 -4570 149 -4569
rect -467 -4572 149 -4570
rect -467 -4573 -453 -4572
rect -450 -4573 -443 -4572
rect -450 -4594 -446 -4573
rect -426 -4594 -422 -4572
rect -402 -4594 -398 -4572
rect -378 -4594 -374 -4572
rect -2393 -4596 -357 -4594
rect -2371 -4618 -2366 -4596
rect -2348 -4618 -2343 -4596
rect -2325 -4618 -2320 -4596
rect -2072 -4598 -2036 -4597
rect -2072 -4604 -2054 -4598
rect -2309 -4612 -2301 -4604
rect -2317 -4618 -2309 -4612
rect -2092 -4613 -2062 -4608
rect -2000 -4617 -1992 -4596
rect -1938 -4597 -1906 -4596
rect -1920 -4598 -1906 -4597
rect -1806 -4604 -1680 -4598
rect -1854 -4613 -1806 -4608
rect -1655 -4612 -1647 -4604
rect -1982 -4617 -1966 -4616
rect -2000 -4618 -1966 -4617
rect -1846 -4618 -1806 -4615
rect -1663 -4618 -1655 -4612
rect -1642 -4618 -1637 -4596
rect -1619 -4618 -1614 -4596
rect -1530 -4618 -1526 -4596
rect -1506 -4618 -1502 -4596
rect -1482 -4618 -1478 -4596
rect -1458 -4618 -1454 -4596
rect -1434 -4618 -1430 -4596
rect -1410 -4618 -1406 -4596
rect -1386 -4618 -1382 -4596
rect -1362 -4618 -1358 -4596
rect -1338 -4618 -1334 -4596
rect -1314 -4618 -1310 -4596
rect -1290 -4618 -1286 -4596
rect -1266 -4618 -1262 -4596
rect -1242 -4618 -1238 -4596
rect -1218 -4618 -1214 -4596
rect -1194 -4618 -1190 -4596
rect -1170 -4617 -1166 -4596
rect -1146 -4597 -1142 -4596
rect -1181 -4618 -1149 -4617
rect -2393 -4620 -1149 -4618
rect -2371 -4642 -2366 -4620
rect -2348 -4642 -2343 -4620
rect -2325 -4642 -2320 -4620
rect -2000 -4622 -1966 -4620
rect -2309 -4640 -2301 -4632
rect -2062 -4633 -2054 -4626
rect -2092 -4640 -2084 -4633
rect -2062 -4640 -2026 -4638
rect -2317 -4642 -2309 -4640
rect -2062 -4642 -2012 -4640
rect -2000 -4642 -1992 -4622
rect -1982 -4623 -1966 -4622
rect -1846 -4624 -1806 -4620
rect -1846 -4631 -1798 -4626
rect -1806 -4633 -1798 -4631
rect -1854 -4635 -1846 -4633
rect -1854 -4640 -1806 -4635
rect -1655 -4640 -1647 -4632
rect -1864 -4642 -1796 -4641
rect -1663 -4642 -1655 -4640
rect -1642 -4642 -1637 -4620
rect -1619 -4642 -1614 -4620
rect -1530 -4642 -1526 -4620
rect -1506 -4642 -1502 -4620
rect -1482 -4642 -1478 -4620
rect -1458 -4621 -1454 -4620
rect -2393 -4644 -1461 -4642
rect -2371 -4690 -2366 -4644
rect -2348 -4690 -2343 -4644
rect -2325 -4690 -2320 -4644
rect -2317 -4648 -2309 -4644
rect -2062 -4648 -2054 -4644
rect -2154 -4652 -2138 -4650
rect -2057 -4652 -2054 -4648
rect -2292 -4658 -2054 -4652
rect -2052 -4658 -2044 -4648
rect -2092 -4674 -2062 -4672
rect -2094 -4678 -2062 -4674
rect -2000 -4690 -1992 -4644
rect -1846 -4651 -1806 -4644
rect -1663 -4648 -1655 -4644
rect -1846 -4658 -1680 -4652
rect -1854 -4674 -1806 -4672
rect -1854 -4678 -1680 -4674
rect -1642 -4690 -1637 -4644
rect -1619 -4690 -1614 -4644
rect -1530 -4690 -1526 -4644
rect -1506 -4690 -1502 -4644
rect -1482 -4690 -1478 -4644
rect -1475 -4645 -1461 -4644
rect -1458 -4669 -1451 -4621
rect -1458 -4690 -1454 -4669
rect -1434 -4690 -1430 -4620
rect -1410 -4690 -1406 -4620
rect -1386 -4690 -1382 -4620
rect -1362 -4690 -1358 -4620
rect -1338 -4690 -1334 -4620
rect -1314 -4690 -1310 -4620
rect -1290 -4690 -1286 -4620
rect -1266 -4690 -1262 -4620
rect -1242 -4690 -1238 -4620
rect -1218 -4690 -1214 -4620
rect -1194 -4690 -1190 -4620
rect -1181 -4627 -1176 -4620
rect -1170 -4627 -1166 -4620
rect -1163 -4621 -1149 -4620
rect -1146 -4621 -1139 -4597
rect -1171 -4641 -1166 -4627
rect -1181 -4666 -1147 -4665
rect -1146 -4666 -1142 -4621
rect -1122 -4666 -1118 -4596
rect -1098 -4666 -1094 -4596
rect -1074 -4666 -1070 -4596
rect -1050 -4666 -1046 -4596
rect -1026 -4666 -1022 -4596
rect -1002 -4666 -998 -4596
rect -978 -4666 -974 -4596
rect -954 -4666 -950 -4596
rect -930 -4666 -926 -4596
rect -906 -4666 -902 -4596
rect -882 -4666 -878 -4596
rect -858 -4666 -854 -4596
rect -834 -4666 -830 -4596
rect -810 -4666 -806 -4596
rect -786 -4666 -782 -4596
rect -762 -4666 -758 -4596
rect -738 -4666 -734 -4596
rect -714 -4666 -710 -4596
rect -701 -4651 -696 -4641
rect -690 -4651 -686 -4596
rect -691 -4665 -686 -4651
rect -666 -4666 -662 -4596
rect -642 -4666 -638 -4596
rect -618 -4666 -614 -4596
rect -594 -4666 -590 -4596
rect -570 -4666 -566 -4596
rect -546 -4666 -542 -4596
rect -522 -4666 -518 -4596
rect -498 -4666 -494 -4596
rect -474 -4666 -470 -4596
rect -450 -4666 -446 -4596
rect -426 -4666 -422 -4596
rect -402 -4666 -398 -4596
rect -378 -4666 -374 -4596
rect -371 -4597 -357 -4596
rect -354 -4597 -347 -4573
rect -354 -4666 -350 -4597
rect -330 -4666 -326 -4572
rect -306 -4666 -302 -4572
rect -282 -4666 -278 -4572
rect -258 -4666 -254 -4572
rect -234 -4666 -230 -4572
rect -210 -4666 -206 -4572
rect -186 -4666 -182 -4572
rect -162 -4666 -158 -4572
rect -138 -4666 -134 -4572
rect -114 -4666 -110 -4572
rect -90 -4666 -86 -4572
rect -66 -4666 -62 -4572
rect -42 -4666 -38 -4572
rect -18 -4666 -14 -4572
rect 6 -4666 10 -4572
rect 30 -4666 34 -4572
rect 54 -4666 58 -4572
rect 78 -4666 82 -4572
rect 102 -4666 106 -4572
rect 115 -4579 120 -4572
rect 126 -4579 130 -4572
rect 125 -4593 130 -4579
rect 115 -4603 120 -4593
rect 125 -4617 130 -4603
rect 126 -4665 130 -4617
rect 115 -4666 147 -4665
rect -1181 -4668 147 -4666
rect -1181 -4675 -1176 -4668
rect -1171 -4689 -1166 -4675
rect -1170 -4690 -1166 -4689
rect -1146 -4690 -1142 -4668
rect -1122 -4690 -1118 -4668
rect -1098 -4690 -1094 -4668
rect -1074 -4690 -1070 -4668
rect -1050 -4690 -1046 -4668
rect -1026 -4690 -1022 -4668
rect -1002 -4690 -998 -4668
rect -978 -4690 -974 -4668
rect -954 -4690 -950 -4668
rect -930 -4690 -926 -4668
rect -906 -4690 -902 -4668
rect -882 -4690 -878 -4668
rect -858 -4690 -854 -4668
rect -834 -4690 -830 -4668
rect -810 -4690 -806 -4668
rect -786 -4690 -782 -4668
rect -762 -4690 -758 -4668
rect -738 -4690 -734 -4668
rect -714 -4690 -710 -4668
rect -701 -4690 -667 -4689
rect -2393 -4692 -667 -4690
rect -2371 -4738 -2366 -4692
rect -2348 -4738 -2343 -4692
rect -2325 -4738 -2320 -4692
rect -2309 -4708 -2301 -4698
rect -2317 -4714 -2309 -4708
rect -2097 -4714 -2095 -4705
rect -2309 -4736 -2301 -4726
rect -2097 -4728 -2095 -4724
rect -2292 -4729 -2095 -4728
rect -2097 -4731 -2095 -4729
rect -2084 -4736 -2083 -4693
rect -2069 -4700 -2054 -4698
rect -2054 -4716 -2018 -4714
rect -2054 -4718 -2004 -4716
rect -2059 -4722 -2045 -4718
rect -2054 -4724 -2049 -4722
rect -2317 -4738 -2309 -4736
rect -2084 -4738 -2054 -4736
rect -2044 -4738 -2039 -4724
rect -2025 -4734 -2014 -4728
rect -2000 -4734 -1992 -4692
rect -1920 -4694 -1906 -4692
rect -1977 -4709 -1929 -4703
rect -1655 -4708 -1647 -4698
rect -1977 -4719 -1966 -4709
rect -1663 -4714 -1655 -4708
rect -1977 -4731 -1929 -4729
rect -2033 -4738 -1992 -4734
rect -1655 -4736 -1647 -4726
rect -1663 -4738 -1655 -4736
rect -1642 -4738 -1637 -4692
rect -1619 -4738 -1614 -4692
rect -1530 -4738 -1526 -4692
rect -1506 -4738 -1502 -4692
rect -1482 -4738 -1478 -4692
rect -1458 -4738 -1454 -4692
rect -1434 -4738 -1430 -4692
rect -1410 -4738 -1406 -4692
rect -1386 -4738 -1382 -4692
rect -1362 -4738 -1358 -4692
rect -1338 -4738 -1334 -4692
rect -1314 -4738 -1310 -4692
rect -1290 -4738 -1286 -4692
rect -1266 -4738 -1262 -4692
rect -1242 -4738 -1238 -4692
rect -1218 -4738 -1214 -4692
rect -1194 -4738 -1190 -4692
rect -1170 -4738 -1166 -4692
rect -1146 -4693 -1142 -4692
rect -1146 -4717 -1139 -4693
rect -1122 -4738 -1118 -4692
rect -1098 -4738 -1094 -4692
rect -1074 -4738 -1070 -4692
rect -1050 -4738 -1046 -4692
rect -1026 -4738 -1022 -4692
rect -1002 -4738 -998 -4692
rect -978 -4738 -974 -4692
rect -954 -4738 -950 -4692
rect -930 -4738 -926 -4692
rect -906 -4738 -902 -4692
rect -882 -4738 -878 -4692
rect -858 -4738 -854 -4692
rect -834 -4738 -830 -4692
rect -810 -4738 -806 -4692
rect -786 -4738 -782 -4692
rect -762 -4738 -758 -4692
rect -738 -4737 -734 -4692
rect -749 -4738 -715 -4737
rect -2393 -4740 -715 -4738
rect -2371 -4858 -2366 -4740
rect -2348 -4858 -2343 -4740
rect -2325 -4774 -2320 -4740
rect -2317 -4742 -2309 -4740
rect -2084 -4753 -2083 -4740
rect -2084 -4754 -2054 -4753
rect -2325 -4782 -2317 -4774
rect -2325 -4802 -2320 -4782
rect -2317 -4790 -2309 -4782
rect -2117 -4791 -2095 -4781
rect -2045 -4784 -2037 -4770
rect -2325 -4818 -2317 -4802
rect -2325 -4834 -2320 -4818
rect -2309 -4830 -2301 -4818
rect -2317 -4834 -2309 -4830
rect -2117 -4832 -2095 -4825
rect -2069 -4826 -2041 -4818
rect -2017 -4820 -2015 -4818
rect -2325 -4846 -2317 -4834
rect -2125 -4841 -2095 -4834
rect -2047 -4836 -2011 -4834
rect -2059 -4838 -2011 -4836
rect -2000 -4838 -1992 -4740
rect -1663 -4742 -1655 -4740
rect -1969 -4791 -1929 -4779
rect -1671 -4782 -1663 -4774
rect -1663 -4790 -1655 -4782
rect -1671 -4818 -1663 -4802
rect -1655 -4830 -1647 -4818
rect -1663 -4834 -1655 -4830
rect -2125 -4843 -2117 -4841
rect -2059 -4842 -2045 -4838
rect -2021 -4841 -1992 -4838
rect -1977 -4841 -1929 -4834
rect -2325 -4858 -2320 -4846
rect -2309 -4858 -2301 -4846
rect -2131 -4851 -2129 -4846
rect -2125 -4849 -2095 -4843
rect -2021 -4848 -2009 -4844
rect -2125 -4851 -2117 -4849
rect -2133 -4858 -2129 -4851
rect -2117 -4858 -2087 -4851
rect -2025 -4854 -2021 -4848
rect -2000 -4854 -1992 -4841
rect -1969 -4849 -1929 -4843
rect -1671 -4846 -1663 -4834
rect -2033 -4858 -1992 -4854
rect -1969 -4858 -1921 -4851
rect -1655 -4858 -1647 -4846
rect -1642 -4858 -1637 -4740
rect -1619 -4858 -1614 -4740
rect -1530 -4858 -1526 -4740
rect -1506 -4858 -1502 -4740
rect -1482 -4858 -1478 -4740
rect -1458 -4858 -1454 -4740
rect -1434 -4858 -1430 -4740
rect -1410 -4858 -1406 -4740
rect -1386 -4858 -1382 -4740
rect -1362 -4858 -1358 -4740
rect -1338 -4858 -1334 -4740
rect -1314 -4858 -1310 -4740
rect -1290 -4858 -1286 -4740
rect -1266 -4858 -1262 -4740
rect -1242 -4858 -1238 -4740
rect -1218 -4858 -1214 -4740
rect -1194 -4858 -1190 -4740
rect -1170 -4858 -1166 -4740
rect -1146 -4762 -1139 -4741
rect -1122 -4762 -1118 -4740
rect -1098 -4762 -1094 -4740
rect -1074 -4762 -1070 -4740
rect -1050 -4762 -1046 -4740
rect -1026 -4762 -1022 -4740
rect -1002 -4762 -998 -4740
rect -978 -4761 -974 -4740
rect -989 -4762 -955 -4761
rect -1163 -4764 -955 -4762
rect -1163 -4765 -1149 -4764
rect -1146 -4765 -1139 -4764
rect -1146 -4858 -1142 -4765
rect -1122 -4858 -1118 -4764
rect -1098 -4857 -1094 -4764
rect -1109 -4858 -1075 -4857
rect -2393 -4860 -1075 -4858
rect -2371 -4954 -2366 -4860
rect -2348 -4954 -2343 -4860
rect -2325 -4862 -2320 -4860
rect -2317 -4862 -2309 -4860
rect -2131 -4862 -2129 -4860
rect -2125 -4862 -2095 -4860
rect -2325 -4874 -2317 -4862
rect -2117 -4867 -2095 -4862
rect -2325 -4894 -2320 -4874
rect -2325 -4902 -2317 -4894
rect -2325 -4922 -2320 -4902
rect -2317 -4910 -2309 -4902
rect -2117 -4911 -2095 -4901
rect -2045 -4904 -2037 -4890
rect -2325 -4936 -2317 -4922
rect -2325 -4952 -2320 -4936
rect -2317 -4938 -2309 -4936
rect -2309 -4950 -2301 -4938
rect -2109 -4939 -2079 -4938
rect -2317 -4952 -2309 -4950
rect -2325 -4954 -2317 -4952
rect -2109 -4953 -2087 -4939
rect -2015 -4952 -2001 -4947
rect -2000 -4952 -1992 -4860
rect -1663 -4862 -1655 -4860
rect -1671 -4874 -1663 -4862
rect -1969 -4911 -1929 -4899
rect -1671 -4902 -1663 -4894
rect -1663 -4910 -1655 -4902
rect -1671 -4936 -1663 -4922
rect -1663 -4938 -1655 -4936
rect -1655 -4950 -1647 -4938
rect -1663 -4952 -1655 -4950
rect -2109 -4954 -2079 -4953
rect -2033 -4954 -1992 -4952
rect -1864 -4954 -1680 -4953
rect -1671 -4954 -1663 -4952
rect -1642 -4954 -1637 -4860
rect -1619 -4954 -1614 -4860
rect -1530 -4954 -1526 -4860
rect -1506 -4954 -1502 -4860
rect -1482 -4954 -1478 -4860
rect -1458 -4954 -1454 -4860
rect -1434 -4954 -1430 -4860
rect -1410 -4954 -1406 -4860
rect -1386 -4954 -1382 -4860
rect -1362 -4954 -1358 -4860
rect -1338 -4954 -1334 -4860
rect -1314 -4954 -1310 -4860
rect -1290 -4954 -1286 -4860
rect -1266 -4954 -1262 -4860
rect -1242 -4953 -1238 -4860
rect -1253 -4954 -1219 -4953
rect -2393 -4956 -1219 -4954
rect -2371 -4978 -2366 -4956
rect -2348 -4978 -2343 -4956
rect -2325 -4964 -2317 -4956
rect -2109 -4961 -2087 -4956
rect -2117 -4963 -2085 -4961
rect -2325 -4978 -2320 -4964
rect -2317 -4966 -2309 -4964
rect -2309 -4978 -2301 -4966
rect -2023 -4973 -2021 -4964
rect -2037 -4974 -2021 -4973
rect -2051 -4976 -2021 -4974
rect -2074 -4978 -2021 -4976
rect -2000 -4978 -1992 -4956
rect -1969 -4963 -1921 -4961
rect -1671 -4964 -1663 -4956
rect -1663 -4966 -1655 -4964
rect -1655 -4978 -1647 -4966
rect -1642 -4978 -1637 -4956
rect -1619 -4978 -1614 -4956
rect -1530 -4978 -1526 -4956
rect -1506 -4978 -1502 -4956
rect -1482 -4978 -1478 -4956
rect -1458 -4978 -1454 -4956
rect -1434 -4978 -1430 -4956
rect -1410 -4978 -1406 -4956
rect -1386 -4978 -1382 -4956
rect -1362 -4978 -1358 -4956
rect -1338 -4978 -1334 -4956
rect -1314 -4978 -1310 -4956
rect -1290 -4978 -1286 -4956
rect -1266 -4978 -1262 -4956
rect -1253 -4963 -1248 -4956
rect -1242 -4963 -1238 -4956
rect -1243 -4977 -1238 -4963
rect -1242 -4978 -1238 -4977
rect -1218 -4978 -1214 -4860
rect -1194 -4978 -1190 -4860
rect -1170 -4978 -1166 -4860
rect -1146 -4978 -1142 -4860
rect -1122 -4978 -1118 -4860
rect -1109 -4867 -1104 -4860
rect -1098 -4867 -1094 -4860
rect -1099 -4881 -1094 -4867
rect -1109 -4906 -1075 -4905
rect -1074 -4906 -1070 -4764
rect -1050 -4906 -1046 -4764
rect -1026 -4906 -1022 -4764
rect -1013 -4891 -1008 -4881
rect -1002 -4891 -998 -4764
rect -989 -4771 -984 -4764
rect -978 -4771 -974 -4764
rect -979 -4785 -974 -4771
rect -989 -4786 -955 -4785
rect -954 -4786 -950 -4740
rect -930 -4786 -926 -4740
rect -906 -4786 -902 -4740
rect -882 -4786 -878 -4740
rect -858 -4786 -854 -4740
rect -834 -4786 -830 -4740
rect -810 -4786 -806 -4740
rect -786 -4786 -782 -4740
rect -762 -4786 -758 -4740
rect -749 -4747 -744 -4740
rect -738 -4747 -734 -4740
rect -739 -4761 -734 -4747
rect -738 -4786 -734 -4761
rect -714 -4786 -710 -4692
rect -701 -4699 -696 -4692
rect -691 -4713 -686 -4699
rect -690 -4786 -686 -4713
rect -666 -4717 -662 -4668
rect -666 -4741 -659 -4717
rect -989 -4788 -669 -4786
rect -989 -4795 -984 -4788
rect -979 -4809 -974 -4795
rect -1003 -4905 -998 -4891
rect -978 -4906 -974 -4809
rect -954 -4837 -950 -4788
rect -954 -4885 -947 -4837
rect -954 -4906 -950 -4885
rect -930 -4906 -926 -4788
rect -906 -4906 -902 -4788
rect -882 -4906 -878 -4788
rect -858 -4906 -854 -4788
rect -834 -4906 -830 -4788
rect -810 -4906 -806 -4788
rect -786 -4906 -782 -4788
rect -762 -4906 -758 -4788
rect -738 -4906 -734 -4788
rect -714 -4813 -710 -4788
rect -714 -4837 -707 -4813
rect -714 -4906 -710 -4837
rect -690 -4906 -686 -4788
rect -683 -4789 -669 -4788
rect -666 -4789 -659 -4765
rect -666 -4906 -662 -4789
rect -642 -4906 -638 -4668
rect -618 -4906 -614 -4668
rect -594 -4906 -590 -4668
rect -570 -4906 -566 -4668
rect -546 -4906 -542 -4668
rect -522 -4906 -518 -4668
rect -498 -4906 -494 -4668
rect -474 -4906 -470 -4668
rect -450 -4906 -446 -4668
rect -426 -4906 -422 -4668
rect -402 -4906 -398 -4668
rect -378 -4906 -374 -4668
rect -354 -4906 -350 -4668
rect -330 -4906 -326 -4668
rect -306 -4906 -302 -4668
rect -282 -4906 -278 -4668
rect -258 -4906 -254 -4668
rect -234 -4906 -230 -4668
rect -210 -4906 -206 -4668
rect -186 -4906 -182 -4668
rect -162 -4906 -158 -4668
rect -138 -4906 -134 -4668
rect -114 -4906 -110 -4668
rect -90 -4906 -86 -4668
rect -66 -4906 -62 -4668
rect -42 -4906 -38 -4668
rect -18 -4906 -14 -4668
rect 6 -4906 10 -4668
rect 30 -4906 34 -4668
rect 54 -4906 58 -4668
rect 78 -4906 82 -4668
rect 91 -4795 96 -4785
rect 102 -4795 106 -4668
rect 115 -4675 120 -4668
rect 126 -4675 130 -4668
rect 133 -4669 147 -4668
rect 125 -4689 130 -4675
rect 139 -4679 147 -4675
rect 133 -4689 139 -4679
rect 101 -4809 106 -4795
rect 91 -4819 96 -4809
rect 101 -4833 106 -4819
rect 102 -4905 106 -4833
rect 91 -4906 123 -4905
rect -1109 -4908 123 -4906
rect -1109 -4915 -1104 -4908
rect -1099 -4929 -1094 -4915
rect -1098 -4978 -1094 -4929
rect -1074 -4933 -1070 -4908
rect -1074 -4957 -1067 -4933
rect -1050 -4978 -1046 -4908
rect -1026 -4978 -1022 -4908
rect -1013 -4963 -1008 -4953
rect -978 -4957 -974 -4908
rect -1003 -4977 -998 -4963
rect -989 -4967 -981 -4963
rect -995 -4977 -989 -4967
rect -1002 -4978 -998 -4977
rect -2393 -4980 -981 -4978
rect -2371 -5026 -2366 -4980
rect -2348 -5026 -2343 -4980
rect -2325 -4992 -2317 -4980
rect -2117 -4987 -2087 -4983
rect -2325 -5012 -2320 -4992
rect -2317 -4994 -2309 -4992
rect -2325 -5020 -2317 -5012
rect -2101 -5017 -2071 -5014
rect -2325 -5026 -2320 -5020
rect -2317 -5026 -2309 -5020
rect -2000 -5022 -1992 -4980
rect -1969 -4987 -1921 -4983
rect -1864 -4987 -1680 -4982
rect -1671 -4992 -1663 -4980
rect -1663 -4994 -1655 -4992
rect -1854 -5008 -1680 -5004
rect -1846 -5017 -1798 -5014
rect -2079 -5023 -2043 -5022
rect -2007 -5023 -1991 -5022
rect -2079 -5024 -2071 -5023
rect -2079 -5026 -2029 -5024
rect -2011 -5026 -1991 -5023
rect -1846 -5025 -1806 -5019
rect -1671 -5020 -1663 -5012
rect -1864 -5026 -1796 -5025
rect -1663 -5026 -1655 -5020
rect -1642 -5026 -1637 -4980
rect -1619 -5026 -1614 -4980
rect -1530 -5026 -1526 -4980
rect -1506 -5026 -1502 -4980
rect -1482 -5026 -1478 -4980
rect -1458 -5026 -1454 -4980
rect -1434 -5026 -1430 -4980
rect -1410 -5026 -1406 -4980
rect -1386 -5026 -1382 -4980
rect -1362 -5026 -1358 -4980
rect -1338 -5025 -1334 -4980
rect -1349 -5026 -1315 -5025
rect -2393 -5028 -1315 -5026
rect -2371 -5074 -2366 -5028
rect -2348 -5074 -2343 -5028
rect -2325 -5040 -2320 -5028
rect -2079 -5030 -2071 -5028
rect -2072 -5032 -2071 -5030
rect -2109 -5037 -2101 -5032
rect -2101 -5039 -2079 -5037
rect -2069 -5039 -2068 -5032
rect -2325 -5048 -2317 -5040
rect -2079 -5044 -2071 -5039
rect -2325 -5068 -2320 -5048
rect -2317 -5056 -2309 -5048
rect -2074 -5053 -2071 -5044
rect -2069 -5048 -2068 -5044
rect -2109 -5062 -2079 -5059
rect -2325 -5074 -2317 -5068
rect -2000 -5074 -1992 -5028
rect -1846 -5030 -1806 -5028
rect -1854 -5035 -1806 -5031
rect -1854 -5037 -1846 -5035
rect -1846 -5039 -1806 -5037
rect -1806 -5041 -1798 -5039
rect -1846 -5044 -1798 -5041
rect -1846 -5057 -1806 -5046
rect -1671 -5048 -1663 -5040
rect -1663 -5056 -1655 -5048
rect -1854 -5062 -1680 -5058
rect -1671 -5074 -1663 -5068
rect -1642 -5074 -1637 -5028
rect -1619 -5074 -1614 -5028
rect -1530 -5074 -1526 -5028
rect -1506 -5074 -1502 -5028
rect -1482 -5074 -1478 -5028
rect -1458 -5074 -1454 -5028
rect -1434 -5074 -1430 -5028
rect -1410 -5074 -1406 -5028
rect -1386 -5074 -1382 -5028
rect -1362 -5074 -1358 -5028
rect -1349 -5035 -1344 -5028
rect -1338 -5035 -1334 -5028
rect -1339 -5049 -1334 -5035
rect -1349 -5050 -1315 -5049
rect -1314 -5050 -1310 -4980
rect -1290 -5050 -1286 -4980
rect -1266 -5050 -1262 -4980
rect -1242 -5050 -1238 -4980
rect -1218 -5029 -1214 -4980
rect -1349 -5052 -1221 -5050
rect -1349 -5059 -1344 -5052
rect -1339 -5073 -1334 -5059
rect -1338 -5074 -1334 -5073
rect -1314 -5074 -1310 -5052
rect -1290 -5074 -1286 -5052
rect -1266 -5074 -1262 -5052
rect -1242 -5074 -1238 -5052
rect -1235 -5053 -1221 -5052
rect -1218 -5053 -1211 -5029
rect -1218 -5074 -1214 -5053
rect -1194 -5074 -1190 -4980
rect -1170 -5074 -1166 -4980
rect -1146 -5074 -1142 -4980
rect -1122 -5074 -1118 -4980
rect -1098 -5074 -1094 -4980
rect -1074 -5002 -1067 -4981
rect -1050 -5002 -1046 -4980
rect -1026 -5002 -1022 -4980
rect -1002 -5002 -998 -4980
rect -995 -4981 -981 -4980
rect -978 -4981 -971 -4957
rect -954 -5002 -950 -4908
rect -930 -5002 -926 -4908
rect -906 -5002 -902 -4908
rect -882 -5002 -878 -4908
rect -858 -5002 -854 -4908
rect -834 -5002 -830 -4908
rect -810 -5002 -806 -4908
rect -786 -5002 -782 -4908
rect -762 -5002 -758 -4908
rect -738 -5002 -734 -4908
rect -714 -5002 -710 -4908
rect -690 -5002 -686 -4908
rect -666 -5002 -662 -4908
rect -642 -5002 -638 -4908
rect -618 -5002 -614 -4908
rect -594 -5002 -590 -4908
rect -570 -5002 -566 -4908
rect -557 -4987 -552 -4977
rect -546 -4987 -542 -4908
rect -547 -5001 -542 -4987
rect -522 -5002 -518 -4908
rect -498 -5002 -494 -4908
rect -474 -5002 -470 -4908
rect -450 -5002 -446 -4908
rect -426 -5002 -422 -4908
rect -402 -5002 -398 -4908
rect -378 -5002 -374 -4908
rect -354 -5002 -350 -4908
rect -330 -5002 -326 -4908
rect -306 -5002 -302 -4908
rect -282 -5002 -278 -4908
rect -269 -4939 -264 -4929
rect -258 -4939 -254 -4908
rect -259 -4953 -254 -4939
rect -269 -4987 -264 -4977
rect -259 -5001 -254 -4987
rect -234 -5001 -230 -4908
rect -258 -5002 -254 -5001
rect -245 -5002 -211 -5001
rect -1091 -5004 -211 -5002
rect -1091 -5005 -1077 -5004
rect -1074 -5005 -1067 -5004
rect -1074 -5074 -1070 -5005
rect -1050 -5074 -1046 -5004
rect -1026 -5074 -1022 -5004
rect -1002 -5074 -998 -5004
rect -978 -5050 -971 -5029
rect -954 -5050 -950 -5004
rect -930 -5050 -926 -5004
rect -906 -5050 -902 -5004
rect -882 -5050 -878 -5004
rect -858 -5050 -854 -5004
rect -834 -5050 -830 -5004
rect -810 -5050 -806 -5004
rect -786 -5050 -782 -5004
rect -762 -5050 -758 -5004
rect -738 -5050 -734 -5004
rect -714 -5050 -710 -5004
rect -690 -5050 -686 -5004
rect -666 -5050 -662 -5004
rect -642 -5050 -638 -5004
rect -618 -5050 -614 -5004
rect -594 -5050 -590 -5004
rect -570 -5050 -566 -5004
rect -557 -5026 -523 -5025
rect -522 -5026 -518 -5004
rect -498 -5026 -494 -5004
rect -474 -5026 -470 -5004
rect -450 -5026 -446 -5004
rect -426 -5026 -422 -5004
rect -402 -5026 -398 -5004
rect -378 -5026 -374 -5004
rect -354 -5026 -350 -5004
rect -330 -5026 -326 -5004
rect -306 -5026 -302 -5004
rect -282 -5026 -278 -5004
rect -258 -5026 -254 -5004
rect -245 -5011 -240 -5004
rect -234 -5005 -230 -5004
rect -234 -5011 -227 -5005
rect -235 -5025 -227 -5011
rect -557 -5028 -237 -5026
rect -557 -5035 -552 -5028
rect -547 -5049 -542 -5035
rect -546 -5050 -542 -5049
rect -522 -5050 -518 -5028
rect -498 -5050 -494 -5028
rect -474 -5050 -470 -5028
rect -450 -5050 -446 -5028
rect -426 -5050 -422 -5028
rect -402 -5050 -398 -5028
rect -378 -5050 -374 -5028
rect -354 -5050 -350 -5028
rect -330 -5050 -326 -5028
rect -306 -5050 -302 -5028
rect -282 -5050 -278 -5028
rect -258 -5050 -254 -5028
rect -251 -5029 -237 -5028
rect -210 -5050 -206 -4908
rect -186 -5050 -182 -4908
rect -162 -5050 -158 -4908
rect -138 -5050 -134 -4908
rect -114 -5050 -110 -4908
rect -90 -5050 -86 -4908
rect -66 -5050 -62 -4908
rect -42 -5050 -38 -4908
rect -18 -5050 -14 -4908
rect 6 -5049 10 -4908
rect 19 -5035 24 -5025
rect 30 -5035 34 -4908
rect 43 -4987 48 -4977
rect 54 -4987 58 -4908
rect 67 -4963 72 -4953
rect 78 -4963 82 -4908
rect 91 -4915 96 -4908
rect 102 -4915 106 -4908
rect 109 -4909 123 -4908
rect 101 -4929 106 -4915
rect 77 -4977 82 -4963
rect 53 -5001 58 -4987
rect 29 -5049 34 -5035
rect -5 -5050 29 -5049
rect -995 -5052 29 -5050
rect -995 -5053 -981 -5052
rect -978 -5053 -971 -5052
rect -978 -5074 -974 -5053
rect -954 -5073 -950 -5052
rect -965 -5074 -931 -5073
rect -2393 -5076 -931 -5074
rect -2371 -5098 -2366 -5076
rect -2348 -5098 -2343 -5076
rect -2325 -5084 -2317 -5076
rect -2325 -5098 -2320 -5084
rect -2309 -5096 -2301 -5084
rect -2092 -5093 -2062 -5088
rect -2000 -5096 -1992 -5076
rect -2317 -5098 -2309 -5096
rect -2000 -5098 -1983 -5096
rect -1906 -5098 -1904 -5076
rect -1806 -5084 -1680 -5078
rect -1671 -5084 -1663 -5076
rect -1854 -5093 -1806 -5088
rect -1846 -5098 -1806 -5095
rect -1655 -5096 -1647 -5084
rect -1663 -5098 -1655 -5096
rect -1642 -5098 -1637 -5076
rect -1619 -5098 -1614 -5076
rect -1530 -5098 -1526 -5076
rect -1506 -5098 -1502 -5076
rect -1482 -5098 -1478 -5076
rect -1458 -5098 -1454 -5076
rect -1434 -5098 -1430 -5076
rect -1410 -5098 -1406 -5076
rect -1386 -5098 -1382 -5076
rect -1362 -5098 -1358 -5076
rect -1338 -5098 -1334 -5076
rect -1314 -5098 -1310 -5076
rect -1290 -5098 -1286 -5076
rect -1266 -5098 -1262 -5076
rect -1242 -5098 -1238 -5076
rect -1218 -5098 -1214 -5076
rect -1194 -5098 -1190 -5076
rect -1170 -5098 -1166 -5076
rect -1146 -5097 -1142 -5076
rect -1157 -5098 -1123 -5097
rect -2393 -5100 -1123 -5098
rect -2371 -5122 -2366 -5100
rect -2348 -5122 -2343 -5100
rect -2325 -5112 -2317 -5100
rect -2071 -5104 -2062 -5100
rect -2013 -5102 -1983 -5100
rect -2000 -5103 -1983 -5102
rect -2325 -5122 -2320 -5112
rect -2309 -5122 -2301 -5112
rect -2100 -5113 -2092 -5106
rect -2064 -5108 -2062 -5105
rect -2061 -5113 -2059 -5108
rect -2071 -5118 -2062 -5113
rect -2071 -5120 -2026 -5118
rect -2066 -5122 -2012 -5120
rect -2000 -5122 -1992 -5103
rect -1906 -5105 -1904 -5100
rect -1846 -5104 -1806 -5100
rect -1846 -5111 -1798 -5106
rect -1806 -5113 -1798 -5111
rect -1671 -5112 -1663 -5100
rect -1854 -5115 -1846 -5113
rect -1854 -5120 -1806 -5115
rect -1864 -5122 -1796 -5121
rect -1655 -5122 -1647 -5112
rect -1642 -5122 -1637 -5100
rect -1619 -5122 -1614 -5100
rect -1530 -5122 -1526 -5100
rect -1506 -5122 -1502 -5100
rect -1482 -5122 -1478 -5100
rect -1458 -5122 -1454 -5100
rect -1434 -5122 -1430 -5100
rect -1410 -5122 -1406 -5100
rect -1386 -5122 -1382 -5100
rect -1362 -5122 -1358 -5100
rect -1338 -5122 -1334 -5100
rect -1314 -5101 -1310 -5100
rect -2393 -5124 -1317 -5122
rect -2371 -5170 -2366 -5124
rect -2348 -5170 -2343 -5124
rect -2325 -5128 -2320 -5124
rect -2317 -5128 -2309 -5124
rect -2325 -5140 -2317 -5128
rect -2066 -5129 -2062 -5124
rect -2147 -5132 -2134 -5130
rect -2292 -5138 -2071 -5132
rect -2325 -5160 -2320 -5140
rect -2092 -5154 -2062 -5152
rect -2094 -5158 -2062 -5154
rect -2325 -5170 -2317 -5160
rect -2095 -5168 -2084 -5164
rect -2000 -5167 -1992 -5124
rect -1846 -5131 -1806 -5124
rect -1663 -5128 -1655 -5124
rect -1846 -5138 -1680 -5132
rect -1671 -5140 -1663 -5128
rect -1854 -5154 -1806 -5152
rect -1854 -5158 -1680 -5154
rect -2119 -5170 -2069 -5168
rect -2054 -5170 -1892 -5167
rect -1671 -5170 -1663 -5160
rect -1642 -5170 -1637 -5124
rect -1619 -5170 -1614 -5124
rect -1530 -5170 -1526 -5124
rect -1506 -5170 -1502 -5124
rect -1482 -5170 -1478 -5124
rect -1458 -5170 -1454 -5124
rect -1434 -5170 -1430 -5124
rect -1410 -5170 -1406 -5124
rect -1386 -5170 -1382 -5124
rect -1362 -5170 -1358 -5124
rect -1338 -5170 -1334 -5124
rect -1331 -5125 -1317 -5124
rect -1314 -5149 -1307 -5101
rect -1314 -5170 -1310 -5149
rect -1290 -5170 -1286 -5100
rect -1266 -5170 -1262 -5100
rect -1242 -5170 -1238 -5100
rect -1218 -5170 -1214 -5100
rect -1194 -5170 -1190 -5100
rect -1170 -5170 -1166 -5100
rect -1157 -5107 -1152 -5100
rect -1146 -5107 -1142 -5100
rect -1147 -5121 -1142 -5107
rect -1157 -5146 -1123 -5145
rect -1122 -5146 -1118 -5076
rect -1098 -5146 -1094 -5076
rect -1074 -5146 -1070 -5076
rect -1050 -5146 -1046 -5076
rect -1026 -5146 -1022 -5076
rect -1002 -5146 -998 -5076
rect -978 -5146 -974 -5076
rect -965 -5083 -960 -5076
rect -954 -5083 -950 -5076
rect -955 -5097 -950 -5083
rect -965 -5098 -931 -5097
rect -930 -5098 -926 -5052
rect -906 -5098 -902 -5052
rect -882 -5098 -878 -5052
rect -858 -5098 -854 -5052
rect -834 -5098 -830 -5052
rect -810 -5098 -806 -5052
rect -786 -5098 -782 -5052
rect -762 -5098 -758 -5052
rect -738 -5098 -734 -5052
rect -714 -5098 -710 -5052
rect -690 -5098 -686 -5052
rect -666 -5098 -662 -5052
rect -642 -5098 -638 -5052
rect -618 -5098 -614 -5052
rect -594 -5098 -590 -5052
rect -570 -5098 -566 -5052
rect -546 -5098 -542 -5052
rect -522 -5053 -518 -5052
rect -522 -5077 -515 -5053
rect -498 -5098 -494 -5052
rect -474 -5098 -470 -5052
rect -450 -5098 -446 -5052
rect -426 -5098 -422 -5052
rect -402 -5098 -398 -5052
rect -378 -5098 -374 -5052
rect -354 -5098 -350 -5052
rect -330 -5098 -326 -5052
rect -306 -5098 -302 -5052
rect -282 -5098 -278 -5052
rect -258 -5098 -254 -5052
rect -245 -5074 -211 -5073
rect -210 -5074 -206 -5052
rect -186 -5074 -182 -5052
rect -162 -5074 -158 -5052
rect -138 -5074 -134 -5052
rect -114 -5074 -110 -5052
rect -90 -5074 -86 -5052
rect -66 -5074 -62 -5052
rect -42 -5074 -38 -5052
rect -18 -5073 -14 -5052
rect -5 -5059 0 -5052
rect 6 -5059 10 -5052
rect 5 -5073 10 -5059
rect -29 -5074 5 -5073
rect -245 -5076 5 -5074
rect -245 -5077 -237 -5076
rect -210 -5077 -206 -5076
rect -245 -5083 -240 -5077
rect -235 -5097 -230 -5083
rect -221 -5087 -213 -5083
rect -227 -5097 -221 -5087
rect -234 -5098 -230 -5097
rect -965 -5100 -213 -5098
rect -965 -5107 -960 -5100
rect -955 -5121 -950 -5107
rect -954 -5146 -950 -5121
rect -930 -5146 -926 -5100
rect -906 -5146 -902 -5100
rect -882 -5146 -878 -5100
rect -858 -5146 -854 -5100
rect -834 -5146 -830 -5100
rect -810 -5146 -806 -5100
rect -786 -5146 -782 -5100
rect -762 -5146 -758 -5100
rect -738 -5146 -734 -5100
rect -714 -5146 -710 -5100
rect -690 -5146 -686 -5100
rect -666 -5146 -662 -5100
rect -642 -5146 -638 -5100
rect -618 -5146 -614 -5100
rect -594 -5146 -590 -5100
rect -570 -5146 -566 -5100
rect -546 -5146 -542 -5100
rect -522 -5122 -515 -5101
rect -498 -5122 -494 -5100
rect -474 -5122 -470 -5100
rect -450 -5122 -446 -5100
rect -426 -5121 -422 -5100
rect -437 -5122 -403 -5121
rect -539 -5124 -403 -5122
rect -539 -5125 -525 -5124
rect -522 -5125 -515 -5124
rect -522 -5146 -518 -5125
rect -498 -5146 -494 -5124
rect -474 -5146 -470 -5124
rect -450 -5146 -446 -5124
rect -437 -5131 -432 -5124
rect -426 -5131 -422 -5124
rect -427 -5145 -422 -5131
rect -402 -5146 -398 -5100
rect -378 -5146 -374 -5100
rect -354 -5146 -350 -5100
rect -330 -5146 -326 -5100
rect -306 -5146 -302 -5100
rect -282 -5146 -278 -5100
rect -258 -5146 -254 -5100
rect -234 -5146 -230 -5100
rect -227 -5101 -213 -5100
rect -210 -5101 -203 -5077
rect -186 -5146 -182 -5076
rect -162 -5146 -158 -5076
rect -138 -5146 -134 -5076
rect -114 -5146 -110 -5076
rect -90 -5146 -86 -5076
rect -66 -5145 -62 -5076
rect -53 -5107 -48 -5097
rect -42 -5107 -38 -5076
rect -29 -5083 -24 -5076
rect -18 -5083 -14 -5076
rect -19 -5097 -14 -5083
rect -43 -5121 -38 -5107
rect -77 -5146 -43 -5145
rect -1157 -5148 -43 -5146
rect -1157 -5155 -1152 -5148
rect -1147 -5169 -1142 -5155
rect -1146 -5170 -1142 -5169
rect -1122 -5170 -1118 -5148
rect -1098 -5170 -1094 -5148
rect -1074 -5170 -1070 -5148
rect -1050 -5170 -1046 -5148
rect -1026 -5170 -1022 -5148
rect -1002 -5170 -998 -5148
rect -978 -5170 -974 -5148
rect -954 -5170 -950 -5148
rect -930 -5149 -926 -5148
rect -2393 -5172 -933 -5170
rect -2371 -5194 -2366 -5172
rect -2348 -5194 -2343 -5172
rect -2325 -5176 -2317 -5172
rect -2325 -5192 -2320 -5176
rect -2309 -5188 -2301 -5176
rect -2095 -5178 -2084 -5172
rect -2054 -5173 -1906 -5172
rect -2054 -5174 -2036 -5173
rect -2084 -5180 -2079 -5178
rect -2317 -5192 -2309 -5188
rect -2092 -5189 -2079 -5182
rect -2000 -5186 -1992 -5173
rect -1920 -5174 -1906 -5173
rect -1671 -5176 -1663 -5172
rect -1846 -5180 -1806 -5178
rect -1854 -5186 -1806 -5182
rect -2054 -5189 -1982 -5186
rect -1966 -5189 -1806 -5186
rect -1655 -5188 -1647 -5176
rect -2003 -5192 -1992 -5189
rect -1904 -5191 -1902 -5189
rect -1854 -5191 -1846 -5189
rect -2325 -5194 -2317 -5192
rect -2033 -5194 -1992 -5192
rect -1854 -5193 -1806 -5191
rect -1663 -5192 -1655 -5188
rect -1864 -5194 -1796 -5193
rect -1671 -5194 -1663 -5192
rect -1642 -5194 -1637 -5172
rect -1619 -5194 -1614 -5172
rect -1530 -5194 -1526 -5172
rect -1506 -5194 -1502 -5172
rect -1482 -5194 -1478 -5172
rect -1458 -5194 -1454 -5172
rect -1434 -5194 -1430 -5172
rect -1410 -5194 -1406 -5172
rect -1386 -5194 -1382 -5172
rect -1362 -5194 -1358 -5172
rect -1338 -5193 -1334 -5172
rect -1349 -5194 -1315 -5193
rect -2393 -5196 -1315 -5194
rect -2371 -5218 -2366 -5196
rect -2348 -5218 -2343 -5196
rect -2325 -5204 -2317 -5196
rect -2079 -5199 -2018 -5196
rect -2003 -5197 -1966 -5196
rect -2000 -5198 -1982 -5197
rect -2000 -5199 -1992 -5198
rect -2084 -5203 -2009 -5199
rect -2028 -5204 -2009 -5203
rect -2000 -5203 -1854 -5199
rect -1846 -5203 -1798 -5196
rect -2325 -5218 -2320 -5204
rect -2309 -5216 -2301 -5204
rect -2028 -5206 -2018 -5204
rect -2092 -5216 -2084 -5209
rect -2023 -5213 -2014 -5206
rect -2000 -5213 -1992 -5203
rect -1671 -5204 -1663 -5196
rect -1846 -5207 -1806 -5205
rect -1854 -5213 -1806 -5209
rect -2054 -5216 -1806 -5213
rect -1655 -5216 -1647 -5204
rect -2317 -5218 -2309 -5216
rect -2054 -5218 -2024 -5216
rect -2000 -5218 -1992 -5216
rect -1663 -5218 -1655 -5216
rect -1642 -5218 -1637 -5196
rect -1619 -5218 -1614 -5196
rect -1530 -5218 -1526 -5196
rect -1506 -5218 -1502 -5196
rect -1482 -5218 -1478 -5196
rect -1458 -5218 -1454 -5196
rect -1434 -5218 -1430 -5196
rect -1410 -5218 -1406 -5196
rect -1386 -5218 -1382 -5196
rect -1362 -5217 -1358 -5196
rect -1349 -5203 -1344 -5196
rect -1338 -5203 -1334 -5196
rect -1339 -5217 -1334 -5203
rect -1373 -5218 -1315 -5217
rect -1314 -5218 -1310 -5172
rect -1290 -5218 -1286 -5172
rect -1266 -5218 -1262 -5172
rect -1242 -5218 -1238 -5172
rect -1218 -5218 -1214 -5172
rect -1194 -5218 -1190 -5172
rect -1170 -5218 -1166 -5172
rect -1146 -5218 -1142 -5172
rect -1122 -5173 -1118 -5172
rect -1122 -5197 -1115 -5173
rect -1098 -5218 -1094 -5172
rect -1074 -5218 -1070 -5172
rect -1050 -5218 -1046 -5172
rect -1026 -5218 -1022 -5172
rect -1002 -5218 -998 -5172
rect -978 -5218 -974 -5172
rect -954 -5218 -950 -5172
rect -947 -5173 -933 -5172
rect -930 -5197 -923 -5149
rect -930 -5218 -926 -5197
rect -906 -5218 -902 -5148
rect -882 -5218 -878 -5148
rect -858 -5218 -854 -5148
rect -834 -5218 -830 -5148
rect -810 -5218 -806 -5148
rect -786 -5218 -782 -5148
rect -762 -5218 -758 -5148
rect -738 -5218 -734 -5148
rect -714 -5218 -710 -5148
rect -690 -5218 -686 -5148
rect -666 -5218 -662 -5148
rect -642 -5218 -638 -5148
rect -618 -5218 -614 -5148
rect -594 -5218 -590 -5148
rect -570 -5218 -566 -5148
rect -546 -5218 -542 -5148
rect -522 -5218 -518 -5148
rect -498 -5218 -494 -5148
rect -474 -5218 -470 -5148
rect -450 -5218 -446 -5148
rect -437 -5194 -403 -5193
rect -402 -5194 -398 -5148
rect -378 -5194 -374 -5148
rect -354 -5194 -350 -5148
rect -330 -5194 -326 -5148
rect -306 -5194 -302 -5148
rect -282 -5194 -278 -5148
rect -258 -5194 -254 -5148
rect -234 -5194 -230 -5148
rect -210 -5169 -203 -5149
rect -221 -5170 -187 -5169
rect -227 -5172 -187 -5170
rect -227 -5173 -213 -5172
rect -210 -5173 -203 -5172
rect -221 -5179 -216 -5173
rect -210 -5179 -206 -5173
rect -211 -5193 -206 -5179
rect -186 -5194 -182 -5148
rect -162 -5194 -158 -5148
rect -138 -5194 -134 -5148
rect -114 -5194 -110 -5148
rect -90 -5193 -86 -5148
rect -77 -5155 -72 -5148
rect -66 -5155 -62 -5148
rect -67 -5169 -62 -5155
rect -101 -5194 -67 -5193
rect -437 -5196 -67 -5194
rect -437 -5203 -432 -5196
rect -402 -5197 -398 -5196
rect -427 -5217 -422 -5203
rect -413 -5207 -405 -5203
rect -419 -5217 -413 -5207
rect -426 -5218 -422 -5217
rect -2393 -5220 -2064 -5218
rect -2060 -5220 -405 -5218
rect -2371 -5266 -2366 -5220
rect -2348 -5266 -2343 -5220
rect -2325 -5232 -2317 -5220
rect -2060 -5223 -2054 -5220
rect -2084 -5230 -2054 -5223
rect -2050 -5226 -2044 -5224
rect -2325 -5252 -2320 -5232
rect -2064 -5234 -2054 -5230
rect -2325 -5260 -2317 -5252
rect -2101 -5257 -2071 -5254
rect -2325 -5266 -2320 -5260
rect -2317 -5266 -2309 -5260
rect -2000 -5262 -1992 -5220
rect -1846 -5221 -1806 -5220
rect -1846 -5230 -1798 -5223
rect -1671 -5232 -1663 -5220
rect -1846 -5234 -1806 -5232
rect -1854 -5248 -1680 -5244
rect -1846 -5257 -1798 -5254
rect -2079 -5263 -2043 -5262
rect -2007 -5263 -1991 -5262
rect -2079 -5264 -2071 -5263
rect -2079 -5266 -2029 -5264
rect -2011 -5266 -1991 -5263
rect -1846 -5265 -1806 -5259
rect -1671 -5260 -1663 -5252
rect -1864 -5266 -1796 -5265
rect -1663 -5266 -1655 -5260
rect -1642 -5266 -1637 -5220
rect -1619 -5266 -1614 -5220
rect -1530 -5266 -1526 -5220
rect -1506 -5266 -1502 -5220
rect -1493 -5251 -1488 -5241
rect -1482 -5251 -1478 -5220
rect -1483 -5265 -1478 -5251
rect -1482 -5266 -1478 -5265
rect -1458 -5266 -1454 -5220
rect -1434 -5266 -1430 -5220
rect -1410 -5266 -1406 -5220
rect -1386 -5266 -1382 -5220
rect -1373 -5227 -1368 -5220
rect -1362 -5227 -1358 -5220
rect -1349 -5227 -1344 -5220
rect -1363 -5241 -1358 -5227
rect -1339 -5241 -1334 -5227
rect -1373 -5251 -1368 -5241
rect -1363 -5265 -1358 -5251
rect -1362 -5266 -1358 -5265
rect -1338 -5266 -1334 -5241
rect -1314 -5266 -1310 -5220
rect -1290 -5266 -1286 -5220
rect -1266 -5266 -1262 -5220
rect -1242 -5266 -1238 -5220
rect -1218 -5266 -1214 -5220
rect -1194 -5266 -1190 -5220
rect -1170 -5266 -1166 -5220
rect -1146 -5266 -1142 -5220
rect -1122 -5242 -1115 -5221
rect -1098 -5242 -1094 -5220
rect -1074 -5242 -1070 -5220
rect -1050 -5242 -1046 -5220
rect -1026 -5242 -1022 -5220
rect -1002 -5242 -998 -5220
rect -978 -5242 -974 -5220
rect -954 -5242 -950 -5220
rect -930 -5242 -926 -5220
rect -906 -5242 -902 -5220
rect -882 -5242 -878 -5220
rect -858 -5242 -854 -5220
rect -834 -5242 -830 -5220
rect -810 -5242 -806 -5220
rect -786 -5242 -782 -5220
rect -762 -5242 -758 -5220
rect -738 -5242 -734 -5220
rect -714 -5242 -710 -5220
rect -690 -5242 -686 -5220
rect -666 -5242 -662 -5220
rect -642 -5242 -638 -5220
rect -618 -5242 -614 -5220
rect -594 -5242 -590 -5220
rect -570 -5242 -566 -5220
rect -546 -5242 -542 -5220
rect -522 -5242 -518 -5220
rect -498 -5242 -494 -5220
rect -474 -5242 -470 -5220
rect -450 -5242 -446 -5220
rect -426 -5242 -422 -5220
rect -419 -5221 -405 -5220
rect -402 -5221 -395 -5197
rect -378 -5242 -374 -5196
rect -354 -5242 -350 -5196
rect -330 -5242 -326 -5196
rect -306 -5242 -302 -5196
rect -282 -5242 -278 -5196
rect -258 -5242 -254 -5196
rect -234 -5242 -230 -5196
rect -186 -5242 -182 -5196
rect -162 -5242 -158 -5196
rect -138 -5241 -134 -5196
rect -125 -5227 -120 -5217
rect -114 -5227 -110 -5196
rect -101 -5203 -96 -5196
rect -90 -5203 -86 -5196
rect -91 -5217 -86 -5203
rect -115 -5241 -110 -5227
rect -149 -5242 -115 -5241
rect -1139 -5244 -115 -5242
rect -1139 -5245 -1125 -5244
rect -1122 -5245 -1115 -5244
rect -1122 -5266 -1118 -5245
rect -1098 -5266 -1094 -5244
rect -1074 -5266 -1070 -5244
rect -1050 -5266 -1046 -5244
rect -1026 -5266 -1022 -5244
rect -1002 -5266 -998 -5244
rect -978 -5266 -974 -5244
rect -954 -5266 -950 -5244
rect -930 -5266 -926 -5244
rect -906 -5266 -902 -5244
rect -882 -5265 -878 -5244
rect -893 -5266 -859 -5265
rect -2393 -5268 -859 -5266
rect -2371 -5314 -2366 -5268
rect -2348 -5314 -2343 -5268
rect -2325 -5280 -2320 -5268
rect -2079 -5270 -2071 -5268
rect -2072 -5272 -2071 -5270
rect -2109 -5277 -2101 -5272
rect -2101 -5279 -2079 -5277
rect -2069 -5279 -2068 -5272
rect -2325 -5288 -2317 -5280
rect -2079 -5284 -2071 -5279
rect -2325 -5308 -2320 -5288
rect -2317 -5296 -2309 -5288
rect -2074 -5293 -2071 -5284
rect -2069 -5288 -2068 -5284
rect -2109 -5302 -2079 -5299
rect -2325 -5314 -2317 -5308
rect -2000 -5314 -1992 -5268
rect -1846 -5270 -1806 -5268
rect -1854 -5275 -1806 -5271
rect -1854 -5277 -1846 -5275
rect -1846 -5279 -1806 -5277
rect -1806 -5281 -1798 -5279
rect -1846 -5284 -1798 -5281
rect -1846 -5297 -1806 -5286
rect -1671 -5288 -1663 -5280
rect -1663 -5296 -1655 -5288
rect -1854 -5302 -1680 -5298
rect -1671 -5314 -1663 -5308
rect -1642 -5314 -1637 -5268
rect -1619 -5314 -1614 -5268
rect -1530 -5314 -1526 -5268
rect -1506 -5314 -1502 -5268
rect -1482 -5314 -1478 -5268
rect -1458 -5314 -1454 -5268
rect -1434 -5314 -1430 -5268
rect -1410 -5314 -1406 -5268
rect -1386 -5314 -1382 -5268
rect -1362 -5314 -1358 -5268
rect -1338 -5293 -1334 -5268
rect -1314 -5269 -1310 -5268
rect -1338 -5314 -1331 -5293
rect -1314 -5314 -1307 -5269
rect -1290 -5314 -1286 -5268
rect -1266 -5314 -1262 -5268
rect -1242 -5314 -1238 -5268
rect -1218 -5314 -1214 -5268
rect -1194 -5314 -1190 -5268
rect -1170 -5314 -1166 -5268
rect -1146 -5314 -1142 -5268
rect -1122 -5314 -1118 -5268
rect -1098 -5314 -1094 -5268
rect -1074 -5314 -1070 -5268
rect -1050 -5314 -1046 -5268
rect -1026 -5314 -1022 -5268
rect -1002 -5314 -998 -5268
rect -978 -5314 -974 -5268
rect -954 -5314 -950 -5268
rect -930 -5314 -926 -5268
rect -906 -5314 -902 -5268
rect -893 -5275 -888 -5268
rect -882 -5275 -878 -5268
rect -883 -5289 -878 -5275
rect -893 -5299 -888 -5289
rect -883 -5313 -878 -5299
rect -882 -5314 -878 -5313
rect -858 -5314 -854 -5244
rect -834 -5314 -830 -5244
rect -810 -5314 -806 -5244
rect -786 -5314 -782 -5244
rect -762 -5314 -758 -5244
rect -738 -5314 -734 -5244
rect -714 -5314 -710 -5244
rect -690 -5314 -686 -5244
rect -666 -5314 -662 -5244
rect -642 -5313 -638 -5244
rect -653 -5314 -619 -5313
rect -2393 -5316 -1341 -5314
rect -2371 -5338 -2366 -5316
rect -2348 -5338 -2343 -5316
rect -2325 -5324 -2317 -5316
rect -2325 -5338 -2320 -5324
rect -2309 -5336 -2301 -5324
rect -2092 -5333 -2062 -5328
rect -2000 -5336 -1992 -5316
rect -2317 -5338 -2309 -5336
rect -2000 -5338 -1983 -5336
rect -1906 -5338 -1904 -5316
rect -1806 -5324 -1680 -5318
rect -1671 -5324 -1663 -5316
rect -1854 -5333 -1806 -5328
rect -1846 -5338 -1806 -5335
rect -1655 -5336 -1647 -5324
rect -1663 -5338 -1655 -5336
rect -1642 -5338 -1637 -5316
rect -1619 -5338 -1614 -5316
rect -1530 -5338 -1526 -5316
rect -1506 -5338 -1502 -5316
rect -1482 -5338 -1478 -5316
rect -1458 -5317 -1454 -5316
rect -2393 -5340 -1461 -5338
rect -2371 -5362 -2366 -5340
rect -2348 -5362 -2343 -5340
rect -2325 -5352 -2317 -5340
rect -2071 -5344 -2062 -5340
rect -2013 -5342 -1983 -5340
rect -2000 -5343 -1983 -5342
rect -2325 -5362 -2320 -5352
rect -2309 -5362 -2301 -5352
rect -2100 -5353 -2092 -5346
rect -2064 -5348 -2062 -5345
rect -2061 -5353 -2059 -5348
rect -2071 -5358 -2062 -5353
rect -2071 -5360 -2026 -5358
rect -2066 -5362 -2012 -5360
rect -2000 -5362 -1992 -5343
rect -1906 -5345 -1904 -5340
rect -1846 -5344 -1806 -5340
rect -1846 -5351 -1798 -5346
rect -1806 -5353 -1798 -5351
rect -1671 -5352 -1663 -5340
rect -1854 -5355 -1846 -5353
rect -1854 -5360 -1806 -5355
rect -1864 -5362 -1796 -5361
rect -1655 -5362 -1647 -5352
rect -1642 -5362 -1637 -5340
rect -1619 -5362 -1614 -5340
rect -1530 -5362 -1526 -5340
rect -1506 -5362 -1502 -5340
rect -1482 -5362 -1478 -5340
rect -1475 -5341 -1461 -5340
rect -1458 -5341 -1451 -5317
rect -1458 -5362 -1454 -5341
rect -1434 -5362 -1430 -5316
rect -1410 -5362 -1406 -5316
rect -1386 -5362 -1382 -5316
rect -1362 -5362 -1358 -5316
rect -1355 -5317 -1341 -5316
rect -1338 -5316 -619 -5314
rect -1338 -5317 -1317 -5316
rect -1314 -5317 -1307 -5316
rect -1338 -5338 -1331 -5317
rect -1314 -5338 -1310 -5317
rect -1290 -5338 -1286 -5316
rect -1266 -5338 -1262 -5316
rect -1242 -5338 -1238 -5316
rect -1218 -5338 -1214 -5316
rect -1194 -5338 -1190 -5316
rect -1170 -5338 -1166 -5316
rect -1146 -5338 -1142 -5316
rect -1122 -5338 -1118 -5316
rect -1098 -5338 -1094 -5316
rect -1074 -5338 -1070 -5316
rect -1050 -5338 -1046 -5316
rect -1026 -5338 -1022 -5316
rect -1002 -5338 -998 -5316
rect -978 -5338 -974 -5316
rect -954 -5338 -950 -5316
rect -930 -5338 -926 -5316
rect -906 -5338 -902 -5316
rect -882 -5338 -878 -5316
rect -858 -5338 -854 -5316
rect -834 -5338 -830 -5316
rect -810 -5337 -806 -5316
rect -821 -5338 -787 -5337
rect -1355 -5340 -787 -5338
rect -1355 -5341 -1341 -5340
rect -1338 -5341 -1331 -5340
rect -1338 -5362 -1334 -5341
rect -1314 -5362 -1310 -5340
rect -1290 -5362 -1286 -5340
rect -1266 -5362 -1262 -5340
rect -1242 -5362 -1238 -5340
rect -1218 -5362 -1214 -5340
rect -1194 -5362 -1190 -5340
rect -1170 -5362 -1166 -5340
rect -1146 -5362 -1142 -5340
rect -1122 -5362 -1118 -5340
rect -1098 -5362 -1094 -5340
rect -1074 -5362 -1070 -5340
rect -1050 -5362 -1046 -5340
rect -1026 -5362 -1022 -5340
rect -1002 -5362 -998 -5340
rect -978 -5361 -974 -5340
rect -989 -5362 -955 -5361
rect -2393 -5364 -955 -5362
rect -2371 -5410 -2366 -5364
rect -2348 -5410 -2343 -5364
rect -2325 -5368 -2320 -5364
rect -2317 -5368 -2309 -5364
rect -2325 -5380 -2317 -5368
rect -2066 -5369 -2062 -5364
rect -2147 -5372 -2134 -5370
rect -2292 -5378 -2071 -5372
rect -2325 -5410 -2320 -5380
rect -2092 -5394 -2062 -5392
rect -2094 -5398 -2062 -5394
rect -2000 -5410 -1992 -5364
rect -1846 -5371 -1806 -5364
rect -1663 -5368 -1655 -5364
rect -1846 -5378 -1680 -5372
rect -1671 -5380 -1663 -5368
rect -1854 -5394 -1806 -5392
rect -1854 -5398 -1680 -5394
rect -1926 -5410 -1892 -5407
rect -1642 -5410 -1637 -5364
rect -1619 -5410 -1614 -5364
rect -1530 -5410 -1526 -5364
rect -1506 -5410 -1502 -5364
rect -1482 -5410 -1478 -5364
rect -1458 -5410 -1454 -5364
rect -1434 -5410 -1430 -5364
rect -1410 -5410 -1406 -5364
rect -1386 -5410 -1382 -5364
rect -1362 -5410 -1358 -5364
rect -1338 -5410 -1334 -5364
rect -1314 -5410 -1310 -5364
rect -1290 -5410 -1286 -5364
rect -1266 -5410 -1262 -5364
rect -1242 -5410 -1238 -5364
rect -1218 -5410 -1214 -5364
rect -1194 -5410 -1190 -5364
rect -1170 -5410 -1166 -5364
rect -1146 -5410 -1142 -5364
rect -1122 -5410 -1118 -5364
rect -1098 -5410 -1094 -5364
rect -1074 -5410 -1070 -5364
rect -1050 -5410 -1046 -5364
rect -1026 -5410 -1022 -5364
rect -1002 -5410 -998 -5364
rect -989 -5371 -984 -5364
rect -978 -5371 -974 -5364
rect -979 -5385 -974 -5371
rect -989 -5395 -984 -5385
rect -979 -5409 -974 -5395
rect -978 -5410 -974 -5409
rect -954 -5410 -950 -5340
rect -930 -5410 -926 -5340
rect -906 -5410 -902 -5340
rect -882 -5410 -878 -5340
rect -858 -5341 -854 -5340
rect -858 -5386 -851 -5341
rect -834 -5386 -830 -5340
rect -821 -5347 -816 -5340
rect -810 -5347 -806 -5340
rect -811 -5361 -806 -5347
rect -821 -5371 -816 -5361
rect -811 -5385 -806 -5371
rect -810 -5386 -806 -5385
rect -786 -5386 -782 -5316
rect -762 -5386 -758 -5316
rect -738 -5386 -734 -5316
rect -714 -5386 -710 -5316
rect -690 -5386 -686 -5316
rect -666 -5386 -662 -5316
rect -653 -5323 -648 -5316
rect -642 -5323 -638 -5316
rect -643 -5337 -638 -5323
rect -653 -5338 -619 -5337
rect -618 -5338 -614 -5244
rect -594 -5338 -590 -5244
rect -570 -5338 -566 -5244
rect -546 -5338 -542 -5244
rect -522 -5338 -518 -5244
rect -498 -5338 -494 -5244
rect -474 -5338 -470 -5244
rect -450 -5338 -446 -5244
rect -426 -5338 -422 -5244
rect -402 -5290 -395 -5269
rect -378 -5290 -374 -5244
rect -354 -5290 -350 -5244
rect -330 -5290 -326 -5244
rect -306 -5290 -302 -5244
rect -282 -5290 -278 -5244
rect -258 -5290 -254 -5244
rect -234 -5290 -230 -5244
rect -186 -5245 -182 -5244
rect -221 -5268 -189 -5265
rect -221 -5275 -216 -5268
rect -203 -5269 -189 -5268
rect -186 -5269 -179 -5245
rect -173 -5275 -168 -5265
rect -162 -5275 -158 -5244
rect -149 -5251 -144 -5244
rect -138 -5251 -134 -5244
rect -139 -5265 -134 -5251
rect -211 -5289 -206 -5275
rect -163 -5289 -158 -5275
rect -210 -5290 -206 -5289
rect -197 -5290 -163 -5289
rect -419 -5292 -163 -5290
rect -419 -5293 -405 -5292
rect -402 -5293 -395 -5292
rect -402 -5338 -398 -5293
rect -378 -5338 -374 -5292
rect -354 -5338 -350 -5292
rect -330 -5338 -326 -5292
rect -306 -5338 -302 -5292
rect -282 -5338 -278 -5292
rect -258 -5338 -254 -5292
rect -234 -5338 -230 -5292
rect -210 -5337 -206 -5292
rect -221 -5338 -187 -5337
rect -653 -5340 -187 -5338
rect -653 -5347 -648 -5340
rect -643 -5361 -638 -5347
rect -642 -5386 -638 -5361
rect -618 -5386 -614 -5340
rect -594 -5386 -590 -5340
rect -570 -5386 -566 -5340
rect -546 -5386 -542 -5340
rect -522 -5386 -518 -5340
rect -498 -5386 -494 -5340
rect -474 -5386 -470 -5340
rect -450 -5386 -446 -5340
rect -426 -5386 -422 -5340
rect -402 -5386 -398 -5340
rect -378 -5386 -374 -5340
rect -354 -5386 -350 -5340
rect -330 -5386 -326 -5340
rect -306 -5386 -302 -5340
rect -282 -5386 -278 -5340
rect -258 -5385 -254 -5340
rect -245 -5371 -240 -5361
rect -234 -5371 -230 -5340
rect -221 -5347 -216 -5340
rect -210 -5347 -206 -5340
rect -211 -5361 -206 -5347
rect -197 -5351 -189 -5347
rect -203 -5361 -197 -5351
rect -235 -5385 -230 -5371
rect -269 -5386 -235 -5385
rect -875 -5388 -235 -5386
rect -875 -5389 -861 -5388
rect -858 -5389 -851 -5388
rect -858 -5410 -854 -5389
rect -834 -5410 -830 -5388
rect -810 -5410 -806 -5388
rect -786 -5410 -782 -5388
rect -762 -5410 -758 -5388
rect -738 -5410 -734 -5388
rect -714 -5410 -710 -5388
rect -690 -5410 -686 -5388
rect -666 -5410 -662 -5388
rect -642 -5410 -638 -5388
rect -618 -5389 -614 -5388
rect -2393 -5412 -621 -5410
rect -2371 -5434 -2366 -5412
rect -2348 -5434 -2343 -5412
rect -2325 -5434 -2320 -5412
rect -2054 -5413 -1906 -5412
rect -2054 -5414 -2036 -5413
rect -2309 -5428 -2301 -5418
rect -2317 -5434 -2309 -5428
rect -2068 -5429 -2038 -5422
rect -2000 -5430 -1992 -5413
rect -1920 -5414 -1906 -5413
rect -1846 -5420 -1794 -5412
rect -1852 -5427 -1804 -5422
rect -1902 -5429 -1804 -5427
rect -1655 -5428 -1647 -5418
rect -2000 -5432 -1975 -5430
rect -1902 -5431 -1852 -5429
rect -2025 -5434 -1975 -5432
rect -1846 -5434 -1804 -5431
rect -1663 -5434 -1655 -5428
rect -1642 -5434 -1637 -5412
rect -1619 -5434 -1614 -5412
rect -1530 -5434 -1526 -5412
rect -1506 -5434 -1502 -5412
rect -1482 -5434 -1478 -5412
rect -1458 -5434 -1454 -5412
rect -1434 -5434 -1430 -5412
rect -1410 -5434 -1406 -5412
rect -1386 -5434 -1382 -5412
rect -1362 -5434 -1358 -5412
rect -1338 -5434 -1334 -5412
rect -1314 -5434 -1310 -5412
rect -1290 -5434 -1286 -5412
rect -1266 -5434 -1262 -5412
rect -1242 -5434 -1238 -5412
rect -1218 -5434 -1214 -5412
rect -1194 -5434 -1190 -5412
rect -1170 -5434 -1166 -5412
rect -1146 -5433 -1142 -5412
rect -1157 -5434 -1123 -5433
rect -2393 -5436 -1123 -5434
rect -2371 -5458 -2366 -5436
rect -2348 -5458 -2343 -5436
rect -2325 -5458 -2320 -5436
rect -2054 -5437 -2038 -5436
rect -2000 -5437 -1966 -5436
rect -1846 -5437 -1804 -5436
rect -2000 -5438 -1975 -5437
rect -2076 -5446 -2054 -5439
rect -2309 -5456 -2301 -5446
rect -2044 -5449 -2038 -5444
rect -2028 -5446 -2001 -5439
rect -2054 -5456 -2038 -5449
rect -2015 -5447 -2001 -5446
rect -2015 -5456 -2014 -5447
rect -2317 -5458 -2309 -5456
rect -2044 -5458 -2028 -5456
rect -2000 -5458 -1992 -5438
rect -1982 -5439 -1975 -5438
rect -1862 -5439 -1798 -5438
rect -1985 -5446 -1796 -5439
rect -1862 -5447 -1798 -5446
rect -1852 -5456 -1804 -5449
rect -1655 -5456 -1647 -5446
rect -1976 -5458 -1940 -5457
rect -1663 -5458 -1655 -5456
rect -1642 -5458 -1637 -5436
rect -1619 -5458 -1614 -5436
rect -1530 -5458 -1526 -5436
rect -1506 -5458 -1502 -5436
rect -1482 -5458 -1478 -5436
rect -1458 -5458 -1454 -5436
rect -1434 -5458 -1430 -5436
rect -1410 -5458 -1406 -5436
rect -1386 -5458 -1382 -5436
rect -1362 -5458 -1358 -5436
rect -1338 -5458 -1334 -5436
rect -1314 -5458 -1310 -5436
rect -1290 -5458 -1286 -5436
rect -1266 -5458 -1262 -5436
rect -1242 -5458 -1238 -5436
rect -1218 -5458 -1214 -5436
rect -1194 -5458 -1190 -5436
rect -1170 -5458 -1166 -5436
rect -1157 -5443 -1152 -5436
rect -1146 -5443 -1142 -5436
rect -1147 -5457 -1142 -5443
rect -1122 -5458 -1118 -5412
rect -1098 -5458 -1094 -5412
rect -1074 -5458 -1070 -5412
rect -1050 -5458 -1046 -5412
rect -1026 -5458 -1022 -5412
rect -1002 -5458 -998 -5412
rect -978 -5458 -974 -5412
rect -954 -5437 -950 -5412
rect -2393 -5460 -957 -5458
rect -2371 -5530 -2366 -5460
rect -2348 -5530 -2343 -5460
rect -2325 -5494 -2320 -5460
rect -2317 -5462 -2309 -5460
rect -2076 -5473 -2054 -5466
rect -2325 -5502 -2317 -5494
rect -2060 -5500 -2030 -5497
rect -2325 -5522 -2320 -5502
rect -2317 -5510 -2309 -5502
rect -2060 -5513 -2038 -5502
rect -2033 -5509 -2030 -5500
rect -2028 -5504 -2027 -5500
rect -2068 -5518 -2038 -5515
rect -2325 -5530 -2317 -5522
rect -2000 -5530 -1992 -5460
rect -1846 -5464 -1804 -5460
rect -1663 -5462 -1655 -5460
rect -1846 -5474 -1794 -5465
rect -1912 -5485 -1884 -5483
rect -1852 -5491 -1804 -5487
rect -1844 -5500 -1796 -5497
rect -1671 -5502 -1663 -5494
rect -1844 -5513 -1804 -5502
rect -1663 -5510 -1655 -5502
rect -1852 -5518 -1680 -5514
rect -1926 -5530 -1892 -5527
rect -1671 -5530 -1663 -5522
rect -1642 -5530 -1637 -5460
rect -1619 -5530 -1614 -5460
rect -1530 -5530 -1526 -5460
rect -1506 -5530 -1502 -5460
rect -1482 -5530 -1478 -5460
rect -1458 -5530 -1454 -5460
rect -1434 -5530 -1430 -5460
rect -1410 -5530 -1406 -5460
rect -1386 -5530 -1382 -5460
rect -1362 -5530 -1358 -5460
rect -1338 -5530 -1334 -5460
rect -1314 -5530 -1310 -5460
rect -1290 -5530 -1286 -5460
rect -1266 -5530 -1262 -5460
rect -1242 -5530 -1238 -5460
rect -1218 -5530 -1214 -5460
rect -1194 -5530 -1190 -5460
rect -1170 -5530 -1166 -5460
rect -1157 -5506 -1123 -5505
rect -1122 -5506 -1118 -5460
rect -1098 -5506 -1094 -5460
rect -1074 -5506 -1070 -5460
rect -1050 -5506 -1046 -5460
rect -1037 -5491 -1032 -5481
rect -1026 -5491 -1022 -5460
rect -1027 -5505 -1022 -5491
rect -1002 -5506 -998 -5460
rect -978 -5506 -974 -5460
rect -971 -5461 -957 -5460
rect -954 -5485 -947 -5437
rect -954 -5506 -950 -5485
rect -930 -5506 -926 -5412
rect -906 -5506 -902 -5412
rect -882 -5506 -878 -5412
rect -858 -5506 -854 -5412
rect -845 -5467 -840 -5457
rect -834 -5467 -830 -5412
rect -835 -5481 -830 -5467
rect -845 -5482 -811 -5481
rect -810 -5482 -806 -5412
rect -786 -5413 -782 -5412
rect -786 -5461 -779 -5413
rect -786 -5482 -782 -5461
rect -762 -5482 -758 -5412
rect -738 -5482 -734 -5412
rect -714 -5482 -710 -5412
rect -690 -5482 -686 -5412
rect -666 -5482 -662 -5412
rect -642 -5482 -638 -5412
rect -635 -5413 -621 -5412
rect -618 -5437 -611 -5389
rect -618 -5482 -614 -5437
rect -594 -5482 -590 -5388
rect -570 -5482 -566 -5388
rect -546 -5482 -542 -5388
rect -522 -5482 -518 -5388
rect -498 -5482 -494 -5388
rect -474 -5482 -470 -5388
rect -450 -5482 -446 -5388
rect -426 -5482 -422 -5388
rect -402 -5482 -398 -5388
rect -378 -5482 -374 -5388
rect -354 -5482 -350 -5388
rect -330 -5482 -326 -5388
rect -306 -5482 -302 -5388
rect -282 -5482 -278 -5388
rect -269 -5395 -264 -5388
rect -258 -5395 -254 -5388
rect -259 -5409 -254 -5395
rect -269 -5419 -264 -5409
rect -259 -5433 -254 -5419
rect -258 -5481 -254 -5433
rect -269 -5482 -237 -5481
rect -845 -5484 -237 -5482
rect -845 -5491 -840 -5484
rect -835 -5505 -830 -5491
rect -834 -5506 -830 -5505
rect -810 -5506 -806 -5484
rect -786 -5506 -782 -5484
rect -762 -5506 -758 -5484
rect -738 -5506 -734 -5484
rect -714 -5506 -710 -5484
rect -690 -5506 -686 -5484
rect -666 -5506 -662 -5484
rect -642 -5506 -638 -5484
rect -618 -5506 -614 -5484
rect -594 -5506 -590 -5484
rect -570 -5506 -566 -5484
rect -546 -5506 -542 -5484
rect -522 -5506 -518 -5484
rect -498 -5506 -494 -5484
rect -474 -5506 -470 -5484
rect -450 -5506 -446 -5484
rect -426 -5506 -422 -5484
rect -402 -5506 -398 -5484
rect -378 -5506 -374 -5484
rect -354 -5506 -350 -5484
rect -330 -5506 -326 -5484
rect -306 -5506 -302 -5484
rect -282 -5505 -278 -5484
rect -269 -5491 -264 -5484
rect -258 -5491 -254 -5484
rect -251 -5485 -237 -5484
rect -259 -5505 -254 -5491
rect -245 -5495 -237 -5491
rect -251 -5505 -245 -5495
rect -293 -5506 -259 -5505
rect -1157 -5508 -259 -5506
rect -1157 -5515 -1152 -5508
rect -1122 -5509 -1118 -5508
rect -1147 -5529 -1142 -5515
rect -1133 -5519 -1125 -5515
rect -1139 -5529 -1133 -5519
rect -1146 -5530 -1142 -5529
rect -2393 -5532 -1125 -5530
rect -2371 -5554 -2366 -5532
rect -2348 -5554 -2343 -5532
rect -2325 -5538 -2317 -5532
rect -2325 -5554 -2320 -5538
rect -2309 -5550 -2301 -5538
rect -2068 -5549 -2038 -5542
rect -2317 -5554 -2309 -5550
rect -2000 -5552 -1992 -5532
rect -1844 -5540 -1794 -5532
rect -1671 -5538 -1663 -5532
rect -1852 -5549 -1804 -5542
rect -1655 -5550 -1647 -5538
rect -2025 -5553 -1991 -5552
rect -2025 -5554 -1975 -5553
rect -1844 -5554 -1804 -5551
rect -1663 -5554 -1655 -5550
rect -1642 -5554 -1637 -5532
rect -1619 -5554 -1614 -5532
rect -1530 -5554 -1526 -5532
rect -1506 -5554 -1502 -5532
rect -1482 -5554 -1478 -5532
rect -1458 -5554 -1454 -5532
rect -1434 -5554 -1430 -5532
rect -1410 -5554 -1406 -5532
rect -1386 -5554 -1382 -5532
rect -1362 -5554 -1358 -5532
rect -1338 -5554 -1334 -5532
rect -1314 -5554 -1310 -5532
rect -1290 -5554 -1286 -5532
rect -1266 -5553 -1262 -5532
rect -1277 -5554 -1243 -5553
rect -2393 -5556 -1243 -5554
rect -2371 -5578 -2366 -5556
rect -2348 -5578 -2343 -5556
rect -2325 -5566 -2317 -5556
rect -2060 -5566 -2020 -5559
rect -2004 -5564 -2001 -5559
rect -2015 -5566 -2001 -5564
rect -2000 -5566 -1992 -5556
rect -1972 -5558 -1958 -5556
rect -1844 -5557 -1804 -5556
rect -1862 -5559 -1796 -5558
rect -1985 -5561 -1796 -5559
rect -1985 -5566 -1852 -5561
rect -2325 -5578 -2320 -5566
rect -2309 -5578 -2301 -5566
rect -2068 -5576 -2060 -5569
rect -2015 -5576 -1990 -5566
rect -1844 -5567 -1796 -5561
rect -1671 -5566 -1663 -5556
rect -1852 -5576 -1804 -5569
rect -2020 -5578 -2004 -5576
rect -2000 -5578 -1992 -5576
rect -1976 -5578 -1940 -5577
rect -1655 -5578 -1647 -5566
rect -1642 -5578 -1637 -5556
rect -1619 -5578 -1614 -5556
rect -1530 -5578 -1526 -5556
rect -1506 -5578 -1502 -5556
rect -1482 -5578 -1478 -5556
rect -1458 -5578 -1454 -5556
rect -1434 -5578 -1430 -5556
rect -1410 -5578 -1406 -5556
rect -1386 -5578 -1382 -5556
rect -1362 -5578 -1358 -5556
rect -1338 -5578 -1334 -5556
rect -1314 -5578 -1310 -5556
rect -1290 -5578 -1286 -5556
rect -1277 -5563 -1272 -5556
rect -1266 -5563 -1262 -5556
rect -1267 -5577 -1262 -5563
rect -1242 -5578 -1238 -5532
rect -1218 -5578 -1214 -5532
rect -1194 -5578 -1190 -5532
rect -1170 -5578 -1166 -5532
rect -1146 -5578 -1142 -5532
rect -1139 -5533 -1125 -5532
rect -1122 -5533 -1115 -5509
rect -1098 -5578 -1094 -5508
rect -1074 -5578 -1070 -5508
rect -1050 -5578 -1046 -5508
rect -1037 -5539 -1032 -5529
rect -1027 -5553 -1022 -5539
rect -1026 -5578 -1022 -5553
rect -1002 -5557 -998 -5508
rect -2393 -5580 -1005 -5578
rect -2371 -5650 -2366 -5580
rect -2348 -5650 -2343 -5580
rect -2325 -5582 -2320 -5580
rect -2317 -5582 -2309 -5580
rect -2325 -5594 -2317 -5582
rect -2060 -5593 -2030 -5586
rect -2325 -5614 -2320 -5594
rect -2325 -5622 -2317 -5614
rect -2060 -5620 -2030 -5617
rect -2325 -5642 -2320 -5622
rect -2317 -5630 -2309 -5622
rect -2060 -5633 -2038 -5622
rect -2033 -5629 -2030 -5620
rect -2028 -5624 -2027 -5620
rect -2068 -5638 -2038 -5635
rect -2325 -5650 -2317 -5642
rect -2000 -5650 -1992 -5580
rect -1844 -5584 -1804 -5580
rect -1663 -5582 -1655 -5580
rect -1844 -5594 -1794 -5585
rect -1671 -5594 -1663 -5582
rect -1912 -5605 -1884 -5603
rect -1852 -5611 -1804 -5607
rect -1844 -5620 -1796 -5617
rect -1671 -5622 -1663 -5614
rect -1844 -5633 -1804 -5622
rect -1663 -5630 -1655 -5622
rect -1852 -5638 -1680 -5634
rect -1926 -5650 -1892 -5647
rect -1671 -5650 -1663 -5642
rect -1642 -5650 -1637 -5580
rect -1619 -5650 -1614 -5580
rect -1530 -5650 -1526 -5580
rect -1506 -5650 -1502 -5580
rect -1482 -5650 -1478 -5580
rect -1458 -5650 -1454 -5580
rect -1434 -5650 -1430 -5580
rect -1410 -5650 -1406 -5580
rect -1386 -5650 -1382 -5580
rect -1362 -5650 -1358 -5580
rect -1338 -5650 -1334 -5580
rect -1314 -5650 -1310 -5580
rect -1290 -5650 -1286 -5580
rect -1277 -5626 -1243 -5625
rect -1242 -5626 -1238 -5580
rect -1218 -5626 -1214 -5580
rect -1194 -5626 -1190 -5580
rect -1170 -5626 -1166 -5580
rect -1146 -5626 -1142 -5580
rect -1122 -5602 -1115 -5581
rect -1098 -5602 -1094 -5580
rect -1074 -5602 -1070 -5580
rect -1050 -5602 -1046 -5580
rect -1026 -5602 -1022 -5580
rect -1019 -5581 -1005 -5580
rect -1002 -5581 -995 -5557
rect -978 -5602 -974 -5508
rect -954 -5602 -950 -5508
rect -930 -5602 -926 -5508
rect -906 -5602 -902 -5508
rect -882 -5602 -878 -5508
rect -858 -5602 -854 -5508
rect -834 -5602 -830 -5508
rect -810 -5533 -806 -5508
rect -810 -5578 -803 -5533
rect -786 -5578 -782 -5508
rect -762 -5578 -758 -5508
rect -738 -5578 -734 -5508
rect -714 -5578 -710 -5508
rect -690 -5578 -686 -5508
rect -666 -5578 -662 -5508
rect -642 -5578 -638 -5508
rect -618 -5577 -614 -5508
rect -629 -5578 -595 -5577
rect -827 -5580 -595 -5578
rect -827 -5581 -813 -5580
rect -810 -5581 -803 -5580
rect -810 -5602 -806 -5581
rect -786 -5602 -782 -5580
rect -762 -5602 -758 -5580
rect -738 -5602 -734 -5580
rect -714 -5602 -710 -5580
rect -690 -5602 -686 -5580
rect -666 -5602 -662 -5580
rect -642 -5602 -638 -5580
rect -629 -5587 -624 -5580
rect -618 -5587 -614 -5580
rect -619 -5601 -614 -5587
rect -594 -5602 -590 -5508
rect -570 -5602 -566 -5508
rect -546 -5602 -542 -5508
rect -522 -5602 -518 -5508
rect -498 -5602 -494 -5508
rect -474 -5602 -470 -5508
rect -450 -5602 -446 -5508
rect -426 -5602 -422 -5508
rect -402 -5602 -398 -5508
rect -378 -5602 -374 -5508
rect -354 -5602 -350 -5508
rect -330 -5602 -326 -5508
rect -306 -5601 -302 -5508
rect -293 -5515 -288 -5508
rect -282 -5515 -278 -5508
rect -283 -5529 -278 -5515
rect -317 -5602 -283 -5601
rect -1139 -5604 -283 -5602
rect -1139 -5605 -1125 -5604
rect -1122 -5605 -1115 -5604
rect -1122 -5626 -1118 -5605
rect -1098 -5626 -1094 -5604
rect -1074 -5626 -1070 -5604
rect -1050 -5626 -1046 -5604
rect -1026 -5626 -1022 -5604
rect -1277 -5628 -1005 -5626
rect -1277 -5635 -1272 -5628
rect -1242 -5629 -1238 -5628
rect -1267 -5649 -1262 -5635
rect -1253 -5639 -1245 -5635
rect -1259 -5649 -1253 -5639
rect -1266 -5650 -1262 -5649
rect -2393 -5652 -1245 -5650
rect -2371 -5674 -2366 -5652
rect -2348 -5674 -2343 -5652
rect -2325 -5658 -2317 -5652
rect -2325 -5674 -2320 -5658
rect -2309 -5670 -2301 -5658
rect -2068 -5669 -2038 -5662
rect -2317 -5674 -2309 -5670
rect -2000 -5672 -1992 -5652
rect -1844 -5660 -1794 -5652
rect -1671 -5658 -1663 -5652
rect -1852 -5669 -1804 -5662
rect -1655 -5670 -1647 -5658
rect -2025 -5673 -1991 -5672
rect -2025 -5674 -1975 -5673
rect -1844 -5674 -1804 -5671
rect -1663 -5674 -1655 -5670
rect -1642 -5674 -1637 -5652
rect -1619 -5674 -1614 -5652
rect -1530 -5674 -1526 -5652
rect -1506 -5674 -1502 -5652
rect -1482 -5674 -1478 -5652
rect -1458 -5674 -1454 -5652
rect -1434 -5674 -1430 -5652
rect -1410 -5674 -1406 -5652
rect -1386 -5674 -1382 -5652
rect -1362 -5674 -1358 -5652
rect -1338 -5674 -1334 -5652
rect -1314 -5674 -1310 -5652
rect -1290 -5674 -1286 -5652
rect -1266 -5674 -1262 -5652
rect -1259 -5653 -1245 -5652
rect -1242 -5653 -1235 -5629
rect -1218 -5674 -1214 -5628
rect -1194 -5674 -1190 -5628
rect -1170 -5674 -1166 -5628
rect -1146 -5674 -1142 -5628
rect -1122 -5674 -1118 -5628
rect -1098 -5674 -1094 -5628
rect -1074 -5674 -1070 -5628
rect -1050 -5674 -1046 -5628
rect -1026 -5674 -1022 -5628
rect -1019 -5629 -1005 -5628
rect -1002 -5629 -995 -5605
rect -1002 -5674 -998 -5629
rect -978 -5674 -974 -5604
rect -954 -5674 -950 -5604
rect -930 -5674 -926 -5604
rect -906 -5674 -902 -5604
rect -882 -5674 -878 -5604
rect -858 -5674 -854 -5604
rect -834 -5674 -830 -5604
rect -810 -5674 -806 -5604
rect -786 -5674 -782 -5604
rect -762 -5674 -758 -5604
rect -738 -5674 -734 -5604
rect -714 -5674 -710 -5604
rect -690 -5674 -686 -5604
rect -666 -5674 -662 -5604
rect -642 -5674 -638 -5604
rect -629 -5659 -624 -5649
rect -594 -5653 -590 -5604
rect -619 -5673 -614 -5659
rect -605 -5663 -597 -5659
rect -611 -5673 -605 -5663
rect -618 -5674 -614 -5673
rect -605 -5674 -597 -5673
rect -2393 -5676 -597 -5674
rect -2371 -5698 -2366 -5676
rect -2348 -5698 -2343 -5676
rect -2325 -5686 -2317 -5676
rect -2060 -5686 -2020 -5679
rect -2004 -5684 -2001 -5679
rect -2015 -5686 -2001 -5684
rect -2000 -5686 -1992 -5676
rect -1972 -5678 -1958 -5676
rect -1844 -5677 -1804 -5676
rect -1862 -5679 -1796 -5678
rect -1985 -5681 -1796 -5679
rect -1985 -5686 -1852 -5681
rect -2325 -5698 -2320 -5686
rect -2309 -5698 -2301 -5686
rect -2068 -5696 -2060 -5689
rect -2015 -5696 -1990 -5686
rect -1844 -5687 -1796 -5681
rect -1671 -5686 -1663 -5676
rect -1852 -5696 -1804 -5689
rect -2020 -5698 -2004 -5696
rect -2000 -5698 -1992 -5696
rect -1976 -5698 -1940 -5697
rect -1655 -5698 -1647 -5686
rect -1642 -5698 -1637 -5676
rect -1619 -5698 -1614 -5676
rect -1530 -5698 -1526 -5676
rect -1506 -5698 -1502 -5676
rect -1482 -5698 -1478 -5676
rect -1458 -5698 -1454 -5676
rect -1434 -5698 -1430 -5676
rect -1410 -5697 -1406 -5676
rect -1421 -5698 -1387 -5697
rect -2393 -5700 -1387 -5698
rect -2371 -5770 -2366 -5700
rect -2348 -5770 -2343 -5700
rect -2325 -5702 -2320 -5700
rect -2317 -5702 -2309 -5700
rect -2325 -5714 -2317 -5702
rect -2060 -5713 -2030 -5706
rect -2325 -5734 -2320 -5714
rect -2325 -5742 -2317 -5734
rect -2060 -5740 -2030 -5737
rect -2325 -5762 -2320 -5742
rect -2317 -5750 -2309 -5742
rect -2060 -5753 -2038 -5742
rect -2033 -5749 -2030 -5740
rect -2028 -5744 -2027 -5740
rect -2068 -5758 -2038 -5755
rect -2325 -5770 -2317 -5762
rect -2000 -5767 -1992 -5700
rect -1844 -5704 -1804 -5700
rect -1663 -5702 -1655 -5700
rect -1844 -5714 -1794 -5705
rect -1671 -5714 -1663 -5702
rect -1912 -5725 -1884 -5723
rect -1852 -5731 -1804 -5727
rect -1844 -5740 -1796 -5737
rect -1671 -5742 -1663 -5734
rect -1844 -5753 -1804 -5742
rect -1663 -5750 -1655 -5742
rect -1852 -5758 -1680 -5754
rect -2119 -5770 -2069 -5768
rect -2007 -5770 -1977 -5767
rect -1926 -5770 -1892 -5767
rect -1671 -5770 -1663 -5762
rect -1642 -5770 -1637 -5700
rect -1619 -5770 -1614 -5700
rect -1530 -5770 -1526 -5700
rect -1506 -5770 -1502 -5700
rect -1482 -5770 -1478 -5700
rect -1458 -5770 -1454 -5700
rect -1434 -5770 -1430 -5700
rect -1421 -5707 -1416 -5700
rect -1410 -5707 -1406 -5700
rect -1411 -5721 -1406 -5707
rect -1421 -5746 -1387 -5745
rect -1386 -5746 -1382 -5676
rect -1362 -5746 -1358 -5676
rect -1338 -5746 -1334 -5676
rect -1314 -5746 -1310 -5676
rect -1290 -5746 -1286 -5676
rect -1266 -5746 -1262 -5676
rect -1242 -5722 -1235 -5701
rect -1218 -5722 -1214 -5676
rect -1194 -5722 -1190 -5676
rect -1170 -5721 -1166 -5676
rect -1181 -5722 -1147 -5721
rect -1259 -5724 -1147 -5722
rect -1259 -5725 -1245 -5724
rect -1242 -5725 -1235 -5724
rect -1242 -5746 -1238 -5725
rect -1218 -5746 -1214 -5724
rect -1194 -5746 -1190 -5724
rect -1181 -5731 -1176 -5724
rect -1170 -5731 -1166 -5724
rect -1171 -5745 -1166 -5731
rect -1146 -5746 -1142 -5676
rect -1122 -5746 -1118 -5676
rect -1098 -5746 -1094 -5676
rect -1074 -5746 -1070 -5676
rect -1050 -5746 -1046 -5676
rect -1026 -5746 -1022 -5676
rect -1002 -5746 -998 -5676
rect -978 -5746 -974 -5676
rect -954 -5746 -950 -5676
rect -930 -5746 -926 -5676
rect -906 -5746 -902 -5676
rect -882 -5746 -878 -5676
rect -858 -5746 -854 -5676
rect -834 -5746 -830 -5676
rect -810 -5746 -806 -5676
rect -786 -5746 -782 -5676
rect -762 -5746 -758 -5676
rect -738 -5746 -734 -5676
rect -714 -5746 -710 -5676
rect -690 -5746 -686 -5676
rect -666 -5746 -662 -5676
rect -642 -5746 -638 -5676
rect -618 -5746 -614 -5676
rect -611 -5677 -597 -5676
rect -594 -5677 -587 -5653
rect -605 -5698 -571 -5697
rect -570 -5698 -566 -5604
rect -546 -5698 -542 -5604
rect -522 -5698 -518 -5604
rect -498 -5698 -494 -5604
rect -474 -5698 -470 -5604
rect -450 -5698 -446 -5604
rect -426 -5698 -422 -5604
rect -402 -5698 -398 -5604
rect -378 -5698 -374 -5604
rect -354 -5697 -350 -5604
rect -341 -5635 -336 -5625
rect -330 -5635 -326 -5604
rect -317 -5611 -312 -5604
rect -306 -5611 -302 -5604
rect -307 -5625 -302 -5611
rect -331 -5649 -326 -5635
rect -365 -5698 -331 -5697
rect -605 -5700 -331 -5698
rect -1421 -5748 -597 -5746
rect -1421 -5755 -1416 -5748
rect -1411 -5769 -1406 -5755
rect -1410 -5770 -1406 -5769
rect -1386 -5770 -1382 -5748
rect -1362 -5770 -1358 -5748
rect -1338 -5770 -1334 -5748
rect -1314 -5770 -1310 -5748
rect -1290 -5770 -1286 -5748
rect -1266 -5770 -1262 -5748
rect -1242 -5770 -1238 -5748
rect -1218 -5770 -1214 -5748
rect -1194 -5770 -1190 -5748
rect -1146 -5770 -1142 -5748
rect -1122 -5770 -1118 -5748
rect -1098 -5770 -1094 -5748
rect -1074 -5770 -1070 -5748
rect -1050 -5770 -1046 -5748
rect -1026 -5770 -1022 -5748
rect -1002 -5770 -998 -5748
rect -978 -5770 -974 -5748
rect -954 -5770 -950 -5748
rect -930 -5770 -926 -5748
rect -906 -5770 -902 -5748
rect -882 -5770 -878 -5748
rect -858 -5770 -854 -5748
rect -834 -5770 -830 -5748
rect -810 -5770 -806 -5748
rect -786 -5770 -782 -5748
rect -762 -5770 -758 -5748
rect -738 -5770 -734 -5748
rect -714 -5770 -710 -5748
rect -690 -5770 -686 -5748
rect -666 -5770 -662 -5748
rect -642 -5770 -638 -5748
rect -618 -5770 -614 -5748
rect -611 -5749 -597 -5748
rect -594 -5749 -587 -5725
rect -570 -5749 -566 -5700
rect -594 -5769 -590 -5749
rect -605 -5770 -573 -5769
rect -2393 -5772 -573 -5770
rect -2371 -5794 -2366 -5772
rect -2348 -5794 -2343 -5772
rect -2325 -5776 -2317 -5772
rect -2325 -5792 -2320 -5776
rect -2317 -5778 -2309 -5776
rect -2309 -5790 -2301 -5778
rect -2000 -5786 -1992 -5772
rect -1671 -5776 -1663 -5772
rect -1663 -5778 -1655 -5776
rect -1844 -5780 -1806 -5778
rect -1854 -5786 -1806 -5782
rect -2068 -5789 -2060 -5786
rect -2030 -5789 -1958 -5786
rect -1942 -5789 -1806 -5786
rect -2317 -5792 -2309 -5790
rect -2000 -5792 -1992 -5789
rect -1655 -5790 -1647 -5778
rect -2325 -5794 -2317 -5792
rect -2033 -5794 -1992 -5792
rect -1844 -5793 -1806 -5791
rect -1663 -5792 -1655 -5790
rect -1864 -5794 -1796 -5793
rect -1671 -5794 -1663 -5792
rect -1642 -5794 -1637 -5772
rect -1619 -5794 -1614 -5772
rect -1530 -5794 -1526 -5772
rect -1506 -5794 -1502 -5772
rect -1482 -5794 -1478 -5772
rect -1458 -5794 -1454 -5772
rect -1434 -5794 -1430 -5772
rect -1410 -5794 -1406 -5772
rect -1386 -5773 -1382 -5772
rect -2393 -5796 -1389 -5794
rect -2371 -5818 -2366 -5796
rect -2348 -5818 -2343 -5796
rect -2325 -5804 -2317 -5796
rect -2060 -5799 -2030 -5796
rect -2000 -5799 -1992 -5796
rect -1972 -5798 -1958 -5796
rect -1904 -5799 -1798 -5796
rect -2078 -5803 -2020 -5799
rect -2023 -5804 -2020 -5803
rect -2000 -5801 -1798 -5799
rect -2000 -5803 -1854 -5801
rect -1844 -5803 -1798 -5801
rect -2325 -5818 -2320 -5804
rect -2317 -5806 -2309 -5804
rect -2020 -5806 -2004 -5804
rect -2000 -5806 -1992 -5803
rect -1671 -5804 -1663 -5796
rect -2309 -5818 -2301 -5806
rect -2020 -5808 -1992 -5806
rect -1844 -5807 -1806 -5805
rect -1663 -5806 -1655 -5804
rect -2023 -5813 -1992 -5808
rect -1854 -5813 -1806 -5809
rect -2068 -5816 -2060 -5813
rect -2030 -5816 -1806 -5813
rect -2074 -5818 -2060 -5816
rect -2020 -5818 -2004 -5816
rect -2000 -5818 -1992 -5816
rect -1655 -5818 -1647 -5806
rect -1642 -5818 -1637 -5796
rect -1619 -5818 -1614 -5796
rect -1530 -5818 -1526 -5796
rect -1506 -5818 -1502 -5796
rect -1482 -5818 -1478 -5796
rect -1458 -5817 -1454 -5796
rect -1469 -5818 -1435 -5817
rect -2393 -5820 -2060 -5818
rect -2050 -5820 -1435 -5818
rect -2371 -5866 -2366 -5820
rect -2348 -5866 -2343 -5820
rect -2325 -5832 -2317 -5820
rect -2109 -5823 -2108 -5820
rect -2117 -5830 -2108 -5823
rect -2325 -5852 -2320 -5832
rect -2317 -5834 -2309 -5832
rect -2109 -5834 -2108 -5830
rect -2060 -5830 -2030 -5823
rect -2060 -5834 -2034 -5830
rect -2325 -5860 -2317 -5852
rect -2101 -5857 -2071 -5854
rect -2325 -5866 -2320 -5860
rect -2317 -5866 -2309 -5860
rect -2000 -5862 -1992 -5820
rect -1844 -5821 -1806 -5820
rect -1844 -5830 -1798 -5823
rect -1671 -5832 -1663 -5820
rect -1844 -5834 -1806 -5832
rect -1663 -5834 -1655 -5832
rect -1854 -5848 -1680 -5844
rect -1846 -5857 -1798 -5854
rect -2079 -5863 -2043 -5862
rect -2007 -5863 -1991 -5862
rect -2079 -5864 -2071 -5863
rect -2079 -5866 -2029 -5864
rect -2011 -5866 -1991 -5863
rect -1846 -5865 -1806 -5859
rect -1671 -5860 -1663 -5852
rect -1864 -5866 -1796 -5865
rect -1663 -5866 -1655 -5860
rect -1642 -5866 -1637 -5820
rect -1619 -5866 -1614 -5820
rect -1530 -5866 -1526 -5820
rect -1506 -5866 -1502 -5820
rect -1482 -5866 -1478 -5820
rect -1469 -5827 -1464 -5820
rect -1458 -5827 -1454 -5820
rect -1459 -5841 -1454 -5827
rect -1434 -5866 -1430 -5796
rect -1410 -5866 -1406 -5796
rect -1403 -5797 -1389 -5796
rect -1386 -5797 -1379 -5773
rect -1386 -5842 -1379 -5821
rect -1362 -5842 -1358 -5772
rect -1338 -5842 -1334 -5772
rect -1314 -5842 -1310 -5772
rect -1290 -5842 -1286 -5772
rect -1266 -5842 -1262 -5772
rect -1242 -5842 -1238 -5772
rect -1218 -5842 -1214 -5772
rect -1194 -5842 -1190 -5772
rect -1181 -5803 -1176 -5793
rect -1146 -5797 -1142 -5772
rect -1171 -5817 -1166 -5803
rect -1157 -5807 -1149 -5803
rect -1163 -5817 -1157 -5807
rect -1170 -5842 -1166 -5817
rect -1146 -5821 -1139 -5797
rect -1122 -5842 -1118 -5772
rect -1098 -5842 -1094 -5772
rect -1074 -5842 -1070 -5772
rect -1050 -5841 -1046 -5772
rect -1061 -5842 -1027 -5841
rect -1403 -5844 -1027 -5842
rect -1403 -5845 -1389 -5844
rect -1386 -5845 -1379 -5844
rect -1386 -5866 -1382 -5845
rect -1362 -5866 -1358 -5844
rect -1338 -5866 -1334 -5844
rect -1314 -5866 -1310 -5844
rect -1290 -5866 -1286 -5844
rect -1266 -5866 -1262 -5844
rect -1242 -5866 -1238 -5844
rect -1218 -5866 -1214 -5844
rect -1194 -5866 -1190 -5844
rect -1170 -5866 -1166 -5844
rect -1122 -5866 -1118 -5844
rect -1098 -5866 -1094 -5844
rect -1074 -5866 -1070 -5844
rect -1061 -5851 -1056 -5844
rect -1050 -5851 -1046 -5844
rect -1051 -5865 -1046 -5851
rect -1026 -5866 -1022 -5772
rect -1002 -5865 -998 -5772
rect -1013 -5866 -979 -5865
rect -2393 -5868 -979 -5866
rect -2371 -5914 -2366 -5868
rect -2348 -5914 -2343 -5868
rect -2325 -5880 -2320 -5868
rect -2079 -5870 -2071 -5868
rect -2072 -5872 -2071 -5870
rect -2109 -5877 -2101 -5872
rect -2101 -5879 -2079 -5877
rect -2069 -5879 -2068 -5872
rect -2325 -5888 -2317 -5880
rect -2079 -5884 -2071 -5879
rect -2325 -5908 -2320 -5888
rect -2317 -5896 -2309 -5888
rect -2074 -5893 -2071 -5884
rect -2069 -5888 -2068 -5884
rect -2109 -5902 -2079 -5899
rect -2325 -5914 -2317 -5908
rect -2080 -5914 -2071 -5913
rect -2000 -5914 -1992 -5868
rect -1846 -5870 -1806 -5868
rect -1854 -5875 -1806 -5871
rect -1854 -5877 -1846 -5875
rect -1846 -5879 -1806 -5877
rect -1806 -5881 -1798 -5879
rect -1846 -5884 -1798 -5881
rect -1846 -5897 -1806 -5886
rect -1671 -5888 -1663 -5880
rect -1663 -5896 -1655 -5888
rect -1854 -5902 -1680 -5898
rect -1926 -5914 -1892 -5911
rect -1671 -5914 -1663 -5908
rect -1642 -5914 -1637 -5868
rect -1619 -5914 -1614 -5868
rect -1530 -5914 -1526 -5868
rect -1506 -5914 -1502 -5868
rect -1482 -5914 -1478 -5868
rect -1469 -5890 -1435 -5889
rect -1434 -5890 -1430 -5868
rect -1410 -5890 -1406 -5868
rect -1386 -5890 -1382 -5868
rect -1362 -5890 -1358 -5868
rect -1338 -5890 -1334 -5868
rect -1314 -5890 -1310 -5868
rect -1290 -5890 -1286 -5868
rect -1266 -5890 -1262 -5868
rect -1242 -5890 -1238 -5868
rect -1218 -5890 -1214 -5868
rect -1194 -5890 -1190 -5868
rect -1170 -5890 -1166 -5868
rect -1146 -5890 -1139 -5869
rect -1122 -5890 -1118 -5868
rect -1098 -5890 -1094 -5868
rect -1074 -5890 -1070 -5868
rect -1026 -5890 -1022 -5868
rect -1013 -5875 -1008 -5868
rect -1002 -5875 -998 -5868
rect -1003 -5889 -998 -5875
rect -978 -5890 -974 -5772
rect -954 -5890 -950 -5772
rect -930 -5890 -926 -5772
rect -906 -5890 -902 -5772
rect -882 -5890 -878 -5772
rect -858 -5890 -854 -5772
rect -834 -5890 -830 -5772
rect -810 -5890 -806 -5772
rect -786 -5890 -782 -5772
rect -762 -5890 -758 -5772
rect -738 -5890 -734 -5772
rect -714 -5890 -710 -5772
rect -690 -5890 -686 -5772
rect -666 -5890 -662 -5772
rect -642 -5890 -638 -5772
rect -618 -5890 -614 -5772
rect -605 -5779 -600 -5772
rect -594 -5779 -590 -5772
rect -587 -5773 -573 -5772
rect -595 -5793 -590 -5779
rect -581 -5783 -573 -5779
rect -587 -5793 -581 -5783
rect -570 -5794 -563 -5749
rect -546 -5793 -542 -5700
rect -557 -5794 -523 -5793
rect -587 -5796 -523 -5794
rect -587 -5797 -573 -5796
rect -570 -5797 -563 -5796
rect -605 -5827 -600 -5817
rect -595 -5841 -590 -5827
rect -594 -5890 -590 -5841
rect -570 -5845 -566 -5797
rect -557 -5803 -552 -5796
rect -546 -5803 -542 -5796
rect -547 -5817 -542 -5803
rect -557 -5842 -523 -5841
rect -522 -5842 -518 -5700
rect -498 -5842 -494 -5700
rect -474 -5842 -470 -5700
rect -450 -5842 -446 -5700
rect -426 -5841 -422 -5700
rect -413 -5827 -408 -5817
rect -402 -5827 -398 -5700
rect -389 -5755 -384 -5745
rect -378 -5755 -374 -5700
rect -365 -5707 -360 -5700
rect -354 -5707 -350 -5700
rect -355 -5721 -350 -5707
rect -379 -5769 -374 -5755
rect -403 -5841 -398 -5827
rect -437 -5842 -403 -5841
rect -557 -5844 -403 -5842
rect -570 -5869 -563 -5845
rect -557 -5851 -552 -5844
rect -547 -5865 -542 -5851
rect -546 -5890 -542 -5865
rect -522 -5869 -518 -5844
rect -1469 -5892 -525 -5890
rect -1469 -5899 -1464 -5892
rect -1434 -5893 -1430 -5892
rect -1459 -5913 -1454 -5899
rect -1445 -5903 -1437 -5899
rect -1451 -5913 -1445 -5903
rect -1458 -5914 -1454 -5913
rect -2393 -5916 -1437 -5914
rect -2371 -5938 -2366 -5916
rect -2348 -5938 -2343 -5916
rect -2325 -5922 -2317 -5916
rect -2325 -5938 -2320 -5922
rect -2317 -5924 -2309 -5922
rect -2309 -5936 -2301 -5924
rect -2080 -5925 -2071 -5916
rect -2068 -5926 -2059 -5925
rect -2068 -5933 -2038 -5926
rect -2317 -5938 -2309 -5936
rect -2068 -5938 -2059 -5933
rect -2000 -5934 -1992 -5916
rect -1846 -5924 -1794 -5916
rect -1671 -5922 -1663 -5916
rect -1663 -5924 -1655 -5922
rect -1852 -5933 -1804 -5926
rect -2011 -5936 -1983 -5934
rect -2025 -5937 -1983 -5936
rect -2025 -5938 -1975 -5937
rect -1846 -5938 -1804 -5935
rect -1655 -5936 -1647 -5924
rect -1663 -5938 -1655 -5936
rect -1642 -5938 -1637 -5916
rect -1619 -5938 -1614 -5916
rect -1530 -5938 -1526 -5916
rect -1506 -5938 -1502 -5916
rect -1482 -5938 -1478 -5916
rect -1458 -5938 -1454 -5916
rect -1451 -5917 -1437 -5916
rect -1434 -5917 -1427 -5893
rect -1410 -5938 -1406 -5892
rect -1386 -5938 -1382 -5892
rect -1362 -5938 -1358 -5892
rect -1338 -5938 -1334 -5892
rect -1314 -5938 -1310 -5892
rect -1290 -5938 -1286 -5892
rect -1266 -5938 -1262 -5892
rect -1242 -5938 -1238 -5892
rect -1218 -5938 -1214 -5892
rect -1194 -5938 -1190 -5892
rect -1170 -5938 -1166 -5892
rect -1163 -5893 -1149 -5892
rect -1146 -5893 -1139 -5892
rect -1146 -5938 -1142 -5893
rect -1122 -5938 -1118 -5892
rect -1098 -5938 -1094 -5892
rect -1074 -5938 -1070 -5892
rect -1026 -5917 -1022 -5892
rect -1061 -5938 -1029 -5937
rect -2393 -5940 -1029 -5938
rect -2371 -5962 -2366 -5940
rect -2348 -5962 -2343 -5940
rect -2325 -5950 -2317 -5940
rect -2068 -5941 -2038 -5940
rect -2068 -5943 -2059 -5941
rect -2013 -5942 -1983 -5940
rect -1846 -5941 -1804 -5940
rect -2000 -5943 -1983 -5942
rect -1862 -5943 -1798 -5942
rect -2076 -5950 -2068 -5943
rect -2061 -5950 -2045 -5948
rect -2038 -5950 -2001 -5943
rect -2325 -5962 -2320 -5950
rect -2317 -5952 -2309 -5950
rect -2309 -5962 -2301 -5952
rect -2068 -5953 -2045 -5950
rect -2015 -5951 -2001 -5950
rect -2068 -5960 -2038 -5953
rect -2068 -5962 -2045 -5960
rect -2000 -5962 -1992 -5943
rect -1985 -5945 -1796 -5943
rect -1985 -5950 -1852 -5945
rect -1846 -5950 -1796 -5945
rect -1671 -5950 -1663 -5940
rect -1846 -5951 -1798 -5950
rect -1663 -5952 -1655 -5950
rect -1852 -5960 -1804 -5953
rect -1976 -5962 -1940 -5961
rect -1655 -5962 -1647 -5952
rect -1642 -5962 -1637 -5940
rect -1619 -5962 -1614 -5940
rect -1530 -5962 -1526 -5940
rect -1506 -5962 -1502 -5940
rect -1482 -5962 -1478 -5940
rect -1458 -5962 -1454 -5940
rect -1410 -5962 -1406 -5940
rect -1386 -5962 -1382 -5940
rect -1362 -5962 -1358 -5940
rect -1338 -5962 -1334 -5940
rect -1314 -5962 -1310 -5940
rect -1290 -5962 -1286 -5940
rect -1266 -5962 -1262 -5940
rect -1242 -5962 -1238 -5940
rect -1218 -5962 -1214 -5940
rect -1194 -5962 -1190 -5940
rect -1170 -5962 -1166 -5940
rect -1146 -5962 -1142 -5940
rect -1122 -5962 -1118 -5940
rect -1098 -5962 -1094 -5940
rect -1074 -5961 -1070 -5940
rect -1061 -5947 -1056 -5940
rect -1043 -5941 -1029 -5940
rect -1026 -5941 -1019 -5917
rect -978 -5941 -974 -5892
rect -1051 -5961 -1046 -5947
rect -1085 -5962 -1051 -5961
rect -2393 -5964 -1051 -5962
rect -2371 -6405 -2366 -5964
rect -2361 -6385 -2353 -6375
rect -2348 -6385 -2343 -5964
rect -2351 -6401 -2343 -6385
rect -2371 -6431 -2363 -6405
rect -2383 -6603 -2376 -6593
rect -2371 -6603 -2366 -6431
rect -2373 -6614 -2366 -6603
rect -2348 -6614 -2343 -6401
rect -2325 -5966 -2320 -5964
rect -2317 -5966 -2309 -5964
rect -2325 -5978 -2317 -5966
rect -2068 -5970 -2059 -5964
rect -2076 -5977 -2071 -5970
rect -2068 -5978 -2059 -5977
rect -2325 -5998 -2320 -5978
rect -2317 -5980 -2309 -5978
rect -2325 -6006 -2317 -5998
rect -2060 -6004 -2030 -6001
rect -2325 -6026 -2320 -6006
rect -2317 -6014 -2309 -6006
rect -2060 -6017 -2038 -6006
rect -2033 -6013 -2030 -6004
rect -2028 -6008 -2027 -6004
rect -2068 -6022 -2038 -6019
rect -2325 -6042 -2317 -6026
rect -2325 -6119 -2320 -6042
rect -2309 -6054 -2301 -6043
rect -2317 -6059 -2309 -6054
rect -2309 -6082 -2301 -6072
rect -2251 -6078 -2093 -6072
rect -2317 -6088 -2309 -6082
rect -2124 -6085 -2108 -6082
rect -2060 -6085 -2030 -6080
rect -2000 -6081 -1992 -5964
rect -1846 -5968 -1804 -5964
rect -1663 -5966 -1655 -5964
rect -1846 -5978 -1794 -5969
rect -1671 -5978 -1663 -5966
rect -1663 -5980 -1655 -5978
rect -1912 -5989 -1884 -5987
rect -1852 -5995 -1804 -5991
rect -1844 -6004 -1796 -6001
rect -1671 -6006 -1663 -5998
rect -1844 -6017 -1804 -6006
rect -1663 -6014 -1655 -6006
rect -1852 -6022 -1680 -6018
rect -1844 -6044 -1837 -6042
rect -1789 -6044 -1680 -6042
rect -1837 -6053 -1789 -6052
rect -1655 -6054 -1647 -6046
rect -1837 -6068 -1796 -6055
rect -1663 -6062 -1655 -6054
rect -1796 -6078 -1789 -6073
rect -1837 -6080 -1796 -6078
rect -2000 -6084 -1990 -6081
rect -1844 -6082 -1837 -6080
rect -1655 -6082 -1647 -6074
rect -2124 -6098 -2113 -6092
rect -2325 -6129 -2317 -6119
rect -2325 -6148 -2320 -6129
rect -2317 -6135 -2309 -6129
rect -2243 -6146 -2221 -6138
rect -2211 -6146 -2201 -6126
rect -2073 -6146 -2065 -6128
rect -2000 -6146 -1992 -6084
rect -1844 -6085 -1796 -6082
rect -1837 -6098 -1796 -6088
rect -1663 -6090 -1655 -6082
rect -1671 -6130 -1663 -6122
rect -1655 -6130 -1647 -6128
rect -1663 -6138 -1647 -6130
rect -1642 -6138 -1637 -5964
rect -1885 -6146 -1877 -6144
rect -1708 -6146 -1672 -6144
rect -2243 -6147 -2213 -6146
rect -2325 -6157 -2317 -6148
rect -2259 -6153 -2211 -6147
rect -2183 -6153 -1877 -6146
rect -1869 -6153 -1758 -6146
rect -1710 -6152 -1672 -6146
rect -1710 -6153 -1692 -6152
rect -2211 -6157 -2201 -6153
rect -2325 -6177 -2320 -6157
rect -2317 -6164 -2309 -6157
rect -2211 -6164 -2198 -6157
rect -2325 -6185 -2317 -6177
rect -2300 -6184 -2292 -6174
rect -2243 -6183 -2228 -6172
rect -2211 -6180 -2181 -6164
rect -2211 -6183 -2201 -6180
rect -2325 -6205 -2320 -6185
rect -2317 -6193 -2309 -6185
rect -2325 -6213 -2317 -6205
rect -2325 -6233 -2320 -6213
rect -2317 -6221 -2309 -6213
rect -2325 -6242 -2317 -6233
rect -2325 -6261 -2320 -6242
rect -2317 -6249 -2309 -6242
rect -2325 -6270 -2317 -6261
rect -2325 -6290 -2320 -6270
rect -2317 -6277 -2309 -6270
rect -2325 -6298 -2317 -6290
rect -2290 -6297 -2282 -6184
rect -2251 -6194 -2240 -6190
rect -2211 -6194 -2181 -6190
rect -2251 -6197 -2181 -6194
rect -2176 -6204 -2173 -6202
rect -2240 -6211 -2173 -6204
rect -2169 -6209 -2163 -6154
rect -2073 -6190 -2065 -6153
rect -2073 -6194 -2043 -6190
rect -2000 -6194 -1992 -6153
rect -1915 -6184 -1907 -6175
rect -1963 -6190 -1955 -6184
rect -1963 -6194 -1915 -6190
rect -1885 -6194 -1877 -6153
rect -1875 -6158 -1869 -6154
rect -1829 -6176 -1781 -6174
rect -1847 -6180 -1781 -6176
rect -1778 -6180 -1771 -6154
rect -1758 -6161 -1710 -6154
rect -1718 -6168 -1710 -6161
rect -1768 -6178 -1760 -6168
rect -1718 -6170 -1700 -6168
rect -2146 -6197 -2135 -6194
rect -2105 -6197 -2043 -6194
rect -2035 -6197 -1989 -6194
rect -1973 -6197 -1915 -6194
rect -1907 -6197 -1854 -6194
rect -2073 -6199 -2043 -6197
rect -2135 -6211 -2105 -6204
rect -2065 -6206 -2043 -6199
rect -2243 -6222 -2240 -6213
rect -2221 -6219 -2213 -6211
rect -2211 -6219 -2208 -6211
rect -2203 -6218 -2173 -6211
rect -2251 -6229 -2240 -6222
rect -2211 -6222 -2203 -6219
rect -2211 -6229 -2181 -6222
rect -2073 -6229 -2043 -6222
rect -2203 -6252 -2173 -6245
rect -2262 -6270 -2240 -6260
rect -2203 -6261 -2176 -6252
rect -2083 -6263 -2075 -6253
rect -2040 -6263 -2035 -6259
rect -2073 -6275 -2043 -6263
rect -2028 -6275 -2023 -6263
rect -2000 -6270 -1992 -6197
rect -1963 -6200 -1955 -6197
rect -1963 -6201 -1915 -6200
rect -1955 -6211 -1907 -6204
rect -1885 -6208 -1877 -6197
rect -1837 -6202 -1828 -6186
rect -1758 -6193 -1750 -6178
rect -1758 -6194 -1692 -6193
rect -1837 -6204 -1833 -6202
rect -1837 -6206 -1835 -6204
rect -1887 -6211 -1851 -6208
rect -1750 -6211 -1702 -6204
rect -1885 -6216 -1877 -6211
rect -1963 -6229 -1915 -6222
rect -1905 -6261 -1897 -6216
rect -1857 -6234 -1851 -6211
rect -1760 -6219 -1758 -6218
rect -1837 -6229 -1789 -6222
rect -1758 -6228 -1750 -6222
rect -1758 -6229 -1710 -6228
rect -1955 -6264 -1915 -6261
rect -1963 -6270 -1962 -6268
rect -2000 -6273 -1981 -6270
rect -1965 -6273 -1962 -6270
rect -1955 -6270 -1907 -6266
rect -1885 -6270 -1877 -6251
rect -1857 -6264 -1851 -6252
rect -1750 -6256 -1702 -6249
rect -1829 -6264 -1789 -6262
rect -1766 -6266 -1760 -6256
rect -1829 -6270 -1781 -6266
rect -1756 -6270 -1740 -6266
rect -1680 -6270 -1672 -6152
rect -1671 -6158 -1663 -6150
rect -1645 -6154 -1637 -6138
rect -1663 -6166 -1655 -6158
rect -1671 -6186 -1663 -6178
rect -1663 -6194 -1655 -6186
rect -1671 -6214 -1663 -6206
rect -1671 -6230 -1669 -6217
rect -1663 -6222 -1655 -6214
rect -1671 -6242 -1663 -6234
rect -1663 -6250 -1655 -6242
rect -1671 -6270 -1663 -6262
rect -1955 -6273 -1837 -6270
rect -1829 -6273 -1740 -6270
rect -2206 -6283 -2176 -6280
rect -2206 -6286 -2203 -6283
rect -2161 -6285 -2145 -6276
rect -2073 -6278 -2065 -6275
rect -2073 -6279 -2043 -6278
rect -2028 -6279 -2012 -6275
rect -2073 -6286 -2065 -6280
rect -2203 -6287 -2176 -6286
rect -2065 -6287 -2043 -6286
rect -2262 -6293 -2232 -6287
rect -2176 -6293 -2173 -6287
rect -2043 -6293 -2035 -6287
rect -2325 -6318 -2320 -6298
rect -2317 -6306 -2309 -6298
rect -2153 -6299 -2146 -6295
rect -2325 -6326 -2317 -6318
rect -2300 -6322 -2292 -6312
rect -2325 -6346 -2320 -6326
rect -2317 -6334 -2309 -6326
rect -2325 -6354 -2317 -6346
rect -2325 -6374 -2320 -6354
rect -2317 -6362 -2309 -6354
rect -2290 -6355 -2282 -6322
rect -2273 -6326 -2264 -6321
rect -2206 -6326 -2176 -6321
rect -2262 -6333 -2232 -6328
rect -2198 -6337 -2176 -6326
rect -2198 -6351 -2176 -6343
rect -2166 -6359 -2158 -6311
rect -2143 -6315 -2136 -6299
rect -2143 -6326 -2113 -6321
rect -2073 -6326 -2065 -6321
rect -2065 -6328 -2043 -6326
rect -2043 -6333 -2035 -6328
rect -2065 -6354 -2043 -6339
rect -2006 -6355 -2004 -6339
rect -2265 -6369 -2260 -6363
rect -2143 -6369 -2113 -6362
rect -2270 -6370 -2240 -6369
rect -2270 -6373 -2265 -6370
rect -2325 -6382 -2317 -6374
rect -2325 -6402 -2320 -6382
rect -2317 -6390 -2309 -6382
rect -2113 -6385 -2105 -6375
rect -2291 -6397 -2270 -6390
rect -2198 -6392 -2168 -6390
rect -2135 -6391 -2105 -6390
rect -2103 -6391 -2095 -6385
rect -2113 -6392 -2105 -6391
rect -2065 -6392 -2035 -6390
rect -2000 -6392 -1992 -6273
rect -1963 -6280 -1960 -6273
rect -1915 -6277 -1905 -6273
rect -1963 -6281 -1955 -6280
rect -1963 -6287 -1915 -6281
rect -1989 -6314 -1973 -6311
rect -1915 -6314 -1907 -6307
rect -1990 -6349 -1989 -6328
rect -1983 -6392 -1981 -6329
rect -1885 -6338 -1877 -6273
rect -1789 -6278 -1778 -6273
rect -1837 -6281 -1829 -6280
rect -1837 -6287 -1789 -6281
rect -1756 -6282 -1740 -6273
rect -1837 -6297 -1829 -6287
rect -1872 -6316 -1867 -6306
rect -1789 -6314 -1781 -6307
rect -1776 -6314 -1769 -6297
rect -1756 -6304 -1750 -6282
rect -1671 -6286 -1669 -6275
rect -1663 -6278 -1655 -6270
rect -1671 -6298 -1663 -6290
rect -1663 -6306 -1655 -6298
rect -1702 -6316 -1696 -6310
rect -1955 -6340 -1915 -6338
rect -1963 -6342 -1955 -6340
rect -1963 -6349 -1915 -6342
rect -1963 -6357 -1955 -6349
rect -1963 -6358 -1915 -6357
rect -1973 -6364 -1965 -6361
rect -1955 -6364 -1907 -6360
rect -1974 -6367 -1907 -6364
rect -1973 -6371 -1965 -6367
rect -1963 -6371 -1960 -6369
rect -1963 -6375 -1915 -6371
rect -1963 -6383 -1955 -6375
rect -1963 -6387 -1915 -6383
rect -1963 -6390 -1955 -6387
rect -2240 -6397 -2206 -6392
rect -2198 -6397 -2143 -6392
rect -2113 -6397 -1981 -6392
rect -1915 -6397 -1907 -6390
rect -2270 -6402 -2266 -6398
rect -2086 -6401 -2070 -6397
rect -2325 -6410 -2317 -6402
rect -2270 -6409 -2240 -6402
rect -2206 -6409 -2176 -6402
rect -2325 -6430 -2320 -6410
rect -2317 -6418 -2309 -6410
rect -2270 -6414 -2266 -6409
rect -2270 -6418 -2266 -6415
rect -2198 -6418 -2176 -6411
rect -2166 -6418 -2158 -6401
rect -2143 -6409 -2113 -6402
rect -2198 -6427 -2168 -6423
rect -2325 -6438 -2317 -6430
rect -2143 -6432 -2136 -6418
rect -2085 -6423 -2060 -6422
rect -2039 -6423 -2035 -6414
rect -2135 -6430 -2105 -6423
rect -2085 -6430 -2035 -6423
rect -2029 -6430 -2025 -6423
rect -2325 -6451 -2320 -6438
rect -2317 -6446 -2309 -6438
rect -2235 -6448 -2232 -6445
rect -2325 -6477 -2317 -6451
rect -2325 -6486 -2320 -6477
rect -2325 -6494 -2317 -6486
rect -2135 -6494 -2119 -6481
rect -2000 -6489 -1992 -6397
rect -1983 -6415 -1981 -6397
rect -1955 -6415 -1915 -6414
rect -1862 -6418 -1857 -6316
rect -1706 -6320 -1702 -6316
rect -1829 -6332 -1789 -6324
rect -1671 -6326 -1663 -6318
rect -1849 -6340 -1842 -6332
rect -1790 -6340 -1781 -6332
rect -1663 -6334 -1655 -6326
rect -1837 -6349 -1829 -6342
rect -1758 -6349 -1732 -6342
rect -1748 -6358 -1732 -6349
rect -1671 -6354 -1663 -6346
rect -1829 -6367 -1781 -6360
rect -1663 -6362 -1655 -6354
rect -1829 -6373 -1789 -6369
rect -1768 -6372 -1760 -6362
rect -1758 -6373 -1750 -6372
rect -1671 -6382 -1663 -6374
rect -1837 -6385 -1780 -6382
rect -1758 -6388 -1748 -6382
rect -1708 -6388 -1690 -6382
rect -1829 -6397 -1781 -6390
rect -1680 -6399 -1672 -6382
rect -1663 -6390 -1655 -6382
rect -1829 -6408 -1791 -6402
rect -1758 -6408 -1710 -6406
rect -1758 -6415 -1692 -6408
rect -1671 -6410 -1663 -6402
rect -1955 -6426 -1907 -6423
rect -1791 -6426 -1781 -6423
rect -1991 -6430 -1839 -6426
rect -1791 -6430 -1780 -6426
rect -1680 -6433 -1672 -6415
rect -1663 -6418 -1655 -6410
rect -1839 -6443 -1791 -6436
rect -1671 -6438 -1663 -6430
rect -1829 -6449 -1791 -6445
rect -1671 -6448 -1669 -6438
rect -1663 -6446 -1655 -6438
rect -1680 -6464 -1672 -6449
rect -1642 -6464 -1637 -6154
rect -1619 -6204 -1614 -5964
rect -1619 -6230 -1611 -6204
rect -1768 -6480 -1760 -6470
rect -1758 -6487 -1710 -6480
rect -2325 -6514 -2320 -6494
rect -2317 -6502 -2306 -6494
rect -2031 -6497 -1992 -6489
rect -1750 -6491 -1710 -6487
rect -1674 -6492 -1663 -6486
rect -2307 -6510 -2306 -6502
rect -2149 -6499 -2135 -6498
rect -2149 -6503 -2119 -6499
rect -2024 -6508 -2021 -6499
rect -2325 -6522 -2317 -6514
rect -2325 -6570 -2320 -6522
rect -2317 -6530 -2306 -6522
rect -2185 -6524 -2169 -6512
rect -2056 -6515 -2040 -6511
rect -2021 -6515 -2008 -6508
rect -2056 -6526 -2054 -6516
rect -2056 -6527 -2048 -6526
rect -2307 -6566 -2306 -6558
rect -2111 -6559 -2054 -6553
rect -2325 -6578 -2314 -6570
rect -2104 -6577 -2101 -6573
rect -2325 -6598 -2320 -6578
rect -2314 -6586 -2306 -6578
rect -2104 -6580 -2101 -6578
rect -2084 -6580 -2054 -6579
rect -2000 -6580 -1992 -6497
rect -1758 -6498 -1750 -6497
rect -1758 -6499 -1749 -6498
rect -1758 -6500 -1710 -6499
rect -1663 -6502 -1658 -6492
rect -1831 -6510 -1783 -6506
rect -1784 -6523 -1783 -6510
rect -1674 -6520 -1663 -6514
rect -1826 -6525 -1796 -6524
rect -1663 -6530 -1658 -6520
rect -1654 -6524 -1647 -6514
rect -1644 -6538 -1637 -6524
rect -1758 -6556 -1750 -6553
rect -1758 -6559 -1710 -6556
rect -1844 -6571 -1828 -6569
rect -1844 -6572 -1792 -6571
rect -1828 -6573 -1792 -6572
rect -1772 -6573 -1758 -6565
rect -1750 -6568 -1702 -6561
rect -1750 -6576 -1710 -6572
rect -1700 -6576 -1692 -6556
rect -1674 -6564 -1665 -6556
rect -1674 -6576 -1666 -6568
rect -1758 -6580 -1710 -6579
rect -2307 -6594 -2306 -6586
rect -2139 -6590 -2123 -6581
rect -2111 -6586 -2016 -6580
rect -2139 -6597 -2111 -6590
rect -2325 -6606 -2314 -6598
rect -2177 -6604 -2161 -6603
rect -2141 -6604 -2119 -6602
rect -2104 -6604 -2101 -6586
rect -2076 -6597 -2046 -6592
rect -2325 -6614 -2320 -6606
rect -2314 -6614 -2306 -6606
rect -2076 -6608 -2054 -6602
rect -2021 -6605 -2016 -6586
rect -2000 -6586 -1818 -6580
rect -1802 -6586 -1776 -6580
rect -1760 -6586 -1710 -6580
rect -1666 -6584 -1658 -6576
rect -2189 -6614 -2175 -6609
rect -2373 -6616 -2175 -6614
rect -2373 -6617 -2359 -6616
rect -2371 -7029 -2366 -6617
rect -2348 -6669 -2343 -6616
rect -2325 -6626 -2320 -6616
rect -2307 -6622 -2306 -6616
rect -2189 -6617 -2175 -6616
rect -2149 -6618 -2119 -6609
rect -2084 -6610 -2036 -6609
rect -2000 -6610 -1992 -6586
rect -1758 -6588 -1710 -6586
rect -1758 -6590 -1755 -6588
rect -1828 -6597 -1792 -6590
rect -1768 -6599 -1760 -6592
rect -1758 -6597 -1757 -6590
rect -1710 -6591 -1702 -6590
rect -1750 -6597 -1702 -6591
rect -1674 -6592 -1665 -6584
rect -1768 -6602 -1764 -6599
rect -1758 -6602 -1755 -6597
rect -1818 -6610 -1789 -6602
rect -1758 -6609 -1754 -6602
rect -1750 -6607 -1710 -6602
rect -1674 -6604 -1666 -6596
rect -1758 -6610 -1692 -6609
rect -2084 -6612 -1692 -6610
rect -1666 -6612 -1658 -6604
rect -2084 -6615 -1690 -6612
rect -2084 -6618 -2054 -6615
rect -2046 -6617 -1710 -6615
rect -2325 -6634 -2314 -6626
rect -2076 -6627 -2046 -6620
rect -2325 -6654 -2320 -6634
rect -2314 -6642 -2306 -6634
rect -2076 -6635 -2054 -6629
rect -2084 -6639 -2054 -6637
rect -2104 -6642 -2054 -6639
rect -2307 -6650 -2306 -6642
rect -2084 -6645 -2054 -6642
rect -2325 -6666 -2314 -6654
rect -2348 -6693 -2341 -6669
rect -2325 -6683 -2320 -6666
rect -2314 -6670 -2309 -6666
rect -2309 -6682 -2298 -6670
rect -2314 -6683 -2309 -6682
rect -2361 -7009 -2353 -6999
rect -2348 -7009 -2343 -6693
rect -2351 -7025 -2343 -7009
rect -2371 -7055 -2363 -7029
rect -2383 -7227 -2376 -7217
rect -2371 -7227 -2366 -7055
rect -2373 -7238 -2366 -7227
rect -2348 -7238 -2343 -7025
rect -2325 -6695 -2314 -6683
rect -2076 -6694 -2073 -6678
rect -2325 -6712 -2320 -6695
rect -2314 -6698 -2309 -6695
rect -2309 -6710 -2298 -6698
rect -2251 -6702 -2101 -6695
rect -2141 -6709 -2111 -6703
rect -2086 -6705 -2083 -6695
rect -2076 -6709 -2046 -6703
rect -2314 -6712 -2309 -6710
rect -2325 -6724 -2314 -6712
rect -2141 -6721 -2113 -6716
rect -2076 -6721 -2073 -6718
rect -2325 -6743 -2320 -6724
rect -2314 -6726 -2309 -6724
rect -2325 -6753 -2317 -6743
rect -2325 -6772 -2320 -6753
rect -2317 -6759 -2309 -6753
rect -2243 -6770 -2221 -6762
rect -2211 -6770 -2201 -6750
rect -2073 -6770 -2065 -6752
rect -2000 -6770 -1992 -6617
rect -1758 -6618 -1710 -6617
rect -1680 -6620 -1665 -6612
rect -1750 -6627 -1702 -6620
rect -1680 -6624 -1672 -6620
rect -1680 -6629 -1666 -6624
rect -1836 -6633 -1820 -6632
rect -1837 -6637 -1820 -6633
rect -1750 -6635 -1710 -6629
rect -1674 -6632 -1666 -6629
rect -1837 -6644 -1789 -6637
rect -1758 -6638 -1710 -6637
rect -1760 -6641 -1692 -6638
rect -1666 -6640 -1658 -6632
rect -1837 -6645 -1820 -6644
rect -1764 -6645 -1692 -6641
rect -1674 -6645 -1665 -6640
rect -1680 -6648 -1665 -6645
rect -1680 -6676 -1672 -6648
rect -1666 -6668 -1665 -6658
rect -1837 -6678 -1789 -6676
rect -1829 -6692 -1789 -6678
rect -1655 -6680 -1650 -6670
rect -1666 -6686 -1655 -6680
rect -1778 -6694 -1771 -6692
rect -1710 -6694 -1702 -6692
rect -1666 -6696 -1665 -6686
rect -1837 -6702 -1829 -6696
rect -1829 -6703 -1789 -6702
rect -1726 -6703 -1710 -6702
rect -1789 -6705 -1781 -6703
rect -1829 -6709 -1781 -6705
rect -1750 -6709 -1710 -6703
rect -1829 -6721 -1789 -6712
rect -1726 -6718 -1710 -6709
rect -1706 -6718 -1702 -6705
rect -1655 -6708 -1650 -6698
rect -1666 -6714 -1655 -6708
rect -1666 -6724 -1665 -6714
rect -1671 -6754 -1663 -6746
rect -1655 -6754 -1647 -6752
rect -1663 -6762 -1647 -6754
rect -1642 -6762 -1637 -6538
rect -1619 -6540 -1614 -6230
rect -1885 -6770 -1877 -6768
rect -1708 -6770 -1672 -6768
rect -2243 -6771 -2213 -6770
rect -2325 -6781 -2317 -6772
rect -2259 -6777 -2211 -6771
rect -2183 -6777 -1877 -6770
rect -1869 -6777 -1758 -6770
rect -1710 -6776 -1672 -6770
rect -1710 -6777 -1692 -6776
rect -2211 -6781 -2201 -6777
rect -2325 -6801 -2320 -6781
rect -2317 -6788 -2309 -6781
rect -2211 -6788 -2198 -6781
rect -2325 -6809 -2317 -6801
rect -2300 -6808 -2292 -6798
rect -2243 -6807 -2228 -6796
rect -2211 -6804 -2181 -6788
rect -2211 -6807 -2201 -6804
rect -2325 -6829 -2320 -6809
rect -2317 -6817 -2309 -6809
rect -2325 -6837 -2317 -6829
rect -2325 -6857 -2320 -6837
rect -2317 -6845 -2309 -6837
rect -2325 -6866 -2317 -6857
rect -2325 -6885 -2320 -6866
rect -2317 -6873 -2309 -6866
rect -2325 -6894 -2317 -6885
rect -2325 -6914 -2320 -6894
rect -2317 -6901 -2309 -6894
rect -2325 -6922 -2317 -6914
rect -2290 -6921 -2282 -6808
rect -2251 -6818 -2240 -6814
rect -2211 -6818 -2181 -6814
rect -2251 -6821 -2181 -6818
rect -2176 -6828 -2173 -6826
rect -2240 -6835 -2173 -6828
rect -2169 -6833 -2163 -6778
rect -2073 -6814 -2065 -6777
rect -2073 -6818 -2043 -6814
rect -2000 -6818 -1992 -6777
rect -1915 -6808 -1907 -6799
rect -1963 -6814 -1955 -6808
rect -1963 -6818 -1915 -6814
rect -1885 -6818 -1877 -6777
rect -1875 -6782 -1869 -6778
rect -1829 -6800 -1781 -6798
rect -1847 -6804 -1781 -6800
rect -1778 -6804 -1771 -6778
rect -1758 -6785 -1710 -6778
rect -1718 -6792 -1710 -6785
rect -1768 -6802 -1760 -6792
rect -1718 -6794 -1700 -6792
rect -2146 -6821 -2135 -6818
rect -2105 -6821 -2043 -6818
rect -2035 -6821 -1989 -6818
rect -1973 -6821 -1915 -6818
rect -1907 -6821 -1854 -6818
rect -2073 -6823 -2043 -6821
rect -2135 -6835 -2105 -6828
rect -2065 -6830 -2043 -6823
rect -2243 -6846 -2240 -6837
rect -2221 -6843 -2213 -6835
rect -2211 -6843 -2208 -6835
rect -2203 -6842 -2173 -6835
rect -2251 -6853 -2240 -6846
rect -2211 -6846 -2203 -6843
rect -2211 -6853 -2181 -6846
rect -2073 -6853 -2043 -6846
rect -2203 -6876 -2173 -6869
rect -2262 -6894 -2240 -6884
rect -2203 -6885 -2176 -6876
rect -2083 -6887 -2075 -6877
rect -2040 -6887 -2035 -6883
rect -2073 -6899 -2043 -6887
rect -2028 -6899 -2023 -6887
rect -2000 -6894 -1992 -6821
rect -1963 -6824 -1955 -6821
rect -1963 -6825 -1915 -6824
rect -1955 -6835 -1907 -6828
rect -1885 -6832 -1877 -6821
rect -1837 -6826 -1828 -6810
rect -1758 -6817 -1750 -6802
rect -1758 -6818 -1692 -6817
rect -1837 -6828 -1833 -6826
rect -1837 -6830 -1835 -6828
rect -1887 -6835 -1851 -6832
rect -1750 -6835 -1702 -6828
rect -1885 -6840 -1877 -6835
rect -1963 -6853 -1915 -6846
rect -1905 -6885 -1897 -6840
rect -1857 -6858 -1851 -6835
rect -1760 -6843 -1758 -6842
rect -1837 -6853 -1789 -6846
rect -1758 -6852 -1750 -6846
rect -1758 -6853 -1710 -6852
rect -1955 -6888 -1915 -6885
rect -1963 -6894 -1962 -6892
rect -2000 -6897 -1981 -6894
rect -1965 -6897 -1962 -6894
rect -1955 -6894 -1907 -6890
rect -1885 -6894 -1877 -6875
rect -1857 -6888 -1851 -6876
rect -1750 -6880 -1702 -6873
rect -1829 -6888 -1789 -6886
rect -1766 -6890 -1760 -6880
rect -1829 -6894 -1781 -6890
rect -1756 -6894 -1740 -6890
rect -1680 -6894 -1672 -6776
rect -1671 -6782 -1663 -6774
rect -1645 -6778 -1637 -6762
rect -1663 -6790 -1655 -6782
rect -1671 -6810 -1663 -6802
rect -1663 -6818 -1655 -6810
rect -1671 -6838 -1663 -6830
rect -1671 -6854 -1669 -6841
rect -1663 -6846 -1655 -6838
rect -1671 -6866 -1663 -6858
rect -1663 -6874 -1655 -6866
rect -1671 -6894 -1663 -6886
rect -1955 -6897 -1837 -6894
rect -1829 -6897 -1740 -6894
rect -2206 -6907 -2176 -6904
rect -2206 -6910 -2203 -6907
rect -2161 -6909 -2145 -6900
rect -2073 -6902 -2065 -6899
rect -2073 -6903 -2043 -6902
rect -2028 -6903 -2012 -6899
rect -2073 -6910 -2065 -6904
rect -2203 -6911 -2176 -6910
rect -2065 -6911 -2043 -6910
rect -2262 -6917 -2232 -6911
rect -2176 -6917 -2173 -6911
rect -2043 -6917 -2035 -6911
rect -2325 -6942 -2320 -6922
rect -2317 -6930 -2309 -6922
rect -2153 -6923 -2146 -6919
rect -2325 -6950 -2317 -6942
rect -2300 -6946 -2292 -6936
rect -2325 -6970 -2320 -6950
rect -2317 -6958 -2309 -6950
rect -2325 -6978 -2317 -6970
rect -2325 -6998 -2320 -6978
rect -2317 -6986 -2309 -6978
rect -2290 -6979 -2282 -6946
rect -2273 -6950 -2264 -6945
rect -2206 -6950 -2176 -6945
rect -2262 -6957 -2232 -6952
rect -2198 -6961 -2176 -6950
rect -2198 -6975 -2176 -6967
rect -2166 -6983 -2158 -6935
rect -2143 -6939 -2136 -6923
rect -2143 -6950 -2113 -6945
rect -2073 -6950 -2065 -6945
rect -2065 -6952 -2043 -6950
rect -2043 -6957 -2035 -6952
rect -2065 -6978 -2043 -6963
rect -2006 -6979 -2004 -6963
rect -2265 -6993 -2260 -6987
rect -2143 -6993 -2113 -6986
rect -2270 -6994 -2240 -6993
rect -2270 -6997 -2265 -6994
rect -2325 -7006 -2317 -6998
rect -2325 -7026 -2320 -7006
rect -2317 -7014 -2309 -7006
rect -2113 -7009 -2105 -6999
rect -2291 -7021 -2270 -7014
rect -2198 -7016 -2168 -7014
rect -2135 -7015 -2105 -7014
rect -2103 -7015 -2095 -7009
rect -2113 -7016 -2105 -7015
rect -2065 -7016 -2035 -7014
rect -2000 -7016 -1992 -6897
rect -1963 -6904 -1960 -6897
rect -1915 -6901 -1905 -6897
rect -1963 -6905 -1955 -6904
rect -1963 -6911 -1915 -6905
rect -1989 -6938 -1973 -6935
rect -1915 -6938 -1907 -6931
rect -1990 -6973 -1989 -6952
rect -1983 -7016 -1981 -6953
rect -1885 -6962 -1877 -6897
rect -1789 -6902 -1778 -6897
rect -1837 -6905 -1829 -6904
rect -1837 -6911 -1789 -6905
rect -1756 -6906 -1740 -6897
rect -1837 -6921 -1829 -6911
rect -1872 -6940 -1867 -6930
rect -1789 -6938 -1781 -6931
rect -1776 -6938 -1769 -6921
rect -1756 -6928 -1750 -6906
rect -1671 -6910 -1669 -6899
rect -1663 -6902 -1655 -6894
rect -1671 -6922 -1663 -6914
rect -1663 -6930 -1655 -6922
rect -1702 -6940 -1696 -6934
rect -1955 -6964 -1915 -6962
rect -1963 -6966 -1955 -6964
rect -1963 -6973 -1915 -6966
rect -1963 -6981 -1955 -6973
rect -1963 -6982 -1915 -6981
rect -1973 -6988 -1965 -6985
rect -1955 -6988 -1907 -6984
rect -1974 -6991 -1907 -6988
rect -1973 -6995 -1965 -6991
rect -1963 -6995 -1960 -6993
rect -1963 -6999 -1915 -6995
rect -1963 -7007 -1955 -6999
rect -1963 -7011 -1915 -7007
rect -1963 -7014 -1955 -7011
rect -2240 -7021 -2206 -7016
rect -2198 -7021 -2143 -7016
rect -2113 -7021 -1981 -7016
rect -1915 -7021 -1907 -7014
rect -2270 -7026 -2266 -7022
rect -2086 -7025 -2070 -7021
rect -2325 -7034 -2317 -7026
rect -2270 -7033 -2240 -7026
rect -2206 -7033 -2176 -7026
rect -2325 -7054 -2320 -7034
rect -2317 -7042 -2309 -7034
rect -2270 -7038 -2266 -7033
rect -2270 -7042 -2266 -7039
rect -2198 -7042 -2176 -7035
rect -2166 -7042 -2158 -7025
rect -2143 -7033 -2113 -7026
rect -2198 -7051 -2168 -7047
rect -2325 -7062 -2317 -7054
rect -2143 -7056 -2136 -7042
rect -2085 -7047 -2060 -7046
rect -2039 -7047 -2035 -7038
rect -2135 -7054 -2105 -7047
rect -2085 -7054 -2035 -7047
rect -2029 -7054 -2025 -7047
rect -2325 -7075 -2320 -7062
rect -2317 -7070 -2309 -7062
rect -2235 -7072 -2232 -7069
rect -2325 -7101 -2317 -7075
rect -2325 -7110 -2320 -7101
rect -2325 -7118 -2317 -7110
rect -2135 -7118 -2119 -7105
rect -2000 -7113 -1992 -7021
rect -1983 -7039 -1981 -7021
rect -1955 -7039 -1915 -7038
rect -1862 -7042 -1857 -6940
rect -1706 -6944 -1702 -6940
rect -1829 -6956 -1789 -6948
rect -1671 -6950 -1663 -6942
rect -1849 -6964 -1842 -6956
rect -1790 -6964 -1781 -6956
rect -1663 -6958 -1655 -6950
rect -1837 -6973 -1829 -6966
rect -1758 -6973 -1732 -6966
rect -1748 -6982 -1732 -6973
rect -1671 -6978 -1663 -6970
rect -1829 -6991 -1781 -6984
rect -1663 -6986 -1655 -6978
rect -1829 -6997 -1789 -6993
rect -1768 -6996 -1760 -6986
rect -1758 -6997 -1750 -6996
rect -1671 -7006 -1663 -6998
rect -1837 -7009 -1780 -7006
rect -1758 -7012 -1748 -7006
rect -1708 -7012 -1690 -7006
rect -1829 -7021 -1781 -7014
rect -1680 -7023 -1672 -7006
rect -1663 -7014 -1655 -7006
rect -1829 -7032 -1791 -7026
rect -1758 -7032 -1710 -7030
rect -1758 -7039 -1692 -7032
rect -1671 -7034 -1663 -7026
rect -1955 -7050 -1907 -7047
rect -1791 -7050 -1781 -7047
rect -1991 -7054 -1839 -7050
rect -1791 -7054 -1780 -7050
rect -1680 -7057 -1672 -7039
rect -1663 -7042 -1655 -7034
rect -1839 -7067 -1791 -7060
rect -1671 -7062 -1663 -7054
rect -1829 -7073 -1791 -7069
rect -1671 -7072 -1669 -7062
rect -1663 -7070 -1655 -7062
rect -1680 -7088 -1672 -7073
rect -1642 -7088 -1637 -6778
rect -1619 -6614 -1612 -6590
rect -1619 -6828 -1614 -6614
rect -1619 -6854 -1611 -6828
rect -1768 -7104 -1760 -7094
rect -1758 -7111 -1710 -7104
rect -2325 -7138 -2320 -7118
rect -2317 -7126 -2306 -7118
rect -2031 -7121 -1992 -7113
rect -1750 -7115 -1710 -7111
rect -1674 -7116 -1663 -7110
rect -2307 -7134 -2306 -7126
rect -2149 -7123 -2135 -7122
rect -2149 -7127 -2119 -7123
rect -2024 -7132 -2021 -7123
rect -2325 -7146 -2317 -7138
rect -2325 -7194 -2320 -7146
rect -2317 -7154 -2306 -7146
rect -2185 -7148 -2169 -7136
rect -2056 -7139 -2040 -7135
rect -2021 -7139 -2008 -7132
rect -2056 -7150 -2054 -7140
rect -2056 -7151 -2048 -7150
rect -2307 -7190 -2306 -7182
rect -2111 -7183 -2054 -7177
rect -2325 -7202 -2314 -7194
rect -2104 -7201 -2101 -7197
rect -2325 -7222 -2320 -7202
rect -2314 -7210 -2306 -7202
rect -2104 -7204 -2101 -7202
rect -2084 -7204 -2054 -7203
rect -2000 -7204 -1992 -7121
rect -1758 -7122 -1750 -7121
rect -1758 -7123 -1749 -7122
rect -1758 -7124 -1710 -7123
rect -1663 -7126 -1658 -7116
rect -1831 -7134 -1783 -7130
rect -1784 -7147 -1783 -7134
rect -1674 -7144 -1663 -7138
rect -1826 -7149 -1796 -7148
rect -1663 -7154 -1658 -7144
rect -1654 -7148 -1647 -7138
rect -1644 -7162 -1637 -7148
rect -1758 -7180 -1750 -7177
rect -1758 -7183 -1710 -7180
rect -1844 -7195 -1828 -7193
rect -1844 -7196 -1792 -7195
rect -1828 -7197 -1792 -7196
rect -1772 -7197 -1758 -7189
rect -1750 -7192 -1702 -7185
rect -1750 -7200 -1710 -7196
rect -1700 -7200 -1692 -7180
rect -1674 -7188 -1665 -7180
rect -1674 -7200 -1666 -7192
rect -1758 -7204 -1710 -7203
rect -2307 -7218 -2306 -7210
rect -2139 -7214 -2123 -7205
rect -2111 -7210 -2016 -7204
rect -2139 -7221 -2111 -7214
rect -2325 -7230 -2314 -7222
rect -2177 -7228 -2161 -7227
rect -2141 -7228 -2119 -7226
rect -2104 -7228 -2101 -7210
rect -2076 -7221 -2046 -7216
rect -2325 -7238 -2320 -7230
rect -2314 -7238 -2306 -7230
rect -2076 -7232 -2054 -7226
rect -2021 -7229 -2016 -7210
rect -2000 -7210 -1818 -7204
rect -1802 -7210 -1776 -7204
rect -1760 -7210 -1710 -7204
rect -1666 -7208 -1658 -7200
rect -2189 -7238 -2175 -7233
rect -2373 -7240 -2175 -7238
rect -2373 -7241 -2359 -7240
rect -2371 -7402 -2366 -7241
rect -2348 -7293 -2343 -7240
rect -2325 -7250 -2320 -7240
rect -2307 -7246 -2306 -7240
rect -2189 -7241 -2175 -7240
rect -2149 -7242 -2119 -7233
rect -2084 -7234 -2036 -7233
rect -2000 -7234 -1992 -7210
rect -1758 -7212 -1710 -7210
rect -1758 -7214 -1755 -7212
rect -1828 -7221 -1792 -7214
rect -1768 -7223 -1760 -7216
rect -1758 -7221 -1757 -7214
rect -1710 -7215 -1702 -7214
rect -1750 -7221 -1702 -7215
rect -1674 -7216 -1665 -7208
rect -1768 -7226 -1764 -7223
rect -1758 -7226 -1755 -7221
rect -1818 -7234 -1789 -7226
rect -1758 -7233 -1754 -7226
rect -1750 -7231 -1710 -7226
rect -1674 -7228 -1666 -7220
rect -1758 -7234 -1692 -7233
rect -2084 -7236 -1692 -7234
rect -1666 -7236 -1658 -7228
rect -2084 -7239 -1690 -7236
rect -2084 -7242 -2054 -7239
rect -2046 -7241 -1710 -7239
rect -2325 -7258 -2314 -7250
rect -2076 -7251 -2046 -7244
rect -2325 -7278 -2320 -7258
rect -2314 -7266 -2306 -7258
rect -2076 -7259 -2054 -7253
rect -2084 -7263 -2054 -7261
rect -2104 -7266 -2054 -7263
rect -2307 -7274 -2306 -7266
rect -2084 -7269 -2054 -7266
rect -2325 -7290 -2314 -7278
rect -2078 -7283 -2026 -7282
rect -2348 -7317 -2341 -7293
rect -2325 -7306 -2320 -7290
rect -2314 -7294 -2309 -7290
rect -2309 -7306 -2298 -7294
rect -2068 -7295 -2038 -7293
rect -2068 -7297 -2013 -7295
rect -2038 -7302 -2013 -7297
rect -2348 -7402 -2343 -7317
rect -2325 -7318 -2314 -7306
rect -2068 -7309 -2046 -7302
rect -2011 -7311 -2003 -7302
rect -2076 -7318 -2046 -7311
rect -2038 -7312 -2001 -7311
rect -2000 -7312 -1992 -7241
rect -1758 -7242 -1710 -7241
rect -1680 -7244 -1665 -7236
rect -1750 -7251 -1702 -7244
rect -1680 -7248 -1672 -7244
rect -1680 -7253 -1666 -7248
rect -1836 -7257 -1820 -7256
rect -1837 -7261 -1820 -7257
rect -1750 -7259 -1710 -7253
rect -1674 -7256 -1666 -7253
rect -1837 -7268 -1789 -7261
rect -1758 -7262 -1710 -7261
rect -1760 -7265 -1692 -7262
rect -1666 -7264 -1658 -7256
rect -1837 -7269 -1820 -7268
rect -1764 -7269 -1692 -7265
rect -1674 -7269 -1665 -7264
rect -1680 -7272 -1665 -7269
rect -1852 -7297 -1804 -7293
rect -1829 -7309 -1804 -7302
rect -1804 -7311 -1781 -7310
rect -2038 -7314 -1992 -7312
rect -2038 -7318 -2001 -7314
rect -2325 -7334 -2320 -7318
rect -2314 -7322 -2309 -7318
rect -2015 -7319 -2001 -7318
rect -2309 -7334 -2298 -7322
rect -2046 -7327 -2038 -7320
rect -2325 -7346 -2314 -7334
rect -2076 -7345 -2046 -7338
rect -2325 -7366 -2320 -7346
rect -2314 -7350 -2309 -7346
rect -2325 -7374 -2317 -7366
rect -2060 -7372 -2030 -7369
rect -2325 -7402 -2320 -7374
rect -2317 -7382 -2309 -7374
rect -2060 -7385 -2038 -7374
rect -2033 -7381 -2030 -7372
rect -2028 -7376 -2027 -7372
rect -2068 -7390 -2038 -7387
rect -2000 -7402 -1992 -7314
rect -1985 -7318 -1852 -7311
rect -1829 -7318 -1781 -7311
rect -1750 -7315 -1682 -7310
rect -1680 -7315 -1672 -7272
rect -1671 -7290 -1666 -7276
rect -1666 -7292 -1655 -7290
rect -1655 -7304 -1650 -7292
rect -1666 -7306 -1655 -7304
rect -1750 -7318 -1702 -7315
rect -1671 -7318 -1666 -7306
rect -1666 -7320 -1655 -7318
rect -1852 -7327 -1804 -7320
rect -1829 -7336 -1804 -7329
rect -1655 -7332 -1650 -7320
rect -1666 -7334 -1655 -7332
rect -1829 -7345 -1794 -7337
rect -1671 -7346 -1666 -7334
rect -1666 -7348 -1655 -7346
rect -1912 -7357 -1884 -7355
rect -1852 -7363 -1804 -7359
rect -1844 -7372 -1796 -7369
rect -1671 -7374 -1663 -7366
rect -1844 -7385 -1804 -7374
rect -1663 -7382 -1655 -7374
rect -1852 -7390 -1680 -7386
rect -1642 -7402 -1637 -7162
rect -1619 -7164 -1614 -6854
rect -1619 -7238 -1612 -7214
rect -1619 -7402 -1614 -7238
rect -1530 -7402 -1526 -5964
rect -1517 -6187 -1512 -6177
rect -1506 -6187 -1502 -5964
rect -1493 -5995 -1488 -5985
rect -1482 -5995 -1478 -5964
rect -1483 -6009 -1478 -5995
rect -1493 -6010 -1459 -6009
rect -1458 -6010 -1454 -5964
rect -1434 -5989 -1427 -5965
rect -1434 -6010 -1430 -5989
rect -1410 -6010 -1406 -5964
rect -1386 -6010 -1382 -5964
rect -1362 -6010 -1358 -5964
rect -1338 -6010 -1334 -5964
rect -1314 -6010 -1310 -5964
rect -1290 -6010 -1286 -5964
rect -1266 -6010 -1262 -5964
rect -1242 -6010 -1238 -5964
rect -1218 -6010 -1214 -5964
rect -1194 -6010 -1190 -5964
rect -1170 -6010 -1166 -5964
rect -1146 -6010 -1142 -5964
rect -1122 -6010 -1118 -5964
rect -1098 -6010 -1094 -5964
rect -1085 -5971 -1080 -5964
rect -1074 -5971 -1070 -5964
rect -1075 -5985 -1070 -5971
rect -1085 -5986 -1051 -5985
rect -1050 -5986 -1046 -5961
rect -1013 -5964 -981 -5961
rect -1013 -5971 -1008 -5964
rect -995 -5965 -981 -5964
rect -978 -5965 -971 -5941
rect -1003 -5985 -998 -5971
rect -1002 -5986 -998 -5985
rect -954 -5986 -950 -5892
rect -930 -5986 -926 -5892
rect -906 -5986 -902 -5892
rect -893 -5923 -888 -5913
rect -882 -5923 -878 -5892
rect -883 -5937 -878 -5923
rect -858 -5986 -854 -5892
rect -834 -5986 -830 -5892
rect -810 -5986 -806 -5892
rect -797 -5947 -792 -5937
rect -786 -5947 -782 -5892
rect -787 -5961 -782 -5947
rect -762 -5986 -758 -5892
rect -738 -5986 -734 -5892
rect -714 -5986 -710 -5892
rect -690 -5986 -686 -5892
rect -666 -5986 -662 -5892
rect -642 -5986 -638 -5892
rect -618 -5986 -614 -5892
rect -594 -5986 -590 -5892
rect -570 -5917 -563 -5893
rect -570 -5986 -566 -5917
rect -546 -5986 -542 -5892
rect -539 -5893 -525 -5892
rect -522 -5893 -515 -5869
rect -522 -5941 -515 -5917
rect -522 -5986 -518 -5941
rect -498 -5985 -494 -5844
rect -485 -5971 -480 -5961
rect -474 -5971 -470 -5844
rect -461 -5899 -456 -5889
rect -450 -5899 -446 -5844
rect -437 -5851 -432 -5844
rect -426 -5851 -422 -5844
rect -427 -5865 -422 -5851
rect -451 -5913 -446 -5899
rect -475 -5985 -470 -5971
rect -509 -5986 -475 -5985
rect -1085 -5988 -475 -5986
rect -1085 -5995 -1080 -5988
rect -1075 -6009 -1070 -5995
rect -1074 -6010 -1070 -6009
rect -1050 -6010 -1046 -5988
rect -1002 -6010 -998 -5988
rect -954 -6010 -950 -5988
rect -930 -6010 -926 -5988
rect -906 -6010 -902 -5988
rect -858 -5989 -854 -5988
rect -1493 -6012 -861 -6010
rect -1493 -6019 -1488 -6012
rect -1483 -6033 -1478 -6019
rect -1507 -6201 -1502 -6187
rect -1517 -6211 -1512 -6201
rect -1507 -6225 -1502 -6211
rect -1506 -7402 -1502 -6225
rect -1482 -6253 -1478 -6033
rect -1458 -6061 -1454 -6012
rect -1458 -6109 -1451 -6061
rect -1482 -6301 -1475 -6253
rect -1493 -6763 -1488 -6753
rect -1482 -6763 -1478 -6301
rect -1483 -6777 -1478 -6763
rect -1493 -6787 -1488 -6777
rect -1483 -6801 -1478 -6787
rect -1482 -7402 -1478 -6801
rect -1458 -6829 -1454 -6109
rect -1445 -6811 -1440 -6801
rect -1434 -6811 -1430 -6012
rect -1435 -6825 -1430 -6811
rect -1458 -6877 -1451 -6829
rect -1445 -6835 -1440 -6825
rect -1435 -6849 -1430 -6835
rect -1458 -7402 -1454 -6877
rect -1434 -7402 -1430 -6849
rect -1410 -6877 -1406 -6012
rect -1410 -6925 -1403 -6877
rect -1421 -7363 -1416 -7353
rect -1410 -7363 -1406 -6925
rect -1411 -7377 -1406 -7363
rect -1421 -7378 -1387 -7377
rect -1386 -7378 -1382 -6012
rect -1362 -7378 -1358 -6012
rect -1338 -7378 -1334 -6012
rect -1325 -6139 -1320 -6129
rect -1314 -6139 -1310 -6012
rect -1315 -6153 -1310 -6139
rect -1325 -6163 -1320 -6153
rect -1315 -6177 -1310 -6163
rect -1314 -7378 -1310 -6177
rect -1290 -6205 -1286 -6012
rect -1290 -6253 -1283 -6205
rect -1290 -7378 -1286 -6253
rect -1277 -6547 -1272 -6537
rect -1266 -6547 -1262 -6012
rect -1267 -6561 -1262 -6547
rect -1277 -6571 -1272 -6561
rect -1267 -6585 -1262 -6571
rect -1266 -7378 -1262 -6585
rect -1242 -6613 -1238 -6012
rect -1242 -6661 -1235 -6613
rect -1242 -7378 -1238 -6661
rect -1218 -7378 -1214 -6012
rect -1194 -7378 -1190 -6012
rect -1170 -7378 -1166 -6012
rect -1146 -7378 -1142 -6012
rect -1122 -7378 -1118 -6012
rect -1098 -7378 -1094 -6012
rect -1074 -7378 -1070 -6012
rect -1050 -6037 -1046 -6012
rect -1026 -6037 -1019 -6013
rect -1050 -6085 -1043 -6037
rect -1050 -7378 -1046 -6085
rect -1026 -7378 -1022 -6037
rect -1002 -7378 -998 -6012
rect -978 -6061 -971 -6037
rect -978 -7378 -974 -6061
rect -965 -7171 -960 -7161
rect -954 -7171 -950 -6012
rect -955 -7185 -950 -7171
rect -965 -7195 -960 -7185
rect -955 -7209 -950 -7195
rect -954 -7378 -950 -7209
rect -930 -7237 -926 -6012
rect -930 -7282 -923 -7237
rect -906 -7282 -902 -6012
rect -875 -6013 -861 -6012
rect -858 -6013 -851 -5989
rect -893 -6034 -859 -6033
rect -834 -6034 -830 -5988
rect -810 -6034 -806 -5988
rect -762 -6013 -758 -5988
rect -893 -6036 -765 -6034
rect -893 -6043 -888 -6036
rect -883 -6057 -878 -6043
rect -882 -7282 -878 -6057
rect -858 -6133 -851 -6109
rect -858 -7282 -854 -6133
rect -834 -7282 -830 -6036
rect -810 -7282 -806 -6036
rect -779 -6037 -765 -6036
rect -762 -6037 -755 -6013
rect -797 -6058 -763 -6057
rect -738 -6058 -734 -5988
rect -714 -6058 -710 -5988
rect -690 -6058 -686 -5988
rect -666 -6058 -662 -5988
rect -642 -6058 -638 -5988
rect -618 -6058 -614 -5988
rect -594 -6058 -590 -5988
rect -570 -6057 -566 -5988
rect -557 -6043 -552 -6033
rect -546 -6043 -542 -5988
rect -533 -6019 -528 -6009
rect -522 -6019 -518 -5988
rect -509 -5995 -504 -5988
rect -498 -5995 -494 -5988
rect -499 -6009 -494 -5995
rect -523 -6033 -518 -6019
rect -547 -6057 -542 -6043
rect -581 -6058 -547 -6057
rect -797 -6060 -547 -6058
rect -797 -6067 -792 -6060
rect -787 -6081 -782 -6067
rect -786 -7282 -782 -6081
rect -762 -6154 -755 -6133
rect -738 -6154 -734 -6060
rect -714 -6154 -710 -6060
rect -690 -6154 -686 -6060
rect -666 -6154 -662 -6060
rect -642 -6154 -638 -6060
rect -618 -6154 -614 -6060
rect -594 -6153 -590 -6060
rect -581 -6067 -576 -6060
rect -570 -6067 -566 -6060
rect -571 -6081 -566 -6067
rect -605 -6154 -571 -6153
rect -779 -6156 -571 -6154
rect -779 -6157 -765 -6156
rect -762 -6157 -755 -6156
rect -762 -7282 -758 -6157
rect -738 -7282 -734 -6156
rect -725 -7195 -720 -7185
rect -714 -7195 -710 -6156
rect -701 -6835 -696 -6825
rect -690 -6835 -686 -6156
rect -677 -6787 -672 -6777
rect -666 -6787 -662 -6156
rect -653 -6571 -648 -6561
rect -642 -6571 -638 -6156
rect -629 -6211 -624 -6201
rect -618 -6211 -614 -6156
rect -605 -6163 -600 -6156
rect -594 -6163 -590 -6156
rect -595 -6177 -590 -6163
rect -619 -6225 -614 -6211
rect -643 -6585 -638 -6571
rect -667 -6801 -662 -6787
rect -691 -6849 -686 -6835
rect -715 -7209 -710 -7195
rect -725 -7282 -693 -7281
rect -947 -7284 -693 -7282
rect -947 -7285 -933 -7284
rect -930 -7285 -923 -7284
rect -930 -7378 -926 -7285
rect -906 -7378 -902 -7284
rect -893 -7315 -888 -7305
rect -882 -7315 -878 -7284
rect -883 -7329 -878 -7315
rect -893 -7339 -888 -7329
rect -883 -7353 -878 -7339
rect -858 -7342 -854 -7284
rect -892 -7366 -888 -7356
rect -869 -7363 -864 -7353
rect -859 -7366 -854 -7363
rect -882 -7378 -878 -7366
rect -859 -7377 -854 -7376
rect -834 -7378 -830 -7284
rect -810 -7378 -806 -7284
rect -786 -7378 -782 -7284
rect -762 -7378 -758 -7284
rect -738 -7377 -734 -7284
rect -725 -7291 -720 -7284
rect -707 -7285 -693 -7284
rect -715 -7305 -710 -7291
rect -725 -7363 -720 -7353
rect -714 -7363 -710 -7305
rect -715 -7377 -710 -7363
rect -701 -7367 -693 -7363
rect -707 -7377 -701 -7367
rect -749 -7378 -715 -7377
rect -1421 -7380 -715 -7378
rect -1421 -7387 -1416 -7380
rect -1411 -7401 -1406 -7387
rect -1410 -7402 -1406 -7401
rect -1386 -7402 -1382 -7380
rect -1362 -7402 -1358 -7380
rect -1338 -7402 -1334 -7380
rect -1314 -7402 -1310 -7380
rect -1290 -7402 -1286 -7380
rect -1266 -7402 -1262 -7380
rect -1242 -7402 -1238 -7380
rect -1218 -7402 -1214 -7380
rect -1194 -7402 -1190 -7380
rect -1170 -7402 -1166 -7380
rect -1146 -7402 -1142 -7380
rect -1122 -7402 -1118 -7380
rect -1098 -7402 -1094 -7380
rect -1074 -7402 -1070 -7380
rect -1050 -7402 -1046 -7380
rect -1026 -7402 -1022 -7380
rect -1002 -7402 -998 -7380
rect -978 -7402 -974 -7380
rect -954 -7402 -950 -7380
rect -930 -7402 -926 -7380
rect -906 -7402 -902 -7380
rect -882 -7402 -878 -7380
rect -869 -7402 -861 -7401
rect -2393 -7404 -861 -7402
rect -2371 -7426 -2366 -7404
rect -2348 -7426 -2343 -7404
rect -2325 -7426 -2320 -7404
rect -2309 -7422 -2301 -7412
rect -2068 -7421 -2062 -7416
rect -2317 -7426 -2309 -7422
rect -2060 -7426 -2050 -7421
rect -2000 -7426 -1992 -7404
rect -1806 -7412 -1680 -7406
rect -1854 -7421 -1806 -7416
rect -1655 -7422 -1647 -7412
rect -1972 -7426 -1964 -7425
rect -1958 -7426 -1942 -7424
rect -1844 -7426 -1806 -7423
rect -1663 -7426 -1655 -7422
rect -1642 -7426 -1637 -7404
rect -1619 -7426 -1614 -7404
rect -1530 -7426 -1526 -7404
rect -1506 -7426 -1502 -7404
rect -1482 -7426 -1478 -7404
rect -1458 -7426 -1454 -7404
rect -1434 -7426 -1430 -7404
rect -1410 -7426 -1406 -7404
rect -1386 -7426 -1382 -7404
rect -1362 -7426 -1358 -7404
rect -1338 -7426 -1334 -7404
rect -1314 -7426 -1310 -7404
rect -1290 -7426 -1286 -7404
rect -1266 -7426 -1262 -7404
rect -1242 -7426 -1238 -7404
rect -1218 -7426 -1214 -7404
rect -1194 -7426 -1190 -7404
rect -1170 -7426 -1166 -7404
rect -1146 -7426 -1142 -7404
rect -1122 -7426 -1118 -7404
rect -1098 -7426 -1094 -7404
rect -1074 -7426 -1070 -7404
rect -1050 -7426 -1046 -7404
rect -1026 -7426 -1022 -7404
rect -1002 -7426 -998 -7404
rect -978 -7426 -974 -7404
rect -954 -7426 -950 -7404
rect -930 -7426 -926 -7404
rect -906 -7426 -902 -7404
rect -882 -7426 -878 -7404
rect -875 -7405 -861 -7404
rect -859 -7418 -851 -7411
rect -859 -7424 -857 -7418
rect -859 -7425 -851 -7424
rect -2393 -7428 -861 -7426
rect -834 -7428 -830 -7380
rect -2371 -7450 -2366 -7428
rect -2348 -7450 -2343 -7428
rect -2325 -7450 -2320 -7428
rect -2060 -7434 -2050 -7428
rect -2309 -7450 -2301 -7440
rect -2060 -7441 -2030 -7434
rect -2000 -7438 -1992 -7428
rect -1972 -7430 -1942 -7428
rect -1958 -7431 -1942 -7430
rect -1844 -7432 -1806 -7428
rect -2068 -7448 -2062 -7441
rect -2062 -7450 -2036 -7448
rect -2393 -7452 -2036 -7450
rect -2030 -7450 -2012 -7448
rect -2004 -7450 -1990 -7438
rect -1844 -7439 -1798 -7434
rect -1806 -7441 -1798 -7439
rect -1854 -7443 -1844 -7441
rect -1854 -7448 -1806 -7443
rect -1864 -7450 -1796 -7449
rect -1655 -7450 -1647 -7440
rect -1642 -7450 -1637 -7428
rect -1619 -7450 -1614 -7428
rect -1530 -7450 -1526 -7428
rect -1506 -7450 -1502 -7428
rect -1482 -7450 -1478 -7428
rect -1458 -7450 -1454 -7428
rect -1434 -7449 -1430 -7428
rect -1445 -7450 -1411 -7449
rect -2030 -7452 -1411 -7450
rect -2371 -7498 -2366 -7452
rect -2348 -7498 -2343 -7452
rect -2325 -7498 -2320 -7452
rect -2317 -7456 -2309 -7452
rect -2060 -7456 -2050 -7452
rect -2060 -7458 -2036 -7456
rect -2060 -7460 -2030 -7458
rect -2292 -7466 -2030 -7460
rect -2092 -7482 -2062 -7480
rect -2094 -7486 -2062 -7482
rect -2000 -7498 -1992 -7452
rect -1844 -7459 -1806 -7452
rect -1663 -7456 -1655 -7452
rect -1844 -7466 -1680 -7460
rect -1854 -7482 -1806 -7480
rect -1854 -7486 -1680 -7482
rect -1642 -7498 -1637 -7452
rect -1619 -7498 -1614 -7452
rect -1530 -7498 -1526 -7452
rect -1506 -7498 -1502 -7452
rect -1482 -7498 -1478 -7452
rect -1458 -7498 -1454 -7452
rect -1445 -7459 -1440 -7452
rect -1434 -7459 -1430 -7452
rect -1435 -7473 -1430 -7459
rect -1445 -7483 -1440 -7473
rect -1435 -7497 -1430 -7483
rect -1434 -7498 -1430 -7497
rect -1410 -7498 -1406 -7428
rect -1386 -7429 -1382 -7428
rect -1386 -7474 -1379 -7429
rect -1362 -7474 -1358 -7428
rect -1338 -7474 -1334 -7428
rect -1314 -7474 -1310 -7428
rect -1290 -7474 -1286 -7428
rect -1266 -7474 -1262 -7428
rect -1242 -7474 -1238 -7428
rect -1218 -7474 -1214 -7428
rect -1194 -7474 -1190 -7428
rect -1170 -7474 -1166 -7428
rect -1146 -7474 -1142 -7428
rect -1122 -7474 -1118 -7428
rect -1098 -7474 -1094 -7428
rect -1074 -7474 -1070 -7428
rect -1050 -7474 -1046 -7428
rect -1026 -7474 -1022 -7428
rect -1002 -7474 -998 -7428
rect -978 -7474 -974 -7428
rect -954 -7474 -950 -7428
rect -930 -7474 -926 -7428
rect -906 -7474 -902 -7428
rect -882 -7474 -878 -7428
rect -875 -7429 -861 -7428
rect -858 -7429 -851 -7428
rect -858 -7474 -854 -7452
rect -834 -7453 -827 -7429
rect -810 -7474 -806 -7380
rect -786 -7473 -782 -7380
rect -773 -7435 -768 -7425
rect -762 -7435 -758 -7380
rect -749 -7387 -744 -7380
rect -738 -7387 -734 -7380
rect -739 -7401 -734 -7387
rect -763 -7449 -758 -7435
rect -797 -7474 -763 -7473
rect -1403 -7476 -763 -7474
rect -1403 -7477 -1389 -7476
rect -1386 -7477 -1379 -7476
rect -1386 -7498 -1382 -7477
rect -1362 -7498 -1358 -7476
rect -1338 -7498 -1334 -7476
rect -1314 -7498 -1310 -7476
rect -1290 -7498 -1286 -7476
rect -1266 -7498 -1262 -7476
rect -1242 -7498 -1238 -7476
rect -1218 -7498 -1214 -7476
rect -1194 -7498 -1190 -7476
rect -1170 -7498 -1166 -7476
rect -1146 -7498 -1142 -7476
rect -1122 -7498 -1118 -7476
rect -1098 -7498 -1094 -7476
rect -1074 -7498 -1070 -7476
rect -1050 -7498 -1046 -7476
rect -1026 -7498 -1022 -7476
rect -1002 -7498 -998 -7476
rect -978 -7498 -974 -7476
rect -954 -7498 -950 -7476
rect -930 -7498 -926 -7476
rect -906 -7498 -902 -7476
rect -882 -7498 -878 -7476
rect -858 -7498 -854 -7476
rect -2393 -7500 -837 -7498
rect -2371 -7522 -2366 -7500
rect -2348 -7522 -2343 -7500
rect -2325 -7522 -2320 -7500
rect -2072 -7502 -2036 -7501
rect -2072 -7508 -2054 -7502
rect -2309 -7516 -2301 -7508
rect -2317 -7522 -2309 -7516
rect -2092 -7517 -2062 -7512
rect -2000 -7521 -1992 -7500
rect -1938 -7501 -1906 -7500
rect -1920 -7502 -1906 -7501
rect -1806 -7508 -1680 -7502
rect -1854 -7517 -1806 -7512
rect -1655 -7516 -1647 -7508
rect -1982 -7521 -1966 -7520
rect -2000 -7522 -1966 -7521
rect -1846 -7522 -1806 -7519
rect -1663 -7522 -1655 -7516
rect -1642 -7522 -1637 -7500
rect -1619 -7522 -1614 -7500
rect -1530 -7522 -1526 -7500
rect -1506 -7522 -1502 -7500
rect -1482 -7522 -1478 -7500
rect -1458 -7522 -1454 -7500
rect -1434 -7522 -1430 -7500
rect -1410 -7522 -1406 -7500
rect -1386 -7522 -1382 -7500
rect -1362 -7522 -1358 -7500
rect -1338 -7522 -1334 -7500
rect -1314 -7522 -1310 -7500
rect -1290 -7522 -1286 -7500
rect -1266 -7522 -1262 -7500
rect -1242 -7522 -1238 -7500
rect -1218 -7522 -1214 -7500
rect -1194 -7522 -1190 -7500
rect -1170 -7522 -1166 -7500
rect -1146 -7522 -1142 -7500
rect -1122 -7522 -1118 -7500
rect -1098 -7522 -1094 -7500
rect -1074 -7522 -1070 -7500
rect -1050 -7522 -1046 -7500
rect -1026 -7522 -1022 -7500
rect -1002 -7522 -998 -7500
rect -978 -7522 -974 -7500
rect -954 -7522 -950 -7500
rect -930 -7522 -926 -7500
rect -906 -7521 -902 -7500
rect -917 -7522 -883 -7521
rect -2393 -7524 -883 -7522
rect -2371 -7546 -2366 -7524
rect -2348 -7546 -2343 -7524
rect -2325 -7546 -2320 -7524
rect -2000 -7526 -1966 -7524
rect -2309 -7544 -2301 -7536
rect -2062 -7537 -2054 -7530
rect -2092 -7544 -2084 -7537
rect -2062 -7544 -2026 -7542
rect -2317 -7546 -2309 -7544
rect -2062 -7546 -2012 -7544
rect -2000 -7546 -1992 -7526
rect -1982 -7527 -1966 -7526
rect -1846 -7528 -1806 -7524
rect -1846 -7535 -1798 -7530
rect -1806 -7537 -1798 -7535
rect -1854 -7539 -1846 -7537
rect -1854 -7544 -1806 -7539
rect -1655 -7544 -1647 -7536
rect -1864 -7546 -1796 -7545
rect -1663 -7546 -1655 -7544
rect -1642 -7546 -1637 -7524
rect -1619 -7546 -1614 -7524
rect -1530 -7546 -1526 -7524
rect -1506 -7546 -1502 -7524
rect -1482 -7546 -1478 -7524
rect -1458 -7546 -1454 -7524
rect -1434 -7546 -1430 -7524
rect -1410 -7525 -1406 -7524
rect -2393 -7548 -1413 -7546
rect -2371 -7594 -2366 -7548
rect -2348 -7594 -2343 -7548
rect -2325 -7584 -2320 -7548
rect -2317 -7552 -2309 -7548
rect -2062 -7552 -2054 -7548
rect -2154 -7556 -2138 -7554
rect -2057 -7556 -2054 -7552
rect -2292 -7562 -2054 -7556
rect -2052 -7562 -2044 -7552
rect -2092 -7578 -2062 -7576
rect -2094 -7582 -2062 -7578
rect -2325 -7594 -2317 -7584
rect -2095 -7592 -2084 -7588
rect -2000 -7591 -1992 -7548
rect -1846 -7555 -1806 -7548
rect -1663 -7552 -1655 -7548
rect -1846 -7562 -1680 -7556
rect -1854 -7578 -1806 -7576
rect -1854 -7582 -1680 -7578
rect -2119 -7594 -2069 -7592
rect -2054 -7594 -1892 -7591
rect -1671 -7594 -1663 -7584
rect -1642 -7594 -1637 -7548
rect -1619 -7594 -1614 -7548
rect -1530 -7593 -1526 -7548
rect -1541 -7594 -1507 -7593
rect -2393 -7596 -1507 -7594
rect -2371 -7618 -2366 -7596
rect -2348 -7618 -2343 -7596
rect -2325 -7600 -2317 -7596
rect -2325 -7616 -2320 -7600
rect -2309 -7612 -2301 -7600
rect -2095 -7602 -2084 -7596
rect -2054 -7597 -1906 -7596
rect -2054 -7598 -2036 -7597
rect -2084 -7604 -2079 -7602
rect -2317 -7616 -2309 -7612
rect -2092 -7613 -2079 -7606
rect -2000 -7610 -1992 -7597
rect -1920 -7598 -1906 -7597
rect -1671 -7600 -1663 -7596
rect -1846 -7604 -1806 -7602
rect -1854 -7610 -1806 -7606
rect -2054 -7613 -1982 -7610
rect -1966 -7613 -1806 -7610
rect -1655 -7612 -1647 -7600
rect -2003 -7616 -1992 -7613
rect -1904 -7615 -1902 -7613
rect -1854 -7615 -1846 -7613
rect -2325 -7618 -2317 -7616
rect -2033 -7618 -1992 -7616
rect -1854 -7617 -1806 -7615
rect -1663 -7616 -1655 -7612
rect -1864 -7618 -1796 -7617
rect -1671 -7618 -1663 -7616
rect -1642 -7618 -1637 -7596
rect -1619 -7618 -1614 -7596
rect -1541 -7603 -1536 -7596
rect -1530 -7603 -1526 -7596
rect -1531 -7617 -1526 -7603
rect -1506 -7618 -1502 -7548
rect -1482 -7618 -1478 -7548
rect -1458 -7618 -1454 -7548
rect -1434 -7617 -1430 -7548
rect -1427 -7549 -1413 -7548
rect -1410 -7573 -1403 -7525
rect -1445 -7618 -1411 -7617
rect -2393 -7620 -1411 -7618
rect -2371 -7642 -2366 -7620
rect -2348 -7642 -2343 -7620
rect -2325 -7628 -2317 -7620
rect -2079 -7623 -2018 -7620
rect -2003 -7621 -1966 -7620
rect -2000 -7622 -1982 -7621
rect -2000 -7623 -1992 -7622
rect -2084 -7627 -2009 -7623
rect -2028 -7628 -2009 -7627
rect -2000 -7627 -1854 -7623
rect -1846 -7627 -1798 -7620
rect -2325 -7642 -2320 -7628
rect -2309 -7640 -2301 -7628
rect -2028 -7630 -2018 -7628
rect -2092 -7640 -2084 -7633
rect -2023 -7637 -2014 -7630
rect -2000 -7637 -1992 -7627
rect -1671 -7628 -1663 -7620
rect -1846 -7631 -1806 -7629
rect -1854 -7637 -1806 -7633
rect -2054 -7640 -1806 -7637
rect -1655 -7640 -1647 -7628
rect -2317 -7642 -2309 -7640
rect -2054 -7642 -2024 -7640
rect -2000 -7642 -1992 -7640
rect -1663 -7642 -1655 -7640
rect -1642 -7642 -1637 -7620
rect -1619 -7642 -1614 -7620
rect -1506 -7642 -1502 -7620
rect -1482 -7642 -1478 -7620
rect -1458 -7642 -1454 -7620
rect -1445 -7627 -1440 -7620
rect -1434 -7627 -1430 -7620
rect -1435 -7641 -1430 -7627
rect -1410 -7642 -1406 -7573
rect -1386 -7642 -1382 -7524
rect -1362 -7642 -1358 -7524
rect -1338 -7642 -1334 -7524
rect -1314 -7641 -1310 -7524
rect -1325 -7642 -1291 -7641
rect -2393 -7644 -2064 -7642
rect -2060 -7644 -1291 -7642
rect -2371 -7690 -2366 -7644
rect -2348 -7690 -2343 -7644
rect -2325 -7656 -2317 -7644
rect -2060 -7647 -2054 -7644
rect -2084 -7654 -2054 -7647
rect -2050 -7650 -2044 -7648
rect -2325 -7676 -2320 -7656
rect -2064 -7658 -2054 -7654
rect -2325 -7684 -2317 -7676
rect -2101 -7681 -2071 -7678
rect -2325 -7690 -2320 -7684
rect -2317 -7690 -2309 -7684
rect -2000 -7686 -1992 -7644
rect -1846 -7645 -1806 -7644
rect -1846 -7654 -1798 -7647
rect -1671 -7656 -1663 -7644
rect -1846 -7658 -1806 -7656
rect -1854 -7672 -1680 -7668
rect -1846 -7681 -1798 -7678
rect -2079 -7687 -2043 -7686
rect -2007 -7687 -1991 -7686
rect -2079 -7688 -2071 -7687
rect -2079 -7690 -2029 -7688
rect -2011 -7690 -1991 -7687
rect -1846 -7689 -1806 -7683
rect -1671 -7684 -1663 -7676
rect -1864 -7690 -1796 -7689
rect -1663 -7690 -1655 -7684
rect -1642 -7690 -1637 -7644
rect -1619 -7690 -1614 -7644
rect -1506 -7669 -1502 -7644
rect -2393 -7692 -1509 -7690
rect -2371 -7738 -2366 -7692
rect -2348 -7738 -2343 -7692
rect -2325 -7704 -2320 -7692
rect -2079 -7694 -2071 -7692
rect -2072 -7696 -2071 -7694
rect -2109 -7701 -2101 -7696
rect -2101 -7703 -2079 -7701
rect -2069 -7703 -2068 -7696
rect -2325 -7712 -2317 -7704
rect -2079 -7708 -2071 -7703
rect -2325 -7732 -2320 -7712
rect -2317 -7720 -2309 -7712
rect -2074 -7717 -2071 -7708
rect -2069 -7712 -2068 -7708
rect -2109 -7726 -2079 -7723
rect -2325 -7738 -2317 -7732
rect -2119 -7738 -2069 -7736
rect -2056 -7738 -2026 -7735
rect -2000 -7738 -1992 -7692
rect -1846 -7694 -1806 -7692
rect -1854 -7699 -1806 -7695
rect -1854 -7701 -1846 -7699
rect -1846 -7703 -1806 -7701
rect -1806 -7705 -1798 -7703
rect -1846 -7708 -1798 -7705
rect -1846 -7721 -1806 -7710
rect -1671 -7712 -1663 -7704
rect -1663 -7720 -1655 -7712
rect -1854 -7726 -1680 -7722
rect -1926 -7738 -1892 -7735
rect -1671 -7738 -1663 -7732
rect -1642 -7738 -1637 -7692
rect -1619 -7738 -1614 -7692
rect -1523 -7693 -1509 -7692
rect -1506 -7693 -1499 -7669
rect -1541 -7714 -1507 -7713
rect -1482 -7714 -1478 -7644
rect -1469 -7675 -1464 -7665
rect -1458 -7675 -1454 -7644
rect -1445 -7675 -1440 -7665
rect -1459 -7689 -1454 -7675
rect -1435 -7689 -1430 -7675
rect -1434 -7714 -1430 -7689
rect -1410 -7693 -1406 -7644
rect -1541 -7716 -1413 -7714
rect -1541 -7723 -1536 -7716
rect -1531 -7737 -1526 -7723
rect -1530 -7738 -1526 -7737
rect -1482 -7738 -1478 -7716
rect -1434 -7738 -1430 -7716
rect -1427 -7717 -1413 -7716
rect -1410 -7717 -1403 -7693
rect -1386 -7738 -1382 -7644
rect -1362 -7738 -1358 -7644
rect -1338 -7737 -1334 -7644
rect -1325 -7651 -1320 -7644
rect -1314 -7651 -1310 -7644
rect -1315 -7665 -1310 -7651
rect -1290 -7717 -1286 -7524
rect -1349 -7738 -1293 -7737
rect -2393 -7740 -1293 -7738
rect -2371 -7762 -2366 -7740
rect -2348 -7762 -2343 -7740
rect -2325 -7744 -2317 -7740
rect -2325 -7760 -2320 -7744
rect -2317 -7748 -2309 -7744
rect -2309 -7760 -2301 -7748
rect -2109 -7757 -2079 -7750
rect -2000 -7751 -1992 -7740
rect -1671 -7744 -1663 -7740
rect -1846 -7748 -1806 -7746
rect -1663 -7748 -1655 -7744
rect -2009 -7754 -1992 -7751
rect -1854 -7754 -1806 -7750
rect -2071 -7757 -1992 -7754
rect -1983 -7757 -1806 -7754
rect -2009 -7760 -1992 -7757
rect -2325 -7762 -2317 -7760
rect -2033 -7762 -1992 -7760
rect -1846 -7761 -1806 -7759
rect -1655 -7760 -1647 -7748
rect -1864 -7762 -1796 -7761
rect -1671 -7762 -1663 -7760
rect -1642 -7762 -1637 -7740
rect -1619 -7762 -1614 -7740
rect -1530 -7762 -1526 -7740
rect -1482 -7762 -1478 -7740
rect -1434 -7741 -1430 -7740
rect -1434 -7762 -1427 -7741
rect -1410 -7762 -1403 -7741
rect -1386 -7762 -1382 -7740
rect -1362 -7762 -1358 -7740
rect -1349 -7747 -1344 -7740
rect -1338 -7747 -1334 -7740
rect -1325 -7747 -1320 -7740
rect -1307 -7741 -1293 -7740
rect -1290 -7741 -1283 -7717
rect -1339 -7761 -1334 -7747
rect -1315 -7761 -1310 -7747
rect -1314 -7762 -1310 -7761
rect -1266 -7762 -1262 -7524
rect -1242 -7762 -1238 -7524
rect -1218 -7762 -1214 -7524
rect -1194 -7762 -1190 -7524
rect -1170 -7761 -1166 -7524
rect -1181 -7762 -1147 -7761
rect -2393 -7764 -1437 -7762
rect -2371 -7786 -2366 -7764
rect -2348 -7786 -2343 -7764
rect -2325 -7772 -2317 -7764
rect -2079 -7767 -2035 -7764
rect -2013 -7766 -1992 -7764
rect -2000 -7767 -1992 -7766
rect -1904 -7767 -1798 -7764
rect -2101 -7771 -2009 -7767
rect -2023 -7772 -2009 -7771
rect -2000 -7769 -1798 -7767
rect -2000 -7771 -1854 -7769
rect -1846 -7771 -1798 -7769
rect -2325 -7786 -2320 -7772
rect -2317 -7776 -2309 -7772
rect -2309 -7786 -2301 -7776
rect -2109 -7784 -2101 -7777
rect -2023 -7781 -2021 -7772
rect -2000 -7781 -1992 -7771
rect -1671 -7772 -1663 -7764
rect -1846 -7775 -1806 -7773
rect -1663 -7776 -1655 -7772
rect -1854 -7781 -1806 -7777
rect -2071 -7784 -1806 -7781
rect -2074 -7786 -2031 -7784
rect -2000 -7786 -1992 -7784
rect -1655 -7786 -1647 -7776
rect -1642 -7786 -1637 -7764
rect -1619 -7786 -1614 -7764
rect -1530 -7786 -1526 -7764
rect -1482 -7786 -1478 -7764
rect -1451 -7765 -1437 -7764
rect -1434 -7764 -1147 -7762
rect -1434 -7765 -1413 -7764
rect -1410 -7765 -1403 -7764
rect -1410 -7786 -1406 -7765
rect -1386 -7786 -1382 -7764
rect -1362 -7786 -1358 -7764
rect -1314 -7786 -1310 -7764
rect -1266 -7786 -1262 -7764
rect -1242 -7786 -1238 -7764
rect -1218 -7786 -1214 -7764
rect -1194 -7786 -1190 -7764
rect -1181 -7771 -1176 -7764
rect -1170 -7771 -1166 -7764
rect -1171 -7785 -1166 -7771
rect -1146 -7786 -1142 -7524
rect -1122 -7786 -1118 -7524
rect -1098 -7786 -1094 -7524
rect -1074 -7786 -1070 -7524
rect -1050 -7786 -1046 -7524
rect -1026 -7786 -1022 -7524
rect -1002 -7785 -998 -7524
rect -989 -7699 -984 -7689
rect -978 -7699 -974 -7524
rect -965 -7555 -960 -7545
rect -954 -7555 -950 -7524
rect -955 -7569 -950 -7555
rect -965 -7570 -931 -7569
rect -930 -7570 -926 -7524
rect -917 -7531 -912 -7524
rect -906 -7531 -902 -7524
rect -907 -7545 -902 -7531
rect -917 -7555 -912 -7545
rect -907 -7569 -902 -7555
rect -906 -7570 -902 -7569
rect -882 -7570 -878 -7500
rect -858 -7570 -854 -7500
rect -851 -7501 -837 -7500
rect -834 -7501 -827 -7477
rect -834 -7570 -830 -7501
rect -810 -7569 -806 -7476
rect -797 -7483 -792 -7476
rect -786 -7483 -782 -7476
rect -787 -7497 -782 -7483
rect -797 -7507 -792 -7497
rect -787 -7521 -782 -7507
rect -797 -7555 -792 -7545
rect -786 -7555 -782 -7521
rect -787 -7569 -782 -7555
rect -773 -7559 -765 -7555
rect -779 -7569 -773 -7559
rect -821 -7570 -787 -7569
rect -965 -7572 -787 -7570
rect -965 -7579 -960 -7572
rect -955 -7593 -950 -7579
rect -979 -7713 -974 -7699
rect -989 -7762 -955 -7761
rect -954 -7762 -950 -7593
rect -930 -7621 -926 -7572
rect -930 -7666 -923 -7621
rect -906 -7666 -902 -7572
rect -882 -7597 -878 -7572
rect -882 -7645 -875 -7597
rect -882 -7666 -878 -7645
rect -858 -7666 -854 -7572
rect -834 -7665 -830 -7572
rect -821 -7579 -816 -7572
rect -810 -7579 -806 -7572
rect -811 -7593 -806 -7579
rect -845 -7666 -811 -7665
rect -947 -7668 -811 -7666
rect -947 -7669 -933 -7668
rect -930 -7669 -923 -7668
rect -930 -7762 -926 -7669
rect -906 -7761 -902 -7668
rect -893 -7747 -888 -7737
rect -882 -7747 -878 -7668
rect -869 -7723 -864 -7713
rect -858 -7723 -854 -7668
rect -845 -7675 -840 -7668
rect -834 -7675 -830 -7668
rect -835 -7689 -830 -7675
rect -859 -7737 -854 -7723
rect -883 -7761 -878 -7747
rect -917 -7762 -883 -7761
rect -989 -7764 -883 -7762
rect -989 -7771 -984 -7764
rect -954 -7765 -950 -7764
rect -979 -7785 -974 -7771
rect -965 -7775 -957 -7771
rect -971 -7785 -965 -7775
rect -1013 -7786 -979 -7785
rect -2393 -7788 -979 -7786
rect -2371 -7834 -2366 -7788
rect -2348 -7834 -2343 -7788
rect -2325 -7800 -2317 -7788
rect -2074 -7791 -2071 -7788
rect -2101 -7798 -2071 -7791
rect -2325 -7820 -2320 -7800
rect -2317 -7804 -2309 -7800
rect -2064 -7802 -2061 -7794
rect -2325 -7828 -2317 -7820
rect -2101 -7825 -2071 -7822
rect -2325 -7834 -2320 -7828
rect -2317 -7834 -2309 -7828
rect -2000 -7830 -1992 -7788
rect -1846 -7789 -1806 -7788
rect -1846 -7798 -1798 -7791
rect -1671 -7800 -1663 -7788
rect -1846 -7802 -1806 -7800
rect -1663 -7804 -1655 -7800
rect -1854 -7816 -1680 -7812
rect -1846 -7825 -1798 -7822
rect -2079 -7831 -2043 -7830
rect -2007 -7831 -1991 -7830
rect -2079 -7832 -2071 -7831
rect -2079 -7834 -2029 -7832
rect -2011 -7834 -1991 -7831
rect -1846 -7833 -1806 -7827
rect -1671 -7828 -1663 -7820
rect -1864 -7834 -1796 -7833
rect -1663 -7834 -1655 -7828
rect -1642 -7834 -1637 -7788
rect -1619 -7834 -1614 -7788
rect -1530 -7834 -1526 -7788
rect -1506 -7810 -1499 -7789
rect -1482 -7810 -1478 -7788
rect -1410 -7810 -1406 -7788
rect -1386 -7810 -1382 -7788
rect -1362 -7810 -1358 -7788
rect -1314 -7810 -1310 -7788
rect -1266 -7810 -1262 -7788
rect -1242 -7810 -1238 -7788
rect -1218 -7810 -1214 -7788
rect -1194 -7810 -1190 -7788
rect -1181 -7810 -1147 -7809
rect -1523 -7812 -1147 -7810
rect -1523 -7813 -1509 -7812
rect -1506 -7813 -1499 -7812
rect -1506 -7834 -1502 -7813
rect -1482 -7834 -1478 -7812
rect -1410 -7834 -1406 -7812
rect -1386 -7834 -1382 -7812
rect -1362 -7834 -1358 -7812
rect -1314 -7813 -1310 -7812
rect -1314 -7834 -1307 -7813
rect -1290 -7833 -1283 -7813
rect -1301 -7834 -1267 -7833
rect -2393 -7836 -1317 -7834
rect -2371 -7882 -2366 -7836
rect -2348 -7882 -2343 -7836
rect -2325 -7848 -2320 -7836
rect -2079 -7838 -2071 -7836
rect -2072 -7840 -2071 -7838
rect -2109 -7845 -2101 -7840
rect -2101 -7847 -2079 -7845
rect -2069 -7847 -2068 -7840
rect -2325 -7856 -2317 -7848
rect -2079 -7852 -2071 -7847
rect -2325 -7876 -2320 -7856
rect -2317 -7864 -2309 -7856
rect -2074 -7861 -2071 -7852
rect -2069 -7856 -2068 -7852
rect -2109 -7870 -2079 -7867
rect -2325 -7882 -2317 -7876
rect -2119 -7882 -2069 -7880
rect -2056 -7882 -2026 -7879
rect -2000 -7882 -1992 -7836
rect -1846 -7838 -1806 -7836
rect -1854 -7843 -1806 -7839
rect -1854 -7845 -1846 -7843
rect -1846 -7847 -1806 -7845
rect -1806 -7849 -1798 -7847
rect -1846 -7852 -1798 -7849
rect -1846 -7865 -1806 -7854
rect -1671 -7856 -1663 -7848
rect -1663 -7864 -1655 -7856
rect -1854 -7870 -1680 -7866
rect -1926 -7882 -1892 -7879
rect -1671 -7882 -1663 -7876
rect -1642 -7882 -1637 -7836
rect -1619 -7882 -1614 -7836
rect -1530 -7882 -1526 -7836
rect -1506 -7882 -1502 -7836
rect -1482 -7882 -1478 -7836
rect -1469 -7858 -1435 -7857
rect -1410 -7858 -1406 -7836
rect -1386 -7858 -1382 -7836
rect -1362 -7858 -1358 -7836
rect -1331 -7837 -1317 -7836
rect -1314 -7836 -1267 -7834
rect -1314 -7837 -1293 -7836
rect -1290 -7837 -1283 -7836
rect -1301 -7843 -1296 -7837
rect -1290 -7843 -1286 -7837
rect -1291 -7857 -1286 -7843
rect -1266 -7858 -1262 -7812
rect -1242 -7858 -1238 -7812
rect -1218 -7858 -1214 -7812
rect -1194 -7858 -1190 -7812
rect -1181 -7819 -1176 -7812
rect -1171 -7833 -1166 -7819
rect -1146 -7822 -1142 -7788
rect -1157 -7834 -1123 -7833
rect -1122 -7834 -1118 -7788
rect -1098 -7834 -1094 -7788
rect -1074 -7834 -1070 -7788
rect -1050 -7834 -1046 -7788
rect -1026 -7834 -1022 -7788
rect -1013 -7795 -1008 -7788
rect -1002 -7795 -998 -7788
rect -1003 -7809 -998 -7795
rect -1013 -7810 -979 -7809
rect -978 -7810 -974 -7785
rect -954 -7789 -947 -7765
rect -930 -7809 -926 -7764
rect -917 -7771 -912 -7764
rect -906 -7771 -902 -7764
rect -907 -7785 -902 -7771
rect -941 -7810 -907 -7809
rect -1013 -7812 -907 -7810
rect -1013 -7819 -1008 -7812
rect -1003 -7833 -998 -7819
rect -1002 -7834 -998 -7833
rect -978 -7834 -974 -7812
rect -941 -7819 -936 -7812
rect -930 -7819 -926 -7812
rect -931 -7833 -926 -7819
rect -965 -7834 -931 -7833
rect -1157 -7836 -931 -7834
rect -1180 -7846 -1176 -7836
rect -1157 -7843 -1152 -7836
rect -1170 -7858 -1166 -7846
rect -1147 -7857 -1139 -7843
rect -1469 -7860 -1149 -7858
rect -1469 -7867 -1464 -7860
rect -1459 -7881 -1454 -7867
rect -1458 -7882 -1454 -7881
rect -1410 -7882 -1406 -7860
rect -1386 -7882 -1382 -7860
rect -1362 -7882 -1358 -7860
rect -1301 -7882 -1267 -7881
rect -2393 -7884 -1267 -7882
rect -2371 -7906 -2366 -7884
rect -2348 -7906 -2343 -7884
rect -2325 -7888 -2317 -7884
rect -2325 -7904 -2320 -7888
rect -2317 -7892 -2309 -7888
rect -2309 -7904 -2301 -7892
rect -2109 -7901 -2079 -7894
rect -2000 -7895 -1992 -7884
rect -1671 -7888 -1663 -7884
rect -1846 -7892 -1806 -7890
rect -1663 -7892 -1655 -7888
rect -2009 -7898 -1992 -7895
rect -1854 -7898 -1806 -7894
rect -2071 -7901 -1992 -7898
rect -1983 -7901 -1806 -7898
rect -2009 -7904 -1992 -7901
rect -2325 -7906 -2317 -7904
rect -2033 -7906 -1992 -7904
rect -1846 -7905 -1806 -7903
rect -1655 -7904 -1647 -7892
rect -1864 -7906 -1796 -7905
rect -1671 -7906 -1663 -7904
rect -1642 -7906 -1637 -7884
rect -1619 -7906 -1614 -7884
rect -1530 -7906 -1526 -7884
rect -1506 -7906 -1502 -7884
rect -1482 -7906 -1478 -7884
rect -1458 -7906 -1454 -7884
rect -1410 -7906 -1406 -7884
rect -1386 -7906 -1382 -7884
rect -1362 -7906 -1358 -7884
rect -1301 -7891 -1296 -7884
rect -1291 -7905 -1286 -7891
rect -1266 -7894 -1262 -7860
rect -1242 -7906 -1238 -7860
rect -1218 -7906 -1214 -7860
rect -1194 -7906 -1190 -7860
rect -1170 -7906 -1166 -7860
rect -1163 -7861 -1149 -7860
rect -1157 -7882 -1123 -7881
rect -1122 -7882 -1118 -7836
rect -1098 -7882 -1094 -7836
rect -1074 -7882 -1070 -7836
rect -1050 -7882 -1046 -7836
rect -1026 -7882 -1022 -7836
rect -1002 -7881 -998 -7836
rect -989 -7867 -984 -7857
rect -978 -7861 -974 -7836
rect -954 -7843 -947 -7837
rect -955 -7857 -947 -7843
rect -971 -7860 -955 -7857
rect -971 -7861 -957 -7860
rect -978 -7867 -971 -7861
rect -979 -7881 -971 -7867
rect -1013 -7882 -981 -7881
rect -1157 -7884 -981 -7882
rect -1147 -7905 -1139 -7891
rect -2393 -7908 -1149 -7906
rect -1122 -7908 -1118 -7884
rect -2371 -7930 -2366 -7908
rect -2348 -7930 -2343 -7908
rect -2325 -7916 -2317 -7908
rect -2079 -7911 -2035 -7908
rect -2013 -7910 -1992 -7908
rect -2000 -7911 -1992 -7910
rect -1904 -7911 -1798 -7908
rect -2101 -7915 -2009 -7911
rect -2023 -7916 -2009 -7915
rect -2000 -7913 -1798 -7911
rect -2000 -7915 -1854 -7913
rect -1846 -7915 -1798 -7913
rect -2325 -7930 -2320 -7916
rect -2317 -7920 -2309 -7916
rect -2309 -7930 -2301 -7920
rect -2109 -7928 -2101 -7921
rect -2023 -7925 -2021 -7916
rect -2000 -7925 -1992 -7915
rect -1671 -7916 -1663 -7908
rect -1846 -7919 -1806 -7917
rect -1663 -7920 -1655 -7916
rect -1854 -7925 -1806 -7921
rect -2071 -7928 -1806 -7925
rect -2074 -7930 -2031 -7928
rect -2000 -7930 -1992 -7928
rect -1655 -7930 -1647 -7920
rect -1642 -7930 -1637 -7908
rect -1619 -7930 -1614 -7908
rect -1530 -7930 -1526 -7908
rect -1506 -7930 -1502 -7908
rect -1482 -7930 -1478 -7908
rect -1458 -7930 -1454 -7908
rect -1410 -7930 -1406 -7908
rect -1386 -7930 -1382 -7908
rect -1362 -7930 -1358 -7908
rect -2393 -7932 -1269 -7930
rect -2371 -7978 -2366 -7932
rect -2348 -7978 -2343 -7932
rect -2325 -7944 -2317 -7932
rect -2074 -7935 -2071 -7932
rect -2101 -7942 -2071 -7935
rect -2325 -7964 -2320 -7944
rect -2317 -7948 -2309 -7944
rect -2064 -7946 -2061 -7938
rect -2325 -7972 -2317 -7964
rect -2101 -7969 -2071 -7966
rect -2325 -7978 -2320 -7972
rect -2317 -7978 -2309 -7972
rect -2000 -7974 -1992 -7932
rect -1846 -7933 -1806 -7932
rect -1846 -7942 -1798 -7935
rect -1671 -7944 -1663 -7932
rect -1846 -7946 -1806 -7944
rect -1663 -7948 -1655 -7944
rect -1854 -7960 -1680 -7956
rect -1846 -7969 -1798 -7966
rect -2079 -7975 -2043 -7974
rect -2007 -7975 -1991 -7974
rect -2079 -7976 -2071 -7975
rect -2079 -7978 -2029 -7976
rect -2011 -7978 -1991 -7975
rect -1846 -7977 -1806 -7971
rect -1671 -7972 -1663 -7964
rect -1864 -7978 -1796 -7977
rect -1663 -7978 -1655 -7972
rect -1642 -7978 -1637 -7932
rect -1619 -7978 -1614 -7932
rect -1589 -7978 -1555 -7977
rect -2393 -7980 -1555 -7978
rect -2371 -8026 -2366 -7980
rect -2348 -8026 -2343 -7980
rect -2325 -7992 -2320 -7980
rect -2079 -7982 -2071 -7980
rect -2072 -7984 -2071 -7982
rect -2109 -7989 -2101 -7984
rect -2101 -7991 -2079 -7989
rect -2069 -7991 -2068 -7984
rect -2325 -8000 -2317 -7992
rect -2079 -7996 -2071 -7991
rect -2325 -8020 -2320 -8000
rect -2317 -8008 -2309 -8000
rect -2074 -8005 -2071 -7996
rect -2069 -8000 -2068 -7996
rect -2109 -8014 -2079 -8011
rect -2325 -8026 -2317 -8020
rect -2080 -8026 -2071 -8025
rect -2000 -8026 -1992 -7980
rect -1846 -7982 -1806 -7980
rect -1854 -7987 -1806 -7983
rect -1854 -7989 -1846 -7987
rect -1846 -7991 -1806 -7989
rect -1806 -7993 -1798 -7991
rect -1846 -7996 -1798 -7993
rect -1846 -8009 -1806 -7998
rect -1671 -8000 -1663 -7992
rect -1663 -8008 -1655 -8000
rect -1854 -8014 -1680 -8010
rect -1926 -8026 -1892 -8023
rect -1671 -8026 -1663 -8020
rect -1642 -8026 -1637 -7980
rect -1619 -8026 -1614 -7980
rect -1565 -8002 -1531 -8001
rect -1530 -8002 -1526 -7932
rect -1506 -8002 -1502 -7932
rect -1482 -8002 -1478 -7932
rect -1458 -8002 -1454 -7932
rect -1434 -7954 -1427 -7933
rect -1410 -7954 -1406 -7932
rect -1386 -7954 -1382 -7932
rect -1362 -7954 -1358 -7932
rect -1283 -7933 -1269 -7932
rect -1242 -7954 -1238 -7908
rect -1218 -7954 -1214 -7908
rect -1194 -7954 -1190 -7908
rect -1170 -7954 -1166 -7908
rect -1163 -7909 -1149 -7908
rect -1146 -7909 -1139 -7908
rect -1122 -7930 -1115 -7909
rect -1098 -7929 -1094 -7884
rect -1109 -7930 -1075 -7929
rect -1139 -7932 -1075 -7930
rect -1146 -7954 -1142 -7932
rect -1139 -7933 -1125 -7932
rect -1122 -7933 -1115 -7932
rect -1109 -7939 -1104 -7932
rect -1098 -7939 -1094 -7932
rect -1099 -7953 -1094 -7939
rect -1109 -7954 -1075 -7953
rect -1451 -7956 -1075 -7954
rect -1451 -7957 -1437 -7956
rect -1434 -7957 -1427 -7956
rect -1434 -8002 -1430 -7957
rect -1410 -8002 -1406 -7956
rect -1386 -8002 -1382 -7956
rect -1362 -8002 -1358 -7956
rect -1349 -7978 -1315 -7977
rect -1349 -7980 -1269 -7978
rect -1242 -7980 -1238 -7956
rect -1349 -7987 -1344 -7980
rect -1283 -7981 -1269 -7980
rect -1339 -8001 -1334 -7987
rect -1338 -8002 -1334 -8001
rect -1218 -8002 -1214 -7956
rect -1194 -8002 -1190 -7956
rect -1170 -8002 -1166 -7956
rect -1146 -8002 -1142 -7956
rect -1122 -7978 -1115 -7957
rect -1109 -7963 -1104 -7956
rect -1099 -7977 -1094 -7963
rect -1074 -7966 -1070 -7884
rect -1061 -7915 -1056 -7905
rect -1050 -7915 -1046 -7884
rect -1051 -7929 -1046 -7915
rect -1060 -7942 -1056 -7932
rect -1026 -7942 -1022 -7884
rect -1013 -7891 -1008 -7884
rect -1002 -7891 -998 -7884
rect -995 -7885 -981 -7884
rect -1003 -7905 -998 -7891
rect -989 -7895 -981 -7891
rect -995 -7905 -989 -7895
rect -1109 -7978 -1075 -7977
rect -1139 -7980 -1075 -7978
rect -1139 -7981 -1125 -7980
rect -1122 -7981 -1115 -7980
rect -1122 -8001 -1118 -7981
rect -1109 -7987 -1104 -7980
rect -1099 -8001 -1094 -7987
rect -1050 -7990 -1046 -7942
rect -1133 -8002 -1099 -8001
rect -1565 -8004 -1099 -8002
rect -1530 -8026 -1526 -8004
rect -1506 -8026 -1502 -8004
rect -1482 -8026 -1478 -8004
rect -1458 -8026 -1454 -8004
rect -1434 -8026 -1430 -8004
rect -1410 -8026 -1406 -8004
rect -1386 -8025 -1382 -8004
rect -1397 -8026 -1363 -8025
rect -2393 -8028 -1363 -8026
rect -2371 -8050 -2366 -8028
rect -2348 -8050 -2343 -8028
rect -2325 -8034 -2317 -8028
rect -2325 -8050 -2320 -8034
rect -2317 -8036 -2309 -8034
rect -2309 -8048 -2301 -8036
rect -2080 -8037 -2071 -8028
rect -2068 -8038 -2059 -8037
rect -2068 -8045 -2038 -8038
rect -2317 -8050 -2309 -8048
rect -2068 -8050 -2059 -8045
rect -2000 -8046 -1992 -8028
rect -1846 -8036 -1794 -8028
rect -1671 -8034 -1663 -8028
rect -1663 -8036 -1655 -8034
rect -1852 -8045 -1804 -8038
rect -2011 -8048 -1983 -8046
rect -2025 -8049 -1983 -8048
rect -2025 -8050 -1975 -8049
rect -1846 -8050 -1804 -8047
rect -1655 -8048 -1647 -8036
rect -1663 -8050 -1655 -8048
rect -1642 -8050 -1637 -8028
rect -1619 -8050 -1614 -8028
rect -1530 -8050 -1526 -8028
rect -1506 -8050 -1502 -8028
rect -1482 -8050 -1478 -8028
rect -1458 -8050 -1454 -8028
rect -1434 -8050 -1430 -8028
rect -1410 -8050 -1406 -8028
rect -1397 -8035 -1392 -8028
rect -1386 -8035 -1382 -8028
rect -1387 -8049 -1382 -8035
rect -1397 -8050 -1363 -8049
rect -1362 -8050 -1358 -8004
rect -1338 -8050 -1334 -8004
rect -1277 -8026 -1243 -8025
rect -1218 -8026 -1214 -8004
rect -1194 -8026 -1190 -8004
rect -1170 -8026 -1166 -8004
rect -1146 -8025 -1142 -8004
rect -1133 -8011 -1128 -8004
rect -1122 -8011 -1118 -8004
rect -1123 -8025 -1118 -8011
rect -1157 -8026 -1123 -8025
rect -1277 -8028 -1123 -8026
rect -1300 -8038 -1296 -8028
rect -1290 -8050 -1286 -8038
rect -1277 -8050 -1243 -8049
rect -2393 -8052 -1243 -8050
rect -2371 -8074 -2366 -8052
rect -2348 -8074 -2343 -8052
rect -2325 -8062 -2317 -8052
rect -2068 -8053 -2038 -8052
rect -2068 -8055 -2059 -8053
rect -2013 -8054 -1983 -8052
rect -1846 -8053 -1804 -8052
rect -2000 -8055 -1983 -8054
rect -1862 -8055 -1798 -8054
rect -2076 -8062 -2068 -8055
rect -2061 -8062 -2045 -8060
rect -2038 -8062 -2001 -8055
rect -2325 -8074 -2320 -8062
rect -2317 -8064 -2309 -8062
rect -2309 -8074 -2301 -8064
rect -2068 -8065 -2045 -8062
rect -2015 -8063 -2001 -8062
rect -2068 -8072 -2038 -8065
rect -2068 -8074 -2045 -8072
rect -2000 -8074 -1992 -8055
rect -1985 -8057 -1796 -8055
rect -1985 -8062 -1852 -8057
rect -1846 -8062 -1796 -8057
rect -1671 -8062 -1663 -8052
rect -1846 -8063 -1798 -8062
rect -1663 -8064 -1655 -8062
rect -1852 -8072 -1804 -8065
rect -1976 -8074 -1940 -8073
rect -1655 -8074 -1647 -8064
rect -1642 -8074 -1637 -8052
rect -1619 -8074 -1614 -8052
rect -1554 -8066 -1547 -8053
rect -2393 -8076 -1557 -8074
rect -1530 -8076 -1526 -8052
rect -2371 -8146 -2366 -8076
rect -2348 -8146 -2343 -8076
rect -2325 -8078 -2320 -8076
rect -2317 -8078 -2309 -8076
rect -2325 -8090 -2317 -8078
rect -2068 -8082 -2059 -8076
rect -2076 -8089 -2071 -8082
rect -2068 -8090 -2059 -8089
rect -2325 -8110 -2320 -8090
rect -2317 -8092 -2309 -8090
rect -2325 -8118 -2317 -8110
rect -2060 -8116 -2030 -8113
rect -2325 -8146 -2320 -8118
rect -2317 -8126 -2309 -8118
rect -2060 -8129 -2038 -8118
rect -2033 -8125 -2030 -8116
rect -2028 -8120 -2027 -8116
rect -2068 -8134 -2038 -8131
rect -2000 -8146 -1992 -8076
rect -1846 -8080 -1804 -8076
rect -1663 -8078 -1655 -8076
rect -1846 -8090 -1794 -8081
rect -1671 -8090 -1663 -8078
rect -1663 -8092 -1655 -8090
rect -1912 -8101 -1884 -8099
rect -1852 -8107 -1804 -8103
rect -1844 -8116 -1796 -8113
rect -1671 -8118 -1663 -8110
rect -1844 -8129 -1804 -8118
rect -1663 -8126 -1655 -8118
rect -1852 -8134 -1680 -8130
rect -1642 -8146 -1637 -8076
rect -1619 -8146 -1614 -8076
rect -1571 -8077 -1557 -8076
rect -1554 -8077 -1547 -8076
rect -1530 -8097 -1523 -8077
rect -1541 -8098 -1507 -8097
rect -1547 -8100 -1507 -8098
rect -1547 -8101 -1533 -8100
rect -1530 -8101 -1523 -8100
rect -1541 -8107 -1536 -8101
rect -1530 -8107 -1526 -8101
rect -1531 -8121 -1526 -8107
rect -1541 -8122 -1507 -8121
rect -1506 -8122 -1502 -8052
rect -1482 -8122 -1478 -8052
rect -1458 -8122 -1454 -8052
rect -1434 -8122 -1430 -8052
rect -1410 -8122 -1406 -8052
rect -1397 -8059 -1392 -8052
rect -1387 -8073 -1382 -8059
rect -1386 -8122 -1382 -8073
rect -1362 -8101 -1358 -8052
rect -1541 -8124 -1365 -8122
rect -1541 -8131 -1536 -8124
rect -1531 -8145 -1526 -8131
rect -1530 -8146 -1526 -8145
rect -1506 -8146 -1502 -8124
rect -1482 -8146 -1478 -8124
rect -1458 -8146 -1454 -8124
rect -1434 -8146 -1430 -8124
rect -1410 -8146 -1406 -8124
rect -1386 -8146 -1382 -8124
rect -1379 -8125 -1365 -8124
rect -1362 -8145 -1355 -8101
rect -1373 -8146 -1339 -8145
rect -2393 -8148 -1339 -8146
rect -2371 -8170 -2366 -8148
rect -2348 -8170 -2343 -8148
rect -2325 -8170 -2320 -8148
rect -2309 -8166 -2301 -8156
rect -2068 -8165 -2062 -8160
rect -2317 -8170 -2309 -8166
rect -2060 -8170 -2050 -8165
rect -2000 -8170 -1992 -8148
rect -1806 -8156 -1680 -8150
rect -1854 -8165 -1806 -8160
rect -1655 -8166 -1647 -8156
rect -1972 -8170 -1964 -8169
rect -1958 -8170 -1942 -8168
rect -1844 -8170 -1806 -8167
rect -1663 -8170 -1655 -8166
rect -1642 -8170 -1637 -8148
rect -1619 -8170 -1614 -8148
rect -1530 -8170 -1526 -8148
rect -1506 -8170 -1502 -8148
rect -1482 -8170 -1478 -8148
rect -1458 -8170 -1454 -8148
rect -1434 -8170 -1430 -8148
rect -1410 -8170 -1406 -8148
rect -1386 -8169 -1382 -8148
rect -1379 -8149 -1365 -8148
rect -1362 -8149 -1355 -8148
rect -1373 -8155 -1368 -8149
rect -1362 -8155 -1358 -8149
rect -1363 -8169 -1358 -8155
rect -1397 -8170 -1339 -8169
rect -1338 -8170 -1334 -8052
rect -1314 -8074 -1307 -8053
rect -1290 -8074 -1286 -8052
rect -1218 -8074 -1214 -8028
rect -1194 -8074 -1190 -8028
rect -1170 -8073 -1166 -8028
rect -1157 -8035 -1152 -8028
rect -1146 -8035 -1142 -8028
rect -1147 -8049 -1142 -8035
rect -1181 -8074 -1147 -8073
rect -1331 -8076 -1147 -8074
rect -1331 -8077 -1317 -8076
rect -1314 -8077 -1307 -8076
rect -1314 -8170 -1310 -8077
rect -1290 -8170 -1286 -8076
rect -1253 -8098 -1219 -8097
rect -1218 -8098 -1214 -8076
rect -1194 -8097 -1190 -8076
rect -1181 -8083 -1176 -8076
rect -1170 -8083 -1166 -8076
rect -1171 -8097 -1166 -8083
rect -1205 -8098 -1171 -8097
rect -1253 -8100 -1171 -8098
rect -1243 -8112 -1235 -8107
rect -1243 -8120 -1241 -8112
rect -1243 -8121 -1235 -8120
rect -1253 -8122 -1219 -8121
rect -1259 -8124 -1219 -8122
rect -1266 -8169 -1262 -8124
rect -1259 -8125 -1245 -8124
rect -1243 -8138 -1235 -8131
rect -1218 -8134 -1214 -8100
rect -1205 -8107 -1200 -8100
rect -1194 -8107 -1190 -8100
rect -1195 -8121 -1190 -8107
rect -1243 -8144 -1241 -8138
rect -1243 -8145 -1235 -8144
rect -1277 -8170 -1243 -8169
rect -2393 -8172 -1243 -8170
rect -2371 -8194 -2366 -8172
rect -2348 -8194 -2343 -8172
rect -2325 -8194 -2320 -8172
rect -2060 -8178 -2050 -8172
rect -2309 -8194 -2301 -8184
rect -2060 -8185 -2030 -8178
rect -2000 -8182 -1992 -8172
rect -1972 -8174 -1942 -8172
rect -1958 -8175 -1942 -8174
rect -1844 -8176 -1806 -8172
rect -2068 -8192 -2062 -8185
rect -2062 -8194 -2036 -8192
rect -2393 -8196 -2036 -8194
rect -2030 -8194 -2012 -8192
rect -2004 -8194 -1990 -8182
rect -1844 -8183 -1798 -8178
rect -1806 -8185 -1798 -8183
rect -1854 -8187 -1844 -8185
rect -1854 -8192 -1806 -8187
rect -1864 -8194 -1796 -8193
rect -1655 -8194 -1647 -8184
rect -1642 -8194 -1637 -8172
rect -1619 -8194 -1614 -8172
rect -1530 -8194 -1526 -8172
rect -1506 -8173 -1502 -8172
rect -2030 -8196 -1509 -8194
rect -2371 -8613 -2366 -8196
rect -2361 -8593 -2353 -8583
rect -2348 -8593 -2343 -8196
rect -2351 -8609 -2343 -8593
rect -2371 -8639 -2363 -8613
rect -2383 -8811 -2376 -8801
rect -2371 -8811 -2366 -8639
rect -2373 -8822 -2366 -8811
rect -2348 -8822 -2343 -8609
rect -2325 -8327 -2320 -8196
rect -2317 -8200 -2309 -8196
rect -2060 -8200 -2050 -8196
rect -2060 -8202 -2036 -8200
rect -2060 -8204 -2030 -8202
rect -2292 -8210 -2030 -8204
rect -2092 -8226 -2062 -8224
rect -2094 -8230 -2062 -8226
rect -2309 -8260 -2301 -8251
rect -2317 -8267 -2309 -8260
rect -2309 -8288 -2301 -8280
rect -2251 -8286 -2093 -8280
rect -2317 -8296 -2309 -8288
rect -2154 -8293 -2138 -8290
rect -2084 -8293 -2054 -8288
rect -2143 -8306 -2138 -8300
rect -2325 -8337 -2317 -8327
rect -2325 -8356 -2320 -8337
rect -2317 -8343 -2309 -8337
rect -2243 -8354 -2221 -8346
rect -2211 -8354 -2201 -8334
rect -2073 -8354 -2065 -8336
rect -2000 -8354 -1992 -8196
rect -1844 -8203 -1806 -8196
rect -1663 -8200 -1655 -8196
rect -1844 -8210 -1680 -8204
rect -1854 -8226 -1806 -8224
rect -1854 -8230 -1680 -8226
rect -1915 -8260 -1906 -8250
rect -1846 -8252 -1837 -8250
rect -1790 -8252 -1680 -8250
rect -1655 -8260 -1647 -8254
rect -1905 -8269 -1896 -8260
rect -1837 -8261 -1790 -8260
rect -1837 -8276 -1798 -8263
rect -1663 -8270 -1655 -8260
rect -1798 -8286 -1790 -8281
rect -1837 -8288 -1798 -8286
rect -1655 -8288 -1647 -8282
rect -1846 -8290 -1837 -8288
rect -1846 -8293 -1798 -8290
rect -1837 -8306 -1798 -8296
rect -1663 -8298 -1655 -8288
rect -1671 -8338 -1663 -8330
rect -1655 -8338 -1647 -8336
rect -1663 -8346 -1647 -8338
rect -1642 -8346 -1637 -8196
rect -1885 -8354 -1877 -8352
rect -1708 -8354 -1672 -8352
rect -2243 -8355 -2213 -8354
rect -2325 -8365 -2317 -8356
rect -2259 -8361 -2211 -8355
rect -2183 -8361 -1877 -8354
rect -1869 -8361 -1758 -8354
rect -1710 -8360 -1672 -8354
rect -1710 -8361 -1692 -8360
rect -2211 -8365 -2201 -8361
rect -2325 -8385 -2320 -8365
rect -2317 -8372 -2309 -8365
rect -2211 -8372 -2198 -8365
rect -2325 -8393 -2317 -8385
rect -2300 -8392 -2292 -8382
rect -2243 -8391 -2228 -8380
rect -2211 -8388 -2181 -8372
rect -2211 -8391 -2201 -8388
rect -2325 -8413 -2320 -8393
rect -2317 -8401 -2309 -8393
rect -2325 -8421 -2317 -8413
rect -2325 -8441 -2320 -8421
rect -2317 -8429 -2309 -8421
rect -2325 -8450 -2317 -8441
rect -2325 -8469 -2320 -8450
rect -2317 -8457 -2309 -8450
rect -2325 -8478 -2317 -8469
rect -2325 -8498 -2320 -8478
rect -2317 -8485 -2309 -8478
rect -2325 -8506 -2317 -8498
rect -2290 -8505 -2282 -8392
rect -2251 -8402 -2240 -8398
rect -2211 -8402 -2181 -8398
rect -2251 -8405 -2181 -8402
rect -2176 -8412 -2173 -8410
rect -2240 -8419 -2173 -8412
rect -2169 -8417 -2163 -8362
rect -2073 -8398 -2065 -8361
rect -2073 -8402 -2043 -8398
rect -2000 -8402 -1992 -8361
rect -1915 -8392 -1907 -8383
rect -1963 -8398 -1955 -8392
rect -1963 -8402 -1915 -8398
rect -1885 -8402 -1877 -8361
rect -1875 -8366 -1869 -8362
rect -1829 -8384 -1781 -8382
rect -1847 -8388 -1781 -8384
rect -1778 -8388 -1771 -8362
rect -1758 -8369 -1710 -8362
rect -1718 -8376 -1710 -8369
rect -1768 -8386 -1760 -8376
rect -1718 -8378 -1700 -8376
rect -2146 -8405 -2135 -8402
rect -2105 -8405 -2043 -8402
rect -2035 -8405 -1989 -8402
rect -1973 -8405 -1915 -8402
rect -1907 -8405 -1854 -8402
rect -2073 -8407 -2043 -8405
rect -2135 -8419 -2105 -8412
rect -2065 -8414 -2043 -8407
rect -2243 -8430 -2240 -8421
rect -2221 -8427 -2213 -8419
rect -2211 -8427 -2208 -8419
rect -2203 -8426 -2173 -8419
rect -2251 -8437 -2240 -8430
rect -2211 -8430 -2203 -8427
rect -2211 -8437 -2181 -8430
rect -2073 -8437 -2043 -8430
rect -2203 -8460 -2173 -8453
rect -2262 -8478 -2240 -8468
rect -2203 -8469 -2176 -8460
rect -2083 -8471 -2075 -8461
rect -2040 -8471 -2035 -8467
rect -2073 -8483 -2043 -8471
rect -2028 -8483 -2023 -8471
rect -2000 -8478 -1992 -8405
rect -1963 -8408 -1955 -8405
rect -1963 -8409 -1915 -8408
rect -1955 -8419 -1907 -8412
rect -1885 -8416 -1877 -8405
rect -1837 -8410 -1828 -8394
rect -1758 -8401 -1750 -8386
rect -1758 -8402 -1692 -8401
rect -1837 -8412 -1833 -8410
rect -1837 -8414 -1835 -8412
rect -1887 -8419 -1851 -8416
rect -1750 -8419 -1702 -8412
rect -1885 -8424 -1877 -8419
rect -1963 -8437 -1915 -8430
rect -1905 -8469 -1897 -8424
rect -1857 -8442 -1851 -8419
rect -1760 -8427 -1758 -8426
rect -1837 -8437 -1789 -8430
rect -1758 -8436 -1750 -8430
rect -1758 -8437 -1710 -8436
rect -1955 -8472 -1915 -8469
rect -1963 -8478 -1962 -8476
rect -2000 -8481 -1981 -8478
rect -1965 -8481 -1962 -8478
rect -1955 -8478 -1907 -8474
rect -1885 -8478 -1877 -8459
rect -1857 -8472 -1851 -8460
rect -1750 -8464 -1702 -8457
rect -1829 -8472 -1789 -8470
rect -1766 -8474 -1760 -8464
rect -1829 -8478 -1781 -8474
rect -1756 -8478 -1740 -8474
rect -1680 -8478 -1672 -8360
rect -1671 -8366 -1663 -8358
rect -1645 -8362 -1637 -8346
rect -1663 -8374 -1655 -8366
rect -1671 -8394 -1663 -8386
rect -1663 -8402 -1655 -8394
rect -1671 -8422 -1663 -8414
rect -1671 -8438 -1669 -8425
rect -1663 -8430 -1655 -8422
rect -1671 -8450 -1663 -8442
rect -1663 -8458 -1655 -8450
rect -1671 -8478 -1663 -8470
rect -1955 -8481 -1837 -8478
rect -1829 -8481 -1740 -8478
rect -2206 -8491 -2176 -8488
rect -2206 -8494 -2203 -8491
rect -2161 -8493 -2145 -8484
rect -2073 -8486 -2065 -8483
rect -2073 -8487 -2043 -8486
rect -2028 -8487 -2012 -8483
rect -2073 -8494 -2065 -8488
rect -2203 -8495 -2176 -8494
rect -2065 -8495 -2043 -8494
rect -2262 -8501 -2232 -8495
rect -2176 -8501 -2173 -8495
rect -2043 -8501 -2035 -8495
rect -2325 -8526 -2320 -8506
rect -2317 -8514 -2309 -8506
rect -2153 -8507 -2146 -8503
rect -2325 -8534 -2317 -8526
rect -2300 -8530 -2292 -8520
rect -2325 -8554 -2320 -8534
rect -2317 -8542 -2309 -8534
rect -2325 -8562 -2317 -8554
rect -2325 -8582 -2320 -8562
rect -2317 -8570 -2309 -8562
rect -2290 -8563 -2282 -8530
rect -2273 -8534 -2264 -8529
rect -2206 -8534 -2176 -8529
rect -2262 -8541 -2232 -8536
rect -2198 -8545 -2176 -8534
rect -2198 -8559 -2176 -8551
rect -2166 -8567 -2158 -8519
rect -2143 -8523 -2136 -8507
rect -2143 -8534 -2113 -8529
rect -2073 -8534 -2065 -8529
rect -2065 -8536 -2043 -8534
rect -2043 -8541 -2035 -8536
rect -2065 -8562 -2043 -8547
rect -2006 -8563 -2004 -8547
rect -2265 -8577 -2260 -8571
rect -2143 -8577 -2113 -8570
rect -2270 -8578 -2240 -8577
rect -2270 -8581 -2265 -8578
rect -2325 -8590 -2317 -8582
rect -2325 -8610 -2320 -8590
rect -2317 -8598 -2309 -8590
rect -2113 -8593 -2105 -8583
rect -2291 -8605 -2270 -8598
rect -2198 -8600 -2168 -8598
rect -2135 -8599 -2105 -8598
rect -2103 -8599 -2095 -8593
rect -2113 -8600 -2105 -8599
rect -2065 -8600 -2035 -8598
rect -2000 -8600 -1992 -8481
rect -1963 -8488 -1960 -8481
rect -1915 -8485 -1905 -8481
rect -1963 -8489 -1955 -8488
rect -1963 -8495 -1915 -8489
rect -1989 -8522 -1973 -8519
rect -1915 -8522 -1907 -8515
rect -1990 -8557 -1989 -8536
rect -1983 -8600 -1981 -8537
rect -1885 -8546 -1877 -8481
rect -1789 -8486 -1778 -8481
rect -1837 -8489 -1829 -8488
rect -1837 -8495 -1789 -8489
rect -1756 -8490 -1740 -8481
rect -1837 -8505 -1829 -8495
rect -1872 -8524 -1867 -8514
rect -1789 -8522 -1781 -8515
rect -1776 -8522 -1769 -8505
rect -1756 -8512 -1750 -8490
rect -1671 -8494 -1669 -8483
rect -1663 -8486 -1655 -8478
rect -1671 -8506 -1663 -8498
rect -1663 -8514 -1655 -8506
rect -1702 -8524 -1696 -8518
rect -1955 -8548 -1915 -8546
rect -1963 -8550 -1955 -8548
rect -1963 -8557 -1915 -8550
rect -1963 -8565 -1955 -8557
rect -1963 -8566 -1915 -8565
rect -1973 -8572 -1965 -8569
rect -1955 -8572 -1907 -8568
rect -1974 -8575 -1907 -8572
rect -1973 -8579 -1965 -8575
rect -1963 -8579 -1960 -8577
rect -1963 -8583 -1915 -8579
rect -1963 -8591 -1955 -8583
rect -1963 -8595 -1915 -8591
rect -1963 -8598 -1955 -8595
rect -2240 -8605 -2206 -8600
rect -2198 -8605 -2143 -8600
rect -2113 -8605 -1981 -8600
rect -1915 -8605 -1907 -8598
rect -2270 -8610 -2266 -8606
rect -2086 -8609 -2070 -8605
rect -2325 -8618 -2317 -8610
rect -2270 -8617 -2240 -8610
rect -2206 -8617 -2176 -8610
rect -2325 -8638 -2320 -8618
rect -2317 -8626 -2309 -8618
rect -2270 -8622 -2266 -8617
rect -2270 -8626 -2266 -8623
rect -2198 -8626 -2176 -8619
rect -2166 -8626 -2158 -8609
rect -2143 -8617 -2113 -8610
rect -2198 -8635 -2168 -8631
rect -2325 -8646 -2317 -8638
rect -2143 -8640 -2136 -8626
rect -2085 -8631 -2060 -8630
rect -2039 -8631 -2035 -8622
rect -2135 -8638 -2105 -8631
rect -2085 -8638 -2035 -8631
rect -2029 -8638 -2025 -8631
rect -2325 -8659 -2320 -8646
rect -2317 -8654 -2309 -8646
rect -2235 -8656 -2232 -8653
rect -2325 -8685 -2317 -8659
rect -2325 -8694 -2320 -8685
rect -2325 -8702 -2317 -8694
rect -2135 -8702 -2119 -8689
rect -2000 -8697 -1992 -8605
rect -1983 -8623 -1981 -8605
rect -1955 -8623 -1915 -8622
rect -1862 -8626 -1857 -8524
rect -1706 -8528 -1702 -8524
rect -1829 -8540 -1789 -8532
rect -1671 -8534 -1663 -8526
rect -1849 -8548 -1842 -8540
rect -1790 -8548 -1781 -8540
rect -1663 -8542 -1655 -8534
rect -1837 -8557 -1829 -8550
rect -1758 -8557 -1732 -8550
rect -1748 -8566 -1732 -8557
rect -1671 -8562 -1663 -8554
rect -1829 -8575 -1781 -8568
rect -1663 -8570 -1655 -8562
rect -1829 -8581 -1789 -8577
rect -1768 -8580 -1760 -8570
rect -1758 -8581 -1750 -8580
rect -1671 -8590 -1663 -8582
rect -1837 -8593 -1780 -8590
rect -1758 -8596 -1748 -8590
rect -1708 -8596 -1690 -8590
rect -1829 -8605 -1781 -8598
rect -1680 -8607 -1672 -8590
rect -1663 -8598 -1655 -8590
rect -1829 -8616 -1791 -8610
rect -1758 -8616 -1710 -8614
rect -1758 -8623 -1692 -8616
rect -1671 -8618 -1663 -8610
rect -1955 -8634 -1907 -8631
rect -1791 -8634 -1781 -8631
rect -1991 -8638 -1839 -8634
rect -1791 -8638 -1780 -8634
rect -1680 -8641 -1672 -8623
rect -1663 -8626 -1655 -8618
rect -1839 -8651 -1791 -8644
rect -1671 -8646 -1663 -8638
rect -1829 -8657 -1791 -8653
rect -1671 -8656 -1669 -8646
rect -1663 -8654 -1655 -8646
rect -1680 -8672 -1672 -8657
rect -1642 -8672 -1637 -8362
rect -1619 -8412 -1614 -8196
rect -1541 -8347 -1536 -8337
rect -1530 -8347 -1526 -8196
rect -1523 -8197 -1509 -8196
rect -1531 -8361 -1526 -8347
rect -1506 -8221 -1499 -8173
rect -1541 -8371 -1536 -8361
rect -1531 -8385 -1526 -8371
rect -1619 -8438 -1611 -8412
rect -1768 -8688 -1760 -8678
rect -1758 -8695 -1710 -8688
rect -2325 -8722 -2320 -8702
rect -2317 -8710 -2306 -8702
rect -2031 -8705 -1992 -8697
rect -1750 -8699 -1710 -8695
rect -1674 -8700 -1663 -8694
rect -2307 -8718 -2306 -8710
rect -2149 -8707 -2135 -8706
rect -2149 -8711 -2119 -8707
rect -2024 -8716 -2021 -8707
rect -2325 -8730 -2317 -8722
rect -2325 -8778 -2320 -8730
rect -2317 -8738 -2306 -8730
rect -2185 -8732 -2169 -8720
rect -2056 -8723 -2040 -8719
rect -2021 -8723 -2008 -8716
rect -2056 -8734 -2054 -8724
rect -2056 -8735 -2048 -8734
rect -2307 -8774 -2306 -8766
rect -2111 -8767 -2054 -8761
rect -2325 -8786 -2314 -8778
rect -2104 -8785 -2101 -8781
rect -2325 -8806 -2320 -8786
rect -2314 -8794 -2306 -8786
rect -2104 -8788 -2101 -8786
rect -2084 -8788 -2054 -8787
rect -2000 -8788 -1992 -8705
rect -1758 -8706 -1750 -8705
rect -1758 -8707 -1749 -8706
rect -1758 -8708 -1710 -8707
rect -1663 -8710 -1658 -8700
rect -1831 -8718 -1783 -8714
rect -1784 -8731 -1783 -8718
rect -1674 -8728 -1663 -8722
rect -1826 -8733 -1796 -8732
rect -1663 -8738 -1658 -8728
rect -1654 -8732 -1647 -8722
rect -1644 -8746 -1637 -8732
rect -1758 -8764 -1750 -8761
rect -1758 -8767 -1710 -8764
rect -1844 -8779 -1828 -8777
rect -1844 -8780 -1792 -8779
rect -1828 -8781 -1792 -8780
rect -1772 -8781 -1758 -8773
rect -1750 -8776 -1702 -8769
rect -1750 -8784 -1710 -8780
rect -1700 -8784 -1692 -8764
rect -1674 -8772 -1665 -8764
rect -1674 -8784 -1666 -8776
rect -1758 -8788 -1710 -8787
rect -2307 -8802 -2306 -8794
rect -2139 -8798 -2123 -8789
rect -2111 -8794 -2016 -8788
rect -2139 -8805 -2111 -8798
rect -2325 -8814 -2314 -8806
rect -2177 -8812 -2161 -8811
rect -2141 -8812 -2119 -8810
rect -2104 -8812 -2101 -8794
rect -2076 -8805 -2046 -8800
rect -2325 -8822 -2320 -8814
rect -2314 -8822 -2306 -8814
rect -2076 -8816 -2054 -8810
rect -2021 -8813 -2016 -8794
rect -2000 -8794 -1818 -8788
rect -1802 -8794 -1776 -8788
rect -1760 -8794 -1710 -8788
rect -1666 -8792 -1658 -8784
rect -2189 -8822 -2175 -8817
rect -2373 -8824 -2175 -8822
rect -2373 -8825 -2359 -8824
rect -2371 -9237 -2366 -8825
rect -2348 -8877 -2343 -8824
rect -2325 -8834 -2320 -8824
rect -2307 -8830 -2306 -8824
rect -2189 -8825 -2175 -8824
rect -2149 -8826 -2119 -8817
rect -2084 -8818 -2036 -8817
rect -2000 -8818 -1992 -8794
rect -1758 -8796 -1710 -8794
rect -1758 -8798 -1755 -8796
rect -1828 -8805 -1792 -8798
rect -1768 -8807 -1760 -8800
rect -1758 -8805 -1757 -8798
rect -1710 -8799 -1702 -8798
rect -1750 -8805 -1702 -8799
rect -1674 -8800 -1665 -8792
rect -1768 -8810 -1764 -8807
rect -1758 -8810 -1755 -8805
rect -1818 -8818 -1789 -8810
rect -1758 -8817 -1754 -8810
rect -1750 -8815 -1710 -8810
rect -1674 -8812 -1666 -8804
rect -1758 -8818 -1692 -8817
rect -2084 -8820 -1692 -8818
rect -1666 -8820 -1658 -8812
rect -2084 -8823 -1690 -8820
rect -2084 -8826 -2054 -8823
rect -2046 -8825 -1710 -8823
rect -2325 -8842 -2314 -8834
rect -2076 -8835 -2046 -8828
rect -2325 -8862 -2320 -8842
rect -2314 -8850 -2306 -8842
rect -2076 -8843 -2054 -8837
rect -2084 -8847 -2054 -8845
rect -2104 -8850 -2054 -8847
rect -2307 -8858 -2306 -8850
rect -2084 -8853 -2054 -8850
rect -2325 -8874 -2314 -8862
rect -2348 -8901 -2341 -8877
rect -2325 -8891 -2320 -8874
rect -2314 -8878 -2309 -8874
rect -2309 -8890 -2298 -8878
rect -2314 -8891 -2309 -8890
rect -2361 -9217 -2353 -9207
rect -2348 -9217 -2343 -8901
rect -2351 -9233 -2343 -9217
rect -2371 -9263 -2363 -9237
rect -2383 -9435 -2376 -9425
rect -2371 -9435 -2366 -9263
rect -2373 -9446 -2366 -9435
rect -2348 -9446 -2343 -9233
rect -2325 -8903 -2314 -8891
rect -2076 -8902 -2073 -8886
rect -2325 -8920 -2320 -8903
rect -2314 -8906 -2309 -8903
rect -2309 -8918 -2298 -8906
rect -2251 -8910 -2101 -8903
rect -2141 -8917 -2111 -8911
rect -2086 -8913 -2083 -8903
rect -2076 -8917 -2046 -8911
rect -2314 -8920 -2309 -8918
rect -2325 -8932 -2314 -8920
rect -2141 -8929 -2113 -8924
rect -2076 -8929 -2073 -8926
rect -2325 -8951 -2320 -8932
rect -2314 -8934 -2309 -8932
rect -2325 -8961 -2317 -8951
rect -2325 -8980 -2320 -8961
rect -2317 -8967 -2309 -8961
rect -2243 -8978 -2221 -8970
rect -2211 -8978 -2201 -8958
rect -2073 -8978 -2065 -8960
rect -2000 -8978 -1992 -8825
rect -1758 -8826 -1710 -8825
rect -1680 -8828 -1665 -8820
rect -1750 -8835 -1702 -8828
rect -1680 -8832 -1672 -8828
rect -1680 -8837 -1666 -8832
rect -1836 -8841 -1820 -8840
rect -1837 -8845 -1820 -8841
rect -1750 -8843 -1710 -8837
rect -1674 -8840 -1666 -8837
rect -1837 -8852 -1789 -8845
rect -1758 -8846 -1710 -8845
rect -1760 -8849 -1692 -8846
rect -1666 -8848 -1658 -8840
rect -1837 -8853 -1820 -8852
rect -1764 -8853 -1692 -8849
rect -1674 -8853 -1665 -8848
rect -1680 -8856 -1665 -8853
rect -1680 -8884 -1672 -8856
rect -1666 -8876 -1665 -8866
rect -1837 -8886 -1789 -8884
rect -1829 -8900 -1789 -8886
rect -1655 -8888 -1650 -8878
rect -1666 -8894 -1655 -8888
rect -1778 -8902 -1771 -8900
rect -1710 -8902 -1702 -8900
rect -1666 -8904 -1665 -8894
rect -1837 -8910 -1829 -8904
rect -1829 -8911 -1789 -8910
rect -1726 -8911 -1710 -8910
rect -1789 -8913 -1781 -8911
rect -1829 -8917 -1781 -8913
rect -1750 -8917 -1710 -8911
rect -1829 -8929 -1789 -8920
rect -1726 -8926 -1710 -8917
rect -1706 -8926 -1702 -8913
rect -1655 -8916 -1650 -8906
rect -1666 -8922 -1655 -8916
rect -1666 -8932 -1665 -8922
rect -1671 -8962 -1663 -8954
rect -1655 -8962 -1647 -8960
rect -1663 -8970 -1647 -8962
rect -1642 -8970 -1637 -8746
rect -1619 -8748 -1614 -8438
rect -1885 -8978 -1877 -8976
rect -1708 -8978 -1672 -8976
rect -2243 -8979 -2213 -8978
rect -2325 -8989 -2317 -8980
rect -2259 -8985 -2211 -8979
rect -2183 -8985 -1877 -8978
rect -1869 -8985 -1758 -8978
rect -1710 -8984 -1672 -8978
rect -1710 -8985 -1692 -8984
rect -2211 -8989 -2201 -8985
rect -2325 -9009 -2320 -8989
rect -2317 -8996 -2309 -8989
rect -2211 -8996 -2198 -8989
rect -2325 -9017 -2317 -9009
rect -2300 -9016 -2292 -9006
rect -2243 -9015 -2228 -9004
rect -2211 -9012 -2181 -8996
rect -2211 -9015 -2201 -9012
rect -2325 -9037 -2320 -9017
rect -2317 -9025 -2309 -9017
rect -2325 -9045 -2317 -9037
rect -2325 -9065 -2320 -9045
rect -2317 -9053 -2309 -9045
rect -2325 -9074 -2317 -9065
rect -2325 -9093 -2320 -9074
rect -2317 -9081 -2309 -9074
rect -2325 -9102 -2317 -9093
rect -2325 -9122 -2320 -9102
rect -2317 -9109 -2309 -9102
rect -2325 -9130 -2317 -9122
rect -2290 -9129 -2282 -9016
rect -2251 -9026 -2240 -9022
rect -2211 -9026 -2181 -9022
rect -2251 -9029 -2181 -9026
rect -2176 -9036 -2173 -9034
rect -2240 -9043 -2173 -9036
rect -2169 -9041 -2163 -8986
rect -2073 -9022 -2065 -8985
rect -2073 -9026 -2043 -9022
rect -2000 -9026 -1992 -8985
rect -1915 -9016 -1907 -9007
rect -1963 -9022 -1955 -9016
rect -1963 -9026 -1915 -9022
rect -1885 -9026 -1877 -8985
rect -1875 -8990 -1869 -8986
rect -1829 -9008 -1781 -9006
rect -1847 -9012 -1781 -9008
rect -1778 -9012 -1771 -8986
rect -1758 -8993 -1710 -8986
rect -1718 -9000 -1710 -8993
rect -1768 -9010 -1760 -9000
rect -1718 -9002 -1700 -9000
rect -2146 -9029 -2135 -9026
rect -2105 -9029 -2043 -9026
rect -2035 -9029 -1989 -9026
rect -1973 -9029 -1915 -9026
rect -1907 -9029 -1854 -9026
rect -2073 -9031 -2043 -9029
rect -2135 -9043 -2105 -9036
rect -2065 -9038 -2043 -9031
rect -2243 -9054 -2240 -9045
rect -2221 -9051 -2213 -9043
rect -2211 -9051 -2208 -9043
rect -2203 -9050 -2173 -9043
rect -2251 -9061 -2240 -9054
rect -2211 -9054 -2203 -9051
rect -2211 -9061 -2181 -9054
rect -2073 -9061 -2043 -9054
rect -2203 -9084 -2173 -9077
rect -2262 -9102 -2240 -9092
rect -2203 -9093 -2176 -9084
rect -2083 -9095 -2075 -9085
rect -2040 -9095 -2035 -9091
rect -2073 -9107 -2043 -9095
rect -2028 -9107 -2023 -9095
rect -2000 -9102 -1992 -9029
rect -1963 -9032 -1955 -9029
rect -1963 -9033 -1915 -9032
rect -1955 -9043 -1907 -9036
rect -1885 -9040 -1877 -9029
rect -1837 -9034 -1828 -9018
rect -1758 -9025 -1750 -9010
rect -1758 -9026 -1692 -9025
rect -1837 -9036 -1833 -9034
rect -1837 -9038 -1835 -9036
rect -1887 -9043 -1851 -9040
rect -1750 -9043 -1702 -9036
rect -1885 -9048 -1877 -9043
rect -1963 -9061 -1915 -9054
rect -1905 -9093 -1897 -9048
rect -1857 -9066 -1851 -9043
rect -1760 -9051 -1758 -9050
rect -1837 -9061 -1789 -9054
rect -1758 -9060 -1750 -9054
rect -1758 -9061 -1710 -9060
rect -1955 -9096 -1915 -9093
rect -1963 -9102 -1962 -9100
rect -2000 -9105 -1981 -9102
rect -1965 -9105 -1962 -9102
rect -1955 -9102 -1907 -9098
rect -1885 -9102 -1877 -9083
rect -1857 -9096 -1851 -9084
rect -1750 -9088 -1702 -9081
rect -1829 -9096 -1789 -9094
rect -1766 -9098 -1760 -9088
rect -1829 -9102 -1781 -9098
rect -1756 -9102 -1740 -9098
rect -1680 -9102 -1672 -8984
rect -1671 -8990 -1663 -8982
rect -1645 -8986 -1637 -8970
rect -1663 -8998 -1655 -8990
rect -1671 -9018 -1663 -9010
rect -1663 -9026 -1655 -9018
rect -1671 -9046 -1663 -9038
rect -1671 -9062 -1669 -9049
rect -1663 -9054 -1655 -9046
rect -1671 -9074 -1663 -9066
rect -1663 -9082 -1655 -9074
rect -1671 -9102 -1663 -9094
rect -1955 -9105 -1837 -9102
rect -1829 -9105 -1740 -9102
rect -2206 -9115 -2176 -9112
rect -2206 -9118 -2203 -9115
rect -2161 -9117 -2145 -9108
rect -2073 -9110 -2065 -9107
rect -2073 -9111 -2043 -9110
rect -2028 -9111 -2012 -9107
rect -2073 -9118 -2065 -9112
rect -2203 -9119 -2176 -9118
rect -2065 -9119 -2043 -9118
rect -2262 -9125 -2232 -9119
rect -2176 -9125 -2173 -9119
rect -2043 -9125 -2035 -9119
rect -2325 -9150 -2320 -9130
rect -2317 -9138 -2309 -9130
rect -2153 -9131 -2146 -9127
rect -2325 -9158 -2317 -9150
rect -2300 -9154 -2292 -9144
rect -2325 -9178 -2320 -9158
rect -2317 -9166 -2309 -9158
rect -2325 -9186 -2317 -9178
rect -2325 -9206 -2320 -9186
rect -2317 -9194 -2309 -9186
rect -2290 -9187 -2282 -9154
rect -2273 -9158 -2264 -9153
rect -2206 -9158 -2176 -9153
rect -2262 -9165 -2232 -9160
rect -2198 -9169 -2176 -9158
rect -2198 -9183 -2176 -9175
rect -2166 -9191 -2158 -9143
rect -2143 -9147 -2136 -9131
rect -2143 -9158 -2113 -9153
rect -2073 -9158 -2065 -9153
rect -2065 -9160 -2043 -9158
rect -2043 -9165 -2035 -9160
rect -2065 -9186 -2043 -9171
rect -2006 -9187 -2004 -9171
rect -2265 -9201 -2260 -9195
rect -2143 -9201 -2113 -9194
rect -2270 -9202 -2240 -9201
rect -2270 -9205 -2265 -9202
rect -2325 -9214 -2317 -9206
rect -2325 -9234 -2320 -9214
rect -2317 -9222 -2309 -9214
rect -2113 -9217 -2105 -9207
rect -2291 -9229 -2270 -9222
rect -2198 -9224 -2168 -9222
rect -2135 -9223 -2105 -9222
rect -2103 -9223 -2095 -9217
rect -2113 -9224 -2105 -9223
rect -2065 -9224 -2035 -9222
rect -2000 -9224 -1992 -9105
rect -1963 -9112 -1960 -9105
rect -1915 -9109 -1905 -9105
rect -1963 -9113 -1955 -9112
rect -1963 -9119 -1915 -9113
rect -1989 -9146 -1973 -9143
rect -1915 -9146 -1907 -9139
rect -1990 -9181 -1989 -9160
rect -1983 -9224 -1981 -9161
rect -1885 -9170 -1877 -9105
rect -1789 -9110 -1778 -9105
rect -1837 -9113 -1829 -9112
rect -1837 -9119 -1789 -9113
rect -1756 -9114 -1740 -9105
rect -1837 -9129 -1829 -9119
rect -1872 -9148 -1867 -9138
rect -1789 -9146 -1781 -9139
rect -1776 -9146 -1769 -9129
rect -1756 -9136 -1750 -9114
rect -1671 -9118 -1669 -9107
rect -1663 -9110 -1655 -9102
rect -1671 -9130 -1663 -9122
rect -1663 -9138 -1655 -9130
rect -1702 -9148 -1696 -9142
rect -1955 -9172 -1915 -9170
rect -1963 -9174 -1955 -9172
rect -1963 -9181 -1915 -9174
rect -1963 -9189 -1955 -9181
rect -1963 -9190 -1915 -9189
rect -1973 -9196 -1965 -9193
rect -1955 -9196 -1907 -9192
rect -1974 -9199 -1907 -9196
rect -1973 -9203 -1965 -9199
rect -1963 -9203 -1960 -9201
rect -1963 -9207 -1915 -9203
rect -1963 -9215 -1955 -9207
rect -1963 -9219 -1915 -9215
rect -1963 -9222 -1955 -9219
rect -2240 -9229 -2206 -9224
rect -2198 -9229 -2143 -9224
rect -2113 -9229 -1981 -9224
rect -1915 -9229 -1907 -9222
rect -2270 -9234 -2266 -9230
rect -2086 -9233 -2070 -9229
rect -2325 -9242 -2317 -9234
rect -2270 -9241 -2240 -9234
rect -2206 -9241 -2176 -9234
rect -2325 -9262 -2320 -9242
rect -2317 -9250 -2309 -9242
rect -2270 -9246 -2266 -9241
rect -2270 -9250 -2266 -9247
rect -2198 -9250 -2176 -9243
rect -2166 -9250 -2158 -9233
rect -2143 -9241 -2113 -9234
rect -2198 -9259 -2168 -9255
rect -2325 -9270 -2317 -9262
rect -2143 -9264 -2136 -9250
rect -2085 -9255 -2060 -9254
rect -2039 -9255 -2035 -9246
rect -2135 -9262 -2105 -9255
rect -2085 -9262 -2035 -9255
rect -2029 -9262 -2025 -9255
rect -2325 -9283 -2320 -9270
rect -2317 -9278 -2309 -9270
rect -2235 -9280 -2232 -9277
rect -2325 -9309 -2317 -9283
rect -2325 -9318 -2320 -9309
rect -2325 -9326 -2317 -9318
rect -2135 -9326 -2119 -9313
rect -2000 -9321 -1992 -9229
rect -1983 -9247 -1981 -9229
rect -1955 -9247 -1915 -9246
rect -1862 -9250 -1857 -9148
rect -1706 -9152 -1702 -9148
rect -1829 -9164 -1789 -9156
rect -1671 -9158 -1663 -9150
rect -1849 -9172 -1842 -9164
rect -1790 -9172 -1781 -9164
rect -1663 -9166 -1655 -9158
rect -1837 -9181 -1829 -9174
rect -1758 -9181 -1732 -9174
rect -1748 -9190 -1732 -9181
rect -1671 -9186 -1663 -9178
rect -1829 -9199 -1781 -9192
rect -1663 -9194 -1655 -9186
rect -1829 -9205 -1789 -9201
rect -1768 -9204 -1760 -9194
rect -1758 -9205 -1750 -9204
rect -1671 -9214 -1663 -9206
rect -1837 -9217 -1780 -9214
rect -1758 -9220 -1748 -9214
rect -1708 -9220 -1690 -9214
rect -1829 -9229 -1781 -9222
rect -1680 -9231 -1672 -9214
rect -1663 -9222 -1655 -9214
rect -1829 -9240 -1791 -9234
rect -1758 -9240 -1710 -9238
rect -1758 -9247 -1692 -9240
rect -1671 -9242 -1663 -9234
rect -1955 -9258 -1907 -9255
rect -1791 -9258 -1781 -9255
rect -1991 -9262 -1839 -9258
rect -1791 -9262 -1780 -9258
rect -1680 -9265 -1672 -9247
rect -1663 -9250 -1655 -9242
rect -1839 -9275 -1791 -9268
rect -1671 -9270 -1663 -9262
rect -1829 -9281 -1791 -9277
rect -1671 -9280 -1669 -9270
rect -1663 -9278 -1655 -9270
rect -1680 -9296 -1672 -9281
rect -1642 -9296 -1637 -8986
rect -1619 -8822 -1612 -8798
rect -1619 -9036 -1614 -8822
rect -1619 -9062 -1611 -9036
rect -1768 -9312 -1760 -9302
rect -1758 -9319 -1710 -9312
rect -2325 -9346 -2320 -9326
rect -2317 -9334 -2306 -9326
rect -2031 -9329 -1992 -9321
rect -1750 -9323 -1710 -9319
rect -1674 -9324 -1663 -9318
rect -2307 -9342 -2306 -9334
rect -2149 -9331 -2135 -9330
rect -2149 -9335 -2119 -9331
rect -2024 -9340 -2021 -9331
rect -2325 -9354 -2317 -9346
rect -2325 -9402 -2320 -9354
rect -2317 -9362 -2306 -9354
rect -2185 -9356 -2169 -9344
rect -2056 -9347 -2040 -9343
rect -2021 -9347 -2008 -9340
rect -2056 -9358 -2054 -9348
rect -2056 -9359 -2048 -9358
rect -2307 -9398 -2306 -9390
rect -2111 -9391 -2054 -9385
rect -2325 -9410 -2314 -9402
rect -2104 -9409 -2101 -9405
rect -2325 -9430 -2320 -9410
rect -2314 -9418 -2306 -9410
rect -2104 -9412 -2101 -9410
rect -2084 -9412 -2054 -9411
rect -2000 -9412 -1992 -9329
rect -1758 -9330 -1750 -9329
rect -1758 -9331 -1749 -9330
rect -1758 -9332 -1710 -9331
rect -1663 -9334 -1658 -9324
rect -1831 -9342 -1783 -9338
rect -1784 -9355 -1783 -9342
rect -1674 -9352 -1663 -9346
rect -1826 -9357 -1796 -9356
rect -1663 -9362 -1658 -9352
rect -1654 -9356 -1647 -9346
rect -1644 -9370 -1637 -9356
rect -1758 -9388 -1750 -9385
rect -1758 -9391 -1710 -9388
rect -1844 -9403 -1828 -9401
rect -1844 -9404 -1792 -9403
rect -1828 -9405 -1792 -9404
rect -1772 -9405 -1758 -9397
rect -1750 -9400 -1702 -9393
rect -1750 -9408 -1710 -9404
rect -1700 -9408 -1692 -9388
rect -1674 -9396 -1665 -9388
rect -1674 -9408 -1666 -9400
rect -1758 -9412 -1710 -9411
rect -2307 -9426 -2306 -9418
rect -2139 -9422 -2123 -9413
rect -2111 -9418 -2016 -9412
rect -2139 -9429 -2111 -9422
rect -2325 -9438 -2314 -9430
rect -2177 -9436 -2161 -9435
rect -2141 -9436 -2119 -9434
rect -2104 -9436 -2101 -9418
rect -2076 -9429 -2046 -9424
rect -2325 -9446 -2320 -9438
rect -2314 -9446 -2306 -9438
rect -2076 -9440 -2054 -9434
rect -2021 -9437 -2016 -9418
rect -2000 -9418 -1818 -9412
rect -1802 -9418 -1776 -9412
rect -1760 -9418 -1710 -9412
rect -1666 -9416 -1658 -9408
rect -2189 -9446 -2175 -9441
rect -2373 -9448 -2175 -9446
rect -2373 -9449 -2359 -9448
rect -2371 -9861 -2366 -9449
rect -2348 -9501 -2343 -9448
rect -2325 -9458 -2320 -9448
rect -2307 -9454 -2306 -9448
rect -2189 -9449 -2175 -9448
rect -2149 -9450 -2119 -9441
rect -2084 -9442 -2036 -9441
rect -2000 -9442 -1992 -9418
rect -1758 -9420 -1710 -9418
rect -1758 -9422 -1755 -9420
rect -1828 -9429 -1792 -9422
rect -1768 -9431 -1760 -9424
rect -1758 -9429 -1757 -9422
rect -1710 -9423 -1702 -9422
rect -1750 -9429 -1702 -9423
rect -1674 -9424 -1665 -9416
rect -1768 -9434 -1764 -9431
rect -1758 -9434 -1755 -9429
rect -1818 -9442 -1789 -9434
rect -1758 -9441 -1754 -9434
rect -1750 -9439 -1710 -9434
rect -1674 -9436 -1666 -9428
rect -1758 -9442 -1692 -9441
rect -2084 -9444 -1692 -9442
rect -1666 -9444 -1658 -9436
rect -2084 -9447 -1690 -9444
rect -2084 -9450 -2054 -9447
rect -2046 -9449 -1710 -9447
rect -2325 -9466 -2314 -9458
rect -2076 -9459 -2046 -9452
rect -2325 -9486 -2320 -9466
rect -2314 -9474 -2306 -9466
rect -2076 -9467 -2054 -9461
rect -2084 -9471 -2054 -9469
rect -2104 -9474 -2054 -9471
rect -2307 -9482 -2306 -9474
rect -2084 -9477 -2054 -9474
rect -2325 -9498 -2314 -9486
rect -2348 -9525 -2341 -9501
rect -2325 -9515 -2320 -9498
rect -2314 -9502 -2309 -9498
rect -2309 -9514 -2298 -9502
rect -2314 -9515 -2309 -9514
rect -2361 -9841 -2353 -9831
rect -2348 -9841 -2343 -9525
rect -2351 -9857 -2343 -9841
rect -2371 -9887 -2363 -9861
rect -2383 -10059 -2376 -10049
rect -2371 -10059 -2366 -9887
rect -2373 -10070 -2366 -10059
rect -2348 -10070 -2343 -9857
rect -2325 -9527 -2314 -9515
rect -2076 -9526 -2073 -9510
rect -2325 -9544 -2320 -9527
rect -2314 -9530 -2309 -9527
rect -2309 -9542 -2298 -9530
rect -2251 -9534 -2101 -9527
rect -2141 -9541 -2111 -9535
rect -2086 -9537 -2083 -9527
rect -2076 -9541 -2046 -9535
rect -2314 -9544 -2309 -9542
rect -2325 -9556 -2314 -9544
rect -2141 -9553 -2113 -9548
rect -2076 -9553 -2073 -9550
rect -2325 -9575 -2320 -9556
rect -2314 -9558 -2309 -9556
rect -2325 -9585 -2317 -9575
rect -2325 -9604 -2320 -9585
rect -2317 -9591 -2309 -9585
rect -2243 -9602 -2221 -9594
rect -2211 -9602 -2201 -9582
rect -2073 -9602 -2065 -9584
rect -2000 -9602 -1992 -9449
rect -1758 -9450 -1710 -9449
rect -1680 -9452 -1665 -9444
rect -1750 -9459 -1702 -9452
rect -1680 -9456 -1672 -9452
rect -1680 -9461 -1666 -9456
rect -1836 -9465 -1820 -9464
rect -1837 -9469 -1820 -9465
rect -1750 -9467 -1710 -9461
rect -1674 -9464 -1666 -9461
rect -1837 -9476 -1789 -9469
rect -1758 -9470 -1710 -9469
rect -1760 -9473 -1692 -9470
rect -1666 -9472 -1658 -9464
rect -1837 -9477 -1820 -9476
rect -1764 -9477 -1692 -9473
rect -1674 -9477 -1665 -9472
rect -1680 -9480 -1665 -9477
rect -1680 -9508 -1672 -9480
rect -1666 -9500 -1665 -9490
rect -1837 -9510 -1789 -9508
rect -1829 -9524 -1789 -9510
rect -1655 -9512 -1650 -9502
rect -1666 -9518 -1655 -9512
rect -1778 -9526 -1771 -9524
rect -1710 -9526 -1702 -9524
rect -1666 -9528 -1665 -9518
rect -1837 -9534 -1829 -9528
rect -1829 -9535 -1789 -9534
rect -1726 -9535 -1710 -9534
rect -1789 -9537 -1781 -9535
rect -1829 -9541 -1781 -9537
rect -1750 -9541 -1710 -9535
rect -1829 -9553 -1789 -9544
rect -1726 -9550 -1710 -9541
rect -1706 -9550 -1702 -9537
rect -1655 -9540 -1650 -9530
rect -1666 -9546 -1655 -9540
rect -1666 -9556 -1665 -9546
rect -1671 -9586 -1663 -9578
rect -1655 -9586 -1647 -9584
rect -1663 -9594 -1647 -9586
rect -1642 -9594 -1637 -9370
rect -1619 -9372 -1614 -9062
rect -1885 -9602 -1877 -9600
rect -1708 -9602 -1672 -9600
rect -2243 -9603 -2213 -9602
rect -2325 -9613 -2317 -9604
rect -2259 -9609 -2211 -9603
rect -2183 -9609 -1877 -9602
rect -1869 -9609 -1758 -9602
rect -1710 -9608 -1672 -9602
rect -1710 -9609 -1692 -9608
rect -2211 -9613 -2201 -9609
rect -2325 -9633 -2320 -9613
rect -2317 -9620 -2309 -9613
rect -2211 -9620 -2198 -9613
rect -2325 -9641 -2317 -9633
rect -2300 -9640 -2292 -9630
rect -2243 -9639 -2228 -9628
rect -2211 -9636 -2181 -9620
rect -2211 -9639 -2201 -9636
rect -2325 -9661 -2320 -9641
rect -2317 -9649 -2309 -9641
rect -2325 -9669 -2317 -9661
rect -2325 -9689 -2320 -9669
rect -2317 -9677 -2309 -9669
rect -2325 -9698 -2317 -9689
rect -2325 -9717 -2320 -9698
rect -2317 -9705 -2309 -9698
rect -2325 -9726 -2317 -9717
rect -2325 -9746 -2320 -9726
rect -2317 -9733 -2309 -9726
rect -2325 -9754 -2317 -9746
rect -2290 -9753 -2282 -9640
rect -2251 -9650 -2240 -9646
rect -2211 -9650 -2181 -9646
rect -2251 -9653 -2181 -9650
rect -2176 -9660 -2173 -9658
rect -2240 -9667 -2173 -9660
rect -2169 -9665 -2163 -9610
rect -2073 -9646 -2065 -9609
rect -2073 -9650 -2043 -9646
rect -2000 -9650 -1992 -9609
rect -1915 -9640 -1907 -9631
rect -1963 -9646 -1955 -9640
rect -1963 -9650 -1915 -9646
rect -1885 -9650 -1877 -9609
rect -1875 -9614 -1869 -9610
rect -1829 -9632 -1781 -9630
rect -1847 -9636 -1781 -9632
rect -1778 -9636 -1771 -9610
rect -1758 -9617 -1710 -9610
rect -1718 -9624 -1710 -9617
rect -1768 -9634 -1760 -9624
rect -1718 -9626 -1700 -9624
rect -2146 -9653 -2135 -9650
rect -2105 -9653 -2043 -9650
rect -2035 -9653 -1989 -9650
rect -1973 -9653 -1915 -9650
rect -1907 -9653 -1854 -9650
rect -2073 -9655 -2043 -9653
rect -2135 -9667 -2105 -9660
rect -2065 -9662 -2043 -9655
rect -2243 -9678 -2240 -9669
rect -2221 -9675 -2213 -9667
rect -2211 -9675 -2208 -9667
rect -2203 -9674 -2173 -9667
rect -2251 -9685 -2240 -9678
rect -2211 -9678 -2203 -9675
rect -2211 -9685 -2181 -9678
rect -2073 -9685 -2043 -9678
rect -2203 -9708 -2173 -9701
rect -2262 -9726 -2240 -9716
rect -2203 -9717 -2176 -9708
rect -2083 -9719 -2075 -9709
rect -2040 -9719 -2035 -9715
rect -2073 -9731 -2043 -9719
rect -2028 -9731 -2023 -9719
rect -2000 -9726 -1992 -9653
rect -1963 -9656 -1955 -9653
rect -1963 -9657 -1915 -9656
rect -1955 -9667 -1907 -9660
rect -1885 -9664 -1877 -9653
rect -1837 -9658 -1828 -9642
rect -1758 -9649 -1750 -9634
rect -1758 -9650 -1692 -9649
rect -1837 -9660 -1833 -9658
rect -1837 -9662 -1835 -9660
rect -1887 -9667 -1851 -9664
rect -1750 -9667 -1702 -9660
rect -1885 -9672 -1877 -9667
rect -1963 -9685 -1915 -9678
rect -1905 -9717 -1897 -9672
rect -1857 -9690 -1851 -9667
rect -1760 -9675 -1758 -9674
rect -1837 -9685 -1789 -9678
rect -1758 -9684 -1750 -9678
rect -1758 -9685 -1710 -9684
rect -1955 -9720 -1915 -9717
rect -1963 -9726 -1962 -9724
rect -2000 -9729 -1981 -9726
rect -1965 -9729 -1962 -9726
rect -1955 -9726 -1907 -9722
rect -1885 -9726 -1877 -9707
rect -1857 -9720 -1851 -9708
rect -1750 -9712 -1702 -9705
rect -1829 -9720 -1789 -9718
rect -1766 -9722 -1760 -9712
rect -1829 -9726 -1781 -9722
rect -1756 -9726 -1740 -9722
rect -1680 -9726 -1672 -9608
rect -1671 -9614 -1663 -9606
rect -1645 -9610 -1637 -9594
rect -1663 -9622 -1655 -9614
rect -1671 -9642 -1663 -9634
rect -1663 -9650 -1655 -9642
rect -1671 -9670 -1663 -9662
rect -1671 -9686 -1669 -9673
rect -1663 -9678 -1655 -9670
rect -1671 -9698 -1663 -9690
rect -1663 -9706 -1655 -9698
rect -1671 -9726 -1663 -9718
rect -1955 -9729 -1837 -9726
rect -1829 -9729 -1740 -9726
rect -2206 -9739 -2176 -9736
rect -2206 -9742 -2203 -9739
rect -2161 -9741 -2145 -9732
rect -2073 -9734 -2065 -9731
rect -2073 -9735 -2043 -9734
rect -2028 -9735 -2012 -9731
rect -2073 -9742 -2065 -9736
rect -2203 -9743 -2176 -9742
rect -2065 -9743 -2043 -9742
rect -2262 -9749 -2232 -9743
rect -2176 -9749 -2173 -9743
rect -2043 -9749 -2035 -9743
rect -2325 -9774 -2320 -9754
rect -2317 -9762 -2309 -9754
rect -2153 -9755 -2146 -9751
rect -2325 -9782 -2317 -9774
rect -2300 -9778 -2292 -9768
rect -2325 -9802 -2320 -9782
rect -2317 -9790 -2309 -9782
rect -2325 -9810 -2317 -9802
rect -2325 -9830 -2320 -9810
rect -2317 -9818 -2309 -9810
rect -2290 -9811 -2282 -9778
rect -2273 -9782 -2264 -9777
rect -2206 -9782 -2176 -9777
rect -2262 -9789 -2232 -9784
rect -2198 -9793 -2176 -9782
rect -2198 -9807 -2176 -9799
rect -2166 -9815 -2158 -9767
rect -2143 -9771 -2136 -9755
rect -2143 -9782 -2113 -9777
rect -2073 -9782 -2065 -9777
rect -2065 -9784 -2043 -9782
rect -2043 -9789 -2035 -9784
rect -2065 -9810 -2043 -9795
rect -2006 -9811 -2004 -9795
rect -2265 -9825 -2260 -9819
rect -2143 -9825 -2113 -9818
rect -2270 -9826 -2240 -9825
rect -2270 -9829 -2265 -9826
rect -2325 -9838 -2317 -9830
rect -2325 -9858 -2320 -9838
rect -2317 -9846 -2309 -9838
rect -2113 -9841 -2105 -9831
rect -2291 -9853 -2270 -9846
rect -2198 -9848 -2168 -9846
rect -2135 -9847 -2105 -9846
rect -2103 -9847 -2095 -9841
rect -2113 -9848 -2105 -9847
rect -2065 -9848 -2035 -9846
rect -2000 -9848 -1992 -9729
rect -1963 -9736 -1960 -9729
rect -1915 -9733 -1905 -9729
rect -1963 -9737 -1955 -9736
rect -1963 -9743 -1915 -9737
rect -1989 -9770 -1973 -9767
rect -1915 -9770 -1907 -9763
rect -1990 -9805 -1989 -9784
rect -1983 -9848 -1981 -9785
rect -1885 -9794 -1877 -9729
rect -1789 -9734 -1778 -9729
rect -1837 -9737 -1829 -9736
rect -1837 -9743 -1789 -9737
rect -1756 -9738 -1740 -9729
rect -1837 -9753 -1829 -9743
rect -1872 -9772 -1867 -9762
rect -1789 -9770 -1781 -9763
rect -1776 -9770 -1769 -9753
rect -1756 -9760 -1750 -9738
rect -1671 -9742 -1669 -9731
rect -1663 -9734 -1655 -9726
rect -1671 -9754 -1663 -9746
rect -1663 -9762 -1655 -9754
rect -1702 -9772 -1696 -9766
rect -1955 -9796 -1915 -9794
rect -1963 -9798 -1955 -9796
rect -1963 -9805 -1915 -9798
rect -1963 -9813 -1955 -9805
rect -1963 -9814 -1915 -9813
rect -1973 -9820 -1965 -9817
rect -1955 -9820 -1907 -9816
rect -1974 -9823 -1907 -9820
rect -1973 -9827 -1965 -9823
rect -1963 -9827 -1960 -9825
rect -1963 -9831 -1915 -9827
rect -1963 -9839 -1955 -9831
rect -1963 -9843 -1915 -9839
rect -1963 -9846 -1955 -9843
rect -2240 -9853 -2206 -9848
rect -2198 -9853 -2143 -9848
rect -2113 -9853 -1981 -9848
rect -1915 -9853 -1907 -9846
rect -2270 -9858 -2266 -9854
rect -2086 -9857 -2070 -9853
rect -2325 -9866 -2317 -9858
rect -2270 -9865 -2240 -9858
rect -2206 -9865 -2176 -9858
rect -2325 -9886 -2320 -9866
rect -2317 -9874 -2309 -9866
rect -2270 -9870 -2266 -9865
rect -2270 -9874 -2266 -9871
rect -2198 -9874 -2176 -9867
rect -2166 -9874 -2158 -9857
rect -2143 -9865 -2113 -9858
rect -2198 -9883 -2168 -9879
rect -2325 -9894 -2317 -9886
rect -2143 -9888 -2136 -9874
rect -2085 -9879 -2060 -9878
rect -2039 -9879 -2035 -9870
rect -2135 -9886 -2105 -9879
rect -2085 -9886 -2035 -9879
rect -2029 -9886 -2025 -9879
rect -2325 -9907 -2320 -9894
rect -2317 -9902 -2309 -9894
rect -2235 -9904 -2232 -9901
rect -2325 -9933 -2317 -9907
rect -2325 -9942 -2320 -9933
rect -2325 -9950 -2317 -9942
rect -2135 -9950 -2119 -9937
rect -2000 -9945 -1992 -9853
rect -1983 -9871 -1981 -9853
rect -1955 -9871 -1915 -9870
rect -1862 -9874 -1857 -9772
rect -1706 -9776 -1702 -9772
rect -1829 -9788 -1789 -9780
rect -1671 -9782 -1663 -9774
rect -1849 -9796 -1842 -9788
rect -1790 -9796 -1781 -9788
rect -1663 -9790 -1655 -9782
rect -1837 -9805 -1829 -9798
rect -1758 -9805 -1732 -9798
rect -1748 -9814 -1732 -9805
rect -1671 -9810 -1663 -9802
rect -1829 -9823 -1781 -9816
rect -1663 -9818 -1655 -9810
rect -1829 -9829 -1789 -9825
rect -1768 -9828 -1760 -9818
rect -1758 -9829 -1750 -9828
rect -1671 -9838 -1663 -9830
rect -1837 -9841 -1780 -9838
rect -1758 -9844 -1748 -9838
rect -1708 -9844 -1690 -9838
rect -1829 -9853 -1781 -9846
rect -1680 -9855 -1672 -9838
rect -1663 -9846 -1655 -9838
rect -1829 -9864 -1791 -9858
rect -1758 -9864 -1710 -9862
rect -1758 -9871 -1692 -9864
rect -1671 -9866 -1663 -9858
rect -1955 -9882 -1907 -9879
rect -1791 -9882 -1781 -9879
rect -1991 -9886 -1839 -9882
rect -1791 -9886 -1780 -9882
rect -1680 -9889 -1672 -9871
rect -1663 -9874 -1655 -9866
rect -1839 -9899 -1791 -9892
rect -1671 -9894 -1663 -9886
rect -1829 -9905 -1791 -9901
rect -1671 -9904 -1669 -9894
rect -1663 -9902 -1655 -9894
rect -1680 -9920 -1672 -9905
rect -1642 -9920 -1637 -9610
rect -1619 -9446 -1612 -9422
rect -1619 -9660 -1614 -9446
rect -1619 -9686 -1611 -9660
rect -1554 -9674 -1547 -9661
rect -1530 -9684 -1526 -8385
rect -1506 -8413 -1502 -8221
rect -1506 -8461 -1499 -8413
rect -1554 -9685 -1547 -9684
rect -1768 -9936 -1760 -9926
rect -1758 -9943 -1710 -9936
rect -2325 -9970 -2320 -9950
rect -2317 -9958 -2306 -9950
rect -2031 -9953 -1992 -9945
rect -1750 -9947 -1710 -9943
rect -1674 -9948 -1663 -9942
rect -2307 -9966 -2306 -9958
rect -2149 -9955 -2135 -9954
rect -2149 -9959 -2119 -9955
rect -2024 -9964 -2021 -9955
rect -2325 -9978 -2317 -9970
rect -2325 -10026 -2320 -9978
rect -2317 -9986 -2306 -9978
rect -2185 -9980 -2169 -9968
rect -2056 -9971 -2040 -9967
rect -2021 -9971 -2008 -9964
rect -2056 -9982 -2054 -9972
rect -2056 -9983 -2048 -9982
rect -2307 -10022 -2306 -10014
rect -2111 -10015 -2054 -10009
rect -2325 -10034 -2314 -10026
rect -2104 -10033 -2101 -10029
rect -2325 -10054 -2320 -10034
rect -2314 -10042 -2306 -10034
rect -2104 -10036 -2101 -10034
rect -2084 -10036 -2054 -10035
rect -2000 -10036 -1992 -9953
rect -1758 -9954 -1750 -9953
rect -1758 -9955 -1749 -9954
rect -1758 -9956 -1710 -9955
rect -1663 -9958 -1658 -9948
rect -1831 -9966 -1783 -9962
rect -1784 -9979 -1783 -9966
rect -1674 -9976 -1663 -9970
rect -1826 -9981 -1796 -9980
rect -1663 -9986 -1658 -9976
rect -1654 -9980 -1647 -9970
rect -1644 -9994 -1637 -9980
rect -1758 -10012 -1750 -10009
rect -1758 -10015 -1710 -10012
rect -1844 -10027 -1828 -10025
rect -1844 -10028 -1792 -10027
rect -1828 -10029 -1792 -10028
rect -1772 -10029 -1758 -10021
rect -1750 -10024 -1702 -10017
rect -1750 -10032 -1710 -10028
rect -1700 -10032 -1692 -10012
rect -1674 -10020 -1665 -10012
rect -1674 -10032 -1666 -10024
rect -1758 -10036 -1710 -10035
rect -2307 -10050 -2306 -10042
rect -2139 -10046 -2123 -10037
rect -2111 -10042 -2016 -10036
rect -2139 -10053 -2111 -10046
rect -2325 -10062 -2314 -10054
rect -2177 -10060 -2161 -10059
rect -2141 -10060 -2119 -10058
rect -2104 -10060 -2101 -10042
rect -2076 -10053 -2046 -10048
rect -2325 -10070 -2320 -10062
rect -2314 -10070 -2306 -10062
rect -2076 -10064 -2054 -10058
rect -2021 -10061 -2016 -10042
rect -2000 -10042 -1818 -10036
rect -1802 -10042 -1776 -10036
rect -1760 -10042 -1710 -10036
rect -1666 -10040 -1658 -10032
rect -2189 -10070 -2175 -10065
rect -2373 -10072 -2175 -10070
rect -2373 -10073 -2359 -10072
rect -2371 -10485 -2366 -10073
rect -2348 -10125 -2343 -10072
rect -2325 -10082 -2320 -10072
rect -2307 -10078 -2306 -10072
rect -2189 -10073 -2175 -10072
rect -2149 -10074 -2119 -10065
rect -2084 -10066 -2036 -10065
rect -2000 -10066 -1992 -10042
rect -1758 -10044 -1710 -10042
rect -1758 -10046 -1755 -10044
rect -1828 -10053 -1792 -10046
rect -1768 -10055 -1760 -10048
rect -1758 -10053 -1757 -10046
rect -1710 -10047 -1702 -10046
rect -1750 -10053 -1702 -10047
rect -1674 -10048 -1665 -10040
rect -1768 -10058 -1764 -10055
rect -1758 -10058 -1755 -10053
rect -1818 -10066 -1789 -10058
rect -1758 -10065 -1754 -10058
rect -1750 -10063 -1710 -10058
rect -1674 -10060 -1666 -10052
rect -1758 -10066 -1692 -10065
rect -2084 -10068 -1692 -10066
rect -1666 -10068 -1658 -10060
rect -2084 -10071 -1690 -10068
rect -2084 -10074 -2054 -10071
rect -2046 -10073 -1710 -10071
rect -2325 -10090 -2314 -10082
rect -2076 -10083 -2046 -10076
rect -2325 -10110 -2320 -10090
rect -2314 -10098 -2306 -10090
rect -2076 -10091 -2054 -10085
rect -2084 -10095 -2054 -10093
rect -2104 -10098 -2054 -10095
rect -2307 -10106 -2306 -10098
rect -2084 -10101 -2054 -10098
rect -2325 -10122 -2314 -10110
rect -2348 -10149 -2341 -10125
rect -2325 -10139 -2320 -10122
rect -2314 -10126 -2309 -10122
rect -2309 -10138 -2298 -10126
rect -2314 -10139 -2309 -10138
rect -2361 -10465 -2353 -10455
rect -2348 -10465 -2343 -10149
rect -2351 -10481 -2343 -10465
rect -2371 -10511 -2363 -10485
rect -2383 -10683 -2376 -10673
rect -2371 -10683 -2366 -10511
rect -2373 -10694 -2366 -10683
rect -2348 -10694 -2343 -10481
rect -2325 -10151 -2314 -10139
rect -2076 -10150 -2073 -10134
rect -2325 -10168 -2320 -10151
rect -2314 -10154 -2309 -10151
rect -2309 -10166 -2298 -10154
rect -2251 -10158 -2101 -10151
rect -2141 -10165 -2111 -10159
rect -2086 -10161 -2083 -10151
rect -2076 -10165 -2046 -10159
rect -2314 -10168 -2309 -10166
rect -2325 -10180 -2314 -10168
rect -2141 -10177 -2113 -10172
rect -2076 -10177 -2073 -10174
rect -2325 -10199 -2320 -10180
rect -2314 -10182 -2309 -10180
rect -2325 -10209 -2317 -10199
rect -2325 -10228 -2320 -10209
rect -2317 -10215 -2309 -10209
rect -2243 -10226 -2221 -10218
rect -2211 -10226 -2201 -10206
rect -2073 -10226 -2065 -10208
rect -2000 -10226 -1992 -10073
rect -1758 -10074 -1710 -10073
rect -1680 -10076 -1665 -10068
rect -1750 -10083 -1702 -10076
rect -1680 -10080 -1672 -10076
rect -1680 -10085 -1666 -10080
rect -1836 -10089 -1820 -10088
rect -1837 -10093 -1820 -10089
rect -1750 -10091 -1710 -10085
rect -1674 -10088 -1666 -10085
rect -1837 -10100 -1789 -10093
rect -1758 -10094 -1710 -10093
rect -1760 -10097 -1692 -10094
rect -1666 -10096 -1658 -10088
rect -1837 -10101 -1820 -10100
rect -1764 -10101 -1692 -10097
rect -1674 -10101 -1665 -10096
rect -1680 -10104 -1665 -10101
rect -1680 -10132 -1672 -10104
rect -1666 -10124 -1665 -10114
rect -1837 -10134 -1789 -10132
rect -1829 -10148 -1789 -10134
rect -1655 -10136 -1650 -10126
rect -1666 -10142 -1655 -10136
rect -1778 -10150 -1771 -10148
rect -1710 -10150 -1702 -10148
rect -1666 -10152 -1665 -10142
rect -1837 -10158 -1829 -10152
rect -1829 -10159 -1789 -10158
rect -1726 -10159 -1710 -10158
rect -1789 -10161 -1781 -10159
rect -1829 -10165 -1781 -10161
rect -1750 -10165 -1710 -10159
rect -1829 -10177 -1789 -10168
rect -1726 -10174 -1710 -10165
rect -1706 -10174 -1702 -10161
rect -1655 -10164 -1650 -10154
rect -1666 -10170 -1655 -10164
rect -1666 -10180 -1665 -10170
rect -1671 -10210 -1663 -10202
rect -1655 -10210 -1647 -10208
rect -1663 -10218 -1647 -10210
rect -1642 -10218 -1637 -9994
rect -1619 -9996 -1614 -9686
rect -1530 -9709 -1523 -9685
rect -1885 -10226 -1877 -10224
rect -1708 -10226 -1672 -10224
rect -2243 -10227 -2213 -10226
rect -2325 -10237 -2317 -10228
rect -2259 -10233 -2211 -10227
rect -2183 -10233 -1877 -10226
rect -1869 -10233 -1758 -10226
rect -1710 -10232 -1672 -10226
rect -1710 -10233 -1692 -10232
rect -2211 -10237 -2201 -10233
rect -2325 -10257 -2320 -10237
rect -2317 -10244 -2309 -10237
rect -2211 -10244 -2198 -10237
rect -2325 -10265 -2317 -10257
rect -2300 -10264 -2292 -10254
rect -2243 -10263 -2228 -10252
rect -2211 -10260 -2181 -10244
rect -2211 -10263 -2201 -10260
rect -2325 -10285 -2320 -10265
rect -2317 -10273 -2309 -10265
rect -2325 -10293 -2317 -10285
rect -2325 -10313 -2320 -10293
rect -2317 -10301 -2309 -10293
rect -2325 -10322 -2317 -10313
rect -2325 -10341 -2320 -10322
rect -2317 -10329 -2309 -10322
rect -2325 -10350 -2317 -10341
rect -2325 -10370 -2320 -10350
rect -2317 -10357 -2309 -10350
rect -2325 -10378 -2317 -10370
rect -2290 -10377 -2282 -10264
rect -2251 -10274 -2240 -10270
rect -2211 -10274 -2181 -10270
rect -2251 -10277 -2181 -10274
rect -2176 -10284 -2173 -10282
rect -2240 -10291 -2173 -10284
rect -2169 -10289 -2163 -10234
rect -2073 -10270 -2065 -10233
rect -2073 -10274 -2043 -10270
rect -2000 -10274 -1992 -10233
rect -1915 -10264 -1907 -10255
rect -1963 -10270 -1955 -10264
rect -1963 -10274 -1915 -10270
rect -1885 -10274 -1877 -10233
rect -1875 -10238 -1869 -10234
rect -1829 -10256 -1781 -10254
rect -1847 -10260 -1781 -10256
rect -1778 -10260 -1771 -10234
rect -1758 -10241 -1710 -10234
rect -1718 -10248 -1710 -10241
rect -1768 -10258 -1760 -10248
rect -1718 -10250 -1700 -10248
rect -2146 -10277 -2135 -10274
rect -2105 -10277 -2043 -10274
rect -2035 -10277 -1989 -10274
rect -1973 -10277 -1915 -10274
rect -1907 -10277 -1854 -10274
rect -2073 -10279 -2043 -10277
rect -2135 -10291 -2105 -10284
rect -2065 -10286 -2043 -10279
rect -2243 -10302 -2240 -10293
rect -2221 -10299 -2213 -10291
rect -2211 -10299 -2208 -10291
rect -2203 -10298 -2173 -10291
rect -2251 -10309 -2240 -10302
rect -2211 -10302 -2203 -10299
rect -2211 -10309 -2181 -10302
rect -2073 -10309 -2043 -10302
rect -2203 -10332 -2173 -10325
rect -2262 -10350 -2240 -10340
rect -2203 -10341 -2176 -10332
rect -2083 -10343 -2075 -10333
rect -2040 -10343 -2035 -10339
rect -2073 -10355 -2043 -10343
rect -2028 -10355 -2023 -10343
rect -2000 -10350 -1992 -10277
rect -1963 -10280 -1955 -10277
rect -1963 -10281 -1915 -10280
rect -1955 -10291 -1907 -10284
rect -1885 -10288 -1877 -10277
rect -1837 -10282 -1828 -10266
rect -1758 -10273 -1750 -10258
rect -1758 -10274 -1692 -10273
rect -1837 -10284 -1833 -10282
rect -1837 -10286 -1835 -10284
rect -1887 -10291 -1851 -10288
rect -1750 -10291 -1702 -10284
rect -1885 -10296 -1877 -10291
rect -1963 -10309 -1915 -10302
rect -1905 -10341 -1897 -10296
rect -1857 -10314 -1851 -10291
rect -1760 -10299 -1758 -10298
rect -1837 -10309 -1789 -10302
rect -1758 -10308 -1750 -10302
rect -1758 -10309 -1710 -10308
rect -1955 -10344 -1915 -10341
rect -1963 -10350 -1962 -10348
rect -2000 -10353 -1981 -10350
rect -1965 -10353 -1962 -10350
rect -1955 -10350 -1907 -10346
rect -1885 -10350 -1877 -10331
rect -1857 -10344 -1851 -10332
rect -1750 -10336 -1702 -10329
rect -1829 -10344 -1789 -10342
rect -1766 -10346 -1760 -10336
rect -1829 -10350 -1781 -10346
rect -1756 -10350 -1740 -10346
rect -1680 -10350 -1672 -10232
rect -1671 -10238 -1663 -10230
rect -1645 -10234 -1637 -10218
rect -1663 -10246 -1655 -10238
rect -1671 -10266 -1663 -10258
rect -1663 -10274 -1655 -10266
rect -1671 -10294 -1663 -10286
rect -1671 -10310 -1669 -10297
rect -1663 -10302 -1655 -10294
rect -1671 -10322 -1663 -10314
rect -1663 -10330 -1655 -10322
rect -1671 -10350 -1663 -10342
rect -1955 -10353 -1837 -10350
rect -1829 -10353 -1740 -10350
rect -2206 -10363 -2176 -10360
rect -2206 -10366 -2203 -10363
rect -2161 -10365 -2145 -10356
rect -2073 -10358 -2065 -10355
rect -2073 -10359 -2043 -10358
rect -2028 -10359 -2012 -10355
rect -2073 -10366 -2065 -10360
rect -2203 -10367 -2176 -10366
rect -2065 -10367 -2043 -10366
rect -2262 -10373 -2232 -10367
rect -2176 -10373 -2173 -10367
rect -2043 -10373 -2035 -10367
rect -2325 -10398 -2320 -10378
rect -2317 -10386 -2309 -10378
rect -2153 -10379 -2146 -10375
rect -2325 -10406 -2317 -10398
rect -2300 -10402 -2292 -10392
rect -2325 -10426 -2320 -10406
rect -2317 -10414 -2309 -10406
rect -2325 -10434 -2317 -10426
rect -2325 -10454 -2320 -10434
rect -2317 -10442 -2309 -10434
rect -2290 -10435 -2282 -10402
rect -2273 -10406 -2264 -10401
rect -2206 -10406 -2176 -10401
rect -2262 -10413 -2232 -10408
rect -2198 -10417 -2176 -10406
rect -2198 -10431 -2176 -10423
rect -2166 -10439 -2158 -10391
rect -2143 -10395 -2136 -10379
rect -2143 -10406 -2113 -10401
rect -2073 -10406 -2065 -10401
rect -2065 -10408 -2043 -10406
rect -2043 -10413 -2035 -10408
rect -2065 -10434 -2043 -10419
rect -2006 -10435 -2004 -10419
rect -2265 -10449 -2260 -10443
rect -2143 -10449 -2113 -10442
rect -2270 -10450 -2240 -10449
rect -2270 -10453 -2265 -10450
rect -2325 -10462 -2317 -10454
rect -2325 -10482 -2320 -10462
rect -2317 -10470 -2309 -10462
rect -2113 -10465 -2105 -10455
rect -2291 -10477 -2270 -10470
rect -2198 -10472 -2168 -10470
rect -2135 -10471 -2105 -10470
rect -2103 -10471 -2095 -10465
rect -2113 -10472 -2105 -10471
rect -2065 -10472 -2035 -10470
rect -2000 -10472 -1992 -10353
rect -1963 -10360 -1960 -10353
rect -1915 -10357 -1905 -10353
rect -1963 -10361 -1955 -10360
rect -1963 -10367 -1915 -10361
rect -1989 -10394 -1973 -10391
rect -1915 -10394 -1907 -10387
rect -1990 -10429 -1989 -10408
rect -1983 -10472 -1981 -10409
rect -1885 -10418 -1877 -10353
rect -1789 -10358 -1778 -10353
rect -1837 -10361 -1829 -10360
rect -1837 -10367 -1789 -10361
rect -1756 -10362 -1740 -10353
rect -1837 -10377 -1829 -10367
rect -1872 -10396 -1867 -10386
rect -1789 -10394 -1781 -10387
rect -1776 -10394 -1769 -10377
rect -1756 -10384 -1750 -10362
rect -1671 -10366 -1669 -10355
rect -1663 -10358 -1655 -10350
rect -1671 -10378 -1663 -10370
rect -1663 -10386 -1655 -10378
rect -1702 -10396 -1696 -10390
rect -1955 -10420 -1915 -10418
rect -1963 -10422 -1955 -10420
rect -1963 -10429 -1915 -10422
rect -1963 -10437 -1955 -10429
rect -1963 -10438 -1915 -10437
rect -1973 -10444 -1965 -10441
rect -1955 -10444 -1907 -10440
rect -1974 -10447 -1907 -10444
rect -1973 -10451 -1965 -10447
rect -1963 -10451 -1960 -10449
rect -1963 -10455 -1915 -10451
rect -1963 -10463 -1955 -10455
rect -1963 -10467 -1915 -10463
rect -1963 -10470 -1955 -10467
rect -2240 -10477 -2206 -10472
rect -2198 -10477 -2143 -10472
rect -2113 -10477 -1981 -10472
rect -1915 -10477 -1907 -10470
rect -2270 -10482 -2266 -10478
rect -2086 -10481 -2070 -10477
rect -2325 -10490 -2317 -10482
rect -2270 -10489 -2240 -10482
rect -2206 -10489 -2176 -10482
rect -2325 -10510 -2320 -10490
rect -2317 -10498 -2309 -10490
rect -2270 -10494 -2266 -10489
rect -2270 -10498 -2266 -10495
rect -2198 -10498 -2176 -10491
rect -2166 -10498 -2158 -10481
rect -2143 -10489 -2113 -10482
rect -2198 -10507 -2168 -10503
rect -2325 -10518 -2317 -10510
rect -2143 -10512 -2136 -10498
rect -2085 -10503 -2060 -10502
rect -2039 -10503 -2035 -10494
rect -2135 -10510 -2105 -10503
rect -2085 -10510 -2035 -10503
rect -2029 -10510 -2025 -10503
rect -2325 -10531 -2320 -10518
rect -2317 -10526 -2309 -10518
rect -2235 -10528 -2232 -10525
rect -2325 -10557 -2317 -10531
rect -2325 -10566 -2320 -10557
rect -2325 -10574 -2317 -10566
rect -2135 -10574 -2119 -10561
rect -2000 -10569 -1992 -10477
rect -1983 -10495 -1981 -10477
rect -1955 -10495 -1915 -10494
rect -1862 -10498 -1857 -10396
rect -1706 -10400 -1702 -10396
rect -1829 -10412 -1789 -10404
rect -1671 -10406 -1663 -10398
rect -1849 -10420 -1842 -10412
rect -1790 -10420 -1781 -10412
rect -1663 -10414 -1655 -10406
rect -1837 -10429 -1829 -10422
rect -1758 -10429 -1732 -10422
rect -1748 -10438 -1732 -10429
rect -1671 -10434 -1663 -10426
rect -1829 -10447 -1781 -10440
rect -1663 -10442 -1655 -10434
rect -1829 -10453 -1789 -10449
rect -1768 -10452 -1760 -10442
rect -1758 -10453 -1750 -10452
rect -1671 -10462 -1663 -10454
rect -1837 -10465 -1780 -10462
rect -1758 -10468 -1748 -10462
rect -1708 -10468 -1690 -10462
rect -1829 -10477 -1781 -10470
rect -1680 -10479 -1672 -10462
rect -1663 -10470 -1655 -10462
rect -1829 -10488 -1791 -10482
rect -1758 -10488 -1710 -10486
rect -1758 -10495 -1692 -10488
rect -1671 -10490 -1663 -10482
rect -1955 -10506 -1907 -10503
rect -1791 -10506 -1781 -10503
rect -1991 -10510 -1839 -10506
rect -1791 -10510 -1780 -10506
rect -1680 -10513 -1672 -10495
rect -1663 -10498 -1655 -10490
rect -1839 -10523 -1791 -10516
rect -1671 -10518 -1663 -10510
rect -1829 -10529 -1791 -10525
rect -1671 -10528 -1669 -10518
rect -1663 -10526 -1655 -10518
rect -1680 -10544 -1672 -10529
rect -1642 -10544 -1637 -10234
rect -1619 -10070 -1612 -10046
rect -1619 -10284 -1614 -10070
rect -1530 -10246 -1526 -9709
rect -1517 -10003 -1512 -9993
rect -1506 -10003 -1502 -8461
rect -1493 -9019 -1488 -9009
rect -1482 -9019 -1478 -8172
rect -1469 -8203 -1464 -8193
rect -1458 -8203 -1454 -8172
rect -1459 -8217 -1454 -8203
rect -1469 -8218 -1435 -8217
rect -1434 -8218 -1430 -8172
rect -1410 -8218 -1406 -8172
rect -1397 -8179 -1392 -8172
rect -1386 -8179 -1382 -8172
rect -1373 -8179 -1368 -8172
rect -1387 -8193 -1382 -8179
rect -1363 -8193 -1358 -8179
rect -1397 -8203 -1392 -8193
rect -1387 -8217 -1382 -8203
rect -1386 -8218 -1382 -8217
rect -1362 -8218 -1358 -8193
rect -1338 -8218 -1334 -8172
rect -1314 -8217 -1310 -8172
rect -1301 -8203 -1296 -8193
rect -1290 -8203 -1286 -8172
rect -1277 -8179 -1272 -8172
rect -1266 -8179 -1262 -8172
rect -1267 -8193 -1262 -8179
rect -1253 -8186 -1248 -8183
rect -1291 -8217 -1286 -8203
rect -1325 -8218 -1291 -8217
rect -1469 -8220 -1291 -8218
rect -1469 -8227 -1464 -8220
rect -1459 -8241 -1454 -8227
rect -1469 -8755 -1464 -8745
rect -1458 -8755 -1454 -8241
rect -1459 -8769 -1454 -8755
rect -1434 -8269 -1430 -8220
rect -1434 -8317 -1427 -8269
rect -1469 -8779 -1464 -8769
rect -1459 -8793 -1454 -8779
rect -1469 -8971 -1464 -8961
rect -1458 -8971 -1454 -8793
rect -1459 -8985 -1454 -8971
rect -1434 -8821 -1430 -8317
rect -1434 -8869 -1427 -8821
rect -1469 -8995 -1464 -8985
rect -1459 -9009 -1454 -8995
rect -1483 -9033 -1478 -9019
rect -1493 -9043 -1488 -9033
rect -1483 -9057 -1478 -9043
rect -1493 -9379 -1488 -9369
rect -1482 -9379 -1478 -9057
rect -1483 -9393 -1478 -9379
rect -1458 -9085 -1454 -9009
rect -1445 -9043 -1440 -9033
rect -1434 -9037 -1430 -8869
rect -1421 -8995 -1416 -8985
rect -1410 -8995 -1406 -8220
rect -1397 -8395 -1392 -8385
rect -1386 -8395 -1382 -8220
rect -1387 -8409 -1382 -8395
rect -1362 -8245 -1358 -8220
rect -1338 -8221 -1334 -8220
rect -1362 -8293 -1355 -8245
rect -1338 -8269 -1331 -8221
rect -1325 -8227 -1320 -8220
rect -1314 -8227 -1310 -8220
rect -1315 -8241 -1310 -8227
rect -1396 -8422 -1392 -8412
rect -1362 -8422 -1358 -8293
rect -1349 -8371 -1344 -8361
rect -1338 -8371 -1334 -8269
rect -1339 -8385 -1334 -8371
rect -1397 -8779 -1392 -8769
rect -1386 -8779 -1382 -8422
rect -1387 -8793 -1382 -8779
rect -1411 -9009 -1406 -8995
rect -1434 -9043 -1427 -9037
rect -1435 -9057 -1427 -9043
rect -1458 -9133 -1451 -9085
rect -1492 -9406 -1488 -9396
rect -1458 -9406 -1454 -9133
rect -1493 -9619 -1488 -9609
rect -1482 -9619 -1478 -9406
rect -1483 -9633 -1478 -9619
rect -1507 -10017 -1502 -10003
rect -1619 -10310 -1611 -10284
rect -1554 -10298 -1547 -10285
rect -1554 -10309 -1547 -10308
rect -1768 -10560 -1760 -10550
rect -1758 -10567 -1710 -10560
rect -2325 -10594 -2320 -10574
rect -2317 -10582 -2306 -10574
rect -2031 -10577 -1992 -10569
rect -1750 -10571 -1710 -10567
rect -1674 -10572 -1663 -10566
rect -2307 -10590 -2306 -10582
rect -2149 -10579 -2135 -10578
rect -2149 -10583 -2119 -10579
rect -2024 -10588 -2021 -10579
rect -2325 -10602 -2317 -10594
rect -2325 -10650 -2320 -10602
rect -2317 -10610 -2306 -10602
rect -2185 -10604 -2169 -10592
rect -2056 -10595 -2040 -10591
rect -2021 -10595 -2008 -10588
rect -2056 -10606 -2054 -10596
rect -2056 -10607 -2048 -10606
rect -2307 -10646 -2306 -10638
rect -2111 -10639 -2054 -10633
rect -2325 -10658 -2314 -10650
rect -2104 -10657 -2101 -10653
rect -2325 -10678 -2320 -10658
rect -2314 -10666 -2306 -10658
rect -2104 -10660 -2101 -10658
rect -2084 -10660 -2054 -10659
rect -2000 -10660 -1992 -10577
rect -1758 -10578 -1750 -10577
rect -1758 -10579 -1749 -10578
rect -1758 -10580 -1710 -10579
rect -1663 -10582 -1658 -10572
rect -1831 -10590 -1783 -10586
rect -1784 -10603 -1783 -10590
rect -1674 -10600 -1663 -10594
rect -1826 -10605 -1796 -10604
rect -1663 -10610 -1658 -10600
rect -1654 -10604 -1647 -10594
rect -1644 -10618 -1637 -10604
rect -1758 -10636 -1750 -10633
rect -1758 -10639 -1710 -10636
rect -1844 -10651 -1828 -10649
rect -1844 -10652 -1792 -10651
rect -1828 -10653 -1792 -10652
rect -1772 -10653 -1758 -10645
rect -1750 -10648 -1702 -10641
rect -1750 -10656 -1710 -10652
rect -1700 -10656 -1692 -10636
rect -1674 -10644 -1665 -10636
rect -1674 -10656 -1666 -10648
rect -1758 -10660 -1710 -10659
rect -2307 -10674 -2306 -10666
rect -2139 -10670 -2123 -10661
rect -2111 -10666 -2016 -10660
rect -2139 -10677 -2111 -10670
rect -2325 -10686 -2314 -10678
rect -2177 -10684 -2161 -10683
rect -2141 -10684 -2119 -10682
rect -2104 -10684 -2101 -10666
rect -2076 -10677 -2046 -10672
rect -2325 -10694 -2320 -10686
rect -2314 -10694 -2306 -10686
rect -2076 -10688 -2054 -10682
rect -2021 -10685 -2016 -10666
rect -2000 -10666 -1818 -10660
rect -1802 -10666 -1776 -10660
rect -1760 -10666 -1710 -10660
rect -1666 -10664 -1658 -10656
rect -2189 -10694 -2175 -10689
rect -2373 -10696 -2175 -10694
rect -2373 -10697 -2359 -10696
rect -2371 -10736 -2366 -10697
rect -2348 -10736 -2343 -10696
rect -2325 -10706 -2320 -10696
rect -2307 -10702 -2306 -10696
rect -2189 -10697 -2175 -10696
rect -2149 -10698 -2119 -10689
rect -2084 -10690 -2036 -10689
rect -2000 -10690 -1992 -10666
rect -1758 -10668 -1710 -10666
rect -1758 -10670 -1755 -10668
rect -1828 -10677 -1792 -10670
rect -1768 -10679 -1760 -10672
rect -1758 -10677 -1757 -10670
rect -1710 -10671 -1702 -10670
rect -1750 -10677 -1702 -10671
rect -1674 -10672 -1665 -10664
rect -1768 -10682 -1764 -10679
rect -1758 -10682 -1755 -10677
rect -1818 -10690 -1789 -10682
rect -1758 -10689 -1754 -10682
rect -1750 -10687 -1710 -10682
rect -1674 -10684 -1666 -10676
rect -1758 -10690 -1692 -10689
rect -2084 -10692 -1692 -10690
rect -1666 -10692 -1658 -10684
rect -2084 -10695 -1690 -10692
rect -2084 -10698 -2054 -10695
rect -2046 -10697 -1710 -10695
rect -2325 -10714 -2314 -10706
rect -2076 -10707 -2046 -10700
rect -2325 -10736 -2320 -10714
rect -2314 -10722 -2306 -10714
rect -2076 -10715 -2054 -10709
rect -2084 -10719 -2054 -10717
rect -2104 -10722 -2054 -10719
rect -2307 -10730 -2306 -10722
rect -2084 -10725 -2054 -10722
rect -2000 -10736 -1992 -10697
rect -1758 -10698 -1710 -10697
rect -1680 -10700 -1665 -10692
rect -1750 -10707 -1702 -10700
rect -1680 -10704 -1672 -10700
rect -1680 -10709 -1666 -10704
rect -1836 -10713 -1820 -10712
rect -1837 -10717 -1820 -10713
rect -1750 -10715 -1710 -10709
rect -1674 -10712 -1666 -10709
rect -1837 -10724 -1789 -10717
rect -1758 -10718 -1710 -10717
rect -1760 -10721 -1692 -10718
rect -1666 -10720 -1658 -10712
rect -1837 -10725 -1820 -10724
rect -1764 -10725 -1692 -10721
rect -1674 -10725 -1665 -10720
rect -1680 -10728 -1665 -10725
rect -1680 -10736 -1672 -10728
rect -1642 -10736 -1637 -10618
rect -1619 -10620 -1614 -10310
rect -1619 -10694 -1612 -10670
rect -1619 -10736 -1614 -10694
use Datapath/datapath datapath_0
timestamp 1394841956
transform -1 0 32539 0 -1 21385
box -48 0 25445 21228
use Control/control_ROUTED control_ROUTED_0
timestamp 1394990067
transform 0 1 -1578 1 0 -10760
box 24 -823 66735 31762
use Control/control_ROUTED control_ROUTED_1
timestamp 1394990067
transform 0 1 -1570 1 0 -10836
box 24 -823 66735 31762
<< end >>
