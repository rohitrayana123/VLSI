magic
tech c035u
timestamp 1393855782
<< metal1 >>
rect 3541 1464 4583 1474
rect 3421 1442 4487 1452
rect 3181 1420 4295 1430
rect 2941 1399 4103 1409
rect 2821 1377 4007 1387
rect 709 1355 1103 1365
rect 3661 1355 3911 1365
rect 3925 1355 4679 1365
rect 829 1333 1079 1343
rect 1165 1333 1320 1343
rect 1381 1333 1439 1343
rect 3301 1333 3815 1343
rect 3829 1333 4391 1343
rect 925 1311 960 1321
rect 1045 1311 1199 1321
rect 1285 1311 1415 1321
rect 1765 1311 1799 1321
rect 2029 1311 2303 1321
rect 3061 1311 3719 1321
rect 3733 1311 4199 1321
rect 4429 1311 6239 1321
rect 517 1289 671 1299
rect 685 1289 863 1299
rect 877 1289 2903 1299
rect 2917 1289 3143 1299
rect 3157 1289 3383 1299
rect 3397 1289 3623 1299
rect 3637 1289 4799 1299
rect 4813 1289 5135 1299
rect 397 1267 1343 1277
rect 1357 1267 2999 1277
rect 3013 1267 3119 1277
rect 3133 1267 3479 1277
rect 3493 1267 3599 1277
rect 3613 1267 4775 1277
rect 4789 1267 5015 1277
rect 5029 1267 5111 1277
rect 5125 1267 5759 1277
rect 5773 1267 6743 1277
rect 277 1245 647 1255
rect 661 1245 983 1255
rect 997 1245 1559 1255
rect 1573 1245 3215 1255
rect 3229 1245 3335 1255
rect 3349 1245 3455 1255
rect 3469 1245 3575 1255
rect 3589 1245 6719 1255
rect 6949 1245 7007 1255
rect 157 1223 791 1233
rect 805 1223 1223 1233
rect 1237 1223 2663 1233
rect 2677 1223 4751 1233
rect 4837 1223 4870 1233
rect 5197 1223 5255 1233
rect 5701 1223 5879 1233
rect 5941 1223 5975 1233
rect 6085 1223 6119 1233
rect 6133 1223 6335 1233
rect 6349 1223 6455 1233
rect 6469 1223 6575 1233
rect 6805 1223 6983 1233
rect 37 1201 1535 1211
rect 1549 1201 2543 1211
rect 2557 1201 2639 1211
rect 2653 1201 4895 1211
rect 5077 1201 5231 1211
rect 5317 1201 5351 1211
rect 5821 1201 5855 1211
rect 5869 1201 7031 1211
rect 7093 1201 7127 1211
rect 85 382 623 392
rect 637 382 1247 392
rect 1261 382 5375 392
rect 5389 382 5999 392
rect 6013 382 7151 392
rect 205 360 2567 370
rect 2581 360 4991 370
rect 5005 360 6023 370
rect 6037 360 6695 370
rect 6709 360 6839 370
rect 325 338 767 348
rect 781 338 887 348
rect 901 338 1583 348
rect 1597 338 2735 348
rect 2749 338 2855 348
rect 2869 338 2975 348
rect 2989 338 3095 348
rect 3109 338 5399 348
rect 5413 338 5615 348
rect 5629 338 5735 348
rect 5749 338 6863 348
rect 445 316 2759 326
rect 2773 316 2879 326
rect 2893 316 3239 326
rect 3253 316 3359 326
rect 3997 316 4079 326
rect 4093 316 4175 326
rect 4189 316 4271 326
rect 4285 316 4367 326
rect 4381 316 4463 326
rect 4477 316 4559 326
rect 4573 316 4655 326
rect 4982 316 5447 326
rect 6181 316 6215 326
rect 565 294 743 304
rect 757 294 2783 304
rect 2797 294 3023 304
rect 3037 294 3263 304
rect 3277 294 3503 304
rect 3517 294 5639 304
rect 5653 294 6887 304
rect 181 272 1487 282
rect 1501 272 1823 282
rect 1837 272 2183 282
rect 2701 271 3695 281
rect 3709 271 3791 281
rect 3805 271 3887 281
rect 5625 272 6287 282
rect 1645 250 1703 260
rect 2605 249 3983 259
rect 4185 250 4319 260
rect 5413 250 6407 260
rect 210 227 3743 237
rect 3853 227 5519 237
rect 5821 228 6527 238
rect 349 205 1919 215
rect 2077 205 4171 215
rect 4525 205 6695 215
rect 517 183 1991 193
rect 2725 183 4607 193
rect 6181 183 6647 193
rect 541 161 2207 171
rect 3061 161 4703 171
rect 6541 161 7199 171
rect 613 139 2375 149
rect 3181 139 5495 149
rect 829 117 2423 127
rect 3229 117 4415 127
rect 973 95 4943 105
rect 1309 73 4031 83
rect 4957 71 5611 81
rect 1669 51 4127 61
rect 2413 29 4223 39
rect 3397 7 3935 17
<< m2contact >>
rect 3527 1462 3541 1476
rect 4583 1462 4597 1476
rect 3407 1440 3421 1454
rect 4487 1440 4501 1454
rect 3167 1419 3181 1433
rect 4295 1418 4309 1432
rect 2927 1397 2941 1411
rect 4103 1396 4117 1410
rect 2807 1375 2821 1389
rect 4007 1375 4021 1389
rect 695 1353 709 1367
rect 1103 1353 1117 1367
rect 3647 1353 3661 1367
rect 3911 1353 3925 1367
rect 4679 1353 4693 1367
rect 815 1331 829 1345
rect 1079 1331 1093 1345
rect 1151 1331 1165 1345
rect 1320 1331 1334 1345
rect 1367 1331 1381 1345
rect 1439 1331 1453 1345
rect 3287 1331 3301 1345
rect 3815 1331 3829 1345
rect 4391 1331 4405 1345
rect 911 1309 925 1323
rect 960 1309 974 1323
rect 1031 1309 1045 1323
rect 1199 1309 1213 1323
rect 1271 1309 1285 1323
rect 1415 1309 1429 1323
rect 1751 1309 1765 1323
rect 1799 1309 1813 1323
rect 2015 1309 2029 1323
rect 2303 1309 2317 1323
rect 3047 1309 3061 1323
rect 3719 1309 3733 1323
rect 4199 1309 4213 1323
rect 4415 1309 4429 1323
rect 6239 1309 6253 1323
rect 503 1287 517 1301
rect 671 1287 685 1301
rect 863 1287 877 1301
rect 2903 1287 2917 1301
rect 3143 1287 3157 1301
rect 3383 1287 3397 1301
rect 3623 1287 3637 1301
rect 4799 1287 4813 1301
rect 5135 1287 5149 1301
rect 383 1265 397 1279
rect 1343 1265 1357 1279
rect 2999 1265 3013 1279
rect 3119 1265 3133 1279
rect 3479 1265 3493 1279
rect 3599 1265 3613 1279
rect 4775 1265 4789 1279
rect 5015 1265 5029 1279
rect 5111 1265 5125 1279
rect 5759 1265 5773 1279
rect 6743 1265 6757 1279
rect 263 1243 277 1257
rect 647 1243 661 1257
rect 983 1243 997 1257
rect 1559 1243 1573 1257
rect 3215 1243 3229 1257
rect 3335 1243 3349 1257
rect 3455 1243 3469 1257
rect 3575 1243 3589 1257
rect 6719 1243 6733 1257
rect 6935 1243 6949 1257
rect 7007 1243 7021 1257
rect 143 1221 157 1235
rect 791 1221 805 1235
rect 1223 1221 1237 1235
rect 2663 1221 2677 1235
rect 4751 1221 4765 1235
rect 4823 1221 4837 1235
rect 4870 1221 4884 1235
rect 5183 1221 5197 1235
rect 5255 1221 5269 1235
rect 5687 1221 5701 1235
rect 5879 1221 5893 1235
rect 5927 1221 5941 1235
rect 5975 1221 5989 1235
rect 6071 1221 6085 1235
rect 6119 1221 6133 1235
rect 6335 1221 6349 1235
rect 6455 1221 6469 1235
rect 6575 1221 6589 1235
rect 6791 1221 6805 1235
rect 6983 1221 6997 1235
rect 23 1199 37 1213
rect 1535 1199 1549 1213
rect 2543 1199 2557 1213
rect 2639 1199 2653 1213
rect 4895 1199 4909 1213
rect 5063 1199 5077 1213
rect 5231 1199 5245 1213
rect 5303 1199 5317 1213
rect 5351 1199 5365 1213
rect 5807 1199 5821 1213
rect 5855 1199 5869 1213
rect 7031 1199 7045 1213
rect 7079 1199 7093 1213
rect 7127 1199 7141 1213
rect 71 380 85 394
rect 623 380 637 394
rect 1247 380 1261 394
rect 5375 380 5389 394
rect 5999 380 6013 394
rect 7151 380 7165 394
rect 191 358 205 372
rect 2567 358 2581 372
rect 4991 358 5005 372
rect 6023 358 6037 372
rect 6695 358 6709 372
rect 6839 358 6853 372
rect 311 336 325 350
rect 767 336 781 350
rect 887 336 901 350
rect 1583 336 1597 350
rect 2735 336 2749 350
rect 2855 336 2869 350
rect 2975 336 2989 350
rect 3095 336 3109 350
rect 5399 336 5413 350
rect 5615 336 5629 350
rect 5735 336 5749 350
rect 6863 336 6877 350
rect 431 314 445 328
rect 2759 314 2773 328
rect 2879 314 2893 328
rect 3239 314 3253 328
rect 3359 314 3373 328
rect 3983 314 3997 328
rect 4079 314 4093 328
rect 4175 314 4189 328
rect 4271 314 4285 328
rect 4367 314 4381 328
rect 4463 314 4477 328
rect 4559 314 4573 328
rect 4655 314 4669 328
rect 4968 314 4982 328
rect 5447 314 5461 328
rect 6167 314 6181 328
rect 6215 314 6229 328
rect 551 292 565 306
rect 743 292 757 306
rect 2783 292 2797 306
rect 3023 292 3037 306
rect 3263 292 3277 306
rect 3503 292 3517 306
rect 5639 292 5653 306
rect 6887 291 6901 305
rect 167 270 181 284
rect 1487 270 1501 284
rect 1823 270 1837 284
rect 2183 270 2197 284
rect 2687 269 2701 283
rect 3695 269 3709 283
rect 3791 269 3805 283
rect 3887 269 3901 283
rect 5611 270 5625 284
rect 6287 270 6301 284
rect 1631 248 1645 262
rect 1703 248 1717 262
rect 2591 247 2605 261
rect 3983 247 3997 261
rect 4171 248 4185 262
rect 4319 248 4333 262
rect 5399 248 5413 262
rect 6407 248 6421 262
rect 196 225 210 239
rect 3743 225 3757 239
rect 3839 225 3853 239
rect 5519 225 5533 239
rect 5807 226 5821 240
rect 6527 226 6541 240
rect 335 203 349 217
rect 1919 203 1933 217
rect 2063 203 2077 217
rect 4171 203 4185 217
rect 4511 203 4525 217
rect 6695 203 6709 217
rect 503 181 517 195
rect 1991 181 2005 195
rect 2711 181 2725 195
rect 4607 181 4621 195
rect 6167 181 6181 195
rect 6647 181 6661 195
rect 527 159 541 173
rect 2207 159 2221 173
rect 3047 159 3061 173
rect 4703 159 4717 173
rect 6527 159 6541 173
rect 7199 159 7213 173
rect 599 137 613 151
rect 2375 137 2389 151
rect 3167 137 3181 151
rect 5495 137 5509 151
rect 815 115 829 129
rect 2423 115 2437 129
rect 3215 115 3229 129
rect 4415 115 4429 129
rect 959 93 973 107
rect 4943 93 4957 107
rect 1295 71 1309 85
rect 4031 71 4045 85
rect 4943 69 4957 83
rect 5611 69 5625 83
rect 1655 49 1669 63
rect 4127 49 4141 63
rect 2399 27 2413 41
rect 4223 27 4237 41
rect 3383 5 3397 19
rect 3935 5 3949 19
<< metal2 >>
rect 24 1213 36 1481
rect 144 1235 156 1481
rect 264 1257 276 1481
rect 384 1279 396 1481
rect 504 1301 516 1481
rect 24 1196 36 1199
rect 144 1196 156 1221
rect 264 1196 276 1243
rect 384 1196 396 1265
rect 504 1196 516 1287
rect 648 1196 660 1243
rect 672 1196 684 1287
rect 696 1196 708 1353
rect 792 1196 804 1221
rect 816 1196 828 1331
rect 864 1196 876 1287
rect 912 1196 924 1309
rect 960 1196 972 1309
rect 984 1196 996 1243
rect 1032 1196 1044 1309
rect 1080 1196 1092 1331
rect 1104 1196 1116 1353
rect 1152 1196 1164 1331
rect 1200 1196 1212 1309
rect 1224 1196 1236 1221
rect 1272 1196 1284 1309
rect 1320 1196 1332 1331
rect 1344 1196 1356 1265
rect 1368 1196 1380 1331
rect 1416 1196 1428 1309
rect 1440 1196 1452 1331
rect 1536 1196 1548 1199
rect 1560 1196 1572 1243
rect 1680 1196 1692 1481
rect 1752 1196 1764 1309
rect 1800 1196 1812 1309
rect 2016 1196 2028 1309
rect 2112 1196 2124 1481
rect 2304 1323 2316 1481
rect 2304 1196 2316 1309
rect 2376 1196 2388 1481
rect 2472 1196 2484 1481
rect 2544 1196 2556 1199
rect 2640 1196 2652 1199
rect 2664 1196 2676 1221
rect 2808 1196 2820 1375
rect 2904 1196 2916 1287
rect 2928 1196 2940 1397
rect 3000 1196 3012 1265
rect 3048 1196 3060 1309
rect 3120 1196 3132 1265
rect 3144 1196 3156 1287
rect 3168 1196 3180 1419
rect 3216 1196 3228 1243
rect 3288 1196 3300 1331
rect 3336 1196 3348 1243
rect 3384 1196 3396 1287
rect 3408 1196 3420 1440
rect 3456 1196 3468 1243
rect 3480 1196 3492 1265
rect 3528 1196 3540 1462
rect 3576 1196 3588 1243
rect 3600 1196 3612 1265
rect 3624 1196 3636 1287
rect 3648 1196 3660 1353
rect 3720 1196 3732 1309
rect 3816 1196 3828 1331
rect 3912 1196 3924 1353
rect 4008 1196 4020 1375
rect 4104 1196 4116 1396
rect 4200 1196 4212 1309
rect 4296 1196 4308 1418
rect 4392 1196 4404 1331
rect 4416 1196 4428 1309
rect 4488 1196 4500 1440
rect 4584 1196 4596 1462
rect 4680 1196 4692 1353
rect 4752 1196 4764 1221
rect 4776 1196 4788 1265
rect 4800 1196 4812 1287
rect 4824 1196 4836 1221
rect 4872 1196 4884 1221
rect 4896 1196 4908 1199
rect 5016 1196 5028 1265
rect 5064 1196 5076 1199
rect 5112 1196 5124 1265
rect 5136 1196 5148 1287
rect 5184 1196 5196 1221
rect 5232 1196 5244 1199
rect 5256 1196 5268 1221
rect 5304 1196 5316 1199
rect 5352 1196 5364 1199
rect 5688 1196 5700 1221
rect 5760 1196 5772 1265
rect 5808 1196 5820 1199
rect 5856 1196 5868 1199
rect 5880 1196 5892 1221
rect 5928 1196 5940 1221
rect 5976 1196 5988 1221
rect 6072 1196 6084 1221
rect 6120 1196 6132 1221
rect 6144 1196 6156 1481
rect 6240 1196 6252 1309
rect 6336 1196 6348 1221
rect 6360 1196 6372 1481
rect 6456 1196 6468 1221
rect 6480 1196 6492 1481
rect 6576 1196 6588 1221
rect 6600 1196 6612 1481
rect 6720 1196 6732 1243
rect 6744 1196 6756 1265
rect 6792 1196 6804 1221
rect 6936 1196 6948 1243
rect 6984 1196 6996 1221
rect 7008 1196 7020 1243
rect 7032 1196 7044 1199
rect 7080 1196 7092 1199
rect 7128 1196 7140 1199
rect 72 394 84 397
rect 192 372 204 397
rect 312 350 324 397
rect 432 328 444 397
rect 552 306 564 397
rect 624 394 636 397
rect 744 306 756 397
rect 768 350 780 397
rect 888 350 900 397
rect 1248 394 1260 397
rect 1488 284 1500 397
rect 1584 350 1596 397
rect 168 0 180 270
rect 1632 262 1644 397
rect 1704 262 1716 397
rect 1824 284 1836 397
rect 197 0 209 225
rect 1920 217 1932 397
rect 336 0 348 203
rect 1992 195 2004 397
rect 2184 284 2196 397
rect 504 0 516 181
rect 528 0 540 159
rect 600 0 612 137
rect 816 0 828 115
rect 960 0 972 93
rect 1296 0 1308 71
rect 1656 0 1668 49
rect 2064 0 2076 203
rect 2208 173 2220 397
rect 2376 151 2388 397
rect 2424 129 2436 397
rect 2568 372 2580 397
rect 2592 261 2604 397
rect 2688 283 2700 397
rect 2736 350 2748 397
rect 2760 328 2772 397
rect 2784 306 2796 397
rect 2856 350 2868 397
rect 2880 328 2892 397
rect 2976 350 2988 397
rect 3024 306 3036 397
rect 3096 350 3108 397
rect 3240 328 3252 397
rect 3264 306 3276 397
rect 3360 328 3372 397
rect 3504 306 3516 397
rect 3696 283 3708 397
rect 3744 239 3756 397
rect 3792 283 3804 397
rect 3840 239 3852 397
rect 3888 283 3900 397
rect 2400 0 2412 27
rect 2712 0 2724 181
rect 3048 0 3060 159
rect 3168 0 3180 137
rect 3216 0 3228 115
rect 3936 19 3948 397
rect 3984 328 3996 397
rect 3984 261 3996 314
rect 4032 85 4044 397
rect 4080 328 4092 397
rect 4128 63 4140 397
rect 4176 328 4188 397
rect 4172 217 4184 248
rect 4224 41 4236 397
rect 4272 328 4284 397
rect 4320 262 4332 397
rect 4368 328 4380 397
rect 4416 129 4428 397
rect 4464 328 4476 397
rect 4512 217 4524 397
rect 4560 328 4572 397
rect 4608 195 4620 397
rect 4656 328 4668 397
rect 4704 173 4716 397
rect 4944 107 4956 397
rect 4992 372 5004 397
rect 5376 394 5388 397
rect 5400 350 5412 397
rect 5448 328 5460 397
rect 3384 0 3396 5
rect 4944 0 4956 69
rect 4969 0 4981 314
rect 5400 0 5412 248
rect 5496 151 5508 397
rect 5520 239 5532 397
rect 5568 0 5580 397
rect 5616 350 5628 397
rect 5640 306 5652 397
rect 5736 350 5748 397
rect 6000 394 6012 397
rect 6024 372 6036 397
rect 6168 328 6180 397
rect 6216 328 6228 397
rect 6288 284 6300 397
rect 5612 83 5624 270
rect 6408 262 6420 397
rect 6528 240 6540 397
rect 5808 0 5820 226
rect 6648 195 6660 397
rect 6696 372 6708 397
rect 6840 372 6852 397
rect 6864 350 6876 397
rect 6888 305 6900 397
rect 7152 394 7164 397
rect 6168 0 6180 181
rect 6528 0 6540 159
rect 6696 0 6708 203
rect 7200 173 7212 397
use inv inv_0
timestamp 1386238110
transform 1 0 0 0 1 397
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 120 0 1 397
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 240 0 1 397
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 360 0 1 397
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 480 0 1 397
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 600 0 1 397
box 0 0 120 799
use nand3 nand3_1
timestamp 1386234893
transform 1 0 720 0 1 397
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 840 0 1 397
box 0 0 96 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 936 0 1 397
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 1056 0 1 397
box 0 0 120 799
use nand3 nand3_2
timestamp 1386234893
transform 1 0 1176 0 1 397
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1296 0 1 397
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 1392 0 1 397
box 0 0 120 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 1512 0 1 397
box 0 0 144 799
use and2 and2_4
timestamp 1386234845
transform 1 0 1656 0 1 397
box 0 0 120 799
use xor2 xor2_3
timestamp 1386237344
transform 1 0 1776 0 1 397
box 0 0 192 799
use xor2 xor2_4
timestamp 1386237344
transform 1 0 1968 0 1 397
box 0 0 192 799
use xor2 xor2_5
timestamp 1386237344
transform 1 0 2160 0 1 397
box 0 0 192 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 2352 0 1 397
box 0 0 48 799
use inv inv_6
timestamp 1386238110
transform 1 0 2400 0 1 397
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 2520 0 1 397
box 0 0 96 799
use nand2 nand2_3
timestamp 1386234792
transform 1 0 2616 0 1 397
box 0 0 96 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 2712 0 1 397
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 2832 0 1 397
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 2952 0 1 397
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 3072 0 1 397
box 0 0 120 799
use nand3 nand3_8
timestamp 1386234893
transform 1 0 3192 0 1 397
box 0 0 120 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 3312 0 1 397
box 0 0 120 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 3432 0 1 397
box 0 0 120 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 3552 0 1 397
box 0 0 120 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 3672 0 1 397
box 0 0 96 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 3768 0 1 397
box 0 0 96 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 3864 0 1 397
box 0 0 96 799
use nand2 nand2_7
timestamp 1386234792
transform 1 0 3960 0 1 397
box 0 0 96 799
use nand2 nand2_8
timestamp 1386234792
transform 1 0 4056 0 1 397
box 0 0 96 799
use nand2 nand2_9
timestamp 1386234792
transform 1 0 4152 0 1 397
box 0 0 96 799
use nand2 nand2_10
timestamp 1386234792
transform 1 0 4248 0 1 397
box 0 0 96 799
use nand2 nand2_11
timestamp 1386234792
transform 1 0 4344 0 1 397
box 0 0 96 799
use nand2 nand2_12
timestamp 1386234792
transform 1 0 4440 0 1 397
box 0 0 96 799
use nand2 nand2_13
timestamp 1386234792
transform 1 0 4536 0 1 397
box 0 0 96 799
use nand2 nand2_14
timestamp 1386234792
transform 1 0 4632 0 1 397
box 0 0 96 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 4728 0 1 397
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 4848 0 1 397
box 0 0 120 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 4968 0 1 397
box 0 0 120 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 5088 0 1 397
box 0 0 120 799
use nor2 nor2_6
timestamp 1386235306
transform 1 0 5208 0 1 397
box 0 0 120 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 5328 0 1 397
box 0 0 144 799
use and2 and2_3
timestamp 1386234845
transform 1 0 5472 0 1 397
box 0 0 120 799
use nor2 nor2_7
timestamp 1386235306
transform 1 0 5592 0 1 397
box 0 0 120 799
use nor2 nor2_8
timestamp 1386235306
transform 1 0 5712 0 1 397
box 0 0 120 799
use nor2 nor2_9
timestamp 1386235306
transform 1 0 5832 0 1 397
box 0 0 120 799
use nor3 nor3_2
timestamp 1386235396
transform 1 0 5952 0 1 397
box 0 0 144 799
use nand2 nand2_15
timestamp 1386234792
transform 1 0 6096 0 1 397
box 0 0 96 799
use nor2 nor2_10
timestamp 1386235306
transform 1 0 6192 0 1 397
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 6312 0 1 397
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 6432 0 1 397
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 6552 0 1 397
box 0 0 120 799
use nor3 nor3_3
timestamp 1386235396
transform 1 0 6672 0 1 397
box 0 0 144 799
use nor3 nor3_4
timestamp 1386235396
transform 1 0 6816 0 1 397
box 0 0 144 799
use nor3 nor3_5
timestamp 1386235396
transform 1 0 6960 0 1 397
box 0 0 144 799
use nor2 nor2_11
timestamp 1386235306
transform 1 0 7104 0 1 397
box 0 0 120 799
<< labels >>
rlabel metal1 336 344 336 344 1 nC
rlabel metal1 579 297 579 297 1 nE
rlabel metal1 104 386 104 386 1 nA
rlabel metal1 210 364 210 364 1 nB
rlabel metal1 459 319 459 319 1 nD
rlabel metal2 24 1481 36 1481 5 OpCode[4]
rlabel metal2 144 1481 156 1481 5 OpCode[3]
rlabel metal2 264 1481 276 1481 5 OpCode[2]
rlabel metal2 384 1481 396 1481 5 OpCode[1]
rlabel metal2 504 1481 516 1481 5 OpCode[0]
rlabel metal2 2472 1481 2484 1481 5 Z
rlabel metal2 2376 1481 2388 1481 5 N
rlabel metal2 2112 1481 2124 1481 5 V
rlabel metal2 1680 1481 1692 1481 5 Cin
rlabel metal2 2304 1481 2316 1481 5 C
rlabel metal2 6600 1481 6612 1481 5 imm4[0]
rlabel metal2 6480 1481 6492 1481 5 imm4[1]
rlabel metal2 6360 1481 6372 1481 5 imm4[2]
rlabel metal2 6144 1481 6156 1481 5 imm4[3]
rlabel metal2 6077 1198 6077 1198 1 N
rlabel metal1 5334 231 5334 231 1 ShSign
rlabel metal2 5568 0 5580 0 1 ShInBit
rlabel metal2 2712 0 2724 0 1 NAND
rlabel metal2 168 0 180 0 1 SUB
rlabel metal2 197 0 209 0 1 ZeroA
rlabel metal2 336 0 348 0 1 CIn_slice
rlabel metal2 504 0 516 0 1 LastCIn
rlabel metal2 528 0 540 0 1 COut
rlabel metal2 600 0 612 0 1 N
rlabel metal2 816 0 828 0 1 nZ
rlabel metal2 960 0 972 0 1 FAOut
rlabel metal2 1296 0 1308 0 1 AND
rlabel metal2 1656 0 1668 0 1 OR
rlabel metal2 2064 0 2076 0 1 XOR
rlabel metal2 2400 0 2412 0 1 NOT
rlabel metal2 3384 0 3396 0 1 ShL
rlabel metal2 4969 0 4981 0 1 ShR
rlabel metal2 6528 0 6540 0 1 ShOut
rlabel metal2 3168 0 3180 0 1 ASign
rlabel metal2 3216 0 3228 0 1 ShB
rlabel metal2 4944 0 4956 0 1 Sh8
rlabel metal2 5400 0 5412 0 1 Sh4
rlabel metal2 5808 0 5820 0 1 Sh2
rlabel metal2 6168 0 6180 0 1 Sh1
rlabel metal2 3048 0 3060 0 1 NOR
rlabel metal2 6696 0 6708 0 1 LLI
<< end >>
