magic
tech c035u
timestamp 1394479763
<< checkpaint >>
rect 6212 -435 8824 2342
<< metal1 >>
rect 4693 1025 6455 1035
rect 4237 1003 5999 1013
rect 3589 981 5351 991
rect 5390 980 5975 990
rect 5989 980 6431 990
rect 6445 981 6791 991
rect 3565 958 4199 968
rect 4213 958 4655 968
rect 4669 958 5015 968
rect 5053 959 6815 969
rect 445 936 647 946
rect 709 938 839 948
rect 3637 936 4031 946
rect 4285 936 4487 946
rect 4741 936 4847 946
rect 5413 936 5807 946
rect 6061 936 6263 946
rect 6517 937 6623 947
rect 6877 936 6935 946
rect 277 914 575 924
rect 685 914 695 924
rect 781 913 911 923
rect 925 914 1055 924
rect 1357 914 1391 924
rect 1693 914 1751 924
rect 2101 914 2159 924
rect 2437 914 2495 924
rect 2773 914 2807 924
rect 3109 914 3143 924
rect 3685 914 3695 924
rect 3733 914 3743 924
rect 3781 914 3791 924
rect 3829 914 3839 924
rect 3877 914 3887 924
rect 3925 914 3935 924
rect 3973 914 3983 924
rect 4333 914 4343 924
rect 4381 914 4391 924
rect 4429 914 4439 924
rect 4789 914 4799 924
rect 5101 917 5159 927
rect 5341 914 5375 924
rect 5437 914 5447 924
rect 5485 914 5495 924
rect 5533 914 5543 924
rect 5581 914 5591 924
rect 5629 914 5639 924
rect 5677 914 5687 924
rect 5725 914 5735 924
rect 5773 914 5879 924
rect 6085 914 6095 924
rect 6133 914 6143 924
rect 6181 914 6191 924
rect 6229 914 6335 924
rect 6541 915 6551 925
rect 6589 914 6695 924
rect 6901 914 7007 924
rect 0 892 311 902
rect 325 892 1295 902
rect 1309 892 1631 902
rect 1645 892 1991 902
rect 2005 892 2735 902
rect 2749 892 3047 902
rect 3061 892 3455 902
rect 3469 892 7296 902
rect 0 870 191 880
rect 205 870 1271 880
rect 1285 870 1607 880
rect 1621 870 1967 880
rect 1981 870 2375 880
rect 2389 870 2711 880
rect 2725 870 3023 880
rect 3037 870 3335 880
rect 3349 870 3407 880
rect 3493 870 3647 880
rect 3661 870 4055 880
rect 4141 870 4295 880
rect 4309 870 4511 880
rect 4597 870 4751 880
rect 4765 870 4871 880
rect 4957 870 5183 880
rect 5269 870 5831 880
rect 5917 870 6287 880
rect 6374 870 6647 880
rect 6733 870 6959 880
rect 7045 870 7103 880
rect 133 51 215 61
rect 949 44 983 54
rect 1213 51 1535 61
rect 1549 51 1895 61
rect 1909 51 2303 61
rect 2317 51 2639 61
rect 2653 51 2951 61
rect 2965 51 3287 61
rect 3301 51 7247 61
rect 7261 51 7296 61
rect 7488 51 7511 61
rect 7669 51 7704 61
rect 3661 29 3671 39
rect 3709 29 3719 39
rect 3757 29 3767 39
rect 3805 29 3815 39
rect 3853 29 3863 39
rect 3901 29 3911 39
rect 3949 29 3959 39
rect 3997 29 4103 39
rect 4309 29 4319 39
rect 4357 29 4367 39
rect 4405 29 4415 39
rect 4453 29 4559 39
rect 4765 29 4775 39
rect 4813 29 4919 39
rect 5197 29 5231 39
rect 5341 29 5376 39
rect 5461 29 5471 39
rect 5509 29 5519 39
rect 5557 29 5567 39
rect 5605 29 5615 39
rect 5653 29 5663 39
rect 5701 29 5711 39
rect 5749 29 5759 39
rect 6109 29 6119 39
rect 6157 29 6167 39
rect 6205 29 6215 39
rect 6565 29 6575 39
rect 6901 29 6959 39
rect 5437 7 5831 17
rect 6085 7 6287 17
rect 6541 7 6647 17
<< m2contact >>
rect 4679 1023 4693 1037
rect 6455 1023 6469 1037
rect 4223 1001 4237 1015
rect 5999 1001 6013 1015
rect 3575 978 3589 992
rect 5351 979 5365 993
rect 5376 979 5390 993
rect 5975 979 5989 993
rect 6431 979 6445 993
rect 6791 979 6805 993
rect 3551 956 3565 970
rect 4199 956 4213 970
rect 4655 956 4669 970
rect 5015 956 5029 970
rect 5039 956 5053 970
rect 6815 957 6829 971
rect 431 935 445 949
rect 647 934 661 948
rect 695 936 709 950
rect 839 936 853 950
rect 3623 934 3637 948
rect 4031 934 4045 948
rect 4271 934 4285 948
rect 4487 934 4501 948
rect 4727 934 4741 948
rect 4847 934 4861 948
rect 5399 934 5413 948
rect 5807 934 5821 948
rect 6047 934 6061 948
rect 6263 934 6277 948
rect 6503 935 6517 949
rect 6623 935 6637 949
rect 6863 934 6877 948
rect 6935 934 6949 948
rect 263 912 277 926
rect 575 912 589 926
rect 671 912 685 926
rect 695 912 709 926
rect 767 912 781 926
rect 911 912 925 926
rect 1055 912 1069 926
rect 1343 912 1357 926
rect 1391 912 1405 926
rect 1679 912 1693 926
rect 1751 912 1765 926
rect 2087 912 2101 926
rect 2159 912 2173 926
rect 2423 912 2437 926
rect 2495 912 2509 926
rect 2759 912 2773 926
rect 2807 912 2821 926
rect 3095 912 3109 926
rect 3143 912 3157 926
rect 3671 912 3685 926
rect 3695 912 3709 926
rect 3719 912 3733 926
rect 3743 912 3757 926
rect 3767 912 3781 926
rect 3791 912 3805 926
rect 3815 912 3829 926
rect 3839 912 3853 926
rect 3863 912 3877 926
rect 3887 912 3901 926
rect 3911 912 3925 926
rect 3935 912 3949 926
rect 3959 912 3973 926
rect 3983 912 3997 926
rect 4319 912 4333 926
rect 4343 912 4357 926
rect 4367 912 4381 926
rect 4391 912 4405 926
rect 4415 912 4429 926
rect 4439 912 4453 926
rect 4775 912 4789 926
rect 4799 912 4813 926
rect 5087 916 5101 930
rect 5159 916 5173 930
rect 5327 912 5341 926
rect 5375 912 5389 926
rect 5423 912 5437 926
rect 5447 912 5461 926
rect 5471 912 5485 926
rect 5495 912 5509 926
rect 5519 912 5533 926
rect 5543 912 5557 926
rect 5567 912 5581 926
rect 5591 912 5605 926
rect 5615 912 5629 926
rect 5639 912 5653 926
rect 5663 912 5677 926
rect 5687 912 5701 926
rect 5711 912 5725 926
rect 5735 912 5749 926
rect 5759 912 5773 926
rect 5879 912 5893 926
rect 6071 912 6085 926
rect 6095 912 6109 926
rect 6119 912 6133 926
rect 6143 912 6157 926
rect 6167 912 6181 926
rect 6191 912 6205 926
rect 6215 912 6229 926
rect 6335 912 6349 926
rect 6527 913 6541 927
rect 6551 913 6565 927
rect 6575 913 6589 927
rect 6695 912 6709 926
rect 6887 912 6901 926
rect 7007 912 7021 926
rect 311 890 325 904
rect 1295 890 1309 904
rect 1631 890 1645 904
rect 1991 890 2005 904
rect 2735 890 2749 904
rect 3047 890 3061 904
rect 3455 890 3469 904
rect 191 868 205 882
rect 1271 868 1285 882
rect 1607 868 1621 882
rect 1967 868 1981 882
rect 2375 868 2389 882
rect 2711 868 2725 882
rect 3023 868 3037 882
rect 3335 868 3349 882
rect 3407 868 3421 882
rect 3479 868 3493 882
rect 3647 868 3661 882
rect 4055 868 4069 882
rect 4127 868 4141 882
rect 4295 868 4309 882
rect 4511 868 4525 882
rect 4583 868 4597 882
rect 4751 868 4765 882
rect 4871 868 4885 882
rect 4943 868 4957 882
rect 5183 868 5197 882
rect 5255 868 5269 882
rect 5831 868 5845 882
rect 5903 868 5917 882
rect 6287 868 6301 882
rect 6360 868 6374 882
rect 6647 868 6661 882
rect 6719 868 6733 882
rect 6959 868 6973 882
rect 7031 868 7045 882
rect 7103 868 7117 882
rect 119 49 133 63
rect 215 49 229 63
rect 935 42 949 56
rect 983 42 997 56
rect 1199 49 1213 63
rect 1535 49 1549 63
rect 1895 49 1909 63
rect 2303 49 2317 63
rect 2639 49 2653 63
rect 2951 49 2965 63
rect 3287 49 3301 63
rect 7247 49 7261 63
rect 7511 49 7525 63
rect 7655 49 7669 63
rect 3647 27 3661 41
rect 3671 27 3685 41
rect 3695 27 3709 41
rect 3719 27 3733 41
rect 3743 27 3757 41
rect 3767 27 3781 41
rect 3791 27 3805 41
rect 3815 27 3829 41
rect 3839 27 3853 41
rect 3863 27 3877 41
rect 3887 27 3901 41
rect 3911 27 3925 41
rect 3935 27 3949 41
rect 3959 27 3973 41
rect 3983 27 3997 41
rect 4103 27 4117 41
rect 4295 27 4309 41
rect 4319 27 4333 41
rect 4343 27 4357 41
rect 4367 27 4381 41
rect 4391 27 4405 41
rect 4415 27 4429 41
rect 4439 27 4453 41
rect 4559 27 4573 41
rect 4751 27 4765 41
rect 4775 27 4789 41
rect 4799 27 4813 41
rect 4919 27 4933 41
rect 5183 27 5197 41
rect 5231 27 5245 41
rect 5327 27 5341 41
rect 5376 27 5390 41
rect 5447 27 5461 41
rect 5471 27 5485 41
rect 5495 27 5509 41
rect 5519 27 5533 41
rect 5543 27 5557 41
rect 5567 27 5581 41
rect 5591 27 5605 41
rect 5615 27 5629 41
rect 5639 27 5653 41
rect 5663 27 5677 41
rect 5687 27 5701 41
rect 5711 27 5725 41
rect 5735 27 5749 41
rect 5759 27 5773 41
rect 6095 27 6109 41
rect 6119 27 6133 41
rect 6143 27 6157 41
rect 6167 27 6181 41
rect 6191 27 6205 41
rect 6215 27 6229 41
rect 6551 27 6565 41
rect 6575 27 6589 41
rect 6887 27 6901 41
rect 6959 27 6973 41
rect 5423 5 5437 19
rect 5831 5 5845 19
rect 6071 5 6085 19
rect 6287 5 6301 19
rect 6527 5 6541 19
rect 6647 5 6661 19
<< metal2 >>
rect 72 865 84 1042
rect 192 865 204 868
rect 264 865 276 912
rect 312 865 324 890
rect 336 865 348 1042
rect 432 865 444 935
rect 504 865 516 1042
rect 576 865 588 912
rect 648 865 660 934
rect 672 926 684 1042
rect 696 950 708 1042
rect 768 926 780 1042
rect 696 865 708 912
rect 768 865 780 912
rect 840 865 852 936
rect 912 865 924 912
rect 984 865 996 1042
rect 1056 865 1068 912
rect 1128 865 1140 1042
rect 1272 865 1284 868
rect 1296 865 1308 890
rect 1344 865 1356 912
rect 1392 865 1404 912
rect 1464 865 1476 1042
rect 1608 865 1620 868
rect 1632 865 1644 890
rect 1680 865 1692 912
rect 1752 865 1764 912
rect 1824 865 1836 1042
rect 1968 865 1980 868
rect 1992 865 2004 890
rect 2088 865 2100 912
rect 2160 865 2172 912
rect 2232 865 2244 1042
rect 2376 865 2388 868
rect 2424 865 2436 912
rect 2496 865 2508 912
rect 2568 865 2580 1042
rect 2712 865 2724 868
rect 2736 865 2748 890
rect 2760 865 2772 912
rect 2808 865 2820 912
rect 2880 865 2892 1042
rect 3024 865 3036 868
rect 3048 865 3060 890
rect 3096 865 3108 912
rect 3144 865 3156 912
rect 3216 865 3228 1042
rect 3336 882 3348 1042
rect 3384 865 3396 1042
rect 3552 970 3564 1042
rect 3408 865 3420 868
rect 3456 865 3468 890
rect 3480 865 3492 868
rect 3552 865 3564 956
rect 3576 865 3588 978
rect 3624 865 3636 934
rect 3648 882 3660 1042
rect 3696 926 3708 1042
rect 3744 926 3756 1042
rect 3792 926 3804 1042
rect 3840 926 3852 1042
rect 3888 926 3900 1042
rect 3936 926 3948 1042
rect 3984 926 3996 1042
rect 3672 865 3684 912
rect 3720 865 3732 912
rect 3768 865 3780 912
rect 3816 865 3828 912
rect 3864 865 3876 912
rect 3912 865 3924 912
rect 3960 865 3972 912
rect 4032 865 4044 934
rect 4056 865 4068 868
rect 4128 865 4140 868
rect 4200 865 4212 956
rect 4224 865 4236 1001
rect 4272 865 4284 934
rect 4296 882 4308 1042
rect 4344 926 4356 1042
rect 4392 926 4404 1042
rect 4440 926 4452 1042
rect 4320 865 4332 912
rect 4368 865 4380 912
rect 4416 865 4428 912
rect 4488 865 4500 934
rect 4512 865 4524 868
rect 4584 865 4596 868
rect 4656 865 4668 956
rect 4680 865 4692 1023
rect 4728 865 4740 934
rect 4752 882 4764 1042
rect 4800 926 4812 1042
rect 4776 865 4788 912
rect 4848 865 4860 934
rect 4872 865 4884 868
rect 4944 865 4956 868
rect 5016 865 5028 956
rect 5040 865 5052 956
rect 5088 865 5100 916
rect 5160 865 5172 916
rect 5184 882 5196 1042
rect 5352 993 5364 1042
rect 5377 993 5389 1042
rect 5184 865 5196 868
rect 5256 865 5268 868
rect 5328 865 5340 912
rect 5352 865 5364 979
rect 5377 926 5389 979
rect 5400 865 5412 934
rect 5424 926 5436 1042
rect 5472 926 5484 1042
rect 5520 926 5532 1042
rect 5568 926 5580 1042
rect 5616 926 5628 1042
rect 5664 926 5676 1042
rect 5712 926 5724 1042
rect 5760 926 5772 1042
rect 6000 1015 6012 1042
rect 5448 865 5460 912
rect 5496 865 5508 912
rect 5544 865 5556 912
rect 5592 865 5604 912
rect 5640 865 5652 912
rect 5688 865 5700 912
rect 5736 865 5748 912
rect 5808 865 5820 934
rect 5832 865 5844 868
rect 5880 865 5892 912
rect 5904 865 5916 868
rect 5976 865 5988 979
rect 6000 865 6012 1001
rect 6048 865 6060 934
rect 6072 926 6084 1042
rect 6120 926 6132 1042
rect 6168 926 6180 1042
rect 6216 926 6228 1042
rect 6456 1037 6468 1042
rect 6096 865 6108 912
rect 6144 865 6156 912
rect 6192 865 6204 912
rect 6264 865 6276 934
rect 6288 865 6300 868
rect 6336 865 6348 912
rect 6360 865 6372 868
rect 6432 865 6444 979
rect 6456 865 6468 1023
rect 6504 865 6516 935
rect 6528 927 6540 1042
rect 6576 927 6588 1042
rect 6552 865 6564 913
rect 6624 865 6636 935
rect 6648 865 6660 868
rect 6696 865 6708 912
rect 6720 865 6732 868
rect 6792 865 6804 979
rect 6816 971 6828 1042
rect 6816 865 6828 957
rect 6864 865 6876 934
rect 6888 926 6900 1042
rect 6936 865 6948 934
rect 6960 865 6972 868
rect 7008 865 7020 912
rect 7032 865 7044 868
rect 7104 865 7116 868
rect 7176 865 7188 1042
rect 7512 865 7524 1042
rect 7584 865 7596 1042
rect 24 0 36 66
rect 72 0 84 66
rect 120 63 132 66
rect 216 63 228 66
rect 336 0 348 66
rect 504 0 516 66
rect 696 0 708 66
rect 936 56 948 66
rect 984 0 996 42
rect 1128 0 1140 66
rect 1200 63 1212 66
rect 1464 0 1476 66
rect 1536 63 1548 66
rect 1824 0 1836 66
rect 1896 63 1908 66
rect 2232 0 2244 66
rect 2304 63 2316 66
rect 2568 0 2580 66
rect 2640 63 2652 66
rect 2880 0 2892 66
rect 2952 63 2964 66
rect 3216 0 3228 66
rect 3288 63 3300 66
rect 3384 0 3396 66
rect 3552 0 3564 66
rect 3672 41 3684 66
rect 3720 41 3732 66
rect 3768 41 3780 66
rect 3816 41 3828 66
rect 3864 41 3876 66
rect 3912 41 3924 66
rect 3960 41 3972 66
rect 4104 41 4116 66
rect 4320 41 4332 66
rect 4368 41 4380 66
rect 4416 41 4428 66
rect 4560 41 4572 66
rect 4776 41 4788 66
rect 4920 41 4932 66
rect 5232 41 5244 66
rect 5328 41 5340 66
rect 3648 0 3660 27
rect 3696 0 3708 27
rect 3744 0 3756 27
rect 3792 0 3804 27
rect 3840 0 3852 27
rect 3888 0 3900 27
rect 3936 0 3948 27
rect 3984 0 3996 27
rect 4296 0 4308 27
rect 4344 0 4356 27
rect 4392 0 4404 27
rect 4440 0 4452 27
rect 4752 0 4764 27
rect 4800 0 4812 27
rect 5184 0 5196 27
rect 5352 0 5364 66
rect 5448 41 5460 66
rect 5496 41 5508 66
rect 5544 41 5556 66
rect 5592 41 5604 66
rect 5640 41 5652 66
rect 5688 41 5700 66
rect 5736 41 5748 66
rect 5377 0 5389 27
rect 5424 0 5436 5
rect 5472 0 5484 27
rect 5520 0 5532 27
rect 5568 0 5580 27
rect 5616 0 5628 27
rect 5664 0 5676 27
rect 5712 0 5724 27
rect 5760 0 5772 27
rect 5832 19 5844 66
rect 6000 0 6012 66
rect 6096 41 6108 66
rect 6144 41 6156 66
rect 6192 41 6204 66
rect 6072 0 6084 5
rect 6120 0 6132 27
rect 6168 0 6180 27
rect 6216 0 6228 27
rect 6288 19 6300 66
rect 6456 0 6468 66
rect 6552 41 6564 66
rect 6528 0 6540 5
rect 6576 0 6588 27
rect 6648 19 6660 66
rect 6816 0 6828 66
rect 6960 41 6972 66
rect 6888 0 6900 27
rect 7176 0 7188 66
rect 7248 63 7260 66
rect 7512 63 7524 66
rect 7584 0 7596 66
rect 7656 63 7668 66
use tielow  tielow_0
timestamp 1386086605
transform 1 0 0 0 1 66
box 0 0 48 799
use inv  inv_1
timestamp 1386238110
transform 1 0 48 0 1 66
box 0 0 120 799
use and2  and2_0
timestamp 1386234845
transform 1 0 168 0 1 66
box 0 0 120 799
use xor2  xor2_0
timestamp 1386237344
transform 1 0 288 0 1 66
box 0 0 192 799
use rowcrosser  rowcrosser_0
timestamp 1386086759
transform 1 0 480 0 1 66
box 0 0 48 799
use fulladder  fulladder_0
timestamp 1386234928
transform 1 0 528 0 1 66
box 0 0 360 799
use or2  or2_0
timestamp 1386235472
transform 1 0 888 0 1 66
box 0 0 144 799
use trisbuf  trisbuf_0
timestamp 1386237216
transform 1 0 1032 0 1 66
box 0 0 216 799
use and2  and2_1
timestamp 1386234845
transform 1 0 1248 0 1 66
box 0 0 120 799
use trisbuf  trisbuf_1
timestamp 1386237216
transform 1 0 1368 0 1 66
box 0 0 216 799
use or2  or2_1
timestamp 1386235472
transform 1 0 1584 0 1 66
box 0 0 144 799
use trisbuf  trisbuf_2
timestamp 1386237216
transform 1 0 1728 0 1 66
box 0 0 216 799
use xor2  xor2_1
timestamp 1386237344
transform 1 0 1944 0 1 66
box 0 0 192 799
use trisbuf  trisbuf_3
timestamp 1386237216
transform 1 0 2136 0 1 66
box 0 0 216 799
use inv  inv_0
timestamp 1386238110
transform 1 0 2352 0 1 66
box 0 0 120 799
use trisbuf  trisbuf_4
timestamp 1386237216
transform 1 0 2472 0 1 66
box 0 0 216 799
use nand2  nand2_0
timestamp 1386234792
transform 1 0 2688 0 1 66
box 0 0 96 799
use trisbuf  trisbuf_5
timestamp 1386237216
transform 1 0 2784 0 1 66
box 0 0 216 799
use nor2  nor2_0
timestamp 1386235306
transform 1 0 3000 0 1 66
box 0 0 120 799
use trisbuf  trisbuf_6
timestamp 1386237216
transform 1 0 3120 0 1 66
box 0 0 216 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 3336 0 1 66
box 0 0 192 799
use and2  and2_2
timestamp 1386234845
transform 1 0 3528 0 1 66
box 0 0 120 799
use rowcrosser  rowcrosser_1
timestamp 1386086759
transform 1 0 3648 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_2
timestamp 1386086759
transform 1 0 3696 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_3
timestamp 1386086759
transform 1 0 3744 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_14
timestamp 1386086759
transform 1 0 3792 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_16
timestamp 1386086759
transform 1 0 3840 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_17
timestamp 1386086759
transform 1 0 3888 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_18
timestamp 1386086759
transform 1 0 3936 0 1 66
box 0 0 48 799
use mux2  mux2_1
timestamp 1386235218
transform 1 0 3984 0 1 66
box 0 0 192 799
use and2  and2_3
timestamp 1386234845
transform 1 0 4176 0 1 66
box 0 0 120 799
use rowcrosser  rowcrosser_13
timestamp 1386086759
transform 1 0 4296 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_7
timestamp 1386086759
transform 1 0 4344 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_10
timestamp 1386086759
transform 1 0 4392 0 1 66
box 0 0 48 799
use mux2  mux2_4
timestamp 1386235218
transform 1 0 4440 0 1 66
box 0 0 192 799
use and2  and2_4
timestamp 1386234845
transform 1 0 4632 0 1 66
box 0 0 120 799
use rowcrosser  rowcrosser_9
timestamp 1386086759
transform 1 0 4752 0 1 66
box 0 0 48 799
use mux2  mux2_3
timestamp 1386235218
transform 1 0 4800 0 1 66
box 0 0 192 799
use and2  and2_5
timestamp 1386234845
transform 1 0 4992 0 1 66
box 0 0 120 799
use mux2  mux2_5
timestamp 1386235218
transform 1 0 5112 0 1 66
box 0 0 192 799
use and2  and2_6
timestamp 1386234845
transform 1 0 5304 0 1 66
box 0 0 120 799
use rowcrosser  rowcrosser_4
timestamp 1386086759
transform 1 0 5424 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_5
timestamp 1386086759
transform 1 0 5472 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_6
timestamp 1386086759
transform 1 0 5520 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_19
timestamp 1386086759
transform 1 0 5568 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_20
timestamp 1386086759
transform 1 0 5616 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_21
timestamp 1386086759
transform 1 0 5664 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_22
timestamp 1386086759
transform 1 0 5712 0 1 66
box 0 0 48 799
use mux2  mux2_2
timestamp 1386235218
transform 1 0 5760 0 1 66
box 0 0 192 799
use and2  and2_7
timestamp 1386234845
transform 1 0 5952 0 1 66
box 0 0 120 799
use rowcrosser  rowcrosser_8
timestamp 1386086759
transform 1 0 6072 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_11
timestamp 1386086759
transform 1 0 6120 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_12
timestamp 1386086759
transform 1 0 6168 0 1 66
box 0 0 48 799
use mux2  mux2_6
timestamp 1386235218
transform 1 0 6216 0 1 66
box 0 0 192 799
use and2  and2_8
timestamp 1386234845
transform 1 0 6408 0 1 66
box 0 0 120 799
use rowcrosser  rowcrosser_15
timestamp 1386086759
transform 1 0 6528 0 1 66
box 0 0 48 799
use mux2  mux2_7
timestamp 1386235218
transform 1 0 6576 0 1 66
box 0 0 192 799
use and2  and2_9
timestamp 1386234845
transform 1 0 6768 0 1 66
box 0 0 120 799
use mux2  mux2_8
timestamp 1386235218
transform 1 0 6888 0 1 66
box 0 0 192 799
use trisbuf  trisbuf_7
timestamp 1386237216
transform 1 0 7080 0 1 66
box 0 0 216 799
use trisbuf  trisbuf_8
timestamp 1386237216
transform 1 0 7488 0 1 66
box 0 0 216 799
<< labels >>
rlabel metal2 696 0 708 0 1 CIn_Slice
rlabel metal2 672 1042 684 1042 5 CIn_Slice
rlabel metal2 984 0 996 0 1 nZ_prev
rlabel metal2 336 0 348 0 1 SUB
rlabel metal2 3384 0 3396 0 1 ShB
rlabel metal2 3552 0 3564 0 1 ShL
rlabel metal2 3216 0 3228 0 1 NOR
rlabel metal2 2880 0 2892 0 1 NAND
rlabel metal2 2568 0 2580 0 1 NOT
rlabel metal2 2232 0 2244 0 1 XOR
rlabel metal2 1824 0 1836 0 1 OR
rlabel metal2 1464 0 1476 0 1 AND
rlabel metal2 504 0 516 0 1 CIn
rlabel metal2 1128 0 1140 0 1 FAOut
rlabel metal2 3552 1042 3564 1042 5 ShL
rlabel metal2 3648 1042 3660 1042 5 Sh8A_L
rlabel metal2 3744 1042 3756 1042 5 Sh8C_L
rlabel metal2 1128 1042 1140 1042 5 FAOut
rlabel metal2 984 1042 996 1042 5 nZ
rlabel metal2 336 1042 348 1042 5 SUB
rlabel metal2 1464 1042 1476 1042 5 AND
rlabel metal2 1824 1042 1836 1042 5 OR
rlabel metal2 2232 1042 2244 1042 5 XOR
rlabel metal2 2568 1042 2580 1042 5 NOT
rlabel metal2 2880 1042 2892 1042 5 NAND
rlabel metal2 3216 1042 3228 1042 5 NOR
rlabel metal2 3384 1042 3396 1042 5 ShB
rlabel metal2 696 1042 708 1042 5 COut
rlabel metal2 768 1042 780 1042 5 Sum
rlabel metal2 504 1042 516 1042 5 CIn
rlabel metal2 3336 1042 3348 1042 5 A
rlabel metal1 557 917 557 917 1 FA_1
rlabel metal1 634 941 634 941 1 FA_2
rlabel metal2 72 0 84 0 1 ZeroA
rlabel metal2 72 1042 84 1042 5 ZeroA
rlabel metal1 0 892 0 902 3 B
rlabel metal1 0 870 0 880 3 A
rlabel metal2 3696 0 3708 0 1 Sh8B_L
rlabel metal2 3744 0 3756 0 1 Sh8C_L
rlabel metal2 3792 1042 3804 1042 5 Sh8D_L
rlabel metal2 3648 0 3660 0 1 Sh8A_L
rlabel metal2 3696 1042 3708 1042 5 Sh8B_L
rlabel metal2 5760 1042 5772 1042 5 Sh8H_R
rlabel metal2 5712 1042 5724 1042 5 Sh8G_R
rlabel metal2 5664 1042 5676 1042 5 Sh8F_R
rlabel metal2 5616 1042 5628 1042 5 Sh8E_R
rlabel metal2 5568 1042 5580 1042 5 Sh8D_R
rlabel metal2 5760 0 5772 0 1 Sh8G_R
rlabel metal2 5712 0 5724 0 1 Sh8F_R
rlabel metal2 5664 0 5676 0 1 Sh8E_R
rlabel metal2 5616 0 5628 0 1 Sh8D_R
rlabel metal2 5568 0 5580 0 1 Sh8C_R
rlabel metal2 6000 0 6012 0 1 Sh4
rlabel metal2 6000 1042 6012 1042 5 Sh4
rlabel metal2 6816 0 6828 0 1 Sh1
rlabel metal2 6456 0 6468 0 1 Sh2
rlabel metal2 7176 0 7188 0 1 ShOut
rlabel metal2 6120 1042 6132 1042 5 Sh4A_R
rlabel metal2 6168 1042 6180 1042 5 Sh4B_R
rlabel metal2 6216 1042 6228 1042 5 Sh4C_R
rlabel metal2 6528 1042 6540 1042 5 Sh2A_R
rlabel metal2 6576 1042 6588 1042 5 Sh2B_R
rlabel metal2 7176 1042 7188 1042 5 ShOut
rlabel metal2 6456 1042 6468 1042 5 Sh2
rlabel metal2 6816 1042 6828 1042 5 Sh1
rlabel metal2 6216 0 6228 0 1 Sh4B_R
rlabel metal2 6168 0 6180 0 1 Sh4A_R
rlabel metal2 6120 0 6132 0 1 Sh4Z_R
rlabel metal2 6528 0 6540 0 1 Sh2Z_R
rlabel metal2 6576 0 6588 0 1 Sh2A_R
rlabel metal2 6888 0 6900 0 1 Sh1_R_Out
rlabel metal2 6888 1042 6900 1042 5 Sh1_R_In
rlabel metal2 7584 1042 7596 1042 5 ALUEnable
rlabel metal1 7704 51 7704 61 7 ALU_Out
rlabel metal2 7584 0 7596 0 1 ALUEnable
rlabel metal1 7296 51 7296 61 1 LLI_In
rlabel metal1 7296 892 7296 902 1 B
rlabel metal1 7488 51 7488 61 1 LLI_Out
rlabel metal2 6072 0 6084 0 1 Sh4Y_L
rlabel metal2 6072 1042 6084 1042 5 Sh4Z_R
rlabel metal2 3984 0 3996 0 1 Sh8H_L
rlabel metal2 4296 1042 4308 1042 5 Sh4Z_L
rlabel metal2 4344 1042 4356 1042 5 Sh4A_L
rlabel metal2 4296 0 4308 0 1 Sh4A_L
rlabel metal2 5352 0 5364 0 1 Sh8
rlabel metal2 5377 0 5389 0 1 ShR
rlabel metal2 5377 1042 5389 1042 5 ShR
rlabel metal2 4752 1042 4764 1042 5 Sh2A_L
rlabel metal2 4800 1042 4812 1042 5 Sh2B_L
rlabel metal2 4392 1042 4404 1042 5 Sh4B_L
rlabel metal2 4440 1042 4452 1042 5 Sh4C_L
rlabel metal2 5424 1042 5436 1042 5 Sh8A_R
rlabel metal2 5472 1042 5484 1042 5 Sh8B_R
rlabel metal2 5520 1042 5532 1042 5 Sh8C_R
rlabel metal2 5352 1042 5364 1042 5 Sh8
rlabel metal2 4752 0 4764 0 1 Sh2B_L
rlabel metal2 4800 0 4812 0 1 Sh2C_L
rlabel metal2 4344 0 4356 0 1 Sh4B_L
rlabel metal2 4392 0 4404 0 1 Sh4C_L
rlabel metal2 4440 0 4452 0 1 Sh4D_L
rlabel metal2 5520 0 5532 0 1 Sh8B_R
rlabel metal2 5472 0 5484 0 1 Sh8A_R
rlabel metal2 5424 0 5436 0 1 Sh8Z_R
rlabel metal2 5184 0 5196 0 1 Sh1_L_In
rlabel metal2 5184 1042 5196 1042 5 Sh1_L_Out
rlabel metal2 3888 1042 3900 1042 5 Sh8F_L
rlabel metal2 3840 1042 3852 1042 5 Sh8E_L
rlabel metal2 3936 1042 3948 1042 5 Sh8G_L
rlabel metal2 3984 1042 3996 1042 5 Sh8H_L
rlabel metal2 3792 0 3804 0 1 Sh8D_L
rlabel metal2 3840 0 3852 0 1 Sh8E_L
rlabel metal2 3888 0 3900 0 1 Sh8F_L
rlabel metal2 3936 0 3948 0 1 Sh8G_L
rlabel metal2 7512 1042 7524 1042 5 AluOut
<< end >>
