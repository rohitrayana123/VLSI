magic
tech c035u
timestamp 1394620980
<< metal1 >>
rect 1573 1159 3023 1169
rect 3037 1159 20040 1169
rect 12709 1003 12744 1013
rect 12517 981 12744 991
rect 0 95 2903 105
rect 2917 95 3071 105
rect 3085 95 20040 105
rect 0 73 12623 83
rect 2629 51 12479 61
rect 12109 29 12431 39
rect 12325 7 12671 17
<< m2contact >>
rect 1559 1157 1573 1171
rect 3023 1157 3037 1171
rect 12695 1001 12709 1015
rect 12503 979 12517 993
rect 2903 93 2917 107
rect 3071 93 3085 107
rect 12623 71 12637 85
rect 2615 49 2629 63
rect 12479 49 12493 63
rect 12095 27 12109 41
rect 12431 27 12445 41
rect 12311 5 12325 19
rect 12671 5 12685 19
<< metal2 >>
rect 216 1153 228 1176
rect 360 1153 372 1176
rect 576 1153 588 1176
rect 1320 1153 1332 1176
rect 1488 1153 1500 1176
rect 1560 1153 1572 1157
rect 1872 1153 1884 1176
rect 2088 1153 2100 1176
rect 2832 1153 2844 1176
rect 3000 976 3012 1176
rect 3024 976 3036 1157
rect 3096 1153 3180 1165
rect 3216 1153 3228 1176
rect 3960 1153 3972 1176
rect 4176 1153 4188 1176
rect 4368 1153 4380 1176
rect 5112 1153 5124 1176
rect 5328 1153 5340 1176
rect 5520 1153 5532 1176
rect 6264 1153 6276 1176
rect 6480 1153 6492 1176
rect 6672 1153 6684 1176
rect 7416 1153 7428 1176
rect 7632 1153 7644 1176
rect 7824 1153 7836 1176
rect 8568 1153 8580 1176
rect 8784 1153 8796 1176
rect 8976 1153 8988 1176
rect 9720 1153 9732 1176
rect 9936 1153 9948 1176
rect 10128 1153 10140 1176
rect 10872 1153 10884 1176
rect 11088 1153 11100 1176
rect 11280 1153 11292 1176
rect 12024 1153 12036 1176
rect 12240 1153 12252 1176
rect 3096 976 3108 1153
rect 12408 976 12420 1176
rect 12504 976 12516 979
rect 12600 976 12612 1176
rect 12816 1153 12828 1176
rect 13080 1153 13092 1176
rect 13248 1153 13260 1176
rect 13416 1153 13428 1176
rect 13440 1153 13452 1176
rect 13512 1153 13524 1176
rect 13728 1153 13740 1176
rect 13872 1153 13884 1176
rect 14208 1153 14220 1176
rect 14568 1153 14580 1176
rect 14976 1153 14988 1176
rect 15312 1153 15324 1176
rect 15624 1153 15636 1176
rect 15960 1153 15972 1176
rect 16080 1153 16092 1176
rect 16128 1153 16140 1176
rect 16296 1153 16308 1176
rect 16392 1153 16404 1176
rect 16440 1153 16452 1176
rect 16488 1153 16500 1176
rect 16536 1153 16548 1176
rect 16584 1153 16596 1176
rect 16632 1153 16644 1176
rect 16680 1153 16692 1176
rect 16728 1153 16740 1176
rect 17040 1153 17052 1176
rect 17088 1153 17100 1176
rect 17136 1153 17148 1176
rect 17184 1153 17196 1176
rect 17496 1153 17508 1176
rect 17544 1153 17556 1176
rect 17928 1153 17940 1176
rect 18096 1153 18108 1176
rect 18121 1153 18133 1176
rect 18168 1153 18180 1176
rect 18216 1153 18228 1176
rect 18264 1153 18276 1176
rect 18312 1153 18324 1176
rect 18360 1153 18372 1176
rect 18408 1153 18420 1176
rect 18456 1153 18468 1176
rect 18504 1153 18516 1176
rect 18744 1153 18756 1176
rect 18816 1153 18828 1176
rect 18864 1153 18876 1176
rect 18912 1153 18924 1176
rect 18960 1153 18972 1176
rect 19200 1153 19212 1176
rect 19272 1153 19284 1176
rect 19320 1153 19332 1176
rect 19560 1153 19572 1176
rect 19632 1153 19644 1176
rect 19920 1153 19932 1176
rect 12696 976 12708 1001
rect 216 0 228 111
rect 360 0 372 111
rect 576 0 588 111
rect 1320 0 1332 111
rect 1488 0 1500 111
rect 1872 0 1884 111
rect 2088 0 2100 111
rect 2616 63 2628 111
rect 2832 0 2844 111
rect 2904 107 2916 111
rect 3000 0 3012 177
rect 3072 107 3084 177
rect 3216 0 3228 111
rect 3960 0 3972 111
rect 4176 0 4188 111
rect 4368 0 4380 111
rect 5112 0 5124 111
rect 5328 0 5340 111
rect 5520 0 5532 111
rect 6264 0 6276 111
rect 6480 0 6492 111
rect 6672 0 6684 111
rect 7416 0 7428 111
rect 7632 0 7644 111
rect 7824 0 7836 111
rect 8568 0 8580 111
rect 8784 0 8796 111
rect 8976 0 8988 111
rect 9720 0 9732 111
rect 9936 0 9948 111
rect 10128 0 10140 111
rect 10872 0 10884 111
rect 11088 0 11100 111
rect 11280 0 11292 111
rect 12024 0 12036 111
rect 12096 41 12108 111
rect 12240 0 12252 111
rect 12312 19 12324 111
rect 12408 0 12420 177
rect 12432 41 12444 177
rect 12480 63 12492 177
rect 12600 0 12612 177
rect 12624 85 12636 177
rect 12672 19 12684 177
rect 12816 0 12828 111
rect 13080 0 13092 111
rect 13248 0 13260 111
rect 13440 0 13452 111
rect 13728 0 13740 111
rect 13872 0 13884 111
rect 14208 0 14220 111
rect 14568 0 14580 111
rect 14976 0 14988 111
rect 15312 0 15324 111
rect 15624 0 15636 111
rect 15960 0 15972 111
rect 16128 0 16140 111
rect 16296 0 16308 111
rect 16392 0 16404 111
rect 16440 0 16452 111
rect 16488 0 16500 111
rect 16536 0 16548 111
rect 16584 0 16596 111
rect 16632 0 16644 111
rect 16680 0 16692 111
rect 16728 0 16740 111
rect 17040 0 17052 111
rect 17088 0 17100 111
rect 17136 0 17148 111
rect 17184 0 17196 111
rect 17496 0 17508 111
rect 17544 0 17556 111
rect 17928 0 17940 111
rect 18096 0 18108 111
rect 18121 0 18133 111
rect 18168 0 18180 111
rect 18216 0 18228 111
rect 18264 0 18276 111
rect 18312 0 18324 111
rect 18360 0 18372 111
rect 18408 0 18420 111
rect 18456 0 18468 111
rect 18504 0 18516 111
rect 18744 0 18756 111
rect 18816 0 18828 111
rect 18864 0 18876 111
rect 18912 0 18924 111
rect 18960 0 18972 111
rect 19200 0 19212 111
rect 19272 0 19284 111
rect 19320 0 19332 111
rect 19560 0 19572 111
rect 19632 0 19644 111
rect 19920 0 19932 111
use Pc_slice Pc_slice_0
timestamp 1394475379
transform 1 0 0 0 1 111
box 0 0 2952 1042
use mux2 mux2_0
timestamp 1386235218
transform 1 0 2952 0 1 177
box 0 0 192 799
use regBlock_slice regBlock_slice_0
timestamp 1394620980
transform 1 0 3144 0 1 111
box 0 0 9216 1042
use mux2 mux2_1
timestamp 1386235218
transform 1 0 12360 0 1 177
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 12552 0 1 177
box 0 0 192 799
use ALUSlice ALUSlice_0
timestamp 1394559926
transform 1 0 12744 0 1 111
box 0 0 7296 1042
<< labels >>
rlabel metal1 3096 100 3096 100 1 SysBus
rlabel metal1 12353 34 12353 34 1 Rd1
rlabel metal1 12355 11 12355 11 1 Rd2
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 2088 0 2100 0 1 PcWe
rlabel metal2 2832 0 2844 0 1 PcEn
rlabel metal2 3000 0 3012 0 1 WdSel
rlabel metal2 3960 0 3972 0 1 Rs1[0]
rlabel metal2 4368 0 4380 0 1 Rw[1]
rlabel metal2 5112 0 5124 0 1 Rs1[1]
rlabel metal2 5328 0 5340 0 1 Rs2[1]
rlabel metal2 5520 0 5532 0 1 Rw[2]
rlabel metal2 6264 0 6276 0 1 Rs1[2]
rlabel metal2 6480 0 6492 0 1 Rs2[2]
rlabel metal2 6672 0 6684 0 1 Rw[3]
rlabel metal2 7416 0 7428 0 1 Rs1[3]
rlabel metal2 7632 0 7644 0 1 Rs2[3]
rlabel metal2 7824 0 7836 0 1 Rw[4]
rlabel metal2 8568 0 8580 0 1 Rs1[4]
rlabel metal2 8784 0 8796 0 1 Rs2[4]
rlabel metal2 8976 0 8988 0 1 Rw[5]
rlabel metal2 9720 0 9732 0 1 Rs1[5]
rlabel metal2 9936 0 9948 0 1 Rs2[5]
rlabel metal2 10128 0 10140 0 1 Rw[6]
rlabel metal2 10872 0 10884 0 1 Rs1[6]
rlabel metal2 11088 0 11100 0 1 Rs2[6]
rlabel metal2 11280 0 11292 0 1 Rw[7]
rlabel metal2 12024 0 12036 0 1 Rs1[7]
rlabel metal2 12240 0 12252 0 1 Rs2[7]
rlabel metal1 12352 100 12352 100 1 SysBus
rlabel metal1 12353 78 12353 78 1 Imm
rlabel metal1 12354 56 12354 56 1 Pc
rlabel metal2 3216 0 3228 0 1 Rw[0]
rlabel metal2 4176 0 4188 0 1 Rs2[0]
rlabel metal1 0 95 0 105 1 SysBus
rlabel metal1 0 73 0 83 1 Imm
rlabel metal2 12240 1176 12252 1176 5 Rs2[7]
rlabel metal2 12024 1176 12036 1176 5 Rs1[7]
rlabel metal2 11280 1176 11292 1176 5 Rw[7]
rlabel metal2 11088 1176 11100 1176 5 Rs2[6]
rlabel metal2 10872 1176 10884 1176 5 Rs1[6]
rlabel metal2 10128 1176 10140 1176 5 Rw[6]
rlabel metal2 9720 1176 9732 1176 5 Rs1[5]
rlabel metal2 9936 1176 9948 1176 5 Rs2[5]
rlabel metal2 8976 1176 8988 1176 5 Rw[5]
rlabel metal2 8784 1176 8796 1176 5 Rs2[4]
rlabel metal2 8568 1176 8580 1176 5 Rs1[4]
rlabel metal2 7824 1176 7836 1176 5 Rw[4]
rlabel metal2 7632 1176 7644 1176 5 Rs2[3]
rlabel metal2 7416 1176 7428 1176 5 Rs1[3]
rlabel metal2 6672 1176 6684 1176 5 Rw[3]
rlabel metal2 6480 1176 6492 1176 5 Rs2[2]
rlabel metal2 6264 1176 6276 1176 5 Rs1[2]
rlabel metal2 5520 1176 5532 1176 5 Rw[2]
rlabel metal2 5328 1176 5340 1176 5 Rs2[1]
rlabel metal2 5112 1176 5124 1176 5 Rs1[1]
rlabel metal2 4368 1176 4380 1176 5 Rw[1]
rlabel metal2 4176 1176 4188 1176 5 Rs2[0]
rlabel metal2 3960 1176 3972 1176 5 Rs1[0]
rlabel metal2 3216 1176 3228 1176 5 Rw[0]
rlabel metal2 3000 1176 3012 1176 5 WdSel
rlabel metal2 2832 1176 2844 1176 5 PcEn
rlabel metal2 2088 1176 2100 1176 5 PcWe
rlabel metal2 1872 1176 1884 1176 5 PcSel[1]
rlabel metal2 1488 1176 1500 1176 5 PcSel[0]
rlabel metal2 1320 1176 1332 1176 5 LrEn
rlabel metal2 576 1176 588 1176 5 LrWe
rlabel metal2 360 1176 372 1176 5 LrSel
rlabel metal2 216 1176 228 1176 5 PcIncCout
rlabel metal2 12600 0 12612 0 1 Op2Sel
rlabel metal2 12408 0 12420 0 1 Op1Sel
rlabel metal1 12733 99 12733 99 1 SysBus
rlabel metal2 12408 1176 12420 1176 5 Op1Sel
rlabel metal2 12600 1176 12612 1176 5 Op2Sel
rlabel metal1 12750 1164 12750 1164 6 AluOut
rlabel metal2 13440 0 13452 0 1 CIn_Slice
rlabel metal2 13728 0 13740 0 1 nZ_prev
rlabel metal2 13080 0 13092 0 1 SUB
rlabel metal2 16128 0 16140 0 1 ShB
rlabel metal2 16296 0 16308 0 1 ShL
rlabel metal2 15960 0 15972 0 1 NOR
rlabel metal2 15624 0 15636 0 1 NAND
rlabel metal2 15312 0 15324 0 1 NOT
rlabel metal2 14976 0 14988 0 1 XOR
rlabel metal2 14568 0 14580 0 1 OR
rlabel metal2 14208 0 14220 0 1 AND
rlabel metal2 13248 0 13260 0 1 CIn
rlabel metal2 13872 0 13884 0 1 FAOut
rlabel metal2 12816 0 12828 0 1 ZeroA
rlabel metal2 16440 0 16452 0 1 Sh8B_L
rlabel metal2 16488 0 16500 0 1 Sh8C_L
rlabel metal2 16392 0 16404 0 1 Sh8A_L
rlabel metal2 18504 0 18516 0 1 Sh8G_R
rlabel metal2 18456 0 18468 0 1 Sh8F_R
rlabel metal2 18408 0 18420 0 1 Sh8E_R
rlabel metal2 18360 0 18372 0 1 Sh8D_R
rlabel metal2 18312 0 18324 0 1 Sh8C_R
rlabel metal2 18744 0 18756 0 1 Sh4
rlabel metal2 19560 0 19572 0 1 Sh1
rlabel metal2 19200 0 19212 0 1 Sh2
rlabel metal2 19920 0 19932 0 1 ShOut
rlabel metal2 18960 0 18972 0 1 Sh4B_R
rlabel metal2 18912 0 18924 0 1 Sh4A_R
rlabel metal2 18864 0 18876 0 1 Sh4Z_R
rlabel metal2 19272 0 19284 0 1 Sh2Z_R
rlabel metal2 19320 0 19332 0 1 Sh2A_R
rlabel metal2 19632 0 19644 0 1 Sh1_R_Out
rlabel metal2 18816 0 18828 0 1 Sh4Y_L
rlabel metal2 16728 0 16740 0 1 Sh8H_L
rlabel metal2 17040 0 17052 0 1 Sh4A_L
rlabel metal2 18096 0 18108 0 1 Sh8
rlabel metal2 18121 0 18133 0 1 ShR
rlabel metal2 17496 0 17508 0 1 Sh2B_L
rlabel metal2 17544 0 17556 0 1 Sh2C_L
rlabel metal2 17088 0 17100 0 1 Sh4B_L
rlabel metal2 17136 0 17148 0 1 Sh4C_L
rlabel metal2 17184 0 17196 0 1 Sh4D_L
rlabel metal2 18264 0 18276 0 1 Sh8B_R
rlabel metal2 18216 0 18228 0 1 Sh8A_R
rlabel metal2 18168 0 18180 0 1 Sh8Z_R
rlabel metal2 17928 0 17940 0 1 Sh1_L_In
rlabel metal2 16536 0 16548 0 1 Sh8D_L
rlabel metal2 16584 0 16596 0 1 Sh8E_L
rlabel metal2 16632 0 16644 0 1 Sh8F_L
rlabel metal2 16680 0 16692 0 1 Sh8G_L
rlabel metal2 13416 1176 13428 1176 5 CIn_Slice
rlabel metal2 16296 1176 16308 1176 5 ShL
rlabel metal2 13872 1176 13884 1176 5 FAOut
rlabel metal2 13728 1176 13740 1176 5 nZ
rlabel metal2 13080 1176 13092 1176 5 SUB
rlabel metal2 14208 1176 14220 1176 5 AND
rlabel metal2 14568 1176 14580 1176 5 OR
rlabel metal2 14976 1176 14988 1176 5 XOR
rlabel metal2 15312 1176 15324 1176 5 NOT
rlabel metal2 15624 1176 15636 1176 5 NAND
rlabel metal2 15960 1176 15972 1176 5 NOR
rlabel metal2 16128 1176 16140 1176 5 ShB
rlabel metal2 13440 1176 13452 1176 5 COut
rlabel metal2 13512 1176 13524 1176 5 Sum
rlabel metal2 13248 1176 13260 1176 5 CIn
rlabel metal2 12816 1176 12828 1176 5 ZeroA
rlabel metal2 18504 1176 18516 1176 5 Sh8H_R
rlabel metal2 18456 1176 18468 1176 5 Sh8G_R
rlabel metal2 18408 1176 18420 1176 5 Sh8F_R
rlabel metal2 18360 1176 18372 1176 5 Sh8E_R
rlabel metal2 18312 1176 18324 1176 5 Sh8D_R
rlabel metal2 18744 1176 18756 1176 5 Sh4
rlabel metal2 18864 1176 18876 1176 5 Sh4A_R
rlabel metal2 18912 1176 18924 1176 5 Sh4B_R
rlabel metal2 18960 1176 18972 1176 5 Sh4C_R
rlabel metal2 19272 1176 19284 1176 5 Sh2A_R
rlabel metal2 19320 1176 19332 1176 5 Sh2B_R
rlabel metal2 19920 1176 19932 1176 5 ShOut
rlabel metal2 19200 1176 19212 1176 5 Sh2
rlabel metal2 19560 1176 19572 1176 5 Sh1
rlabel metal2 18816 1176 18828 1176 5 Sh4Z_R
rlabel metal2 17040 1176 17052 1176 5 Sh4Z_L
rlabel metal2 17088 1176 17100 1176 5 Sh4A_L
rlabel metal2 18121 1176 18133 1176 5 ShR
rlabel metal2 17496 1176 17508 1176 5 Sh2A_L
rlabel metal2 17544 1176 17556 1176 5 Sh2B_L
rlabel metal2 17136 1176 17148 1176 5 Sh4B_L
rlabel metal2 17184 1176 17196 1176 5 Sh4C_L
rlabel metal2 18168 1176 18180 1176 5 Sh8A_R
rlabel metal2 18216 1176 18228 1176 5 Sh8B_R
rlabel metal2 18264 1176 18276 1176 5 Sh8C_R
rlabel metal2 18096 1176 18108 1176 5 Sh8
rlabel metal2 17928 1176 17940 1176 5 Sh1_L_Out
rlabel metal2 16080 1176 16092 1176 5 A
rlabel metal1 20040 1159 20040 1169 7 AluOut
rlabel metal1 20040 95 20040 105 7 SysBus
rlabel metal2 16440 1176 16452 1176 5 Sh8A_L
rlabel metal2 16536 1176 16548 1176 5 Sh8C_L
rlabel metal2 16584 1176 16596 1176 5 Sh8D_L
rlabel metal2 16488 1176 16500 1176 5 Sh8B_L
rlabel metal2 16680 1176 16692 1176 5 Sh8F_L
rlabel metal2 16632 1176 16644 1176 5 Sh8E_L
rlabel metal2 16728 1176 16740 1176 5 Sh8G_L
rlabel metal2 16392 1176 16404 1176 5 Sh8Z_L
rlabel metal2 19632 1176 19644 1176 5 Sh1_R_in
rlabel metal1 12643 983 12643 983 1 Op1
rlabel metal1 12721 1008 12721 1008 1 Op2
<< end >>
