magic
tech c035u
timestamp 1396389552
<< metal1 >>
rect 0 96 1469 106
rect 0 29 1469 39
<< metal2 >>
rect 5 911 205 1111
rect 221 911 233 1111
rect 245 911 257 1111
rect 269 911 281 1111
rect 293 911 305 1111
rect 5 0 205 112
rect 221 0 233 112
rect 245 0 257 112
rect 269 0 281 112
rect 293 0 305 112
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 5 0 1 112
box 0 0 1464 799
<< labels >>
rlabel metal2 5 1111 205 1111 5 Vdd!
rlabel metal2 221 1111 233 1111 5 SDO
rlabel metal2 245 1111 257 1111 5 Test
rlabel metal2 269 1111 281 1111 5 Clock
rlabel metal2 293 1111 305 1111 5 nReset
rlabel metal1 0 29 0 39 3 SysBus
rlabel metal1 0 96 0 106 3 Ir
rlabel metal1 1469 96 1469 106 7 Ir
rlabel metal1 1469 29 1469 39 7 SysBus
rlabel metal2 5 0 205 0 1 Vdd!
rlabel metal2 221 0 233 0 1 SDI
rlabel metal2 245 0 257 0 1 Test
rlabel metal2 269 0 281 0 1 Clock
rlabel metal2 293 0 305 0 1 nReset
<< end >>
