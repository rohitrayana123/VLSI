magic
tech c035u
timestamp 1396388721
<< nwell >>
rect 1464 665 3504 1063
rect 15073 665 15696 1063
rect 23352 665 24696 1063
<< pwell >>
rect 1464 264 3504 665
rect 15073 271 15696 665
rect 23352 264 24696 665
<< pohmic >>
rect 1464 340 1470 350
rect 3498 340 3504 350
rect 15073 340 15078 350
rect 15690 340 15696 350
rect 23352 340 23356 350
rect 24690 340 24696 350
<< nohmic >>
rect 1464 1000 1470 1010
rect 3500 1000 3504 1010
rect 15073 1000 15078 1010
rect 15690 1000 15696 1010
rect 23352 1000 23356 1010
rect 24690 1000 24696 1010
<< psubstratetap >>
rect 1470 340 3498 356
rect 15078 340 15690 356
rect 23356 340 24690 356
<< nsubstratetap >>
rect 1470 994 3500 1010
rect 15078 994 15690 1010
rect 23356 994 24690 1010
<< metal1 >>
rect 4405 1267 5591 1277
rect 4453 1245 5543 1255
rect 5798 1249 5856 1259
rect 4069 1223 5159 1233
rect 5774 1227 5856 1237
rect 4021 1201 5207 1211
rect 5245 1201 5351 1211
rect 5437 1201 5760 1211
rect 5821 1204 5856 1214
rect 3589 1179 4823 1189
rect 4861 1179 4967 1189
rect 5053 1179 5784 1189
rect 15073 1178 15696 1188
rect 3637 1157 4775 1167
rect 4957 1157 5327 1167
rect 5341 1157 5711 1167
rect 15073 1156 15696 1166
rect 3805 1135 4175 1145
rect 4189 1135 4559 1145
rect 4765 1135 5135 1145
rect 5149 1135 5519 1145
rect 5629 1135 5735 1145
rect 15073 1134 15696 1144
rect 3901 1113 5856 1123
rect 15073 1112 15696 1122
rect 3661 1091 3815 1101
rect 4093 1091 4199 1101
rect 4285 1091 5856 1101
rect 15073 1090 15696 1100
rect 3565 1069 3983 1079
rect 3997 1069 4367 1079
rect 4477 1068 4583 1078
rect 4669 1068 5856 1078
rect 15073 1068 15696 1078
rect 1464 1046 3504 1056
rect 15073 1046 15696 1056
rect 23352 1046 24696 1056
rect 1464 1023 3504 1033
rect 15073 1023 15696 1033
rect 23352 1023 24696 1033
rect 1464 994 1470 1010
rect 3500 994 3504 1010
rect 1464 985 3504 994
rect 15073 994 15078 1010
rect 15690 994 15696 1010
rect 15073 985 15696 994
rect 23352 994 23356 1010
rect 24690 994 24696 1010
rect 23352 985 24696 994
rect 1464 356 3504 365
rect 1464 340 1470 356
rect 3498 340 3504 356
rect 15073 356 15696 365
rect 15073 340 15078 356
rect 15690 340 15696 356
rect 23352 356 24696 365
rect 23352 340 23356 356
rect 24690 340 24696 356
rect 1464 317 3504 327
rect 15073 317 15696 327
rect 1464 294 3504 304
rect 15073 294 15696 304
rect 1464 271 3504 281
rect 15073 271 15696 281
rect 23352 249 23999 259
<< m2contact >>
rect 4391 1265 4405 1279
rect 5591 1265 5605 1279
rect 4439 1243 4453 1257
rect 5543 1243 5557 1257
rect 5784 1247 5798 1261
rect 4055 1221 4069 1235
rect 5159 1221 5173 1235
rect 5760 1226 5774 1240
rect 4007 1199 4021 1213
rect 5207 1199 5221 1213
rect 5231 1199 5245 1213
rect 5351 1199 5365 1213
rect 5423 1199 5437 1213
rect 5760 1199 5774 1213
rect 5807 1202 5821 1216
rect 3575 1178 3589 1192
rect 4823 1177 4837 1191
rect 4847 1177 4861 1191
rect 4967 1177 4981 1191
rect 5039 1177 5053 1191
rect 5784 1177 5798 1191
rect 3623 1155 3637 1169
rect 4775 1155 4789 1169
rect 4943 1155 4957 1169
rect 5327 1155 5341 1169
rect 5711 1155 5725 1169
rect 3791 1133 3805 1147
rect 4175 1133 4189 1147
rect 4559 1133 4573 1147
rect 4751 1133 4765 1147
rect 5135 1133 5149 1147
rect 5519 1133 5533 1147
rect 5615 1133 5629 1147
rect 5735 1133 5749 1147
rect 3887 1111 3901 1125
rect 3647 1089 3661 1103
rect 3815 1089 3829 1103
rect 4079 1089 4093 1103
rect 4199 1089 4213 1103
rect 4271 1089 4285 1103
rect 3551 1067 3565 1081
rect 3983 1067 3997 1081
rect 4367 1067 4381 1081
rect 4463 1066 4477 1080
rect 4583 1066 4597 1080
rect 4655 1066 4669 1080
rect 23999 247 24013 261
<< metal2 >>
rect 0 1063 200 1302
rect 216 1063 228 1302
rect 240 1063 252 1302
rect 264 1063 276 1302
rect 288 1063 300 1302
rect 3552 1081 3564 1302
rect 3576 1192 3588 1302
rect 3552 1063 3564 1067
rect 3576 1063 3588 1178
rect 3624 1169 3636 1302
rect 3624 1063 3636 1155
rect 3792 1147 3804 1302
rect 4008 1213 4020 1302
rect 4056 1235 4068 1302
rect 4392 1279 4404 1302
rect 3648 1063 3660 1089
rect 3792 1063 3804 1133
rect 3816 1063 3828 1089
rect 3888 1063 3900 1111
rect 3984 1063 3996 1067
rect 4008 1063 4020 1199
rect 4056 1063 4068 1221
rect 4080 1063 4092 1089
rect 4176 1063 4188 1133
rect 4200 1063 4212 1089
rect 4272 1063 4284 1089
rect 4368 1063 4380 1067
rect 4392 1063 4404 1265
rect 4440 1257 4452 1302
rect 4440 1063 4452 1243
rect 4752 1147 4764 1302
rect 4464 1063 4476 1066
rect 4560 1063 4572 1133
rect 4584 1063 4596 1066
rect 4656 1063 4668 1066
rect 4752 1063 4764 1133
rect 4776 1063 4788 1155
rect 4824 1063 4836 1177
rect 4848 1063 4860 1177
rect 4944 1169 4956 1302
rect 5978 1290 5990 1302
rect 6532 1290 6544 1302
rect 6556 1290 6568 1302
rect 6580 1290 6592 1302
rect 13969 1290 13981 1302
rect 13993 1290 14005 1302
rect 14185 1290 14197 1302
rect 14233 1290 14245 1302
rect 14377 1290 14389 1302
rect 14569 1290 14581 1302
rect 14761 1290 14773 1302
rect 14953 1290 14965 1302
rect 4944 1063 4956 1155
rect 4968 1063 4980 1177
rect 5040 1063 5052 1177
rect 5136 1063 5148 1133
rect 5160 1063 5172 1221
rect 5208 1063 5220 1199
rect 5232 1063 5244 1199
rect 5328 1063 5340 1155
rect 5352 1063 5364 1199
rect 5424 1063 5436 1199
rect 5520 1063 5532 1133
rect 5544 1063 5556 1243
rect 5592 1063 5604 1265
rect 5761 1213 5773 1226
rect 5785 1191 5797 1247
rect 16752 1239 16764 1302
rect 16944 1239 16956 1302
rect 17016 1239 17028 1302
rect 17112 1239 17124 1302
rect 21768 1239 21780 1302
rect 21960 1239 21972 1302
rect 22080 1239 22092 1302
rect 22200 1239 22212 1302
rect 23280 1239 23292 1302
rect 5616 1063 5628 1133
rect 5712 1063 5724 1155
rect 5736 1063 5748 1133
rect 5808 1063 5820 1202
rect 24816 1063 25016 1302
rect 0 0 200 264
rect 216 0 228 264
rect 240 0 252 264
rect 264 0 276 264
rect 288 0 300 264
rect 3720 254 3732 264
rect 3864 254 3876 264
rect 4104 254 4116 255
rect 4248 254 4260 264
rect 4632 254 4644 264
rect 5016 254 5028 264
rect 5256 254 5268 255
rect 5400 254 5412 264
rect 5784 254 5796 264
rect 3720 242 5796 254
rect 5928 0 5940 159
rect 6672 0 6684 159
rect 6888 0 6900 159
rect 7080 0 7092 159
rect 7824 0 7836 159
rect 8040 0 8052 159
rect 8232 0 8244 159
rect 8976 0 8988 159
rect 9192 0 9204 159
rect 9384 0 9396 159
rect 10128 0 10140 159
rect 10344 0 10356 159
rect 10536 0 10548 159
rect 11280 0 11292 159
rect 11496 0 11508 159
rect 11688 0 11700 159
rect 12432 0 12444 159
rect 12648 0 12660 159
rect 12840 0 12852 159
rect 13584 0 13596 159
rect 13800 0 13812 159
rect 13992 0 14004 159
rect 14736 0 14748 159
rect 14952 0 14964 159
rect 24000 0 24012 247
rect 24816 0 25016 264
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 0 0 1 264
box 0 0 1464 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 3504 0 1 264
box 0 0 192 799
use tiehigh tiehigh_3
timestamp 1386086759
transform 1 0 3696 0 1 264
box 0 0 48 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 3744 0 1 264
box 0 0 192 799
use mux2 mux2_8
timestamp 1386235218
transform 1 0 3936 0 1 264
box 0 0 192 799
use mux2 mux2_9
timestamp 1386235218
transform 1 0 4128 0 1 264
box 0 0 192 799
use mux2 mux2_10
timestamp 1386235218
transform 1 0 4320 0 1 264
box 0 0 192 799
use mux2 mux2_11
timestamp 1386235218
transform 1 0 4512 0 1 264
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4704 0 1 264
box 0 0 192 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 4896 0 1 264
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 5088 0 1 264
box 0 0 192 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 5280 0 1 264
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 5472 0 1 264
box 0 0 192 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 5664 0 1 264
box 0 0 192 799
use regBlock_decoder regBlock_decoder_0
timestamp 1395339189
transform 1 0 5856 0 1 159
box 0 0 9217 1131
use ALUDecoder_new ALUDecoder_new_0
timestamp 1396388070
transform 1 0 15696 0 1 0
box 0 0 7656 1239
use rightend rightend_0
timestamp 1386235834
transform 1 0 24696 0 1 264
box 0 0 320 799
<< labels >>
rlabel metal2 240 1302 252 1302 1 Test
rlabel metal2 264 1302 276 1302 1 Clock
rlabel metal2 288 1302 300 1302 1 nReset
rlabel metal2 0 1302 200 1302 5 Vdd!
rlabel metal2 216 1302 228 1302 5 SDO
rlabel metal2 24816 1302 25016 1302 1 GND!
rlabel metal1 5853 1209 5853 1209 1 Rw0
rlabel metal1 5852 1231 5852 1231 1 Rw1
rlabel metal1 5847 1251 5847 1251 1 Rw2
rlabel metal1 15661 1071 15661 1071 1 AOp0
rlabel metal1 15662 1093 15662 1093 1 AOp1
rlabel metal1 15662 1114 15662 1114 1 AOp2
rlabel metal1 15662 1139 15662 1139 1 AOp3
rlabel metal1 15661 1159 15661 1159 1 AOp4
rlabel metal1 15660 1182 15660 1182 1 ACin
rlabel metal2 4056 1302 4068 1302 5 Ir[6]
rlabel metal2 4008 1302 4020 1302 5 Ir[9]
rlabel metal2 3624 1302 3636 1302 5 Ir[7]
rlabel metal2 3576 1302 3588 1302 5 Ir[10]
rlabel metal2 3792 1302 3804 1302 5 Rs1Sel[1]
rlabel metal2 3552 1302 3564 1302 5 Rs1Sel[0]
rlabel metal2 4392 1302 4404 1302 5 Ir[8]
rlabel metal2 4440 1302 4452 1302 5 Ir[5]
rlabel metal2 4752 1302 4764 1302 5 RwSel[0]
rlabel metal2 4944 1302 4956 1302 5 RwSel[1]
rlabel metal2 13969 1302 13981 1302 1 AluOR[1]
rlabel metal2 13993 1302 14005 1302 5 Ir[15]
rlabel metal2 14185 1302 14197 1302 5 Ir[14]
rlabel metal2 14233 1302 14245 1302 1 AluOR[0]
rlabel metal2 14377 1302 14389 1302 5 Ir[13]
rlabel metal2 14569 1302 14581 1302 5 Ir[12]
rlabel metal2 14761 1302 14773 1302 5 Ir[11]
rlabel metal2 14953 1302 14965 1302 5 Cin
rlabel metal2 6580 1302 6592 1302 5 Ir[4]
rlabel metal2 6556 1302 6568 1302 5 Ir[3]
rlabel metal2 6532 1302 6544 1302 5 Ir[2]
rlabel metal2 23280 1302 23292 1302 5 ALUOutEn
rlabel metal2 5978 1302 5990 1302 5 RegWe
rlabel metal2 17016 1302 17028 1302 5 Flags[3]
rlabel metal2 16944 1302 16956 1302 5 Flags[1]
rlabel metal2 16752 1302 16764 1302 5 Flags[2]
rlabel metal2 21768 1302 21780 1302 5 Ir[3]
rlabel metal2 21960 1302 21972 1302 5 Ir[2]
rlabel metal2 22080 1302 22092 1302 5 Ir[1]
rlabel metal2 22200 1302 22212 1302 5 Ir[0]
rlabel metal2 17112 1302 17124 1302 5 Flags[0]
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 10344 0 10356 0 1 Rs2[3]
rlabel metal2 7824 0 7836 0 1 Rs1[1]
rlabel metal2 7080 0 7092 0 1 Rw[1]
rlabel metal2 14952 0 14964 0 1 Rs2[7]
rlabel metal2 14736 0 14748 0 1 Rs1[7]
rlabel metal2 13992 0 14004 0 1 Rw[7]
rlabel metal2 13800 0 13812 0 1 Rs2[6]
rlabel metal2 13584 0 13596 0 1 Rs1[6]
rlabel metal2 12840 0 12852 0 1 Rw[6]
rlabel metal2 12648 0 12660 0 1 Rs2[5]
rlabel metal2 12432 0 12444 0 1 Rs1[5]
rlabel metal2 11688 0 11700 0 1 Rw[5]
rlabel metal2 11496 0 11508 0 1 Rs2[4]
rlabel metal2 11280 0 11292 0 1 Rs1[4]
rlabel metal2 10536 0 10548 0 1 Rw[4]
rlabel metal2 10128 0 10140 0 1 Rs1[3]
rlabel metal2 9384 0 9396 0 1 Rw[3]
rlabel metal2 9192 0 9204 0 1 Rs2[2]
rlabel metal2 8976 0 8988 0 1 Rs1[2]
rlabel metal2 8232 0 8244 0 1 Rw[2]
rlabel metal2 8040 0 8052 0 1 Rs2[1]
rlabel metal2 6888 0 6900 0 1 Rs2[0]
rlabel metal2 6672 0 6684 0 1 Rs1[0]
rlabel metal2 5928 0 5940 0 1 Rw[0]
rlabel metal2 24818 0 25016 0 1 GND!
rlabel metal2 24000 0 24012 0 1 ALUOutEn
<< end >>
