magic
tech c035u
timestamp 1394307496
use slice17 slice17_0
timestamp 1394305018
transform 1 0 4334 0 1 17264
box -4329 0 10503 1795
use Datapath_slice Datapath_slice_0
array 0 0 14841 0 15 1079
timestamp 1394307282
transform 1 0 0 0 1 0
box 0 0 14841 1079
<< end >>
