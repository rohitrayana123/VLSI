magic
tech c035u
timestamp 1395422998
<< metal1 >>
rect 6816 41410 6826 41452
rect 6864 41410 6874 41452
rect 6816 41400 6874 41410
rect 5828 40416 5890 40426
rect 5880 40402 5890 40416
rect 6816 40405 6826 41400
rect 6912 40405 6922 41452
rect 10848 41266 10858 41452
rect 10896 41293 10906 41452
rect 14976 41437 14986 41452
rect 15024 41437 15034 41452
rect 19104 41437 19114 41452
rect 19152 41437 19162 41452
rect 19296 41437 19306 41452
rect 27360 41437 27370 41452
rect 27408 41437 27418 41452
rect 27552 41410 27562 41452
rect 31488 41437 31498 41452
rect 31536 41437 31546 41452
rect 11472 41400 27562 41410
rect 11472 41341 11482 41400
rect 31680 41410 31690 41452
rect 35616 41437 35626 41452
rect 35664 41413 35674 41452
rect 35808 41437 35818 41452
rect 27589 41400 31690 41410
rect 31717 41400 35639 41410
rect 35688 41400 36658 41410
rect 11496 41376 27407 41386
rect 11496 41341 11506 41376
rect 27445 41376 31487 41386
rect 31501 41376 35615 41386
rect 35688 41386 35698 41400
rect 35629 41376 35698 41386
rect 35712 41376 35807 41386
rect 11520 41352 15023 41362
rect 11520 41341 11530 41352
rect 15061 41352 35663 41362
rect 35712 41362 35722 41376
rect 36648 41386 36658 41400
rect 36648 41376 36682 41386
rect 35688 41352 35722 41362
rect 36504 41352 36658 41362
rect 11557 41328 31535 41338
rect 31560 41328 31703 41338
rect 31560 41314 31570 41328
rect 35688 41338 35698 41352
rect 35653 41328 35698 41338
rect 11448 41304 31570 41314
rect 11448 41293 11458 41304
rect 11581 41280 19151 41290
rect 19189 41280 27575 41290
rect 10848 41256 14975 41266
rect 10896 40405 10906 41231
rect 5880 40392 5903 40402
rect 11424 40378 11434 41256
rect 15013 41256 19103 41266
rect 19117 41256 27359 41266
rect 27373 41256 27431 41266
rect 11592 41232 19295 41242
rect 5828 40368 11434 40378
rect 5880 35722 5890 40368
rect 5904 35749 5914 40343
rect 6816 39778 6826 40343
rect 6912 39805 6922 40343
rect 10896 39805 10906 40343
rect 11448 39994 11458 41231
rect 11437 39984 11458 39994
rect 11472 39970 11482 41231
rect 11496 39973 11506 41231
rect 11520 39973 11530 41231
rect 11544 39973 11554 41231
rect 11568 39973 11578 41231
rect 11592 39973 11602 41232
rect 11616 41208 19175 41218
rect 11616 39973 11626 41208
rect 11640 41184 15047 41194
rect 11640 39973 11650 41184
rect 11664 41160 14999 41170
rect 11664 39973 11674 41160
rect 11413 39960 11482 39970
rect 11389 39936 11698 39946
rect 11352 39912 11495 39922
rect 11352 39898 11362 39912
rect 11688 39922 11698 39936
rect 11688 39912 11746 39922
rect 11293 39888 11362 39898
rect 11448 39888 11711 39898
rect 11376 39874 11386 39887
rect 11448 39877 11458 39888
rect 11736 39898 11746 39912
rect 11736 39888 11770 39898
rect 11269 39864 11386 39874
rect 11485 39864 11746 39874
rect 11232 39840 11279 39850
rect 11232 39805 11242 39840
rect 11317 39840 11698 39850
rect 11280 39816 11663 39826
rect 11280 39805 11290 39816
rect 11688 39805 11698 39840
rect 11341 39792 11663 39802
rect 11712 39802 11722 39839
rect 11736 39829 11746 39864
rect 11760 39850 11770 39888
rect 14976 39877 14986 41135
rect 27133 39936 29002 39946
rect 26413 39912 28967 39922
rect 28992 39922 29002 39936
rect 28992 39912 29170 39922
rect 26149 39888 29135 39898
rect 29160 39898 29170 39912
rect 29160 39888 29279 39898
rect 36504 39877 36514 41352
rect 36648 39877 36658 41352
rect 36672 40642 36682 41376
rect 36672 40632 40916 40642
rect 40848 40621 40858 40632
rect 40824 40584 40916 40594
rect 40824 40477 40834 40584
rect 40848 40477 40858 40559
rect 40800 40440 40916 40450
rect 18157 39864 29351 39874
rect 11760 39840 36671 39850
rect 17125 39816 29231 39826
rect 29269 39816 29303 39826
rect 29341 39816 36527 39826
rect 36661 39816 36719 39826
rect 11712 39792 11759 39802
rect 16933 39792 28943 39802
rect 28981 39792 36647 39802
rect 36685 39792 36754 39802
rect 36744 39781 36754 39792
rect 6816 39768 11711 39778
rect 11749 39768 36706 39778
rect 11208 39744 11303 39754
rect 5880 35712 5938 35722
rect 5828 35688 5890 35698
rect 5880 35677 5890 35688
rect 5928 35650 5938 35712
rect 5828 35640 5938 35650
rect 5880 30997 5890 35615
rect 5904 30997 5914 35615
rect 5928 30994 5938 35640
rect 5928 30984 5962 30994
rect 5828 30960 5938 30970
rect 5928 30949 5938 30960
rect 5952 30922 5962 30984
rect 5828 30912 5962 30922
rect 5880 26317 5890 30887
rect 5904 26317 5914 30887
rect 5928 26317 5938 30887
rect 5828 26280 5962 26290
rect 5880 21685 5890 26255
rect 5904 21685 5914 26255
rect 5928 21685 5938 26255
rect 5952 21685 5962 26280
rect 5828 21648 5986 21658
rect 5880 16957 5890 21623
rect 5904 18010 5914 21623
rect 5928 18058 5938 21623
rect 5952 18226 5962 21623
rect 5976 18634 5986 21648
rect 6912 18661 6922 39743
rect 10896 22621 10906 39743
rect 11208 39733 11218 39744
rect 11365 39744 11735 39754
rect 11773 39744 11794 39754
rect 11317 39720 11759 39730
rect 11784 39730 11794 39744
rect 15973 39744 29255 39754
rect 29293 39744 36671 39754
rect 36696 39754 36706 39768
rect 36696 39744 36802 39754
rect 36792 39733 36802 39744
rect 11784 39720 36767 39730
rect 11173 39696 11471 39706
rect 40800 39706 40810 40440
rect 11509 39696 40810 39706
rect 11136 39672 11231 39682
rect 11136 39637 11146 39672
rect 11389 39672 12071 39682
rect 15733 39672 29327 39682
rect 29365 39672 36695 39682
rect 36733 39672 36839 39682
rect 11184 39648 11639 39658
rect 11184 39610 11194 39648
rect 11773 39648 12191 39658
rect 14976 39658 14986 39671
rect 14976 39648 29218 39658
rect 11232 39624 11615 39634
rect 11232 39613 11242 39624
rect 11125 39600 11194 39610
rect 11485 39600 11591 39610
rect 11664 39589 11674 39647
rect 11101 39576 11567 39586
rect 11688 39586 11698 39647
rect 11712 39610 11722 39647
rect 11736 39634 11746 39647
rect 11736 39624 29183 39634
rect 29208 39634 29218 39648
rect 29245 39648 36719 39658
rect 36757 39648 36863 39658
rect 29208 39624 36503 39634
rect 36541 39624 36743 39634
rect 36781 39624 36898 39634
rect 11712 39600 12047 39610
rect 12085 39600 29279 39610
rect 29317 39600 36815 39610
rect 36888 39610 36898 39624
rect 36888 39600 36911 39610
rect 11688 39576 28919 39586
rect 28957 39576 36767 39586
rect 36805 39576 36946 39586
rect 36936 39565 36946 39576
rect 11077 39552 11135 39562
rect 11197 39552 36887 39562
rect 11040 39528 11087 39538
rect 11040 36797 11050 39528
rect 40824 39538 40834 40415
rect 11149 39528 40834 39538
rect 11088 39504 11543 39514
rect 11064 36797 11074 39503
rect 11088 36797 11098 39504
rect 11677 39504 12178 39514
rect 12168 39493 12178 39504
rect 12205 39504 29122 39514
rect 29112 39493 29122 39504
rect 29149 39504 36802 39514
rect 11112 36797 11122 39479
rect 11136 36797 11146 39479
rect 11160 36797 11170 39479
rect 11184 36797 11194 39479
rect 11208 36797 11218 39479
rect 11232 36797 11242 39479
rect 11256 36797 11266 39479
rect 11280 36797 11290 39479
rect 11304 36797 11314 39479
rect 11328 36797 11338 39479
rect 11352 36797 11362 39479
rect 11376 36797 11386 39479
rect 11400 36797 11410 39479
rect 11424 36797 11434 39479
rect 11448 36797 11458 39479
rect 11472 36767 11482 39479
rect 11496 36773 11506 39479
rect 11520 36773 11530 39479
rect 11016 36757 11482 36767
rect 11016 36706 11026 36757
rect 11485 36734 11572 36744
rect 11544 36706 11572 36712
rect 11016 36702 11572 36706
rect 11016 36696 11554 36702
rect 11053 36678 11554 36682
rect 11053 36672 11572 36678
rect 11544 36668 11572 36672
rect 11064 35605 11074 36647
rect 11088 35605 11098 36647
rect 11112 35605 11122 36647
rect 11136 35605 11146 36647
rect 11160 35605 11170 36647
rect 11184 35605 11194 36647
rect 11208 35605 11218 36647
rect 11232 35605 11242 36647
rect 11256 35605 11266 36647
rect 11280 35605 11290 36647
rect 11304 35605 11314 36647
rect 11328 35605 11338 36647
rect 11352 35605 11362 36647
rect 11376 35605 11386 36647
rect 11400 35578 11410 36647
rect 11424 35597 11434 36647
rect 11448 35597 11458 36647
rect 11472 35597 11482 36647
rect 11496 35597 11506 36647
rect 11520 35597 11530 36647
rect 11040 35568 11410 35578
rect 11040 35530 11050 35568
rect 11544 35558 11572 35568
rect 11544 35557 11554 35558
rect 11413 35547 11554 35557
rect 11544 35530 11572 35536
rect 11040 35526 11572 35530
rect 11040 35520 11554 35526
rect 11077 35502 11554 35506
rect 11077 35496 11572 35502
rect 11544 35492 11572 35496
rect 11088 34429 11098 35471
rect 11112 34429 11122 35471
rect 11136 34429 11146 35471
rect 11160 34429 11170 35471
rect 11184 34429 11194 35471
rect 11208 34429 11218 35471
rect 11232 34402 11242 35471
rect 11256 34437 11266 35471
rect 11280 34437 11290 35471
rect 11304 34437 11314 35471
rect 11328 34437 11338 35471
rect 11352 34437 11362 35471
rect 11376 34437 11386 35471
rect 11400 34437 11410 35471
rect 11424 34437 11434 35471
rect 11448 34437 11458 35471
rect 11472 34437 11482 35471
rect 11496 34437 11506 35471
rect 11520 34437 11530 35471
rect 11064 34392 11242 34402
rect 11064 34354 11074 34392
rect 11544 34382 11572 34392
rect 11544 34380 11554 34382
rect 11245 34370 11554 34380
rect 11544 34354 11572 34360
rect 11064 34350 11572 34354
rect 11064 34344 11554 34350
rect 11101 34326 11554 34330
rect 11101 34320 11572 34326
rect 11544 34316 11572 34320
rect 11112 33253 11122 34295
rect 11136 33253 11146 34295
rect 11160 33253 11170 34295
rect 11184 33253 11194 34295
rect 11208 33253 11218 34295
rect 11232 33253 11242 34295
rect 11256 33253 11266 34295
rect 11280 33253 11290 34295
rect 11304 33253 11314 34295
rect 11328 33253 11338 34295
rect 11352 33253 11362 34295
rect 11376 33253 11386 34295
rect 11400 33253 11410 34295
rect 11424 33227 11434 34295
rect 11448 33229 11458 34295
rect 11472 33229 11482 34295
rect 11496 33229 11506 34295
rect 11520 33229 11530 34295
rect 11088 33217 11434 33227
rect 11088 33178 11098 33217
rect 11544 33206 11572 33216
rect 11544 33204 11554 33206
rect 11437 33194 11554 33204
rect 11544 33178 11572 33184
rect 11088 33174 11572 33178
rect 11088 33168 11554 33174
rect 11125 33150 11554 33154
rect 11125 33144 11572 33150
rect 11544 33140 11572 33144
rect 11136 32077 11146 33119
rect 11160 32077 11170 33119
rect 11184 32077 11194 33119
rect 11208 32077 11218 33119
rect 11232 32077 11242 33119
rect 11256 32077 11266 33119
rect 11280 32077 11290 33119
rect 11304 32077 11314 33119
rect 11328 32077 11338 33119
rect 11352 32077 11362 33119
rect 11376 32077 11386 33119
rect 11400 32077 11410 33119
rect 11424 32077 11434 33119
rect 11448 32077 11458 33119
rect 11472 32077 11482 33119
rect 11496 32051 11506 33119
rect 11520 32053 11530 33119
rect 11112 32041 11506 32051
rect 11112 32002 11122 32041
rect 11544 32030 11572 32040
rect 11544 32028 11554 32030
rect 11509 32018 11554 32028
rect 11544 32002 11572 32008
rect 11112 31998 11572 32002
rect 11112 31992 11554 31998
rect 11149 31974 11554 31978
rect 11149 31968 11572 31974
rect 11544 31964 11572 31968
rect 11160 30901 11170 31943
rect 11184 30901 11194 31943
rect 11208 30901 11218 31943
rect 11232 30901 11242 31943
rect 11256 30901 11266 31943
rect 11280 30901 11290 31943
rect 11304 30901 11314 31943
rect 11328 30901 11338 31943
rect 11352 30901 11362 31943
rect 11376 30901 11386 31943
rect 11400 30901 11410 31943
rect 11424 30901 11434 31943
rect 11448 30875 11458 31943
rect 11472 30877 11482 31943
rect 11496 30877 11506 31943
rect 11520 30877 11530 31943
rect 11136 30865 11458 30875
rect 11136 30826 11146 30865
rect 11544 30854 11572 30864
rect 11544 30852 11554 30854
rect 11461 30842 11554 30852
rect 11544 30826 11572 30832
rect 11136 30822 11572 30826
rect 11136 30816 11554 30822
rect 11173 30798 11554 30802
rect 11173 30792 11572 30798
rect 11544 30788 11572 30792
rect 11184 29753 11194 30767
rect 11208 29753 11218 30767
rect 11232 29753 11242 30767
rect 11256 29726 11266 30767
rect 11280 29729 11290 30767
rect 11304 29729 11314 30767
rect 11328 29729 11338 30767
rect 11352 29729 11362 30767
rect 11376 29729 11386 30767
rect 11400 29729 11410 30767
rect 11424 29729 11434 30767
rect 11448 29729 11458 30767
rect 11472 29729 11482 30767
rect 11496 29729 11506 30767
rect 11520 29729 11530 30767
rect 11160 29716 11266 29726
rect 11160 29656 11170 29716
rect 11269 29678 11572 29688
rect 11160 29646 11572 29656
rect 11197 29622 11554 29626
rect 11197 29616 11572 29622
rect 11544 29612 11572 29616
rect 11208 28549 11218 29591
rect 11232 28549 11242 29591
rect 11256 28549 11266 29591
rect 11280 28549 11290 29591
rect 11304 28549 11314 29591
rect 11328 28549 11338 29591
rect 11352 28549 11362 29591
rect 11376 28549 11386 29591
rect 11400 28549 11410 29591
rect 11424 28549 11434 29591
rect 11448 28549 11458 29591
rect 11472 28549 11482 29591
rect 11496 28549 11506 29591
rect 11520 28525 11530 29591
rect 11197 28515 11530 28525
rect 11173 28488 11447 28498
rect 11544 28502 11572 28512
rect 11544 28501 11554 28502
rect 11533 28491 11554 28501
rect 11136 28464 11303 28474
rect 11136 27349 11146 28464
rect 11544 28474 11572 28480
rect 11461 28470 11572 28474
rect 11461 28464 11554 28470
rect 11304 28446 11554 28450
rect 11304 28440 11572 28446
rect 11160 27322 11170 28439
rect 11184 27325 11194 28439
rect 11208 27325 11218 28439
rect 11232 27325 11242 28439
rect 11256 27325 11266 28439
rect 11280 27325 11290 28439
rect 11304 27325 11314 28440
rect 11544 28436 11572 28440
rect 11328 27325 11338 28415
rect 11352 27325 11362 28415
rect 11376 27325 11386 28415
rect 11400 27325 11410 28415
rect 11424 27325 11434 28415
rect 11448 27325 11458 28415
rect 11472 27325 11482 28415
rect 11496 27325 11506 28415
rect 11520 27325 11530 28415
rect 11125 27312 11170 27322
rect 11544 27298 11572 27304
rect 11088 27294 11572 27298
rect 11088 27288 11554 27294
rect 11088 26173 11098 27288
rect 11160 27270 11554 27274
rect 11160 27264 11572 27270
rect 11112 26173 11122 27263
rect 11136 26173 11146 27263
rect 11160 26173 11170 27264
rect 11544 27260 11572 27264
rect 11184 26173 11194 27239
rect 11208 26173 11218 27239
rect 11232 26173 11242 27239
rect 11256 26173 11266 27239
rect 11280 26173 11290 27239
rect 11304 26173 11314 27239
rect 11328 26173 11338 27239
rect 11352 26173 11362 27239
rect 11376 26146 11386 27239
rect 11400 26149 11410 27239
rect 11424 26149 11434 27239
rect 11448 26149 11458 27239
rect 11472 26149 11482 27239
rect 11496 26149 11506 27239
rect 11520 26149 11530 27239
rect 11077 26136 11386 26146
rect 11040 26112 11351 26122
rect 11040 24997 11050 26112
rect 11544 26122 11572 26128
rect 11389 26118 11572 26122
rect 11389 26112 11554 26118
rect 11352 26094 11554 26098
rect 11352 26088 11572 26094
rect 11064 24997 11074 26087
rect 11088 24997 11098 26087
rect 11112 24997 11122 26087
rect 11136 24997 11146 26087
rect 11160 24997 11170 26087
rect 11184 24997 11194 26087
rect 11208 24997 11218 26087
rect 11232 24997 11242 26087
rect 11256 24997 11266 26087
rect 11280 24997 11290 26087
rect 11304 24997 11314 26087
rect 11328 24970 11338 26087
rect 11352 24973 11362 26088
rect 11544 26084 11572 26088
rect 11376 24973 11386 26063
rect 11400 24973 11410 26063
rect 11424 24973 11434 26063
rect 11448 24973 11458 26063
rect 11472 24973 11482 26063
rect 11496 24973 11506 26063
rect 11520 24973 11530 26063
rect 11016 24960 11338 24970
rect 11016 24949 11026 24960
rect 11544 24946 11572 24952
rect 11341 24942 11572 24946
rect 11341 24936 11554 24942
rect 10992 24918 11554 24922
rect 10992 24912 11572 24918
rect 10992 23818 11002 24912
rect 11544 24908 11572 24912
rect 11016 23821 11026 24887
rect 11040 23821 11050 24887
rect 11064 23821 11074 24887
rect 11088 23821 11098 24887
rect 11112 23821 11122 24887
rect 11136 23821 11146 24887
rect 11160 23821 11170 24887
rect 11184 23821 11194 24887
rect 11208 23821 11218 24887
rect 11232 23821 11242 24887
rect 11256 23821 11266 24887
rect 11280 23821 11290 24887
rect 11304 23821 11314 24887
rect 11328 23821 11338 24887
rect 11352 23821 11362 24887
rect 10981 23808 11002 23818
rect 11376 23794 11386 24887
rect 11400 23797 11410 24887
rect 11424 23797 11434 24887
rect 11448 23797 11458 24887
rect 11472 23797 11482 24887
rect 11496 23797 11506 24887
rect 11520 23797 11530 24887
rect 10944 23784 11386 23794
rect 10944 22645 10954 23784
rect 11544 23770 11572 23776
rect 10992 23766 11572 23770
rect 10992 23760 11554 23766
rect 10968 22645 10978 23759
rect 10992 22645 11002 23760
rect 11376 23742 11554 23746
rect 11376 23736 11572 23742
rect 11016 22645 11026 23735
rect 11040 22645 11050 23735
rect 11064 22645 11074 23735
rect 11088 22645 11098 23735
rect 11112 22645 11122 23735
rect 11136 22645 11146 23735
rect 11160 22645 11170 23735
rect 11184 22645 11194 23735
rect 11208 22645 11218 23735
rect 11232 22645 11242 23735
rect 11256 22645 11266 23735
rect 11280 22645 11290 23735
rect 11304 22645 11314 23735
rect 11328 22645 11338 23735
rect 11352 22618 11362 23735
rect 11376 22621 11386 23736
rect 11544 23732 11572 23736
rect 11400 22621 11410 23711
rect 11424 22621 11434 23711
rect 11448 22621 11458 23711
rect 11472 22621 11482 23711
rect 11496 22621 11506 23711
rect 11520 22621 11530 23711
rect 10933 22608 11362 22618
rect 10872 22584 11231 22594
rect 10872 21469 10882 22584
rect 11544 22594 11572 22600
rect 11365 22590 11572 22594
rect 11365 22584 11554 22590
rect 11232 22566 11554 22570
rect 11232 22560 11572 22566
rect 10896 21469 10906 22559
rect 10920 21469 10930 22559
rect 10944 21469 10954 22559
rect 10968 21469 10978 22559
rect 10992 21442 11002 22559
rect 11016 21445 11026 22559
rect 11040 21445 11050 22559
rect 11064 21445 11074 22559
rect 11088 21445 11098 22559
rect 11112 21445 11122 22559
rect 11136 21445 11146 22559
rect 11160 21445 11170 22559
rect 11184 21445 11194 22559
rect 11208 21445 11218 22559
rect 11232 21445 11242 22560
rect 11544 22556 11572 22560
rect 11256 21445 11266 22535
rect 11280 21445 11290 22535
rect 11304 21445 11314 22535
rect 11328 21445 11338 22535
rect 11352 21445 11362 22535
rect 11376 21445 11386 22535
rect 11400 21445 11410 22535
rect 11424 21445 11434 22535
rect 11448 21445 11458 22535
rect 11472 21445 11482 22535
rect 11496 21445 11506 22535
rect 11520 21445 11530 22535
rect 10861 21432 11002 21442
rect 10824 21408 10919 21418
rect 10824 20293 10834 21408
rect 11544 21418 11572 21424
rect 11005 21414 11572 21418
rect 11005 21408 11554 21414
rect 10920 21390 11554 21394
rect 10920 21384 11572 21390
rect 10848 20293 10858 21383
rect 10872 20293 10882 21383
rect 10896 20293 10906 21383
rect 10920 20293 10930 21384
rect 11544 21380 11572 21384
rect 10944 20266 10954 21359
rect 10968 20269 10978 21359
rect 10992 20269 11002 21359
rect 11016 20269 11026 21359
rect 11040 20269 11050 21359
rect 11064 20269 11074 21359
rect 11088 20269 11098 21359
rect 11112 20269 11122 21359
rect 11136 20269 11146 21359
rect 11160 20269 11170 21359
rect 11184 20269 11194 21359
rect 11208 20269 11218 21359
rect 11232 20269 11242 21359
rect 11256 20269 11266 21359
rect 11280 20269 11290 21359
rect 11304 20269 11314 21359
rect 11328 20269 11338 21359
rect 11352 20269 11362 21359
rect 11376 20269 11386 21359
rect 11400 20269 11410 21359
rect 11424 20269 11434 21359
rect 11448 20269 11458 21359
rect 11472 20269 11482 21359
rect 11496 20269 11506 21359
rect 11520 20269 11530 21359
rect 10813 20256 10954 20266
rect 10776 20232 10871 20242
rect 10776 19117 10786 20232
rect 11544 20242 11572 20248
rect 10957 20238 11572 20242
rect 10957 20232 11554 20238
rect 10872 20214 11554 20218
rect 10872 20208 11572 20214
rect 10800 19117 10810 20207
rect 10824 19117 10834 20207
rect 10848 19117 10858 20207
rect 10872 19117 10882 20208
rect 11544 20204 11572 20208
rect 10896 19117 10906 20183
rect 10920 19117 10930 20183
rect 10944 19117 10954 20183
rect 10968 19117 10978 20183
rect 10992 19117 11002 20183
rect 11016 19117 11026 20183
rect 11040 19117 11050 20183
rect 11064 19117 11074 20183
rect 11088 19117 11098 20183
rect 11112 19090 11122 20183
rect 11136 19093 11146 20183
rect 11160 19093 11170 20183
rect 11184 19093 11194 20183
rect 11208 19093 11218 20183
rect 11232 19093 11242 20183
rect 11256 19093 11266 20183
rect 11280 19093 11290 20183
rect 11304 19093 11314 20183
rect 11328 19093 11338 20183
rect 11352 19093 11362 20183
rect 11376 19093 11386 20183
rect 11400 19093 11410 20183
rect 11424 19093 11434 20183
rect 11448 19093 11458 20183
rect 11472 19093 11482 20183
rect 11496 19093 11506 20183
rect 11520 19093 11530 20183
rect 10765 19080 11122 19090
rect 10728 19056 10823 19066
rect 10728 18826 10738 19056
rect 11544 19066 11572 19072
rect 11125 19062 11572 19066
rect 11125 19056 11554 19062
rect 10824 19038 11554 19042
rect 10824 19032 11572 19038
rect 10752 18853 10762 19031
rect 10776 18853 10786 19031
rect 10800 18853 10810 19031
rect 10824 18853 10834 19032
rect 11544 19028 11572 19032
rect 10848 18853 10858 19007
rect 10872 18853 10882 19007
rect 10896 18853 10906 19007
rect 10920 18853 10930 19007
rect 10944 18853 10954 19007
rect 10968 18853 10978 19007
rect 10992 18853 11002 19007
rect 11016 18853 11026 19007
rect 11040 18853 11050 19007
rect 11064 18853 11074 19007
rect 11088 18853 11098 19007
rect 11112 18853 11122 19007
rect 11136 18853 11146 19007
rect 11160 18853 11170 19007
rect 11184 18853 11194 19007
rect 11208 18853 11218 19007
rect 11232 18853 11242 19007
rect 11256 18853 11266 19007
rect 11280 18853 11290 19007
rect 11304 18853 11314 19007
rect 11328 18853 11338 19007
rect 11352 18853 11362 19007
rect 11376 18853 11386 19007
rect 11400 18853 11410 19007
rect 11424 18853 11434 19007
rect 11448 18853 11458 19007
rect 11472 18853 11482 19007
rect 11496 18853 11506 19007
rect 11520 18853 11530 19007
rect 36648 18853 36658 39479
rect 36672 18853 36682 39479
rect 36696 18853 36706 39479
rect 36720 18853 36730 39479
rect 36744 18853 36754 39479
rect 36768 18853 36778 39479
rect 36792 18850 36802 39504
rect 36816 18877 36826 39503
rect 36840 26314 36850 39503
rect 36864 30994 36874 39503
rect 36888 31138 36898 39503
rect 36912 35722 36922 39503
rect 36936 35866 36946 39503
rect 40848 35914 40858 40415
rect 40848 35904 40916 35914
rect 40848 35893 40858 35904
rect 36936 35856 40916 35866
rect 40848 35749 40858 35831
rect 36912 35712 40916 35722
rect 40848 31186 40858 35687
rect 40848 31176 40916 31186
rect 40848 31165 40858 31176
rect 36888 31128 40916 31138
rect 40848 31021 40858 31103
rect 36864 30984 40916 30994
rect 40848 26341 40858 30959
rect 36840 26304 40871 26314
rect 36792 18840 36874 18850
rect 36864 18829 36874 18840
rect 10728 18816 36839 18826
rect 10765 18792 36922 18802
rect 36912 18781 36922 18792
rect 11461 18768 36887 18778
rect 10776 18730 10786 18767
rect 11461 18744 12234 18754
rect 12949 18744 36167 18754
rect 36517 18744 36791 18754
rect 36853 18744 36946 18754
rect 36936 18733 36946 18744
rect 10776 18720 36839 18730
rect 11557 18696 12047 18706
rect 12085 18696 12210 18706
rect 14533 18696 27719 18706
rect 27757 18696 35423 18706
rect 36805 18696 36970 18706
rect 10800 18682 10810 18695
rect 10800 18672 36802 18682
rect 11581 18648 12186 18658
rect 14544 18648 27743 18658
rect 5976 18624 12162 18634
rect 11592 18600 12071 18610
rect 6912 18253 6922 18599
rect 10896 18562 10906 18599
rect 10008 18552 10906 18562
rect 10008 18538 10018 18552
rect 9744 18528 10018 18538
rect 9744 18514 9754 18528
rect 10045 18528 10823 18538
rect 9720 18504 9754 18514
rect 9720 18490 9730 18504
rect 10848 18514 10858 18527
rect 9781 18504 10858 18514
rect 9696 18480 9730 18490
rect 9696 18466 9706 18480
rect 10872 18490 10882 18527
rect 9757 18480 10882 18490
rect 9672 18456 9706 18466
rect 9672 18442 9682 18456
rect 10920 18466 10930 18599
rect 9733 18456 10930 18466
rect 9648 18432 9682 18442
rect 9648 18418 9658 18432
rect 10944 18442 10954 18599
rect 9709 18432 10954 18442
rect 9600 18408 9658 18418
rect 9600 18394 9610 18408
rect 10968 18418 10978 18599
rect 9685 18408 10978 18418
rect 9576 18384 9610 18394
rect 9576 18370 9586 18384
rect 10992 18394 11002 18599
rect 9637 18384 11002 18394
rect 9552 18360 9586 18370
rect 9552 18346 9562 18360
rect 11016 18370 11026 18599
rect 9613 18360 11026 18370
rect 9504 18336 9562 18346
rect 9504 18322 9514 18336
rect 11040 18346 11050 18599
rect 9589 18336 11050 18346
rect 9480 18312 9514 18322
rect 9480 18298 9490 18312
rect 11064 18322 11074 18599
rect 9541 18312 11074 18322
rect 11088 18322 11098 18599
rect 11112 18349 11122 18599
rect 11136 18349 11146 18599
rect 11160 18349 11170 18599
rect 11184 18349 11194 18599
rect 11208 18349 11218 18599
rect 11232 18349 11242 18599
rect 11256 18349 11266 18599
rect 11280 18349 11290 18599
rect 11304 18349 11314 18599
rect 11328 18349 11338 18599
rect 11352 18349 11362 18599
rect 11376 18349 11386 18599
rect 11400 18349 11410 18599
rect 11424 18349 11434 18599
rect 11448 18349 11458 18599
rect 11472 18349 11482 18599
rect 11496 18349 11506 18599
rect 11520 18349 11530 18599
rect 11544 18349 11554 18599
rect 11568 18349 11578 18599
rect 11592 18349 11602 18600
rect 11088 18312 11626 18322
rect 11616 18301 11626 18312
rect 9456 18288 9490 18298
rect 9456 18274 9466 18288
rect 9517 18288 11111 18298
rect 9432 18264 9466 18274
rect 9432 18250 9442 18264
rect 11136 18274 11146 18287
rect 9493 18264 11146 18274
rect 11160 18274 11170 18287
rect 11160 18264 11650 18274
rect 11640 18253 11650 18264
rect 12936 18253 12946 18647
rect 13512 18253 13522 18647
rect 13704 18253 13714 18647
rect 14496 18274 14506 18647
rect 14520 18301 14530 18647
rect 14544 18301 14554 18648
rect 16992 18624 27479 18634
rect 15048 18274 15058 18623
rect 15264 18298 15274 18623
rect 16008 18322 16018 18623
rect 16176 18346 16186 18623
rect 16560 18370 16570 18623
rect 16752 18394 16762 18623
rect 16968 18442 16978 18623
rect 16992 18469 17002 18624
rect 20688 18600 27287 18610
rect 17712 18442 17722 18599
rect 17880 18466 17890 18599
rect 20688 18469 20698 18600
rect 17880 18456 18599 18466
rect 16968 18432 17026 18442
rect 17712 18432 22114 18442
rect 16981 18408 16991 18418
rect 17016 18418 17026 18432
rect 17016 18408 22079 18418
rect 22104 18418 22114 18432
rect 22104 18408 23783 18418
rect 16752 18384 25319 18394
rect 16560 18360 26865 18370
rect 16176 18336 26889 18346
rect 16008 18312 29937 18322
rect 15264 18288 30009 18298
rect 14496 18264 14578 18274
rect 15048 18264 31522 18274
rect 9421 18240 9442 18250
rect 9469 18240 11183 18250
rect 14509 18240 14543 18250
rect 14568 18250 14578 18264
rect 14568 18240 18575 18250
rect 18613 18240 29961 18250
rect 30023 18240 31487 18250
rect 31512 18250 31522 18264
rect 31512 18240 33023 18250
rect 36648 18250 36658 18647
rect 36672 18277 36682 18647
rect 36696 18277 36706 18647
rect 36720 18274 36730 18647
rect 36744 18298 36754 18647
rect 36768 18322 36778 18647
rect 36792 18346 36802 18672
rect 36816 18370 36826 18671
rect 36840 18394 36850 18671
rect 36864 18418 36874 18671
rect 36888 18442 36898 18671
rect 36912 18466 36922 18671
rect 36936 18490 36946 18671
rect 36960 18514 36970 18696
rect 36960 18504 37847 18514
rect 36936 18480 38183 18490
rect 36912 18456 38207 18466
rect 36888 18432 38231 18442
rect 36864 18408 38255 18418
rect 36840 18384 38279 18394
rect 36816 18360 38303 18370
rect 36792 18336 38327 18346
rect 36768 18312 38351 18322
rect 36744 18288 38399 18298
rect 36720 18264 38423 18274
rect 36648 18240 38519 18250
rect 5952 18216 10055 18226
rect 11544 18226 11554 18239
rect 10069 18216 11554 18226
rect 11616 18226 11626 18239
rect 11616 18216 36658 18226
rect 36648 18205 36658 18216
rect 36709 18216 38543 18226
rect 9384 18192 9407 18202
rect 6912 18085 6922 18191
rect 9384 18181 9394 18192
rect 9445 18192 11207 18202
rect 11544 18192 11663 18202
rect 11232 18178 11242 18191
rect 9421 18168 11242 18178
rect 11256 18178 11266 18191
rect 11544 18178 11554 18192
rect 13717 18192 34559 18202
rect 36672 18202 36682 18215
rect 36672 18192 38567 18202
rect 11256 18168 11554 18178
rect 11653 18168 38591 18178
rect 9373 18144 11279 18154
rect 11317 18144 11615 18154
rect 13525 18144 36095 18154
rect 36661 18144 38639 18154
rect 9349 18120 11327 18130
rect 11509 18120 11639 18130
rect 11664 18130 11674 18143
rect 11664 18120 38495 18130
rect 38533 18120 38674 18130
rect 11352 18106 11362 18119
rect 9325 18096 11362 18106
rect 11376 18082 11386 18119
rect 9301 18072 11386 18082
rect 11400 18082 11410 18119
rect 38664 18109 38674 18120
rect 11509 18096 11591 18106
rect 11629 18096 38626 18106
rect 11400 18072 11591 18082
rect 11653 18072 38519 18082
rect 38616 18082 38626 18096
rect 38616 18072 38698 18082
rect 5928 18048 10103 18058
rect 11437 18048 38626 18058
rect 9253 18024 10031 18034
rect 10080 18024 11567 18034
rect 5904 18000 9551 18010
rect 10080 18010 10090 18024
rect 11605 18024 38482 18034
rect 9661 18000 10090 18010
rect 6840 17976 10055 17986
rect 6840 16957 6850 17976
rect 10080 17986 10090 18000
rect 10117 18000 10173 18010
rect 10259 18000 11447 18010
rect 11485 18000 38458 18010
rect 10080 17976 10210 17986
rect 10056 17965 10066 17975
rect 10200 17965 10210 17976
rect 10224 17976 11495 17986
rect 10224 17965 10234 17976
rect 11533 17976 38386 17986
rect 6912 17722 6922 17951
rect 9240 17749 9250 17951
rect 9288 17892 9298 17951
rect 9312 17892 9322 17951
rect 9336 17892 9346 17951
rect 9360 17892 9370 17951
rect 9384 17892 9394 17951
rect 9408 17892 9418 17951
rect 9432 17892 9442 17951
rect 9456 17892 9466 17951
rect 9480 17892 9490 17951
rect 9504 17892 9514 17951
rect 9528 17892 9538 17951
rect 9552 17865 9562 17951
rect 9264 17855 9562 17865
rect 9264 17817 9274 17855
rect 9576 17841 9586 17951
rect 9565 17831 9586 17841
rect 9600 17820 9610 17951
rect 9624 17820 9634 17951
rect 9648 17820 9658 17951
rect 9672 17820 9682 17951
rect 9696 17820 9706 17951
rect 9720 17820 9730 17951
rect 9744 17820 9754 17951
rect 9768 17820 9778 17951
rect 9264 17807 9575 17817
rect 9469 17772 9791 17782
rect 38184 17761 38194 17951
rect 38208 17761 38218 17951
rect 38232 17761 38242 17951
rect 38256 17761 38266 17951
rect 38280 17761 38290 17951
rect 38304 17761 38314 17951
rect 38328 17761 38338 17951
rect 38352 17761 38362 17951
rect 38376 17761 38386 17976
rect 38400 17761 38410 17975
rect 38424 17761 38434 17975
rect 38448 17761 38458 18000
rect 38472 17761 38482 18024
rect 38496 17761 38506 18023
rect 38520 17761 38530 18023
rect 38544 17761 38554 18023
rect 9397 17748 9791 17758
rect 6912 17712 9791 17722
rect 38568 17734 38578 18023
rect 38592 17986 38602 18023
rect 38616 18013 38626 18048
rect 38640 18010 38650 18047
rect 38688 18034 38698 18072
rect 40848 18058 40858 26279
rect 40765 18048 40858 18058
rect 38688 18024 40799 18034
rect 38640 18000 40823 18010
rect 38592 17976 40858 17986
rect 38173 17724 38578 17734
rect 38173 17700 38543 17710
rect 9240 16957 9250 17687
rect 9288 16957 9298 17687
rect 9312 16957 9322 17687
rect 9336 16957 9346 17687
rect 9360 16957 9370 17687
rect 9408 16957 9418 17687
rect 9432 16957 9442 17687
rect 9480 16957 9490 17687
rect 9504 16957 9514 17687
rect 9528 16957 9538 17687
rect 9552 16957 9562 17687
rect 9576 16957 9586 17687
rect 9600 16957 9610 17687
rect 9624 16957 9634 17687
rect 9648 16930 9658 17687
rect 5828 16920 9658 16930
rect 5880 13229 5890 16895
rect 6840 13261 6850 16895
rect 9240 13261 9250 16895
rect 9288 13261 9298 16895
rect 9312 13261 9322 16895
rect 9336 13261 9346 16895
rect 9360 13261 9370 16895
rect 9408 13261 9418 16895
rect 9432 13261 9442 16895
rect 9480 13261 9490 16895
rect 9504 13261 9514 16895
rect 9528 13261 9538 16895
rect 9552 13261 9562 16895
rect 9576 13306 9586 16895
rect 9600 13333 9610 16895
rect 9624 13333 9634 16895
rect 9672 13357 9682 17687
rect 9696 13357 9706 17687
rect 9720 13357 9730 17687
rect 9744 13330 9754 17687
rect 9661 13320 9754 13330
rect 9576 13296 9743 13306
rect 9768 13282 9778 17687
rect 38173 17676 38351 17686
rect 38173 17652 38303 17662
rect 38424 17638 38434 17675
rect 38173 17628 38434 17638
rect 38448 17617 38458 17675
rect 38472 17617 38482 17675
rect 38496 17617 38506 17675
rect 38520 17617 38530 17675
rect 38616 17617 38626 17951
rect 38173 17604 38399 17614
rect 38664 17590 38674 17951
rect 38173 17580 38674 17590
rect 9576 13272 9778 13282
rect 9576 13261 9586 13272
rect 9757 13243 9791 13253
rect 5880 13219 9791 13229
rect 5828 12192 5890 12202
rect 5880 8962 5890 12192
rect 6840 8989 6850 13190
rect 9240 8989 9250 13195
rect 9288 8989 9298 13195
rect 9312 8989 9322 13195
rect 9336 8989 9346 13195
rect 9360 13181 9370 13195
rect 9757 13195 9791 13205
rect 9360 13171 9791 13181
rect 9408 8989 9418 13140
rect 9432 9178 9442 13140
rect 9480 9226 9490 13140
rect 9504 9253 9514 13140
rect 9528 9253 9538 13140
rect 9552 9253 9562 13140
rect 9576 9253 9586 13140
rect 9600 9253 9610 13140
rect 9624 9253 9634 13140
rect 9648 9253 9658 13140
rect 9672 9253 9682 13140
rect 9696 9253 9706 13140
rect 9720 9253 9730 13140
rect 9744 9253 9754 13140
rect 9768 9253 9778 13171
rect 38184 11677 38194 17555
rect 38208 11677 38218 17555
rect 38232 16786 38242 17555
rect 38256 16813 38266 17555
rect 38280 16813 38290 17555
rect 38328 16813 38338 17555
rect 38376 16813 38386 17555
rect 38448 16813 38458 17555
rect 38472 16813 38482 17555
rect 38496 16813 38506 17555
rect 38520 16813 38530 17555
rect 38616 16813 38626 17555
rect 40752 16978 40762 17951
rect 40800 17002 40810 17951
rect 40824 17005 40834 17951
rect 40848 17005 40858 17976
rect 40789 16992 40810 17002
rect 40752 16968 40916 16978
rect 40800 16957 40810 16968
rect 40776 16930 40786 16943
rect 40776 16920 40916 16930
rect 40800 16813 40810 16895
rect 40824 16813 40834 16895
rect 40848 16813 40858 16895
rect 38232 16776 40916 16786
rect 38256 11650 38266 16751
rect 38173 11640 38266 11650
rect 38184 11144 38194 11615
rect 38208 11144 38218 11615
rect 38280 11144 38290 16751
rect 38328 11144 38338 16751
rect 38376 11144 38386 16751
rect 38448 11144 38458 16751
rect 38472 11144 38482 16751
rect 38496 11144 38506 16751
rect 38520 11117 38530 16751
rect 38173 11107 38530 11117
rect 38173 11083 38495 11093
rect 38184 9301 38194 11058
rect 38208 9301 38218 11058
rect 38280 9301 38290 11058
rect 38328 9301 38338 11058
rect 38376 9276 38386 11058
rect 38173 9266 38386 9276
rect 38173 9243 38207 9253
rect 9480 9216 9791 9226
rect 38448 9229 38458 11058
rect 38173 9219 38458 9229
rect 9565 9192 9791 9202
rect 38472 9205 38482 11058
rect 38173 9195 38482 9205
rect 9432 9168 9791 9178
rect 38616 9181 38626 16751
rect 40800 12298 40810 16751
rect 40824 12301 40834 16751
rect 40776 12288 40810 12298
rect 40776 12250 40786 12288
rect 40848 12274 40858 16751
rect 40813 12264 40858 12274
rect 40776 12240 40916 12250
rect 40776 12226 40786 12240
rect 40776 12216 40847 12226
rect 40813 12192 40916 12202
rect 40824 12058 40834 12167
rect 40848 12085 40858 12167
rect 40824 12048 40916 12058
rect 38173 9171 38626 9181
rect 9541 9144 9791 9154
rect 38173 9147 38279 9157
rect 9504 8989 9514 9143
rect 9576 9082 9586 9119
rect 9576 9072 9791 9082
rect 10222 9082 10232 9095
rect 9912 9072 10232 9082
rect 9661 9048 9815 9058
rect 9600 8989 9610 9047
rect 9624 8989 9634 9047
rect 9733 9024 9839 9034
rect 9672 8986 9682 9023
rect 9696 9010 9706 9023
rect 9696 9000 9863 9010
rect 9672 8976 9887 8986
rect 9912 8962 9922 9072
rect 10246 9058 10256 9095
rect 5880 8952 9922 8962
rect 9936 9048 10256 9058
rect 9637 8928 9922 8938
rect 6840 7501 6850 8927
rect 9240 7501 9250 8927
rect 9288 7501 9298 8927
rect 9312 7501 9322 8927
rect 9336 7501 9346 8927
rect 9408 7501 9418 8927
rect 9504 7501 9514 8927
rect 9600 8890 9610 8927
rect 9912 8917 9922 8928
rect 9936 8917 9946 9048
rect 9960 9024 10173 9034
rect 9960 8890 9970 9024
rect 9600 8880 9970 8890
rect 9936 8842 9946 8855
rect 9720 8832 9946 8842
rect 9720 7474 9730 8832
rect 5828 7464 9730 7474
rect 6840 6565 6850 7439
rect 9240 6586 9250 7439
rect 9288 6634 9298 7439
rect 9312 6706 9322 7439
rect 9336 6733 9346 7439
rect 9408 6733 9418 7439
rect 9504 6733 9514 7439
rect 9744 6733 9754 8807
rect 9768 6733 9778 8807
rect 9792 6733 9802 8807
rect 9816 6733 9826 8807
rect 9840 6730 9850 8807
rect 9864 6754 9874 8807
rect 9888 6778 9898 8807
rect 9912 6802 9922 8807
rect 38184 7474 38194 9119
rect 38328 7501 38338 9143
rect 40848 7522 40858 12023
rect 40848 7512 40916 7522
rect 38184 7464 40916 7474
rect 38328 7330 38338 7439
rect 38328 7320 40916 7330
rect 9912 6792 10943 6802
rect 9888 6768 11087 6778
rect 9864 6744 15047 6754
rect 9840 6720 15215 6730
rect 9312 6696 19199 6706
rect 9829 6672 15191 6682
rect 15229 6672 19319 6682
rect 9768 6658 9778 6671
rect 9768 6648 11111 6658
rect 11125 6648 15239 6658
rect 15253 6648 19367 6658
rect 19381 6648 27455 6658
rect 9288 6624 9767 6634
rect 9805 6624 27610 6634
rect 9421 6600 27575 6610
rect 27600 6610 27610 6624
rect 27600 6600 31559 6610
rect 9240 6576 11063 6586
rect 11101 6576 31727 6586
rect 9349 6552 35687 6562
rect 6816 6528 9743 6538
rect 6816 6514 6826 6528
rect 9781 6528 31703 6538
rect 31741 6528 35831 6538
rect 6792 6504 6826 6514
rect 6792 6450 6802 6504
rect 6853 6504 6898 6514
rect 6840 6450 6850 6503
rect 6888 6450 6898 6504
rect 9517 6504 10930 6514
rect 10920 6450 10930 6504
rect 10957 6504 19186 6514
rect 11064 6450 11074 6479
rect 11112 6450 11122 6479
rect 15048 6450 15058 6479
rect 15192 6450 15202 6479
rect 15240 6450 15250 6479
rect 19176 6450 19186 6504
rect 19213 6504 27442 6514
rect 19320 6450 19330 6479
rect 19368 6450 19378 6479
rect 27432 6450 27442 6504
rect 27469 6504 35890 6514
rect 27576 6450 27586 6479
rect 27624 6450 27634 6504
rect 31560 6450 31570 6479
rect 31704 6450 31714 6479
rect 31752 6450 31762 6504
rect 35688 6450 35698 6479
rect 35832 6450 35842 6479
rect 35880 6450 35890 6504
<< m2contact >>
rect 14975 41423 14989 41437
rect 15023 41423 15037 41437
rect 19103 41423 19117 41437
rect 19151 41423 19165 41437
rect 19295 41423 19309 41437
rect 27359 41423 27373 41437
rect 27407 41423 27421 41437
rect 31487 41423 31501 41437
rect 31535 41423 31549 41437
rect 27575 41399 27589 41413
rect 35615 41423 35629 41437
rect 35807 41423 35821 41437
rect 31703 41399 31717 41413
rect 35639 41399 35653 41413
rect 35663 41399 35677 41413
rect 27407 41375 27421 41389
rect 27431 41375 27445 41389
rect 31487 41375 31501 41389
rect 35615 41375 35629 41389
rect 15023 41351 15037 41365
rect 15047 41351 15061 41365
rect 35663 41351 35677 41365
rect 35807 41375 35821 41389
rect 11471 41327 11485 41341
rect 11495 41327 11509 41341
rect 11519 41327 11533 41341
rect 11543 41327 11557 41341
rect 31535 41327 31549 41341
rect 31703 41327 31717 41341
rect 35639 41327 35653 41341
rect 10895 41279 10909 41293
rect 11447 41279 11461 41293
rect 11567 41279 11581 41293
rect 19151 41279 19165 41293
rect 19175 41279 19189 41293
rect 27575 41279 27589 41293
rect 10895 41231 10909 41245
rect 5903 40391 5917 40405
rect 6815 40391 6829 40405
rect 6911 40391 6925 40405
rect 10895 40391 10909 40405
rect 14975 41255 14989 41269
rect 14999 41255 15013 41269
rect 19103 41255 19117 41269
rect 27359 41255 27373 41269
rect 27431 41255 27445 41269
rect 11447 41231 11461 41245
rect 11471 41231 11485 41245
rect 11495 41231 11509 41245
rect 11519 41231 11533 41245
rect 11543 41231 11557 41245
rect 11567 41231 11581 41245
rect 5903 40343 5917 40357
rect 6815 40343 6829 40357
rect 6911 40343 6925 40357
rect 10895 40343 10909 40357
rect 11423 39983 11437 39997
rect 11399 39959 11413 39973
rect 19295 41231 19309 41245
rect 19175 41207 19189 41221
rect 15047 41183 15061 41197
rect 14999 41159 15013 41173
rect 14975 41135 14989 41149
rect 11495 39959 11509 39973
rect 11519 39959 11533 39973
rect 11543 39959 11557 39973
rect 11567 39959 11581 39973
rect 11591 39959 11605 39973
rect 11615 39959 11629 39973
rect 11639 39959 11653 39973
rect 11663 39959 11677 39973
rect 11375 39935 11389 39949
rect 11279 39887 11293 39901
rect 11495 39911 11509 39925
rect 11375 39887 11389 39901
rect 11255 39863 11269 39877
rect 11711 39887 11725 39901
rect 11447 39863 11461 39877
rect 11471 39863 11485 39877
rect 11279 39839 11293 39853
rect 11303 39839 11317 39853
rect 11663 39815 11677 39829
rect 11711 39839 11725 39853
rect 6911 39791 6925 39805
rect 10895 39791 10909 39805
rect 11231 39791 11245 39805
rect 11279 39791 11293 39805
rect 11327 39791 11341 39805
rect 11663 39791 11677 39805
rect 11687 39791 11701 39805
rect 27119 39935 27133 39949
rect 26399 39911 26413 39925
rect 28967 39911 28981 39925
rect 26135 39887 26149 39901
rect 29135 39887 29149 39901
rect 29279 39887 29293 39901
rect 40847 40607 40861 40621
rect 40847 40559 40861 40573
rect 40823 40463 40837 40477
rect 40847 40463 40861 40477
rect 14975 39863 14989 39877
rect 18143 39863 18157 39877
rect 29351 39863 29365 39877
rect 36503 39863 36517 39877
rect 36647 39863 36661 39877
rect 36671 39839 36685 39853
rect 11735 39815 11749 39829
rect 17111 39815 17125 39829
rect 29231 39815 29245 39829
rect 29255 39815 29269 39829
rect 29303 39815 29317 39829
rect 29327 39815 29341 39829
rect 36527 39815 36541 39829
rect 36647 39815 36661 39829
rect 36719 39815 36733 39829
rect 11759 39791 11773 39805
rect 16919 39791 16933 39805
rect 28943 39791 28957 39805
rect 28967 39791 28981 39805
rect 36647 39791 36661 39805
rect 36671 39791 36685 39805
rect 11711 39767 11725 39781
rect 11735 39767 11749 39781
rect 6911 39743 6925 39757
rect 10895 39743 10909 39757
rect 5903 35735 5917 35749
rect 5879 35663 5893 35677
rect 5879 35615 5893 35629
rect 5903 35615 5917 35629
rect 5879 30983 5893 30997
rect 5903 30983 5917 30997
rect 5927 30935 5941 30949
rect 5879 30887 5893 30901
rect 5903 30887 5917 30901
rect 5927 30887 5941 30901
rect 5879 26303 5893 26317
rect 5903 26303 5917 26317
rect 5927 26303 5941 26317
rect 5879 26255 5893 26269
rect 5903 26255 5917 26269
rect 5927 26255 5941 26269
rect 5879 21671 5893 21685
rect 5903 21671 5917 21685
rect 5927 21671 5941 21685
rect 5951 21671 5965 21685
rect 5879 21623 5893 21637
rect 5903 21623 5917 21637
rect 5927 21623 5941 21637
rect 5951 21623 5965 21637
rect 11303 39743 11317 39757
rect 11351 39743 11365 39757
rect 11735 39743 11749 39757
rect 11759 39743 11773 39757
rect 11207 39719 11221 39733
rect 11303 39719 11317 39733
rect 11759 39719 11773 39733
rect 15959 39743 15973 39757
rect 29255 39743 29269 39757
rect 29279 39743 29293 39757
rect 36671 39743 36685 39757
rect 36743 39767 36757 39781
rect 36767 39719 36781 39733
rect 36791 39719 36805 39733
rect 11159 39695 11173 39709
rect 11471 39695 11485 39709
rect 11495 39695 11509 39709
rect 40823 40415 40837 40429
rect 40847 40415 40861 40429
rect 11231 39671 11245 39685
rect 11375 39671 11389 39685
rect 12071 39671 12085 39685
rect 14975 39671 14989 39685
rect 15719 39671 15733 39685
rect 29327 39671 29341 39685
rect 29351 39671 29365 39685
rect 36695 39671 36709 39685
rect 36719 39671 36733 39685
rect 36839 39671 36853 39685
rect 11135 39623 11149 39637
rect 11111 39599 11125 39613
rect 11639 39647 11653 39661
rect 11663 39647 11677 39661
rect 11687 39647 11701 39661
rect 11711 39647 11725 39661
rect 11735 39647 11749 39661
rect 11759 39647 11773 39661
rect 12191 39647 12205 39661
rect 11615 39623 11629 39637
rect 11231 39599 11245 39613
rect 11471 39599 11485 39613
rect 11591 39599 11605 39613
rect 11087 39575 11101 39589
rect 11567 39575 11581 39589
rect 11663 39575 11677 39589
rect 29183 39623 29197 39637
rect 29231 39647 29245 39661
rect 36719 39647 36733 39661
rect 36743 39647 36757 39661
rect 36863 39647 36877 39661
rect 36503 39623 36517 39637
rect 36527 39623 36541 39637
rect 36743 39623 36757 39637
rect 36767 39623 36781 39637
rect 12047 39599 12061 39613
rect 12071 39599 12085 39613
rect 29279 39599 29293 39613
rect 29303 39599 29317 39613
rect 36815 39599 36829 39613
rect 36911 39599 36925 39613
rect 28919 39575 28933 39589
rect 28943 39575 28957 39589
rect 36767 39575 36781 39589
rect 36791 39575 36805 39589
rect 11063 39551 11077 39565
rect 11135 39551 11149 39565
rect 11183 39551 11197 39565
rect 36887 39551 36901 39565
rect 36935 39551 36949 39565
rect 11087 39527 11101 39541
rect 11135 39527 11149 39541
rect 11063 39503 11077 39517
rect 11543 39503 11557 39517
rect 11663 39503 11677 39517
rect 12191 39503 12205 39517
rect 29135 39503 29149 39517
rect 11111 39479 11125 39493
rect 11135 39479 11149 39493
rect 11159 39479 11173 39493
rect 11183 39479 11197 39493
rect 11207 39479 11221 39493
rect 11231 39479 11245 39493
rect 11255 39479 11269 39493
rect 11279 39479 11293 39493
rect 11303 39479 11317 39493
rect 11327 39479 11341 39493
rect 11351 39479 11365 39493
rect 11375 39479 11389 39493
rect 11399 39479 11413 39493
rect 11423 39479 11437 39493
rect 11447 39479 11461 39493
rect 11471 39479 11485 39493
rect 11495 39479 11509 39493
rect 11519 39479 11533 39493
rect 12167 39479 12181 39493
rect 29111 39479 29125 39493
rect 36647 39479 36661 39493
rect 36671 39479 36685 39493
rect 36695 39479 36709 39493
rect 36719 39479 36733 39493
rect 36743 39479 36757 39493
rect 36767 39479 36781 39493
rect 11039 36783 11053 36797
rect 11063 36783 11077 36797
rect 11087 36783 11101 36797
rect 11111 36783 11125 36797
rect 11135 36783 11149 36797
rect 11159 36783 11173 36797
rect 11183 36783 11197 36797
rect 11207 36783 11221 36797
rect 11231 36783 11245 36797
rect 11255 36783 11269 36797
rect 11279 36783 11293 36797
rect 11303 36783 11317 36797
rect 11327 36783 11341 36797
rect 11351 36783 11365 36797
rect 11375 36783 11389 36797
rect 11399 36783 11413 36797
rect 11423 36783 11437 36797
rect 11447 36783 11461 36797
rect 11495 36759 11509 36773
rect 11519 36759 11533 36773
rect 11471 36733 11485 36747
rect 11039 36671 11053 36685
rect 11063 36647 11077 36661
rect 11087 36647 11101 36661
rect 11111 36647 11125 36661
rect 11135 36647 11149 36661
rect 11159 36647 11173 36661
rect 11183 36647 11197 36661
rect 11207 36647 11221 36661
rect 11231 36647 11245 36661
rect 11255 36647 11269 36661
rect 11279 36647 11293 36661
rect 11303 36647 11317 36661
rect 11327 36647 11341 36661
rect 11351 36647 11365 36661
rect 11375 36647 11389 36661
rect 11399 36647 11413 36661
rect 11423 36647 11437 36661
rect 11447 36647 11461 36661
rect 11471 36647 11485 36661
rect 11495 36647 11509 36661
rect 11519 36647 11533 36661
rect 11063 35591 11077 35605
rect 11087 35591 11101 35605
rect 11111 35591 11125 35605
rect 11135 35591 11149 35605
rect 11159 35591 11173 35605
rect 11183 35591 11197 35605
rect 11207 35591 11221 35605
rect 11231 35591 11245 35605
rect 11255 35591 11269 35605
rect 11279 35591 11293 35605
rect 11303 35591 11317 35605
rect 11327 35591 11341 35605
rect 11351 35591 11365 35605
rect 11375 35591 11389 35605
rect 11423 35583 11437 35597
rect 11447 35583 11461 35597
rect 11471 35583 11485 35597
rect 11495 35583 11509 35597
rect 11519 35583 11533 35597
rect 11399 35543 11413 35557
rect 11063 35495 11077 35509
rect 11087 35471 11101 35485
rect 11111 35471 11125 35485
rect 11135 35471 11149 35485
rect 11159 35471 11173 35485
rect 11183 35471 11197 35485
rect 11207 35471 11221 35485
rect 11231 35471 11245 35485
rect 11255 35471 11269 35485
rect 11279 35471 11293 35485
rect 11303 35471 11317 35485
rect 11327 35471 11341 35485
rect 11351 35471 11365 35485
rect 11375 35471 11389 35485
rect 11399 35471 11413 35485
rect 11423 35471 11437 35485
rect 11447 35471 11461 35485
rect 11471 35471 11485 35485
rect 11495 35471 11509 35485
rect 11519 35471 11533 35485
rect 11087 34415 11101 34429
rect 11111 34415 11125 34429
rect 11135 34415 11149 34429
rect 11159 34415 11173 34429
rect 11183 34415 11197 34429
rect 11207 34415 11221 34429
rect 11255 34423 11269 34437
rect 11279 34423 11293 34437
rect 11303 34423 11317 34437
rect 11327 34423 11341 34437
rect 11351 34423 11365 34437
rect 11375 34423 11389 34437
rect 11399 34423 11413 34437
rect 11423 34423 11437 34437
rect 11447 34423 11461 34437
rect 11471 34423 11485 34437
rect 11495 34423 11509 34437
rect 11519 34423 11533 34437
rect 11231 34367 11245 34381
rect 11087 34319 11101 34333
rect 11111 34295 11125 34309
rect 11135 34295 11149 34309
rect 11159 34295 11173 34309
rect 11183 34295 11197 34309
rect 11207 34295 11221 34309
rect 11231 34295 11245 34309
rect 11255 34295 11269 34309
rect 11279 34295 11293 34309
rect 11303 34295 11317 34309
rect 11327 34295 11341 34309
rect 11351 34295 11365 34309
rect 11375 34295 11389 34309
rect 11399 34295 11413 34309
rect 11423 34295 11437 34309
rect 11447 34295 11461 34309
rect 11471 34295 11485 34309
rect 11495 34295 11509 34309
rect 11519 34295 11533 34309
rect 11111 33239 11125 33253
rect 11135 33239 11149 33253
rect 11159 33239 11173 33253
rect 11183 33239 11197 33253
rect 11207 33239 11221 33253
rect 11231 33239 11245 33253
rect 11255 33239 11269 33253
rect 11279 33239 11293 33253
rect 11303 33239 11317 33253
rect 11327 33239 11341 33253
rect 11351 33239 11365 33253
rect 11375 33239 11389 33253
rect 11399 33239 11413 33253
rect 11447 33215 11461 33229
rect 11471 33215 11485 33229
rect 11495 33215 11509 33229
rect 11519 33215 11533 33229
rect 11423 33193 11437 33207
rect 11111 33143 11125 33157
rect 11135 33119 11149 33133
rect 11159 33119 11173 33133
rect 11183 33119 11197 33133
rect 11207 33119 11221 33133
rect 11231 33119 11245 33133
rect 11255 33119 11269 33133
rect 11279 33119 11293 33133
rect 11303 33119 11317 33133
rect 11327 33119 11341 33133
rect 11351 33119 11365 33133
rect 11375 33119 11389 33133
rect 11399 33119 11413 33133
rect 11423 33119 11437 33133
rect 11447 33119 11461 33133
rect 11471 33119 11485 33133
rect 11495 33119 11509 33133
rect 11519 33119 11533 33133
rect 11135 32063 11149 32077
rect 11159 32063 11173 32077
rect 11183 32063 11197 32077
rect 11207 32063 11221 32077
rect 11231 32063 11245 32077
rect 11255 32063 11269 32077
rect 11279 32063 11293 32077
rect 11303 32063 11317 32077
rect 11327 32063 11341 32077
rect 11351 32063 11365 32077
rect 11375 32063 11389 32077
rect 11399 32063 11413 32077
rect 11423 32063 11437 32077
rect 11447 32063 11461 32077
rect 11471 32063 11485 32077
rect 11519 32039 11533 32053
rect 11495 32017 11509 32031
rect 11135 31967 11149 31981
rect 11159 31943 11173 31957
rect 11183 31943 11197 31957
rect 11207 31943 11221 31957
rect 11231 31943 11245 31957
rect 11255 31943 11269 31957
rect 11279 31943 11293 31957
rect 11303 31943 11317 31957
rect 11327 31943 11341 31957
rect 11351 31943 11365 31957
rect 11375 31943 11389 31957
rect 11399 31943 11413 31957
rect 11423 31943 11437 31957
rect 11447 31943 11461 31957
rect 11471 31943 11485 31957
rect 11495 31943 11509 31957
rect 11519 31943 11533 31957
rect 11159 30887 11173 30901
rect 11183 30887 11197 30901
rect 11207 30887 11221 30901
rect 11231 30887 11245 30901
rect 11255 30887 11269 30901
rect 11279 30887 11293 30901
rect 11303 30887 11317 30901
rect 11327 30887 11341 30901
rect 11351 30887 11365 30901
rect 11375 30887 11389 30901
rect 11399 30887 11413 30901
rect 11423 30887 11437 30901
rect 11471 30863 11485 30877
rect 11495 30863 11509 30877
rect 11519 30863 11533 30877
rect 11447 30841 11461 30855
rect 11159 30791 11173 30805
rect 11183 30767 11197 30781
rect 11207 30767 11221 30781
rect 11231 30767 11245 30781
rect 11255 30767 11269 30781
rect 11279 30767 11293 30781
rect 11303 30767 11317 30781
rect 11327 30767 11341 30781
rect 11351 30767 11365 30781
rect 11375 30767 11389 30781
rect 11399 30767 11413 30781
rect 11423 30767 11437 30781
rect 11447 30767 11461 30781
rect 11471 30767 11485 30781
rect 11495 30767 11509 30781
rect 11519 30767 11533 30781
rect 11183 29739 11197 29753
rect 11207 29739 11221 29753
rect 11231 29739 11245 29753
rect 11279 29715 11293 29729
rect 11303 29715 11317 29729
rect 11327 29715 11341 29729
rect 11351 29715 11365 29729
rect 11375 29715 11389 29729
rect 11399 29715 11413 29729
rect 11423 29715 11437 29729
rect 11447 29715 11461 29729
rect 11471 29715 11485 29729
rect 11495 29715 11509 29729
rect 11519 29715 11533 29729
rect 11255 29677 11269 29691
rect 11183 29615 11197 29629
rect 11207 29591 11221 29605
rect 11231 29591 11245 29605
rect 11255 29591 11269 29605
rect 11279 29591 11293 29605
rect 11303 29591 11317 29605
rect 11327 29591 11341 29605
rect 11351 29591 11365 29605
rect 11375 29591 11389 29605
rect 11399 29591 11413 29605
rect 11423 29591 11437 29605
rect 11447 29591 11461 29605
rect 11471 29591 11485 29605
rect 11495 29591 11509 29605
rect 11519 29591 11533 29605
rect 11207 28535 11221 28549
rect 11231 28535 11245 28549
rect 11255 28535 11269 28549
rect 11279 28535 11293 28549
rect 11303 28535 11317 28549
rect 11327 28535 11341 28549
rect 11351 28535 11365 28549
rect 11375 28535 11389 28549
rect 11399 28535 11413 28549
rect 11423 28535 11437 28549
rect 11447 28535 11461 28549
rect 11471 28535 11485 28549
rect 11495 28535 11509 28549
rect 11183 28514 11197 28528
rect 11159 28487 11173 28501
rect 11447 28487 11461 28501
rect 11519 28490 11533 28504
rect 11303 28463 11317 28477
rect 11447 28463 11461 28477
rect 11159 28439 11173 28453
rect 11183 28439 11197 28453
rect 11207 28439 11221 28453
rect 11231 28439 11245 28453
rect 11255 28439 11269 28453
rect 11279 28439 11293 28453
rect 11135 27335 11149 27349
rect 11111 27311 11125 27325
rect 11327 28415 11341 28429
rect 11351 28415 11365 28429
rect 11375 28415 11389 28429
rect 11399 28415 11413 28429
rect 11423 28415 11437 28429
rect 11447 28415 11461 28429
rect 11471 28415 11485 28429
rect 11495 28415 11509 28429
rect 11519 28415 11533 28429
rect 11183 27311 11197 27325
rect 11207 27311 11221 27325
rect 11231 27311 11245 27325
rect 11255 27311 11269 27325
rect 11279 27311 11293 27325
rect 11303 27311 11317 27325
rect 11327 27311 11341 27325
rect 11351 27311 11365 27325
rect 11375 27311 11389 27325
rect 11399 27311 11413 27325
rect 11423 27311 11437 27325
rect 11447 27311 11461 27325
rect 11471 27311 11485 27325
rect 11495 27311 11509 27325
rect 11519 27311 11533 27325
rect 11111 27263 11125 27277
rect 11135 27263 11149 27277
rect 11183 27239 11197 27253
rect 11207 27239 11221 27253
rect 11231 27239 11245 27253
rect 11255 27239 11269 27253
rect 11279 27239 11293 27253
rect 11303 27239 11317 27253
rect 11327 27239 11341 27253
rect 11351 27239 11365 27253
rect 11375 27239 11389 27253
rect 11399 27239 11413 27253
rect 11423 27239 11437 27253
rect 11447 27239 11461 27253
rect 11471 27239 11485 27253
rect 11495 27239 11509 27253
rect 11519 27239 11533 27253
rect 11087 26159 11101 26173
rect 11111 26159 11125 26173
rect 11135 26159 11149 26173
rect 11159 26159 11173 26173
rect 11183 26159 11197 26173
rect 11207 26159 11221 26173
rect 11231 26159 11245 26173
rect 11255 26159 11269 26173
rect 11279 26159 11293 26173
rect 11303 26159 11317 26173
rect 11327 26159 11341 26173
rect 11351 26159 11365 26173
rect 11063 26135 11077 26149
rect 11399 26135 11413 26149
rect 11423 26135 11437 26149
rect 11447 26135 11461 26149
rect 11471 26135 11485 26149
rect 11495 26135 11509 26149
rect 11519 26135 11533 26149
rect 11351 26111 11365 26125
rect 11375 26111 11389 26125
rect 11063 26087 11077 26101
rect 11087 26087 11101 26101
rect 11111 26087 11125 26101
rect 11135 26087 11149 26101
rect 11159 26087 11173 26101
rect 11183 26087 11197 26101
rect 11207 26087 11221 26101
rect 11231 26087 11245 26101
rect 11255 26087 11269 26101
rect 11279 26087 11293 26101
rect 11303 26087 11317 26101
rect 11327 26087 11341 26101
rect 11039 24983 11053 24997
rect 11063 24983 11077 24997
rect 11087 24983 11101 24997
rect 11111 24983 11125 24997
rect 11135 24983 11149 24997
rect 11159 24983 11173 24997
rect 11183 24983 11197 24997
rect 11207 24983 11221 24997
rect 11231 24983 11245 24997
rect 11255 24983 11269 24997
rect 11279 24983 11293 24997
rect 11303 24983 11317 24997
rect 11375 26063 11389 26077
rect 11399 26063 11413 26077
rect 11423 26063 11437 26077
rect 11447 26063 11461 26077
rect 11471 26063 11485 26077
rect 11495 26063 11509 26077
rect 11519 26063 11533 26077
rect 11351 24959 11365 24973
rect 11375 24959 11389 24973
rect 11399 24959 11413 24973
rect 11423 24959 11437 24973
rect 11447 24959 11461 24973
rect 11471 24959 11485 24973
rect 11495 24959 11509 24973
rect 11519 24959 11533 24973
rect 11015 24935 11029 24949
rect 11327 24935 11341 24949
rect 10967 23807 10981 23821
rect 11015 24887 11029 24901
rect 11039 24887 11053 24901
rect 11063 24887 11077 24901
rect 11087 24887 11101 24901
rect 11111 24887 11125 24901
rect 11135 24887 11149 24901
rect 11159 24887 11173 24901
rect 11183 24887 11197 24901
rect 11207 24887 11221 24901
rect 11231 24887 11245 24901
rect 11255 24887 11269 24901
rect 11279 24887 11293 24901
rect 11303 24887 11317 24901
rect 11327 24887 11341 24901
rect 11351 24887 11365 24901
rect 11375 24887 11389 24901
rect 11399 24887 11413 24901
rect 11423 24887 11437 24901
rect 11447 24887 11461 24901
rect 11471 24887 11485 24901
rect 11495 24887 11509 24901
rect 11519 24887 11533 24901
rect 11015 23807 11029 23821
rect 11039 23807 11053 23821
rect 11063 23807 11077 23821
rect 11087 23807 11101 23821
rect 11111 23807 11125 23821
rect 11135 23807 11149 23821
rect 11159 23807 11173 23821
rect 11183 23807 11197 23821
rect 11207 23807 11221 23821
rect 11231 23807 11245 23821
rect 11255 23807 11269 23821
rect 11279 23807 11293 23821
rect 11303 23807 11317 23821
rect 11327 23807 11341 23821
rect 11351 23807 11365 23821
rect 11399 23783 11413 23797
rect 11423 23783 11437 23797
rect 11447 23783 11461 23797
rect 11471 23783 11485 23797
rect 11495 23783 11509 23797
rect 11519 23783 11533 23797
rect 10967 23759 10981 23773
rect 11015 23735 11029 23749
rect 11039 23735 11053 23749
rect 11063 23735 11077 23749
rect 11087 23735 11101 23749
rect 11111 23735 11125 23749
rect 11135 23735 11149 23749
rect 11159 23735 11173 23749
rect 11183 23735 11197 23749
rect 11207 23735 11221 23749
rect 11231 23735 11245 23749
rect 11255 23735 11269 23749
rect 11279 23735 11293 23749
rect 11303 23735 11317 23749
rect 11327 23735 11341 23749
rect 11351 23735 11365 23749
rect 10943 22631 10957 22645
rect 10967 22631 10981 22645
rect 10991 22631 11005 22645
rect 11015 22631 11029 22645
rect 11039 22631 11053 22645
rect 11063 22631 11077 22645
rect 11087 22631 11101 22645
rect 11111 22631 11125 22645
rect 11135 22631 11149 22645
rect 11159 22631 11173 22645
rect 11183 22631 11197 22645
rect 11207 22631 11221 22645
rect 11231 22631 11245 22645
rect 11255 22631 11269 22645
rect 11279 22631 11293 22645
rect 11303 22631 11317 22645
rect 11327 22631 11341 22645
rect 10895 22607 10909 22621
rect 10919 22607 10933 22621
rect 11399 23711 11413 23725
rect 11423 23711 11437 23725
rect 11447 23711 11461 23725
rect 11471 23711 11485 23725
rect 11495 23711 11509 23725
rect 11519 23711 11533 23725
rect 11375 22607 11389 22621
rect 11399 22607 11413 22621
rect 11423 22607 11437 22621
rect 11447 22607 11461 22621
rect 11471 22607 11485 22621
rect 11495 22607 11509 22621
rect 11519 22607 11533 22621
rect 11231 22583 11245 22597
rect 11351 22583 11365 22597
rect 10895 22559 10909 22573
rect 10919 22559 10933 22573
rect 10943 22559 10957 22573
rect 10967 22559 10981 22573
rect 10991 22559 11005 22573
rect 11015 22559 11029 22573
rect 11039 22559 11053 22573
rect 11063 22559 11077 22573
rect 11087 22559 11101 22573
rect 11111 22559 11125 22573
rect 11135 22559 11149 22573
rect 11159 22559 11173 22573
rect 11183 22559 11197 22573
rect 11207 22559 11221 22573
rect 10871 21455 10885 21469
rect 10895 21455 10909 21469
rect 10919 21455 10933 21469
rect 10943 21455 10957 21469
rect 10967 21455 10981 21469
rect 10847 21431 10861 21445
rect 11255 22535 11269 22549
rect 11279 22535 11293 22549
rect 11303 22535 11317 22549
rect 11327 22535 11341 22549
rect 11351 22535 11365 22549
rect 11375 22535 11389 22549
rect 11399 22535 11413 22549
rect 11423 22535 11437 22549
rect 11447 22535 11461 22549
rect 11471 22535 11485 22549
rect 11495 22535 11509 22549
rect 11519 22535 11533 22549
rect 11015 21431 11029 21445
rect 11039 21431 11053 21445
rect 11063 21431 11077 21445
rect 11087 21431 11101 21445
rect 11111 21431 11125 21445
rect 11135 21431 11149 21445
rect 11159 21431 11173 21445
rect 11183 21431 11197 21445
rect 11207 21431 11221 21445
rect 11231 21431 11245 21445
rect 11255 21431 11269 21445
rect 11279 21431 11293 21445
rect 11303 21431 11317 21445
rect 11327 21431 11341 21445
rect 11351 21431 11365 21445
rect 11375 21431 11389 21445
rect 11399 21431 11413 21445
rect 11423 21431 11437 21445
rect 11447 21431 11461 21445
rect 11471 21431 11485 21445
rect 11495 21431 11509 21445
rect 11519 21431 11533 21445
rect 10919 21407 10933 21421
rect 10991 21407 11005 21421
rect 10847 21383 10861 21397
rect 10871 21383 10885 21397
rect 10895 21383 10909 21397
rect 10943 21359 10957 21373
rect 10967 21359 10981 21373
rect 10991 21359 11005 21373
rect 11015 21359 11029 21373
rect 11039 21359 11053 21373
rect 11063 21359 11077 21373
rect 11087 21359 11101 21373
rect 11111 21359 11125 21373
rect 11135 21359 11149 21373
rect 11159 21359 11173 21373
rect 11183 21359 11197 21373
rect 11207 21359 11221 21373
rect 11231 21359 11245 21373
rect 11255 21359 11269 21373
rect 11279 21359 11293 21373
rect 11303 21359 11317 21373
rect 11327 21359 11341 21373
rect 11351 21359 11365 21373
rect 11375 21359 11389 21373
rect 11399 21359 11413 21373
rect 11423 21359 11437 21373
rect 11447 21359 11461 21373
rect 11471 21359 11485 21373
rect 11495 21359 11509 21373
rect 11519 21359 11533 21373
rect 10823 20279 10837 20293
rect 10847 20279 10861 20293
rect 10871 20279 10885 20293
rect 10895 20279 10909 20293
rect 10919 20279 10933 20293
rect 10799 20255 10813 20269
rect 10967 20255 10981 20269
rect 10991 20255 11005 20269
rect 11015 20255 11029 20269
rect 11039 20255 11053 20269
rect 11063 20255 11077 20269
rect 11087 20255 11101 20269
rect 11111 20255 11125 20269
rect 11135 20255 11149 20269
rect 11159 20255 11173 20269
rect 11183 20255 11197 20269
rect 11207 20255 11221 20269
rect 11231 20255 11245 20269
rect 11255 20255 11269 20269
rect 11279 20255 11293 20269
rect 11303 20255 11317 20269
rect 11327 20255 11341 20269
rect 11351 20255 11365 20269
rect 11375 20255 11389 20269
rect 11399 20255 11413 20269
rect 11423 20255 11437 20269
rect 11447 20255 11461 20269
rect 11471 20255 11485 20269
rect 11495 20255 11509 20269
rect 11519 20255 11533 20269
rect 10871 20231 10885 20245
rect 10943 20231 10957 20245
rect 10799 20207 10813 20221
rect 10823 20207 10837 20221
rect 10847 20207 10861 20221
rect 10895 20183 10909 20197
rect 10919 20183 10933 20197
rect 10943 20183 10957 20197
rect 10967 20183 10981 20197
rect 10991 20183 11005 20197
rect 11015 20183 11029 20197
rect 11039 20183 11053 20197
rect 11063 20183 11077 20197
rect 11087 20183 11101 20197
rect 11111 20183 11125 20197
rect 11135 20183 11149 20197
rect 11159 20183 11173 20197
rect 11183 20183 11197 20197
rect 11207 20183 11221 20197
rect 11231 20183 11245 20197
rect 11255 20183 11269 20197
rect 11279 20183 11293 20197
rect 11303 20183 11317 20197
rect 11327 20183 11341 20197
rect 11351 20183 11365 20197
rect 11375 20183 11389 20197
rect 11399 20183 11413 20197
rect 11423 20183 11437 20197
rect 11447 20183 11461 20197
rect 11471 20183 11485 20197
rect 11495 20183 11509 20197
rect 11519 20183 11533 20197
rect 10775 19103 10789 19117
rect 10799 19103 10813 19117
rect 10823 19103 10837 19117
rect 10847 19103 10861 19117
rect 10871 19103 10885 19117
rect 10895 19103 10909 19117
rect 10919 19103 10933 19117
rect 10943 19103 10957 19117
rect 10967 19103 10981 19117
rect 10991 19103 11005 19117
rect 11015 19103 11029 19117
rect 11039 19103 11053 19117
rect 11063 19103 11077 19117
rect 11087 19103 11101 19117
rect 10751 19079 10765 19093
rect 11135 19079 11149 19093
rect 11159 19079 11173 19093
rect 11183 19079 11197 19093
rect 11207 19079 11221 19093
rect 11231 19079 11245 19093
rect 11255 19079 11269 19093
rect 11279 19079 11293 19093
rect 11303 19079 11317 19093
rect 11327 19079 11341 19093
rect 11351 19079 11365 19093
rect 11375 19079 11389 19093
rect 11399 19079 11413 19093
rect 11423 19079 11437 19093
rect 11447 19079 11461 19093
rect 11471 19079 11485 19093
rect 11495 19079 11509 19093
rect 11519 19079 11533 19093
rect 10823 19055 10837 19069
rect 11111 19055 11125 19069
rect 10751 19031 10765 19045
rect 10775 19031 10789 19045
rect 10799 19031 10813 19045
rect 10847 19007 10861 19021
rect 10871 19007 10885 19021
rect 10895 19007 10909 19021
rect 10919 19007 10933 19021
rect 10943 19007 10957 19021
rect 10967 19007 10981 19021
rect 10991 19007 11005 19021
rect 11015 19007 11029 19021
rect 11039 19007 11053 19021
rect 11063 19007 11077 19021
rect 11087 19007 11101 19021
rect 11111 19007 11125 19021
rect 11135 19007 11149 19021
rect 11159 19007 11173 19021
rect 11183 19007 11197 19021
rect 11207 19007 11221 19021
rect 11231 19007 11245 19021
rect 11255 19007 11269 19021
rect 11279 19007 11293 19021
rect 11303 19007 11317 19021
rect 11327 19007 11341 19021
rect 11351 19007 11365 19021
rect 11375 19007 11389 19021
rect 11399 19007 11413 19021
rect 11423 19007 11437 19021
rect 11447 19007 11461 19021
rect 11471 19007 11485 19021
rect 11495 19007 11509 19021
rect 11519 19007 11533 19021
rect 10751 18839 10765 18853
rect 10775 18839 10789 18853
rect 10799 18839 10813 18853
rect 10823 18839 10837 18853
rect 10847 18839 10861 18853
rect 10871 18839 10885 18853
rect 10895 18839 10909 18853
rect 10919 18839 10933 18853
rect 10943 18839 10957 18853
rect 10967 18839 10981 18853
rect 10991 18839 11005 18853
rect 11015 18839 11029 18853
rect 11039 18839 11053 18853
rect 11063 18839 11077 18853
rect 11087 18839 11101 18853
rect 11111 18839 11125 18853
rect 11135 18839 11149 18853
rect 11159 18839 11173 18853
rect 11183 18839 11197 18853
rect 11207 18839 11221 18853
rect 11231 18839 11245 18853
rect 11255 18839 11269 18853
rect 11279 18839 11293 18853
rect 11303 18839 11317 18853
rect 11327 18839 11341 18853
rect 11351 18839 11365 18853
rect 11375 18839 11389 18853
rect 11399 18839 11413 18853
rect 11423 18839 11437 18853
rect 11447 18839 11461 18853
rect 11471 18839 11485 18853
rect 11495 18839 11509 18853
rect 11519 18839 11533 18853
rect 36647 18839 36661 18853
rect 36671 18839 36685 18853
rect 36695 18839 36709 18853
rect 36719 18839 36733 18853
rect 36743 18839 36757 18853
rect 36767 18839 36781 18853
rect 36815 39503 36829 39517
rect 36839 39503 36853 39517
rect 36863 39503 36877 39517
rect 36887 39503 36901 39517
rect 36911 39503 36925 39517
rect 36935 39503 36949 39517
rect 40847 35879 40861 35893
rect 40847 35831 40861 35845
rect 40847 35735 40861 35749
rect 40847 35687 40861 35701
rect 40847 31151 40861 31165
rect 40847 31103 40861 31117
rect 40847 31007 40861 31021
rect 40847 30959 40861 30973
rect 40847 26327 40861 26341
rect 40871 26303 40885 26317
rect 40847 26279 40861 26293
rect 36815 18863 36829 18877
rect 36839 18815 36853 18829
rect 36863 18815 36877 18829
rect 10751 18791 10765 18805
rect 10775 18767 10789 18781
rect 11447 18767 11461 18781
rect 36887 18767 36901 18781
rect 36911 18767 36925 18781
rect 11447 18743 11461 18757
rect 12234 18743 12248 18757
rect 12935 18743 12949 18757
rect 36167 18743 36181 18757
rect 36503 18743 36517 18757
rect 36791 18743 36805 18757
rect 36839 18743 36853 18757
rect 36839 18719 36853 18733
rect 36935 18719 36949 18733
rect 10799 18695 10813 18709
rect 11543 18695 11557 18709
rect 12047 18695 12061 18709
rect 12071 18695 12085 18709
rect 12210 18695 12224 18709
rect 14519 18695 14533 18709
rect 27719 18695 27733 18709
rect 27743 18695 27757 18709
rect 35423 18695 35437 18709
rect 36791 18695 36805 18709
rect 6911 18647 6925 18661
rect 11567 18647 11581 18661
rect 12186 18647 12200 18661
rect 12935 18647 12949 18661
rect 13511 18647 13525 18661
rect 13703 18647 13717 18661
rect 14495 18647 14509 18661
rect 14519 18647 14533 18661
rect 12162 18623 12176 18637
rect 6911 18599 6925 18613
rect 10895 18599 10909 18613
rect 10919 18599 10933 18613
rect 10943 18599 10957 18613
rect 10967 18599 10981 18613
rect 10991 18599 11005 18613
rect 11015 18599 11029 18613
rect 11039 18599 11053 18613
rect 11063 18599 11077 18613
rect 11087 18599 11101 18613
rect 11111 18599 11125 18613
rect 11135 18599 11149 18613
rect 11159 18599 11173 18613
rect 11183 18599 11197 18613
rect 11207 18599 11221 18613
rect 11231 18599 11245 18613
rect 11255 18599 11269 18613
rect 11279 18599 11293 18613
rect 11303 18599 11317 18613
rect 11327 18599 11341 18613
rect 11351 18599 11365 18613
rect 11375 18599 11389 18613
rect 11399 18599 11413 18613
rect 11423 18599 11437 18613
rect 11447 18599 11461 18613
rect 11471 18599 11485 18613
rect 11495 18599 11509 18613
rect 11519 18599 11533 18613
rect 11543 18599 11557 18613
rect 11567 18599 11581 18613
rect 10031 18527 10045 18541
rect 10823 18527 10837 18541
rect 10847 18527 10861 18541
rect 10871 18527 10885 18541
rect 9767 18503 9781 18517
rect 9743 18479 9757 18493
rect 9719 18455 9733 18469
rect 9695 18431 9709 18445
rect 9671 18407 9685 18421
rect 9623 18383 9637 18397
rect 9599 18359 9613 18373
rect 9575 18335 9589 18349
rect 9527 18311 9541 18325
rect 12071 18599 12085 18613
rect 11111 18335 11125 18349
rect 11135 18335 11149 18349
rect 11159 18335 11173 18349
rect 11183 18335 11197 18349
rect 11207 18335 11221 18349
rect 11231 18335 11245 18349
rect 11255 18335 11269 18349
rect 11279 18335 11293 18349
rect 11303 18335 11317 18349
rect 11327 18335 11341 18349
rect 11351 18335 11365 18349
rect 11375 18335 11389 18349
rect 11399 18335 11413 18349
rect 11423 18335 11437 18349
rect 11447 18335 11461 18349
rect 11471 18335 11485 18349
rect 11495 18335 11509 18349
rect 11519 18335 11533 18349
rect 11543 18335 11557 18349
rect 11567 18335 11581 18349
rect 11591 18335 11605 18349
rect 9503 18287 9517 18301
rect 11111 18287 11125 18301
rect 11135 18287 11149 18301
rect 11159 18287 11173 18301
rect 11615 18287 11629 18301
rect 6911 18239 6925 18253
rect 9407 18239 9421 18253
rect 9479 18263 9493 18277
rect 27743 18647 27757 18661
rect 36647 18647 36661 18661
rect 36671 18647 36685 18661
rect 36695 18647 36709 18661
rect 36719 18647 36733 18661
rect 36743 18647 36757 18661
rect 36767 18647 36781 18661
rect 15047 18623 15061 18637
rect 15263 18623 15277 18637
rect 16007 18623 16021 18637
rect 16175 18623 16189 18637
rect 16559 18623 16573 18637
rect 16751 18623 16765 18637
rect 16967 18623 16981 18637
rect 14519 18287 14533 18301
rect 14543 18287 14557 18301
rect 27479 18623 27493 18637
rect 17711 18599 17725 18613
rect 17879 18599 17893 18613
rect 16991 18455 17005 18469
rect 27287 18599 27301 18613
rect 18599 18455 18613 18469
rect 20687 18455 20701 18469
rect 16967 18407 16981 18421
rect 16991 18407 17005 18421
rect 22079 18407 22093 18421
rect 23783 18407 23797 18421
rect 25319 18383 25333 18397
rect 26865 18359 26879 18373
rect 26889 18335 26903 18349
rect 29937 18311 29951 18325
rect 30009 18287 30023 18301
rect 9455 18239 9469 18253
rect 11183 18239 11197 18253
rect 11543 18239 11557 18253
rect 11615 18239 11629 18253
rect 11639 18239 11653 18253
rect 12935 18239 12949 18253
rect 13511 18239 13525 18253
rect 13703 18239 13717 18253
rect 14495 18239 14509 18253
rect 14543 18239 14557 18253
rect 18575 18239 18589 18253
rect 18599 18239 18613 18253
rect 29961 18239 29975 18253
rect 30009 18239 30023 18253
rect 31487 18239 31501 18253
rect 33023 18239 33037 18253
rect 36671 18263 36685 18277
rect 36695 18263 36709 18277
rect 36815 18671 36829 18685
rect 36839 18671 36853 18685
rect 36863 18671 36877 18685
rect 36887 18671 36901 18685
rect 36911 18671 36925 18685
rect 36935 18671 36949 18685
rect 37847 18503 37861 18517
rect 38183 18479 38197 18493
rect 38207 18455 38221 18469
rect 38231 18431 38245 18445
rect 38255 18407 38269 18421
rect 38279 18383 38293 18397
rect 38303 18359 38317 18373
rect 38327 18335 38341 18349
rect 38351 18311 38365 18325
rect 38399 18287 38413 18301
rect 38423 18263 38437 18277
rect 38519 18239 38533 18253
rect 10055 18215 10069 18229
rect 36671 18215 36685 18229
rect 36695 18215 36709 18229
rect 38543 18215 38557 18229
rect 6911 18191 6925 18205
rect 9407 18191 9421 18205
rect 9431 18191 9445 18205
rect 11207 18191 11221 18205
rect 11231 18191 11245 18205
rect 11255 18191 11269 18205
rect 9383 18167 9397 18181
rect 9407 18167 9421 18181
rect 11663 18191 11677 18205
rect 13703 18191 13717 18205
rect 34559 18191 34573 18205
rect 36647 18191 36661 18205
rect 38567 18191 38581 18205
rect 11639 18167 11653 18181
rect 38591 18167 38605 18181
rect 9359 18143 9373 18157
rect 11279 18143 11293 18157
rect 11303 18143 11317 18157
rect 11615 18143 11629 18157
rect 11663 18143 11677 18157
rect 13511 18143 13525 18157
rect 36095 18143 36109 18157
rect 36647 18143 36661 18157
rect 38639 18143 38653 18157
rect 9335 18119 9349 18133
rect 11327 18119 11341 18133
rect 11351 18119 11365 18133
rect 11375 18119 11389 18133
rect 11399 18119 11413 18133
rect 11495 18119 11509 18133
rect 11639 18119 11653 18133
rect 38495 18119 38509 18133
rect 38519 18119 38533 18133
rect 9311 18095 9325 18109
rect 6911 18071 6925 18085
rect 9287 18071 9301 18085
rect 11495 18095 11509 18109
rect 11591 18095 11605 18109
rect 11615 18095 11629 18109
rect 11591 18071 11605 18085
rect 11639 18071 11653 18085
rect 38519 18071 38533 18085
rect 38663 18095 38677 18109
rect 10103 18047 10117 18061
rect 11423 18047 11437 18061
rect 9239 18023 9253 18037
rect 10031 18023 10045 18037
rect 9551 17999 9565 18013
rect 9647 17999 9661 18013
rect 11567 18023 11581 18037
rect 11591 18023 11605 18037
rect 10055 17975 10069 17989
rect 10103 17999 10117 18013
rect 10173 17999 10187 18013
rect 10245 17999 10259 18013
rect 11447 17999 11461 18013
rect 11471 17999 11485 18013
rect 11495 17975 11509 17989
rect 11519 17975 11533 17989
rect 6911 17951 6925 17965
rect 9239 17951 9253 17965
rect 9287 17951 9301 17965
rect 9311 17951 9325 17965
rect 9335 17951 9349 17965
rect 9359 17951 9373 17965
rect 9383 17951 9397 17965
rect 9407 17951 9421 17965
rect 9431 17951 9445 17965
rect 9455 17951 9469 17965
rect 9479 17951 9493 17965
rect 9503 17951 9517 17965
rect 9527 17951 9541 17965
rect 9551 17951 9565 17965
rect 9575 17951 9589 17965
rect 9599 17951 9613 17965
rect 9623 17951 9637 17965
rect 9647 17951 9661 17965
rect 9671 17951 9685 17965
rect 9695 17951 9709 17965
rect 9719 17951 9733 17965
rect 9743 17951 9757 17965
rect 9767 17951 9781 17965
rect 10055 17951 10069 17965
rect 10197 17951 10211 17965
rect 10221 17951 10235 17965
rect 38183 17951 38197 17965
rect 38207 17951 38221 17965
rect 38231 17951 38245 17965
rect 38255 17951 38269 17965
rect 38279 17951 38293 17965
rect 38303 17951 38317 17965
rect 38327 17951 38341 17965
rect 38351 17951 38365 17965
rect 9287 17878 9301 17892
rect 9311 17878 9325 17892
rect 9335 17878 9349 17892
rect 9359 17878 9373 17892
rect 9383 17878 9397 17892
rect 9407 17878 9421 17892
rect 9431 17878 9445 17892
rect 9455 17878 9469 17892
rect 9479 17878 9493 17892
rect 9503 17878 9517 17892
rect 9527 17878 9541 17892
rect 9551 17830 9565 17844
rect 9575 17806 9589 17820
rect 9599 17806 9613 17820
rect 9623 17806 9637 17820
rect 9647 17806 9661 17820
rect 9671 17806 9685 17820
rect 9695 17806 9709 17820
rect 9719 17806 9733 17820
rect 9743 17806 9757 17820
rect 9767 17806 9781 17820
rect 9455 17771 9469 17785
rect 9791 17771 9805 17785
rect 38399 17975 38413 17989
rect 38423 17975 38437 17989
rect 38495 18023 38509 18037
rect 38519 18023 38533 18037
rect 38543 18023 38557 18037
rect 38567 18023 38581 18037
rect 38591 18023 38605 18037
rect 9239 17735 9253 17749
rect 9383 17746 9397 17760
rect 9791 17747 9805 17761
rect 38183 17747 38197 17761
rect 38207 17747 38221 17761
rect 38231 17747 38245 17761
rect 38255 17747 38269 17761
rect 38279 17747 38293 17761
rect 38303 17747 38317 17761
rect 38327 17747 38341 17761
rect 38351 17747 38365 17761
rect 38375 17747 38389 17761
rect 38399 17747 38413 17761
rect 38423 17747 38437 17761
rect 38447 17747 38461 17761
rect 38471 17747 38485 17761
rect 38495 17747 38509 17761
rect 38519 17747 38533 17761
rect 38543 17747 38557 17761
rect 9791 17711 9805 17725
rect 38159 17723 38173 17737
rect 38639 18047 38653 18061
rect 38615 17999 38629 18013
rect 40751 18047 40765 18061
rect 40799 18023 40813 18037
rect 40823 17999 40837 18013
rect 38615 17951 38629 17965
rect 38663 17951 38677 17965
rect 40751 17951 40765 17965
rect 40799 17951 40813 17965
rect 40823 17951 40837 17965
rect 9239 17687 9253 17701
rect 9287 17687 9301 17701
rect 9311 17687 9325 17701
rect 9335 17687 9349 17701
rect 9359 17687 9373 17701
rect 9407 17687 9421 17701
rect 9431 17687 9445 17701
rect 9479 17687 9493 17701
rect 9503 17687 9517 17701
rect 9527 17687 9541 17701
rect 9551 17687 9565 17701
rect 9575 17687 9589 17701
rect 9599 17687 9613 17701
rect 9623 17687 9637 17701
rect 9647 17687 9661 17701
rect 9671 17687 9685 17701
rect 9695 17687 9709 17701
rect 9719 17687 9733 17701
rect 9743 17687 9757 17701
rect 9767 17687 9781 17701
rect 38159 17699 38173 17713
rect 38543 17699 38557 17713
rect 5879 16943 5893 16957
rect 6839 16943 6853 16957
rect 9239 16943 9253 16957
rect 9287 16943 9301 16957
rect 9311 16943 9325 16957
rect 9335 16943 9349 16957
rect 9359 16943 9373 16957
rect 9407 16943 9421 16957
rect 9431 16943 9445 16957
rect 9479 16943 9493 16957
rect 9503 16943 9517 16957
rect 9527 16943 9541 16957
rect 9551 16943 9565 16957
rect 9575 16943 9589 16957
rect 9599 16943 9613 16957
rect 9623 16943 9637 16957
rect 5879 16895 5893 16909
rect 6839 16895 6853 16909
rect 9239 16895 9253 16909
rect 9287 16895 9301 16909
rect 9311 16895 9325 16909
rect 9335 16895 9349 16909
rect 9359 16895 9373 16909
rect 9407 16895 9421 16909
rect 9431 16895 9445 16909
rect 9479 16895 9493 16909
rect 9503 16895 9517 16909
rect 9527 16895 9541 16909
rect 9551 16895 9565 16909
rect 9575 16895 9589 16909
rect 9599 16895 9613 16909
rect 9623 16895 9637 16909
rect 9671 13343 9685 13357
rect 9695 13343 9709 13357
rect 9719 13343 9733 13357
rect 9599 13319 9613 13333
rect 9623 13319 9637 13333
rect 9647 13319 9661 13333
rect 9743 13295 9757 13309
rect 38159 17675 38173 17689
rect 38351 17675 38365 17689
rect 38423 17675 38437 17689
rect 38447 17675 38461 17689
rect 38471 17675 38485 17689
rect 38495 17675 38509 17689
rect 38519 17675 38533 17689
rect 38159 17651 38173 17665
rect 38303 17651 38317 17665
rect 38159 17627 38173 17641
rect 38159 17603 38173 17617
rect 38399 17603 38413 17617
rect 38447 17603 38461 17617
rect 38471 17603 38485 17617
rect 38495 17603 38509 17617
rect 38519 17603 38533 17617
rect 38615 17603 38629 17617
rect 38159 17579 38173 17593
rect 38183 17555 38197 17569
rect 38207 17555 38221 17569
rect 38231 17555 38245 17569
rect 38255 17555 38269 17569
rect 38279 17555 38293 17569
rect 38327 17555 38341 17569
rect 38375 17555 38389 17569
rect 38447 17555 38461 17569
rect 38471 17555 38485 17569
rect 38495 17555 38509 17569
rect 38519 17555 38533 17569
rect 38615 17555 38629 17569
rect 6839 13247 6853 13261
rect 9239 13247 9253 13261
rect 9287 13247 9301 13261
rect 9311 13247 9325 13261
rect 9335 13247 9349 13261
rect 9359 13247 9373 13261
rect 9407 13247 9421 13261
rect 9431 13247 9445 13261
rect 9479 13247 9493 13261
rect 9503 13247 9517 13261
rect 9527 13247 9541 13261
rect 9551 13247 9565 13261
rect 9575 13247 9589 13261
rect 9743 13242 9757 13256
rect 9791 13242 9805 13256
rect 9791 13218 9805 13232
rect 6839 13190 6853 13204
rect 9239 13195 9253 13209
rect 9287 13195 9301 13209
rect 9311 13195 9325 13209
rect 9335 13195 9349 13209
rect 9359 13195 9373 13209
rect 9743 13194 9757 13208
rect 9791 13194 9805 13208
rect 9407 13140 9421 13154
rect 9431 13140 9445 13154
rect 9479 13140 9493 13154
rect 9503 13140 9517 13154
rect 9527 13140 9541 13154
rect 9551 13140 9565 13154
rect 9575 13140 9589 13154
rect 9599 13140 9613 13154
rect 9623 13140 9637 13154
rect 9647 13140 9661 13154
rect 9671 13140 9685 13154
rect 9695 13140 9709 13154
rect 9719 13140 9733 13154
rect 9743 13140 9757 13154
rect 9791 13170 9805 13184
rect 40775 16991 40789 17005
rect 40823 16991 40837 17005
rect 40847 16991 40861 17005
rect 40775 16943 40789 16957
rect 40799 16943 40813 16957
rect 40799 16895 40813 16909
rect 40823 16895 40837 16909
rect 40847 16895 40861 16909
rect 38255 16799 38269 16813
rect 38279 16799 38293 16813
rect 38327 16799 38341 16813
rect 38375 16799 38389 16813
rect 38447 16799 38461 16813
rect 38471 16799 38485 16813
rect 38495 16799 38509 16813
rect 38519 16799 38533 16813
rect 38615 16799 38629 16813
rect 40799 16799 40813 16813
rect 40823 16799 40837 16813
rect 40847 16799 40861 16813
rect 38255 16751 38269 16765
rect 38279 16751 38293 16765
rect 38327 16751 38341 16765
rect 38375 16751 38389 16765
rect 38447 16751 38461 16765
rect 38471 16751 38485 16765
rect 38495 16751 38509 16765
rect 38519 16751 38533 16765
rect 38615 16751 38629 16765
rect 40799 16751 40813 16765
rect 40823 16751 40837 16765
rect 40847 16751 40861 16765
rect 38183 11663 38197 11677
rect 38207 11663 38221 11677
rect 38159 11639 38173 11653
rect 38183 11615 38197 11629
rect 38207 11615 38221 11629
rect 38183 11130 38197 11144
rect 38207 11130 38221 11144
rect 38279 11130 38293 11144
rect 38327 11130 38341 11144
rect 38375 11130 38389 11144
rect 38447 11130 38461 11144
rect 38471 11130 38485 11144
rect 38495 11130 38509 11144
rect 38159 11106 38173 11120
rect 38159 11082 38173 11096
rect 38495 11082 38509 11096
rect 38183 11058 38197 11072
rect 38207 11058 38221 11072
rect 38279 11058 38293 11072
rect 38327 11058 38341 11072
rect 38375 11058 38389 11072
rect 38447 11058 38461 11072
rect 38471 11058 38485 11072
rect 38183 9287 38197 9301
rect 38207 9287 38221 9301
rect 38279 9287 38293 9301
rect 38327 9287 38341 9301
rect 38159 9265 38173 9279
rect 9503 9239 9517 9253
rect 9527 9239 9541 9253
rect 9551 9239 9565 9253
rect 9575 9239 9589 9253
rect 9599 9239 9613 9253
rect 9623 9239 9637 9253
rect 9647 9239 9661 9253
rect 9671 9239 9685 9253
rect 9695 9239 9709 9253
rect 9719 9239 9733 9253
rect 9743 9239 9757 9253
rect 9767 9239 9781 9253
rect 38159 9241 38173 9255
rect 38207 9242 38221 9256
rect 9791 9216 9805 9230
rect 38159 9217 38173 9231
rect 9551 9191 9565 9205
rect 9791 9192 9805 9206
rect 38159 9193 38173 9207
rect 9791 9168 9805 9182
rect 38159 9169 38173 9183
rect 40823 12287 40837 12301
rect 40799 12263 40813 12277
rect 40847 12215 40861 12229
rect 40799 12191 40813 12205
rect 40823 12167 40837 12181
rect 40847 12167 40861 12181
rect 40847 12071 40861 12085
rect 40847 12023 40861 12037
rect 9503 9143 9517 9157
rect 9527 9143 9541 9157
rect 9791 9144 9805 9158
rect 38159 9145 38173 9159
rect 38279 9146 38293 9160
rect 38327 9143 38341 9157
rect 9575 9119 9589 9133
rect 38183 9119 38197 9133
rect 10221 9095 10235 9109
rect 10245 9095 10259 9109
rect 9791 9071 9805 9085
rect 9599 9047 9613 9061
rect 9623 9047 9637 9061
rect 9647 9047 9661 9061
rect 9815 9047 9829 9061
rect 9671 9023 9685 9037
rect 9695 9023 9709 9037
rect 9719 9023 9733 9037
rect 9839 9023 9853 9037
rect 6839 8975 6853 8989
rect 9239 8975 9253 8989
rect 9287 8975 9301 8989
rect 9311 8975 9325 8989
rect 9335 8975 9349 8989
rect 9407 8975 9421 8989
rect 9503 8975 9517 8989
rect 9599 8975 9613 8989
rect 9623 8975 9637 8989
rect 9863 8999 9877 9013
rect 9887 8975 9901 8989
rect 6839 8927 6853 8941
rect 9239 8927 9253 8941
rect 9287 8927 9301 8941
rect 9311 8927 9325 8941
rect 9335 8927 9349 8941
rect 9407 8927 9421 8941
rect 9503 8927 9517 8941
rect 9599 8927 9613 8941
rect 9623 8927 9637 8941
rect 9911 8903 9925 8917
rect 9935 8903 9949 8917
rect 10173 9023 10187 9037
rect 9935 8855 9949 8869
rect 6839 7487 6853 7501
rect 9239 7487 9253 7501
rect 9287 7487 9301 7501
rect 9311 7487 9325 7501
rect 9335 7487 9349 7501
rect 9407 7487 9421 7501
rect 9503 7487 9517 7501
rect 9743 8807 9757 8821
rect 9767 8807 9781 8821
rect 9791 8807 9805 8821
rect 9815 8807 9829 8821
rect 9839 8807 9853 8821
rect 9863 8807 9877 8821
rect 9887 8807 9901 8821
rect 9911 8807 9925 8821
rect 6839 7439 6853 7453
rect 9239 7439 9253 7453
rect 9287 7439 9301 7453
rect 9311 7439 9325 7453
rect 9335 7439 9349 7453
rect 9407 7439 9421 7453
rect 9503 7439 9517 7453
rect 9335 6719 9349 6733
rect 9407 6719 9421 6733
rect 9503 6719 9517 6733
rect 9743 6719 9757 6733
rect 9767 6719 9781 6733
rect 9791 6719 9805 6733
rect 9815 6719 9829 6733
rect 38327 7487 38341 7501
rect 38327 7439 38341 7453
rect 10943 6791 10957 6805
rect 11087 6767 11101 6781
rect 15047 6743 15061 6757
rect 15215 6719 15229 6733
rect 19199 6695 19213 6709
rect 9767 6671 9781 6685
rect 9815 6671 9829 6685
rect 15191 6671 15205 6685
rect 15215 6671 15229 6685
rect 19319 6671 19333 6685
rect 11111 6647 11125 6661
rect 15239 6647 15253 6661
rect 19367 6647 19381 6661
rect 27455 6647 27469 6661
rect 9767 6623 9781 6637
rect 9791 6623 9805 6637
rect 9407 6599 9421 6613
rect 27575 6599 27589 6613
rect 31559 6599 31573 6613
rect 11063 6575 11077 6589
rect 11087 6575 11101 6589
rect 31727 6575 31741 6589
rect 6839 6551 6853 6565
rect 9335 6551 9349 6565
rect 35687 6551 35701 6565
rect 9743 6527 9757 6541
rect 9767 6527 9781 6541
rect 31703 6527 31717 6541
rect 31727 6527 31741 6541
rect 35831 6527 35845 6541
rect 6839 6503 6853 6517
rect 9503 6503 9517 6517
rect 10943 6503 10957 6517
rect 11063 6479 11077 6493
rect 11111 6479 11125 6493
rect 15047 6479 15061 6493
rect 15191 6479 15205 6493
rect 15239 6479 15253 6493
rect 19199 6503 19213 6517
rect 19319 6479 19333 6493
rect 19367 6479 19381 6493
rect 27455 6503 27469 6517
rect 27575 6479 27589 6493
rect 31559 6479 31573 6493
rect 31703 6479 31717 6493
rect 35687 6479 35701 6493
rect 35831 6479 35845 6493
<< metal2 >>
rect 10896 41245 10908 41279
rect 11448 41245 11460 41279
rect 11472 41245 11484 41327
rect 11496 41245 11508 41327
rect 11520 41245 11532 41327
rect 11544 41245 11556 41327
rect 11568 41245 11580 41279
rect 14976 41269 14988 41423
rect 15024 41365 15036 41423
rect 14976 41149 14988 41255
rect 15000 41173 15012 41255
rect 15048 41197 15060 41351
rect 19104 41269 19116 41423
rect 19152 41293 19164 41423
rect 19176 41221 19188 41279
rect 19296 41245 19308 41423
rect 27360 41269 27372 41423
rect 27408 41389 27420 41423
rect 27432 41269 27444 41375
rect 27576 41293 27588 41399
rect 31488 41389 31500 41423
rect 31536 41341 31548 41423
rect 31704 41341 31716 41399
rect 35616 41389 35628 41423
rect 35640 41341 35652 41399
rect 35664 41365 35676 41399
rect 35808 41389 35820 41423
rect 40848 40573 40860 40607
rect 40824 40429 40836 40463
rect 40848 40429 40860 40463
rect 5904 40357 5916 40391
rect 6816 40357 6828 40391
rect 6912 40357 6924 40391
rect 10896 40357 10908 40391
rect 11376 39901 11388 39935
rect 6912 39757 6924 39791
rect 10896 39757 10908 39791
rect 11064 39517 11076 39551
rect 11088 39541 11100 39575
rect 11112 39493 11124 39599
rect 11136 39565 11148 39623
rect 11136 39493 11148 39527
rect 11160 39493 11172 39695
rect 11184 39493 11196 39551
rect 11208 39493 11220 39719
rect 11232 39685 11244 39791
rect 11232 39493 11244 39599
rect 11256 39493 11268 39863
rect 11280 39853 11292 39887
rect 11280 39493 11292 39791
rect 11304 39757 11316 39839
rect 11304 39493 11316 39719
rect 11328 39493 11340 39791
rect 11352 39493 11364 39743
rect 11376 39493 11388 39671
rect 11400 39493 11412 39959
rect 11424 39493 11436 39983
rect 11496 39925 11508 39959
rect 11448 39493 11460 39863
rect 11472 39709 11484 39863
rect 11472 39493 11484 39599
rect 11496 39493 11508 39695
rect 11520 39493 11532 39959
rect 11544 39517 11556 39959
rect 11568 39589 11580 39959
rect 11592 39613 11604 39959
rect 11616 39637 11628 39959
rect 11640 39661 11652 39959
rect 11664 39829 11676 39959
rect 11712 39853 11724 39887
rect 11664 39661 11676 39791
rect 11688 39661 11700 39791
rect 11736 39781 11748 39815
rect 11712 39661 11724 39767
rect 11760 39757 11772 39791
rect 11736 39661 11748 39743
rect 11760 39661 11772 39719
rect 14976 39685 14988 39863
rect 12072 39613 12084 39671
rect 11664 39517 11676 39575
rect 12048 39456 12060 39599
rect 12192 39517 12204 39647
rect 12163 39479 12167 39493
rect 15720 39492 15732 39671
rect 15960 39492 15972 39743
rect 16920 39492 16932 39791
rect 17112 39492 17124 39815
rect 18144 39492 18156 39863
rect 26136 39492 26148 39887
rect 26400 39492 26412 39911
rect 27120 39492 27132 39935
rect 28968 39805 28980 39911
rect 28944 39589 28956 39791
rect 28920 39492 28932 39575
rect 29136 39517 29148 39887
rect 29232 39661 29244 39815
rect 29256 39757 29268 39815
rect 29280 39757 29292 39887
rect 15715 39480 15732 39492
rect 15955 39480 15972 39492
rect 16915 39480 16932 39492
rect 17107 39480 17124 39492
rect 18141 39480 18156 39492
rect 26132 39480 26148 39492
rect 26396 39480 26412 39492
rect 27116 39480 27132 39492
rect 28915 39480 28932 39492
rect 12163 39456 12175 39479
rect 15715 39456 15727 39480
rect 15955 39456 15967 39480
rect 16915 39456 16927 39480
rect 17107 39456 17119 39480
rect 18141 39456 18153 39480
rect 26132 39456 26144 39480
rect 26396 39456 26408 39480
rect 27116 39456 27128 39480
rect 28915 39456 28927 39480
rect 29107 39479 29111 39493
rect 29184 39492 29196 39623
rect 29304 39613 29316 39815
rect 29328 39685 29340 39815
rect 29352 39685 29364 39863
rect 36504 39637 36516 39863
rect 36648 39829 36660 39863
rect 36528 39637 36540 39815
rect 36672 39805 36684 39839
rect 29280 39492 29292 39599
rect 29179 39480 29196 39492
rect 29275 39480 29292 39492
rect 29107 39456 29119 39479
rect 29179 39456 29191 39480
rect 29275 39456 29287 39480
rect 36504 39456 36516 39623
rect 36648 39493 36660 39791
rect 36672 39493 36684 39743
rect 36720 39685 36732 39815
rect 36696 39493 36708 39671
rect 36744 39661 36756 39767
rect 36720 39493 36732 39647
rect 36768 39637 36780 39719
rect 36744 39493 36756 39623
rect 36792 39589 36804 39719
rect 36768 39493 36780 39575
rect 36816 39517 36828 39599
rect 36840 39517 36852 39671
rect 36864 39517 36876 39647
rect 36888 39517 36900 39551
rect 36912 39517 36924 39599
rect 36936 39517 36948 39551
rect 11040 36685 11052 36783
rect 11064 36661 11076 36783
rect 11088 36661 11100 36783
rect 11112 36661 11124 36783
rect 11136 36661 11148 36783
rect 11160 36661 11172 36783
rect 11184 36661 11196 36783
rect 11208 36661 11220 36783
rect 11232 36661 11244 36783
rect 11256 36661 11268 36783
rect 11280 36661 11292 36783
rect 11304 36661 11316 36783
rect 11328 36661 11340 36783
rect 11352 36661 11364 36783
rect 11376 36661 11388 36783
rect 11400 36661 11412 36783
rect 11424 36661 11436 36783
rect 11448 36661 11460 36783
rect 11472 36661 11484 36733
rect 11496 36661 11508 36759
rect 11520 36661 11532 36759
rect 40848 35845 40860 35879
rect 5880 35629 5892 35663
rect 5904 35629 5916 35735
rect 40848 35701 40860 35735
rect 11064 35509 11076 35591
rect 11088 35485 11100 35591
rect 11112 35485 11124 35591
rect 11136 35485 11148 35591
rect 11160 35485 11172 35591
rect 11184 35485 11196 35591
rect 11208 35485 11220 35591
rect 11232 35485 11244 35591
rect 11256 35485 11268 35591
rect 11280 35485 11292 35591
rect 11304 35485 11316 35591
rect 11328 35485 11340 35591
rect 11352 35485 11364 35591
rect 11376 35485 11388 35591
rect 11400 35485 11412 35543
rect 11424 35485 11436 35583
rect 11448 35485 11460 35583
rect 11472 35485 11484 35583
rect 11496 35485 11508 35583
rect 11520 35485 11532 35583
rect 11088 34333 11100 34415
rect 11112 34309 11124 34415
rect 11136 34309 11148 34415
rect 11160 34309 11172 34415
rect 11184 34309 11196 34415
rect 11208 34309 11220 34415
rect 11232 34309 11244 34367
rect 11256 34309 11268 34423
rect 11280 34309 11292 34423
rect 11304 34309 11316 34423
rect 11328 34309 11340 34423
rect 11352 34309 11364 34423
rect 11376 34309 11388 34423
rect 11400 34309 11412 34423
rect 11424 34309 11436 34423
rect 11448 34309 11460 34423
rect 11472 34309 11484 34423
rect 11496 34309 11508 34423
rect 11520 34309 11532 34423
rect 11112 33157 11124 33239
rect 11136 33133 11148 33239
rect 11160 33133 11172 33239
rect 11184 33133 11196 33239
rect 11208 33133 11220 33239
rect 11232 33133 11244 33239
rect 11256 33133 11268 33239
rect 11280 33133 11292 33239
rect 11304 33133 11316 33239
rect 11328 33133 11340 33239
rect 11352 33133 11364 33239
rect 11376 33133 11388 33239
rect 11400 33133 11412 33239
rect 11424 33133 11436 33193
rect 11448 33133 11460 33215
rect 11472 33133 11484 33215
rect 11496 33133 11508 33215
rect 11520 33133 11532 33215
rect 11136 31981 11148 32063
rect 11160 31957 11172 32063
rect 11184 31957 11196 32063
rect 11208 31957 11220 32063
rect 11232 31957 11244 32063
rect 11256 31957 11268 32063
rect 11280 31957 11292 32063
rect 11304 31957 11316 32063
rect 11328 31957 11340 32063
rect 11352 31957 11364 32063
rect 11376 31957 11388 32063
rect 11400 31957 11412 32063
rect 11424 31957 11436 32063
rect 11448 31957 11460 32063
rect 11472 31957 11484 32063
rect 11496 31957 11508 32017
rect 11520 31957 11532 32039
rect 40848 31117 40860 31151
rect 5880 30901 5892 30983
rect 5904 30901 5916 30983
rect 40848 30973 40860 31007
rect 5928 30901 5940 30935
rect 11160 30805 11172 30887
rect 11184 30781 11196 30887
rect 11208 30781 11220 30887
rect 11232 30781 11244 30887
rect 11256 30781 11268 30887
rect 11280 30781 11292 30887
rect 11304 30781 11316 30887
rect 11328 30781 11340 30887
rect 11352 30781 11364 30887
rect 11376 30781 11388 30887
rect 11400 30781 11412 30887
rect 11424 30781 11436 30887
rect 11448 30781 11460 30841
rect 11472 30781 11484 30863
rect 11496 30781 11508 30863
rect 11520 30781 11532 30863
rect 11184 29629 11196 29739
rect 11208 29605 11220 29739
rect 11232 29605 11244 29739
rect 11256 29605 11268 29677
rect 11280 29605 11292 29715
rect 11304 29605 11316 29715
rect 11328 29605 11340 29715
rect 11352 29605 11364 29715
rect 11376 29605 11388 29715
rect 11400 29605 11412 29715
rect 11424 29605 11436 29715
rect 11448 29605 11460 29715
rect 11472 29605 11484 29715
rect 11496 29605 11508 29715
rect 11520 29605 11532 29715
rect 11160 28453 11172 28487
rect 11184 28453 11196 28514
rect 11208 28453 11220 28535
rect 11232 28453 11244 28535
rect 11256 28453 11268 28535
rect 11280 28453 11292 28535
rect 11304 28477 11316 28535
rect 11328 28429 11340 28535
rect 11352 28429 11364 28535
rect 11376 28429 11388 28535
rect 11400 28429 11412 28535
rect 11424 28429 11436 28535
rect 11448 28501 11460 28535
rect 11448 28429 11460 28463
rect 11472 28429 11484 28535
rect 11496 28429 11508 28535
rect 11520 28429 11532 28490
rect 11112 27277 11124 27311
rect 11136 27277 11148 27335
rect 11184 27253 11196 27311
rect 11208 27253 11220 27311
rect 11232 27253 11244 27311
rect 11256 27253 11268 27311
rect 11280 27253 11292 27311
rect 11304 27253 11316 27311
rect 11328 27253 11340 27311
rect 11352 27253 11364 27311
rect 11376 27253 11388 27311
rect 11400 27253 11412 27311
rect 11424 27253 11436 27311
rect 11448 27253 11460 27311
rect 11472 27253 11484 27311
rect 11496 27253 11508 27311
rect 11520 27253 11532 27311
rect 5880 26269 5892 26303
rect 5904 26269 5916 26303
rect 5928 26269 5940 26303
rect 40848 26293 40860 26327
rect 40885 26304 40916 26316
rect 11064 26101 11076 26135
rect 11088 26101 11100 26159
rect 11112 26101 11124 26159
rect 11136 26101 11148 26159
rect 11160 26101 11172 26159
rect 11184 26101 11196 26159
rect 11208 26101 11220 26159
rect 11232 26101 11244 26159
rect 11256 26101 11268 26159
rect 11280 26101 11292 26159
rect 11304 26101 11316 26159
rect 11328 26101 11340 26159
rect 11352 26125 11364 26159
rect 11376 26077 11388 26111
rect 11400 26077 11412 26135
rect 11424 26077 11436 26135
rect 11448 26077 11460 26135
rect 11472 26077 11484 26135
rect 11496 26077 11508 26135
rect 11520 26077 11532 26135
rect 11016 24901 11028 24935
rect 11040 24901 11052 24983
rect 11064 24901 11076 24983
rect 11088 24901 11100 24983
rect 11112 24901 11124 24983
rect 11136 24901 11148 24983
rect 11160 24901 11172 24983
rect 11184 24901 11196 24983
rect 11208 24901 11220 24983
rect 11232 24901 11244 24983
rect 11256 24901 11268 24983
rect 11280 24901 11292 24983
rect 11304 24901 11316 24983
rect 11328 24901 11340 24935
rect 11352 24901 11364 24959
rect 11376 24901 11388 24959
rect 11400 24901 11412 24959
rect 11424 24901 11436 24959
rect 11448 24901 11460 24959
rect 11472 24901 11484 24959
rect 11496 24901 11508 24959
rect 11520 24901 11532 24959
rect 10968 23773 10980 23807
rect 11016 23749 11028 23807
rect 11040 23749 11052 23807
rect 11064 23749 11076 23807
rect 11088 23749 11100 23807
rect 11112 23749 11124 23807
rect 11136 23749 11148 23807
rect 11160 23749 11172 23807
rect 11184 23749 11196 23807
rect 11208 23749 11220 23807
rect 11232 23749 11244 23807
rect 11256 23749 11268 23807
rect 11280 23749 11292 23807
rect 11304 23749 11316 23807
rect 11328 23749 11340 23807
rect 11352 23749 11364 23807
rect 11400 23725 11412 23783
rect 11424 23725 11436 23783
rect 11448 23725 11460 23783
rect 11472 23725 11484 23783
rect 11496 23725 11508 23783
rect 11520 23725 11532 23783
rect 10896 22573 10908 22607
rect 10920 22573 10932 22607
rect 10944 22573 10956 22631
rect 10968 22573 10980 22631
rect 10992 22573 11004 22631
rect 11016 22573 11028 22631
rect 11040 22573 11052 22631
rect 11064 22573 11076 22631
rect 11088 22573 11100 22631
rect 11112 22573 11124 22631
rect 11136 22573 11148 22631
rect 11160 22573 11172 22631
rect 11184 22573 11196 22631
rect 11208 22573 11220 22631
rect 11232 22597 11244 22631
rect 11256 22549 11268 22631
rect 11280 22549 11292 22631
rect 11304 22549 11316 22631
rect 11328 22549 11340 22631
rect 11352 22549 11364 22583
rect 11376 22549 11388 22607
rect 11400 22549 11412 22607
rect 11424 22549 11436 22607
rect 11448 22549 11460 22607
rect 11472 22549 11484 22607
rect 11496 22549 11508 22607
rect 11520 22549 11532 22607
rect 5880 21637 5892 21671
rect 5904 21637 5916 21671
rect 5928 21637 5940 21671
rect 5952 21637 5964 21671
rect 10848 21397 10860 21431
rect 10872 21397 10884 21455
rect 10896 21397 10908 21455
rect 10920 21421 10932 21455
rect 10944 21373 10956 21455
rect 10968 21373 10980 21455
rect 10992 21373 11004 21407
rect 11016 21373 11028 21431
rect 11040 21373 11052 21431
rect 11064 21373 11076 21431
rect 11088 21373 11100 21431
rect 11112 21373 11124 21431
rect 11136 21373 11148 21431
rect 11160 21373 11172 21431
rect 11184 21373 11196 21431
rect 11208 21373 11220 21431
rect 11232 21373 11244 21431
rect 11256 21373 11268 21431
rect 11280 21373 11292 21431
rect 11304 21373 11316 21431
rect 11328 21373 11340 21431
rect 11352 21373 11364 21431
rect 11376 21373 11388 21431
rect 11400 21373 11412 21431
rect 11424 21373 11436 21431
rect 11448 21373 11460 21431
rect 11472 21373 11484 21431
rect 11496 21373 11508 21431
rect 11520 21373 11532 21431
rect 10800 20221 10812 20255
rect 10824 20221 10836 20279
rect 10848 20221 10860 20279
rect 10872 20245 10884 20279
rect 10896 20197 10908 20279
rect 10920 20197 10932 20279
rect 10944 20197 10956 20231
rect 10968 20197 10980 20255
rect 10992 20197 11004 20255
rect 11016 20197 11028 20255
rect 11040 20197 11052 20255
rect 11064 20197 11076 20255
rect 11088 20197 11100 20255
rect 11112 20197 11124 20255
rect 11136 20197 11148 20255
rect 11160 20197 11172 20255
rect 11184 20197 11196 20255
rect 11208 20197 11220 20255
rect 11232 20197 11244 20255
rect 11256 20197 11268 20255
rect 11280 20197 11292 20255
rect 11304 20197 11316 20255
rect 11328 20197 11340 20255
rect 11352 20197 11364 20255
rect 11376 20197 11388 20255
rect 11400 20197 11412 20255
rect 11424 20197 11436 20255
rect 11448 20197 11460 20255
rect 11472 20197 11484 20255
rect 11496 20197 11508 20255
rect 11520 20197 11532 20255
rect 10752 19045 10764 19079
rect 10776 19045 10788 19103
rect 10800 19045 10812 19103
rect 10824 19069 10836 19103
rect 10848 19021 10860 19103
rect 10872 19021 10884 19103
rect 10896 19021 10908 19103
rect 10920 19021 10932 19103
rect 10944 19021 10956 19103
rect 10968 19021 10980 19103
rect 10992 19021 11004 19103
rect 11016 19021 11028 19103
rect 11040 19021 11052 19103
rect 11064 19021 11076 19103
rect 11088 19021 11100 19103
rect 11112 19021 11124 19055
rect 11136 19021 11148 19079
rect 11160 19021 11172 19079
rect 11184 19021 11196 19079
rect 11208 19021 11220 19079
rect 11232 19021 11244 19079
rect 11256 19021 11268 19079
rect 11280 19021 11292 19079
rect 11304 19021 11316 19079
rect 11328 19021 11340 19079
rect 11352 19021 11364 19079
rect 11376 19021 11388 19079
rect 11400 19021 11412 19079
rect 11424 19021 11436 19079
rect 11448 19021 11460 19079
rect 11472 19021 11484 19079
rect 11496 19021 11508 19079
rect 11520 19021 11532 19079
rect 10752 18805 10764 18839
rect 10776 18781 10788 18839
rect 10800 18709 10812 18839
rect 6912 18613 6924 18647
rect 10824 18541 10836 18839
rect 10848 18541 10860 18839
rect 10872 18541 10884 18839
rect 10896 18613 10908 18839
rect 10920 18613 10932 18839
rect 10944 18613 10956 18839
rect 10968 18613 10980 18839
rect 10992 18613 11004 18839
rect 11016 18613 11028 18839
rect 11040 18613 11052 18839
rect 11064 18613 11076 18839
rect 11088 18613 11100 18839
rect 11112 18613 11124 18839
rect 11136 18613 11148 18839
rect 11160 18613 11172 18839
rect 11184 18613 11196 18839
rect 11208 18613 11220 18839
rect 11232 18613 11244 18839
rect 11256 18613 11268 18839
rect 11280 18613 11292 18839
rect 11304 18613 11316 18839
rect 11328 18613 11340 18839
rect 11352 18613 11364 18839
rect 11376 18613 11388 18839
rect 11400 18613 11412 18839
rect 11424 18613 11436 18839
rect 11448 18781 11460 18839
rect 11448 18613 11460 18743
rect 11472 18613 11484 18839
rect 11496 18613 11508 18839
rect 11520 18613 11532 18839
rect 12048 18709 12060 18884
rect 11544 18613 11556 18695
rect 11568 18613 11580 18647
rect 12072 18613 12084 18695
rect 12163 18637 12175 18884
rect 12187 18661 12199 18884
rect 12211 18709 12223 18884
rect 12235 18757 12247 18884
rect 13507 18852 13519 18884
rect 13699 18852 13711 18884
rect 14491 18852 14503 18884
rect 15043 18852 15055 18884
rect 15259 18852 15271 18884
rect 16003 18852 16015 18884
rect 16171 18852 16183 18884
rect 16555 18852 16567 18884
rect 16747 18852 16759 18884
rect 16963 18852 16975 18884
rect 17707 18852 17719 18884
rect 17875 18852 17887 18884
rect 27283 18852 27295 18884
rect 27475 18852 27487 18884
rect 27715 18852 27727 18884
rect 35419 18852 35431 18884
rect 36163 18852 36175 18884
rect 13507 18840 13524 18852
rect 13699 18840 13716 18852
rect 14491 18840 14508 18852
rect 15043 18840 15060 18852
rect 15259 18840 15276 18852
rect 16003 18840 16020 18852
rect 16171 18840 16188 18852
rect 16555 18840 16572 18852
rect 16747 18840 16764 18852
rect 16963 18840 16980 18852
rect 17707 18840 17724 18852
rect 17875 18840 17892 18852
rect 27283 18840 27300 18852
rect 27475 18840 27492 18852
rect 27715 18840 27732 18852
rect 35419 18840 35436 18852
rect 36163 18840 36180 18852
rect 12936 18661 12948 18743
rect 13512 18661 13524 18840
rect 13704 18661 13716 18840
rect 14496 18661 14508 18840
rect 14520 18661 14532 18695
rect 15048 18637 15060 18840
rect 15264 18637 15276 18840
rect 16008 18637 16020 18840
rect 16176 18637 16188 18840
rect 16560 18637 16572 18840
rect 16752 18637 16764 18840
rect 16968 18637 16980 18840
rect 17712 18613 17724 18840
rect 17880 18613 17892 18840
rect 27288 18613 27300 18840
rect 27480 18637 27492 18840
rect 27720 18709 27732 18840
rect 35424 18709 35436 18840
rect 36168 18757 36180 18840
rect 36504 18757 36516 18884
rect 27744 18661 27756 18695
rect 36648 18661 36660 18839
rect 36672 18661 36684 18839
rect 36696 18661 36708 18839
rect 36720 18661 36732 18839
rect 36744 18661 36756 18839
rect 36768 18661 36780 18839
rect 36792 18709 36804 18743
rect 36816 18685 36828 18863
rect 36840 18757 36852 18815
rect 36840 18685 36852 18719
rect 36864 18685 36876 18815
rect 36888 18685 36900 18767
rect 36912 18685 36924 18767
rect 36936 18685 36948 18719
rect 6912 18205 6924 18239
rect 9408 18205 9420 18239
rect 6912 17965 6924 18071
rect 9240 17965 9252 18023
rect 9288 17965 9300 18071
rect 9312 17965 9324 18095
rect 9336 17965 9348 18119
rect 9360 17965 9372 18143
rect 9384 17965 9396 18167
rect 9408 17965 9420 18167
rect 9432 17965 9444 18191
rect 9456 17965 9468 18239
rect 9480 17965 9492 18263
rect 9504 17965 9516 18287
rect 9528 17965 9540 18311
rect 9552 17965 9564 17999
rect 9576 17965 9588 18335
rect 9600 17965 9612 18359
rect 9624 17965 9636 18383
rect 9648 17965 9660 17999
rect 9672 17965 9684 18407
rect 9696 17965 9708 18431
rect 9720 17965 9732 18455
rect 9744 17965 9756 18479
rect 9768 17965 9780 18503
rect 10032 18037 10044 18527
rect 16992 18421 17004 18455
rect 11112 18301 11124 18335
rect 11136 18301 11148 18335
rect 11160 18301 11172 18335
rect 11184 18253 11196 18335
rect 10056 17989 10068 18215
rect 11208 18205 11220 18335
rect 11232 18205 11244 18335
rect 11256 18205 11268 18335
rect 11280 18157 11292 18335
rect 11304 18157 11316 18335
rect 11328 18133 11340 18335
rect 11352 18133 11364 18335
rect 11376 18133 11388 18335
rect 11400 18133 11412 18335
rect 11424 18061 11436 18335
rect 10104 18013 10116 18047
rect 11448 18013 11460 18335
rect 11472 18013 11484 18335
rect 11496 18133 11508 18335
rect 10056 17939 10068 17951
rect 10174 17939 10186 17999
rect 10198 17939 10210 17951
rect 10222 17939 10234 17951
rect 10246 17939 10258 17999
rect 11496 17989 11508 18095
rect 11520 17989 11532 18335
rect 11544 18253 11556 18335
rect 11568 18037 11580 18335
rect 11592 18109 11604 18335
rect 11616 18253 11628 18287
rect 11640 18181 11652 18239
rect 11664 18157 11676 18191
rect 11616 18109 11628 18143
rect 11640 18085 11652 18119
rect 11592 18037 11604 18071
rect 12936 17964 12948 18239
rect 13512 18157 13524 18239
rect 13704 18205 13716 18239
rect 14496 17964 14508 18239
rect 12936 17952 12958 17964
rect 12946 17939 12958 17952
rect 14494 17952 14508 17964
rect 14520 17964 14532 18287
rect 14544 18253 14556 18287
rect 16968 17964 16980 18407
rect 18600 18253 18612 18455
rect 18576 17964 18588 18239
rect 20688 17964 20700 18455
rect 14520 17952 14542 17964
rect 16968 17952 16990 17964
rect 18576 17952 18598 17964
rect 14494 17939 14506 17952
rect 14530 17939 14542 17952
rect 16978 17939 16990 17952
rect 18586 17939 18598 17952
rect 20686 17952 20700 17964
rect 22080 17964 22092 18407
rect 23784 17964 23796 18407
rect 22080 17952 22102 17964
rect 20686 17939 20698 17952
rect 22090 17939 22102 17952
rect 23782 17952 23796 17964
rect 25320 17964 25332 18383
rect 25320 17952 25342 17964
rect 23782 17939 23794 17952
rect 25330 17939 25342 17952
rect 26866 17939 26878 18359
rect 26890 17939 26902 18335
rect 29938 17939 29950 18311
rect 30010 18253 30022 18287
rect 29962 17939 29974 18239
rect 31488 17964 31500 18239
rect 33024 17964 33036 18239
rect 36672 18229 36684 18263
rect 36696 18229 36708 18263
rect 34560 17964 34572 18191
rect 36648 18157 36660 18191
rect 36096 17964 36108 18143
rect 31488 17952 31510 17964
rect 33024 17952 33046 17964
rect 34560 17952 34582 17964
rect 36096 17952 36118 17964
rect 31498 17939 31510 17952
rect 33034 17939 33046 17952
rect 34570 17939 34582 17952
rect 36106 17939 36118 17952
rect 37848 17939 37860 18503
rect 38184 17965 38196 18479
rect 38208 17965 38220 18455
rect 38232 17965 38244 18431
rect 38256 17965 38268 18407
rect 38280 17965 38292 18383
rect 38304 17965 38316 18359
rect 38328 17965 38340 18335
rect 38352 17965 38364 18311
rect 38400 17989 38412 18287
rect 38424 17989 38436 18263
rect 38520 18133 38532 18239
rect 38496 18037 38508 18119
rect 38520 18037 38532 18071
rect 38544 18037 38556 18215
rect 38568 18037 38580 18191
rect 38592 18037 38604 18167
rect 38640 18061 38652 18143
rect 38616 17965 38628 17999
rect 38664 17965 38676 18095
rect 40752 17965 40764 18047
rect 40800 17965 40812 18023
rect 40824 17965 40836 17999
rect 9240 17701 9252 17735
rect 9288 17701 9300 17878
rect 9312 17701 9324 17878
rect 9336 17701 9348 17878
rect 9360 17701 9372 17878
rect 9384 17760 9396 17878
rect 9408 17701 9420 17878
rect 9432 17701 9444 17878
rect 9456 17785 9468 17878
rect 9480 17701 9492 17878
rect 9504 17701 9516 17878
rect 9528 17701 9540 17878
rect 9552 17701 9564 17830
rect 9576 17701 9588 17806
rect 9600 17701 9612 17806
rect 9624 17701 9636 17806
rect 9648 17701 9660 17806
rect 9672 17701 9684 17806
rect 9696 17701 9708 17806
rect 9720 17701 9732 17806
rect 9744 17701 9756 17806
rect 9768 17701 9780 17806
rect 9805 17772 9835 17784
rect 9805 17748 9835 17760
rect 9792 17725 9835 17736
rect 9805 17724 9835 17725
rect 38146 17724 38159 17736
rect 38146 17700 38159 17712
rect 38146 17676 38159 17688
rect 38146 17652 38159 17664
rect 38146 17628 38159 17640
rect 38146 17604 38159 17616
rect 38146 17580 38159 17592
rect 38184 17569 38196 17747
rect 38208 17569 38220 17747
rect 38232 17569 38244 17747
rect 38256 17569 38268 17747
rect 38280 17569 38292 17747
rect 38304 17665 38316 17747
rect 38328 17569 38340 17747
rect 38352 17689 38364 17747
rect 38376 17569 38388 17747
rect 38400 17617 38412 17747
rect 38424 17689 38436 17747
rect 38448 17689 38460 17747
rect 38472 17689 38484 17747
rect 38496 17689 38508 17747
rect 38520 17689 38532 17747
rect 38544 17713 38556 17747
rect 38448 17569 38460 17603
rect 38472 17569 38484 17603
rect 38496 17569 38508 17603
rect 38520 17569 38532 17603
rect 38616 17569 38628 17603
rect 40776 16957 40788 16991
rect 5880 16909 5892 16943
rect 6840 16909 6852 16943
rect 9240 16909 9252 16943
rect 9288 16909 9300 16943
rect 9312 16909 9324 16943
rect 9336 16909 9348 16943
rect 9360 16909 9372 16943
rect 9408 16909 9420 16943
rect 9432 16909 9444 16943
rect 9480 16909 9492 16943
rect 9504 16909 9516 16943
rect 9528 16909 9540 16943
rect 9552 16909 9564 16943
rect 9576 16909 9588 16943
rect 9600 16909 9612 16943
rect 9624 16909 9636 16943
rect 40800 16909 40812 16943
rect 40824 16909 40836 16991
rect 40848 16909 40860 16991
rect 38256 16765 38268 16799
rect 38280 16765 38292 16799
rect 38328 16765 38340 16799
rect 38376 16765 38388 16799
rect 38448 16765 38460 16799
rect 38472 16765 38484 16799
rect 38496 16765 38508 16799
rect 38520 16765 38532 16799
rect 38616 16765 38628 16799
rect 40800 16765 40812 16799
rect 40824 16765 40836 16799
rect 40848 16765 40860 16799
rect 6840 13204 6852 13247
rect 9240 13209 9252 13247
rect 9288 13209 9300 13247
rect 9312 13209 9324 13247
rect 9336 13209 9348 13247
rect 9360 13209 9372 13247
rect 9408 13154 9420 13247
rect 9432 13154 9444 13247
rect 9480 13154 9492 13247
rect 9504 13154 9516 13247
rect 9528 13154 9540 13247
rect 9552 13154 9564 13247
rect 9576 13154 9588 13247
rect 9600 13154 9612 13319
rect 9624 13154 9636 13319
rect 9648 13154 9660 13319
rect 9672 13154 9684 13343
rect 9696 13154 9708 13343
rect 9720 13154 9732 13343
rect 9744 13256 9756 13295
rect 9805 13243 9835 13255
rect 9805 13219 9835 13231
rect 9805 13195 9835 13207
rect 9744 13154 9756 13194
rect 9805 13171 9835 13183
rect 40800 12205 40812 12263
rect 40824 12181 40836 12287
rect 40848 12181 40860 12215
rect 40848 12037 40860 12071
rect 38146 11639 38159 11647
rect 38146 11635 38173 11639
rect 38184 11629 38196 11663
rect 38208 11629 38220 11663
rect 38146 11107 38159 11119
rect 38146 11083 38159 11095
rect 38184 11072 38196 11130
rect 38208 11072 38220 11130
rect 38280 11072 38292 11130
rect 38328 11072 38340 11130
rect 38376 11072 38388 11130
rect 38448 11072 38460 11130
rect 38472 11072 38484 11130
rect 38496 11096 38508 11130
rect 38146 9266 38159 9278
rect 38146 9242 38159 9254
rect 9504 9157 9516 9239
rect 9528 9157 9540 9239
rect 9552 9205 9564 9239
rect 9576 9133 9588 9239
rect 9600 9061 9612 9239
rect 9624 9061 9636 9239
rect 9648 9061 9660 9239
rect 9672 9037 9684 9239
rect 9696 9037 9708 9239
rect 9720 9037 9732 9239
rect 6840 8941 6852 8975
rect 9240 8941 9252 8975
rect 9288 8941 9300 8975
rect 9312 8941 9324 8975
rect 9336 8941 9348 8975
rect 9408 8941 9420 8975
rect 9504 8941 9516 8975
rect 9600 8941 9612 8975
rect 9624 8941 9636 8975
rect 9744 8821 9756 9239
rect 9768 8821 9780 9239
rect 9805 9218 9835 9230
rect 38146 9218 38159 9230
rect 9805 9194 9835 9206
rect 38146 9194 38159 9206
rect 9805 9170 9835 9182
rect 38146 9170 38159 9182
rect 9805 9146 9835 9158
rect 38146 9146 38159 9158
rect 9792 8821 9804 9071
rect 9816 8821 9828 9047
rect 10174 9037 10186 9140
rect 10222 9109 10234 9140
rect 10246 9109 10258 9140
rect 38184 9133 38196 9287
rect 38208 9256 38220 9287
rect 38280 9160 38292 9287
rect 38328 9157 38340 9287
rect 9840 8821 9852 9023
rect 9864 8821 9876 8999
rect 9888 8821 9900 8975
rect 9912 8821 9924 8903
rect 9936 8869 9948 8903
rect 6840 7453 6852 7487
rect 9240 7453 9252 7487
rect 9288 7453 9300 7487
rect 9312 7453 9324 7487
rect 9336 7453 9348 7487
rect 9408 7453 9420 7487
rect 9504 7453 9516 7487
rect 38328 7453 38340 7487
rect 9336 6565 9348 6719
rect 9408 6613 9420 6719
rect 6840 6517 6852 6551
rect 9504 6517 9516 6719
rect 9744 6541 9756 6719
rect 9768 6685 9780 6719
rect 9792 6637 9804 6719
rect 9816 6685 9828 6719
rect 9768 6541 9780 6623
rect 10944 6517 10956 6791
rect 11088 6589 11100 6767
rect 11064 6493 11076 6575
rect 11112 6493 11124 6647
rect 15048 6493 15060 6743
rect 15216 6685 15228 6719
rect 15192 6493 15204 6671
rect 15240 6493 15252 6647
rect 19200 6517 19212 6695
rect 19320 6493 19332 6671
rect 19368 6493 19380 6647
rect 27456 6517 27468 6647
rect 27576 6493 27588 6599
rect 31560 6493 31572 6599
rect 31728 6541 31740 6575
rect 31704 6493 31716 6527
rect 35688 6493 35700 6551
rect 35832 6493 35844 6527
<< metal4 >>
rect 6080 46264 7640 47824
rect 10208 46264 11768 47824
rect 14336 46264 15896 47824
rect 18464 46264 20024 47824
rect 22592 46264 24152 47824
rect 26720 46264 28280 47824
rect 30848 46264 32408 47824
rect 34976 46264 36536 47824
rect 39104 46264 40664 47824
rect -544 39726 1016 41286
rect 45728 39726 47288 41286
rect -544 34996 1016 36556
rect 45728 34996 47288 36556
rect -544 30266 1016 31826
rect 45728 30266 47288 31826
rect -544 25536 1016 27096
rect 45728 25536 47288 27096
rect -544 20806 1016 22366
rect 45728 20806 47288 22366
rect -544 16076 1016 17636
rect 45728 16076 47288 17636
rect -544 11346 1016 12906
rect 45728 11346 47288 12906
rect -544 6616 1016 8176
rect 45728 6616 47288 8176
rect 6080 78 7640 1638
rect 10208 78 11768 1638
rect 14336 78 15896 1638
rect 18464 78 20024 1638
rect 22592 78 24152 1638
rect 26720 78 28280 1638
rect 30848 78 32408 1638
rect 34976 78 36536 1638
rect 39104 78 40664 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 -622 -1 0 47902
box 0 0 6450 6450
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform 0 -1 5914 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform 0 -1 6000 1 0 41452
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 7720 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform 0 -1 7806 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform 0 -1 7892 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform 0 -1 7978 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform 0 -1 8064 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform 0 -1 8150 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform 0 -1 8236 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform 0 -1 8322 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform 0 -1 8408 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform 0 -1 8494 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform 0 -1 8580 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform 0 -1 8666 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform 0 -1 8752 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform 0 -1 8838 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform 0 -1 8924 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform 0 -1 9010 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform 0 -1 9096 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform 0 -1 9182 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform 0 -1 9268 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform 0 -1 9354 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform 0 -1 9440 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform 0 -1 9526 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform 0 -1 9612 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform 0 -1 9698 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform 0 -1 9784 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform 0 -1 9870 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform 0 -1 9956 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform 0 -1 10042 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform 0 -1 10128 1 0 41452
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 11848 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform 0 -1 11934 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform 0 -1 12020 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform 0 -1 12106 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform 0 -1 12192 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform 0 -1 12278 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform 0 -1 12364 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform 0 -1 12450 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform 0 -1 12536 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform 0 -1 12622 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform 0 -1 12708 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform 0 -1 12794 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform 0 -1 12880 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform 0 -1 12966 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform 0 -1 13052 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform 0 -1 13138 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform 0 -1 13224 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform 0 -1 13310 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform 0 -1 13396 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform 0 -1 13482 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform 0 -1 13568 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform 0 -1 13654 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform 0 -1 13740 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform 0 -1 13826 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform 0 -1 13912 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform 0 -1 13998 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform 0 -1 14084 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform 0 -1 14170 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform 0 -1 14256 1 0 41452
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 15976 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform 0 -1 16062 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform 0 -1 16148 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform 0 -1 16234 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform 0 -1 16320 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform 0 -1 16406 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform 0 -1 16492 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform 0 -1 16578 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform 0 -1 16664 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform 0 -1 16750 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform 0 -1 16836 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform 0 -1 16922 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform 0 -1 17008 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform 0 -1 17094 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform 0 -1 17180 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform 0 -1 17266 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform 0 -1 17352 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform 0 -1 17438 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform 0 -1 17524 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform 0 -1 17610 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform 0 -1 17696 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform 0 -1 17782 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform 0 -1 17868 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform 0 -1 17954 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform 0 -1 18040 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform 0 -1 18126 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform 0 -1 18212 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform 0 -1 18298 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform 0 -1 18384 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 20104 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform 0 -1 20190 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform 0 -1 20276 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform 0 -1 20362 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform 0 -1 20448 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform 0 -1 20534 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform 0 -1 20620 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform 0 -1 20706 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform 0 -1 20792 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform 0 -1 20878 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform 0 -1 20964 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform 0 -1 21050 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform 0 -1 21136 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform 0 -1 21222 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform 0 -1 21308 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform 0 -1 21394 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform 0 -1 21480 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform 0 -1 21566 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform 0 -1 21652 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform 0 -1 21738 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform 0 -1 21824 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform 0 -1 21910 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform 0 -1 21996 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform 0 -1 22082 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform 0 -1 22168 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform 0 -1 22254 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform 0 -1 22340 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform 0 -1 22426 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform 0 -1 22512 1 0 41452
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 24232 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform 0 -1 24318 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform 0 -1 24404 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform 0 -1 24490 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform 0 -1 24576 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform 0 -1 24662 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform 0 -1 24748 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform 0 -1 24834 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform 0 -1 24920 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform 0 -1 25006 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform 0 -1 25092 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform 0 -1 25178 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform 0 -1 25264 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform 0 -1 25350 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform 0 -1 25436 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform 0 -1 25522 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform 0 -1 25608 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform 0 -1 25694 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform 0 -1 25780 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform 0 -1 25866 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform 0 -1 25952 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform 0 -1 26038 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform 0 -1 26124 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform 0 -1 26210 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform 0 -1 26296 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform 0 -1 26382 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 26468 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 26554 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 26640 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 28360 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 28446 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 28532 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 28618 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 28704 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 28790 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 28876 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 28962 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 29048 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 29134 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 29220 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 29306 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 29392 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 29478 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 29564 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 29650 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 29736 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 29822 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 0 -1 29908 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 0 -1 29994 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 0 -1 30080 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 0 -1 30166 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 0 -1 30252 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 0 -1 30338 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 0 -1 30424 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 0 -1 30510 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 0 -1 30596 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 0 -1 30682 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 0 -1 30768 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 32488 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 0 -1 32574 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 0 -1 32660 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 0 -1 32746 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 0 -1 32832 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 32918 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 33004 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 33090 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 33176 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 33262 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 33348 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 33434 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 33520 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 33606 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 33692 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 33778 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 33864 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 33950 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 34036 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 34122 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 34208 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 34294 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 34380 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 34466 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 34552 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 34638 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 34724 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 34810 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 34896 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 36616 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 36702 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 36788 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 36874 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 36960 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 37046 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 37132 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 37218 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 37304 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 37390 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 37476 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 37562 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 37648 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 37734 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 37820 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 37906 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 37992 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 38078 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 38164 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 38250 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 38336 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 38422 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 38508 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 38594 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 38680 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 38766 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 38852 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 38938 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 39024 1 0 41452
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 40744 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 40830 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 40916 1 0 41452
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 47366 0 -1 47902
box 0 0 6450 6450
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 5828 0 -1 41452
box 0 0 6450 86
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 5828 0 -1 41366
box 0 0 6450 1720
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 5828 0 -1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 5828 0 -1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 5828 0 -1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 1 0 40916 0 1 41366
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 40916 0 1 39646
box 0 0 6450 1720
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 1 0 40916 0 1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 1 0 40916 0 1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 5828 0 -1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 5828 0 -1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 5828 0 -1 39216
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 5828 0 -1 39130
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 5828 0 -1 39044
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 5828 0 -1 38958
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 5828 0 -1 38872
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 5828 0 -1 38786
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 5828 0 -1 38700
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 5828 0 -1 38614
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 5828 0 -1 38528
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform -1 0 5828 0 -1 38442
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform -1 0 5828 0 -1 38356
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform -1 0 5828 0 -1 38270
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform -1 0 5828 0 -1 38184
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform -1 0 5828 0 -1 38098
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform -1 0 5828 0 -1 38012
box 0 0 6450 86
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform -1 0 5828 0 -1 37926
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform -1 0 5828 0 -1 37840
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform -1 0 5828 0 -1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform -1 0 5828 0 -1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform -1 0 5828 0 -1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform -1 0 5828 0 -1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform -1 0 5828 0 -1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform -1 0 5828 0 -1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform -1 0 5828 0 -1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform -1 0 5828 0 -1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform -1 0 5828 0 -1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform -1 0 5828 0 -1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform -1 0 5828 0 -1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform -1 0 5828 0 -1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform -1 0 5828 0 -1 36722
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 5828 0 -1 36636
box 0 0 6450 1720
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform -1 0 5828 0 -1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform -1 0 5828 0 -1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform -1 0 5828 0 -1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform -1 0 5828 0 -1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform -1 0 5828 0 -1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform -1 0 5828 0 -1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform -1 0 5828 0 -1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform -1 0 5828 0 -1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform -1 0 5828 0 -1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform -1 0 5828 0 -1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform -1 0 5828 0 -1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform -1 0 5828 0 -1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform -1 0 5828 0 -1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform -1 0 5828 0 -1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform -1 0 5828 0 -1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform -1 0 5828 0 -1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform -1 0 5828 0 -1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform -1 0 5828 0 -1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform -1 0 5828 0 -1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform -1 0 5828 0 -1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform -1 0 5828 0 -1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform -1 0 5828 0 -1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform -1 0 5828 0 -1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform -1 0 5828 0 -1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform -1 0 5828 0 -1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform -1 0 5828 0 -1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform -1 0 5828 0 -1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform -1 0 5828 0 -1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform -1 0 5828 0 -1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform -1 0 5828 0 -1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform -1 0 5828 0 -1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform -1 0 5828 0 -1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform -1 0 5828 0 -1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform -1 0 5828 0 -1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform -1 0 5828 0 -1 31992
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 5828 0 -1 31906
box 0 0 6450 1720
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform -1 0 5828 0 -1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform -1 0 5828 0 -1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform -1 0 5828 0 -1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform -1 0 5828 0 -1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform -1 0 5828 0 -1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform -1 0 5828 0 -1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform -1 0 5828 0 -1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform -1 0 5828 0 -1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform -1 0 5828 0 -1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform -1 0 5828 0 -1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform -1 0 5828 0 -1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform -1 0 5828 0 -1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform -1 0 5828 0 -1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform -1 0 5828 0 -1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_788
timestamp 1300117811
transform -1 0 5828 0 -1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_789
timestamp 1300117811
transform -1 0 5828 0 -1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_790
timestamp 1300117811
transform -1 0 5828 0 -1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_791
timestamp 1300117811
transform -1 0 5828 0 -1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_792
timestamp 1300117811
transform -1 0 5828 0 -1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_793
timestamp 1300117811
transform -1 0 5828 0 -1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_794
timestamp 1300117811
transform -1 0 5828 0 -1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_795
timestamp 1300117811
transform -1 0 5828 0 -1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_796
timestamp 1300117811
transform -1 0 5828 0 -1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_797
timestamp 1300117811
transform -1 0 5828 0 -1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_798
timestamp 1300117811
transform -1 0 5828 0 -1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_799
timestamp 1300117811
transform -1 0 5828 0 -1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_800
timestamp 1300117811
transform -1 0 5828 0 -1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_801
timestamp 1300117811
transform -1 0 5828 0 -1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_802
timestamp 1300117811
transform -1 0 5828 0 -1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_803
timestamp 1300117811
transform -1 0 5828 0 -1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_804
timestamp 1300117811
transform -1 0 5828 0 -1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_805
timestamp 1300117811
transform -1 0 5828 0 -1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_806
timestamp 1300117811
transform -1 0 5828 0 -1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_807
timestamp 1300117811
transform -1 0 5828 0 -1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_808
timestamp 1300117811
transform -1 0 5828 0 -1 27262
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 5828 0 -1 27176
box 0 0 6450 1720
use fillpp_mt fillpp_mt_809
timestamp 1300117811
transform -1 0 5828 0 -1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_810
timestamp 1300117811
transform -1 0 5828 0 -1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_811
timestamp 1300117811
transform -1 0 5828 0 -1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_812
timestamp 1300117811
transform -1 0 5828 0 -1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_813
timestamp 1300117811
transform -1 0 5828 0 -1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_814
timestamp 1300117811
transform -1 0 5828 0 -1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_815
timestamp 1300117811
transform -1 0 5828 0 -1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_816
timestamp 1300117811
transform -1 0 5828 0 -1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_817
timestamp 1300117811
transform -1 0 5828 0 -1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_818
timestamp 1300117811
transform -1 0 5828 0 -1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_819
timestamp 1300117811
transform -1 0 5828 0 -1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_820
timestamp 1300117811
transform -1 0 5828 0 -1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_821
timestamp 1300117811
transform -1 0 5828 0 -1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_822
timestamp 1300117811
transform -1 0 5828 0 -1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_823
timestamp 1300117811
transform -1 0 5828 0 -1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_824
timestamp 1300117811
transform -1 0 5828 0 -1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_825
timestamp 1300117811
transform -1 0 5828 0 -1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_826
timestamp 1300117811
transform -1 0 5828 0 -1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_827
timestamp 1300117811
transform -1 0 5828 0 -1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_828
timestamp 1300117811
transform -1 0 5828 0 -1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_829
timestamp 1300117811
transform -1 0 5828 0 -1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_830
timestamp 1300117811
transform -1 0 5828 0 -1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_831
timestamp 1300117811
transform -1 0 5828 0 -1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_832
timestamp 1300117811
transform -1 0 5828 0 -1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_833
timestamp 1300117811
transform -1 0 5828 0 -1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_834
timestamp 1300117811
transform -1 0 5828 0 -1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_835
timestamp 1300117811
transform -1 0 5828 0 -1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_836
timestamp 1300117811
transform -1 0 5828 0 -1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_837
timestamp 1300117811
transform -1 0 5828 0 -1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_838
timestamp 1300117811
transform -1 0 5828 0 -1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_839
timestamp 1300117811
transform -1 0 5828 0 -1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_840
timestamp 1300117811
transform -1 0 5828 0 -1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_841
timestamp 1300117811
transform -1 0 5828 0 -1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_842
timestamp 1300117811
transform -1 0 5828 0 -1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_843
timestamp 1300117811
transform -1 0 5828 0 -1 22532
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 5828 0 -1 22446
box 0 0 6450 1720
use fillpp_mt fillpp_mt_844
timestamp 1300117811
transform -1 0 5828 0 -1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_845
timestamp 1300117811
transform -1 0 5828 0 -1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_846
timestamp 1300117811
transform -1 0 5828 0 -1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_847
timestamp 1300117811
transform -1 0 5828 0 -1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_848
timestamp 1300117811
transform -1 0 5828 0 -1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_849
timestamp 1300117811
transform -1 0 5828 0 -1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_850
timestamp 1300117811
transform -1 0 5828 0 -1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_851
timestamp 1300117811
transform -1 0 5828 0 -1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_852
timestamp 1300117811
transform -1 0 5828 0 -1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_853
timestamp 1300117811
transform -1 0 5828 0 -1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_854
timestamp 1300117811
transform -1 0 5828 0 -1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_855
timestamp 1300117811
transform -1 0 5828 0 -1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_856
timestamp 1300117811
transform -1 0 5828 0 -1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_857
timestamp 1300117811
transform -1 0 5828 0 -1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_858
timestamp 1300117811
transform -1 0 5828 0 -1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_859
timestamp 1300117811
transform -1 0 5828 0 -1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_860
timestamp 1300117811
transform -1 0 5828 0 -1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_861
timestamp 1300117811
transform -1 0 5828 0 -1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_862
timestamp 1300117811
transform -1 0 5828 0 -1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_863
timestamp 1300117811
transform -1 0 5828 0 -1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_864
timestamp 1300117811
transform -1 0 5828 0 -1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_865
timestamp 1300117811
transform -1 0 5828 0 -1 18920
box 0 0 6450 86
use datapath datapath_0
timestamp 1395340701
transform 1 0 11158 0 1 18841
box 414 43 25445 20615
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 1 0 40916 0 1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 1 0 40916 0 1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 1 0 40916 0 1 39216
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 1 0 40916 0 1 39130
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 1 0 40916 0 1 39044
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 1 0 40916 0 1 38958
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 1 0 40916 0 1 38872
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 1 0 40916 0 1 38786
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 1 0 40916 0 1 38700
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 1 0 40916 0 1 38614
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 1 0 40916 0 1 38528
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 1 0 40916 0 1 38442
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 1 0 40916 0 1 38356
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 1 0 40916 0 1 38270
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 1 0 40916 0 1 38184
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 1 0 40916 0 1 38098
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 1 0 40916 0 1 38012
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 1 0 40916 0 1 37926
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 1 0 40916 0 1 37840
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 1 0 40916 0 1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 1 0 40916 0 1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 1 0 40916 0 1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 1 0 40916 0 1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 1 0 40916 0 1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 1 0 40916 0 1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 1 0 40916 0 1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 1 0 40916 0 1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 1 0 40916 0 1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 1 0 40916 0 1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 1 0 40916 0 1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 1 0 40916 0 1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 1 0 40916 0 1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 1 0 40916 0 1 36636
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 40916 0 1 34916
box 0 0 6450 1720
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 1 0 40916 0 1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 1 0 40916 0 1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 1 0 40916 0 1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 1 0 40916 0 1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 1 0 40916 0 1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 1 0 40916 0 1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 1 0 40916 0 1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 1 0 40916 0 1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 1 0 40916 0 1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 1 0 40916 0 1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 1 0 40916 0 1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 1 0 40916 0 1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 1 0 40916 0 1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 1 0 40916 0 1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 1 0 40916 0 1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 1 0 40916 0 1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 1 0 40916 0 1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 1 0 40916 0 1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 1 0 40916 0 1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 1 0 40916 0 1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 1 0 40916 0 1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 1 0 40916 0 1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 1 0 40916 0 1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 1 0 40916 0 1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 1 0 40916 0 1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 1 0 40916 0 1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 1 0 40916 0 1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 1 0 40916 0 1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 1 0 40916 0 1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 1 0 40916 0 1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 1 0 40916 0 1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 1 0 40916 0 1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 1 0 40916 0 1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 1 0 40916 0 1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 1 0 40916 0 1 31906
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 40916 0 1 30186
box 0 0 6450 1720
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 1 0 40916 0 1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 1 0 40916 0 1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 1 0 40916 0 1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 1 0 40916 0 1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 1 0 40916 0 1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 1 0 40916 0 1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 1 0 40916 0 1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 1 0 40916 0 1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 1 0 40916 0 1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 1 0 40916 0 1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 40916 0 1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 40916 0 1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 40916 0 1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 40916 0 1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 40916 0 1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 40916 0 1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 40916 0 1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 40916 0 1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 40916 0 1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 40916 0 1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 40916 0 1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 40916 0 1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 40916 0 1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 40916 0 1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 40916 0 1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 40916 0 1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 40916 0 1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 40916 0 1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 40916 0 1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 40916 0 1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 40916 0 1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 40916 0 1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 40916 0 1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 40916 0 1 27262
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 40916 0 1 27176
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 40916 0 1 25456
box 0 0 6450 1720
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 40916 0 1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 40916 0 1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 40916 0 1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 40916 0 1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 40916 0 1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 40916 0 1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 40916 0 1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 40916 0 1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 40916 0 1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 40916 0 1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 40916 0 1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 40916 0 1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 40916 0 1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 40916 0 1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 40916 0 1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 40916 0 1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 40916 0 1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 40916 0 1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 40916 0 1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 40916 0 1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 40916 0 1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 40916 0 1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 40916 0 1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 40916 0 1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 40916 0 1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 40916 0 1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 40916 0 1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 40916 0 1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 40916 0 1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 40916 0 1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 40916 0 1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 40916 0 1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 40916 0 1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 40916 0 1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 40916 0 1 22446
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 40916 0 1 20726
box 0 0 6450 1720
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 40916 0 1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 40916 0 1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 40916 0 1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 40916 0 1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 40916 0 1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 40916 0 1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 40916 0 1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 40916 0 1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 40916 0 1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 40916 0 1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 40916 0 1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 40916 0 1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 40916 0 1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 40916 0 1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 40916 0 1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 40916 0 1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 40916 0 1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 40916 0 1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 40916 0 1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 40916 0 1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 40916 0 1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_866
timestamp 1300117811
transform -1 0 5828 0 -1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_867
timestamp 1300117811
transform -1 0 5828 0 -1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_868
timestamp 1300117811
transform -1 0 5828 0 -1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_869
timestamp 1300117811
transform -1 0 5828 0 -1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_870
timestamp 1300117811
transform -1 0 5828 0 -1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_871
timestamp 1300117811
transform -1 0 5828 0 -1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_872
timestamp 1300117811
transform -1 0 5828 0 -1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_873
timestamp 1300117811
transform -1 0 5828 0 -1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_874
timestamp 1300117811
transform -1 0 5828 0 -1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_875
timestamp 1300117811
transform -1 0 5828 0 -1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_876
timestamp 1300117811
transform -1 0 5828 0 -1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 40916 0 1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 40916 0 1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 40916 0 1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 40916 0 1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 40916 0 1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 40916 0 1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 40916 0 1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 40916 0 1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 40916 0 1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 40916 0 1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 40916 0 1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_877
timestamp 1300117811
transform -1 0 5828 0 -1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_878
timestamp 1300117811
transform -1 0 5828 0 -1 17802
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 5828 0 -1 17716
box 0 0 6450 1720
use fillpp_mt fillpp_mt_879
timestamp 1300117811
transform -1 0 5828 0 -1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_880
timestamp 1300117811
transform -1 0 5828 0 -1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_881
timestamp 1300117811
transform -1 0 5828 0 -1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_882
timestamp 1300117811
transform -1 0 5828 0 -1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_883
timestamp 1300117811
transform -1 0 5828 0 -1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_884
timestamp 1300117811
transform -1 0 5828 0 -1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_885
timestamp 1300117811
transform -1 0 5828 0 -1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_886
timestamp 1300117811
transform -1 0 5828 0 -1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_887
timestamp 1300117811
transform -1 0 5828 0 -1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_888
timestamp 1300117811
transform -1 0 5828 0 -1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_889
timestamp 1300117811
transform -1 0 5828 0 -1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_890
timestamp 1300117811
transform -1 0 5828 0 -1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_891
timestamp 1300117811
transform -1 0 5828 0 -1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_892
timestamp 1300117811
transform -1 0 5828 0 -1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_893
timestamp 1300117811
transform -1 0 5828 0 -1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_894
timestamp 1300117811
transform -1 0 5828 0 -1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_895
timestamp 1300117811
transform -1 0 5828 0 -1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_896
timestamp 1300117811
transform -1 0 5828 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_897
timestamp 1300117811
transform -1 0 5828 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_898
timestamp 1300117811
transform -1 0 5828 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_899
timestamp 1300117811
transform -1 0 5828 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_900
timestamp 1300117811
transform -1 0 5828 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_901
timestamp 1300117811
transform -1 0 5828 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_902
timestamp 1300117811
transform -1 0 5828 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_903
timestamp 1300117811
transform -1 0 5828 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_904
timestamp 1300117811
transform -1 0 5828 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_905
timestamp 1300117811
transform -1 0 5828 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_906
timestamp 1300117811
transform -1 0 5828 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_907
timestamp 1300117811
transform -1 0 5828 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_908
timestamp 1300117811
transform -1 0 5828 0 -1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_909
timestamp 1300117811
transform -1 0 5828 0 -1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_910
timestamp 1300117811
transform -1 0 5828 0 -1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_911
timestamp 1300117811
transform -1 0 5828 0 -1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_912
timestamp 1300117811
transform -1 0 5828 0 -1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_913
timestamp 1300117811
transform -1 0 5828 0 -1 13072
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 5828 0 -1 12986
box 0 0 6450 1720
use fillpp_mt fillpp_mt_914
timestamp 1300117811
transform -1 0 5828 0 -1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_915
timestamp 1300117811
transform -1 0 5828 0 -1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_916
timestamp 1300117811
transform -1 0 5828 0 -1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_917
timestamp 1300117811
transform -1 0 5828 0 -1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_918
timestamp 1300117811
transform -1 0 5828 0 -1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_919
timestamp 1300117811
transform -1 0 5828 0 -1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_920
timestamp 1300117811
transform -1 0 5828 0 -1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_921
timestamp 1300117811
transform -1 0 5828 0 -1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_922
timestamp 1300117811
transform -1 0 5828 0 -1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_923
timestamp 1300117811
transform -1 0 5828 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_924
timestamp 1300117811
transform -1 0 5828 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_925
timestamp 1300117811
transform -1 0 5828 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_926
timestamp 1300117811
transform -1 0 5828 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_927
timestamp 1300117811
transform -1 0 5828 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_928
timestamp 1300117811
transform -1 0 5828 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_929
timestamp 1300117811
transform -1 0 5828 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_930
timestamp 1300117811
transform -1 0 5828 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_931
timestamp 1300117811
transform -1 0 5828 0 -1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_932
timestamp 1300117811
transform -1 0 5828 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_933
timestamp 1300117811
transform -1 0 5828 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_934
timestamp 1300117811
transform -1 0 5828 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_935
timestamp 1300117811
transform -1 0 5828 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_936
timestamp 1300117811
transform -1 0 5828 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_937
timestamp 1300117811
transform -1 0 5828 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_938
timestamp 1300117811
transform -1 0 5828 0 -1 9202
box 0 0 6450 86
use control control_0
timestamp 1395422108
transform 1 0 9835 0 1 9140
box 0 0 28311 8799
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 40916 0 1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 40916 0 1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 40916 0 1 17716
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 40916 0 1 15996
box 0 0 6450 1720
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 40916 0 1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 40916 0 1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 40916 0 1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 40916 0 1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 40916 0 1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 40916 0 1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 40916 0 1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 40916 0 1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 40916 0 1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 40916 0 1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 40916 0 1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 40916 0 1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 40916 0 1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 40916 0 1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 40916 0 1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 40916 0 1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 40916 0 1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 40916 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 40916 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 40916 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 40916 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 40916 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 40916 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 40916 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 40916 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 40916 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 40916 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 40916 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 40916 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 40916 0 1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 40916 0 1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 40916 0 1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 40916 0 1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 40916 0 1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 40916 0 1 12986
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 40916 0 1 11266
box 0 0 6450 1720
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 40916 0 1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 40916 0 1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 40916 0 1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 40916 0 1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 40916 0 1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 40916 0 1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 40916 0 1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 40916 0 1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 40916 0 1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 40916 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 40916 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 40916 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 40916 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 40916 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 40916 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 40916 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 40916 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 40916 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 40916 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 40916 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 40916 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 40916 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 40916 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 40916 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_939
timestamp 1300117811
transform -1 0 5828 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_940
timestamp 1300117811
transform -1 0 5828 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_941
timestamp 1300117811
transform -1 0 5828 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_942
timestamp 1300117811
transform -1 0 5828 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_943
timestamp 1300117811
transform -1 0 5828 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_944
timestamp 1300117811
transform -1 0 5828 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_945
timestamp 1300117811
transform -1 0 5828 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_946
timestamp 1300117811
transform -1 0 5828 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_947
timestamp 1300117811
transform -1 0 5828 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_948
timestamp 1300117811
transform -1 0 5828 0 -1 8342
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 5828 0 -1 8256
box 0 0 6450 1720
use fillpp_mt fillpp_mt_949
timestamp 1300117811
transform -1 0 5828 0 -1 6536
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 40916 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 40916 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 40916 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 40916 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 40916 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 40916 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 40916 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 40916 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 40916 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 40916 0 1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 40916 0 1 8256
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 40916 0 1 6536
box 0 0 6450 1720
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 40916 0 1 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 -622 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 5828 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 5914 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6000 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 7720 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 7806 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 7892 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 7978 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8064 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8150 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8236 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8322 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 8408 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 8494 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 8580 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 8666 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 8752 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 8838 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 8924 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9010 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9096 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9182 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9268 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9354 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 9440 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 9526 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 9612 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 9698 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 9784 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 9870 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 9956 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 10042 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10128 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 11848 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 11934 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 12020 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 12106 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 12192 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12278 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12364 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 12450 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 12536 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 12622 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 12708 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 12794 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 12880 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 12966 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 13052 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 13138 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 13224 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 13310 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 13396 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 13482 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 13568 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 13654 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 13740 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 13826 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 13912 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 13998 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 14084 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 14170 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 14256 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 15976 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 16062 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 16148 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 16234 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 16320 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 16406 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 16492 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 16578 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 16664 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 16750 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 16836 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 16922 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 17008 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 17094 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 17180 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 17266 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 17352 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 17438 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 17524 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 17610 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 17696 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 17782 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 17868 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 17954 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 18040 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 18126 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 18212 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 18298 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 18384 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 20104 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 20190 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 20276 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 20362 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 20448 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 20534 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 20620 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 20706 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 20792 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 20878 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 20964 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 21050 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 21136 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 21222 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 21308 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 21394 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 21480 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 21566 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 21652 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 21738 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 21824 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 21910 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 21996 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 22082 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 22168 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 22254 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 22340 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 22426 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 22512 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 24232 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 24318 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 24404 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 24490 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 24576 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 24662 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 24748 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 24834 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 24920 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 25006 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 25092 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 25178 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 25264 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 25350 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 25436 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 25522 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 25608 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 25694 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 25780 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 25866 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 25952 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 26038 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 26124 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 26210 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 26296 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 26382 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 26468 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 26554 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 26640 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 28360 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 28446 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 28532 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 28618 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 28704 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 28790 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 28876 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 28962 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 29048 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 29134 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 29220 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 29306 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 29392 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 29478 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 29564 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 29650 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 29736 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 29822 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 29908 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 29994 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 30080 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 30166 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 30252 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 30338 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 30424 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 30510 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 30596 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 30682 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 30768 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 0 1 32488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 0 1 32574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 0 1 32660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 0 1 32746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 0 1 32832 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 0 1 32918 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 0 1 33004 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 0 1 33090 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 0 1 33176 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 0 1 33262 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 0 1 33348 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 0 1 33434 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 0 1 33520 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 0 1 33606 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 0 1 33692 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 0 1 33778 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 0 1 33864 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 0 1 33950 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 0 1 34036 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 0 1 34122 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 0 1 34208 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 0 1 34294 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 0 1 34380 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 0 1 34466 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 0 1 34552 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 0 1 34638 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 0 1 34724 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 0 1 34810 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 34896 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 0 1 36616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 0 1 36702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 0 1 36788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 0 1 36874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 0 1 36960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 0 1 37046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 0 1 37132 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 0 1 37218 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 0 1 37304 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 0 1 37390 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 0 1 37476 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 0 1 37562 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 0 1 37648 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 0 1 37734 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 0 1 37820 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 0 1 37906 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 0 1 37992 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 0 1 38078 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 0 1 38164 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 0 1 38250 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 0 1 38336 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 0 1 38422 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 0 1 38508 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 0 1 38594 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 0 1 38680 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 0 1 38766 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 0 1 38852 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 0 1 38938 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 39024 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 0 1 40744 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 0 1 40830 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 47366 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 6080 78 7640 1638 0 nIRQ
rlabel metal4 10208 78 11768 1638 0 Data[0]
rlabel metal4 14336 78 15896 1638 0 Data[1]
rlabel metal4 18464 78 20024 1638 0 Data[2]
rlabel metal4 22592 78 24152 1638 0 vdde!
rlabel metal4 26720 78 28280 1638 0 Data[3]
rlabel metal4 30848 78 32408 1638 0 Data[4]
rlabel metal4 34976 78 36536 1638 0 Data[5]
rlabel metal4 39104 78 40664 1638 0 gnde!
rlabel metal4 45728 6616 47288 8176 0 Data[6]
rlabel metal4 45728 11346 47288 12906 0 Data[7]
rlabel metal4 45728 16076 47288 17636 0 Data[8]
rlabel metal4 45728 20806 47288 22366 0 gnde!
rlabel metal4 45728 25536 47288 27096 0 GND!
rlabel metal4 45728 30266 47288 31826 0 Data[9]
rlabel metal4 45728 34996 47288 36556 0 Data[10]
rlabel metal4 45728 39726 47288 41286 0 Data[11]
rlabel metal4 39104 46264 40664 47824 0 vdde!
rlabel metal4 34976 46264 36536 47824 0 Data[12]
rlabel metal4 30848 46264 32408 47824 0 Data[13]
rlabel metal4 26720 46264 28280 47824 0 Data[14]
rlabel metal4 22592 46264 24152 47824 0 gnde!
rlabel metal4 18464 46264 20024 47824 0 Data[15]
rlabel metal4 14336 46264 15896 47824 0 ALE
rlabel metal4 10208 46264 11768 47824 0 nME
rlabel metal4 6080 46264 7640 47824 0 nWait
rlabel metal4 -544 39726 1016 41286 0 nOE
rlabel metal4 -544 34996 1016 36556 0 RnW
rlabel metal4 -544 30266 1016 31826 0 SDO
rlabel metal4 -544 25536 1016 27096 0 Vdd!
rlabel metal4 -544 20806 1016 22366 0 SDI
rlabel metal4 -544 16076 1016 17636 0 Test
rlabel metal4 -544 11346 1016 12906 0 Clock
rlabel metal4 -544 6616 1016 8176 0 nReset
<< end >>
