magic
tech c035u
timestamp 1393856096
<< error_s >>
rect 3935 2045 3949 2050
use ALUDecoder ALUDecoder_0
timestamp 1393855782
transform 1 0 0 0 1 2040
box 0 0 7224 1481
use ALU ALU_1
timestamp 1393852311
transform 1 0 0 0 1 998
box 0 0 6648 1042
use LLIcell_U LLIcell_U_0
timestamp 1393855556
transform 1 0 6648 0 1 998
box 0 0 192 1042
use ALU ALU_0
timestamp 1393852311
transform 1 0 0 0 1 -44
box 0 0 6648 1042
use LLIcell_L LLIcell_L_0
timestamp 1393855517
transform 1 0 6648 0 1 -44
box 0 0 192 1042
<< end >>
