magic
tech c035u
timestamp 1396394133
<< metal1 >>
rect 0 1094 23 1104
rect 0 97 23 107
rect 973 95 1837 105
rect 0 29 887 39
rect 901 29 1103 39
rect 1117 29 1463 39
rect 1477 29 1837 39
<< m2contact >>
rect 23 1092 37 1106
rect 23 95 37 109
rect 959 93 973 107
rect 887 27 901 41
rect 1103 27 1117 41
rect 1463 27 1477 41
<< metal2 >>
rect 24 911 36 1092
rect 72 911 84 1111
rect 600 911 756 923
rect 816 911 828 1111
rect 1032 911 1044 1111
rect 1224 982 1236 1111
rect 1176 970 1236 982
rect 1176 911 1188 970
rect 1272 960 1284 1111
rect 1224 948 1284 960
rect 1224 911 1236 948
rect 1320 938 1332 1111
rect 1272 926 1332 938
rect 1272 911 1284 926
rect 1392 911 1404 1111
rect 1632 911 1832 1111
rect 24 109 36 112
rect 72 0 84 112
rect 816 0 828 112
rect 888 41 900 112
rect 960 107 972 200
rect 1032 0 1044 112
rect 1104 41 1116 112
rect 1176 0 1188 112
rect 1224 0 1236 112
rect 1272 0 1284 113
rect 1320 0 1332 112
rect 1392 0 1404 112
rect 1464 41 1476 112
rect 1632 0 1832 112
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 112
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 720 0 1 112
box 0 0 216 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 936 0 1 112
box 0 0 216 799
use rowcrosser rowcrosser_0
array 0 2 48 0 0 799
timestamp 1386086759
transform 1 0 1152 0 1 112
box 0 0 48 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 1296 0 1 112
box 0 0 216 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 1512 0 1 112
box 0 0 320 799
<< labels >>
rlabel metal2 816 1111 828 1111 5 AluEn
rlabel metal2 72 1111 84 1111 5 AluWe
rlabel metal1 0 1094 0 1104 3 AluOut
rlabel metal2 654 915 654 915 1 AluRegOut
rlabel metal1 0 97 0 107 3 AluOut
rlabel metal1 0 29 0 39 3 DataOut
rlabel metal1 1837 29 1837 39 7 DataOut
rlabel metal2 1320 1111 1332 1111 5 StatusReg[1]
rlabel metal2 1272 1111 1284 1111 5 StatusReg[2]
rlabel metal2 1224 1111 1236 1111 5 StatusReg[3]
rlabel metal2 1392 1111 1404 1111 5 StatusRegEn
rlabel metal2 1632 1111 1832 1111 5 GND!
rlabel metal2 1032 1111 1044 1111 5 MemEn
rlabel metal2 72 0 84 0 1 AluWe
rlabel metal2 816 0 828 0 1 AluEn
rlabel metal2 1224 0 1236 0 1 StatusReg[2]
rlabel metal2 1272 0 1284 0 1 StatusReg[1]
rlabel metal2 1320 0 1332 0 1 StatusReg[0]
rlabel metal2 1176 0 1188 0 1 StatusReg[3]
rlabel metal2 1392 0 1404 0 1 StatusRegEn
rlabel metal2 1632 0 1832 0 1 GND!
rlabel metal2 1032 0 1044 0 1 MemEn
rlabel metal1 1837 95 1837 105 7 DataIn
<< end >>
