magic
tech c035u
timestamp 1395569717
<< checkpaint >>
rect 0 0 27110 20800
rect 20800 -1257 27110 0
rect 20800 -1300 26696 -1257
<< metal1 >>
rect 19 20557 14582 20567
rect 42 20533 14775 20543
rect 65 20509 14967 20519
rect 88 20485 15159 20495
rect 111 20461 15351 20471
rect 134 20437 4166 20447
rect 157 20413 4598 20423
rect 180 20389 4982 20399
rect 203 20365 4214 20375
rect 226 20341 4646 20351
rect 249 20317 5030 20327
rect 272 20293 7170 20303
rect 295 20269 7146 20279
rect 7160 20269 22358 20279
rect 318 20245 7122 20255
rect 7136 20245 22550 20255
rect 341 20221 22670 20231
rect 364 20197 22790 20207
rect 23583 18848 23775 18858
rect 3100 18737 3111 18747
rect 0 17850 5 17860
rect 19 17850 370 17860
rect 0 17818 370 17828
rect 0 17784 370 17794
rect 3063 17784 3111 17794
rect 23583 17784 23775 17794
rect 3063 17762 3111 17772
rect 23583 17672 23775 17682
rect 3100 17561 3111 17571
rect 0 16674 28 16684
rect 42 16674 370 16684
rect 0 16642 370 16652
rect 0 16608 370 16618
rect 3063 16608 3111 16618
rect 23583 16608 23775 16618
rect 3063 16586 3111 16596
rect 23583 16496 23775 16506
rect 3100 16385 3111 16395
rect 0 15498 51 15508
rect 65 15498 370 15508
rect 0 15466 370 15476
rect 0 15432 370 15442
rect 3063 15432 3111 15442
rect 23583 15432 23775 15442
rect 3063 15410 3111 15420
rect 23583 15320 23775 15330
rect 3100 15209 3111 15219
rect 0 14322 74 14332
rect 88 14322 370 14332
rect 0 14290 370 14300
rect 0 14256 370 14266
rect 3063 14256 3111 14266
rect 23583 14256 23775 14266
rect 3063 14234 3111 14244
rect 23583 14144 23775 14154
rect 3100 14033 3111 14043
rect 0 13146 97 13156
rect 111 13146 370 13156
rect 0 13114 370 13124
rect 0 13080 370 13090
rect 3063 13080 3111 13090
rect 23583 13080 23775 13090
rect 3063 13058 3111 13068
rect 23583 12968 23775 12978
rect 3100 12857 3111 12867
rect 0 11970 120 11980
rect 134 11970 370 11980
rect 0 11938 370 11948
rect 0 11904 370 11914
rect 3063 11904 3111 11914
rect 23583 11904 23775 11914
rect 3063 11882 3111 11892
rect 23583 11792 23775 11802
rect 3100 11681 3111 11691
rect 0 10794 143 10804
rect 157 10794 370 10804
rect 0 10762 370 10772
rect 0 10728 370 10738
rect 3063 10728 3111 10738
rect 23583 10728 23775 10738
rect 3063 10706 3111 10716
rect 23583 10616 23775 10626
rect 3100 10505 3111 10515
rect 0 9618 166 9628
rect 180 9618 370 9628
rect 0 9586 370 9596
rect 0 9552 370 9562
rect 3063 9552 3111 9562
rect 23583 9552 23775 9562
rect 3063 9530 3111 9540
rect 23583 9440 23775 9450
rect 3100 9329 3111 9339
rect 0 8442 189 8452
rect 203 8442 370 8452
rect 0 8410 370 8420
rect 0 8376 370 8386
rect 3063 8376 3111 8386
rect 23583 8376 23775 8386
rect 3063 8354 3111 8364
rect 23583 8264 23775 8274
rect 3100 8153 3111 8163
rect 0 7266 212 7276
rect 226 7266 370 7276
rect 0 7234 370 7244
rect 0 7200 370 7210
rect 3063 7200 3111 7210
rect 23583 7200 23775 7210
rect 3063 7178 3111 7188
rect 23583 7088 23775 7098
rect 3100 6977 3111 6987
rect 0 6090 235 6100
rect 249 6090 370 6100
rect 0 6058 370 6068
rect 0 6024 370 6034
rect 3063 6024 3111 6034
rect 23583 6024 23775 6034
rect 3063 6002 3111 6012
rect 23583 5912 23775 5922
rect 3100 5801 3111 5811
rect 0 4914 258 4924
rect 272 4914 370 4924
rect 0 4882 370 4892
rect 0 4848 370 4858
rect 3063 4848 3111 4858
rect 23583 4848 23775 4858
rect 3063 4826 3111 4836
rect 23583 4736 23775 4746
rect 3100 4625 3111 4635
rect 0 3738 281 3748
rect 295 3738 370 3748
rect 0 3706 370 3716
rect 0 3672 370 3682
rect 3063 3672 3111 3682
rect 23583 3672 23775 3682
rect 3063 3650 3111 3660
rect 23583 3560 23775 3570
rect 3100 3449 3111 3459
rect 0 2562 304 2572
rect 318 2562 370 2572
rect 0 2530 370 2540
rect 0 2496 370 2506
rect 3063 2496 3111 2506
rect 23583 2496 23775 2506
rect 3063 2474 3111 2484
rect 23583 2384 23775 2394
rect 3100 2273 3111 2283
rect 0 1386 327 1396
rect 341 1386 370 1396
rect 0 1354 370 1364
rect 0 1320 370 1330
rect 3063 1320 3111 1330
rect 23583 1320 23775 1330
rect 3063 1298 3111 1308
rect 23583 1208 23775 1218
rect 3100 1097 3111 1107
rect 0 210 350 220
rect 364 210 370 220
rect 0 178 370 188
rect 0 144 370 154
rect 3063 144 3111 154
rect 23583 144 23775 154
rect 3063 122 3111 132
rect 2060 29 17270 39
rect 17284 29 19934 39
rect 19948 29 19981 39
rect 19995 29 20030 39
rect 20044 29 20078 39
rect 20092 29 20126 39
rect 20140 29 20174 39
rect 20188 29 20222 39
rect 20236 29 20270 39
rect 20284 29 20582 39
rect 20596 29 20630 39
rect 20644 29 20677 39
rect 20691 29 20726 39
rect 20740 29 21038 39
rect 21052 29 21086 39
rect 21100 29 21470 39
rect 21484 29 25191 39
rect 575 8 3326 18
<< m2contact >>
rect 5 20555 19 20569
rect 14582 20556 14596 20570
rect 28 20531 42 20545
rect 14775 20531 14789 20545
rect 51 20507 65 20521
rect 14967 20507 14981 20521
rect 74 20483 88 20497
rect 15159 20483 15173 20497
rect 97 20459 111 20473
rect 15351 20459 15365 20474
rect 120 20435 134 20449
rect 4166 20435 4180 20449
rect 143 20411 157 20425
rect 4598 20411 4612 20425
rect 166 20387 180 20401
rect 4982 20387 4996 20401
rect 189 20363 203 20377
rect 4214 20363 4228 20377
rect 212 20339 226 20353
rect 4646 20339 4660 20353
rect 235 20315 249 20329
rect 5030 20315 5044 20329
rect 258 20291 272 20305
rect 7170 20291 7184 20305
rect 281 20267 295 20281
rect 7146 20267 7160 20281
rect 22358 20267 22372 20281
rect 304 20243 318 20257
rect 7122 20243 7136 20257
rect 22550 20242 22564 20256
rect 327 20219 341 20233
rect 22670 20219 22684 20233
rect 350 20195 364 20209
rect 22790 20195 22804 20209
rect 3086 18735 3100 18749
rect 5 17848 19 17862
rect 3086 17559 3100 17573
rect 28 16672 42 16686
rect 3086 16383 3100 16397
rect 51 15496 65 15510
rect 3086 15207 3100 15221
rect 74 14320 88 14334
rect 3086 14031 3100 14045
rect 97 13144 111 13158
rect 3086 12855 3100 12869
rect 120 11968 134 11982
rect 3086 11679 3100 11693
rect 143 10792 157 10806
rect 3086 10503 3100 10517
rect 166 9616 180 9630
rect 3086 9327 3100 9341
rect 189 8440 203 8454
rect 3086 8151 3100 8165
rect 212 7264 226 7278
rect 3086 6975 3100 6989
rect 235 6088 249 6102
rect 3086 5799 3100 5813
rect 258 4912 272 4926
rect 3086 4623 3100 4637
rect 281 3736 295 3750
rect 3086 3447 3100 3461
rect 304 2560 318 2574
rect 3086 2271 3100 2285
rect 327 1384 341 1398
rect 3086 1095 3100 1109
rect 350 208 364 222
rect 17270 27 17284 41
rect 19934 27 19948 41
rect 19981 27 19995 41
rect 20030 27 20044 41
rect 20078 27 20092 41
rect 20126 27 20140 41
rect 20174 27 20188 41
rect 20222 27 20236 41
rect 20270 27 20284 41
rect 20582 27 20596 41
rect 20630 27 20644 41
rect 20677 27 20691 41
rect 20726 27 20740 41
rect 21038 27 21052 41
rect 21086 27 21100 41
rect 21470 27 21484 41
rect 25191 27 25205 41
rect 561 6 575 20
rect 3326 5 3340 19
<< metal2 >>
rect 6 17862 18 20555
rect 29 16686 41 20531
rect 52 15510 64 20507
rect 75 14334 87 20483
rect 98 13158 110 20459
rect 121 11982 133 20435
rect 144 10806 156 20411
rect 167 9630 179 20387
rect 190 8454 202 20363
rect 213 7278 225 20339
rect 236 6102 248 20315
rect 259 4926 271 20291
rect 282 3750 294 20267
rect 305 2574 317 20243
rect 328 1398 340 20219
rect 351 222 363 20195
rect 375 20186 575 20572
rect 591 20186 603 20572
rect 615 20186 627 20572
rect 639 20186 651 20572
rect 663 20186 675 20572
rect 4143 20186 4155 20572
rect 4167 20186 4179 20435
rect 4215 20186 4227 20363
rect 4383 20186 4395 20572
rect 4599 20186 4611 20411
rect 4647 20186 4659 20339
rect 4983 20186 4995 20387
rect 5031 20186 5043 20315
rect 5343 20186 5355 20572
rect 5535 20186 5547 20572
rect 6569 20186 6581 20572
rect 7123 20186 7135 20243
rect 7147 20186 7159 20267
rect 7171 20186 7183 20291
rect 14560 20186 14572 20572
rect 14584 20186 14596 20556
rect 14776 20186 14788 20531
rect 14824 20186 14836 20572
rect 14968 20186 14980 20507
rect 15160 20186 15172 20483
rect 15352 20186 15364 20459
rect 15544 20186 15556 20572
rect 17343 20186 17355 20572
rect 17535 20186 17547 20572
rect 17607 20186 17619 20572
rect 17703 20186 17715 20572
rect 22359 20186 22371 20267
rect 22551 20186 22563 20242
rect 22671 20186 22683 20219
rect 22791 20186 22803 20195
rect 25191 20186 25391 20572
rect 23631 18842 23643 18865
rect 3087 18665 3099 18735
rect 23631 17666 23643 17800
rect 3087 17489 3099 17559
rect 23631 16490 23643 16624
rect 3087 16313 3099 16383
rect 23631 15314 23643 15448
rect 3087 15137 3099 15207
rect 23631 14138 23643 14272
rect 3087 13961 3099 14031
rect 23631 12962 23643 13096
rect 3087 12785 3099 12855
rect 23631 11786 23643 11920
rect 3087 11609 3099 11679
rect 23631 10610 23643 10744
rect 3087 10433 3099 10503
rect 23631 9434 23643 9568
rect 3087 9257 3099 9327
rect 23631 8258 23643 8392
rect 3087 8081 3099 8151
rect 23631 7082 23643 7216
rect 3087 6905 3099 6975
rect 23631 5906 23643 6040
rect 3087 5729 3099 5799
rect 23631 4730 23643 4864
rect 3087 4553 3099 4623
rect 23631 3554 23643 3688
rect 3087 3377 3099 3447
rect 23631 2378 23643 2512
rect 3087 2201 3099 2271
rect 23631 1202 23643 1336
rect 3087 1025 3099 1095
rect 23631 49 23643 160
rect 375 20 575 49
rect 375 6 561 20
rect 375 0 575 6
rect 591 0 603 49
rect 615 0 627 49
rect 639 0 651 49
rect 663 0 675 49
rect 1935 0 1947 49
rect 2127 0 2139 49
rect 2919 0 2931 49
rect 3327 19 3339 49
rect 3471 0 3483 49
rect 3687 0 3699 49
rect 4431 0 4443 49
rect 4599 0 4611 49
rect 4983 0 4995 49
rect 5175 0 5187 49
rect 5391 0 5403 49
rect 6135 0 6147 49
rect 6303 0 6315 49
rect 15711 0 15723 49
rect 15903 0 15915 49
rect 16143 0 16155 49
rect 16791 43 16803 49
rect 16983 43 16995 49
rect 16791 31 16995 43
rect 17271 41 17283 49
rect 19935 41 19947 49
rect 19983 41 19995 49
rect 20031 41 20043 49
rect 20079 41 20091 49
rect 20127 41 20139 49
rect 20175 41 20187 49
rect 20223 41 20235 49
rect 20271 41 20283 49
rect 20583 41 20595 49
rect 20631 41 20643 49
rect 20679 41 20691 49
rect 20727 41 20739 49
rect 21039 41 21051 49
rect 21087 41 21099 49
rect 21471 41 21483 49
rect 23847 0 23859 49
rect 24591 0 24603 49
rect 24735 0 24747 49
rect 24783 0 24795 49
rect 24831 0 24843 49
rect 24879 0 24891 49
rect 24951 0 24963 49
rect 25191 41 25391 49
rect 25205 27 25391 41
rect 25191 0 25391 27
use slice17 slice17_0
timestamp 1395569125
transform 1 0 375 0 1 18865
box 0 0 25016 1321
use leftbuf_slice leftbuf_slice_0
array 0 0 1685 0 15 1176
timestamp 1394551156
transform 1 0 370 0 1 55
box 0 -6 1685 1170
use IrAA IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 2055 0 1 9568
box 0 -111 1008 1065
use tielow tielow_0
timestamp 1386086605
transform 1 0 3063 0 1 17866
box 0 0 48 799
use tielow tielow_1
timestamp 1386086605
transform 1 0 3063 0 1 16690
box 0 0 48 799
use tielow tielow_2
timestamp 1386086605
transform 1 0 3063 0 1 15514
box 0 0 48 799
use tielow tielow_3
timestamp 1386086605
transform 1 0 3063 0 1 14338
box 0 0 48 799
use tielow tielow_4
timestamp 1386086605
transform 1 0 3063 0 1 13162
box 0 0 48 799
use tielow tielow_5
timestamp 1386086605
transform 1 0 3063 0 1 11986
box 0 0 48 799
use tielow tielow_6
timestamp 1386086605
transform 1 0 3063 0 1 10810
box 0 0 48 799
use tielow tielow_7
timestamp 1386086605
transform 1 0 3063 0 1 9634
box 0 0 48 799
use IrBA IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 2055 0 1 6040
box 0 -111 1008 1065
use tielow tielow_8
timestamp 1386086605
transform 1 0 3063 0 1 8458
box 0 0 48 799
use tielow tielow_9
timestamp 1386086605
transform 1 0 3063 0 1 7282
box 0 0 48 799
use tielow tielow_10
timestamp 1386086605
transform 1 0 3063 0 1 6106
box 0 0 48 799
use IrBB IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 2055 0 1 161
box 0 -112 1008 1064
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 3063 0 1 4930
box 0 0 48 799
use tielow tielow_12
timestamp 1386086605
transform 1 0 3063 0 1 3754
box 0 0 48 799
use tielow tielow_13
timestamp 1386086605
transform 1 0 3063 0 1 2578
box 0 0 48 799
use tielow tielow_14
timestamp 1386086605
transform 1 0 3063 0 1 1402
box 0 0 48 799
use tielow tielow_15
timestamp 1386086605
transform 1 0 3063 0 1 226
box 0 0 48 799
use Datapath_slice Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394725603
transform 1 0 3111 0 1 49
box 0 0 20472 1176
use LLIcell_U LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1394841956
transform 1 0 23583 0 1 9568
box 0 0 192 1042
use LLIcell_L LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23583 0 1 160
box 0 0 192 1042
use Datapath_end_high Datapath_end_high_0
array 0 0 1621 0 11 1176
timestamp 1395569595
transform 1 0 23775 0 1 4753
box 0 0 1621 1176
use Datapath_end_low Datapath_end_low_0
array 0 0 1616 0 3 1176
timestamp 1395569514
transform 1 0 23775 0 1 49
box 0 0 1621 1176
<< labels >>
rlabel metal1 23679 1214 23679 1214 1 Aluout[0]
rlabel metal2 11 20260 11 20260 1 Ir[15]
rlabel metal2 35 20259 35 20259 1 Ir[14]
rlabel metal2 58 20259 58 20259 1 Ir[13]
rlabel metal2 81 20260 81 20260 1 Ir[12]
rlabel metal2 104 20260 104 20260 1 Ir[11]
rlabel metal2 127 20259 127 20259 1 Ir[10]
rlabel metal2 150 20260 150 20260 1 Ir[9]
rlabel metal2 173 20260 173 20260 1 Ir[8]
rlabel metal2 196 20262 196 20262 1 Ir[7]
rlabel metal2 219 20263 219 20263 1 Ir[6]
rlabel metal2 242 20264 242 20264 1 Ir[5]
rlabel metal2 265 20265 265 20265 1 Ir[4]
rlabel metal2 288 20264 288 20264 1 Ir[3]
rlabel metal2 22797 20190 22797 20190 1 Ir[0]
rlabel metal2 22676 20212 22676 20212 1 Ir[1]
rlabel metal2 22556 20237 22556 20237 1 Ir[2]
rlabel metal2 22365 20262 22365 20262 1 Ir[3]
rlabel metal2 14973 20501 14973 20501 1 Ir[13]
rlabel metal2 15166 20477 15166 20477 1 Ir[12]
rlabel metal2 15358 20452 15358 20452 1 Ir[11]
rlabel metal2 14780 20524 14780 20524 1 Ir[14]
rlabel metal2 14589 20549 14589 20549 1 Ir[15]
rlabel metal2 7127 20235 7127 20235 1 Ir[2]
rlabel metal2 7153 20259 7153 20259 1 Ir[3]
rlabel metal2 7176 20283 7176 20283 1 Ir[4]
rlabel metal2 4221 20355 4221 20355 1 Ir[7]
rlabel metal2 4172 20428 4172 20428 1 Ir[10]
rlabel metal2 4653 20332 4653 20332 1 Ir[6]
rlabel metal2 4604 20403 4604 20403 1 Ir[9]
rlabel metal2 4988 20380 4988 20380 1 Ir[8]
rlabel metal2 5038 20309 5038 20309 1 Ir[5]
rlabel metal1 0 144 0 154 3 SysBus[0]
rlabel metal1 0 1320 0 1330 3 SysBus[1]
rlabel metal1 0 2496 0 2506 3 SysBus[2]
rlabel metal1 0 3672 0 3682 3 SysBus[3]
rlabel metal1 0 4848 0 4858 3 SysBus[4]
rlabel metal1 0 6024 0 6034 3 SysBus[5]
rlabel metal1 0 7200 0 7210 3 SysBus[6]
rlabel metal1 0 8376 0 8386 3 SysBus[7]
rlabel metal1 0 9552 0 9562 3 SysBus[8]
rlabel metal1 0 10728 0 10738 3 SysBus[9]
rlabel metal1 0 11904 0 11914 3 SysBus[10]
rlabel metal1 0 13080 0 13090 3 SysBus[11]
rlabel metal1 0 14256 0 14266 3 SysBus[12]
rlabel metal1 0 15432 0 15442 3 SysBus[13]
rlabel metal1 0 16608 0 16618 3 SysBus[14]
rlabel metal1 0 17784 0 17794 3 SysBus[15]
rlabel metal1 0 210 0 220 3 Ir[0]
rlabel metal1 0 1386 0 1396 3 Ir[1]
rlabel metal1 0 2562 0 2572 3 Ir[2]
rlabel metal1 0 3738 0 3748 3 Ir[3]
rlabel metal1 0 4914 0 4924 3 Ir[4]
rlabel metal1 0 6090 0 6100 3 Ir[5]
rlabel metal1 0 7266 0 7276 3 Ir[6]
rlabel metal1 0 8442 0 8452 3 Ir[7]
rlabel metal1 0 9618 0 9628 3 Ir[8]
rlabel metal1 0 10794 0 10804 3 Ir[9]
rlabel metal1 0 11970 0 11980 3 Ir[10]
rlabel metal1 0 13146 0 13156 3 Ir[11]
rlabel metal1 0 14322 0 14332 3 Ir[12]
rlabel metal1 0 15498 0 15508 3 Ir[13]
rlabel metal1 0 16674 0 16684 3 Ir[14]
rlabel metal1 0 17850 0 17860 3 Ir[15]
rlabel metal1 0 178 0 188 3 DataIn[0]
rlabel metal1 0 17818 0 17828 3 DataIn[15]
rlabel metal1 0 16642 0 16652 3 DataIn[14]
rlabel metal1 0 15466 0 15476 3 DataIn[13]
rlabel metal1 0 14290 0 14300 3 DataIn[12]
rlabel metal1 0 13114 0 13124 3 DataIn[11]
rlabel metal1 0 11938 0 11948 3 DataIn[10]
rlabel metal1 0 10762 0 10772 3 DataIn[9]
rlabel metal1 0 9586 0 9596 3 DataIn[8]
rlabel metal1 0 8410 0 8420 3 DataIn[7]
rlabel metal1 0 7234 0 7244 3 DataIn[6]
rlabel metal1 0 6058 0 6068 3 DataIn[5]
rlabel metal1 0 4882 0 4892 3 DataIn[4]
rlabel metal1 0 3706 0 3716 3 DataIn[3]
rlabel metal1 0 2530 0 2540 3 DataIn[2]
rlabel metal1 0 1354 0 1364 3 DataIn[1]
rlabel metal2 6569 20572 6581 20572 5 RegWe
rlabel metal2 591 20572 603 20572 5 SDO
rlabel metal2 375 20572 575 20572 5 Vdd!
rlabel metal2 663 20572 675 20572 1 nReset
rlabel metal2 639 20572 651 20572 1 Clock
rlabel metal2 615 20572 627 20572 1 Test
rlabel metal2 17703 20572 17715 20572 5 Flags[0]
rlabel metal2 17607 20572 17619 20572 5 Flags[3]
rlabel metal2 17535 20572 17547 20572 5 Flags[1]
rlabel metal2 17343 20572 17355 20572 5 Flags[2]
rlabel metal2 14824 20572 14836 20572 5 AluOR[0]
rlabel metal2 14560 20572 14572 20572 5 AluOR[1]
rlabel metal2 15544 20572 15556 20572 5 CFlag
rlabel metal2 4143 20572 4155 20572 5 Rs1Sel[0]
rlabel metal2 4383 20572 4395 20572 5 Rs1Sel[1]
rlabel metal2 5343 20572 5355 20572 5 RwSel[0]
rlabel metal2 5535 20572 5547 20572 5 RwSel[1]
rlabel metal2 3471 0 3483 0 1 LrSel
rlabel metal2 3687 0 3699 0 1 LrWe
rlabel metal2 4431 0 4443 0 1 LrEn
rlabel metal2 4599 0 4611 0 1 PcSel[0]
rlabel metal2 4983 0 4995 0 1 PcSel[1]
rlabel metal2 23847 0 23859 0 1 AluWe
rlabel metal2 24591 0 24603 0 1 AluEn
rlabel metal2 375 0 575 0 1 Vdd!
rlabel metal2 591 0 603 0 1 SDI
rlabel metal2 615 0 627 0 1 Test
rlabel metal2 639 0 651 0 1 Clock
rlabel metal2 663 0 675 0 1 nReset
rlabel metal2 2919 0 2931 0 1 ImmSel
rlabel metal2 2127 0 2139 0 1 IrWe
rlabel metal2 1935 0 1947 0 1 MemEn
rlabel metal2 5391 0 5403 0 1 PcWe
rlabel metal2 5175 0 5187 0 1 PcSel[2]
rlabel metal2 6135 0 6147 0 1 PcEn
rlabel metal2 6303 0 6315 0 1 WdSel
rlabel metal2 15711 0 15723 0 1 Op1Sel
rlabel metal2 15903 0 15915 0 1 Op2Sel[0]
rlabel metal2 16143 0 16155 0 1 Op2Sel[1]
rlabel metal2 25191 0 25391 0 1 GND!
rlabel metal2 25191 20572 25391 20572 1 GND!
rlabel metal2 24735 0 24747 0 1 StatusReg[0]
rlabel metal2 24783 0 24795 0 1 StatusReg[1]
rlabel metal2 24831 0 24843 0 1 StatusReg[2]
rlabel metal2 24879 0 24891 0 1 StatusReg[3]
rlabel metal2 24951 0 24963 0 1 StatusRegEn
<< end >>
