../behavioural/control.sv