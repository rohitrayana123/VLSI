../../Design/Implementation/verilog/behavioural/aludecoder.sv