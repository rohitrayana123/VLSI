magic
tech c035u
timestamp 1395569514
<< metal1 >>
rect 0 1159 23 1169
rect 0 162 23 172
rect 0 95 887 105
rect 901 95 1247 105
rect 1261 95 1621 105
<< m2contact >>
rect 23 1157 37 1171
rect 23 160 37 174
rect 887 93 901 107
rect 1247 92 1261 106
<< metal2 >>
rect 24 976 36 1157
rect 72 976 84 1176
rect 600 976 756 988
rect 816 976 828 1176
rect 1008 1047 1020 1176
rect 960 1035 1020 1047
rect 960 976 972 1035
rect 1056 1025 1068 1176
rect 1008 1013 1068 1025
rect 1008 976 1020 1013
rect 1104 1003 1116 1176
rect 1056 991 1116 1003
rect 1056 976 1068 991
rect 1176 976 1188 1176
rect 1416 976 1616 1176
rect 24 174 36 177
rect 72 0 84 177
rect 816 0 828 177
rect 888 107 900 177
rect 960 0 972 177
rect 1008 0 1020 177
rect 1056 0 1068 178
rect 1104 0 1116 177
rect 1176 0 1188 177
rect 1248 106 1260 177
rect 1416 0 1616 177
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 177
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 720 0 1 177
box 0 0 216 799
use rowcrosser rowcrosser_0
array 0 2 48 0 0 799
timestamp 1386086759
transform 1 0 936 0 1 177
box 0 0 48 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 1080 0 1 177
box 0 0 216 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 1296 0 1 177
box 0 0 320 799
<< labels >>
rlabel metal2 816 1176 828 1176 5 AluEn
rlabel metal2 72 0 84 0 1 AluWe
rlabel metal2 72 1176 84 1176 5 AluWe
rlabel metal1 0 1159 0 1169 3 AluOut
rlabel metal2 654 980 654 980 1 AluRegOut
rlabel metal2 1416 1176 1616 1176 5 GND!
rlabel metal2 1416 0 1616 0 1 GND!
rlabel metal2 960 0 972 0 1 StatusReg[0]
rlabel metal2 1008 0 1020 0 1 StatusReg[1]
rlabel metal2 1056 0 1068 0 1 StatusReg[2]
rlabel metal2 1104 0 1116 0 1 StatusReg[3]
rlabel metal2 1176 0 1188 0 1 StatusRegEn
rlabel metal2 1008 1176 1020 1176 5 StatusReg[0]
rlabel metal2 1056 1176 1068 1176 5 StatusReg[1]
rlabel metal2 1104 1176 1116 1176 5 StatusReg[2]
rlabel metal2 1176 1176 1188 1176 5 StatusRegEn
rlabel metal1 1621 95 1621 105 7 DataOut
rlabel metal1 0 95 0 105 3 DataOut
rlabel metal2 816 0 828 0 1 AluEn
rlabel metal1 0 162 0 172 3 AluOut
<< end >>
