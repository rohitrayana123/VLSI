../../../Design/Implementation/verilog/behavioural/signExtend.sv