magic
tech c035u
timestamp 1396952988
<< metal1 >>
rect 21120 39730 21130 39773
rect 21168 39730 21178 39773
rect 21120 39720 21178 39730
rect 21120 39226 21130 39720
rect 21216 39253 21226 39773
rect 24552 39757 24562 39773
rect 24600 39730 24610 39773
rect 28080 39757 28090 39773
rect 21480 39720 24610 39730
rect 21480 39706 21490 39720
rect 28128 39730 28138 39773
rect 24637 39720 28138 39730
rect 31584 39730 31594 39773
rect 31632 39757 31642 39773
rect 31776 39757 31786 39773
rect 38640 39730 38650 39773
rect 38688 39757 38698 39773
rect 38832 39757 38842 39773
rect 42168 39730 42178 39773
rect 42216 39757 42226 39773
rect 42360 39757 42370 39773
rect 45696 39733 45706 39773
rect 45744 39757 45754 39773
rect 45888 39757 45898 39773
rect 31584 39720 45695 39730
rect 45720 39720 46991 39730
rect 21456 39696 21490 39706
rect 21456 39685 21466 39696
rect 21517 39696 24551 39706
rect 24565 39696 28079 39706
rect 45720 39706 45730 39720
rect 31645 39696 45730 39706
rect 46837 39696 47050 39706
rect 21493 39672 24623 39682
rect 21432 39648 21503 39658
rect 21432 39253 21442 39648
rect 21456 39253 21466 39623
rect 21480 39253 21490 39623
rect 28080 39589 28090 39695
rect 38701 39672 47015 39682
rect 47040 39682 47050 39696
rect 47040 39672 47063 39682
rect 31776 39589 31786 39671
rect 38845 39648 47087 39658
rect 45901 39624 47122 39634
rect 42216 39589 42226 39623
rect 42360 39589 42370 39623
rect 45696 39610 45706 39623
rect 47112 39613 47122 39624
rect 45696 39600 47039 39610
rect 45757 39576 45767 39586
rect 47029 39576 47135 39586
rect 27888 39552 47015 39562
rect 27888 39469 27898 39552
rect 47125 39552 47159 39562
rect 45757 39528 46871 39538
rect 47005 39528 47207 39538
rect 28080 39469 28090 39527
rect 31776 39469 31786 39527
rect 38869 39504 46991 39514
rect 47029 39504 47231 39514
rect 38664 39480 47015 39490
rect 38664 39469 38674 39480
rect 47053 39480 47255 39490
rect 39037 39456 47183 39466
rect 47221 39456 47279 39466
rect 25464 39432 47039 39442
rect 21120 39216 21514 39226
rect 21408 39192 21431 39202
rect 20207 38832 20266 38842
rect 20256 38818 20266 38832
rect 21216 38821 21226 39191
rect 20256 38808 20279 38818
rect 21408 38794 21418 39192
rect 21504 39202 21514 39216
rect 21504 39192 22007 39202
rect 20207 38784 21418 38794
rect 21432 39168 22138 39178
rect 20256 34810 20266 38784
rect 20280 34837 20290 38759
rect 20256 34800 20314 34810
rect 20207 34776 20266 34786
rect 20256 34765 20266 34776
rect 20304 34738 20314 34800
rect 20207 34728 20314 34738
rect 20256 30781 20266 34703
rect 20280 30781 20290 34703
rect 20304 30781 20314 34728
rect 21216 30781 21226 38759
rect 21432 30754 21442 39168
rect 22128 39157 22138 39168
rect 25464 39157 25474 39432
rect 47101 39432 47303 39442
rect 26856 39408 47111 39418
rect 26856 39373 26866 39408
rect 47173 39408 47338 39418
rect 47328 39397 47338 39408
rect 36144 39384 47218 39394
rect 36144 39373 36154 39384
rect 47208 39373 47218 39384
rect 36877 39360 47159 39370
rect 47256 39370 47266 39383
rect 47256 39360 47351 39370
rect 26664 39336 47255 39346
rect 26664 39277 26674 39336
rect 47293 39336 47375 39346
rect 35880 39312 47087 39322
rect 26856 39277 26866 39311
rect 27888 39277 27898 39311
rect 28080 39277 28090 39311
rect 31776 39277 31786 39311
rect 35880 39277 35890 39312
rect 47149 39312 47399 39322
rect 38928 39288 47279 39298
rect 38928 39277 38938 39288
rect 47317 39288 47423 39298
rect 42373 39264 45743 39274
rect 45781 39264 47314 39274
rect 47304 39253 47314 39264
rect 47389 39264 47447 39274
rect 25704 39240 47135 39250
rect 25704 39157 25714 39240
rect 47352 39250 47362 39263
rect 47352 39240 47506 39250
rect 31789 39216 47482 39226
rect 26664 39157 26674 39215
rect 26856 39157 26866 39215
rect 27888 39157 27898 39215
rect 28080 39178 28090 39215
rect 42229 39192 46858 39202
rect 28080 39168 46823 39178
rect 46848 39178 46858 39192
rect 46885 39192 47386 39202
rect 46848 39168 47362 39178
rect 46824 39157 46834 39167
rect 20207 30744 21442 30754
rect 20304 30706 20314 30719
rect 20207 30696 20314 30706
rect 20256 26794 20266 30671
rect 20280 26821 20290 30671
rect 20256 26784 20314 26794
rect 20207 26760 20266 26770
rect 20256 22834 20266 26760
rect 20280 22861 20290 26759
rect 20304 22861 20314 26784
rect 20256 22824 20338 22834
rect 20207 22800 20266 22810
rect 20256 19594 20266 22800
rect 20280 19618 20290 22799
rect 20304 19645 20314 22799
rect 20328 19642 20338 22824
rect 21216 19645 21226 30719
rect 21456 19666 21466 39143
rect 21445 19656 21466 19666
rect 20328 19632 21119 19642
rect 21480 19642 21490 39143
rect 46992 36469 47002 39143
rect 47016 36469 47026 39143
rect 47040 36469 47050 39143
rect 47064 36469 47074 39143
rect 47088 36469 47098 39143
rect 47112 36469 47122 39143
rect 47136 36469 47146 39143
rect 47160 36469 47170 39143
rect 47184 36469 47194 39143
rect 47208 36469 47218 39143
rect 47232 36469 47242 39143
rect 47256 36469 47266 39143
rect 47280 36469 47290 39143
rect 47304 36469 47314 39143
rect 47328 36469 47338 39143
rect 47352 36469 47362 39168
rect 47376 36469 47386 39192
rect 47400 36469 47410 39191
rect 47424 36469 47434 39191
rect 47448 36469 47458 39191
rect 47472 36442 47482 39216
rect 47496 39034 47506 39240
rect 47496 39024 50307 39034
rect 50256 39013 50266 39024
rect 50232 38976 50307 38986
rect 50232 38866 50242 38976
rect 50256 38869 50266 38951
rect 46968 36440 47482 36442
rect 46943 36432 47482 36440
rect 50208 38856 50242 38866
rect 46943 36430 46978 36432
rect 46943 36370 46978 36374
rect 47448 36370 47458 36407
rect 46943 36364 47458 36370
rect 46968 36360 47458 36364
rect 46992 35365 47002 36335
rect 47016 35365 47026 36335
rect 47040 35365 47050 36335
rect 47064 35365 47074 36335
rect 47088 35365 47098 36335
rect 47112 35365 47122 36335
rect 47136 35365 47146 36335
rect 47160 35365 47170 36335
rect 47184 35365 47194 36335
rect 47208 35365 47218 36335
rect 47232 35365 47242 36335
rect 47256 35365 47266 36335
rect 47280 35365 47290 36335
rect 47304 35365 47314 36335
rect 47328 35365 47338 36335
rect 47352 35365 47362 36335
rect 47376 35365 47386 36335
rect 47400 35365 47410 36335
rect 47424 35338 47434 36335
rect 46968 35329 47434 35338
rect 46943 35328 47434 35329
rect 46943 35319 46978 35328
rect 47400 35266 47410 35303
rect 46968 35263 47410 35266
rect 46943 35256 47410 35263
rect 46943 35253 46978 35256
rect 46992 34237 47002 35231
rect 47016 34237 47026 35231
rect 47040 34237 47050 35231
rect 47064 34237 47074 35231
rect 47088 34237 47098 35231
rect 47112 34237 47122 35231
rect 47136 34237 47146 35231
rect 47160 34237 47170 35231
rect 47184 34237 47194 35231
rect 47208 34237 47218 35231
rect 47232 34237 47242 35231
rect 47256 34237 47266 35231
rect 47280 34237 47290 35231
rect 47304 34237 47314 35231
rect 47328 34237 47338 35231
rect 47352 34237 47362 35231
rect 46943 34210 46978 34218
rect 47376 34210 47386 35231
rect 50208 34978 50218 38856
rect 50232 38832 50307 38842
rect 50232 34981 50242 38832
rect 50256 35002 50266 38807
rect 50256 34992 50307 35002
rect 50256 34981 50266 34992
rect 50184 34968 50218 34978
rect 50184 34861 50194 34968
rect 50208 34944 50307 34954
rect 50208 34861 50218 34944
rect 50232 34834 50242 34919
rect 50256 34837 50266 34919
rect 46943 34208 47386 34210
rect 46968 34200 47386 34208
rect 50160 34824 50242 34834
rect 46943 34142 46978 34152
rect 46968 34138 46978 34142
rect 47352 34138 47362 34175
rect 46968 34128 47362 34138
rect 46992 33133 47002 34103
rect 47016 33133 47026 34103
rect 47040 33133 47050 34103
rect 47064 33133 47074 34103
rect 47088 33133 47098 34103
rect 47112 33133 47122 34103
rect 47136 33133 47146 34103
rect 47160 33133 47170 34103
rect 47184 33133 47194 34103
rect 47208 33133 47218 34103
rect 47232 33133 47242 34103
rect 47256 33133 47266 34103
rect 47280 33133 47290 34103
rect 47304 33133 47314 34103
rect 46943 33106 46978 33107
rect 47328 33106 47338 34103
rect 46943 33097 47338 33106
rect 46968 33096 47338 33097
rect 46943 33034 46978 33041
rect 47304 33034 47314 33071
rect 46943 33031 47314 33034
rect 46968 33024 47314 33031
rect 46992 32029 47002 32999
rect 47016 32029 47026 32999
rect 47040 32029 47050 32999
rect 47064 32029 47074 32999
rect 47088 32029 47098 32999
rect 47112 32029 47122 32999
rect 47136 32029 47146 32999
rect 47160 32029 47170 32999
rect 47184 32029 47194 32999
rect 47208 32029 47218 32999
rect 47232 32029 47242 32999
rect 47256 32029 47266 32999
rect 47280 32029 47290 32999
rect 50160 32002 50170 34824
rect 50232 34800 50307 34810
rect 46968 31996 50170 32002
rect 46943 31992 50170 31996
rect 46943 31986 46978 31992
rect 50184 31930 50194 34799
rect 46943 31920 50194 31930
rect 46992 30901 47002 31895
rect 47016 30901 47026 31895
rect 47040 30901 47050 31895
rect 47064 30901 47074 31895
rect 47088 30901 47098 31895
rect 47112 30901 47122 31895
rect 47136 30901 47146 31895
rect 47160 30901 47170 31895
rect 47184 30901 47194 31895
rect 47208 30901 47218 31895
rect 47232 30901 47242 31895
rect 47256 30901 47266 31895
rect 47280 30901 47290 31895
rect 50208 30973 50218 34799
rect 50232 30946 50242 34800
rect 50256 30970 50266 34775
rect 50256 30960 50307 30970
rect 50256 30949 50266 30960
rect 50184 30936 50242 30946
rect 46943 30875 46978 30885
rect 46968 30874 46978 30875
rect 50184 30874 50194 30936
rect 50232 30912 50307 30922
rect 46968 30864 50194 30874
rect 50208 30826 50218 30911
rect 46968 30819 50218 30826
rect 46943 30816 50218 30819
rect 46943 30809 46978 30816
rect 50232 30805 50242 30912
rect 50256 30805 50266 30887
rect 46992 29797 47002 30791
rect 47016 29797 47026 30791
rect 47040 29797 47050 30791
rect 47064 29797 47074 30791
rect 47088 29797 47098 30791
rect 47112 29797 47122 30791
rect 47136 29797 47146 30791
rect 47160 29797 47170 30791
rect 47184 29797 47194 30791
rect 47208 29797 47218 30791
rect 47232 29797 47242 30791
rect 47256 29797 47266 30791
rect 47280 29797 47290 30791
rect 50208 30768 50307 30778
rect 46943 29770 46978 29774
rect 50208 29770 50218 30768
rect 46943 29764 50218 29770
rect 46968 29760 50218 29764
rect 46943 29698 46978 29708
rect 50232 29698 50242 30743
rect 46968 29688 50242 29698
rect 46992 28693 47002 29663
rect 47016 28690 47026 29663
rect 47040 28717 47050 29663
rect 47064 28717 47074 29663
rect 47088 28717 47098 29663
rect 47112 28717 47122 29663
rect 47136 28717 47146 29663
rect 47160 28717 47170 29663
rect 47184 28717 47194 29663
rect 47208 28717 47218 29663
rect 47232 28717 47242 29663
rect 47256 28717 47266 29663
rect 47280 28717 47290 29663
rect 47016 28680 47314 28690
rect 46968 28663 47026 28666
rect 46943 28656 47026 28663
rect 46943 28653 46978 28656
rect 47016 28645 47026 28656
rect 47304 28645 47314 28680
rect 46992 28618 47002 28631
rect 46992 28608 47338 28618
rect 46943 28594 46978 28597
rect 46943 28587 47002 28594
rect 46968 28584 47002 28587
rect 46992 27565 47002 28584
rect 46943 27542 46978 27552
rect 47016 27562 47026 28583
rect 47040 27589 47050 28583
rect 47064 27589 47074 28583
rect 47088 27589 47098 28583
rect 47112 27589 47122 28583
rect 47136 27589 47146 28583
rect 47160 27589 47170 28583
rect 47184 27589 47194 28583
rect 47208 27589 47218 28583
rect 47232 27589 47242 28583
rect 47256 27589 47266 28583
rect 47280 27589 47290 28583
rect 47304 27589 47314 28583
rect 47328 27589 47338 28608
rect 47016 27552 47362 27562
rect 46968 27538 46978 27542
rect 47352 27541 47362 27552
rect 46968 27528 47026 27538
rect 47016 27517 47026 27528
rect 47064 27514 47074 27527
rect 47064 27504 47386 27514
rect 46968 27486 47074 27490
rect 46943 27480 47074 27486
rect 46943 27476 46978 27480
rect 46992 26461 47002 27455
rect 47016 26461 47026 27455
rect 47040 26461 47050 27455
rect 47064 26461 47074 27480
rect 47088 26461 47098 27479
rect 47112 26461 47122 27479
rect 47136 26461 47146 27479
rect 47160 26461 47170 27479
rect 47184 26458 47194 27479
rect 47208 26485 47218 27479
rect 47232 26485 47242 27479
rect 47256 26485 47266 27479
rect 47280 26485 47290 27479
rect 47304 26485 47314 27479
rect 47328 26485 47338 27479
rect 47352 26485 47362 27479
rect 47376 26794 47386 27504
rect 50256 26821 50266 30743
rect 47376 26784 50279 26794
rect 47184 26448 47386 26458
rect 46943 26434 46978 26441
rect 46943 26431 47194 26434
rect 46968 26424 47194 26431
rect 47184 26413 47194 26424
rect 47376 26413 47386 26448
rect 47040 26386 47050 26399
rect 47040 26376 47410 26386
rect 46943 26365 46978 26375
rect 46968 26362 46978 26365
rect 46968 26352 47050 26362
rect 46992 25357 47002 26327
rect 47016 25357 47026 26327
rect 47040 25357 47050 26352
rect 47064 25357 47074 26351
rect 47088 25357 47098 26351
rect 47112 25354 47122 26351
rect 47136 25381 47146 26351
rect 47160 25381 47170 26351
rect 47184 25381 47194 26351
rect 47208 25381 47218 26351
rect 47232 25381 47242 26351
rect 47256 25381 47266 26351
rect 47280 25381 47290 26351
rect 47304 25381 47314 26351
rect 47328 25381 47338 26351
rect 47352 25381 47362 26351
rect 47376 25381 47386 26351
rect 47400 25381 47410 26376
rect 47112 25344 47434 25354
rect 46943 25320 47122 25330
rect 47112 25285 47122 25320
rect 47136 25285 47146 25319
rect 47160 25285 47170 25319
rect 47184 25285 47194 25319
rect 47208 25282 47218 25319
rect 47424 25309 47434 25344
rect 47208 25272 47458 25282
rect 46943 25258 46978 25264
rect 46943 25254 47218 25258
rect 46968 25248 47218 25254
rect 46992 24253 47002 25223
rect 47016 24253 47026 25223
rect 47040 24253 47050 25223
rect 47064 24253 47074 25223
rect 47088 24253 47098 25223
rect 47112 24253 47122 25223
rect 47136 24253 47146 25223
rect 47160 24250 47170 25223
rect 47184 24277 47194 25223
rect 47208 24277 47218 25248
rect 47232 24277 47242 25247
rect 47256 24277 47266 25247
rect 47280 24277 47290 25247
rect 47304 24277 47314 25247
rect 47328 24277 47338 25247
rect 47352 24277 47362 25247
rect 47376 24277 47386 25247
rect 47400 24277 47410 25247
rect 47424 24277 47434 25247
rect 47448 24277 47458 25272
rect 47160 24240 47482 24250
rect 46968 24219 47170 24226
rect 46943 24216 47170 24219
rect 46943 24209 46978 24216
rect 47160 24181 47170 24216
rect 47184 24181 47194 24215
rect 47208 24181 47218 24215
rect 47232 24181 47242 24215
rect 47256 24178 47266 24215
rect 47472 24205 47482 24240
rect 47256 24168 47506 24178
rect 46968 24153 47266 24154
rect 46943 24144 47266 24153
rect 46943 24143 46978 24144
rect 46992 23125 47002 24119
rect 47016 23125 47026 24119
rect 47040 23125 47050 24119
rect 47064 23125 47074 24119
rect 47088 23122 47098 24119
rect 47112 23149 47122 24119
rect 47136 23149 47146 24119
rect 47160 23149 47170 24119
rect 47184 23149 47194 24119
rect 47208 23149 47218 24119
rect 47232 23149 47242 24119
rect 47256 23149 47266 24144
rect 47280 23149 47290 24143
rect 47304 23149 47314 24143
rect 47328 23149 47338 24143
rect 47352 23149 47362 24143
rect 47376 23149 47386 24143
rect 47400 23149 47410 24143
rect 47424 23149 47434 24143
rect 47448 23149 47458 24143
rect 47472 23149 47482 24143
rect 47496 23149 47506 24168
rect 47088 23112 47530 23122
rect 46943 23098 46978 23108
rect 47520 23101 47530 23112
rect 46968 23088 47098 23098
rect 47088 23077 47098 23088
rect 47280 23074 47290 23087
rect 47280 23064 47554 23074
rect 46968 23042 47290 23050
rect 46943 23040 47290 23042
rect 46943 23032 46978 23040
rect 46992 22021 47002 23015
rect 47016 22021 47026 23015
rect 47040 22021 47050 23015
rect 47064 22021 47074 23015
rect 47088 22021 47098 23015
rect 47112 22021 47122 23015
rect 47136 22021 47146 23015
rect 47160 22021 47170 23015
rect 47184 22021 47194 23015
rect 47208 22021 47218 23015
rect 47232 22021 47242 23015
rect 47256 22021 47266 23015
rect 47280 22021 47290 23040
rect 47304 22021 47314 23039
rect 47328 22021 47338 23039
rect 47352 22021 47362 23039
rect 47376 22021 47386 23039
rect 47400 22021 47410 23039
rect 47424 22021 47434 23039
rect 47448 22021 47458 23039
rect 47472 22021 47482 23039
rect 47496 22021 47506 23039
rect 47520 22021 47530 23039
rect 47544 22021 47554 23064
rect 46943 21994 46978 21997
rect 46943 21987 47578 21994
rect 46968 21984 47578 21987
rect 47568 21973 47578 21984
rect 47136 21946 47146 21959
rect 47136 21936 47602 21946
rect 46943 21922 46978 21931
rect 46943 21921 47146 21922
rect 46968 21912 47146 21921
rect 46992 20917 47002 21887
rect 47016 20917 47026 21887
rect 47040 20917 47050 21887
rect 47064 20917 47074 21887
rect 47088 20917 47098 21887
rect 47112 20917 47122 21887
rect 47136 20917 47146 21912
rect 47160 20917 47170 21911
rect 47184 20917 47194 21911
rect 47208 20917 47218 21911
rect 47232 20917 47242 21911
rect 47256 20917 47266 21911
rect 47280 20917 47290 21911
rect 47304 20917 47314 21911
rect 47328 20917 47338 21911
rect 47352 20917 47362 21911
rect 47376 20917 47386 21911
rect 47400 20917 47410 21911
rect 47424 20917 47434 21911
rect 47448 20917 47458 21911
rect 47472 20917 47482 21911
rect 47496 20917 47506 21911
rect 47520 20917 47530 21911
rect 47544 20917 47554 21911
rect 47568 20917 47578 21911
rect 47592 20917 47602 21936
rect 46968 20886 47626 20890
rect 46943 20880 47626 20886
rect 46943 20876 46978 20880
rect 47616 20869 47626 20880
rect 47352 20842 47362 20855
rect 47352 20832 47650 20842
rect 46943 20818 46978 20820
rect 46943 20810 47362 20818
rect 46968 20808 47362 20810
rect 46992 19789 47002 20783
rect 47016 19789 47026 20783
rect 47040 19789 47050 20783
rect 47064 19789 47074 20783
rect 47088 19789 47098 20783
rect 47112 19789 47122 20783
rect 47136 19789 47146 20783
rect 47160 19789 47170 20783
rect 47184 19786 47194 20783
rect 47208 19813 47218 20783
rect 47232 19813 47242 20783
rect 47256 19813 47266 20783
rect 47280 19813 47290 20783
rect 47304 19813 47314 20783
rect 47328 19813 47338 20783
rect 47352 19813 47362 20808
rect 47376 19813 47386 20807
rect 47400 19813 47410 20807
rect 47424 19813 47434 20807
rect 47448 19813 47458 20807
rect 47472 19813 47482 20807
rect 47496 19813 47506 20807
rect 47520 19813 47530 20807
rect 47544 19813 47554 20807
rect 47568 19813 47578 20807
rect 47592 19813 47602 20807
rect 47616 19813 47626 20807
rect 47640 19813 47650 20832
rect 47184 19776 47674 19786
rect 46943 19765 46978 19775
rect 47664 19765 47674 19776
rect 46968 19762 46978 19765
rect 46968 19752 47183 19762
rect 47173 19728 47698 19738
rect 46968 19709 47170 19714
rect 46943 19704 47170 19709
rect 46943 19699 46978 19704
rect 21397 19632 21490 19642
rect 46992 19621 47002 19679
rect 47016 19621 47026 19679
rect 47040 19621 47050 19679
rect 47064 19621 47074 19679
rect 47088 19621 47098 19679
rect 47112 19621 47122 19679
rect 47136 19621 47146 19679
rect 47160 19621 47170 19704
rect 47184 19621 47194 19703
rect 20280 19608 21479 19618
rect 47208 19618 47218 19703
rect 47232 19645 47242 19703
rect 47256 19645 47266 19703
rect 47280 19645 47290 19703
rect 47304 19645 47314 19703
rect 47328 19645 47338 19703
rect 47352 19645 47362 19703
rect 47376 19645 47386 19703
rect 47400 19645 47410 19703
rect 47424 19645 47434 19703
rect 47448 19645 47458 19703
rect 47472 19645 47482 19703
rect 47496 19645 47506 19703
rect 47520 19645 47530 19703
rect 47544 19645 47554 19703
rect 47568 19645 47578 19703
rect 47592 19645 47602 19703
rect 47616 19645 47626 19703
rect 47640 19645 47650 19703
rect 47664 19642 47674 19703
rect 47688 19666 47698 19728
rect 47688 19656 48479 19666
rect 47664 19632 48791 19642
rect 47208 19608 48815 19618
rect 20256 19584 21503 19594
rect 21596 19584 21762 19594
rect 21752 19573 21762 19584
rect 20317 19560 21727 19570
rect 21133 19536 21582 19546
rect 21664 19536 21786 19546
rect 21776 19525 21786 19536
rect 21229 19512 21655 19522
rect 21120 19488 21582 19498
rect 21120 19069 21130 19488
rect 22008 19498 22018 19607
rect 21596 19488 22018 19498
rect 21397 19464 21594 19474
rect 21445 19440 21466 19450
rect 21456 19114 21466 19440
rect 21480 19141 21490 19439
rect 21504 19141 21514 19439
rect 21584 19141 21594 19464
rect 21608 19138 21618 19463
rect 21632 19165 21642 19463
rect 21656 19165 21666 19463
rect 21680 19165 21690 19463
rect 21704 19165 21714 19463
rect 21728 19165 21738 19463
rect 21752 19165 21762 19463
rect 21776 19162 21786 19463
rect 22008 19189 22018 19488
rect 21776 19152 22223 19162
rect 21608 19128 22247 19138
rect 23448 19138 23458 19607
rect 23448 19128 24119 19138
rect 24240 19138 24250 19607
rect 24792 19162 24802 19607
rect 25008 19186 25018 19607
rect 25008 19176 25031 19186
rect 25752 19186 25762 19607
rect 25752 19176 25847 19186
rect 25920 19186 25930 19607
rect 26304 19210 26314 19607
rect 26496 19234 26506 19607
rect 26496 19224 26687 19234
rect 26712 19234 26722 19607
rect 27456 19258 27466 19607
rect 27456 19248 27503 19258
rect 26712 19224 27551 19234
rect 27624 19234 27634 19607
rect 46128 19594 46138 19607
rect 30792 19584 46138 19594
rect 27624 19224 28607 19234
rect 30792 19213 30802 19584
rect 46320 19594 46330 19607
rect 46368 19594 46378 19607
rect 46416 19594 46426 19607
rect 46165 19584 46330 19594
rect 46344 19584 46378 19594
rect 46392 19584 46426 19594
rect 46488 19594 46498 19607
rect 46488 19584 47218 19594
rect 43104 19560 45167 19570
rect 26304 19200 29207 19210
rect 25920 19176 31319 19186
rect 24792 19152 32242 19162
rect 24240 19128 32207 19138
rect 32232 19138 32242 19152
rect 32232 19128 32975 19138
rect 21456 19104 21607 19114
rect 21765 19104 25823 19114
rect 25861 19104 33335 19114
rect 21549 19080 24095 19090
rect 24133 19080 31295 19090
rect 31333 19080 34991 19090
rect 21480 19066 21490 19079
rect 21480 19056 21535 19066
rect 21693 19056 28583 19066
rect 28621 19056 35026 19066
rect 20256 19032 22168 19042
rect 20256 18805 20266 19032
rect 22261 19032 26663 19042
rect 26701 19032 34967 19042
rect 35016 19042 35026 19056
rect 35016 19032 35807 19042
rect 37032 19042 37042 19559
rect 37224 19066 37234 19559
rect 37224 19056 37415 19066
rect 37464 19066 37474 19559
rect 37464 19056 38039 19066
rect 37032 19032 38266 19042
rect 21645 19008 27479 19018
rect 27517 19008 38231 19018
rect 38256 19018 38266 19032
rect 38256 19008 39082 19018
rect 21504 18994 21514 19007
rect 21504 18984 21679 18994
rect 21717 18984 29183 18994
rect 29221 18984 35783 18994
rect 35821 18984 39047 18994
rect 39072 18994 39082 19008
rect 39072 18984 40655 18994
rect 20280 18960 22144 18970
rect 20280 18778 20290 18960
rect 22237 18960 27527 18970
rect 27565 18960 38015 18970
rect 38053 18960 41471 18970
rect 21573 18936 25018 18946
rect 20207 18768 20290 18778
rect 20256 14722 20266 18743
rect 20207 14712 20266 14722
rect 21120 10717 21130 18935
rect 21537 18922 21547 18935
rect 25008 18925 25018 18936
rect 25045 18936 33322 18946
rect 33312 18925 33322 18936
rect 33349 18936 34954 18946
rect 34944 18925 34954 18936
rect 35005 18936 37402 18946
rect 34968 18925 34978 18935
rect 37392 18925 37402 18936
rect 37429 18936 42082 18946
rect 42072 18925 42082 18936
rect 43104 18925 43114 19560
rect 45205 19560 46271 19570
rect 46344 19570 46354 19584
rect 46296 19560 46354 19570
rect 43926 19536 45911 19546
rect 43926 18925 43936 19536
rect 46296 19546 46306 19560
rect 45949 19536 46306 19546
rect 43950 19512 45191 19522
rect 43950 18925 43960 19512
rect 45558 19512 46151 19522
rect 45558 18925 45568 19512
rect 45582 19488 45935 19498
rect 45582 18925 45592 19488
rect 46392 18925 46402 19584
rect 47208 19573 47218 19584
rect 47653 19584 48839 19594
rect 47616 19570 47626 19583
rect 47616 19560 48863 19570
rect 46824 19546 46834 19559
rect 46824 19536 48455 19546
rect 48493 19536 48887 19546
rect 47605 19512 48911 19522
rect 46992 18946 47002 19511
rect 47016 18970 47026 19511
rect 47040 18994 47050 19511
rect 47064 19018 47074 19511
rect 47088 19042 47098 19511
rect 47112 19066 47122 19511
rect 47136 19090 47146 19511
rect 47160 19114 47170 19511
rect 47184 19138 47194 19511
rect 47208 19165 47218 19511
rect 47232 19162 47242 19511
rect 47256 19186 47266 19511
rect 47280 19210 47290 19511
rect 47304 19234 47314 19511
rect 47328 19258 47338 19511
rect 47352 19282 47362 19511
rect 47376 19306 47386 19511
rect 47400 19330 47410 19511
rect 47424 19354 47434 19511
rect 47448 19378 47458 19511
rect 47472 19402 47482 19511
rect 47496 19426 47506 19511
rect 47520 19450 47530 19511
rect 47544 19474 47554 19511
rect 47568 19498 47578 19511
rect 47568 19488 48935 19498
rect 47544 19464 48959 19474
rect 47520 19440 48983 19450
rect 47496 19416 49007 19426
rect 47472 19392 49031 19402
rect 47448 19368 49055 19378
rect 47424 19344 49079 19354
rect 47400 19320 49103 19330
rect 47376 19296 49127 19306
rect 47352 19272 49151 19282
rect 47328 19248 49175 19258
rect 47304 19224 49199 19234
rect 47280 19200 49223 19210
rect 47256 19176 49247 19186
rect 47232 19152 49271 19162
rect 47184 19128 49295 19138
rect 47160 19104 49319 19114
rect 47136 19080 49343 19090
rect 50256 19090 50266 26759
rect 49381 19080 50266 19090
rect 47112 19056 49415 19066
rect 47088 19032 49463 19042
rect 47064 19008 50159 19018
rect 47040 18984 50207 18994
rect 47016 18960 50231 18970
rect 46992 18936 50266 18946
rect 21537 18912 21706 18922
rect 21597 18888 21641 18898
rect 21609 18749 21619 18863
rect 21631 18773 21641 18888
rect 21696 18805 21706 18912
rect 21631 18763 21743 18773
rect 48792 18752 48802 18906
rect 48816 18752 48826 18906
rect 21609 18739 21743 18749
rect 48840 18749 48850 18906
rect 48864 18776 48874 18906
rect 48888 18776 48898 18906
rect 48912 18776 48922 18906
rect 48936 18776 48946 18906
rect 48960 18776 48970 18906
rect 48984 18797 48994 18906
rect 49008 18824 49018 18906
rect 49032 18824 49042 18906
rect 49056 18869 49066 18906
rect 49416 18872 49426 18906
rect 49056 18859 49391 18869
rect 49464 18850 49474 18906
rect 50160 18853 50170 18911
rect 50208 18877 50218 18911
rect 50232 18877 50242 18911
rect 49056 18835 49079 18845
rect 49056 18824 49066 18835
rect 49381 18835 49450 18845
rect 50256 18850 50266 18936
rect 50197 18840 50266 18850
rect 49440 18826 49450 18835
rect 49093 18811 49391 18821
rect 49440 18816 50307 18826
rect 48984 18787 49402 18797
rect 48997 18763 49055 18773
rect 49392 18773 49402 18787
rect 49368 18763 49402 18773
rect 49368 18752 49378 18763
rect 49416 18752 49426 18810
rect 50136 18802 50146 18816
rect 50136 18792 50255 18802
rect 49464 18752 49474 18786
rect 50197 18768 50307 18778
rect 48840 18739 49055 18749
rect 50256 18730 50266 18743
rect 48781 18715 48839 18725
rect 49516 18725 50266 18730
rect 48853 18720 50266 18725
rect 48853 18715 49526 18720
rect 21648 14316 21658 18714
rect 21672 14343 21682 18714
rect 21696 14343 21706 18714
rect 21720 14343 21730 18714
rect 48781 18691 49367 18701
rect 48781 18667 49079 18677
rect 49272 18653 49282 18666
rect 49416 18656 49426 18690
rect 49464 18656 49474 18690
rect 50160 18661 50170 18695
rect 50208 18661 50218 18695
rect 50232 18661 50242 18695
rect 48781 18643 49282 18653
rect 48781 18619 48983 18629
rect 49516 18629 50307 18634
rect 49069 18624 50307 18629
rect 49069 18619 49526 18624
rect 48792 15133 48802 18594
rect 48816 15133 48826 18594
rect 48840 15133 48850 18594
rect 48864 15133 48874 18594
rect 48888 15133 48898 18594
rect 48912 15133 48922 18594
rect 48936 15133 48946 18594
rect 48960 15133 48970 18594
rect 49008 15106 49018 18618
rect 48781 15096 49018 15106
rect 21648 14306 21743 14316
rect 21709 14282 21743 14292
rect 21672 14266 21682 14281
rect 21672 14256 21706 14266
rect 20207 10680 21682 10690
rect 21120 10429 21130 10655
rect 21672 10429 21682 10680
rect 21696 10429 21706 14256
rect 21720 10435 21730 14257
rect 48792 12183 48802 15071
rect 48816 12183 48826 15071
rect 48840 14794 48850 15071
rect 48864 14821 48874 15071
rect 48888 14821 48898 15071
rect 48912 14821 48922 15071
rect 48936 14821 48946 15071
rect 48960 14821 48970 15071
rect 49032 14821 49042 18618
rect 49104 14821 49114 18594
rect 49128 14821 49138 18594
rect 49152 14821 49162 18594
rect 49176 14821 49186 18594
rect 49200 14821 49210 18594
rect 49224 14821 49234 18594
rect 49248 14821 49258 18594
rect 49296 14821 49306 18594
rect 49320 14821 49330 18594
rect 49344 14821 49354 18594
rect 49416 14821 49426 18594
rect 49464 14821 49474 18594
rect 50160 14821 50170 18599
rect 50208 14821 50218 18599
rect 50232 14821 50242 18599
rect 48840 14784 50307 14794
rect 50256 14773 50266 14784
rect 48864 12183 48874 14759
rect 48888 12183 48898 14759
rect 48912 12156 48922 14759
rect 48936 12159 48946 14759
rect 48960 12159 48970 14759
rect 48781 12146 48922 12156
rect 49032 12157 49042 14759
rect 49104 12132 49114 14759
rect 48781 12122 49114 12132
rect 48781 12098 48959 12108
rect 48792 10546 48802 12073
rect 48816 10573 48826 12073
rect 48864 10573 48874 12073
rect 48888 10573 48898 12073
rect 48936 10573 48946 12073
rect 49032 10573 49042 12095
rect 49128 10573 49138 14759
rect 49152 10573 49162 14759
rect 49176 10573 49186 14759
rect 49200 10573 49210 14759
rect 49224 10573 49234 14759
rect 49248 10573 49258 14759
rect 49296 10573 49306 14759
rect 49320 10573 49330 14759
rect 49344 10573 49354 14759
rect 49416 10573 49426 14759
rect 49464 10573 49474 14759
rect 50160 14746 50170 14759
rect 50160 14736 50307 14746
rect 50208 10690 50218 14711
rect 50232 14602 50242 14711
rect 50256 14629 50266 14711
rect 50232 14592 50307 14602
rect 50256 10738 50266 14567
rect 50256 10728 50307 10738
rect 50256 10717 50266 10728
rect 50208 10680 50307 10690
rect 50256 10573 50266 10655
rect 48792 10536 50307 10546
rect 21720 10425 21743 10435
rect 48816 10414 48826 10511
rect 48864 10414 48874 10511
rect 48888 10414 48898 10511
rect 48936 10414 48946 10511
rect 49032 10414 49042 10511
rect 49128 10414 49138 10511
rect 49152 10414 49162 10511
rect 49176 10414 49186 10511
rect 21072 10392 21743 10402
rect 21072 9759 21082 10392
rect 21685 10368 21730 10378
rect 49200 10387 49210 10511
rect 48781 10377 49210 10387
rect 21120 9826 21130 10367
rect 21696 10210 21706 10343
rect 21720 10234 21730 10368
rect 48781 10353 49175 10363
rect 48781 10329 49127 10339
rect 48781 10305 49031 10315
rect 22200 10234 22210 10247
rect 26208 10234 26218 10247
rect 21720 10224 22210 10234
rect 24744 10224 26218 10234
rect 21696 10200 21730 10210
rect 21720 10186 21730 10200
rect 21744 10200 22127 10210
rect 21744 10186 21754 10200
rect 21720 10176 21754 10186
rect 24744 9949 24754 10224
rect 26208 10042 26218 10224
rect 28285 10224 29591 10234
rect 31813 10224 39239 10234
rect 39277 10224 44783 10234
rect 48888 10234 48898 10280
rect 44821 10224 48898 10234
rect 28128 10200 48863 10210
rect 28128 10069 28138 10200
rect 48936 10189 48946 10280
rect 38869 10176 39263 10186
rect 42253 10176 44807 10186
rect 45925 10176 48815 10186
rect 28272 10069 28282 10175
rect 29592 10162 29602 10175
rect 49152 10162 49162 10328
rect 29592 10152 49162 10162
rect 49224 10141 49234 10511
rect 49248 10141 49258 10511
rect 49296 10141 49306 10511
rect 49320 10141 49330 10511
rect 31656 10128 48935 10138
rect 31656 10069 31666 10128
rect 49344 10114 49354 10511
rect 39253 10104 49354 10114
rect 31800 10069 31810 10103
rect 38856 10069 38866 10103
rect 44797 10080 49223 10090
rect 49320 10042 49330 10079
rect 26208 10032 49330 10042
rect 28128 9949 28138 10007
rect 28272 9949 28282 10007
rect 31656 9949 31666 10007
rect 31800 9949 31810 10007
rect 49416 9997 49426 10511
rect 49464 9970 49474 10511
rect 38712 9960 49474 9970
rect 38712 9949 38722 9960
rect 49296 9922 49306 9935
rect 24600 9912 49306 9922
rect 21120 9816 21178 9826
rect 21120 9759 21130 9816
rect 21168 9759 21178 9816
rect 24600 9759 24610 9912
rect 49416 9901 49426 9935
rect 45960 9888 46031 9898
rect 24744 9759 24754 9887
rect 28128 9853 28138 9887
rect 28272 9853 28282 9887
rect 31656 9853 31666 9887
rect 31800 9853 31810 9887
rect 38712 9853 38722 9887
rect 38856 9853 38866 9887
rect 42240 9853 42250 9887
rect 45960 9874 45970 9888
rect 45781 9864 45970 9874
rect 50256 9874 50266 10511
rect 45997 9864 50266 9874
rect 42397 9840 46018 9850
rect 24792 9816 45983 9826
rect 24792 9759 24802 9816
rect 28128 9759 28138 9791
rect 28272 9759 28282 9791
rect 28320 9759 28330 9816
rect 31656 9759 31666 9791
rect 31800 9759 31810 9791
rect 31848 9759 31858 9816
rect 38712 9759 38722 9791
rect 38856 9759 38866 9791
rect 38904 9759 38914 9816
rect 42240 9759 42250 9791
rect 42384 9759 42394 9791
rect 42432 9759 42442 9816
rect 45768 9759 45778 9791
rect 45912 9759 45922 9791
rect 45960 9759 45970 9816
rect 46008 9826 46018 9840
rect 46045 9840 49415 9850
rect 46008 9816 49247 9826
<< m2contact >>
rect 24551 39743 24565 39757
rect 28079 39743 28093 39757
rect 24623 39719 24637 39733
rect 31631 39743 31645 39757
rect 31775 39743 31789 39757
rect 38687 39743 38701 39757
rect 38831 39743 38845 39757
rect 42215 39743 42229 39757
rect 42359 39743 42373 39757
rect 45743 39743 45757 39757
rect 45887 39743 45901 39757
rect 45695 39719 45709 39733
rect 21503 39695 21517 39709
rect 24551 39695 24565 39709
rect 28079 39695 28093 39709
rect 31631 39695 31645 39709
rect 46991 39719 47005 39733
rect 46823 39695 46837 39709
rect 21455 39671 21469 39685
rect 21479 39671 21493 39685
rect 24623 39671 24637 39685
rect 21503 39647 21517 39661
rect 21455 39623 21469 39637
rect 21479 39623 21493 39637
rect 31775 39671 31789 39685
rect 38687 39671 38701 39685
rect 47015 39671 47029 39685
rect 47063 39671 47077 39685
rect 38831 39647 38845 39661
rect 47087 39647 47101 39661
rect 42215 39623 42229 39637
rect 42359 39623 42373 39637
rect 45695 39623 45709 39637
rect 45887 39623 45901 39637
rect 47039 39599 47053 39613
rect 47111 39599 47125 39613
rect 28079 39575 28093 39589
rect 31775 39575 31789 39589
rect 42215 39575 42229 39589
rect 42359 39575 42373 39589
rect 45743 39575 45757 39589
rect 45767 39575 45781 39589
rect 47015 39575 47029 39589
rect 47135 39575 47149 39589
rect 47015 39551 47029 39565
rect 47111 39551 47125 39565
rect 47159 39551 47173 39565
rect 28079 39527 28093 39541
rect 31775 39527 31789 39541
rect 45743 39527 45757 39541
rect 46871 39527 46885 39541
rect 46991 39527 47005 39541
rect 47207 39527 47221 39541
rect 38855 39503 38869 39517
rect 46991 39503 47005 39517
rect 47015 39503 47029 39517
rect 47231 39503 47245 39517
rect 47015 39479 47029 39493
rect 47039 39479 47053 39493
rect 47255 39479 47269 39493
rect 27887 39455 27901 39469
rect 28079 39455 28093 39469
rect 31775 39455 31789 39469
rect 38663 39455 38677 39469
rect 39023 39455 39037 39469
rect 47183 39455 47197 39469
rect 47207 39455 47221 39469
rect 47279 39455 47293 39469
rect 21215 39239 21229 39253
rect 21431 39239 21445 39253
rect 21455 39239 21469 39253
rect 21479 39239 21493 39253
rect 21215 39191 21229 39205
rect 20279 38807 20293 38821
rect 21215 38807 21229 38821
rect 21431 39191 21445 39205
rect 22007 39191 22021 39205
rect 20279 38759 20293 38773
rect 21215 38759 21229 38773
rect 20279 34823 20293 34837
rect 20255 34751 20269 34765
rect 20255 34703 20269 34717
rect 20279 34703 20293 34717
rect 20255 30767 20269 30781
rect 20279 30767 20293 30781
rect 20303 30767 20317 30781
rect 21215 30767 21229 30781
rect 47039 39431 47053 39445
rect 47087 39431 47101 39445
rect 47303 39431 47317 39445
rect 47111 39407 47125 39421
rect 47159 39407 47173 39421
rect 47255 39383 47269 39397
rect 47327 39383 47341 39397
rect 26855 39359 26869 39373
rect 36143 39359 36157 39373
rect 36863 39359 36877 39373
rect 47159 39359 47173 39373
rect 47207 39359 47221 39373
rect 47351 39359 47365 39373
rect 47255 39335 47269 39349
rect 47279 39335 47293 39349
rect 47375 39335 47389 39349
rect 26855 39311 26869 39325
rect 27887 39311 27901 39325
rect 28079 39311 28093 39325
rect 31775 39311 31789 39325
rect 47087 39311 47101 39325
rect 47135 39311 47149 39325
rect 47399 39311 47413 39325
rect 47279 39287 47293 39301
rect 47303 39287 47317 39301
rect 47423 39287 47437 39301
rect 26663 39263 26677 39277
rect 26855 39263 26869 39277
rect 27887 39263 27901 39277
rect 28079 39263 28093 39277
rect 31775 39263 31789 39277
rect 35879 39263 35893 39277
rect 38927 39263 38941 39277
rect 42359 39263 42373 39277
rect 45743 39263 45757 39277
rect 45767 39263 45781 39277
rect 47351 39263 47365 39277
rect 47375 39263 47389 39277
rect 47447 39263 47461 39277
rect 47135 39239 47149 39253
rect 47303 39239 47317 39253
rect 26663 39215 26677 39229
rect 26855 39215 26869 39229
rect 27887 39215 27901 39229
rect 28079 39215 28093 39229
rect 31775 39215 31789 39229
rect 42215 39191 42229 39205
rect 46823 39167 46837 39181
rect 46871 39191 46885 39205
rect 21455 39143 21469 39157
rect 21479 39143 21493 39157
rect 22127 39143 22141 39157
rect 25463 39143 25477 39157
rect 25703 39143 25717 39157
rect 26663 39143 26677 39157
rect 26855 39143 26869 39157
rect 27887 39143 27901 39157
rect 46823 39143 46837 39157
rect 46991 39143 47005 39157
rect 47015 39143 47029 39157
rect 47039 39143 47053 39157
rect 47063 39143 47077 39157
rect 47087 39143 47101 39157
rect 47111 39143 47125 39157
rect 47135 39143 47149 39157
rect 47159 39143 47173 39157
rect 47183 39143 47197 39157
rect 47207 39143 47221 39157
rect 47231 39143 47245 39157
rect 47255 39143 47269 39157
rect 47279 39143 47293 39157
rect 47303 39143 47317 39157
rect 47327 39143 47341 39157
rect 20303 30719 20317 30733
rect 21215 30719 21229 30733
rect 20255 30671 20269 30685
rect 20279 30671 20293 30685
rect 20279 26807 20293 26821
rect 20279 26759 20293 26773
rect 20279 22847 20293 22861
rect 20303 22847 20317 22861
rect 20279 22799 20293 22813
rect 20303 22799 20317 22813
rect 20303 19631 20317 19645
rect 21431 19655 21445 19669
rect 21119 19631 21133 19645
rect 21215 19631 21229 19645
rect 21383 19631 21397 19645
rect 47399 39191 47413 39205
rect 47423 39191 47437 39205
rect 47447 39191 47461 39205
rect 46991 36455 47005 36469
rect 47015 36455 47029 36469
rect 47039 36455 47053 36469
rect 47063 36455 47077 36469
rect 47087 36455 47101 36469
rect 47111 36455 47125 36469
rect 47135 36455 47149 36469
rect 47159 36455 47173 36469
rect 47183 36455 47197 36469
rect 47207 36455 47221 36469
rect 47231 36455 47245 36469
rect 47255 36455 47269 36469
rect 47279 36455 47293 36469
rect 47303 36455 47317 36469
rect 47327 36455 47341 36469
rect 47351 36455 47365 36469
rect 47375 36455 47389 36469
rect 47399 36455 47413 36469
rect 47423 36455 47437 36469
rect 47447 36455 47461 36469
rect 50255 38999 50269 39013
rect 50255 38951 50269 38965
rect 47447 36407 47461 36421
rect 46991 36335 47005 36349
rect 47015 36335 47029 36349
rect 47039 36335 47053 36349
rect 47063 36335 47077 36349
rect 47087 36335 47101 36349
rect 47111 36335 47125 36349
rect 47135 36335 47149 36349
rect 47159 36335 47173 36349
rect 47183 36335 47197 36349
rect 47207 36335 47221 36349
rect 47231 36335 47245 36349
rect 47255 36335 47269 36349
rect 47279 36335 47293 36349
rect 47303 36335 47317 36349
rect 47327 36335 47341 36349
rect 47351 36335 47365 36349
rect 47375 36335 47389 36349
rect 47399 36335 47413 36349
rect 47423 36335 47437 36349
rect 46991 35351 47005 35365
rect 47015 35351 47029 35365
rect 47039 35351 47053 35365
rect 47063 35351 47077 35365
rect 47087 35351 47101 35365
rect 47111 35351 47125 35365
rect 47135 35351 47149 35365
rect 47159 35351 47173 35365
rect 47183 35351 47197 35365
rect 47207 35351 47221 35365
rect 47231 35351 47245 35365
rect 47255 35351 47269 35365
rect 47279 35351 47293 35365
rect 47303 35351 47317 35365
rect 47327 35351 47341 35365
rect 47351 35351 47365 35365
rect 47375 35351 47389 35365
rect 47399 35351 47413 35365
rect 47399 35303 47413 35317
rect 46991 35231 47005 35245
rect 47015 35231 47029 35245
rect 47039 35231 47053 35245
rect 47063 35231 47077 35245
rect 47087 35231 47101 35245
rect 47111 35231 47125 35245
rect 47135 35231 47149 35245
rect 47159 35231 47173 35245
rect 47183 35231 47197 35245
rect 47207 35231 47221 35245
rect 47231 35231 47245 35245
rect 47255 35231 47269 35245
rect 47279 35231 47293 35245
rect 47303 35231 47317 35245
rect 47327 35231 47341 35245
rect 47351 35231 47365 35245
rect 47375 35231 47389 35245
rect 46991 34223 47005 34237
rect 47015 34223 47029 34237
rect 47039 34223 47053 34237
rect 47063 34223 47077 34237
rect 47087 34223 47101 34237
rect 47111 34223 47125 34237
rect 47135 34223 47149 34237
rect 47159 34223 47173 34237
rect 47183 34223 47197 34237
rect 47207 34223 47221 34237
rect 47231 34223 47245 34237
rect 47255 34223 47269 34237
rect 47279 34223 47293 34237
rect 47303 34223 47317 34237
rect 47327 34223 47341 34237
rect 47351 34223 47365 34237
rect 50255 38855 50269 38869
rect 50255 38807 50269 38821
rect 50231 34967 50245 34981
rect 50255 34967 50269 34981
rect 50231 34919 50245 34933
rect 50255 34919 50269 34933
rect 50183 34847 50197 34861
rect 50207 34847 50221 34861
rect 47351 34175 47365 34189
rect 46991 34103 47005 34117
rect 47015 34103 47029 34117
rect 47039 34103 47053 34117
rect 47063 34103 47077 34117
rect 47087 34103 47101 34117
rect 47111 34103 47125 34117
rect 47135 34103 47149 34117
rect 47159 34103 47173 34117
rect 47183 34103 47197 34117
rect 47207 34103 47221 34117
rect 47231 34103 47245 34117
rect 47255 34103 47269 34117
rect 47279 34103 47293 34117
rect 47303 34103 47317 34117
rect 47327 34103 47341 34117
rect 46991 33119 47005 33133
rect 47015 33119 47029 33133
rect 47039 33119 47053 33133
rect 47063 33119 47077 33133
rect 47087 33119 47101 33133
rect 47111 33119 47125 33133
rect 47135 33119 47149 33133
rect 47159 33119 47173 33133
rect 47183 33119 47197 33133
rect 47207 33119 47221 33133
rect 47231 33119 47245 33133
rect 47255 33119 47269 33133
rect 47279 33119 47293 33133
rect 47303 33119 47317 33133
rect 47303 33071 47317 33085
rect 46991 32999 47005 33013
rect 47015 32999 47029 33013
rect 47039 32999 47053 33013
rect 47063 32999 47077 33013
rect 47087 32999 47101 33013
rect 47111 32999 47125 33013
rect 47135 32999 47149 33013
rect 47159 32999 47173 33013
rect 47183 32999 47197 33013
rect 47207 32999 47221 33013
rect 47231 32999 47245 33013
rect 47255 32999 47269 33013
rect 47279 32999 47293 33013
rect 46991 32015 47005 32029
rect 47015 32015 47029 32029
rect 47039 32015 47053 32029
rect 47063 32015 47077 32029
rect 47087 32015 47101 32029
rect 47111 32015 47125 32029
rect 47135 32015 47149 32029
rect 47159 32015 47173 32029
rect 47183 32015 47197 32029
rect 47207 32015 47221 32029
rect 47231 32015 47245 32029
rect 47255 32015 47269 32029
rect 47279 32015 47293 32029
rect 50255 34823 50269 34837
rect 50183 34799 50197 34813
rect 50207 34799 50221 34813
rect 46991 31895 47005 31909
rect 47015 31895 47029 31909
rect 47039 31895 47053 31909
rect 47063 31895 47077 31909
rect 47087 31895 47101 31909
rect 47111 31895 47125 31909
rect 47135 31895 47149 31909
rect 47159 31895 47173 31909
rect 47183 31895 47197 31909
rect 47207 31895 47221 31909
rect 47231 31895 47245 31909
rect 47255 31895 47269 31909
rect 47279 31895 47293 31909
rect 50207 30959 50221 30973
rect 50255 34775 50269 34789
rect 46991 30887 47005 30901
rect 47015 30887 47029 30901
rect 47039 30887 47053 30901
rect 47063 30887 47077 30901
rect 47087 30887 47101 30901
rect 47111 30887 47125 30901
rect 47135 30887 47149 30901
rect 47159 30887 47173 30901
rect 47183 30887 47197 30901
rect 47207 30887 47221 30901
rect 47231 30887 47245 30901
rect 47255 30887 47269 30901
rect 47279 30887 47293 30901
rect 50255 30935 50269 30949
rect 50207 30911 50221 30925
rect 50255 30887 50269 30901
rect 46991 30791 47005 30805
rect 47015 30791 47029 30805
rect 47039 30791 47053 30805
rect 47063 30791 47077 30805
rect 47087 30791 47101 30805
rect 47111 30791 47125 30805
rect 47135 30791 47149 30805
rect 47159 30791 47173 30805
rect 47183 30791 47197 30805
rect 47207 30791 47221 30805
rect 47231 30791 47245 30805
rect 47255 30791 47269 30805
rect 47279 30791 47293 30805
rect 50231 30791 50245 30805
rect 50255 30791 50269 30805
rect 46991 29783 47005 29797
rect 47015 29783 47029 29797
rect 47039 29783 47053 29797
rect 47063 29783 47077 29797
rect 47087 29783 47101 29797
rect 47111 29783 47125 29797
rect 47135 29783 47149 29797
rect 47159 29783 47173 29797
rect 47183 29783 47197 29797
rect 47207 29783 47221 29797
rect 47231 29783 47245 29797
rect 47255 29783 47269 29797
rect 47279 29783 47293 29797
rect 50231 30743 50245 30757
rect 50255 30743 50269 30757
rect 46991 29663 47005 29677
rect 47015 29663 47029 29677
rect 47039 29663 47053 29677
rect 47063 29663 47077 29677
rect 47087 29663 47101 29677
rect 47111 29663 47125 29677
rect 47135 29663 47149 29677
rect 47159 29663 47173 29677
rect 47183 29663 47197 29677
rect 47207 29663 47221 29677
rect 47231 29663 47245 29677
rect 47255 29663 47269 29677
rect 47279 29663 47293 29677
rect 46991 28679 47005 28693
rect 47039 28703 47053 28717
rect 47063 28703 47077 28717
rect 47087 28703 47101 28717
rect 47111 28703 47125 28717
rect 47135 28703 47149 28717
rect 47159 28703 47173 28717
rect 47183 28703 47197 28717
rect 47207 28703 47221 28717
rect 47231 28703 47245 28717
rect 47255 28703 47269 28717
rect 47279 28703 47293 28717
rect 46991 28631 47005 28645
rect 47015 28631 47029 28645
rect 47303 28631 47317 28645
rect 47015 28583 47029 28597
rect 47039 28583 47053 28597
rect 47063 28583 47077 28597
rect 47087 28583 47101 28597
rect 47111 28583 47125 28597
rect 47135 28583 47149 28597
rect 47159 28583 47173 28597
rect 47183 28583 47197 28597
rect 47207 28583 47221 28597
rect 47231 28583 47245 28597
rect 47255 28583 47269 28597
rect 47279 28583 47293 28597
rect 47303 28583 47317 28597
rect 46991 27551 47005 27565
rect 47039 27575 47053 27589
rect 47063 27575 47077 27589
rect 47087 27575 47101 27589
rect 47111 27575 47125 27589
rect 47135 27575 47149 27589
rect 47159 27575 47173 27589
rect 47183 27575 47197 27589
rect 47207 27575 47221 27589
rect 47231 27575 47245 27589
rect 47255 27575 47269 27589
rect 47279 27575 47293 27589
rect 47303 27575 47317 27589
rect 47327 27575 47341 27589
rect 47063 27527 47077 27541
rect 47351 27527 47365 27541
rect 47015 27503 47029 27517
rect 46991 27455 47005 27469
rect 47015 27455 47029 27469
rect 47039 27455 47053 27469
rect 47087 27479 47101 27493
rect 47111 27479 47125 27493
rect 47135 27479 47149 27493
rect 47159 27479 47173 27493
rect 47183 27479 47197 27493
rect 47207 27479 47221 27493
rect 47231 27479 47245 27493
rect 47255 27479 47269 27493
rect 47279 27479 47293 27493
rect 47303 27479 47317 27493
rect 47327 27479 47341 27493
rect 47351 27479 47365 27493
rect 46991 26447 47005 26461
rect 47015 26447 47029 26461
rect 47039 26447 47053 26461
rect 47063 26447 47077 26461
rect 47087 26447 47101 26461
rect 47111 26447 47125 26461
rect 47135 26447 47149 26461
rect 47159 26447 47173 26461
rect 50255 26807 50269 26821
rect 50279 26783 50293 26797
rect 50255 26759 50269 26773
rect 47207 26471 47221 26485
rect 47231 26471 47245 26485
rect 47255 26471 47269 26485
rect 47279 26471 47293 26485
rect 47303 26471 47317 26485
rect 47327 26471 47341 26485
rect 47351 26471 47365 26485
rect 47039 26399 47053 26413
rect 47183 26399 47197 26413
rect 47375 26399 47389 26413
rect 46991 26327 47005 26341
rect 47015 26327 47029 26341
rect 47063 26351 47077 26365
rect 47087 26351 47101 26365
rect 47111 26351 47125 26365
rect 47135 26351 47149 26365
rect 47159 26351 47173 26365
rect 47183 26351 47197 26365
rect 47207 26351 47221 26365
rect 47231 26351 47245 26365
rect 47255 26351 47269 26365
rect 47279 26351 47293 26365
rect 47303 26351 47317 26365
rect 47327 26351 47341 26365
rect 47351 26351 47365 26365
rect 47375 26351 47389 26365
rect 46991 25343 47005 25357
rect 47015 25343 47029 25357
rect 47039 25343 47053 25357
rect 47063 25343 47077 25357
rect 47087 25343 47101 25357
rect 47135 25367 47149 25381
rect 47159 25367 47173 25381
rect 47183 25367 47197 25381
rect 47207 25367 47221 25381
rect 47231 25367 47245 25381
rect 47255 25367 47269 25381
rect 47279 25367 47293 25381
rect 47303 25367 47317 25381
rect 47327 25367 47341 25381
rect 47351 25367 47365 25381
rect 47375 25367 47389 25381
rect 47399 25367 47413 25381
rect 47135 25319 47149 25333
rect 47159 25319 47173 25333
rect 47183 25319 47197 25333
rect 47207 25319 47221 25333
rect 47111 25271 47125 25285
rect 47135 25271 47149 25285
rect 47159 25271 47173 25285
rect 47183 25271 47197 25285
rect 47423 25295 47437 25309
rect 46991 25223 47005 25237
rect 47015 25223 47029 25237
rect 47039 25223 47053 25237
rect 47063 25223 47077 25237
rect 47087 25223 47101 25237
rect 47111 25223 47125 25237
rect 47135 25223 47149 25237
rect 47159 25223 47173 25237
rect 47183 25223 47197 25237
rect 46991 24239 47005 24253
rect 47015 24239 47029 24253
rect 47039 24239 47053 24253
rect 47063 24239 47077 24253
rect 47087 24239 47101 24253
rect 47111 24239 47125 24253
rect 47135 24239 47149 24253
rect 47231 25247 47245 25261
rect 47255 25247 47269 25261
rect 47279 25247 47293 25261
rect 47303 25247 47317 25261
rect 47327 25247 47341 25261
rect 47351 25247 47365 25261
rect 47375 25247 47389 25261
rect 47399 25247 47413 25261
rect 47423 25247 47437 25261
rect 47183 24263 47197 24277
rect 47207 24263 47221 24277
rect 47231 24263 47245 24277
rect 47255 24263 47269 24277
rect 47279 24263 47293 24277
rect 47303 24263 47317 24277
rect 47327 24263 47341 24277
rect 47351 24263 47365 24277
rect 47375 24263 47389 24277
rect 47399 24263 47413 24277
rect 47423 24263 47437 24277
rect 47447 24263 47461 24277
rect 47183 24215 47197 24229
rect 47207 24215 47221 24229
rect 47231 24215 47245 24229
rect 47255 24215 47269 24229
rect 47159 24167 47173 24181
rect 47183 24167 47197 24181
rect 47207 24167 47221 24181
rect 47231 24167 47245 24181
rect 47471 24191 47485 24205
rect 46991 24119 47005 24133
rect 47015 24119 47029 24133
rect 47039 24119 47053 24133
rect 47063 24119 47077 24133
rect 47087 24119 47101 24133
rect 47111 24119 47125 24133
rect 47135 24119 47149 24133
rect 47159 24119 47173 24133
rect 47183 24119 47197 24133
rect 47207 24119 47221 24133
rect 47231 24119 47245 24133
rect 46991 23111 47005 23125
rect 47015 23111 47029 23125
rect 47039 23111 47053 23125
rect 47063 23111 47077 23125
rect 47279 24143 47293 24157
rect 47303 24143 47317 24157
rect 47327 24143 47341 24157
rect 47351 24143 47365 24157
rect 47375 24143 47389 24157
rect 47399 24143 47413 24157
rect 47423 24143 47437 24157
rect 47447 24143 47461 24157
rect 47471 24143 47485 24157
rect 47111 23135 47125 23149
rect 47135 23135 47149 23149
rect 47159 23135 47173 23149
rect 47183 23135 47197 23149
rect 47207 23135 47221 23149
rect 47231 23135 47245 23149
rect 47255 23135 47269 23149
rect 47279 23135 47293 23149
rect 47303 23135 47317 23149
rect 47327 23135 47341 23149
rect 47351 23135 47365 23149
rect 47375 23135 47389 23149
rect 47399 23135 47413 23149
rect 47423 23135 47437 23149
rect 47447 23135 47461 23149
rect 47471 23135 47485 23149
rect 47495 23135 47509 23149
rect 47279 23087 47293 23101
rect 47519 23087 47533 23101
rect 47087 23063 47101 23077
rect 46991 23015 47005 23029
rect 47015 23015 47029 23029
rect 47039 23015 47053 23029
rect 47063 23015 47077 23029
rect 47087 23015 47101 23029
rect 47111 23015 47125 23029
rect 47135 23015 47149 23029
rect 47159 23015 47173 23029
rect 47183 23015 47197 23029
rect 47207 23015 47221 23029
rect 47231 23015 47245 23029
rect 47255 23015 47269 23029
rect 47303 23039 47317 23053
rect 47327 23039 47341 23053
rect 47351 23039 47365 23053
rect 47375 23039 47389 23053
rect 47399 23039 47413 23053
rect 47423 23039 47437 23053
rect 47447 23039 47461 23053
rect 47471 23039 47485 23053
rect 47495 23039 47509 23053
rect 47519 23039 47533 23053
rect 46991 22007 47005 22021
rect 47015 22007 47029 22021
rect 47039 22007 47053 22021
rect 47063 22007 47077 22021
rect 47087 22007 47101 22021
rect 47111 22007 47125 22021
rect 47135 22007 47149 22021
rect 47159 22007 47173 22021
rect 47183 22007 47197 22021
rect 47207 22007 47221 22021
rect 47231 22007 47245 22021
rect 47255 22007 47269 22021
rect 47279 22007 47293 22021
rect 47303 22007 47317 22021
rect 47327 22007 47341 22021
rect 47351 22007 47365 22021
rect 47375 22007 47389 22021
rect 47399 22007 47413 22021
rect 47423 22007 47437 22021
rect 47447 22007 47461 22021
rect 47471 22007 47485 22021
rect 47495 22007 47509 22021
rect 47519 22007 47533 22021
rect 47543 22007 47557 22021
rect 47135 21959 47149 21973
rect 47567 21959 47581 21973
rect 46991 21887 47005 21901
rect 47015 21887 47029 21901
rect 47039 21887 47053 21901
rect 47063 21887 47077 21901
rect 47087 21887 47101 21901
rect 47111 21887 47125 21901
rect 47159 21911 47173 21925
rect 47183 21911 47197 21925
rect 47207 21911 47221 21925
rect 47231 21911 47245 21925
rect 47255 21911 47269 21925
rect 47279 21911 47293 21925
rect 47303 21911 47317 21925
rect 47327 21911 47341 21925
rect 47351 21911 47365 21925
rect 47375 21911 47389 21925
rect 47399 21911 47413 21925
rect 47423 21911 47437 21925
rect 47447 21911 47461 21925
rect 47471 21911 47485 21925
rect 47495 21911 47509 21925
rect 47519 21911 47533 21925
rect 47543 21911 47557 21925
rect 47567 21911 47581 21925
rect 46991 20903 47005 20917
rect 47015 20903 47029 20917
rect 47039 20903 47053 20917
rect 47063 20903 47077 20917
rect 47087 20903 47101 20917
rect 47111 20903 47125 20917
rect 47135 20903 47149 20917
rect 47159 20903 47173 20917
rect 47183 20903 47197 20917
rect 47207 20903 47221 20917
rect 47231 20903 47245 20917
rect 47255 20903 47269 20917
rect 47279 20903 47293 20917
rect 47303 20903 47317 20917
rect 47327 20903 47341 20917
rect 47351 20903 47365 20917
rect 47375 20903 47389 20917
rect 47399 20903 47413 20917
rect 47423 20903 47437 20917
rect 47447 20903 47461 20917
rect 47471 20903 47485 20917
rect 47495 20903 47509 20917
rect 47519 20903 47533 20917
rect 47543 20903 47557 20917
rect 47567 20903 47581 20917
rect 47591 20903 47605 20917
rect 47351 20855 47365 20869
rect 47615 20855 47629 20869
rect 46991 20783 47005 20797
rect 47015 20783 47029 20797
rect 47039 20783 47053 20797
rect 47063 20783 47077 20797
rect 47087 20783 47101 20797
rect 47111 20783 47125 20797
rect 47135 20783 47149 20797
rect 47159 20783 47173 20797
rect 47183 20783 47197 20797
rect 47207 20783 47221 20797
rect 47231 20783 47245 20797
rect 47255 20783 47269 20797
rect 47279 20783 47293 20797
rect 47303 20783 47317 20797
rect 47327 20783 47341 20797
rect 46991 19775 47005 19789
rect 47015 19775 47029 19789
rect 47039 19775 47053 19789
rect 47063 19775 47077 19789
rect 47087 19775 47101 19789
rect 47111 19775 47125 19789
rect 47135 19775 47149 19789
rect 47159 19775 47173 19789
rect 47375 20807 47389 20821
rect 47399 20807 47413 20821
rect 47423 20807 47437 20821
rect 47447 20807 47461 20821
rect 47471 20807 47485 20821
rect 47495 20807 47509 20821
rect 47519 20807 47533 20821
rect 47543 20807 47557 20821
rect 47567 20807 47581 20821
rect 47591 20807 47605 20821
rect 47615 20807 47629 20821
rect 47207 19799 47221 19813
rect 47231 19799 47245 19813
rect 47255 19799 47269 19813
rect 47279 19799 47293 19813
rect 47303 19799 47317 19813
rect 47327 19799 47341 19813
rect 47351 19799 47365 19813
rect 47375 19799 47389 19813
rect 47399 19799 47413 19813
rect 47423 19799 47437 19813
rect 47447 19799 47461 19813
rect 47471 19799 47485 19813
rect 47495 19799 47509 19813
rect 47519 19799 47533 19813
rect 47543 19799 47557 19813
rect 47567 19799 47581 19813
rect 47591 19799 47605 19813
rect 47615 19799 47629 19813
rect 47639 19799 47653 19813
rect 47183 19751 47197 19765
rect 47663 19751 47677 19765
rect 47159 19727 47173 19741
rect 46991 19679 47005 19693
rect 47015 19679 47029 19693
rect 47039 19679 47053 19693
rect 47063 19679 47077 19693
rect 47087 19679 47101 19693
rect 47111 19679 47125 19693
rect 47135 19679 47149 19693
rect 47183 19703 47197 19717
rect 47207 19703 47221 19717
rect 47231 19703 47245 19717
rect 47255 19703 47269 19717
rect 47279 19703 47293 19717
rect 47303 19703 47317 19717
rect 47327 19703 47341 19717
rect 47351 19703 47365 19717
rect 47375 19703 47389 19717
rect 47399 19703 47413 19717
rect 47423 19703 47437 19717
rect 47447 19703 47461 19717
rect 47471 19703 47485 19717
rect 47495 19703 47509 19717
rect 47519 19703 47533 19717
rect 47543 19703 47557 19717
rect 47567 19703 47581 19717
rect 47591 19703 47605 19717
rect 47615 19703 47629 19717
rect 47639 19703 47653 19717
rect 47663 19703 47677 19717
rect 21479 19607 21493 19621
rect 22007 19607 22021 19621
rect 23447 19607 23461 19621
rect 24239 19607 24253 19621
rect 24791 19607 24805 19621
rect 25007 19607 25021 19621
rect 25751 19607 25765 19621
rect 25919 19607 25933 19621
rect 26303 19607 26317 19621
rect 26495 19607 26509 19621
rect 26711 19607 26725 19621
rect 27455 19607 27469 19621
rect 27623 19607 27637 19621
rect 46127 19607 46141 19621
rect 46319 19607 46333 19621
rect 46367 19607 46381 19621
rect 46415 19607 46429 19621
rect 46487 19607 46501 19621
rect 46991 19607 47005 19621
rect 47015 19607 47029 19621
rect 47039 19607 47053 19621
rect 47063 19607 47077 19621
rect 47087 19607 47101 19621
rect 47111 19607 47125 19621
rect 47135 19607 47149 19621
rect 47159 19607 47173 19621
rect 47183 19607 47197 19621
rect 47231 19631 47245 19645
rect 47255 19631 47269 19645
rect 47279 19631 47293 19645
rect 47303 19631 47317 19645
rect 47327 19631 47341 19645
rect 47351 19631 47365 19645
rect 47375 19631 47389 19645
rect 47399 19631 47413 19645
rect 47423 19631 47437 19645
rect 47447 19631 47461 19645
rect 47471 19631 47485 19645
rect 47495 19631 47509 19645
rect 47519 19631 47533 19645
rect 47543 19631 47557 19645
rect 47567 19631 47581 19645
rect 47591 19631 47605 19645
rect 47615 19631 47629 19645
rect 47639 19631 47653 19645
rect 48479 19655 48493 19669
rect 48791 19631 48805 19645
rect 48815 19607 48829 19621
rect 21503 19583 21517 19597
rect 21582 19582 21596 19596
rect 20303 19559 20317 19573
rect 21727 19559 21741 19573
rect 21751 19559 21765 19573
rect 21119 19535 21133 19549
rect 21582 19535 21596 19549
rect 21650 19535 21664 19549
rect 21215 19511 21229 19525
rect 21655 19511 21669 19525
rect 21775 19511 21789 19525
rect 21582 19487 21596 19501
rect 21383 19463 21397 19477
rect 21431 19439 21445 19453
rect 21479 19439 21493 19453
rect 21503 19439 21517 19453
rect 21604 19463 21618 19477
rect 21628 19463 21642 19477
rect 21655 19463 21669 19477
rect 21679 19463 21693 19477
rect 21703 19463 21717 19477
rect 21727 19463 21741 19477
rect 21751 19463 21765 19477
rect 21775 19463 21789 19477
rect 21479 19127 21493 19141
rect 21503 19127 21517 19141
rect 21583 19127 21597 19141
rect 21631 19151 21645 19165
rect 21655 19151 21669 19165
rect 21679 19151 21693 19165
rect 21703 19151 21717 19165
rect 21727 19151 21741 19165
rect 21751 19151 21765 19165
rect 22007 19175 22021 19189
rect 22223 19151 22237 19165
rect 22247 19127 22261 19141
rect 24119 19127 24133 19141
rect 25031 19175 25045 19189
rect 25847 19175 25861 19189
rect 26687 19223 26701 19237
rect 27503 19247 27517 19261
rect 27551 19223 27565 19237
rect 28607 19223 28621 19237
rect 46151 19583 46165 19597
rect 37031 19559 37045 19573
rect 37223 19559 37237 19573
rect 37463 19559 37477 19573
rect 29207 19199 29221 19213
rect 30791 19199 30805 19213
rect 31319 19175 31333 19189
rect 32207 19127 32221 19141
rect 32975 19127 32989 19141
rect 21607 19103 21621 19117
rect 21751 19103 21765 19117
rect 25823 19103 25837 19117
rect 25847 19103 25861 19117
rect 33335 19103 33349 19117
rect 21479 19079 21493 19093
rect 21535 19079 21549 19093
rect 24095 19079 24109 19093
rect 24119 19079 24133 19093
rect 31295 19079 31309 19093
rect 31319 19079 31333 19093
rect 34991 19079 35005 19093
rect 21119 19055 21133 19069
rect 21535 19055 21549 19069
rect 21679 19055 21693 19069
rect 28583 19055 28597 19069
rect 28607 19055 28621 19069
rect 22168 19031 22182 19045
rect 22247 19031 22261 19045
rect 26663 19031 26677 19045
rect 26687 19031 26701 19045
rect 34967 19031 34981 19045
rect 35807 19031 35821 19045
rect 37415 19055 37429 19069
rect 38039 19055 38053 19069
rect 21503 19007 21517 19021
rect 21631 19007 21645 19021
rect 27479 19007 27493 19021
rect 27503 19007 27517 19021
rect 38231 19007 38245 19021
rect 21679 18983 21693 18997
rect 21703 18983 21717 18997
rect 29183 18983 29197 18997
rect 29207 18983 29221 18997
rect 35783 18983 35797 18997
rect 35807 18983 35821 18997
rect 39047 18983 39061 18997
rect 40655 18983 40669 18997
rect 20255 18791 20269 18805
rect 22144 18959 22158 18973
rect 22223 18959 22237 18973
rect 27527 18959 27541 18973
rect 27551 18959 27565 18973
rect 38015 18959 38029 18973
rect 38039 18959 38053 18973
rect 41471 18959 41485 18973
rect 21119 18935 21133 18949
rect 21535 18935 21549 18949
rect 21559 18935 21573 18949
rect 20255 18743 20269 18757
rect 25031 18935 25045 18949
rect 33335 18935 33349 18949
rect 34967 18935 34981 18949
rect 34991 18935 35005 18949
rect 37415 18935 37429 18949
rect 45167 19559 45181 19573
rect 45191 19559 45205 19573
rect 46271 19559 46285 19573
rect 45911 19535 45925 19549
rect 45935 19535 45949 19549
rect 45191 19511 45205 19525
rect 46151 19511 46165 19525
rect 45935 19487 45949 19501
rect 47615 19583 47629 19597
rect 47639 19583 47653 19597
rect 48839 19583 48853 19597
rect 46823 19559 46837 19573
rect 47207 19559 47221 19573
rect 48863 19559 48877 19573
rect 48455 19535 48469 19549
rect 48479 19535 48493 19549
rect 48887 19535 48901 19549
rect 46991 19511 47005 19525
rect 47015 19511 47029 19525
rect 47039 19511 47053 19525
rect 47063 19511 47077 19525
rect 47087 19511 47101 19525
rect 47111 19511 47125 19525
rect 47135 19511 47149 19525
rect 47159 19511 47173 19525
rect 47183 19511 47197 19525
rect 47207 19511 47221 19525
rect 47231 19511 47245 19525
rect 47255 19511 47269 19525
rect 47279 19511 47293 19525
rect 47303 19511 47317 19525
rect 47327 19511 47341 19525
rect 47351 19511 47365 19525
rect 47375 19511 47389 19525
rect 47399 19511 47413 19525
rect 47423 19511 47437 19525
rect 47447 19511 47461 19525
rect 47471 19511 47485 19525
rect 47495 19511 47509 19525
rect 47519 19511 47533 19525
rect 47543 19511 47557 19525
rect 47567 19511 47581 19525
rect 47591 19511 47605 19525
rect 48911 19511 48925 19525
rect 47207 19151 47221 19165
rect 48935 19487 48949 19501
rect 48959 19463 48973 19477
rect 48983 19439 48997 19453
rect 49007 19415 49021 19429
rect 49031 19391 49045 19405
rect 49055 19367 49069 19381
rect 49079 19343 49093 19357
rect 49103 19319 49117 19333
rect 49127 19295 49141 19309
rect 49151 19271 49165 19285
rect 49175 19247 49189 19261
rect 49199 19223 49213 19237
rect 49223 19199 49237 19213
rect 49247 19175 49261 19189
rect 49271 19151 49285 19165
rect 49295 19127 49309 19141
rect 49319 19103 49333 19117
rect 49343 19079 49357 19093
rect 49367 19079 49381 19093
rect 49415 19055 49429 19069
rect 49463 19031 49477 19045
rect 50159 19007 50173 19021
rect 50207 18983 50221 18997
rect 50231 18959 50245 18973
rect 21583 18887 21597 18901
rect 21607 18863 21621 18877
rect 25007 18911 25021 18925
rect 33311 18911 33325 18925
rect 34943 18911 34957 18925
rect 34967 18911 34981 18925
rect 37391 18911 37405 18925
rect 42071 18911 42085 18925
rect 43103 18911 43117 18925
rect 43924 18911 43938 18925
rect 43948 18911 43962 18925
rect 45556 18911 45570 18925
rect 45580 18911 45594 18925
rect 46391 18911 46405 18925
rect 48791 18906 48805 18920
rect 48815 18906 48829 18920
rect 48839 18906 48853 18920
rect 48863 18906 48877 18920
rect 48887 18906 48901 18920
rect 48911 18906 48925 18920
rect 48935 18906 48949 18920
rect 48959 18906 48973 18920
rect 48983 18906 48997 18920
rect 49007 18906 49021 18920
rect 49031 18906 49045 18920
rect 49055 18906 49069 18920
rect 49415 18906 49429 18920
rect 49463 18906 49477 18920
rect 50159 18911 50173 18925
rect 50207 18911 50221 18925
rect 50231 18911 50245 18925
rect 21695 18791 21709 18805
rect 21743 18762 21757 18776
rect 21743 18738 21757 18752
rect 48791 18738 48805 18752
rect 48815 18738 48829 18752
rect 49391 18858 49405 18872
rect 49415 18858 49429 18872
rect 50207 18863 50221 18877
rect 50231 18863 50245 18877
rect 49079 18834 49093 18848
rect 49367 18834 49381 18848
rect 49463 18836 49477 18850
rect 50159 18839 50173 18853
rect 50183 18839 50197 18853
rect 49007 18810 49021 18824
rect 49031 18810 49045 18824
rect 49055 18810 49069 18824
rect 49079 18810 49093 18824
rect 49391 18810 49405 18824
rect 49415 18810 49429 18824
rect 48863 18762 48877 18776
rect 48887 18762 48901 18776
rect 48911 18762 48925 18776
rect 48935 18762 48949 18776
rect 48959 18762 48973 18776
rect 48983 18762 48997 18776
rect 49055 18762 49069 18776
rect 49463 18786 49477 18800
rect 50255 18791 50269 18805
rect 50183 18767 50197 18781
rect 49055 18738 49069 18752
rect 49367 18738 49381 18752
rect 49415 18738 49429 18752
rect 49463 18738 49477 18752
rect 50255 18743 50269 18757
rect 21647 18714 21661 18728
rect 21671 18714 21685 18728
rect 21695 18714 21709 18728
rect 21719 18714 21733 18728
rect 48767 18714 48781 18728
rect 48839 18714 48853 18728
rect 48767 18690 48781 18704
rect 49367 18690 49381 18704
rect 49415 18690 49429 18704
rect 49463 18690 49477 18704
rect 50159 18695 50173 18709
rect 50207 18695 50221 18709
rect 50231 18695 50245 18709
rect 48767 18666 48781 18680
rect 49079 18666 49093 18680
rect 49271 18666 49285 18680
rect 48767 18642 48781 18656
rect 49415 18642 49429 18656
rect 49463 18642 49477 18656
rect 50159 18647 50173 18661
rect 50207 18647 50221 18661
rect 50231 18647 50245 18661
rect 48767 18618 48781 18632
rect 48983 18618 48997 18632
rect 49007 18618 49021 18632
rect 49031 18618 49045 18632
rect 49055 18618 49069 18632
rect 48791 18594 48805 18608
rect 48815 18594 48829 18608
rect 48839 18594 48853 18608
rect 48863 18594 48877 18608
rect 48887 18594 48901 18608
rect 48911 18594 48925 18608
rect 48935 18594 48949 18608
rect 48959 18594 48973 18608
rect 48791 15119 48805 15133
rect 48815 15119 48829 15133
rect 48839 15119 48853 15133
rect 48863 15119 48877 15133
rect 48887 15119 48901 15133
rect 48911 15119 48925 15133
rect 48935 15119 48949 15133
rect 48959 15119 48973 15133
rect 48767 15095 48781 15109
rect 48791 15071 48805 15085
rect 48815 15071 48829 15085
rect 48839 15071 48853 15085
rect 48863 15071 48877 15085
rect 48887 15071 48901 15085
rect 48911 15071 48925 15085
rect 48935 15071 48949 15085
rect 48959 15071 48973 15085
rect 21671 14329 21685 14343
rect 21695 14329 21709 14343
rect 21719 14329 21733 14343
rect 21743 14305 21757 14319
rect 21671 14281 21685 14295
rect 21695 14281 21709 14295
rect 21743 14281 21757 14295
rect 21719 14257 21733 14271
rect 21119 10703 21133 10717
rect 21119 10655 21133 10669
rect 49103 18594 49117 18608
rect 49127 18594 49141 18608
rect 49151 18594 49165 18608
rect 49175 18594 49189 18608
rect 49199 18594 49213 18608
rect 49223 18594 49237 18608
rect 49247 18594 49261 18608
rect 49295 18594 49309 18608
rect 49319 18594 49333 18608
rect 49343 18594 49357 18608
rect 49415 18594 49429 18608
rect 49463 18594 49477 18608
rect 50159 18599 50173 18613
rect 50207 18599 50221 18613
rect 50231 18599 50245 18613
rect 48863 14807 48877 14821
rect 48887 14807 48901 14821
rect 48911 14807 48925 14821
rect 48935 14807 48949 14821
rect 48959 14807 48973 14821
rect 49031 14807 49045 14821
rect 49103 14807 49117 14821
rect 49127 14807 49141 14821
rect 49151 14807 49165 14821
rect 49175 14807 49189 14821
rect 49199 14807 49213 14821
rect 49223 14807 49237 14821
rect 49247 14807 49261 14821
rect 49295 14807 49309 14821
rect 49319 14807 49333 14821
rect 49343 14807 49357 14821
rect 49415 14807 49429 14821
rect 49463 14807 49477 14821
rect 50159 14807 50173 14821
rect 50207 14807 50221 14821
rect 50231 14807 50245 14821
rect 48863 14759 48877 14773
rect 48887 14759 48901 14773
rect 48911 14759 48925 14773
rect 48935 14759 48949 14773
rect 48959 14759 48973 14773
rect 49031 14759 49045 14773
rect 49103 14759 49117 14773
rect 49127 14759 49141 14773
rect 49151 14759 49165 14773
rect 49175 14759 49189 14773
rect 49199 14759 49213 14773
rect 49223 14759 49237 14773
rect 49247 14759 49261 14773
rect 49295 14759 49309 14773
rect 49319 14759 49333 14773
rect 49343 14759 49357 14773
rect 49415 14759 49429 14773
rect 49463 14759 49477 14773
rect 50159 14759 50173 14773
rect 50255 14759 50269 14773
rect 48791 12169 48805 12183
rect 48815 12169 48829 12183
rect 48863 12169 48877 12183
rect 48887 12169 48901 12183
rect 48767 12145 48781 12159
rect 48935 12145 48949 12159
rect 48959 12145 48973 12159
rect 49031 12143 49045 12157
rect 48767 12121 48781 12135
rect 48767 12097 48781 12111
rect 48959 12097 48973 12111
rect 49031 12095 49045 12109
rect 48791 12073 48805 12087
rect 48815 12073 48829 12087
rect 48863 12073 48877 12087
rect 48887 12073 48901 12087
rect 48935 12073 48949 12087
rect 50207 14711 50221 14725
rect 50231 14711 50245 14725
rect 50255 14711 50269 14725
rect 50255 14615 50269 14629
rect 50255 14567 50269 14581
rect 50255 10703 50269 10717
rect 50255 10655 50269 10669
rect 48815 10559 48829 10573
rect 48863 10559 48877 10573
rect 48887 10559 48901 10573
rect 48935 10559 48949 10573
rect 49031 10559 49045 10573
rect 49127 10559 49141 10573
rect 49151 10559 49165 10573
rect 49175 10559 49189 10573
rect 49199 10559 49213 10573
rect 49223 10559 49237 10573
rect 49247 10559 49261 10573
rect 49295 10559 49309 10573
rect 49319 10559 49333 10573
rect 49343 10559 49357 10573
rect 49415 10559 49429 10573
rect 49463 10559 49477 10573
rect 50255 10559 50269 10573
rect 48815 10511 48829 10525
rect 48863 10511 48877 10525
rect 48887 10511 48901 10525
rect 48935 10511 48949 10525
rect 49031 10511 49045 10525
rect 49127 10511 49141 10525
rect 49151 10511 49165 10525
rect 49175 10511 49189 10525
rect 49199 10511 49213 10525
rect 49223 10511 49237 10525
rect 49247 10511 49261 10525
rect 49295 10511 49309 10525
rect 49319 10511 49333 10525
rect 49343 10511 49357 10525
rect 49415 10511 49429 10525
rect 49463 10511 49477 10525
rect 50255 10511 50269 10525
rect 21119 10415 21133 10429
rect 21671 10415 21685 10429
rect 21695 10415 21709 10429
rect 21743 10424 21757 10438
rect 21743 10391 21757 10405
rect 48815 10400 48829 10414
rect 48863 10400 48877 10414
rect 48887 10400 48901 10414
rect 48935 10400 48949 10414
rect 49031 10400 49045 10414
rect 49127 10400 49141 10414
rect 49151 10400 49165 10414
rect 49175 10400 49189 10414
rect 21119 10367 21133 10381
rect 21671 10367 21685 10381
rect 48767 10376 48781 10390
rect 21695 10343 21709 10357
rect 48767 10352 48781 10366
rect 49175 10352 49189 10366
rect 48767 10328 48781 10342
rect 49127 10328 49141 10342
rect 49151 10328 49165 10342
rect 48767 10304 48781 10318
rect 49031 10304 49045 10318
rect 48887 10280 48901 10294
rect 48935 10280 48949 10294
rect 22199 10247 22213 10261
rect 26207 10247 26221 10261
rect 22127 10199 22141 10213
rect 28271 10223 28285 10237
rect 29591 10223 29605 10237
rect 31799 10223 31813 10237
rect 39239 10223 39253 10237
rect 39263 10223 39277 10237
rect 44783 10223 44797 10237
rect 44807 10223 44821 10237
rect 48863 10199 48877 10213
rect 28271 10175 28285 10189
rect 29591 10175 29605 10189
rect 38855 10175 38869 10189
rect 39263 10175 39277 10189
rect 42239 10175 42253 10189
rect 44807 10175 44821 10189
rect 45911 10175 45925 10189
rect 48815 10175 48829 10189
rect 48935 10175 48949 10189
rect 48935 10127 48949 10141
rect 49223 10127 49237 10141
rect 49247 10127 49261 10141
rect 49295 10127 49309 10141
rect 49319 10127 49333 10141
rect 31799 10103 31813 10117
rect 38855 10103 38869 10117
rect 39239 10103 39253 10117
rect 44783 10079 44797 10093
rect 49223 10079 49237 10093
rect 49319 10079 49333 10093
rect 28127 10055 28141 10069
rect 28271 10055 28285 10069
rect 31655 10055 31669 10069
rect 31799 10055 31813 10069
rect 38855 10055 38869 10069
rect 28127 10007 28141 10021
rect 28271 10007 28285 10021
rect 31655 10007 31669 10021
rect 31799 10007 31813 10021
rect 49415 9983 49429 9997
rect 24743 9935 24757 9949
rect 28127 9935 28141 9949
rect 28271 9935 28285 9949
rect 31655 9935 31669 9949
rect 31799 9935 31813 9949
rect 38711 9935 38725 9949
rect 49295 9935 49309 9949
rect 49415 9935 49429 9949
rect 24743 9887 24757 9901
rect 28127 9887 28141 9901
rect 28271 9887 28285 9901
rect 31655 9887 31669 9901
rect 31799 9887 31813 9901
rect 38711 9887 38725 9901
rect 38855 9887 38869 9901
rect 42239 9887 42253 9901
rect 45767 9863 45781 9877
rect 46031 9887 46045 9901
rect 49415 9887 49429 9901
rect 45983 9863 45997 9877
rect 28127 9839 28141 9853
rect 28271 9839 28285 9853
rect 31655 9839 31669 9853
rect 31799 9839 31813 9853
rect 38711 9839 38725 9853
rect 38855 9839 38869 9853
rect 42239 9839 42253 9853
rect 42383 9839 42397 9853
rect 28127 9791 28141 9805
rect 28271 9791 28285 9805
rect 31655 9791 31669 9805
rect 31799 9791 31813 9805
rect 38711 9791 38725 9805
rect 38855 9791 38869 9805
rect 42239 9791 42253 9805
rect 42383 9791 42397 9805
rect 45767 9791 45781 9805
rect 45911 9791 45925 9805
rect 45983 9815 45997 9829
rect 46031 9839 46045 9853
rect 49415 9839 49429 9853
rect 49247 9815 49261 9829
<< metal2 >>
rect 24552 39709 24564 39743
rect 21456 39637 21468 39671
rect 21480 39637 21492 39671
rect 21504 39661 21516 39695
rect 24624 39685 24636 39719
rect 28080 39709 28092 39743
rect 31632 39709 31644 39743
rect 31776 39685 31788 39743
rect 38688 39685 38700 39743
rect 38832 39661 38844 39743
rect 42216 39637 42228 39743
rect 42360 39637 42372 39743
rect 45696 39637 45708 39719
rect 45744 39589 45756 39743
rect 45888 39637 45900 39743
rect 28080 39541 28092 39575
rect 31776 39541 31788 39575
rect 26856 39325 26868 39359
rect 27888 39325 27900 39455
rect 28080 39325 28092 39455
rect 31776 39325 31788 39455
rect 21216 39205 21228 39239
rect 21432 39205 21444 39239
rect 21456 39157 21468 39239
rect 21480 39157 21492 39239
rect 26664 39229 26676 39263
rect 26856 39229 26868 39263
rect 27888 39229 27900 39263
rect 28080 39229 28092 39263
rect 31776 39229 31788 39263
rect 22008 39133 22020 39191
rect 22121 39143 22127 39157
rect 25457 39143 25463 39157
rect 25697 39143 25703 39157
rect 26657 39143 26663 39157
rect 26849 39143 26855 39157
rect 27883 39143 27887 39157
rect 35880 39156 35892 39263
rect 36144 39156 36156 39359
rect 36864 39156 36876 39359
rect 38664 39156 38676 39455
rect 38856 39156 38868 39503
rect 38928 39156 38940 39263
rect 39024 39156 39036 39455
rect 42216 39205 42228 39575
rect 42360 39277 42372 39575
rect 45744 39277 45756 39527
rect 45768 39277 45780 39575
rect 46824 39181 46836 39695
rect 46992 39541 47004 39719
rect 47016 39589 47028 39671
rect 46872 39205 46884 39527
rect 47016 39517 47028 39551
rect 46992 39157 47004 39503
rect 47040 39493 47052 39599
rect 47016 39157 47028 39479
rect 47040 39157 47052 39431
rect 47064 39157 47076 39671
rect 47088 39445 47100 39647
rect 47112 39565 47124 39599
rect 47088 39157 47100 39311
rect 47112 39157 47124 39407
rect 47136 39325 47148 39575
rect 47160 39421 47172 39551
rect 47208 39469 47220 39527
rect 47136 39157 47148 39239
rect 47160 39157 47172 39359
rect 47184 39157 47196 39455
rect 47208 39157 47220 39359
rect 47232 39157 47244 39503
rect 47256 39397 47268 39479
rect 47280 39349 47292 39455
rect 47256 39157 47268 39335
rect 47304 39301 47316 39431
rect 47280 39157 47292 39287
rect 47304 39157 47316 39239
rect 47328 39157 47340 39383
rect 47352 39277 47364 39359
rect 47376 39277 47388 39335
rect 47400 39205 47412 39311
rect 47424 39205 47436 39287
rect 47448 39205 47460 39263
rect 35874 39144 35892 39156
rect 36138 39144 36156 39156
rect 36858 39144 36876 39156
rect 38657 39144 38676 39156
rect 38849 39144 38868 39156
rect 38921 39144 38940 39156
rect 39017 39144 39036 39156
rect 22121 39133 22133 39143
rect 25457 39133 25469 39143
rect 25697 39133 25709 39143
rect 26657 39133 26669 39143
rect 26849 39133 26861 39143
rect 27883 39133 27895 39143
rect 35874 39133 35886 39144
rect 36138 39133 36150 39144
rect 36858 39133 36870 39144
rect 38657 39133 38669 39144
rect 38849 39133 38861 39144
rect 38921 39133 38933 39144
rect 39017 39133 39029 39144
rect 46824 39133 46836 39143
rect 50256 38965 50268 38999
rect 50256 38821 50268 38855
rect 20280 38773 20292 38807
rect 21216 38773 21228 38807
rect 46992 36349 47004 36455
rect 47016 36349 47028 36455
rect 47040 36349 47052 36455
rect 47064 36349 47076 36455
rect 47088 36349 47100 36455
rect 47112 36349 47124 36455
rect 47136 36349 47148 36455
rect 47160 36349 47172 36455
rect 47184 36349 47196 36455
rect 47208 36349 47220 36455
rect 47232 36349 47244 36455
rect 47256 36349 47268 36455
rect 47280 36349 47292 36455
rect 47304 36349 47316 36455
rect 47328 36349 47340 36455
rect 47352 36349 47364 36455
rect 47376 36349 47388 36455
rect 47400 36349 47412 36455
rect 47424 36349 47436 36455
rect 47448 36421 47460 36455
rect 46992 35245 47004 35351
rect 47016 35245 47028 35351
rect 47040 35245 47052 35351
rect 47064 35245 47076 35351
rect 47088 35245 47100 35351
rect 47112 35245 47124 35351
rect 47136 35245 47148 35351
rect 47160 35245 47172 35351
rect 47184 35245 47196 35351
rect 47208 35245 47220 35351
rect 47232 35245 47244 35351
rect 47256 35245 47268 35351
rect 47280 35245 47292 35351
rect 47304 35245 47316 35351
rect 47328 35245 47340 35351
rect 47352 35245 47364 35351
rect 47376 35245 47388 35351
rect 47400 35317 47412 35351
rect 50232 34933 50244 34967
rect 50256 34933 50268 34967
rect 20256 34717 20268 34751
rect 20280 34717 20292 34823
rect 50184 34813 50196 34847
rect 50208 34813 50220 34847
rect 50256 34789 50268 34823
rect 46992 34117 47004 34223
rect 47016 34117 47028 34223
rect 47040 34117 47052 34223
rect 47064 34117 47076 34223
rect 47088 34117 47100 34223
rect 47112 34117 47124 34223
rect 47136 34117 47148 34223
rect 47160 34117 47172 34223
rect 47184 34117 47196 34223
rect 47208 34117 47220 34223
rect 47232 34117 47244 34223
rect 47256 34117 47268 34223
rect 47280 34117 47292 34223
rect 47304 34117 47316 34223
rect 47328 34117 47340 34223
rect 47352 34189 47364 34223
rect 46992 33013 47004 33119
rect 47016 33013 47028 33119
rect 47040 33013 47052 33119
rect 47064 33013 47076 33119
rect 47088 33013 47100 33119
rect 47112 33013 47124 33119
rect 47136 33013 47148 33119
rect 47160 33013 47172 33119
rect 47184 33013 47196 33119
rect 47208 33013 47220 33119
rect 47232 33013 47244 33119
rect 47256 33013 47268 33119
rect 47280 33013 47292 33119
rect 47304 33085 47316 33119
rect 46992 31909 47004 32015
rect 47016 31909 47028 32015
rect 47040 31909 47052 32015
rect 47064 31909 47076 32015
rect 47088 31909 47100 32015
rect 47112 31909 47124 32015
rect 47136 31909 47148 32015
rect 47160 31909 47172 32015
rect 47184 31909 47196 32015
rect 47208 31909 47220 32015
rect 47232 31909 47244 32015
rect 47256 31909 47268 32015
rect 47280 31909 47292 32015
rect 50208 30925 50220 30959
rect 50256 30901 50268 30935
rect 46992 30805 47004 30887
rect 47016 30805 47028 30887
rect 47040 30805 47052 30887
rect 47064 30805 47076 30887
rect 47088 30805 47100 30887
rect 47112 30805 47124 30887
rect 47136 30805 47148 30887
rect 47160 30805 47172 30887
rect 47184 30805 47196 30887
rect 47208 30805 47220 30887
rect 47232 30805 47244 30887
rect 47256 30805 47268 30887
rect 47280 30805 47292 30887
rect 20256 30685 20268 30767
rect 20280 30685 20292 30767
rect 20304 30733 20316 30767
rect 21216 30733 21228 30767
rect 50232 30757 50244 30791
rect 50256 30757 50268 30791
rect 46992 29677 47004 29783
rect 47016 29677 47028 29783
rect 47040 29677 47052 29783
rect 47064 29677 47076 29783
rect 47088 29677 47100 29783
rect 47112 29677 47124 29783
rect 47136 29677 47148 29783
rect 47160 29677 47172 29783
rect 47184 29677 47196 29783
rect 47208 29677 47220 29783
rect 47232 29677 47244 29783
rect 47256 29677 47268 29783
rect 47280 29677 47292 29783
rect 46992 28645 47004 28679
rect 47016 28597 47028 28631
rect 47040 28597 47052 28703
rect 47064 28597 47076 28703
rect 47088 28597 47100 28703
rect 47112 28597 47124 28703
rect 47136 28597 47148 28703
rect 47160 28597 47172 28703
rect 47184 28597 47196 28703
rect 47208 28597 47220 28703
rect 47232 28597 47244 28703
rect 47256 28597 47268 28703
rect 47280 28597 47292 28703
rect 47304 28597 47316 28631
rect 46992 27469 47004 27551
rect 47016 27469 47028 27503
rect 47040 27469 47052 27575
rect 47064 27541 47076 27575
rect 47088 27493 47100 27575
rect 47112 27493 47124 27575
rect 47136 27493 47148 27575
rect 47160 27493 47172 27575
rect 47184 27493 47196 27575
rect 47208 27493 47220 27575
rect 47232 27493 47244 27575
rect 47256 27493 47268 27575
rect 47280 27493 47292 27575
rect 47304 27493 47316 27575
rect 47328 27493 47340 27575
rect 47352 27493 47364 27527
rect 20280 26773 20292 26807
rect 50256 26773 50268 26807
rect 50293 26784 50307 26796
rect 46992 26341 47004 26447
rect 47016 26341 47028 26447
rect 47040 26413 47052 26447
rect 47064 26365 47076 26447
rect 47088 26365 47100 26447
rect 47112 26365 47124 26447
rect 47136 26365 47148 26447
rect 47160 26365 47172 26447
rect 47184 26365 47196 26399
rect 47208 26365 47220 26471
rect 47232 26365 47244 26471
rect 47256 26365 47268 26471
rect 47280 26365 47292 26471
rect 47304 26365 47316 26471
rect 47328 26365 47340 26471
rect 47352 26365 47364 26471
rect 47376 26365 47388 26399
rect 46992 25237 47004 25343
rect 47016 25237 47028 25343
rect 47040 25237 47052 25343
rect 47064 25237 47076 25343
rect 47088 25237 47100 25343
rect 47136 25333 47148 25367
rect 47160 25333 47172 25367
rect 47184 25333 47196 25367
rect 47208 25333 47220 25367
rect 47112 25237 47124 25271
rect 47136 25237 47148 25271
rect 47160 25237 47172 25271
rect 47184 25237 47196 25271
rect 47232 25261 47244 25367
rect 47256 25261 47268 25367
rect 47280 25261 47292 25367
rect 47304 25261 47316 25367
rect 47328 25261 47340 25367
rect 47352 25261 47364 25367
rect 47376 25261 47388 25367
rect 47400 25261 47412 25367
rect 47424 25261 47436 25295
rect 46992 24133 47004 24239
rect 47016 24133 47028 24239
rect 47040 24133 47052 24239
rect 47064 24133 47076 24239
rect 47088 24133 47100 24239
rect 47112 24133 47124 24239
rect 47136 24133 47148 24239
rect 47184 24229 47196 24263
rect 47208 24229 47220 24263
rect 47232 24229 47244 24263
rect 47256 24229 47268 24263
rect 47160 24133 47172 24167
rect 47184 24133 47196 24167
rect 47208 24133 47220 24167
rect 47232 24133 47244 24167
rect 47280 24157 47292 24263
rect 47304 24157 47316 24263
rect 47328 24157 47340 24263
rect 47352 24157 47364 24263
rect 47376 24157 47388 24263
rect 47400 24157 47412 24263
rect 47424 24157 47436 24263
rect 47448 24157 47460 24263
rect 47472 24157 47484 24191
rect 46992 23029 47004 23111
rect 47016 23029 47028 23111
rect 47040 23029 47052 23111
rect 47064 23029 47076 23111
rect 47088 23029 47100 23063
rect 47112 23029 47124 23135
rect 47136 23029 47148 23135
rect 47160 23029 47172 23135
rect 47184 23029 47196 23135
rect 47208 23029 47220 23135
rect 47232 23029 47244 23135
rect 47256 23029 47268 23135
rect 47280 23101 47292 23135
rect 47304 23053 47316 23135
rect 47328 23053 47340 23135
rect 47352 23053 47364 23135
rect 47376 23053 47388 23135
rect 47400 23053 47412 23135
rect 47424 23053 47436 23135
rect 47448 23053 47460 23135
rect 47472 23053 47484 23135
rect 47496 23053 47508 23135
rect 47520 23053 47532 23087
rect 20280 22813 20292 22847
rect 20304 22813 20316 22847
rect 46992 21901 47004 22007
rect 47016 21901 47028 22007
rect 47040 21901 47052 22007
rect 47064 21901 47076 22007
rect 47088 21901 47100 22007
rect 47112 21901 47124 22007
rect 47136 21973 47148 22007
rect 47160 21925 47172 22007
rect 47184 21925 47196 22007
rect 47208 21925 47220 22007
rect 47232 21925 47244 22007
rect 47256 21925 47268 22007
rect 47280 21925 47292 22007
rect 47304 21925 47316 22007
rect 47328 21925 47340 22007
rect 47352 21925 47364 22007
rect 47376 21925 47388 22007
rect 47400 21925 47412 22007
rect 47424 21925 47436 22007
rect 47448 21925 47460 22007
rect 47472 21925 47484 22007
rect 47496 21925 47508 22007
rect 47520 21925 47532 22007
rect 47544 21925 47556 22007
rect 47568 21925 47580 21959
rect 46992 20797 47004 20903
rect 47016 20797 47028 20903
rect 47040 20797 47052 20903
rect 47064 20797 47076 20903
rect 47088 20797 47100 20903
rect 47112 20797 47124 20903
rect 47136 20797 47148 20903
rect 47160 20797 47172 20903
rect 47184 20797 47196 20903
rect 47208 20797 47220 20903
rect 47232 20797 47244 20903
rect 47256 20797 47268 20903
rect 47280 20797 47292 20903
rect 47304 20797 47316 20903
rect 47328 20797 47340 20903
rect 47352 20869 47364 20903
rect 47376 20821 47388 20903
rect 47400 20821 47412 20903
rect 47424 20821 47436 20903
rect 47448 20821 47460 20903
rect 47472 20821 47484 20903
rect 47496 20821 47508 20903
rect 47520 20821 47532 20903
rect 47544 20821 47556 20903
rect 47568 20821 47580 20903
rect 47592 20821 47604 20903
rect 47616 20821 47628 20855
rect 46992 19693 47004 19775
rect 47016 19693 47028 19775
rect 47040 19693 47052 19775
rect 47064 19693 47076 19775
rect 47088 19693 47100 19775
rect 47112 19693 47124 19775
rect 47136 19693 47148 19775
rect 47160 19741 47172 19775
rect 47184 19717 47196 19751
rect 47208 19717 47220 19799
rect 47232 19717 47244 19799
rect 47256 19717 47268 19799
rect 47280 19717 47292 19799
rect 47304 19717 47316 19799
rect 47328 19717 47340 19799
rect 47352 19717 47364 19799
rect 47376 19717 47388 19799
rect 47400 19717 47412 19799
rect 47424 19717 47436 19799
rect 47448 19717 47460 19799
rect 47472 19717 47484 19799
rect 47496 19717 47508 19799
rect 47520 19717 47532 19799
rect 47544 19717 47556 19799
rect 47568 19717 47580 19799
rect 47592 19717 47604 19799
rect 47616 19717 47628 19799
rect 47640 19717 47652 19799
rect 47664 19717 47676 19751
rect 20304 19573 20316 19631
rect 21120 19549 21132 19631
rect 21216 19525 21228 19631
rect 21384 19477 21396 19631
rect 21432 19453 21444 19655
rect 21480 19453 21492 19607
rect 21504 19453 21516 19583
rect 21480 19093 21492 19127
rect 21120 18949 21132 19055
rect 21504 19021 21516 19127
rect 21536 19093 21548 19643
rect 21536 18949 21548 19055
rect 21559 18949 21571 19643
rect 21582 19596 21594 19643
rect 21605 19630 21618 19643
rect 21583 19501 21595 19535
rect 21606 19477 21618 19630
rect 21628 19477 21640 19643
rect 21651 19549 21663 19643
rect 21674 19582 21686 19643
rect 21697 19620 21709 19643
rect 22008 19621 22020 19643
rect 21697 19608 21716 19620
rect 21674 19570 21692 19582
rect 21656 19477 21668 19511
rect 21680 19477 21692 19570
rect 21704 19477 21716 19608
rect 21728 19477 21740 19559
rect 21752 19477 21764 19559
rect 21776 19477 21788 19511
rect 21584 18901 21596 19127
rect 21608 18877 21620 19103
rect 21632 19021 21644 19151
rect 21656 18951 21668 19151
rect 21680 19069 21692 19151
rect 21704 18997 21716 19151
rect 21648 18935 21668 18951
rect 20256 18757 20268 18791
rect 21648 18728 21660 18935
rect 21680 18912 21692 18983
rect 21728 18947 21740 19151
rect 21752 19117 21764 19151
rect 21672 18900 21692 18912
rect 21720 18935 21740 18947
rect 21672 18728 21684 18900
rect 21696 18728 21708 18791
rect 21720 18728 21732 18935
rect 22008 18882 22020 19175
rect 22121 18882 22133 19643
rect 22145 18973 22157 19643
rect 22169 19045 22181 19643
rect 22145 18882 22157 18959
rect 22169 18882 22181 19031
rect 22193 18882 22205 19643
rect 23441 19621 23453 19643
rect 24233 19621 24245 19643
rect 24785 19621 24797 19643
rect 25001 19621 25013 19643
rect 25745 19621 25757 19643
rect 25913 19621 25925 19643
rect 26297 19621 26309 19643
rect 26489 19621 26501 19643
rect 26705 19621 26717 19643
rect 27449 19621 27461 19643
rect 27617 19621 27629 19643
rect 23441 19607 23447 19621
rect 24233 19607 24239 19621
rect 24785 19607 24791 19621
rect 25001 19607 25007 19621
rect 25745 19607 25751 19621
rect 25913 19607 25919 19621
rect 26297 19607 26303 19621
rect 26489 19607 26495 19621
rect 26705 19607 26711 19621
rect 27449 19607 27455 19621
rect 27617 19607 27623 19621
rect 37025 19620 37037 19643
rect 37217 19620 37229 19643
rect 37457 19620 37469 19643
rect 45161 19620 45173 19643
rect 45905 19620 45917 19643
rect 46121 19621 46133 19643
rect 37025 19608 37044 19620
rect 37217 19608 37236 19620
rect 37457 19608 37476 19620
rect 45161 19608 45180 19620
rect 45905 19608 45924 19620
rect 37032 19573 37044 19608
rect 37224 19573 37236 19608
rect 37464 19573 37476 19608
rect 45168 19573 45180 19608
rect 45192 19525 45204 19559
rect 45912 19549 45924 19608
rect 46121 19607 46127 19621
rect 46265 19620 46277 19643
rect 46313 19621 46325 19643
rect 46361 19621 46373 19643
rect 46409 19621 46421 19643
rect 46481 19621 46493 19643
rect 46265 19608 46284 19620
rect 45936 19501 45948 19535
rect 46152 19525 46164 19583
rect 46272 19573 46284 19608
rect 46313 19607 46319 19621
rect 46361 19607 46367 19621
rect 46409 19607 46415 19621
rect 46481 19607 46487 19621
rect 46824 19573 46836 19643
rect 46992 19525 47004 19607
rect 47016 19525 47028 19607
rect 47040 19525 47052 19607
rect 47064 19525 47076 19607
rect 47088 19525 47100 19607
rect 47112 19525 47124 19607
rect 47136 19525 47148 19607
rect 47160 19525 47172 19607
rect 47184 19525 47196 19607
rect 47208 19525 47220 19559
rect 47232 19525 47244 19631
rect 47256 19525 47268 19631
rect 47280 19525 47292 19631
rect 47304 19525 47316 19631
rect 47328 19525 47340 19631
rect 47352 19525 47364 19631
rect 47376 19525 47388 19631
rect 47400 19525 47412 19631
rect 47424 19525 47436 19631
rect 47448 19525 47460 19631
rect 47472 19525 47484 19631
rect 47496 19525 47508 19631
rect 47520 19525 47532 19631
rect 47544 19525 47556 19631
rect 47568 19525 47580 19631
rect 47592 19525 47604 19631
rect 47616 19597 47628 19631
rect 47640 19597 47652 19631
rect 48480 19549 48492 19655
rect 22224 18973 22236 19151
rect 22248 19045 22260 19127
rect 24120 19093 24132 19127
rect 24096 18924 24108 19079
rect 25032 18949 25044 19175
rect 25848 19117 25860 19175
rect 24096 18912 24113 18924
rect 24101 18882 24113 18912
rect 25001 18911 25007 18925
rect 25824 18924 25836 19103
rect 26688 19045 26700 19223
rect 26664 18924 26676 19031
rect 27504 19021 27516 19247
rect 25824 18912 25841 18924
rect 25001 18882 25013 18911
rect 25829 18882 25841 18912
rect 26657 18912 26676 18924
rect 27480 18924 27492 19007
rect 27552 18973 27564 19223
rect 28608 19069 28620 19223
rect 27528 18924 27540 18959
rect 27480 18912 27497 18924
rect 26657 18882 26669 18912
rect 27485 18882 27497 18912
rect 27521 18912 27540 18924
rect 28584 18924 28596 19055
rect 29208 18997 29220 19199
rect 29184 18924 29196 18983
rect 28584 18912 28601 18924
rect 27521 18882 27533 18912
rect 28589 18882 28601 18912
rect 29177 18912 29196 18924
rect 30792 18924 30804 19199
rect 31320 19093 31332 19175
rect 31296 18924 31308 19079
rect 32208 18924 32220 19127
rect 32976 18924 32988 19127
rect 33336 18949 33348 19103
rect 34968 18949 34980 19031
rect 34992 18949 35004 19079
rect 35808 18997 35820 19031
rect 30792 18912 30809 18924
rect 31296 18912 31313 18924
rect 32208 18912 32225 18924
rect 32976 18912 32993 18924
rect 29177 18882 29189 18912
rect 30797 18882 30809 18912
rect 31301 18882 31313 18912
rect 32213 18882 32225 18912
rect 32981 18882 32993 18912
rect 33325 18911 33329 18925
rect 33317 18882 33329 18911
rect 34937 18911 34943 18925
rect 34981 18911 34985 18925
rect 35784 18924 35796 18983
rect 37416 18949 37428 19055
rect 38040 18973 38052 19055
rect 35784 18912 35801 18924
rect 34937 18882 34949 18911
rect 34973 18882 34985 18911
rect 35789 18882 35801 18912
rect 37405 18911 37409 18925
rect 38016 18924 38028 18959
rect 38232 18924 38244 19007
rect 39048 18924 39060 18983
rect 40656 18924 40668 18983
rect 41472 18924 41484 18959
rect 38016 18912 38033 18924
rect 38232 18912 38249 18924
rect 39048 18912 39065 18924
rect 40656 18912 40673 18924
rect 41472 18912 41489 18924
rect 37397 18882 37409 18911
rect 38021 18882 38033 18912
rect 38237 18882 38249 18912
rect 39053 18882 39065 18912
rect 40661 18882 40673 18912
rect 41477 18882 41489 18912
rect 42085 18911 42089 18925
rect 43117 18911 43121 18925
rect 46405 18911 46409 18925
rect 47208 18924 47220 19151
rect 47208 18912 47225 18924
rect 42077 18882 42089 18911
rect 43109 18882 43121 18911
rect 43925 18882 43937 18911
rect 43949 18882 43961 18911
rect 45557 18882 45569 18911
rect 45581 18882 45593 18911
rect 46397 18882 46409 18911
rect 47213 18882 47225 18912
rect 48456 18882 48468 19535
rect 48792 18920 48804 19631
rect 48816 18920 48828 19607
rect 48840 18920 48852 19583
rect 48864 18920 48876 19559
rect 48888 18920 48900 19535
rect 48912 18920 48924 19511
rect 48936 18920 48948 19487
rect 48960 18920 48972 19463
rect 48984 18920 48996 19439
rect 49008 18920 49020 19415
rect 49032 18920 49044 19391
rect 49056 18920 49068 19367
rect 49080 18848 49092 19343
rect 21757 18763 21782 18775
rect 21757 18739 21782 18751
rect 48735 18715 48767 18727
rect 48735 18691 48767 18703
rect 48735 18667 48767 18679
rect 48735 18643 48767 18655
rect 48735 18619 48767 18631
rect 48792 18608 48804 18738
rect 48816 18608 48828 18738
rect 48840 18608 48852 18714
rect 48864 18608 48876 18762
rect 48888 18608 48900 18762
rect 48912 18608 48924 18762
rect 48936 18608 48948 18762
rect 48960 18608 48972 18762
rect 48984 18632 48996 18762
rect 49008 18632 49020 18810
rect 49032 18632 49044 18810
rect 49056 18776 49068 18810
rect 49056 18632 49068 18738
rect 49080 18680 49092 18810
rect 49104 18608 49116 19319
rect 49128 18608 49140 19295
rect 49152 18608 49164 19271
rect 49176 18608 49188 19247
rect 49200 18608 49212 19223
rect 49224 18608 49236 19199
rect 49248 18608 49260 19175
rect 49272 18680 49284 19151
rect 49296 18608 49308 19127
rect 49320 18608 49332 19103
rect 49344 18608 49356 19079
rect 49368 18848 49380 19079
rect 49416 18920 49428 19055
rect 49464 18920 49476 19031
rect 50160 18925 50172 19007
rect 50208 18925 50220 18983
rect 50232 18925 50244 18959
rect 49392 18824 49404 18858
rect 49416 18824 49428 18858
rect 49464 18800 49476 18836
rect 49368 18704 49380 18738
rect 49416 18704 49428 18738
rect 49464 18704 49476 18738
rect 50160 18709 50172 18839
rect 50184 18781 50196 18839
rect 50208 18709 50220 18863
rect 50232 18709 50244 18863
rect 50256 18757 50268 18791
rect 49416 18608 49428 18642
rect 49464 18608 49476 18642
rect 50160 18613 50172 18647
rect 50208 18613 50220 18647
rect 50232 18613 50244 18647
rect 48735 15109 48781 15110
rect 48735 15098 48767 15109
rect 48792 15085 48804 15119
rect 48816 15085 48828 15119
rect 48840 15085 48852 15119
rect 48864 15085 48876 15119
rect 48888 15085 48900 15119
rect 48912 15085 48924 15119
rect 48936 15085 48948 15119
rect 48960 15085 48972 15119
rect 48864 14773 48876 14807
rect 48888 14773 48900 14807
rect 48912 14773 48924 14807
rect 48936 14773 48948 14807
rect 48960 14773 48972 14807
rect 49032 14773 49044 14807
rect 49104 14773 49116 14807
rect 49128 14773 49140 14807
rect 49152 14773 49164 14807
rect 49176 14773 49188 14807
rect 49200 14773 49212 14807
rect 49224 14773 49236 14807
rect 49248 14773 49260 14807
rect 49296 14773 49308 14807
rect 49320 14773 49332 14807
rect 49344 14773 49356 14807
rect 49416 14773 49428 14807
rect 49464 14773 49476 14807
rect 50160 14773 50172 14807
rect 50208 14725 50220 14807
rect 50232 14725 50244 14807
rect 50256 14725 50268 14759
rect 50256 14581 50268 14615
rect 21672 14295 21684 14329
rect 21696 14295 21708 14329
rect 21720 14271 21732 14329
rect 21757 14306 21782 14318
rect 21757 14282 21782 14294
rect 48735 12146 48767 12158
rect 48735 12122 48767 12134
rect 48735 12098 48767 12110
rect 48792 12087 48804 12169
rect 48816 12087 48828 12169
rect 48864 12087 48876 12169
rect 48888 12087 48900 12169
rect 48936 12087 48948 12145
rect 48960 12111 48972 12145
rect 49032 12109 49044 12143
rect 21120 10669 21132 10703
rect 50256 10669 50268 10703
rect 48816 10525 48828 10559
rect 48864 10525 48876 10559
rect 48888 10525 48900 10559
rect 48936 10525 48948 10559
rect 49032 10525 49044 10559
rect 49128 10525 49140 10559
rect 49152 10525 49164 10559
rect 49176 10525 49188 10559
rect 49200 10525 49212 10559
rect 49224 10525 49236 10559
rect 49248 10525 49260 10559
rect 49296 10525 49308 10559
rect 49320 10525 49332 10559
rect 49344 10525 49356 10559
rect 49416 10525 49428 10559
rect 49464 10525 49476 10559
rect 50256 10525 50268 10559
rect 21757 10425 21782 10437
rect 21120 10381 21132 10415
rect 21672 10381 21684 10415
rect 21696 10357 21708 10415
rect 21743 10405 21782 10413
rect 21757 10401 21782 10405
rect 48735 10377 48767 10389
rect 48735 10353 48767 10365
rect 48735 10329 48767 10341
rect 48735 10305 48767 10317
rect 22121 10260 22133 10294
rect 22193 10261 22205 10294
rect 26213 10261 26225 10294
rect 22121 10248 22140 10260
rect 22128 10213 22140 10248
rect 22193 10247 22199 10261
rect 26221 10247 26225 10261
rect 29597 10260 29609 10294
rect 39245 10260 39257 10294
rect 44789 10260 44801 10294
rect 29592 10248 29609 10260
rect 39240 10248 39257 10260
rect 44784 10248 44801 10260
rect 29592 10237 29604 10248
rect 39240 10237 39252 10248
rect 44784 10237 44796 10248
rect 28272 10189 28284 10223
rect 29592 10189 29604 10223
rect 31800 10117 31812 10223
rect 38856 10117 38868 10175
rect 39240 10117 39252 10223
rect 39264 10189 39276 10223
rect 28128 10021 28140 10055
rect 28272 10021 28284 10055
rect 31656 10021 31668 10055
rect 31800 10021 31812 10055
rect 24744 9901 24756 9935
rect 28128 9901 28140 9935
rect 28272 9901 28284 9935
rect 31656 9901 31668 9935
rect 31800 9901 31812 9935
rect 38712 9901 38724 9935
rect 38856 9901 38868 10055
rect 42240 9901 42252 10175
rect 44784 10093 44796 10223
rect 44808 10189 44820 10223
rect 48816 10189 48828 10400
rect 48864 10213 48876 10400
rect 48888 10294 48900 10400
rect 48936 10294 48948 10400
rect 49032 10318 49044 10400
rect 49128 10342 49140 10400
rect 49152 10342 49164 10400
rect 49176 10366 49188 10400
rect 28128 9805 28140 9839
rect 28272 9805 28284 9839
rect 31656 9805 31668 9839
rect 31800 9805 31812 9839
rect 38712 9805 38724 9839
rect 38856 9805 38868 9839
rect 42240 9805 42252 9839
rect 42384 9805 42396 9839
rect 45768 9805 45780 9863
rect 45912 9805 45924 10175
rect 48936 10141 48948 10175
rect 49224 10093 49236 10127
rect 45984 9829 45996 9863
rect 46032 9853 46044 9887
rect 49248 9829 49260 10127
rect 49296 9949 49308 10127
rect 49320 10093 49332 10127
rect 49416 9949 49428 9983
rect 49416 9853 49428 9887
<< metal4 >>
rect 20373 44585 21933 46145
rect 23899 44585 25459 46145
rect 27425 44585 28985 46145
rect 30951 44585 32511 46145
rect 34477 44585 36037 46145
rect 38003 44585 39563 46145
rect 41529 44585 43089 46145
rect 45055 44585 46615 46145
rect 48581 44585 50141 46145
rect 13835 38133 15395 39693
rect 55119 38133 56679 39693
rect 13835 34091 15395 35651
rect 55119 34091 56679 35651
rect 13835 30049 15395 31609
rect 55119 30049 56679 31609
rect 13835 26007 15395 27567
rect 55119 26007 56679 27567
rect 13835 21965 15395 23525
rect 55119 21965 56679 23525
rect 13835 17923 15395 19483
rect 55119 17923 56679 19483
rect 13835 13881 15395 15441
rect 55119 13881 56679 15441
rect 13835 9839 15395 11399
rect 55119 9839 56679 11399
rect 20373 3387 21933 4947
rect 23899 3387 25459 4947
rect 27425 3387 28985 4947
rect 30951 3387 32511 4947
rect 34477 3387 36037 4947
rect 38003 3387 39563 4947
rect 41529 3387 43089 4947
rect 45055 3387 46615 4947
rect 48581 3387 50141 4947
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 13757 -1 0 46223
box 0 0 6450 6450
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 20293 1 0 39773
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 22013 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 22099 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 22185 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 22271 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 22357 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 22443 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 22529 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 22615 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 22701 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 22787 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 22873 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 22959 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 23045 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 23131 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 23217 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 23303 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 23389 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 23475 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 23561 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 23647 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 23733 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 23819 1 0 39773
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 25539 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 25625 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 25711 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 25797 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 25883 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 25969 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 26055 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 26141 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 26227 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 26313 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 26399 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 26485 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 26571 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 26657 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 26743 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 26829 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 26915 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 27001 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 27087 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 27173 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 27259 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 27345 1 0 39773
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 29065 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 29151 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 29237 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 29323 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 29409 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 29495 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 29581 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 29667 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 29753 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 29839 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 29925 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 30011 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 0 -1 30097 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 0 -1 30183 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 0 -1 30269 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 0 -1 30355 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 0 -1 30441 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 0 -1 30527 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 0 -1 30613 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 0 -1 30699 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 0 -1 30785 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 0 -1 30871 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 32591 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 0 -1 32677 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 0 -1 32763 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 0 -1 32849 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 0 -1 32935 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 0 -1 33021 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 0 -1 33107 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 0 -1 33193 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 0 -1 33279 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 0 -1 33365 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 0 -1 33451 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 0 -1 33537 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 0 -1 33623 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 0 -1 33709 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 0 -1 33795 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 0 -1 33881 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 0 -1 33967 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 0 -1 34053 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 0 -1 34139 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 0 -1 34225 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 0 -1 34311 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 0 -1 34397 1 0 39773
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 36117 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 0 -1 36203 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 0 -1 36289 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 0 -1 36375 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 0 -1 36461 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 0 -1 36547 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 0 -1 36633 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 0 -1 36719 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 0 -1 36805 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 0 -1 36891 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 0 -1 36977 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 0 -1 37063 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 0 -1 37149 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 0 -1 37235 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 0 -1 37321 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 0 -1 37407 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 0 -1 37493 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 0 -1 37579 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 0 -1 37665 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 0 -1 37751 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 0 -1 37837 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 0 -1 37923 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 39643 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 0 -1 39729 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 0 -1 39815 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 0 -1 39901 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 0 -1 39987 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 0 -1 40073 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 0 -1 40159 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 0 -1 40245 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 0 -1 40331 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 0 -1 40417 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 0 -1 40503 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 0 -1 40589 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 0 -1 40675 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 0 -1 40761 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 0 -1 40847 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 0 -1 40933 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 0 -1 41019 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 0 -1 41105 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 0 -1 41191 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 0 -1 41277 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 0 -1 41363 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 0 -1 41449 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 43169 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 0 -1 43255 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 0 -1 43341 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 0 -1 43427 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 0 -1 43513 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 0 -1 43599 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 0 -1 43685 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 0 -1 43771 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 0 -1 43857 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 0 -1 43943 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 0 -1 44029 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 0 -1 44115 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 0 -1 44201 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 0 -1 44287 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 0 -1 44373 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 0 -1 44459 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 0 -1 44545 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 0 -1 44631 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 0 -1 44717 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 0 -1 44803 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 0 -1 44889 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 0 -1 44975 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 46695 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 0 -1 46781 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 0 -1 46867 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 0 -1 46953 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 0 -1 47039 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 0 -1 47125 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 0 -1 47211 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 0 -1 47297 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 0 -1 47383 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 0 -1 47469 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 0 -1 47555 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 0 -1 47641 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 0 -1 47727 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 0 -1 47813 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 0 -1 47899 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 0 -1 47985 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 0 -1 48071 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 0 -1 48157 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 0 -1 48243 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 0 -1 48329 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 0 -1 48415 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 0 -1 48501 1 0 39773
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 50221 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 0 -1 50307 1 0 39773
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 56757 0 -1 46223
box 0 0 6450 6450
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 20207 0 -1 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform -1 0 20207 0 -1 38053
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform -1 0 20207 0 -1 37967
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform -1 0 20207 0 -1 37881
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform -1 0 20207 0 -1 37795
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform -1 0 20207 0 -1 37709
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform -1 0 20207 0 -1 37623
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform -1 0 20207 0 -1 37537
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform -1 0 20207 0 -1 37451
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform -1 0 20207 0 -1 37365
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform -1 0 20207 0 -1 37279
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform -1 0 20207 0 -1 37193
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform -1 0 20207 0 -1 37107
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform -1 0 20207 0 -1 37021
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform -1 0 20207 0 -1 36935
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform -1 0 20207 0 -1 36849
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform -1 0 20207 0 -1 36763
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform -1 0 20207 0 -1 36677
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform -1 0 20207 0 -1 36591
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform -1 0 20207 0 -1 36505
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform -1 0 20207 0 -1 36419
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform -1 0 20207 0 -1 36333
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform -1 0 20207 0 -1 36247
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform -1 0 20207 0 -1 36161
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform -1 0 20207 0 -1 36075
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform -1 0 20207 0 -1 35989
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform -1 0 20207 0 -1 35903
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform -1 0 20207 0 -1 35817
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 20207 0 -1 35731
box 0 0 6450 1720
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform -1 0 20207 0 -1 34011
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform -1 0 20207 0 -1 33925
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform -1 0 20207 0 -1 33839
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform -1 0 20207 0 -1 33753
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform -1 0 20207 0 -1 33667
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform -1 0 20207 0 -1 33581
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform -1 0 20207 0 -1 33495
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform -1 0 20207 0 -1 33409
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform -1 0 20207 0 -1 33323
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform -1 0 20207 0 -1 33237
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform -1 0 20207 0 -1 33151
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform -1 0 20207 0 -1 33065
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform -1 0 20207 0 -1 32979
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform -1 0 20207 0 -1 32893
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform -1 0 20207 0 -1 32807
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform -1 0 20207 0 -1 32721
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform -1 0 20207 0 -1 32635
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform -1 0 20207 0 -1 32549
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform -1 0 20207 0 -1 32463
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform -1 0 20207 0 -1 32377
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform -1 0 20207 0 -1 32291
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform -1 0 20207 0 -1 32205
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform -1 0 20207 0 -1 32119
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform -1 0 20207 0 -1 32033
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform -1 0 20207 0 -1 31947
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform -1 0 20207 0 -1 31861
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform -1 0 20207 0 -1 31775
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 20207 0 -1 31689
box 0 0 6450 1720
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform -1 0 20207 0 -1 29969
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform -1 0 20207 0 -1 29883
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform -1 0 20207 0 -1 29797
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform -1 0 20207 0 -1 29711
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform -1 0 20207 0 -1 29625
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform -1 0 20207 0 -1 29539
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform -1 0 20207 0 -1 29453
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform -1 0 20207 0 -1 29367
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform -1 0 20207 0 -1 29281
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform -1 0 20207 0 -1 29195
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform -1 0 20207 0 -1 29109
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform -1 0 20207 0 -1 29023
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform -1 0 20207 0 -1 28937
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform -1 0 20207 0 -1 28851
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform -1 0 20207 0 -1 28765
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform -1 0 20207 0 -1 28679
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform -1 0 20207 0 -1 28593
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform -1 0 20207 0 -1 28507
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform -1 0 20207 0 -1 28421
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform -1 0 20207 0 -1 28335
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform -1 0 20207 0 -1 28249
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform -1 0 20207 0 -1 28163
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform -1 0 20207 0 -1 28077
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform -1 0 20207 0 -1 27991
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform -1 0 20207 0 -1 27905
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform -1 0 20207 0 -1 27819
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform -1 0 20207 0 -1 27733
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 20207 0 -1 27647
box 0 0 6450 1720
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform -1 0 20207 0 -1 25927
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform -1 0 20207 0 -1 25841
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform -1 0 20207 0 -1 25755
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform -1 0 20207 0 -1 25669
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform -1 0 20207 0 -1 25583
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform -1 0 20207 0 -1 25497
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform -1 0 20207 0 -1 25411
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform -1 0 20207 0 -1 25325
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform -1 0 20207 0 -1 25239
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform -1 0 20207 0 -1 25153
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform -1 0 20207 0 -1 25067
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform -1 0 20207 0 -1 24981
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform -1 0 20207 0 -1 24895
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform -1 0 20207 0 -1 24809
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform -1 0 20207 0 -1 24723
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform -1 0 20207 0 -1 24637
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform -1 0 20207 0 -1 24551
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform -1 0 20207 0 -1 24465
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform -1 0 20207 0 -1 24379
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform -1 0 20207 0 -1 24293
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform -1 0 20207 0 -1 24207
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform -1 0 20207 0 -1 24121
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform -1 0 20207 0 -1 24035
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform -1 0 20207 0 -1 23949
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform -1 0 20207 0 -1 23863
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform -1 0 20207 0 -1 23777
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform -1 0 20207 0 -1 23691
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 20207 0 -1 23605
box 0 0 6450 1720
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform -1 0 20207 0 -1 21885
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform -1 0 20207 0 -1 21799
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform -1 0 20207 0 -1 21713
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform -1 0 20207 0 -1 21627
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform -1 0 20207 0 -1 21541
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform -1 0 20207 0 -1 21455
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform -1 0 20207 0 -1 21369
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform -1 0 20207 0 -1 21283
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform -1 0 20207 0 -1 21197
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform -1 0 20207 0 -1 21111
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform -1 0 20207 0 -1 21025
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform -1 0 20207 0 -1 20939
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform -1 0 20207 0 -1 20853
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform -1 0 20207 0 -1 20767
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform -1 0 20207 0 -1 20681
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform -1 0 20207 0 -1 20595
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform -1 0 20207 0 -1 20509
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform -1 0 20207 0 -1 20423
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform -1 0 20207 0 -1 20337
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform -1 0 20207 0 -1 20251
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform -1 0 20207 0 -1 20165
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform -1 0 20207 0 -1 20079
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform -1 0 20207 0 -1 19993
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform -1 0 20207 0 -1 19907
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform -1 0 20207 0 -1 19821
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform -1 0 20207 0 -1 19735
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform -1 0 20207 0 -1 19649
box 0 0 6450 86
use datapath datapath_0
timestamp 1396952988
transform 1 0 21535 0 1 19643
box 0 0 25408 19490
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 50307 0 1 38053
box 0 0 6450 1720
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 50307 0 1 37967
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 50307 0 1 37881
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 50307 0 1 37795
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 50307 0 1 37709
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 50307 0 1 37623
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 50307 0 1 37537
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 50307 0 1 37451
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 50307 0 1 37365
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 50307 0 1 37279
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 50307 0 1 37193
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 50307 0 1 37107
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 50307 0 1 37021
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 50307 0 1 36935
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 50307 0 1 36849
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 50307 0 1 36763
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 50307 0 1 36677
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 50307 0 1 36591
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 50307 0 1 36505
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 50307 0 1 36419
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 50307 0 1 36333
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 50307 0 1 36247
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 50307 0 1 36161
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 50307 0 1 36075
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 50307 0 1 35989
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 50307 0 1 35903
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 50307 0 1 35817
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 50307 0 1 35731
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 50307 0 1 34011
box 0 0 6450 1720
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 50307 0 1 33925
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 50307 0 1 33839
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 50307 0 1 33753
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 50307 0 1 33667
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 50307 0 1 33581
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 50307 0 1 33495
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 50307 0 1 33409
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 50307 0 1 33323
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 50307 0 1 33237
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 50307 0 1 33151
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 50307 0 1 33065
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 50307 0 1 32979
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 50307 0 1 32893
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 50307 0 1 32807
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 50307 0 1 32721
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 50307 0 1 32635
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 50307 0 1 32549
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 50307 0 1 32463
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 50307 0 1 32377
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 50307 0 1 32291
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 50307 0 1 32205
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 50307 0 1 32119
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 50307 0 1 32033
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 50307 0 1 31947
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 50307 0 1 31861
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 50307 0 1 31775
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 50307 0 1 31689
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 50307 0 1 29969
box 0 0 6450 1720
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 50307 0 1 29883
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 50307 0 1 29797
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 50307 0 1 29711
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 50307 0 1 29625
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 50307 0 1 29539
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 50307 0 1 29453
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 50307 0 1 29367
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 50307 0 1 29281
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 50307 0 1 29195
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 50307 0 1 29109
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 50307 0 1 29023
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 50307 0 1 28937
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 50307 0 1 28851
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 50307 0 1 28765
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 50307 0 1 28679
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 50307 0 1 28593
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 50307 0 1 28507
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 50307 0 1 28421
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 50307 0 1 28335
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 50307 0 1 28249
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 50307 0 1 28163
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 50307 0 1 28077
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 50307 0 1 27991
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 50307 0 1 27905
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 50307 0 1 27819
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 50307 0 1 27733
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 50307 0 1 27647
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 50307 0 1 25927
box 0 0 6450 1720
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 50307 0 1 25841
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 50307 0 1 25755
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 50307 0 1 25669
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 50307 0 1 25583
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 50307 0 1 25497
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 50307 0 1 25411
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 50307 0 1 25325
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 50307 0 1 25239
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 50307 0 1 25153
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 50307 0 1 25067
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 50307 0 1 24981
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 50307 0 1 24895
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 50307 0 1 24809
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 50307 0 1 24723
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 50307 0 1 24637
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 50307 0 1 24551
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 50307 0 1 24465
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 50307 0 1 24379
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 50307 0 1 24293
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 50307 0 1 24207
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 50307 0 1 24121
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 50307 0 1 24035
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 50307 0 1 23949
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 50307 0 1 23863
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 50307 0 1 23777
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 50307 0 1 23691
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 50307 0 1 23605
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 50307 0 1 21885
box 0 0 6450 1720
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 50307 0 1 21799
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 50307 0 1 21713
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 50307 0 1 21627
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 50307 0 1 21541
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 50307 0 1 21455
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 50307 0 1 21369
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 50307 0 1 21283
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 50307 0 1 21197
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 50307 0 1 21111
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 50307 0 1 21025
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 50307 0 1 20939
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 50307 0 1 20853
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 50307 0 1 20767
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 50307 0 1 20681
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 50307 0 1 20595
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 50307 0 1 20509
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 50307 0 1 20423
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 50307 0 1 20337
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 50307 0 1 20251
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 50307 0 1 20165
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 50307 0 1 20079
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 50307 0 1 19993
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 50307 0 1 19907
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 1 0 50307 0 1 19821
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 1 0 50307 0 1 19735
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 1 0 50307 0 1 19649
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 20207 0 -1 19563
box 0 0 6450 1720
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 1 0 50307 0 1 19563
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform -1 0 20207 0 -1 17843
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform -1 0 20207 0 -1 17757
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform -1 0 20207 0 -1 17671
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform -1 0 20207 0 -1 17585
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform -1 0 20207 0 -1 17499
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform -1 0 20207 0 -1 17413
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform -1 0 20207 0 -1 17327
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform -1 0 20207 0 -1 17241
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform -1 0 20207 0 -1 17155
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform -1 0 20207 0 -1 17069
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform -1 0 20207 0 -1 16983
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform -1 0 20207 0 -1 16897
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform -1 0 20207 0 -1 16811
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform -1 0 20207 0 -1 16725
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform -1 0 20207 0 -1 16639
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform -1 0 20207 0 -1 16553
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform -1 0 20207 0 -1 16467
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform -1 0 20207 0 -1 16381
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform -1 0 20207 0 -1 16295
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform -1 0 20207 0 -1 16209
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform -1 0 20207 0 -1 16123
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform -1 0 20207 0 -1 16037
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform -1 0 20207 0 -1 15951
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform -1 0 20207 0 -1 15865
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform -1 0 20207 0 -1 15779
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform -1 0 20207 0 -1 15693
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform -1 0 20207 0 -1 15607
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 20207 0 -1 15521
box 0 0 6450 1720
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform -1 0 20207 0 -1 13801
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform -1 0 20207 0 -1 13715
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform -1 0 20207 0 -1 13629
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform -1 0 20207 0 -1 13543
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform -1 0 20207 0 -1 13457
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform -1 0 20207 0 -1 13371
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform -1 0 20207 0 -1 13285
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform -1 0 20207 0 -1 13199
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform -1 0 20207 0 -1 13113
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform -1 0 20207 0 -1 13027
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform -1 0 20207 0 -1 12941
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform -1 0 20207 0 -1 12855
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 20207 0 -1 12769
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 20207 0 -1 12683
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 20207 0 -1 12597
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 20207 0 -1 12511
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 20207 0 -1 12425
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 20207 0 -1 12339
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 20207 0 -1 12253
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 20207 0 -1 12167
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 20207 0 -1 12081
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 20207 0 -1 11995
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 20207 0 -1 11909
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 20207 0 -1 11823
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 20207 0 -1 11737
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 20207 0 -1 11651
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 20207 0 -1 11565
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 20207 0 -1 11479
box 0 0 6450 1720
use control control_0
timestamp 1396952988
transform 1 0 21782 0 1 10294
box 0 0 26953 8588
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 50307 0 1 17843
box 0 0 6450 1720
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 1 0 50307 0 1 17757
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 1 0 50307 0 1 17671
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 1 0 50307 0 1 17585
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 1 0 50307 0 1 17499
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 1 0 50307 0 1 17413
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 1 0 50307 0 1 17327
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 1 0 50307 0 1 17241
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 1 0 50307 0 1 17155
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 1 0 50307 0 1 17069
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 1 0 50307 0 1 16983
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 1 0 50307 0 1 16897
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 1 0 50307 0 1 16811
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 1 0 50307 0 1 16725
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 1 0 50307 0 1 16639
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 1 0 50307 0 1 16553
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 1 0 50307 0 1 16467
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 1 0 50307 0 1 16381
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 1 0 50307 0 1 16295
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 1 0 50307 0 1 16209
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 1 0 50307 0 1 16123
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 1 0 50307 0 1 16037
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 1 0 50307 0 1 15951
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 1 0 50307 0 1 15865
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 1 0 50307 0 1 15779
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 1 0 50307 0 1 15693
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 1 0 50307 0 1 15607
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 1 0 50307 0 1 15521
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 50307 0 1 13801
box 0 0 6450 1720
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 1 0 50307 0 1 13715
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 1 0 50307 0 1 13629
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 1 0 50307 0 1 13543
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 1 0 50307 0 1 13457
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 1 0 50307 0 1 13371
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 1 0 50307 0 1 13285
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 1 0 50307 0 1 13199
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 1 0 50307 0 1 13113
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 1 0 50307 0 1 13027
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 1 0 50307 0 1 12941
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 1 0 50307 0 1 12855
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 1 0 50307 0 1 12769
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 1 0 50307 0 1 12683
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 1 0 50307 0 1 12597
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 1 0 50307 0 1 12511
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 1 0 50307 0 1 12425
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 1 0 50307 0 1 12339
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 1 0 50307 0 1 12253
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 1 0 50307 0 1 12167
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 1 0 50307 0 1 12081
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 1 0 50307 0 1 11995
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 1 0 50307 0 1 11909
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 1 0 50307 0 1 11823
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 1 0 50307 0 1 11737
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 1 0 50307 0 1 11651
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 1 0 50307 0 1 11565
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 1 0 50307 0 1 11479
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 50307 0 1 9759
box 0 0 6450 1720
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 13757 0 1 3309
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 20207 -1 0 9759
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 20293 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 22013 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 22099 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 22185 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 22271 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 22357 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 22443 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 22529 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 22615 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 22701 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 22787 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 22873 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 22959 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 23045 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 23131 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 23217 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 23303 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 23389 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 23475 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 23561 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 23647 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 23733 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 23819 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 25539 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 25625 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 25711 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 25797 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 25883 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 25969 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 26055 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 26141 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 26227 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 26313 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 26399 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 26485 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 26571 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 26657 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 26743 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 26829 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 26915 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 27001 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 27087 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 27173 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 27259 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 27345 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 29065 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 29151 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 29237 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 29323 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 29409 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 29495 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 29581 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 29667 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 29753 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 29839 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 29925 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 30011 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 30097 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 30183 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 30269 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 30355 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 30441 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 30527 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 30613 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 30699 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 30785 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 30871 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 32591 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 32677 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 32763 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 32849 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 32935 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 33021 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 33107 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 33193 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 33279 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 33365 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 33451 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 33537 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 33623 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 33709 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 33795 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 33881 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 33967 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 34053 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 34139 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 34225 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 34311 -1 0 9759
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 34397 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 36117 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 36203 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 36289 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 36375 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 36461 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 36547 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 36633 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 36719 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 36805 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 36891 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 36977 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 37063 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 37149 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 37235 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 37321 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 37407 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 37493 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 37579 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 37665 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 37751 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 37837 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 37923 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 39643 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 39729 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 39815 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 39901 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 39987 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 40073 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 40159 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 40245 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 40331 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 40417 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 40503 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 40589 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 40675 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 40761 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 40847 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 40933 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 41019 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 41105 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 41191 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 41277 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 41363 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 41449 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 43169 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 43255 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 43341 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 43427 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 43513 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 43599 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 43685 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 43771 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 43857 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 43943 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 44029 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 44115 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 44201 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 44287 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 44373 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 44459 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 44545 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 44631 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 44717 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 44803 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 44889 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 44975 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 46695 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 46781 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 46867 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 46953 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 47039 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 47125 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 47211 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 47297 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 47383 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 47469 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 47555 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 47641 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 47727 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 47813 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 47899 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 47985 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 48071 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 48157 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 48243 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 48329 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 48415 -1 0 9759
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 48501 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 50221 -1 0 9759
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 56757 1 0 3309
box 0 0 6450 6450
<< labels >>
rlabel metal4 20373 3387 21933 4947 0 nIRQ
rlabel metal4 23899 3387 25459 4947 0 Data[0]
rlabel metal4 27425 3387 28985 4947 0 Data[1]
rlabel metal4 30951 3387 32511 4947 0 Data[2]
rlabel metal4 34477 3387 36037 4947 0 vdde!
rlabel metal4 38003 3387 39563 4947 0 Data[3]
rlabel metal4 41529 3387 43089 4947 0 Data[4]
rlabel metal4 45055 3387 46615 4947 0 Data[5]
rlabel metal4 48581 3387 50141 4947 0 gnde!
rlabel metal4 55119 9839 56679 11399 0 Data[6]
rlabel metal4 55119 13881 56679 15441 0 Data[7]
rlabel metal4 55119 17923 56679 19483 0 Data[8]
rlabel metal4 55119 21965 56679 23525 0 gnde!
rlabel metal4 55119 26007 56679 27567 0 GND!
rlabel metal4 55119 30049 56679 31609 0 Data[9]
rlabel metal4 55119 34091 56679 35651 0 Data[10]
rlabel metal4 55119 38133 56679 39693 0 Data[11]
rlabel metal4 48581 44585 50141 46145 0 vdde!
rlabel metal4 45055 44585 46615 46145 0 Data[12]
rlabel metal4 41529 44585 43089 46145 0 Data[13]
rlabel metal4 38003 44585 39563 46145 0 Data[14]
rlabel metal4 34477 44585 36037 46145 0 gnde!
rlabel metal4 30951 44585 32511 46145 0 Data[15]
rlabel metal4 27425 44585 28985 46145 0 ALE
rlabel metal4 23899 44585 25459 46145 0 nME
rlabel metal4 20373 44585 21933 46145 0 nWait
rlabel metal4 13835 38133 15395 39693 0 nOE
rlabel metal4 13835 34091 15395 35651 0 RnW
rlabel metal4 13835 30049 15395 31609 0 SDO
rlabel metal4 13835 26007 15395 27567 0 Vdd!
rlabel metal4 13835 21965 15395 23525 0 SDI
rlabel metal4 13835 17923 15395 19483 0 Test
rlabel metal4 13835 13881 15395 15441 0 Clock
rlabel metal4 13835 9839 15395 11399 0 nReset
<< end >>
