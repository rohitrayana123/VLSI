magic
tech c035u
timestamp 1396308628
<< metal1 >>
rect 1573 1137 3215 1147
rect 3229 1137 20472 1147
rect 12552 1008 12623 1018
rect 12552 986 12863 996
rect 12901 987 13055 997
rect 13141 981 13176 991
rect 12709 959 13176 969
rect 12973 127 13103 137
rect 2821 94 12671 104
rect 0 72 3095 82
rect 3109 72 3263 82
rect 3277 72 20472 82
rect 0 50 12815 60
rect 0 28 20472 38
<< m2contact >>
rect 1559 1135 1573 1149
rect 3215 1135 3229 1149
rect 12623 1006 12637 1020
rect 12863 984 12877 998
rect 12887 983 12901 997
rect 13055 985 13069 999
rect 13127 979 13141 993
rect 12695 957 12709 971
rect 12959 123 12973 137
rect 13103 125 13117 139
rect 2807 93 2821 107
rect 12671 92 12685 106
rect 3095 70 3109 84
rect 3263 70 3277 84
rect 12815 48 12829 62
<< metal2 >>
rect 216 1043 228 1154
rect 360 1043 372 1154
rect 576 1043 588 1154
rect 1320 1043 1332 1154
rect 1488 1043 1500 1154
rect 1560 1043 1572 1135
rect 1872 1043 1884 1154
rect 2064 1043 2076 1154
rect 2280 1043 2292 1154
rect 3024 1043 3036 1154
rect 3192 954 3204 1154
rect 3216 954 3228 1135
rect 3288 1025 3372 1037
rect 3408 1025 3420 1154
rect 4152 1025 4164 1154
rect 4368 1025 4380 1154
rect 4560 1025 4572 1154
rect 5304 1025 5316 1154
rect 5520 1025 5532 1154
rect 5712 1025 5724 1154
rect 6456 1025 6468 1154
rect 6672 1025 6684 1154
rect 6864 1025 6876 1154
rect 7608 1025 7620 1154
rect 7824 1025 7836 1154
rect 8016 1025 8028 1154
rect 8760 1025 8772 1154
rect 8976 1025 8988 1154
rect 9168 1025 9180 1154
rect 9912 1025 9924 1154
rect 10128 1025 10140 1154
rect 10320 1025 10332 1154
rect 11064 1025 11076 1154
rect 11280 1025 11292 1154
rect 11472 1025 11484 1154
rect 12216 1025 12228 1154
rect 12432 1025 12444 1154
rect 3288 954 3300 1025
rect 12600 954 12612 1154
rect 12624 954 12636 1006
rect 12696 954 12708 957
rect 12792 954 12804 1154
rect 12864 954 12876 984
rect 12888 954 12900 983
rect 13032 954 13044 1154
rect 13248 1131 13260 1154
rect 13512 1131 13524 1154
rect 13680 1131 13692 1154
rect 13848 1131 13860 1154
rect 13872 1131 13884 1154
rect 13944 1131 13956 1154
rect 14160 1131 14172 1154
rect 14304 1131 14316 1154
rect 14640 1131 14652 1154
rect 15000 1131 15012 1154
rect 15408 1131 15420 1154
rect 15744 1131 15756 1154
rect 16056 1131 16068 1154
rect 16392 1131 16404 1154
rect 16512 1131 16524 1154
rect 16560 1131 16572 1154
rect 16728 1131 16740 1154
rect 16824 1131 16836 1154
rect 16872 1131 16884 1154
rect 16920 1131 16932 1154
rect 16968 1131 16980 1154
rect 17016 1131 17028 1154
rect 17064 1131 17076 1154
rect 17112 1131 17124 1154
rect 17160 1131 17172 1154
rect 17472 1131 17484 1154
rect 17520 1131 17532 1154
rect 17568 1131 17580 1154
rect 17616 1131 17628 1154
rect 17928 1131 17940 1154
rect 17976 1131 17988 1154
rect 18360 1131 18372 1154
rect 18528 1131 18540 1154
rect 18553 1131 18565 1154
rect 18600 1131 18612 1154
rect 18648 1131 18660 1154
rect 18696 1131 18708 1154
rect 18744 1131 18756 1154
rect 18792 1131 18804 1154
rect 18840 1131 18852 1154
rect 18888 1131 18900 1154
rect 18936 1131 18948 1154
rect 19176 1131 19188 1154
rect 19248 1131 19260 1154
rect 19296 1131 19308 1154
rect 19344 1131 19356 1154
rect 19392 1131 19404 1154
rect 19632 1131 19644 1154
rect 19704 1131 19716 1154
rect 19752 1131 19764 1154
rect 19992 1131 20004 1154
rect 20064 1131 20076 1154
rect 20352 1131 20364 1154
rect 13056 954 13068 985
rect 13128 954 13140 979
rect 216 0 228 126
rect 360 0 372 126
rect 576 0 588 126
rect 1320 0 1332 126
rect 1488 0 1500 126
rect 1872 0 1884 126
rect 2064 0 2076 126
rect 2280 0 2292 126
rect 2808 107 2820 126
rect 3024 0 3036 126
rect 3096 84 3108 126
rect 3192 0 3204 155
rect 3264 84 3276 155
rect 3408 0 3420 111
rect 4152 0 4164 111
rect 4368 0 4380 111
rect 4560 0 4572 111
rect 5304 0 5316 111
rect 5520 0 5532 111
rect 5712 0 5724 111
rect 6456 0 6468 111
rect 6672 0 6684 111
rect 6864 0 6876 111
rect 7608 0 7620 111
rect 7824 0 7836 111
rect 8016 0 8028 111
rect 8760 0 8772 111
rect 8976 0 8988 111
rect 9168 0 9180 111
rect 9912 0 9924 111
rect 10128 0 10140 111
rect 10320 0 10332 111
rect 11064 0 11076 111
rect 11280 0 11292 111
rect 11472 0 11484 111
rect 12216 0 12228 111
rect 12432 0 12444 111
rect 12600 0 12612 155
rect 12672 106 12684 155
rect 12792 0 12804 155
rect 12816 62 12828 155
rect 12960 137 12972 155
rect 13032 0 13044 155
rect 13104 139 13116 155
rect 13248 0 13260 89
rect 13512 0 13524 89
rect 13680 0 13692 89
rect 13872 0 13884 89
rect 14160 0 14172 89
rect 14304 0 14316 89
rect 14640 0 14652 89
rect 15000 0 15012 89
rect 15408 0 15420 89
rect 15744 0 15756 89
rect 16056 0 16068 89
rect 16392 0 16404 89
rect 16560 0 16572 89
rect 16728 0 16740 89
rect 16824 0 16836 89
rect 16872 0 16884 89
rect 16920 0 16932 89
rect 16968 0 16980 89
rect 17016 0 17028 89
rect 17064 0 17076 89
rect 17112 0 17124 89
rect 17160 0 17172 89
rect 17472 0 17484 89
rect 17520 0 17532 89
rect 17568 0 17580 89
rect 17616 0 17628 89
rect 17928 0 17940 89
rect 17976 0 17988 89
rect 18360 0 18372 89
rect 18528 0 18540 89
rect 18553 0 18565 89
rect 18600 0 18612 89
rect 18648 0 18660 89
rect 18696 0 18708 89
rect 18744 0 18756 89
rect 18792 0 18804 89
rect 18840 0 18852 89
rect 18888 0 18900 89
rect 18936 0 18948 89
rect 19176 0 19188 89
rect 19248 0 19260 89
rect 19296 0 19308 89
rect 19344 0 19356 89
rect 19392 0 19404 89
rect 19632 0 19644 89
rect 19704 0 19716 89
rect 19752 0 19764 89
rect 19992 0 20004 89
rect 20064 0 20076 89
rect 20352 0 20364 89
use Pc_slice Pc_slice_0
timestamp 1396307000
transform 1 0 0 0 1 89
box 0 37 3144 954
use mux2 mux2_0
timestamp 1386235218
transform 1 0 3144 0 1 155
box 0 0 192 799
use regBlock_slice regBlock_slice_0
timestamp 1396308165
transform 1 0 3336 0 1 110
box 0 0 9216 915
use mux2 mux2_1
timestamp 1386235218
transform 1 0 12552 0 1 155
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 12744 0 1 155
box 0 0 192 799
use tielow tielow_0
timestamp 1386086605
transform 1 0 12936 0 1 155
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 12984 0 1 155
box 0 0 192 799
use ALUSlice ALUSlice_0
timestamp 1396295595
transform 1 0 13176 0 1 89
box 0 0 7296 1042
<< labels >>
rlabel metal2 12792 1154 12804 1154 5 Op2Sel[0]
rlabel metal2 13032 1154 13044 1154 5 Op2Sel[1]
rlabel metal1 13163 985 13163 985 1 B
rlabel metal2 20064 1154 20076 1154 5 Sh1_R_in
rlabel metal2 16824 1154 16836 1154 5 Sh8Z_L
rlabel metal2 17160 1154 17172 1154 5 Sh8G_L
rlabel metal2 17064 1154 17076 1154 5 Sh8E_L
rlabel metal2 17112 1154 17124 1154 5 Sh8F_L
rlabel metal2 16920 1154 16932 1154 5 Sh8B_L
rlabel metal2 17016 1154 17028 1154 5 Sh8D_L
rlabel metal2 16968 1154 16980 1154 5 Sh8C_L
rlabel metal2 16872 1154 16884 1154 5 Sh8A_L
rlabel metal1 20472 1137 20472 1147 7 AluOut
rlabel metal2 16512 1154 16524 1154 5 A
rlabel metal2 18360 1154 18372 1154 5 Sh1_L_Out
rlabel metal2 18528 1154 18540 1154 5 Sh8
rlabel metal2 18696 1154 18708 1154 5 Sh8C_R
rlabel metal2 18648 1154 18660 1154 5 Sh8B_R
rlabel metal2 18600 1154 18612 1154 5 Sh8A_R
rlabel metal2 17616 1154 17628 1154 5 Sh4C_L
rlabel metal2 17568 1154 17580 1154 5 Sh4B_L
rlabel metal2 17976 1154 17988 1154 5 Sh2B_L
rlabel metal2 17928 1154 17940 1154 5 Sh2A_L
rlabel metal2 18553 1154 18565 1154 5 ShR
rlabel metal2 17520 1154 17532 1154 5 Sh4A_L
rlabel metal2 17472 1154 17484 1154 5 Sh4Z_L
rlabel metal2 19248 1154 19260 1154 5 Sh4Z_R
rlabel metal2 19992 1154 20004 1154 5 Sh1
rlabel metal2 19632 1154 19644 1154 5 Sh2
rlabel metal2 20352 1154 20364 1154 5 ShOut
rlabel metal2 19752 1154 19764 1154 5 Sh2B_R
rlabel metal2 19704 1154 19716 1154 5 Sh2A_R
rlabel metal2 19392 1154 19404 1154 5 Sh4C_R
rlabel metal2 19344 1154 19356 1154 5 Sh4B_R
rlabel metal2 19296 1154 19308 1154 5 Sh4A_R
rlabel metal2 19176 1154 19188 1154 5 Sh4
rlabel metal2 18744 1154 18756 1154 5 Sh8D_R
rlabel metal2 18792 1154 18804 1154 5 Sh8E_R
rlabel metal2 18840 1154 18852 1154 5 Sh8F_R
rlabel metal2 18888 1154 18900 1154 5 Sh8G_R
rlabel metal2 18936 1154 18948 1154 5 Sh8H_R
rlabel metal2 13248 1154 13260 1154 5 ZeroA
rlabel metal2 13680 1154 13692 1154 5 CIn
rlabel metal2 13944 1154 13956 1154 5 Sum
rlabel metal2 13872 1154 13884 1154 5 COut
rlabel metal2 16560 1154 16572 1154 5 ShB
rlabel metal2 16392 1154 16404 1154 5 NOR
rlabel metal2 16056 1154 16068 1154 5 NAND
rlabel metal2 15744 1154 15756 1154 5 NOT
rlabel metal2 15408 1154 15420 1154 5 XOR
rlabel metal2 15000 1154 15012 1154 5 OR
rlabel metal2 14640 1154 14652 1154 5 AND
rlabel metal2 13512 1154 13524 1154 5 SUB
rlabel metal2 14160 1154 14172 1154 5 nZ
rlabel metal2 14304 1154 14316 1154 5 FAOut
rlabel metal2 16728 1154 16740 1154 5 ShL
rlabel metal2 13848 1154 13860 1154 5 CIn_Slice
rlabel metal1 12815 965 12815 965 1 A
rlabel metal1 12942 1142 12942 1142 6 AluOut
rlabel metal2 12600 1154 12612 1154 5 Op1Sel
rlabel metal2 3192 1154 3204 1154 5 WdSel
rlabel metal2 3408 1154 3420 1154 5 Rw[0]
rlabel metal2 4152 1154 4164 1154 5 Rs1[0]
rlabel metal2 4368 1154 4380 1154 5 Rs2[0]
rlabel metal2 4560 1154 4572 1154 5 Rw[1]
rlabel metal2 5304 1154 5316 1154 5 Rs1[1]
rlabel metal2 5520 1154 5532 1154 5 Rs2[1]
rlabel metal2 5712 1154 5724 1154 5 Rw[2]
rlabel metal2 6456 1154 6468 1154 5 Rs1[2]
rlabel metal2 6672 1154 6684 1154 5 Rs2[2]
rlabel metal2 6864 1154 6876 1154 5 Rw[3]
rlabel metal2 7608 1154 7620 1154 5 Rs1[3]
rlabel metal2 7824 1154 7836 1154 5 Rs2[3]
rlabel metal2 8016 1154 8028 1154 5 Rw[4]
rlabel metal2 8760 1154 8772 1154 5 Rs1[4]
rlabel metal2 8976 1154 8988 1154 5 Rs2[4]
rlabel metal2 9168 1154 9180 1154 5 Rw[5]
rlabel metal2 10128 1154 10140 1154 5 Rs2[5]
rlabel metal2 9912 1154 9924 1154 5 Rs1[5]
rlabel metal2 10320 1154 10332 1154 5 Rw[6]
rlabel metal2 11064 1154 11076 1154 5 Rs1[6]
rlabel metal2 11280 1154 11292 1154 5 Rs2[6]
rlabel metal2 11472 1154 11484 1154 5 Rw[7]
rlabel metal2 12216 1154 12228 1154 5 Rs1[7]
rlabel metal2 12432 1154 12444 1154 5 Rs2[7]
rlabel metal2 3024 1154 3036 1154 5 PcEn
rlabel metal2 1872 1154 1884 1154 5 PcSel[1]
rlabel metal2 1488 1154 1500 1154 5 PcSel[0]
rlabel metal2 1320 1154 1332 1154 5 LrEn
rlabel metal2 576 1154 588 1154 5 LrWe
rlabel metal2 360 1154 372 1154 5 LrSel
rlabel metal2 216 1154 228 1154 5 PcIncCout
rlabel metal2 2280 1154 2292 1154 5 PcWe
rlabel metal2 2064 1154 2076 1154 5 PcSel[2]
rlabel metal1 12577 1013 12577 1013 1 Rd1
rlabel metal1 12579 991 12579 991 1 Rd2
rlabel metal2 3294 1031 3294 1031 1 WData
rlabel metal1 12546 99 12546 99 1 Pc
rlabel metal1 20472 72 20472 82 7 SysBus
rlabel metal1 12925 76 12925 76 1 SysBus
rlabel metal1 12544 77 12544 77 1 SysBus
rlabel metal1 3288 77 3288 77 1 SysBus
rlabel metal1 0 72 0 82 1 SysBus
rlabel metal1 12545 55 12545 55 1 Imm
rlabel metal1 0 50 0 60 1 Imm
rlabel metal2 13032 0 13044 0 1 Op2Sel[1]
rlabel metal2 17112 0 17124 0 1 Sh8G_L
rlabel metal2 17064 0 17076 0 1 Sh8F_L
rlabel metal2 17016 0 17028 0 1 Sh8E_L
rlabel metal2 16968 0 16980 0 1 Sh8D_L
rlabel metal2 18360 0 18372 0 1 Sh1_L_In
rlabel metal2 18600 0 18612 0 1 Sh8Z_R
rlabel metal2 18648 0 18660 0 1 Sh8A_R
rlabel metal2 18696 0 18708 0 1 Sh8B_R
rlabel metal2 17616 0 17628 0 1 Sh4D_L
rlabel metal2 17568 0 17580 0 1 Sh4C_L
rlabel metal2 17520 0 17532 0 1 Sh4B_L
rlabel metal2 17976 0 17988 0 1 Sh2C_L
rlabel metal2 17928 0 17940 0 1 Sh2B_L
rlabel metal2 18553 0 18565 0 1 ShR
rlabel metal2 18528 0 18540 0 1 Sh8
rlabel metal2 17472 0 17484 0 1 Sh4A_L
rlabel metal2 17160 0 17172 0 1 Sh8H_L
rlabel metal2 20064 0 20076 0 1 Sh1_R_Out
rlabel metal2 19752 0 19764 0 1 Sh2A_R
rlabel metal2 19704 0 19716 0 1 Sh2Z_R
rlabel metal2 19296 0 19308 0 1 Sh4Z_R
rlabel metal2 19344 0 19356 0 1 Sh4A_R
rlabel metal2 19392 0 19404 0 1 Sh4B_R
rlabel metal2 20352 0 20364 0 1 ShOut
rlabel metal2 19632 0 19644 0 1 Sh2
rlabel metal2 19992 0 20004 0 1 Sh1
rlabel metal2 19176 0 19188 0 1 Sh4
rlabel metal2 18744 0 18756 0 1 Sh8C_R
rlabel metal2 18792 0 18804 0 1 Sh8D_R
rlabel metal2 18840 0 18852 0 1 Sh8E_R
rlabel metal2 18888 0 18900 0 1 Sh8F_R
rlabel metal2 18936 0 18948 0 1 Sh8G_R
rlabel metal2 16824 0 16836 0 1 Sh8A_L
rlabel metal2 16920 0 16932 0 1 Sh8C_L
rlabel metal2 16872 0 16884 0 1 Sh8B_L
rlabel metal2 13248 0 13260 0 1 ZeroA
rlabel metal2 14304 0 14316 0 1 FAOut
rlabel metal2 13680 0 13692 0 1 CIn
rlabel metal2 14640 0 14652 0 1 AND
rlabel metal2 15000 0 15012 0 1 OR
rlabel metal2 15408 0 15420 0 1 XOR
rlabel metal2 15744 0 15756 0 1 NOT
rlabel metal2 16056 0 16068 0 1 NAND
rlabel metal2 16392 0 16404 0 1 NOR
rlabel metal2 16728 0 16740 0 1 ShL
rlabel metal2 16560 0 16572 0 1 ShB
rlabel metal2 13512 0 13524 0 1 SUB
rlabel metal2 14160 0 14172 0 1 nZ_prev
rlabel metal2 13872 0 13884 0 1 CIn_Slice
rlabel metal2 12792 0 12804 0 1 Op2Sel[0]
rlabel metal2 12600 0 12612 0 1 Op1Sel
rlabel metal2 4368 0 4380 0 1 Rs2[0]
rlabel metal2 3408 0 3420 0 1 Rw[0]
rlabel metal2 12432 0 12444 0 1 Rs2[7]
rlabel metal2 12216 0 12228 0 1 Rs1[7]
rlabel metal2 11472 0 11484 0 1 Rw[7]
rlabel metal2 11280 0 11292 0 1 Rs2[6]
rlabel metal2 11064 0 11076 0 1 Rs1[6]
rlabel metal2 10320 0 10332 0 1 Rw[6]
rlabel metal2 10128 0 10140 0 1 Rs2[5]
rlabel metal2 9912 0 9924 0 1 Rs1[5]
rlabel metal2 9168 0 9180 0 1 Rw[5]
rlabel metal2 8976 0 8988 0 1 Rs2[4]
rlabel metal2 8760 0 8772 0 1 Rs1[4]
rlabel metal2 8016 0 8028 0 1 Rw[4]
rlabel metal2 7824 0 7836 0 1 Rs2[3]
rlabel metal2 7608 0 7620 0 1 Rs1[3]
rlabel metal2 6864 0 6876 0 1 Rw[3]
rlabel metal2 6672 0 6684 0 1 Rs2[2]
rlabel metal2 6456 0 6468 0 1 Rs1[2]
rlabel metal2 5712 0 5724 0 1 Rw[2]
rlabel metal2 5520 0 5532 0 1 Rs2[1]
rlabel metal2 5304 0 5316 0 1 Rs1[1]
rlabel metal2 4560 0 4572 0 1 Rw[1]
rlabel metal2 4152 0 4164 0 1 Rs1[0]
rlabel metal2 3192 0 3204 0 1 WdSel
rlabel metal2 3024 0 3036 0 1 PcEn
rlabel metal2 2280 0 2292 0 1 PcWe
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 2064 0 2076 0 1 PcSel[2]
rlabel metal2 19248 0 19260 0 1 Sh4Y_R
rlabel metal1 0 28 0 38 3 DataIn
rlabel metal1 20472 28 20472 38 7 DataIn
<< end >>
