../behavioural/options.sv