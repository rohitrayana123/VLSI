magic
tech c035u
timestamp 1396388820
<< metal1 >>
rect 14 20163 14577 20173
rect 37 20139 14770 20149
rect 60 20115 14962 20125
rect 83 20091 15154 20101
rect 106 20067 15346 20077
rect 129 20043 4161 20053
rect 152 20019 4593 20029
rect 175 19995 4977 20005
rect 198 19971 4209 19981
rect 221 19947 4641 19957
rect 244 19923 5025 19933
rect 267 19899 7165 19909
rect 290 19875 7141 19885
rect 7155 19875 22353 19885
rect 313 19851 7117 19861
rect 7131 19851 22545 19861
rect 336 19827 22665 19837
rect 359 19803 22785 19813
rect 2879 18363 2890 18373
rect 14 17476 365 17486
rect 2842 17409 2890 17419
rect 25391 17409 25408 17419
rect 2842 17387 2890 17397
rect 2842 17365 2890 17375
rect 25391 17365 25408 17375
rect 2879 17209 2890 17219
rect 37 16322 365 16332
rect 2842 16255 2890 16265
rect 25391 16255 25408 16265
rect 2842 16233 2890 16243
rect 2842 16211 2890 16221
rect 25391 16211 25408 16221
rect 2879 16055 2890 16065
rect 60 15168 365 15178
rect 2842 15101 2890 15111
rect 25391 15101 25408 15111
rect 2842 15079 2890 15089
rect 2842 15057 2890 15067
rect 25391 15057 25408 15067
rect 2879 14901 2890 14911
rect 83 14014 365 14024
rect 2842 13947 2890 13957
rect 25391 13947 25408 13957
rect 2842 13925 2890 13935
rect 2842 13903 2890 13913
rect 25391 13903 25408 13913
rect 2879 13747 2890 13757
rect 106 12860 365 12870
rect 2842 12793 2890 12803
rect 25391 12793 25408 12803
rect 2842 12771 2890 12781
rect 2842 12749 2890 12759
rect 25391 12749 25408 12759
rect 2879 12593 2890 12603
rect 129 11706 365 11716
rect 2842 11639 2890 11649
rect 25391 11639 25408 11649
rect 2842 11617 2890 11627
rect 2842 11595 2890 11605
rect 25391 11595 25408 11605
rect 2879 11439 2890 11449
rect 152 10552 365 10562
rect 2842 10485 2890 10495
rect 25391 10485 25408 10495
rect 2842 10463 2890 10473
rect 2842 10441 2890 10451
rect 25391 10441 25408 10451
rect 2879 10285 2890 10295
rect 175 9398 365 9408
rect 2842 9331 2890 9341
rect 25391 9331 25408 9341
rect 2842 9309 2890 9319
rect 2842 9287 2890 9297
rect 25391 9287 25408 9297
rect 2879 9131 2890 9141
rect 198 8244 365 8254
rect 2842 8177 2890 8187
rect 25391 8177 25408 8187
rect 2842 8155 2890 8165
rect 2842 8133 2890 8143
rect 25391 8133 25408 8143
rect 2879 7977 2890 7987
rect 221 7090 365 7100
rect 2842 7023 2890 7033
rect 25391 7023 25408 7033
rect 2842 7001 2890 7011
rect 2842 6979 2890 6989
rect 25391 6979 25408 6989
rect 2879 6823 2890 6833
rect 244 5936 365 5946
rect 2842 5869 2890 5879
rect 25391 5869 25408 5879
rect 2842 5847 2890 5857
rect 2842 5825 2890 5835
rect 25391 5825 25408 5835
rect 2879 5669 2890 5679
rect 267 4782 365 4792
rect 2842 4715 2890 4725
rect 25391 4715 25408 4725
rect 2842 4693 2890 4703
rect 2842 4671 2890 4681
rect 25391 4671 25408 4681
rect 2879 4515 2890 4525
rect 290 3628 365 3638
rect 2842 3561 2890 3571
rect 25391 3561 25408 3571
rect 2842 3539 2890 3549
rect 2842 3517 2890 3527
rect 25391 3517 25408 3527
rect 2879 3361 2890 3371
rect 313 2474 365 2484
rect 2842 2407 2890 2417
rect 25391 2407 25408 2417
rect 2842 2385 2890 2395
rect 2842 2363 2890 2373
rect 25391 2363 25408 2373
rect 2879 2207 2890 2217
rect 336 1320 365 1330
rect 2842 1253 2890 1263
rect 25391 1253 25408 1263
rect 2842 1231 2890 1241
rect 2842 1209 2890 1219
rect 25391 1209 25408 1219
rect 2879 1053 2890 1063
rect 359 166 365 176
rect 2842 99 2890 109
rect 25391 99 25408 109
rect 2842 77 2890 87
rect 2842 55 2890 65
rect 25391 55 25408 65
rect 570 8 3105 18
rect 17063 7 19713 17
rect 19727 7 19760 17
rect 19774 7 19809 17
rect 19823 7 19857 17
rect 19871 7 19905 17
rect 19919 7 19953 17
rect 19967 7 20001 17
rect 20015 7 20049 17
rect 20063 7 20361 17
rect 20375 7 20409 17
rect 20423 7 20456 17
rect 20470 7 20505 17
rect 20519 7 20817 17
rect 20831 7 20865 17
rect 20879 7 21249 17
rect 21263 7 25186 17
<< m2contact >>
rect 0 20161 14 20175
rect 14577 20162 14591 20176
rect 23 20137 37 20151
rect 14770 20137 14784 20151
rect 46 20113 60 20127
rect 14962 20113 14976 20127
rect 69 20089 83 20103
rect 15154 20089 15168 20103
rect 92 20065 106 20079
rect 15346 20065 15360 20080
rect 115 20041 129 20055
rect 4161 20041 4175 20055
rect 138 20017 152 20031
rect 4593 20017 4607 20031
rect 161 19993 175 20007
rect 4977 19993 4991 20007
rect 184 19969 198 19983
rect 4209 19969 4223 19983
rect 207 19945 221 19959
rect 4641 19945 4655 19959
rect 230 19921 244 19935
rect 5025 19921 5039 19935
rect 253 19897 267 19911
rect 7165 19897 7179 19911
rect 276 19873 290 19887
rect 7141 19873 7155 19887
rect 22353 19873 22367 19887
rect 299 19849 313 19863
rect 7117 19849 7131 19863
rect 22545 19848 22559 19862
rect 322 19825 336 19839
rect 22665 19825 22679 19839
rect 345 19801 359 19815
rect 22785 19801 22799 19815
rect 2865 18361 2879 18375
rect 0 17474 14 17488
rect 2865 17207 2879 17221
rect 23 16320 37 16334
rect 2865 16053 2879 16067
rect 46 15166 60 15180
rect 2865 14899 2879 14913
rect 69 14012 83 14026
rect 2865 13745 2879 13759
rect 92 12858 106 12872
rect 2865 12591 2879 12605
rect 115 11704 129 11718
rect 2865 11437 2879 11451
rect 138 10550 152 10564
rect 2865 10283 2879 10297
rect 161 9396 175 9410
rect 2865 9129 2879 9143
rect 184 8242 198 8256
rect 2865 7975 2879 7989
rect 207 7088 221 7102
rect 2865 6821 2879 6835
rect 230 5934 244 5948
rect 2865 5667 2879 5681
rect 253 4780 267 4794
rect 2865 4513 2879 4527
rect 276 3626 290 3640
rect 2865 3359 2879 3373
rect 299 2472 313 2486
rect 2865 2205 2879 2219
rect 322 1318 336 1332
rect 2865 1051 2879 1065
rect 345 164 359 178
rect 556 6 570 20
rect 3105 5 3119 19
rect 17049 5 17063 19
rect 19713 5 19727 19
rect 19760 5 19774 19
rect 19809 5 19823 19
rect 19857 5 19871 19
rect 19905 5 19919 19
rect 19953 5 19967 19
rect 20001 5 20015 19
rect 20049 5 20063 19
rect 20361 5 20375 19
rect 20409 5 20423 19
rect 20456 5 20470 19
rect 20505 5 20519 19
rect 20817 5 20831 19
rect 20865 5 20879 19
rect 21249 5 21263 19
rect 25186 5 25200 19
<< metal2 >>
rect 1 17488 13 20161
rect 1 0 13 17474
rect 24 16334 36 20137
rect 24 0 36 16320
rect 47 15180 59 20113
rect 47 0 59 15166
rect 70 14026 82 20089
rect 70 0 82 14012
rect 93 12872 105 20065
rect 93 0 105 12858
rect 116 11718 128 20041
rect 116 0 128 11704
rect 139 10564 151 20017
rect 139 0 151 10550
rect 162 9410 174 19993
rect 162 0 174 9396
rect 185 8256 197 19969
rect 185 0 197 8242
rect 208 7102 220 19945
rect 208 0 220 7088
rect 231 5948 243 19921
rect 231 0 243 5934
rect 254 4794 266 19897
rect 254 0 266 4780
rect 277 3640 289 19873
rect 277 0 289 3626
rect 300 2486 312 19849
rect 300 0 312 2472
rect 323 1332 335 19825
rect 323 0 335 1318
rect 346 178 358 19801
rect 370 19793 570 20178
rect 586 19793 598 20178
rect 610 19793 622 20178
rect 634 19793 646 20178
rect 658 19793 670 20178
rect 4138 19793 4150 20178
rect 4162 19793 4174 20041
rect 4210 19793 4222 19969
rect 4378 19793 4390 20178
rect 4594 19793 4606 20017
rect 4642 19793 4654 19945
rect 4978 19793 4990 19993
rect 5026 19793 5038 19921
rect 5338 19793 5350 20178
rect 5530 19793 5542 20178
rect 6564 19793 6576 20178
rect 7118 19793 7130 19849
rect 7142 19793 7154 19873
rect 7166 19793 7178 19897
rect 14555 19793 14567 20178
rect 14579 19793 14591 20162
rect 14771 19793 14783 20137
rect 14819 19793 14831 20178
rect 14963 19793 14975 20113
rect 15155 19793 15167 20089
rect 15347 19793 15359 20065
rect 15539 19793 15551 20178
rect 17338 19793 17350 20178
rect 17530 19793 17542 20178
rect 17602 19793 17614 20178
rect 17698 19793 17710 20178
rect 22354 19793 22366 19873
rect 22546 19793 22558 19848
rect 22666 19793 22678 19825
rect 22786 19793 22798 19801
rect 25186 19793 25386 20178
rect 2866 18291 2878 18361
rect 2866 17137 2878 17207
rect 2866 15983 2878 16053
rect 2866 14829 2878 14899
rect 2866 13675 2878 13745
rect 2866 12521 2878 12591
rect 2866 11367 2878 11437
rect 2866 10213 2878 10283
rect 2866 9059 2878 9129
rect 2866 7905 2878 7975
rect 2866 6751 2878 6821
rect 2866 5597 2878 5667
rect 2866 4443 2878 4513
rect 2866 3289 2878 3359
rect 2866 2135 2878 2205
rect 2866 981 2878 1051
rect 346 0 358 164
rect 370 20 570 27
rect 370 6 556 20
rect 370 0 570 6
rect 586 0 598 27
rect 610 0 622 27
rect 634 0 646 27
rect 658 0 670 27
rect 1906 0 1918 27
rect 2698 0 2710 27
rect 3106 19 3118 27
rect 3250 0 3262 27
rect 3466 0 3478 27
rect 4210 0 4222 27
rect 4378 0 4390 27
rect 4762 0 4774 27
rect 4954 0 4966 27
rect 5170 0 5182 27
rect 5914 0 5926 27
rect 6082 0 6094 27
rect 15490 0 15502 27
rect 15682 0 15694 27
rect 15922 0 15934 27
rect 16570 21 16582 27
rect 16762 21 16774 27
rect 16570 9 16774 21
rect 17050 19 17062 27
rect 19714 19 19726 27
rect 19762 19 19774 27
rect 19810 19 19822 27
rect 19858 19 19870 27
rect 19906 19 19918 27
rect 19954 19 19966 27
rect 20002 19 20014 27
rect 20050 19 20062 27
rect 20362 19 20374 27
rect 20410 19 20422 27
rect 20458 19 20470 27
rect 20506 19 20518 27
rect 20818 19 20830 27
rect 20866 19 20878 27
rect 21250 19 21262 27
rect 23626 0 23638 27
rect 24370 0 24382 27
rect 24586 0 24598 27
rect 24730 0 24742 27
rect 24778 0 24790 27
rect 24826 0 24838 27
rect 24874 0 24886 27
rect 24946 0 24958 27
rect 25186 19 25386 27
rect 25200 5 25386 19
rect 25186 0 25386 5
use slice17 slice17_0
timestamp 1396388721
transform 1 0 370 0 1 18491
box 0 0 25016 1302
use leftbuf_slice leftbuf_slice_15
timestamp 1396386414
transform 1 0 365 0 1 17337
box 0 0 1469 1154
use IrAA IrAA_7
timestamp 1396382230
transform 1 0 1834 0 1 17337
box 0 0 1008 1154
use tielow tielow_0
timestamp 1386086605
transform 1 0 2842 0 1 17492
box 0 0 48 799
use leftbuf_slice leftbuf_slice_14
timestamp 1396386414
transform 1 0 365 0 1 16183
box 0 0 1469 1154
use IrAA IrAA_6
timestamp 1396382230
transform 1 0 1834 0 1 16183
box 0 0 1008 1154
use Datapath_slice Datapath_slice_15
timestamp 1396308628
transform 1 0 2890 0 1 17337
box 0 0 20472 1154
use LLIcell_U LLIcell_U_7
timestamp 1396314228
transform 1 0 23362 0 1 17337
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_11
timestamp 1396385716
transform 1 0 23554 0 1 17337
box 0 0 1837 1154
use tielow tielow_1
timestamp 1386086605
transform 1 0 2842 0 1 16338
box 0 0 48 799
use leftbuf_slice leftbuf_slice_13
timestamp 1396386414
transform 1 0 365 0 1 15029
box 0 0 1469 1154
use IrAA IrAA_5
timestamp 1396382230
transform 1 0 1834 0 1 15029
box 0 0 1008 1154
use Datapath_slice Datapath_slice_14
timestamp 1396308628
transform 1 0 2890 0 1 16183
box 0 0 20472 1154
use LLIcell_U LLIcell_U_6
timestamp 1396314228
transform 1 0 23362 0 1 16183
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_10
timestamp 1396385716
transform 1 0 23554 0 1 16183
box 0 0 1837 1154
use tielow tielow_2
timestamp 1386086605
transform 1 0 2842 0 1 15184
box 0 0 48 799
use leftbuf_slice leftbuf_slice_12
timestamp 1396386414
transform 1 0 365 0 1 13875
box 0 0 1469 1154
use IrAA IrAA_4
timestamp 1396382230
transform 1 0 1834 0 1 13875
box 0 0 1008 1154
use Datapath_slice Datapath_slice_13
timestamp 1396308628
transform 1 0 2890 0 1 15029
box 0 0 20472 1154
use LLIcell_U LLIcell_U_5
timestamp 1396314228
transform 1 0 23362 0 1 15029
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_9
timestamp 1396385716
transform 1 0 23554 0 1 15029
box 0 0 1837 1154
use tielow tielow_3
timestamp 1386086605
transform 1 0 2842 0 1 14030
box 0 0 48 799
use leftbuf_slice leftbuf_slice_11
timestamp 1396386414
transform 1 0 365 0 1 12721
box 0 0 1469 1154
use IrAA IrAA_3
timestamp 1396382230
transform 1 0 1834 0 1 12721
box 0 0 1008 1154
use Datapath_slice Datapath_slice_12
timestamp 1396308628
transform 1 0 2890 0 1 13875
box 0 0 20472 1154
use LLIcell_U LLIcell_U_4
timestamp 1396314228
transform 1 0 23362 0 1 13875
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_8
timestamp 1396385716
transform 1 0 23554 0 1 13875
box 0 0 1837 1154
use tielow tielow_4
timestamp 1386086605
transform 1 0 2842 0 1 12876
box 0 0 48 799
use leftbuf_slice leftbuf_slice_10
timestamp 1396386414
transform 1 0 365 0 1 11567
box 0 0 1469 1154
use IrAA IrAA_2
timestamp 1396382230
transform 1 0 1834 0 1 11567
box 0 0 1008 1154
use Datapath_slice Datapath_slice_11
timestamp 1396308628
transform 1 0 2890 0 1 12721
box 0 0 20472 1154
use LLIcell_U LLIcell_U_3
timestamp 1396314228
transform 1 0 23362 0 1 12721
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_7
timestamp 1396385716
transform 1 0 23554 0 1 12721
box 0 0 1837 1154
use tielow tielow_5
timestamp 1386086605
transform 1 0 2842 0 1 11722
box 0 0 48 799
use leftbuf_slice leftbuf_slice_9
timestamp 1396386414
transform 1 0 365 0 1 10413
box 0 0 1469 1154
use IrAA IrAA_1
timestamp 1396382230
transform 1 0 1834 0 1 10413
box 0 0 1008 1154
use Datapath_slice Datapath_slice_10
timestamp 1396308628
transform 1 0 2890 0 1 11567
box 0 0 20472 1154
use LLIcell_U LLIcell_U_2
timestamp 1396314228
transform 1 0 23362 0 1 11567
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_6
timestamp 1396385716
transform 1 0 23554 0 1 11567
box 0 0 1837 1154
use tielow tielow_6
timestamp 1386086605
transform 1 0 2842 0 1 10568
box 0 0 48 799
use leftbuf_slice leftbuf_slice_8
timestamp 1396386414
transform 1 0 365 0 1 9259
box 0 0 1469 1154
use IrAA IrAA_0
timestamp 1396382230
transform 1 0 1834 0 1 9259
box 0 0 1008 1154
use Datapath_slice Datapath_slice_9
timestamp 1396308628
transform 1 0 2890 0 1 10413
box 0 0 20472 1154
use LLIcell_U LLIcell_U_1
timestamp 1396314228
transform 1 0 23362 0 1 10413
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_5
timestamp 1396385716
transform 1 0 23554 0 1 10413
box 0 0 1837 1154
use tielow tielow_7
timestamp 1386086605
transform 1 0 2842 0 1 9414
box 0 0 48 799
use leftbuf_slice leftbuf_slice_7
timestamp 1396386414
transform 1 0 365 0 1 8105
box 0 0 1469 1154
use IrBA IrBA_2
timestamp 1396382245
transform 1 0 1834 0 1 8105
box 0 0 1008 1154
use Datapath_slice Datapath_slice_8
timestamp 1396308628
transform 1 0 2890 0 1 9259
box 0 0 20472 1154
use LLIcell_U LLIcell_U_0
timestamp 1396314228
transform 1 0 23362 0 1 9259
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_4
timestamp 1396385716
transform 1 0 23554 0 1 9259
box 0 0 1837 1154
use tielow tielow_8
timestamp 1386086605
transform 1 0 2842 0 1 8260
box 0 0 48 799
use leftbuf_slice leftbuf_slice_6
timestamp 1396386414
transform 1 0 365 0 1 6951
box 0 0 1469 1154
use IrBA IrBA_1
timestamp 1396382245
transform 1 0 1834 0 1 6951
box 0 0 1008 1154
use Datapath_slice Datapath_slice_7
timestamp 1396308628
transform 1 0 2890 0 1 8105
box 0 0 20472 1154
use LLIcell_L LLIcell_L_7
timestamp 1396313505
transform 1 0 23362 0 1 8105
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_3
timestamp 1396385716
transform 1 0 23554 0 1 8105
box 0 0 1837 1154
use tielow tielow_9
timestamp 1386086605
transform 1 0 2842 0 1 7106
box 0 0 48 799
use leftbuf_slice leftbuf_slice_5
timestamp 1396386414
transform 1 0 365 0 1 5797
box 0 0 1469 1154
use IrBA IrBA_0
timestamp 1396382245
transform 1 0 1834 0 1 5797
box 0 0 1008 1154
use Datapath_slice Datapath_slice_6
timestamp 1396308628
transform 1 0 2890 0 1 6951
box 0 0 20472 1154
use LLIcell_L LLIcell_L_6
timestamp 1396313505
transform 1 0 23362 0 1 6951
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_2
timestamp 1396385716
transform 1 0 23554 0 1 6951
box 0 0 1837 1154
use tielow tielow_10
timestamp 1386086605
transform 1 0 2842 0 1 5952
box 0 0 48 799
use leftbuf_slice leftbuf_slice_4
timestamp 1396386414
transform 1 0 365 0 1 4643
box 0 0 1469 1154
use IrBB IrBB_4
timestamp 1396382275
transform 1 0 1834 0 1 4643
box 0 0 1008 1154
use Datapath_slice Datapath_slice_5
timestamp 1396308628
transform 1 0 2890 0 1 5797
box 0 0 20472 1154
use LLIcell_L LLIcell_L_5
timestamp 1396313505
transform 1 0 23362 0 1 5797
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_1
timestamp 1396385716
transform 1 0 23554 0 1 5797
box 0 0 1837 1154
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 2842 0 1 4798
box 0 0 48 799
use leftbuf_slice leftbuf_slice_3
timestamp 1396386414
transform 1 0 365 0 1 3489
box 0 0 1469 1154
use IrBB IrBB_3
timestamp 1396382275
transform 1 0 1834 0 1 3489
box 0 0 1008 1154
use Datapath_slice Datapath_slice_4
timestamp 1396308628
transform 1 0 2890 0 1 4643
box 0 0 20472 1154
use LLIcell_L LLIcell_L_4
timestamp 1396313505
transform 1 0 23362 0 1 4643
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_0
timestamp 1396385716
transform 1 0 23554 0 1 4643
box 0 0 1837 1154
use tielow tielow_12
timestamp 1386086605
transform 1 0 2842 0 1 3644
box 0 0 48 799
use leftbuf_slice leftbuf_slice_2
timestamp 1396386414
transform 1 0 365 0 1 2335
box 0 0 1469 1154
use IrBB IrBB_2
timestamp 1396382275
transform 1 0 1834 0 1 2335
box 0 0 1008 1154
use Datapath_slice Datapath_slice_3
timestamp 1396308628
transform 1 0 2890 0 1 3489
box 0 0 20472 1154
use LLIcell_L LLIcell_L_3
timestamp 1396313505
transform 1 0 23362 0 1 3489
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_3
timestamp 1396386132
transform 1 0 23554 0 1 3489
box 0 0 1837 1154
use tielow tielow_13
timestamp 1386086605
transform 1 0 2842 0 1 2490
box 0 0 48 799
use leftbuf_slice leftbuf_slice_1
timestamp 1396386414
transform 1 0 365 0 1 1181
box 0 0 1469 1154
use IrBB IrBB_1
timestamp 1396382275
transform 1 0 1834 0 1 1181
box 0 0 1008 1154
use Datapath_slice Datapath_slice_2
timestamp 1396308628
transform 1 0 2890 0 1 2335
box 0 0 20472 1154
use LLIcell_L LLIcell_L_2
timestamp 1396313505
transform 1 0 23362 0 1 2335
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_2
timestamp 1396386132
transform 1 0 23554 0 1 2335
box 0 0 1837 1154
use tielow tielow_14
timestamp 1386086605
transform 1 0 2842 0 1 1336
box 0 0 48 799
use leftbuf_slice leftbuf_slice_0
timestamp 1396386414
transform 1 0 365 0 1 27
box 0 0 1469 1154
use IrBB IrBB_0
timestamp 1396382275
transform 1 0 1834 0 1 27
box 0 0 1008 1154
use Datapath_slice Datapath_slice_1
timestamp 1396308628
transform 1 0 2890 0 1 1181
box 0 0 20472 1154
use LLIcell_L LLIcell_L_1
timestamp 1396313505
transform 1 0 23362 0 1 1181
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_1
timestamp 1396386132
transform 1 0 23554 0 1 1181
box 0 0 1837 1154
use tielow tielow_15
timestamp 1386086605
transform 1 0 2842 0 1 182
box 0 0 48 799
use Datapath_slice Datapath_slice_0
timestamp 1396308628
transform 1 0 2890 0 1 27
box 0 0 20472 1154
use LLIcell_L LLIcell_L_0
timestamp 1396313505
transform 1 0 23362 0 1 27
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_0
timestamp 1396386132
transform 1 0 23554 0 1 27
box 0 0 1837 1154
<< labels >>
rlabel metal2 1 0 13 0 1 Ir[15]
rlabel metal2 24 0 36 0 1 Ir[14]
rlabel metal2 47 0 59 0 1 Ir[13]
rlabel metal2 70 0 82 0 1 Ir[12]
rlabel metal2 93 0 105 0 1 Ir[11]
rlabel metal2 116 0 128 0 1 Ir[10]
rlabel metal2 139 0 151 0 1 Ir[9]
rlabel metal2 162 0 174 0 1 Ir[8]
rlabel metal2 185 0 197 0 1 Ir[7]
rlabel metal2 208 0 220 0 1 Ir[6]
rlabel metal2 231 0 243 0 1 Ir[5]
rlabel metal2 254 0 266 0 1 Ir[4]
rlabel metal2 277 0 289 0 1 Ir[3]
rlabel metal2 300 0 312 0 1 Ir[2]
rlabel metal2 323 0 335 0 1 Ir[1]
rlabel metal2 346 0 358 0 1 Ir[0]
rlabel metal2 658 0 670 0 1 nReset
rlabel metal2 634 0 646 0 1 Clock
rlabel metal2 610 0 622 0 1 Test
rlabel metal2 586 0 598 0 1 SDI
rlabel metal2 370 0 570 0 1 Vdd!
rlabel metal2 24586 0 24598 0 1 MemEn
rlabel metal2 24946 0 24958 0 1 StatusRegEn
rlabel metal2 24730 0 24742 0 1 StatusReg[3]
rlabel metal2 24778 0 24790 0 1 StatusReg[2]
rlabel metal2 24826 0 24838 0 1 StatusReg[1]
rlabel metal2 24874 0 24886 0 1 StatusReg[0]
rlabel metal2 25186 0 25386 0 1 GND!
rlabel metal1 25408 55 25408 65 7 DataIn[0]
rlabel metal1 25408 99 25408 109 7 DataOut[0]
rlabel metal1 25408 17409 25408 17419 7 DataOut[15]
rlabel metal1 25408 17365 25408 17375 7 DataIn[15]
rlabel metal1 25408 16255 25408 16265 7 DataOut[14]
rlabel metal1 25408 16211 25408 16221 7 DataIn[14]
rlabel metal1 25408 15101 25408 15111 7 DataOut[13]
rlabel metal1 25408 15057 25408 15067 7 DataIn[13]
rlabel metal1 25408 13947 25408 13957 7 DataOut[12]
rlabel metal1 25408 13903 25408 13913 7 DataIn[12]
rlabel metal1 25408 12793 25408 12803 7 DataOut[11]
rlabel metal1 25408 12749 25408 12759 7 DataIn[11]
rlabel metal1 25408 11639 25408 11649 7 DataOut[10]
rlabel metal1 25408 11595 25408 11605 7 DataIn[10]
rlabel metal1 25408 10485 25408 10495 7 DataOut[9]
rlabel metal1 25408 10441 25408 10451 7 DataIn[9]
rlabel metal1 25408 9331 25408 9341 7 DataOut[8]
rlabel metal1 25408 9287 25408 9297 7 DataIn[8]
rlabel metal1 25408 8177 25408 8187 7 DataOut[7]
rlabel metal1 25408 8133 25408 8143 7 DataIn[7]
rlabel metal1 25408 7023 25408 7033 7 DataOut[6]
rlabel metal1 25408 6979 25408 6989 7 DataIn[6]
rlabel metal1 25408 5869 25408 5879 7 DataOut[5]
rlabel metal1 25408 5825 25408 5835 7 DataIn[5]
rlabel metal1 25408 4715 25408 4725 7 DataOut[4]
rlabel metal1 25408 4671 25408 4681 7 DataIn[4]
rlabel metal1 25408 3561 25408 3571 7 DataOut[3]
rlabel metal1 25408 3517 25408 3527 7 DataIn[3]
rlabel metal1 25408 2407 25408 2417 7 DataOut[2]
rlabel metal1 25408 2363 25408 2373 7 DataIn[2]
rlabel metal1 25408 1253 25408 1263 7 DataOut[1]
rlabel metal1 25408 1209 25408 1219 7 DataIn[1]
rlabel metal2 4210 0 4222 0 1 LrEn
rlabel metal2 4378 0 4390 0 1 PcSel[0]
rlabel metal2 4762 0 4774 0 1 PcSel[1]
rlabel metal2 23626 0 23638 0 1 AluWe
rlabel metal2 24370 0 24382 0 1 AluEn
rlabel metal2 5170 0 5182 0 1 PcWe
rlabel metal2 4954 0 4966 0 1 PcSel[2]
rlabel metal2 5914 0 5926 0 1 PcEn
rlabel metal2 6082 0 6094 0 1 WdSel
rlabel metal2 15490 0 15502 0 1 Op1Sel
rlabel metal2 15682 0 15694 0 1 Op2Sel[0]
rlabel metal2 15922 0 15934 0 1 Op2Sel[1]
rlabel metal2 1906 0 1918 0 1 IrWe
rlabel metal2 2698 0 2710 0 1 ImmSel
rlabel metal2 3466 0 3478 0 1 LrWe
rlabel metal2 3250 0 3262 0 1 LrSel
rlabel metal2 6 19866 6 19866 1 Ir[15]
rlabel metal2 30 19865 30 19865 1 Ir[14]
rlabel metal2 53 19865 53 19865 1 Ir[13]
rlabel metal2 76 19866 76 19866 1 Ir[12]
rlabel metal2 99 19866 99 19866 1 Ir[11]
rlabel metal2 122 19865 122 19865 1 Ir[10]
rlabel metal2 145 19866 145 19866 1 Ir[9]
rlabel metal2 168 19866 168 19866 1 Ir[8]
rlabel metal2 191 19868 191 19868 1 Ir[7]
rlabel metal2 214 19869 214 19869 1 Ir[6]
rlabel metal2 237 19870 237 19870 1 Ir[5]
rlabel metal2 260 19871 260 19871 1 Ir[4]
rlabel metal2 283 19870 283 19870 1 Ir[3]
rlabel metal2 22792 19796 22792 19796 1 Ir[0]
rlabel metal2 22671 19818 22671 19818 1 Ir[1]
rlabel metal2 22551 19843 22551 19843 1 Ir[2]
rlabel metal2 22360 19868 22360 19868 1 Ir[3]
rlabel metal2 14968 20107 14968 20107 1 Ir[13]
rlabel metal2 15161 20083 15161 20083 1 Ir[12]
rlabel metal2 15353 20058 15353 20058 1 Ir[11]
rlabel metal2 14775 20130 14775 20130 1 Ir[14]
rlabel metal2 14584 20155 14584 20155 1 Ir[15]
rlabel metal2 7122 19841 7122 19841 1 Ir[2]
rlabel metal2 7148 19865 7148 19865 1 Ir[3]
rlabel metal2 7171 19889 7171 19889 1 Ir[4]
rlabel metal2 4216 19961 4216 19961 1 Ir[7]
rlabel metal2 4167 20034 4167 20034 1 Ir[10]
rlabel metal2 4648 19938 4648 19938 1 Ir[6]
rlabel metal2 4599 20009 4599 20009 1 Ir[9]
rlabel metal2 4983 19986 4983 19986 1 Ir[8]
rlabel metal2 5033 19915 5033 19915 1 Ir[5]
rlabel metal2 6564 20178 6576 20178 5 RegWe
rlabel metal2 586 20178 598 20178 5 SDO
rlabel metal2 370 20178 570 20178 5 Vdd!
rlabel metal2 658 20178 670 20178 1 nReset
rlabel metal2 634 20178 646 20178 1 Clock
rlabel metal2 610 20178 622 20178 1 Test
rlabel metal2 17698 20178 17710 20178 5 Flags[0]
rlabel metal2 17602 20178 17614 20178 5 Flags[3]
rlabel metal2 17530 20178 17542 20178 5 Flags[1]
rlabel metal2 17338 20178 17350 20178 5 Flags[2]
rlabel metal2 14819 20178 14831 20178 5 AluOR[0]
rlabel metal2 14555 20178 14567 20178 5 AluOR[1]
rlabel metal2 15539 20178 15551 20178 5 CFlag
rlabel metal2 4138 20178 4150 20178 5 Rs1Sel[0]
rlabel metal2 4378 20178 4390 20178 5 Rs1Sel[1]
rlabel metal2 5338 20178 5350 20178 5 RwSel[0]
rlabel metal2 5530 20178 5542 20178 5 RwSel[1]
rlabel metal2 25186 20178 25386 20178 1 GND!
<< end >>
