magic
tech c035u
timestamp 1395577935
<< error_s >>
rect 10837 8083 10855 8090
<< nwell >>
rect 26979 1313 27531 1711
<< pwell >>
rect 26979 912 27531 1313
<< pohmic >>
rect 26979 988 26985 998
rect 27525 988 27531 998
<< nohmic >>
rect 26979 1648 26985 1658
rect 27525 1648 27531 1658
<< psubstratetap >>
rect 26985 988 27525 1004
<< nsubstratetap >>
rect 26985 1642 27525 1658
<< metal1 >>
rect 16048 9010 16066 9024
rect 9904 8988 16934 8998
rect 7288 8964 18458 8974
rect 3952 8938 3970 8952
rect 4144 8940 23030 8950
rect 2392 8914 2410 8928
rect 3256 8916 27554 8926
rect 2056 8892 24554 8902
rect 84 8868 22778 8878
rect 84 8844 20258 8854
rect 84 8820 11210 8830
rect 12328 8820 17282 8830
rect 17536 8820 26078 8830
rect 27520 8820 27626 8830
rect 2224 8796 13346 8806
rect 13360 8796 18698 8806
rect 18712 8796 27578 8806
rect 3688 8772 27530 8782
rect 27592 8772 27963 8782
rect 6184 8748 17138 8758
rect 19240 8748 19982 8758
rect 22744 8746 22762 8760
rect 25840 8748 27578 8758
rect 27616 8748 27963 8758
rect 7720 8724 23354 8734
rect 27592 8724 27963 8734
rect 9256 8700 19178 8710
rect 27568 8700 27963 8710
rect 9304 8676 27602 8686
rect 27640 8676 27963 8686
rect 10792 8652 11714 8662
rect 12376 8652 27963 8662
rect 13864 8628 14834 8638
rect 15400 8628 21098 8638
rect 27544 8628 27963 8638
rect 13144 7795 13346 7805
rect 13048 7771 13274 7781
rect 13024 7747 13202 7757
rect 13768 7747 13922 7757
rect 20536 7747 20762 7757
rect 20872 7747 21146 7757
rect 12952 7723 19274 7733
rect 19288 7723 19802 7733
rect 19816 7723 24146 7733
rect 12928 7699 15218 7709
rect 15232 7699 18146 7709
rect 18160 7699 19874 7709
rect 19888 7699 20282 7709
rect 20296 7699 20522 7709
rect 20536 7699 20858 7709
rect 20872 7699 23402 7709
rect 12784 7675 14450 7685
rect 24688 7675 24986 7685
rect 11872 7651 11930 7661
rect 12016 7651 12266 7661
rect 12736 7651 18074 7661
rect 18088 7651 23474 7661
rect 23488 7651 23522 7661
rect 23536 7651 24674 7661
rect 11824 7627 12866 7637
rect 12880 7627 26762 7637
rect 11584 7603 11618 7613
rect 11776 7603 21086 7613
rect 11488 7579 11546 7589
rect 11704 7579 13778 7589
rect 11416 7555 13850 7565
rect 11224 7531 11282 7541
rect 11296 7531 23138 7541
rect 11080 7507 27098 7517
rect 11008 7483 23786 7493
rect 10600 7459 11306 7469
rect 11392 7459 22730 7469
rect 10000 7435 10178 7445
rect 10336 7435 25346 7445
rect 9976 7411 14330 7421
rect 14344 7411 18482 7421
rect 9928 7387 26954 7397
rect 9856 7363 16874 7373
rect 9808 7339 10346 7349
rect 10360 7339 13562 7349
rect 13576 7339 17354 7349
rect 17368 7339 19322 7349
rect 19336 7339 20330 7349
rect 21640 7339 21698 7349
rect 9760 7315 18266 7325
rect 18280 7315 26714 7325
rect 9760 7291 9890 7301
rect 9952 7291 14354 7301
rect 14368 7291 16946 7301
rect 16960 7291 21626 7301
rect 9448 7267 13826 7277
rect 13840 7267 14618 7277
rect 9280 7243 11090 7253
rect 11104 7243 15986 7253
rect 16000 7243 17714 7253
rect 17728 7243 24890 7253
rect 9208 7219 18362 7229
rect 18376 7219 19634 7229
rect 19648 7219 20618 7229
rect 9160 7195 17498 7205
rect 24232 7195 24650 7205
rect 9016 7171 22538 7181
rect 22552 7171 24218 7181
rect 8728 7147 8738 7157
rect 8848 7147 10970 7157
rect 11032 7147 11066 7157
rect 11128 7147 21578 7157
rect 8608 7123 21122 7133
rect 8536 7099 14762 7109
rect 8512 7075 9362 7085
rect 9376 7075 17930 7085
rect 17944 7075 22466 7085
rect 22480 7075 23690 7085
rect 8464 7051 10874 7061
rect 10888 7051 12218 7061
rect 12232 7051 15074 7061
rect 8272 7027 14714 7037
rect 17968 7027 19538 7037
rect 7960 7003 17954 7013
rect 7864 6979 10778 6989
rect 10792 6979 14066 6989
rect 7648 6955 13754 6965
rect 7600 6931 12074 6941
rect 12088 6931 13634 6941
rect 13648 6931 17570 6941
rect 7552 6907 9242 6917
rect 9424 6907 12842 6917
rect 12856 6907 13490 6917
rect 13504 6907 13826 6917
rect 13840 6907 27026 6917
rect 7504 6883 8786 6893
rect 8800 6883 25922 6893
rect 7432 6859 8090 6869
rect 8176 6859 8282 6869
rect 8368 6859 19610 6869
rect 7384 6835 12482 6845
rect 12592 6835 21938 6845
rect 7360 6811 8186 6821
rect 8248 6811 27626 6821
rect 7336 6787 26138 6797
rect 7264 6763 19346 6773
rect 7072 6739 13010 6749
rect 13024 6739 16586 6749
rect 7072 6715 23282 6725
rect 7048 6691 15842 6701
rect 7024 6667 7034 6677
rect 7144 6667 12914 6677
rect 12928 6667 23234 6677
rect 6952 6643 16250 6653
rect 16264 6643 25706 6653
rect 6664 6619 23954 6629
rect 6520 6595 25730 6605
rect 6496 6571 21986 6581
rect 6448 6547 20978 6557
rect 6424 6523 16754 6533
rect 17248 6523 17306 6533
rect 18928 6523 20642 6533
rect 6376 6499 6914 6509
rect 6976 6499 18890 6509
rect 6352 6475 17210 6485
rect 17224 6475 20618 6485
rect 6304 6451 14258 6461
rect 14272 6451 16202 6461
rect 16216 6451 19562 6461
rect 6280 6427 11834 6437
rect 11848 6427 13514 6437
rect 13528 6427 17234 6437
rect 17248 6427 25682 6437
rect 25696 6427 26786 6437
rect 6208 6403 18314 6413
rect 18328 6403 18914 6413
rect 19024 6403 25082 6413
rect 6064 6379 20114 6389
rect 23512 6379 23810 6389
rect 5968 6355 13946 6365
rect 18304 6355 24026 6365
rect 5920 6331 6434 6341
rect 6448 6331 8066 6341
rect 8080 6331 14234 6341
rect 18016 6331 24122 6341
rect 5560 6307 7706 6317
rect 7720 6307 14954 6317
rect 14968 6307 26642 6317
rect 5560 6283 10634 6293
rect 10960 6283 17258 6293
rect 17464 6283 24962 6293
rect 5512 6259 12194 6269
rect 12304 6259 13790 6269
rect 17440 6259 21578 6269
rect 21592 6259 25370 6269
rect 5488 6235 8138 6245
rect 8152 6235 19898 6245
rect 21544 6235 26354 6245
rect 5464 6211 10322 6221
rect 10336 6211 19202 6221
rect 19216 6211 19298 6221
rect 19312 6211 21530 6221
rect 21544 6211 23498 6221
rect 5464 6187 27218 6197
rect 5440 6163 14114 6173
rect 15352 6163 15386 6173
rect 17392 6163 20426 6173
rect 20512 6163 20546 6173
rect 5416 6139 24794 6149
rect 5368 6115 9650 6125
rect 9736 6115 17138 6125
rect 17152 6115 21050 6125
rect 21064 6115 23714 6125
rect 23728 6115 25058 6125
rect 25072 6115 26570 6125
rect 5368 6091 16154 6101
rect 17080 6091 23450 6101
rect 5344 6067 21266 6077
rect 5320 6043 25274 6053
rect 5272 6019 19346 6029
rect 19360 6019 24410 6029
rect 5272 5995 16994 6005
rect 17056 5995 26474 6005
rect 5080 5971 26882 5981
rect 5032 5947 10418 5957
rect 10432 5947 20498 5957
rect 4984 5923 15338 5933
rect 16048 5923 26618 5933
rect 4936 5899 24530 5909
rect 4888 5875 19658 5885
rect 4864 5851 5042 5861
rect 5056 5851 9386 5861
rect 9400 5851 9554 5861
rect 9568 5851 10562 5861
rect 10576 5851 11882 5861
rect 11896 5851 13130 5861
rect 13144 5851 20594 5861
rect 20608 5851 22970 5861
rect 22984 5851 23258 5861
rect 23272 5851 26810 5861
rect 4792 5827 4946 5837
rect 4960 5827 6674 5837
rect 6688 5827 25898 5837
rect 4768 5803 9026 5813
rect 9040 5803 10634 5813
rect 10648 5803 11474 5813
rect 11488 5803 16442 5813
rect 16984 5803 24314 5813
rect 4744 5779 8594 5789
rect 8608 5779 9986 5789
rect 10000 5779 21722 5789
rect 4624 5755 5570 5765
rect 5584 5755 21890 5765
rect 4600 5731 7106 5741
rect 7192 5731 25778 5741
rect 4576 5707 20930 5717
rect 4528 5683 19586 5693
rect 26920 5683 27074 5693
rect 4432 5659 26906 5669
rect 4384 5635 20906 5645
rect 4360 5611 11690 5621
rect 11704 5611 15242 5621
rect 15256 5611 23618 5621
rect 4216 5587 7322 5597
rect 7336 5587 13082 5597
rect 13096 5587 23378 5597
rect 4096 5563 11330 5573
rect 11344 5563 15050 5573
rect 15280 5563 19010 5573
rect 4096 5539 25010 5549
rect 4048 5515 5882 5525
rect 5896 5515 23042 5525
rect 23872 5515 23882 5525
rect 4024 5491 6842 5501
rect 6856 5491 10610 5501
rect 10624 5491 16322 5501
rect 16336 5491 18290 5501
rect 18304 5491 20834 5501
rect 20848 5491 23162 5501
rect 23176 5491 23642 5501
rect 23656 5491 24098 5501
rect 24112 5491 24386 5501
rect 24400 5491 26882 5501
rect 26896 5491 27554 5501
rect 4000 5467 6290 5477
rect 6304 5467 7994 5477
rect 8008 5467 8474 5477
rect 8488 5467 17186 5477
rect 17200 5467 23858 5477
rect 3952 5443 6650 5453
rect 6736 5443 7730 5453
rect 7840 5443 7850 5453
rect 7936 5443 7946 5453
rect 8008 5443 8066 5453
rect 8128 5443 10730 5453
rect 10912 5443 13322 5453
rect 13336 5443 23090 5453
rect 3880 5419 13994 5429
rect 15112 5419 20762 5429
rect 3880 5395 19682 5405
rect 3856 5371 4226 5381
rect 4240 5371 7298 5381
rect 7312 5371 7634 5381
rect 7648 5371 7802 5381
rect 7816 5371 8114 5381
rect 8128 5371 8570 5381
rect 8584 5371 14282 5381
rect 14296 5371 16514 5381
rect 16528 5371 16946 5381
rect 16960 5371 23930 5381
rect 23944 5371 24362 5381
rect 3856 5347 6554 5357
rect 6712 5347 10538 5357
rect 10552 5347 14114 5357
rect 14128 5347 18146 5357
rect 3808 5323 7394 5333
rect 7480 5323 19082 5333
rect 20200 5323 20258 5333
rect 3784 5299 7682 5309
rect 7696 5299 26234 5309
rect 3784 5275 6122 5285
rect 6184 5275 17090 5285
rect 17104 5275 18122 5285
rect 20104 5275 27578 5285
rect 3736 5251 12314 5261
rect 12376 5251 12386 5261
rect 12568 5251 13178 5261
rect 14800 5251 24770 5261
rect 3640 5227 14018 5237
rect 14032 5227 17690 5237
rect 17752 5227 27963 5237
rect 3592 5203 20210 5213
rect 22048 5203 22130 5213
rect 3544 5179 11642 5189
rect 11728 5179 15098 5189
rect 15208 5179 22058 5189
rect 3520 5155 5738 5165
rect 5848 5155 17978 5165
rect 17992 5155 21290 5165
rect 21304 5155 25562 5165
rect 25576 5155 25706 5165
rect 3424 5131 25850 5141
rect 3400 5107 25634 5117
rect 3328 5083 7922 5093
rect 7936 5083 8450 5093
rect 8464 5083 9482 5093
rect 9496 5083 11042 5093
rect 11056 5083 18986 5093
rect 20032 5083 20234 5093
rect 20320 5083 20354 5093
rect 20464 5083 20738 5093
rect 21016 5083 26738 5093
rect 3232 5059 6554 5069
rect 6568 5059 11018 5069
rect 11032 5059 19922 5069
rect 19936 5059 21002 5069
rect 22024 5059 27458 5069
rect 3160 5035 19058 5045
rect 19072 5035 22826 5045
rect 3112 5011 4178 5021
rect 4192 5011 17018 5021
rect 17032 5011 17786 5021
rect 17800 5011 26306 5021
rect 3064 4987 27146 4997
rect 3016 4963 3914 4973
rect 3928 4963 13034 4973
rect 14704 4963 24458 4973
rect 24472 4963 25682 4973
rect 2968 4939 16826 4949
rect 16840 4939 21374 4949
rect 21388 4939 24338 4949
rect 2944 4915 27122 4925
rect 2920 4891 20474 4901
rect 21880 4891 22106 4901
rect 22960 4891 23210 4901
rect 23224 4891 23534 4901
rect 2800 4867 24002 4877
rect 2752 4843 8210 4853
rect 8224 4843 20066 4853
rect 20080 4843 20378 4853
rect 20392 4843 22034 4853
rect 22864 4843 23186 4853
rect 23344 4843 23654 4853
rect 2680 4819 4826 4829
rect 4840 4819 7010 4829
rect 7024 4819 10418 4829
rect 10480 4819 13730 4829
rect 13984 4819 21242 4829
rect 21256 4819 23594 4829
rect 23608 4819 24242 4829
rect 24304 4819 24542 4829
rect 24616 4819 24806 4829
rect 25504 4819 25610 4829
rect 25816 4819 25826 4829
rect 25888 4819 26978 4829
rect 2536 4795 6602 4805
rect 6616 4795 16106 4805
rect 16120 4795 19706 4805
rect 19720 4795 24722 4805
rect 24736 4795 27314 4805
rect 2464 4771 8666 4781
rect 8680 4771 9338 4781
rect 9352 4771 13970 4781
rect 13984 4771 14426 4781
rect 14584 4771 17594 4781
rect 17608 4771 26690 4781
rect 26968 4771 27338 4781
rect 2440 4747 14930 4757
rect 14944 4747 24290 4757
rect 24976 4747 25082 4757
rect 26656 4747 26714 4757
rect 2344 4723 23738 4733
rect 24016 4723 26426 4733
rect 26704 4723 26978 4733
rect 2320 4699 2450 4709
rect 2464 4699 4538 4709
rect 4552 4699 4970 4709
rect 4984 4699 8258 4709
rect 8272 4699 10658 4709
rect 10672 4699 10706 4709
rect 10720 4699 12626 4709
rect 12640 4699 14378 4709
rect 14392 4699 14546 4709
rect 14560 4699 18026 4709
rect 18040 4699 20186 4709
rect 20200 4699 25538 4709
rect 2296 4675 11906 4685
rect 12040 4675 21770 4685
rect 22072 4675 27602 4685
rect 2248 4651 23978 4661
rect 2200 4627 7826 4637
rect 7840 4627 11762 4637
rect 11776 4627 11858 4637
rect 11872 4627 23018 4637
rect 2152 4603 21410 4613
rect 2128 4579 5498 4589
rect 5512 4579 19130 4589
rect 19144 4579 23906 4589
rect 23920 4579 23954 4589
rect 23968 4579 24938 4589
rect 24952 4579 25442 4589
rect 2008 4555 10298 4565
rect 10312 4555 18194 4565
rect 18544 4555 24542 4565
rect 1984 4531 9098 4541
rect 9112 4531 18962 4541
rect 18976 4531 21338 4541
rect 23920 4531 24146 4541
rect 1936 4507 15482 4517
rect 15760 4507 24482 4517
rect 1912 4483 22082 4493
rect 1912 4459 24842 4469
rect 1864 4435 2570 4445
rect 2632 4435 8042 4445
rect 8056 4435 9218 4445
rect 9232 4435 17066 4445
rect 17176 4435 17282 4445
rect 18736 4435 25514 4445
rect 1816 4411 7442 4421
rect 7456 4411 10154 4421
rect 10168 4411 10874 4421
rect 10888 4411 20786 4421
rect 20800 4411 20882 4421
rect 20992 4411 21086 4421
rect 21352 4411 21374 4421
rect 1792 4387 6626 4397
rect 6760 4387 12530 4397
rect 12544 4387 13274 4397
rect 13288 4387 19754 4397
rect 20920 4387 24986 4397
rect 1768 4363 3602 4373
rect 3616 4363 9818 4373
rect 9832 4363 12458 4373
rect 12472 4363 20666 4373
rect 1744 4339 4418 4349
rect 4432 4339 5138 4349
rect 5152 4339 14882 4349
rect 14896 4339 20714 4349
rect 20728 4339 27530 4349
rect 1672 4315 19274 4325
rect 1672 4291 4250 4301
rect 4336 4291 5690 4301
rect 5704 4291 8714 4301
rect 8728 4291 12434 4301
rect 12448 4291 16730 4301
rect 16744 4291 20378 4301
rect 1648 4267 19442 4277
rect 1624 4243 3074 4253
rect 3088 4243 3290 4253
rect 3304 4243 5786 4253
rect 5800 4243 13418 4253
rect 13432 4243 14594 4253
rect 14608 4243 22634 4253
rect 22648 4243 24578 4253
rect 84 4219 1682 4229
rect 1744 4219 2546 4229
rect 2632 4219 4442 4229
rect 4456 4219 6698 4229
rect 6712 4219 7130 4229
rect 7144 4219 11978 4229
rect 11992 4219 14210 4229
rect 14224 4219 20834 4229
rect 20848 4219 21074 4229
rect 21088 4219 21650 4229
rect 21664 4219 24602 4229
rect 84 4195 14882 4205
rect 15064 4195 15074 4205
rect 15928 4195 16706 4205
rect 16720 4195 22994 4205
rect 84 4171 8306 4181
rect 8368 4171 26834 4181
rect 84 4147 25394 4157
rect 1624 4123 3458 4133
rect 3472 4123 14810 4133
rect 14872 4123 17834 4133
rect 18784 4123 19226 4133
rect 1888 4099 11906 4109
rect 12112 4099 13706 4109
rect 14248 4099 14258 4109
rect 14800 4099 21554 4109
rect 21568 4099 22682 4109
rect 2104 4075 14978 4085
rect 16528 4075 16586 4085
rect 16672 4075 20954 4085
rect 2272 4051 4994 4061
rect 5008 4051 11594 4061
rect 11608 4051 19466 4061
rect 19480 4051 21218 4061
rect 21232 4051 21818 4061
rect 2320 4027 3746 4037
rect 3760 4027 7658 4037
rect 7672 4027 9122 4037
rect 9136 4027 10298 4037
rect 10312 4027 10514 4037
rect 10528 4027 17906 4037
rect 17920 4027 22658 4037
rect 22672 4027 23330 4037
rect 23344 4027 23618 4037
rect 2392 4003 21026 4013
rect 2488 3979 8162 3989
rect 8248 3979 9530 3989
rect 9616 3979 16898 3989
rect 16912 3979 20738 3989
rect 2512 3955 16826 3965
rect 16840 3955 26090 3965
rect 2560 3931 9530 3941
rect 9544 3931 12482 3941
rect 12496 3931 12650 3941
rect 12664 3931 14402 3941
rect 14416 3931 21938 3941
rect 2584 3907 8018 3917
rect 8032 3907 16754 3917
rect 16768 3907 18650 3917
rect 18664 3907 18866 3917
rect 18880 3907 21866 3917
rect 21880 3907 26186 3917
rect 26200 3907 27002 3917
rect 2680 3883 10274 3893
rect 10288 3883 18002 3893
rect 18952 3883 19178 3893
rect 2776 3859 27963 3869
rect 2800 3835 7898 3845
rect 7912 3835 23570 3845
rect 23584 3835 24842 3845
rect 24856 3835 24914 3845
rect 2824 3811 3962 3821
rect 3976 3811 4394 3821
rect 4408 3811 11258 3821
rect 11272 3811 11570 3821
rect 11584 3811 12170 3821
rect 12184 3811 13610 3821
rect 13624 3811 22946 3821
rect 22960 3811 23402 3821
rect 23416 3811 26210 3821
rect 2848 3787 7466 3797
rect 7528 3787 12794 3797
rect 12808 3787 13202 3797
rect 13216 3787 13226 3797
rect 13240 3787 14426 3797
rect 14440 3787 23834 3797
rect 2872 3763 22970 3773
rect 2920 3739 3458 3749
rect 3472 3739 10682 3749
rect 10696 3739 19970 3749
rect 19984 3739 23114 3749
rect 23128 3739 24806 3749
rect 24820 3739 25034 3749
rect 25048 3739 25802 3749
rect 3208 3715 24122 3725
rect 3352 3691 5282 3701
rect 5344 3691 11522 3701
rect 11536 3691 12098 3701
rect 12160 3691 21362 3701
rect 3424 3667 5810 3677
rect 5824 3667 7946 3677
rect 7960 3667 9506 3677
rect 9520 3667 11618 3677
rect 11632 3667 14402 3677
rect 14416 3667 14594 3677
rect 14608 3667 14666 3677
rect 14680 3667 16970 3677
rect 16984 3667 24266 3677
rect 24280 3667 25250 3677
rect 25264 3667 26546 3677
rect 3664 3643 4682 3653
rect 4696 3643 5114 3653
rect 5128 3643 13946 3653
rect 13960 3643 22322 3653
rect 3760 3619 7106 3629
rect 7120 3619 7610 3629
rect 7624 3619 10850 3629
rect 10864 3619 19154 3629
rect 19168 3619 23354 3629
rect 23368 3619 24434 3629
rect 24448 3619 26666 3629
rect 3832 3595 3938 3605
rect 3952 3595 6818 3605
rect 6832 3595 8330 3605
rect 8344 3595 9890 3605
rect 9904 3595 12242 3605
rect 12256 3595 21458 3605
rect 21472 3595 23786 3605
rect 24448 3595 27194 3605
rect 3904 3571 8762 3581
rect 8920 3571 14822 3581
rect 14836 3571 26594 3581
rect 4168 3547 4658 3557
rect 4672 3547 9698 3557
rect 9712 3547 10274 3557
rect 10288 3547 13658 3557
rect 13672 3547 17810 3557
rect 17824 3547 21554 3557
rect 21568 3547 23426 3557
rect 26608 3547 26618 3557
rect 4216 3523 4298 3533
rect 4312 3523 8930 3533
rect 8944 3523 12746 3533
rect 12760 3523 13154 3533
rect 13168 3523 13466 3533
rect 13480 3523 19370 3533
rect 19384 3523 23534 3533
rect 23548 3523 26330 3533
rect 4312 3499 21962 3509
rect 4456 3475 12410 3485
rect 12424 3475 25106 3485
rect 4480 3451 6482 3461
rect 6544 3451 10370 3461
rect 10384 3451 27050 3461
rect 4528 3427 18050 3437
rect 4552 3403 8282 3413
rect 8392 3403 21434 3413
rect 4576 3379 12338 3389
rect 12352 3379 12674 3389
rect 12688 3379 20162 3389
rect 4648 3355 13514 3365
rect 13528 3355 25154 3365
rect 4672 3331 6938 3341
rect 6952 3331 15002 3341
rect 15016 3331 15122 3341
rect 17104 3331 17258 3341
rect 4720 3307 7226 3317
rect 7240 3307 26546 3317
rect 4768 3283 6722 3293
rect 6736 3283 8666 3293
rect 8680 3283 8738 3293
rect 8752 3283 12578 3293
rect 12592 3283 12818 3293
rect 12832 3283 13106 3293
rect 13120 3283 17882 3293
rect 17896 3283 21962 3293
rect 4816 3259 5210 3269
rect 5224 3259 19514 3269
rect 4864 3235 11786 3245
rect 11800 3235 20690 3245
rect 20704 3235 22586 3245
rect 4888 3211 5162 3221
rect 5176 3211 16850 3221
rect 16864 3211 21314 3221
rect 21328 3211 22922 3221
rect 4936 3187 17330 3197
rect 5104 3163 9602 3173
rect 9616 3163 11138 3173
rect 11152 3163 19994 3173
rect 20008 3163 21842 3173
rect 21856 3163 22562 3173
rect 22576 3163 23882 3173
rect 23896 3163 26330 3173
rect 5128 3139 6386 3149
rect 6472 3139 7802 3149
rect 7816 3139 13898 3149
rect 14296 3139 14450 3149
rect 14680 3139 27362 3149
rect 5200 3115 6866 3125
rect 6880 3115 18098 3125
rect 5416 3091 11954 3101
rect 11968 3091 13298 3101
rect 13600 3091 14186 3101
rect 14200 3091 15026 3101
rect 15040 3091 23522 3101
rect 23536 3091 27410 3101
rect 5536 3067 5618 3077
rect 5632 3067 25466 3077
rect 25480 3067 26522 3077
rect 5680 3043 22490 3053
rect 5704 3019 6074 3029
rect 6160 3019 20330 3029
rect 6016 2995 16154 3005
rect 17224 2995 21410 3005
rect 21424 2995 24650 3005
rect 6040 2971 23066 2981
rect 6064 2947 15386 2957
rect 17296 2947 20570 2957
rect 20584 2947 24386 2957
rect 6112 2923 7034 2933
rect 7048 2923 23042 2933
rect 6232 2899 24050 2909
rect 6616 2875 18866 2885
rect 18880 2875 20954 2885
rect 20968 2875 24746 2885
rect 6640 2851 6674 2861
rect 6784 2851 25994 2861
rect 6808 2827 7538 2837
rect 7552 2827 9578 2837
rect 9592 2827 10490 2837
rect 10504 2827 11642 2837
rect 11656 2827 12674 2837
rect 12688 2827 14498 2837
rect 14512 2827 19442 2837
rect 19456 2827 21194 2837
rect 21208 2827 21746 2837
rect 21760 2827 24074 2837
rect 24088 2827 25586 2837
rect 25600 2827 26378 2837
rect 6832 2803 8642 2813
rect 8656 2803 14306 2813
rect 14320 2803 25490 2813
rect 6904 2779 15026 2789
rect 15040 2779 17306 2789
rect 18112 2779 18122 2789
rect 20584 2779 23654 2789
rect 24088 2779 24242 2789
rect 7216 2755 17642 2765
rect 17656 2755 21914 2765
rect 7240 2731 7850 2741
rect 7864 2731 11354 2741
rect 11368 2731 12266 2741
rect 12280 2731 13346 2741
rect 13360 2731 14474 2741
rect 14488 2731 20306 2741
rect 20320 2731 21842 2741
rect 21856 2731 26282 2741
rect 7264 2707 26402 2717
rect 7360 2683 16370 2693
rect 16384 2683 23978 2693
rect 23992 2683 25610 2693
rect 7384 2659 13682 2669
rect 13744 2659 21146 2669
rect 21208 2659 22898 2669
rect 7696 2635 7706 2645
rect 7768 2635 9674 2645
rect 9688 2635 12818 2645
rect 12832 2635 20810 2645
rect 20824 2635 24170 2645
rect 24184 2635 24866 2645
rect 7744 2611 8618 2621
rect 8944 2611 10106 2621
rect 10216 2611 26858 2621
rect 7888 2587 10010 2597
rect 10024 2587 11546 2597
rect 11560 2587 12770 2597
rect 12784 2587 19490 2597
rect 19504 2587 20162 2597
rect 24184 2587 24458 2597
rect 8056 2563 8138 2573
rect 8440 2563 9482 2573
rect 9496 2563 10922 2573
rect 10936 2563 13874 2573
rect 13888 2563 22730 2573
rect 22744 2563 27434 2573
rect 8488 2539 14738 2549
rect 8536 2515 21170 2525
rect 21184 2515 24626 2525
rect 8584 2491 8594 2501
rect 8968 2491 17474 2501
rect 9064 2467 12002 2477
rect 12136 2467 26042 2477
rect 9352 2443 11066 2453
rect 11080 2443 23690 2453
rect 9520 2419 9554 2429
rect 9640 2419 22442 2429
rect 9592 2395 19106 2405
rect 19120 2395 20258 2405
rect 9712 2371 15146 2381
rect 9808 2347 20234 2357
rect 20248 2347 25226 2357
rect 25240 2347 25778 2357
rect 9832 2323 11498 2333
rect 11512 2323 11930 2333
rect 11944 2323 12362 2333
rect 12376 2323 14522 2333
rect 14536 2323 16562 2333
rect 16576 2323 22346 2333
rect 22360 2323 24194 2333
rect 24208 2323 26114 2333
rect 10048 2299 23738 2309
rect 10048 2275 13922 2285
rect 13936 2275 17114 2285
rect 10072 2251 10130 2261
rect 10216 2251 10802 2261
rect 10816 2251 12170 2261
rect 12184 2251 25826 2261
rect 10096 2227 22274 2237
rect 10456 2203 18842 2213
rect 18856 2203 21770 2213
rect 10720 2179 10730 2189
rect 10816 2179 12050 2189
rect 12064 2179 14642 2189
rect 14752 2179 22178 2189
rect 10936 2155 11114 2165
rect 11128 2155 23810 2165
rect 11008 2131 12962 2141
rect 13072 2131 20546 2141
rect 22192 2131 22778 2141
rect 11056 2107 11090 2117
rect 11176 2107 11978 2117
rect 12064 2107 19394 2117
rect 11080 2083 27506 2093
rect 11176 2059 21698 2069
rect 11440 2035 13250 2045
rect 13264 2035 13442 2045
rect 13456 2035 22106 2045
rect 11560 2011 16034 2021
rect 16048 2011 20354 2021
rect 11608 1987 24506 1997
rect 24520 1987 26522 1997
rect 11896 1963 15314 1973
rect 15328 1963 15890 1973
rect 17128 1963 21482 1973
rect 11968 1939 12194 1949
rect 12304 1939 24698 1949
rect 12208 1915 12386 1925
rect 12616 1915 23306 1925
rect 12424 1891 25970 1901
rect 12760 1867 12794 1877
rect 12880 1867 16778 1877
rect 16792 1867 23762 1877
rect 13000 1843 15362 1853
rect 15376 1843 16538 1853
rect 18856 1843 27266 1853
rect 13168 1819 22130 1829
rect 27640 1819 27963 1829
rect 13696 1795 13790 1805
rect 14320 1795 14618 1805
rect 15160 1795 21674 1805
rect 27616 1795 27963 1805
rect 14488 1771 14822 1781
rect 15904 1771 21722 1781
rect 21736 1771 22778 1781
rect 22792 1771 26930 1781
rect 27592 1771 27963 1781
rect 14536 1747 25322 1757
rect 27568 1747 27963 1757
rect 19408 1723 27074 1733
rect 27544 1723 27963 1733
rect 26979 1694 27531 1704
rect 26979 1671 27531 1681
rect 26979 1642 26985 1658
rect 27525 1642 27531 1658
rect 26979 1633 27531 1642
rect 26979 1004 27531 1013
rect 26979 988 26985 1004
rect 27525 988 27531 1004
rect 14056 890 14618 900
rect 16624 890 24554 900
rect 13984 866 20762 876
rect 20776 866 22370 876
rect 22384 866 22850 876
rect 22864 866 23810 876
rect 23824 866 24626 876
rect 24640 866 27026 876
rect 13792 842 18050 852
rect 13480 818 14066 828
rect 15184 818 22874 828
rect 13384 794 19034 804
rect 13216 770 23546 780
rect 12472 746 15938 756
rect 16480 746 22130 756
rect 12160 722 26810 732
rect 11272 698 22826 708
rect 10384 674 11354 684
rect 11824 674 14690 684
rect 14824 674 22586 684
rect 10360 650 11138 660
rect 11152 650 16346 660
rect 16360 650 27050 660
rect 10240 626 12650 636
rect 12712 626 14090 636
rect 14152 626 25970 636
rect 10120 602 17810 612
rect 22168 602 23642 612
rect 10096 578 15698 588
rect 16432 578 25730 588
rect 8824 554 11666 564
rect 11728 554 24506 564
rect 8800 530 20786 540
rect 21688 530 24986 540
rect 8440 506 19298 516
rect 20464 506 26762 516
rect 8296 482 24938 492
rect 8152 458 16874 468
rect 17416 458 20018 468
rect 20032 458 22226 468
rect 23296 458 24482 468
rect 25024 458 25130 468
rect 7792 434 15218 444
rect 17776 434 22250 444
rect 7432 410 16562 420
rect 7168 386 10754 396
rect 11224 386 20690 396
rect 7048 362 12506 372
rect 12568 362 18410 372
rect 6280 338 13826 348
rect 13840 338 20402 348
rect 20416 338 27002 348
rect 5032 314 5066 324
rect 5584 314 18986 324
rect 4792 290 10514 300
rect 10528 290 13346 300
rect 13360 290 14186 300
rect 14200 290 20546 300
rect 20560 290 22754 300
rect 22768 290 26978 300
rect 4504 266 22394 276
rect 4360 242 6578 252
rect 6856 242 24530 252
rect 4288 218 23426 228
rect 4240 194 19250 204
rect 4000 170 5162 180
rect 5224 170 6338 180
rect 6520 170 21650 180
rect 3616 146 13538 156
rect 13552 146 24314 156
rect 24328 146 27963 156
rect 2896 122 4034 132
rect 4048 122 9842 132
rect 9952 122 19058 132
rect 2848 98 14930 108
rect 27064 98 27963 108
rect 84 74 1778 84
rect 2728 74 14834 84
rect 27040 74 27963 84
rect 84 50 1730 60
rect 2488 50 11690 60
rect 11704 50 14210 60
rect 14224 50 18602 60
rect 18616 50 27963 60
rect 84 26 16130 36
rect 27016 26 27963 36
rect 84 2 26954 12
rect 26992 2 27963 12
<< m2contact >>
rect 16034 9010 16048 9024
rect 9890 8986 9904 9000
rect 16934 8986 16948 9000
rect 7274 8962 7288 8976
rect 18458 8962 18472 8976
rect 3938 8938 3952 8952
rect 4130 8938 4144 8952
rect 23030 8938 23044 8952
rect 2378 8914 2392 8928
rect 3242 8914 3256 8928
rect 27554 8914 27568 8928
rect 2042 8890 2056 8904
rect 24554 8890 24568 8904
rect 70 8866 84 8880
rect 22778 8866 22792 8880
rect 70 8842 84 8856
rect 20258 8842 20272 8856
rect 70 8818 84 8832
rect 11210 8818 11224 8832
rect 12314 8818 12328 8832
rect 17282 8818 17296 8832
rect 17522 8818 17536 8832
rect 26078 8818 26092 8832
rect 27506 8818 27520 8832
rect 27626 8818 27640 8832
rect 2210 8794 2224 8808
rect 13346 8794 13360 8808
rect 18698 8794 18712 8808
rect 27578 8794 27592 8808
rect 3674 8770 3688 8784
rect 27530 8770 27544 8784
rect 27578 8770 27592 8784
rect 27963 8770 27977 8784
rect 6170 8746 6184 8760
rect 17138 8746 17152 8760
rect 19226 8746 19240 8760
rect 19982 8746 19996 8760
rect 22730 8746 22744 8760
rect 25826 8746 25840 8760
rect 27578 8746 27592 8760
rect 27602 8746 27616 8760
rect 27963 8746 27977 8760
rect 7706 8722 7720 8736
rect 23354 8722 23368 8736
rect 27578 8722 27592 8736
rect 27963 8722 27977 8736
rect 9242 8698 9256 8712
rect 19178 8698 19192 8712
rect 27554 8698 27568 8712
rect 27963 8698 27977 8712
rect 9290 8674 9304 8688
rect 27602 8674 27616 8688
rect 27626 8674 27640 8688
rect 27963 8674 27977 8688
rect 10778 8650 10792 8664
rect 11714 8650 11728 8664
rect 12362 8650 12376 8664
rect 27963 8650 27977 8664
rect 13850 8626 13864 8640
rect 14834 8626 14848 8640
rect 15386 8626 15400 8640
rect 21098 8626 21112 8640
rect 27530 8626 27544 8640
rect 27963 8626 27977 8640
rect 13130 7793 13144 7807
rect 13346 7793 13360 7807
rect 13034 7769 13048 7783
rect 13274 7769 13288 7783
rect 13010 7745 13024 7759
rect 13202 7745 13216 7759
rect 13754 7745 13768 7759
rect 13922 7745 13936 7759
rect 20522 7745 20536 7759
rect 20762 7745 20776 7759
rect 20858 7745 20872 7759
rect 21146 7745 21160 7759
rect 12938 7721 12952 7735
rect 19274 7721 19288 7735
rect 19802 7721 19816 7735
rect 24146 7721 24160 7735
rect 12914 7697 12928 7711
rect 15218 7697 15232 7711
rect 18146 7697 18160 7711
rect 19874 7697 19888 7711
rect 20282 7697 20296 7711
rect 20522 7697 20536 7711
rect 20858 7697 20872 7711
rect 23402 7697 23416 7711
rect 12770 7673 12784 7687
rect 14450 7673 14464 7687
rect 24674 7673 24688 7687
rect 24986 7673 25000 7687
rect 11858 7649 11872 7663
rect 11930 7649 11944 7663
rect 12002 7649 12016 7663
rect 12266 7649 12280 7663
rect 12722 7649 12736 7663
rect 18074 7649 18088 7663
rect 23474 7649 23488 7663
rect 23522 7649 23536 7663
rect 24674 7649 24688 7663
rect 11810 7625 11824 7639
rect 12866 7625 12880 7639
rect 26762 7625 26776 7639
rect 11570 7601 11584 7615
rect 11618 7601 11632 7615
rect 11762 7601 11776 7615
rect 21086 7601 21100 7615
rect 11474 7577 11488 7591
rect 11546 7577 11560 7591
rect 11690 7577 11704 7591
rect 13778 7577 13792 7591
rect 11402 7553 11416 7567
rect 13850 7553 13864 7567
rect 11210 7529 11224 7543
rect 11282 7529 11296 7543
rect 23138 7529 23152 7543
rect 11066 7505 11080 7519
rect 27098 7505 27112 7519
rect 10994 7481 11008 7495
rect 23786 7481 23800 7495
rect 10586 7457 10600 7471
rect 11306 7457 11320 7471
rect 11378 7457 11392 7471
rect 22730 7457 22744 7471
rect 9986 7433 10000 7447
rect 10178 7433 10192 7447
rect 10322 7433 10336 7447
rect 25346 7433 25360 7447
rect 9962 7409 9976 7423
rect 14330 7409 14344 7423
rect 18482 7409 18496 7423
rect 9914 7385 9928 7399
rect 26954 7385 26968 7399
rect 9842 7361 9856 7375
rect 16874 7361 16888 7375
rect 9794 7337 9808 7351
rect 10346 7337 10360 7351
rect 13562 7337 13576 7351
rect 17354 7337 17368 7351
rect 19322 7337 19336 7351
rect 20330 7337 20344 7351
rect 21626 7337 21640 7351
rect 21698 7337 21712 7351
rect 9746 7313 9760 7327
rect 18266 7313 18280 7327
rect 26714 7313 26728 7327
rect 9746 7289 9760 7303
rect 9890 7289 9904 7303
rect 9938 7289 9952 7303
rect 14354 7289 14368 7303
rect 16946 7289 16960 7303
rect 21626 7289 21640 7303
rect 9434 7265 9448 7279
rect 13826 7265 13840 7279
rect 14618 7265 14632 7279
rect 9266 7241 9280 7255
rect 11090 7241 11104 7255
rect 15986 7241 16000 7255
rect 17714 7241 17728 7255
rect 24890 7241 24904 7255
rect 9194 7217 9208 7231
rect 18362 7217 18376 7231
rect 19634 7217 19648 7231
rect 20618 7217 20632 7231
rect 9146 7193 9160 7207
rect 17498 7193 17512 7207
rect 24218 7193 24232 7207
rect 24650 7193 24664 7207
rect 9002 7169 9016 7183
rect 22538 7169 22552 7183
rect 24218 7169 24232 7183
rect 8714 7145 8728 7159
rect 8738 7145 8752 7159
rect 8834 7145 8848 7159
rect 10970 7145 10984 7159
rect 11018 7145 11032 7159
rect 11066 7145 11080 7159
rect 11114 7145 11128 7159
rect 21578 7145 21592 7159
rect 8594 7121 8608 7135
rect 21122 7121 21136 7135
rect 8522 7097 8536 7111
rect 14762 7097 14776 7111
rect 8498 7073 8512 7087
rect 9362 7073 9376 7087
rect 17930 7073 17944 7087
rect 22466 7073 22480 7087
rect 23690 7073 23704 7087
rect 8450 7049 8464 7063
rect 10874 7049 10888 7063
rect 12218 7049 12232 7063
rect 15074 7049 15088 7063
rect 8258 7025 8272 7039
rect 14714 7025 14728 7039
rect 17954 7025 17968 7039
rect 19538 7025 19552 7039
rect 7946 7001 7960 7015
rect 17954 7001 17968 7015
rect 7850 6977 7864 6991
rect 10778 6977 10792 6991
rect 14066 6977 14080 6991
rect 7634 6953 7648 6967
rect 13754 6953 13768 6967
rect 7586 6929 7600 6943
rect 12074 6929 12088 6943
rect 13634 6929 13648 6943
rect 17570 6929 17584 6943
rect 7538 6905 7552 6919
rect 9242 6905 9256 6919
rect 9410 6905 9424 6919
rect 12842 6905 12856 6919
rect 13490 6905 13504 6919
rect 13826 6905 13840 6919
rect 27026 6905 27040 6919
rect 7490 6881 7504 6895
rect 8786 6881 8800 6895
rect 25922 6881 25936 6895
rect 7418 6857 7432 6871
rect 8090 6857 8104 6871
rect 8162 6857 8176 6871
rect 8282 6857 8296 6871
rect 8354 6857 8368 6871
rect 19610 6857 19624 6871
rect 7370 6833 7384 6847
rect 12482 6833 12496 6847
rect 12578 6833 12592 6847
rect 21938 6833 21952 6847
rect 7346 6809 7360 6823
rect 8186 6809 8200 6823
rect 8234 6809 8248 6823
rect 27626 6809 27640 6823
rect 7322 6785 7336 6799
rect 26138 6785 26152 6799
rect 7250 6761 7264 6775
rect 19346 6761 19360 6775
rect 7058 6737 7072 6751
rect 13010 6737 13024 6751
rect 16586 6737 16600 6751
rect 7058 6713 7072 6727
rect 23282 6713 23296 6727
rect 7034 6689 7048 6703
rect 15842 6689 15856 6703
rect 7010 6665 7024 6679
rect 7034 6665 7048 6679
rect 7130 6665 7144 6679
rect 12914 6665 12928 6679
rect 23234 6665 23248 6679
rect 6938 6641 6952 6655
rect 16250 6641 16264 6655
rect 25706 6641 25720 6655
rect 6650 6617 6664 6631
rect 23954 6617 23968 6631
rect 6506 6593 6520 6607
rect 25730 6593 25744 6607
rect 6482 6569 6496 6583
rect 21986 6569 22000 6583
rect 6434 6545 6448 6559
rect 20978 6545 20992 6559
rect 6410 6521 6424 6535
rect 16754 6521 16768 6535
rect 17234 6521 17248 6535
rect 17306 6521 17320 6535
rect 18914 6521 18928 6535
rect 20642 6521 20656 6535
rect 6362 6497 6376 6511
rect 6914 6497 6928 6511
rect 6962 6497 6976 6511
rect 18890 6497 18904 6511
rect 6338 6473 6352 6487
rect 17210 6473 17224 6487
rect 20618 6473 20632 6487
rect 6290 6449 6304 6463
rect 14258 6449 14272 6463
rect 16202 6449 16216 6463
rect 19562 6449 19576 6463
rect 6266 6425 6280 6439
rect 11834 6425 11848 6439
rect 13514 6425 13528 6439
rect 17234 6425 17248 6439
rect 25682 6425 25696 6439
rect 26786 6425 26800 6439
rect 6194 6401 6208 6415
rect 18314 6401 18328 6415
rect 18914 6401 18928 6415
rect 19010 6401 19024 6415
rect 25082 6401 25096 6415
rect 6050 6377 6064 6391
rect 20114 6377 20128 6391
rect 23498 6377 23512 6391
rect 23810 6377 23824 6391
rect 5954 6353 5968 6367
rect 13946 6353 13960 6367
rect 18290 6353 18304 6367
rect 24026 6353 24040 6367
rect 5906 6329 5920 6343
rect 6434 6329 6448 6343
rect 8066 6329 8080 6343
rect 14234 6329 14248 6343
rect 18002 6329 18016 6343
rect 24122 6329 24136 6343
rect 5546 6305 5560 6319
rect 7706 6305 7720 6319
rect 14954 6305 14968 6319
rect 26642 6305 26656 6319
rect 5546 6281 5560 6295
rect 10634 6281 10648 6295
rect 10946 6281 10960 6295
rect 17258 6281 17272 6295
rect 17450 6281 17464 6295
rect 24962 6281 24976 6295
rect 5498 6257 5512 6271
rect 12194 6257 12208 6271
rect 12290 6257 12304 6271
rect 13790 6257 13804 6271
rect 17426 6257 17440 6271
rect 21578 6257 21592 6271
rect 25370 6257 25384 6271
rect 5474 6233 5488 6247
rect 8138 6233 8152 6247
rect 19898 6233 19912 6247
rect 21530 6233 21544 6247
rect 26354 6233 26368 6247
rect 5450 6209 5464 6223
rect 10322 6209 10336 6223
rect 19202 6209 19216 6223
rect 19298 6209 19312 6223
rect 21530 6209 21544 6223
rect 23498 6209 23512 6223
rect 5450 6185 5464 6199
rect 27218 6185 27232 6199
rect 5426 6161 5440 6175
rect 14114 6161 14128 6175
rect 15338 6161 15352 6175
rect 15386 6161 15400 6175
rect 17378 6161 17392 6175
rect 20426 6161 20440 6175
rect 20498 6161 20512 6175
rect 20546 6161 20560 6175
rect 5402 6137 5416 6151
rect 24794 6137 24808 6151
rect 5354 6113 5368 6127
rect 9650 6113 9664 6127
rect 9722 6113 9736 6127
rect 17138 6113 17152 6127
rect 21050 6113 21064 6127
rect 23714 6113 23728 6127
rect 25058 6113 25072 6127
rect 26570 6113 26584 6127
rect 5354 6089 5368 6103
rect 16154 6089 16168 6103
rect 17066 6089 17080 6103
rect 23450 6089 23464 6103
rect 5330 6065 5344 6079
rect 21266 6065 21280 6079
rect 5306 6041 5320 6055
rect 25274 6041 25288 6055
rect 5258 6017 5272 6031
rect 19346 6017 19360 6031
rect 24410 6017 24424 6031
rect 5258 5993 5272 6007
rect 16994 5993 17008 6007
rect 17042 5993 17056 6007
rect 26474 5993 26488 6007
rect 5066 5969 5080 5983
rect 26882 5969 26896 5983
rect 5018 5945 5032 5959
rect 10418 5945 10432 5959
rect 20498 5945 20512 5959
rect 4970 5921 4984 5935
rect 15338 5921 15352 5935
rect 16034 5921 16048 5935
rect 26618 5921 26632 5935
rect 4922 5897 4936 5911
rect 24530 5897 24544 5911
rect 4874 5873 4888 5887
rect 19658 5873 19672 5887
rect 4850 5849 4864 5863
rect 5042 5849 5056 5863
rect 9386 5849 9400 5863
rect 9554 5849 9568 5863
rect 10562 5849 10576 5863
rect 11882 5849 11896 5863
rect 13130 5849 13144 5863
rect 20594 5849 20608 5863
rect 22970 5849 22984 5863
rect 23258 5849 23272 5863
rect 26810 5849 26824 5863
rect 4778 5825 4792 5839
rect 4946 5825 4960 5839
rect 6674 5825 6688 5839
rect 25898 5825 25912 5839
rect 4754 5801 4768 5815
rect 9026 5801 9040 5815
rect 10634 5801 10648 5815
rect 11474 5801 11488 5815
rect 16442 5801 16456 5815
rect 16970 5801 16984 5815
rect 24314 5801 24328 5815
rect 4730 5777 4744 5791
rect 8594 5777 8608 5791
rect 9986 5777 10000 5791
rect 21722 5777 21736 5791
rect 4610 5753 4624 5767
rect 5570 5753 5584 5767
rect 21890 5753 21904 5767
rect 4586 5729 4600 5743
rect 7106 5729 7120 5743
rect 7178 5729 7192 5743
rect 25778 5729 25792 5743
rect 4562 5705 4576 5719
rect 20930 5705 20944 5719
rect 4514 5681 4528 5695
rect 19586 5681 19600 5695
rect 26906 5681 26920 5695
rect 27074 5681 27088 5695
rect 4418 5657 4432 5671
rect 26906 5657 26920 5671
rect 4370 5633 4384 5647
rect 20906 5633 20920 5647
rect 4346 5609 4360 5623
rect 11690 5609 11704 5623
rect 15242 5609 15256 5623
rect 23618 5609 23632 5623
rect 4202 5585 4216 5599
rect 7322 5585 7336 5599
rect 13082 5585 13096 5599
rect 23378 5585 23392 5599
rect 4082 5561 4096 5575
rect 11330 5561 11344 5575
rect 15050 5561 15064 5575
rect 15266 5561 15280 5575
rect 19010 5561 19024 5575
rect 4082 5537 4096 5551
rect 25010 5537 25024 5551
rect 4034 5513 4048 5527
rect 5882 5513 5896 5527
rect 23042 5513 23056 5527
rect 23858 5513 23872 5527
rect 23882 5513 23896 5527
rect 4010 5489 4024 5503
rect 6842 5489 6856 5503
rect 10610 5489 10624 5503
rect 16322 5489 16336 5503
rect 18290 5489 18304 5503
rect 20834 5489 20848 5503
rect 23162 5489 23176 5503
rect 23642 5489 23656 5503
rect 24098 5489 24112 5503
rect 24386 5489 24400 5503
rect 26882 5489 26896 5503
rect 27554 5489 27568 5503
rect 3986 5465 4000 5479
rect 6290 5465 6304 5479
rect 7994 5465 8008 5479
rect 8474 5465 8488 5479
rect 17186 5465 17200 5479
rect 23858 5465 23872 5479
rect 3938 5441 3952 5455
rect 6650 5441 6664 5455
rect 6722 5441 6736 5455
rect 7730 5441 7744 5455
rect 7826 5441 7840 5455
rect 7850 5441 7864 5455
rect 7922 5441 7936 5455
rect 7946 5441 7960 5455
rect 7994 5441 8008 5455
rect 8066 5441 8080 5455
rect 8114 5441 8128 5455
rect 10730 5441 10744 5455
rect 10898 5441 10912 5455
rect 13322 5441 13336 5455
rect 23090 5441 23104 5455
rect 3866 5417 3880 5431
rect 13994 5417 14008 5431
rect 15098 5417 15112 5431
rect 20762 5417 20776 5431
rect 3866 5393 3880 5407
rect 19682 5393 19696 5407
rect 3842 5369 3856 5383
rect 4226 5369 4240 5383
rect 7298 5369 7312 5383
rect 7634 5369 7648 5383
rect 7802 5369 7816 5383
rect 8114 5369 8128 5383
rect 8570 5369 8584 5383
rect 14282 5369 14296 5383
rect 16514 5369 16528 5383
rect 16946 5369 16960 5383
rect 23930 5369 23944 5383
rect 24362 5369 24376 5383
rect 3842 5345 3856 5359
rect 6554 5345 6568 5359
rect 6698 5345 6712 5359
rect 10538 5345 10552 5359
rect 14114 5345 14128 5359
rect 18146 5345 18160 5359
rect 3794 5321 3808 5335
rect 7394 5321 7408 5335
rect 7466 5321 7480 5335
rect 19082 5321 19096 5335
rect 20186 5321 20200 5335
rect 20258 5321 20272 5335
rect 3770 5297 3784 5311
rect 7682 5297 7696 5311
rect 26234 5297 26248 5311
rect 3770 5273 3784 5287
rect 6122 5273 6136 5287
rect 6170 5273 6184 5287
rect 17090 5273 17104 5287
rect 18122 5273 18136 5287
rect 20090 5273 20104 5287
rect 27578 5273 27592 5287
rect 3722 5249 3736 5263
rect 12314 5249 12328 5263
rect 12362 5249 12376 5263
rect 12386 5249 12400 5263
rect 12554 5249 12568 5263
rect 13178 5249 13192 5263
rect 14786 5249 14800 5263
rect 24770 5249 24784 5263
rect 3626 5225 3640 5239
rect 14018 5225 14032 5239
rect 17690 5225 17704 5239
rect 17738 5225 17752 5239
rect 27963 5225 27977 5239
rect 3578 5201 3592 5215
rect 20210 5201 20224 5215
rect 22034 5201 22048 5215
rect 22130 5201 22144 5215
rect 3530 5177 3544 5191
rect 11642 5177 11656 5191
rect 11714 5177 11728 5191
rect 15098 5177 15112 5191
rect 15194 5177 15208 5191
rect 22058 5177 22072 5191
rect 3506 5153 3520 5167
rect 5738 5153 5752 5167
rect 5834 5153 5848 5167
rect 17978 5153 17992 5167
rect 21290 5153 21304 5167
rect 25562 5153 25576 5167
rect 25706 5153 25720 5167
rect 3410 5129 3424 5143
rect 25850 5129 25864 5143
rect 3386 5105 3400 5119
rect 25634 5105 25648 5119
rect 3314 5081 3328 5095
rect 7922 5081 7936 5095
rect 8450 5081 8464 5095
rect 9482 5081 9496 5095
rect 11042 5081 11056 5095
rect 18986 5081 19000 5095
rect 20018 5081 20032 5095
rect 20234 5081 20248 5095
rect 20306 5081 20320 5095
rect 20354 5081 20368 5095
rect 20450 5081 20464 5095
rect 20738 5081 20752 5095
rect 21002 5081 21016 5095
rect 26738 5081 26752 5095
rect 3218 5057 3232 5071
rect 6554 5057 6568 5071
rect 11018 5057 11032 5071
rect 19922 5057 19936 5071
rect 21002 5057 21016 5071
rect 22010 5057 22024 5071
rect 27458 5057 27472 5071
rect 3146 5033 3160 5047
rect 19058 5033 19072 5047
rect 22826 5033 22840 5047
rect 3098 5009 3112 5023
rect 4178 5009 4192 5023
rect 17018 5009 17032 5023
rect 17786 5009 17800 5023
rect 26306 5009 26320 5023
rect 3050 4985 3064 4999
rect 27146 4985 27160 4999
rect 3002 4961 3016 4975
rect 3914 4961 3928 4975
rect 13034 4961 13048 4975
rect 14690 4961 14704 4975
rect 24458 4961 24472 4975
rect 25682 4961 25696 4975
rect 2954 4937 2968 4951
rect 16826 4937 16840 4951
rect 21374 4937 21388 4951
rect 24338 4937 24352 4951
rect 2930 4913 2944 4927
rect 27122 4913 27136 4927
rect 2906 4889 2920 4903
rect 20474 4889 20488 4903
rect 21866 4889 21880 4903
rect 22106 4889 22120 4903
rect 22946 4889 22960 4903
rect 23210 4889 23224 4903
rect 23534 4889 23548 4903
rect 2786 4865 2800 4879
rect 24002 4865 24016 4879
rect 2738 4841 2752 4855
rect 8210 4841 8224 4855
rect 20066 4841 20080 4855
rect 20378 4841 20392 4855
rect 22034 4841 22048 4855
rect 22850 4841 22864 4855
rect 23186 4841 23200 4855
rect 23330 4841 23344 4855
rect 23654 4841 23668 4855
rect 2666 4817 2680 4831
rect 4826 4817 4840 4831
rect 7010 4817 7024 4831
rect 10418 4817 10432 4831
rect 10466 4817 10480 4831
rect 13730 4817 13744 4831
rect 13970 4817 13984 4831
rect 21242 4817 21256 4831
rect 23594 4817 23608 4831
rect 24242 4817 24256 4831
rect 24290 4817 24304 4831
rect 24542 4817 24556 4831
rect 24602 4817 24616 4831
rect 24806 4817 24820 4831
rect 25490 4817 25504 4831
rect 25610 4817 25624 4831
rect 25802 4817 25816 4831
rect 25826 4817 25840 4831
rect 25874 4817 25888 4831
rect 26978 4817 26992 4831
rect 2522 4793 2536 4807
rect 6602 4793 6616 4807
rect 16106 4793 16120 4807
rect 19706 4793 19720 4807
rect 24722 4793 24736 4807
rect 27314 4793 27328 4807
rect 2450 4769 2464 4783
rect 8666 4769 8680 4783
rect 9338 4769 9352 4783
rect 13970 4769 13984 4783
rect 14426 4769 14440 4783
rect 14570 4769 14584 4783
rect 17594 4769 17608 4783
rect 26690 4769 26704 4783
rect 26954 4769 26968 4783
rect 27338 4769 27352 4783
rect 2426 4745 2440 4759
rect 14930 4745 14944 4759
rect 24290 4745 24304 4759
rect 24962 4745 24976 4759
rect 25082 4745 25096 4759
rect 26642 4745 26656 4759
rect 26714 4745 26728 4759
rect 2330 4721 2344 4735
rect 23738 4721 23752 4735
rect 24002 4721 24016 4735
rect 26426 4721 26440 4735
rect 26690 4721 26704 4735
rect 26978 4721 26992 4735
rect 2306 4697 2320 4711
rect 2450 4697 2464 4711
rect 4538 4697 4552 4711
rect 4970 4697 4984 4711
rect 8258 4697 8272 4711
rect 10658 4697 10672 4711
rect 10706 4697 10720 4711
rect 12626 4697 12640 4711
rect 14378 4697 14392 4711
rect 14546 4697 14560 4711
rect 18026 4697 18040 4711
rect 20186 4697 20200 4711
rect 25538 4697 25552 4711
rect 2282 4673 2296 4687
rect 11906 4673 11920 4687
rect 12026 4673 12040 4687
rect 21770 4673 21784 4687
rect 22058 4673 22072 4687
rect 27602 4673 27616 4687
rect 2234 4649 2248 4663
rect 23978 4649 23992 4663
rect 2186 4625 2200 4639
rect 7826 4625 7840 4639
rect 11762 4625 11776 4639
rect 11858 4625 11872 4639
rect 23018 4625 23032 4639
rect 2138 4601 2152 4615
rect 21410 4601 21424 4615
rect 2114 4577 2128 4591
rect 5498 4577 5512 4591
rect 19130 4577 19144 4591
rect 23906 4577 23920 4591
rect 23954 4577 23968 4591
rect 24938 4577 24952 4591
rect 25442 4577 25456 4591
rect 1994 4553 2008 4567
rect 10298 4553 10312 4567
rect 18194 4553 18208 4567
rect 18530 4553 18544 4567
rect 24542 4553 24556 4567
rect 1970 4529 1984 4543
rect 9098 4529 9112 4543
rect 18962 4529 18976 4543
rect 21338 4529 21352 4543
rect 23906 4529 23920 4543
rect 24146 4529 24160 4543
rect 1922 4505 1936 4519
rect 15482 4505 15496 4519
rect 15746 4505 15760 4519
rect 24482 4505 24496 4519
rect 1898 4481 1912 4495
rect 22082 4481 22096 4495
rect 1898 4457 1912 4471
rect 24842 4457 24856 4471
rect 1850 4433 1864 4447
rect 2570 4433 2584 4447
rect 2618 4433 2632 4447
rect 8042 4433 8056 4447
rect 9218 4433 9232 4447
rect 17066 4433 17080 4447
rect 17162 4433 17176 4447
rect 17282 4433 17296 4447
rect 18722 4433 18736 4447
rect 25514 4433 25528 4447
rect 1802 4409 1816 4423
rect 7442 4409 7456 4423
rect 10154 4409 10168 4423
rect 10874 4409 10888 4423
rect 20786 4409 20800 4423
rect 20882 4409 20896 4423
rect 20978 4409 20992 4423
rect 21086 4409 21100 4423
rect 21338 4409 21352 4423
rect 21374 4409 21388 4423
rect 1778 4385 1792 4399
rect 6626 4385 6640 4399
rect 6746 4385 6760 4399
rect 12530 4385 12544 4399
rect 13274 4385 13288 4399
rect 19754 4385 19768 4399
rect 20906 4385 20920 4399
rect 24986 4385 25000 4399
rect 1754 4361 1768 4375
rect 3602 4361 3616 4375
rect 9818 4361 9832 4375
rect 12458 4361 12472 4375
rect 20666 4361 20680 4375
rect 1730 4337 1744 4351
rect 4418 4337 4432 4351
rect 5138 4337 5152 4351
rect 14882 4337 14896 4351
rect 20714 4337 20728 4351
rect 27530 4337 27544 4351
rect 1658 4313 1672 4327
rect 19274 4313 19288 4327
rect 1658 4289 1672 4303
rect 4250 4289 4264 4303
rect 4322 4289 4336 4303
rect 5690 4289 5704 4303
rect 8714 4289 8728 4303
rect 12434 4289 12448 4303
rect 16730 4289 16744 4303
rect 20378 4289 20392 4303
rect 1634 4265 1648 4279
rect 19442 4265 19456 4279
rect 1610 4241 1624 4255
rect 3074 4241 3088 4255
rect 3290 4241 3304 4255
rect 5786 4241 5800 4255
rect 13418 4241 13432 4255
rect 14594 4241 14608 4255
rect 22634 4241 22648 4255
rect 24578 4241 24592 4255
rect 70 4217 84 4231
rect 1682 4217 1696 4231
rect 1730 4217 1744 4231
rect 2546 4217 2560 4231
rect 2618 4217 2632 4231
rect 4442 4217 4456 4231
rect 6698 4217 6712 4231
rect 7130 4217 7144 4231
rect 11978 4217 11992 4231
rect 14210 4217 14224 4231
rect 20834 4217 20848 4231
rect 21074 4217 21088 4231
rect 21650 4217 21664 4231
rect 24602 4217 24616 4231
rect 70 4193 84 4207
rect 14882 4193 14896 4207
rect 15050 4193 15064 4207
rect 15074 4193 15088 4207
rect 15914 4193 15928 4207
rect 16706 4193 16720 4207
rect 22994 4193 23008 4207
rect 70 4169 84 4183
rect 8306 4169 8320 4183
rect 8354 4169 8368 4183
rect 26834 4169 26848 4183
rect 70 4145 84 4159
rect 25394 4145 25408 4159
rect 1610 4121 1624 4135
rect 3458 4121 3472 4135
rect 14810 4121 14824 4135
rect 14858 4121 14872 4135
rect 17834 4121 17848 4135
rect 18770 4121 18784 4135
rect 19226 4121 19240 4135
rect 1874 4097 1888 4111
rect 11906 4097 11920 4111
rect 12098 4097 12112 4111
rect 13706 4097 13720 4111
rect 14234 4097 14248 4111
rect 14258 4097 14272 4111
rect 14786 4097 14800 4111
rect 21554 4097 21568 4111
rect 22682 4097 22696 4111
rect 2090 4073 2104 4087
rect 14978 4073 14992 4087
rect 16514 4073 16528 4087
rect 16586 4073 16600 4087
rect 16658 4073 16672 4087
rect 20954 4073 20968 4087
rect 2258 4049 2272 4063
rect 4994 4049 5008 4063
rect 11594 4049 11608 4063
rect 19466 4049 19480 4063
rect 21218 4049 21232 4063
rect 21818 4049 21832 4063
rect 2306 4025 2320 4039
rect 3746 4025 3760 4039
rect 7658 4025 7672 4039
rect 9122 4025 9136 4039
rect 10298 4025 10312 4039
rect 10514 4025 10528 4039
rect 17906 4025 17920 4039
rect 22658 4025 22672 4039
rect 23330 4025 23344 4039
rect 23618 4025 23632 4039
rect 2378 4001 2392 4015
rect 21026 4001 21040 4015
rect 2474 3977 2488 3991
rect 8162 3977 8176 3991
rect 8234 3977 8248 3991
rect 9530 3977 9544 3991
rect 9602 3977 9616 3991
rect 16898 3977 16912 3991
rect 20738 3977 20752 3991
rect 2498 3953 2512 3967
rect 16826 3953 16840 3967
rect 26090 3953 26104 3967
rect 2546 3929 2560 3943
rect 9530 3929 9544 3943
rect 12482 3929 12496 3943
rect 12650 3929 12664 3943
rect 14402 3929 14416 3943
rect 21938 3929 21952 3943
rect 2570 3905 2584 3919
rect 8018 3905 8032 3919
rect 16754 3905 16768 3919
rect 18650 3905 18664 3919
rect 18866 3905 18880 3919
rect 21866 3905 21880 3919
rect 26186 3905 26200 3919
rect 27002 3905 27016 3919
rect 2666 3881 2680 3895
rect 10274 3881 10288 3895
rect 18002 3881 18016 3895
rect 18938 3881 18952 3895
rect 19178 3881 19192 3895
rect 2762 3857 2776 3871
rect 27963 3857 27977 3871
rect 2786 3833 2800 3847
rect 7898 3833 7912 3847
rect 23570 3833 23584 3847
rect 24842 3833 24856 3847
rect 24914 3833 24928 3847
rect 2810 3809 2824 3823
rect 3962 3809 3976 3823
rect 4394 3809 4408 3823
rect 11258 3809 11272 3823
rect 11570 3809 11584 3823
rect 12170 3809 12184 3823
rect 13610 3809 13624 3823
rect 22946 3809 22960 3823
rect 23402 3809 23416 3823
rect 26210 3809 26224 3823
rect 2834 3785 2848 3799
rect 7466 3785 7480 3799
rect 7514 3785 7528 3799
rect 12794 3785 12808 3799
rect 13202 3785 13216 3799
rect 13226 3785 13240 3799
rect 14426 3785 14440 3799
rect 23834 3785 23848 3799
rect 2858 3761 2872 3775
rect 22970 3761 22984 3775
rect 2906 3737 2920 3751
rect 3458 3737 3472 3751
rect 10682 3737 10696 3751
rect 19970 3737 19984 3751
rect 23114 3737 23128 3751
rect 24806 3737 24820 3751
rect 25034 3737 25048 3751
rect 25802 3737 25816 3751
rect 3194 3713 3208 3727
rect 24122 3713 24136 3727
rect 3338 3689 3352 3703
rect 5282 3689 5296 3703
rect 5330 3689 5344 3703
rect 11522 3689 11536 3703
rect 12098 3689 12112 3703
rect 12146 3689 12160 3703
rect 21362 3689 21376 3703
rect 3410 3665 3424 3679
rect 5810 3665 5824 3679
rect 7946 3665 7960 3679
rect 9506 3665 9520 3679
rect 11618 3665 11632 3679
rect 14402 3665 14416 3679
rect 14594 3665 14608 3679
rect 14666 3665 14680 3679
rect 16970 3665 16984 3679
rect 24266 3665 24280 3679
rect 25250 3665 25264 3679
rect 26546 3665 26560 3679
rect 3650 3641 3664 3655
rect 4682 3641 4696 3655
rect 5114 3641 5128 3655
rect 13946 3641 13960 3655
rect 22322 3641 22336 3655
rect 3746 3617 3760 3631
rect 7106 3617 7120 3631
rect 7610 3617 7624 3631
rect 10850 3617 10864 3631
rect 19154 3617 19168 3631
rect 23354 3617 23368 3631
rect 24434 3617 24448 3631
rect 26666 3617 26680 3631
rect 3818 3593 3832 3607
rect 3938 3593 3952 3607
rect 6818 3593 6832 3607
rect 8330 3593 8344 3607
rect 9890 3593 9904 3607
rect 12242 3593 12256 3607
rect 21458 3593 21472 3607
rect 23786 3593 23800 3607
rect 24434 3593 24448 3607
rect 27194 3593 27208 3607
rect 3890 3569 3904 3583
rect 8762 3569 8776 3583
rect 8906 3569 8920 3583
rect 14822 3569 14836 3583
rect 26594 3569 26608 3583
rect 4154 3545 4168 3559
rect 4658 3545 4672 3559
rect 9698 3545 9712 3559
rect 10274 3545 10288 3559
rect 13658 3545 13672 3559
rect 17810 3545 17824 3559
rect 21554 3545 21568 3559
rect 23426 3545 23440 3559
rect 26594 3545 26608 3559
rect 26618 3545 26632 3559
rect 4202 3521 4216 3535
rect 4298 3521 4312 3535
rect 8930 3521 8944 3535
rect 12746 3521 12760 3535
rect 13154 3521 13168 3535
rect 13466 3521 13480 3535
rect 19370 3521 19384 3535
rect 23534 3521 23548 3535
rect 26330 3521 26344 3535
rect 4298 3497 4312 3511
rect 21962 3497 21976 3511
rect 4442 3473 4456 3487
rect 12410 3473 12424 3487
rect 25106 3473 25120 3487
rect 4466 3449 4480 3463
rect 6482 3449 6496 3463
rect 6530 3449 6544 3463
rect 10370 3449 10384 3463
rect 27050 3449 27064 3463
rect 4514 3425 4528 3439
rect 18050 3425 18064 3439
rect 4538 3401 4552 3415
rect 8282 3401 8296 3415
rect 8378 3401 8392 3415
rect 21434 3401 21448 3415
rect 4562 3377 4576 3391
rect 12338 3377 12352 3391
rect 12674 3377 12688 3391
rect 20162 3377 20176 3391
rect 4634 3353 4648 3367
rect 13514 3353 13528 3367
rect 25154 3353 25168 3367
rect 4658 3329 4672 3343
rect 6938 3329 6952 3343
rect 15002 3329 15016 3343
rect 15122 3329 15136 3343
rect 17090 3329 17104 3343
rect 17258 3329 17272 3343
rect 4706 3305 4720 3319
rect 7226 3305 7240 3319
rect 26546 3305 26560 3319
rect 4754 3281 4768 3295
rect 6722 3281 6736 3295
rect 8666 3281 8680 3295
rect 8738 3281 8752 3295
rect 12578 3281 12592 3295
rect 12818 3281 12832 3295
rect 13106 3281 13120 3295
rect 17882 3281 17896 3295
rect 21962 3281 21976 3295
rect 4802 3257 4816 3271
rect 5210 3257 5224 3271
rect 19514 3257 19528 3271
rect 4850 3233 4864 3247
rect 11786 3233 11800 3247
rect 20690 3233 20704 3247
rect 22586 3233 22600 3247
rect 4874 3209 4888 3223
rect 5162 3209 5176 3223
rect 16850 3209 16864 3223
rect 21314 3209 21328 3223
rect 22922 3209 22936 3223
rect 4922 3185 4936 3199
rect 17330 3185 17344 3199
rect 5090 3161 5104 3175
rect 9602 3161 9616 3175
rect 11138 3161 11152 3175
rect 19994 3161 20008 3175
rect 21842 3161 21856 3175
rect 22562 3161 22576 3175
rect 23882 3161 23896 3175
rect 26330 3161 26344 3175
rect 5114 3137 5128 3151
rect 6386 3137 6400 3151
rect 6458 3137 6472 3151
rect 7802 3137 7816 3151
rect 13898 3137 13912 3151
rect 14282 3137 14296 3151
rect 14450 3137 14464 3151
rect 14666 3137 14680 3151
rect 27362 3137 27376 3151
rect 5186 3113 5200 3127
rect 6866 3113 6880 3127
rect 18098 3113 18112 3127
rect 5402 3089 5416 3103
rect 11954 3089 11968 3103
rect 13298 3089 13312 3103
rect 13586 3089 13600 3103
rect 14186 3089 14200 3103
rect 15026 3089 15040 3103
rect 23522 3089 23536 3103
rect 27410 3089 27424 3103
rect 5522 3065 5536 3079
rect 5618 3065 5632 3079
rect 25466 3065 25480 3079
rect 26522 3065 26536 3079
rect 5666 3041 5680 3055
rect 22490 3041 22504 3055
rect 5690 3017 5704 3031
rect 6074 3017 6088 3031
rect 6146 3017 6160 3031
rect 20330 3017 20344 3031
rect 6002 2993 6016 3007
rect 16154 2993 16168 3007
rect 17210 2993 17224 3007
rect 21410 2993 21424 3007
rect 24650 2993 24664 3007
rect 6026 2969 6040 2983
rect 23066 2969 23080 2983
rect 6050 2945 6064 2959
rect 15386 2945 15400 2959
rect 17282 2945 17296 2959
rect 20570 2945 20584 2959
rect 24386 2945 24400 2959
rect 6098 2921 6112 2935
rect 7034 2921 7048 2935
rect 23042 2921 23056 2935
rect 6218 2897 6232 2911
rect 24050 2897 24064 2911
rect 6602 2873 6616 2887
rect 18866 2873 18880 2887
rect 20954 2873 20968 2887
rect 24746 2873 24760 2887
rect 6626 2849 6640 2863
rect 6674 2849 6688 2863
rect 6770 2849 6784 2863
rect 25994 2849 26008 2863
rect 6794 2825 6808 2839
rect 7538 2825 7552 2839
rect 9578 2825 9592 2839
rect 10490 2825 10504 2839
rect 11642 2825 11656 2839
rect 12674 2825 12688 2839
rect 14498 2825 14512 2839
rect 19442 2825 19456 2839
rect 21194 2825 21208 2839
rect 21746 2825 21760 2839
rect 24074 2825 24088 2839
rect 25586 2825 25600 2839
rect 26378 2825 26392 2839
rect 6818 2801 6832 2815
rect 8642 2801 8656 2815
rect 14306 2801 14320 2815
rect 25490 2801 25504 2815
rect 6890 2777 6904 2791
rect 15026 2777 15040 2791
rect 17306 2777 17320 2791
rect 18098 2777 18112 2791
rect 18122 2777 18136 2791
rect 20570 2777 20584 2791
rect 23654 2777 23668 2791
rect 24074 2777 24088 2791
rect 24242 2777 24256 2791
rect 7202 2753 7216 2767
rect 17642 2753 17656 2767
rect 21914 2753 21928 2767
rect 7226 2729 7240 2743
rect 7850 2729 7864 2743
rect 11354 2729 11368 2743
rect 12266 2729 12280 2743
rect 13346 2729 13360 2743
rect 14474 2729 14488 2743
rect 20306 2729 20320 2743
rect 21842 2729 21856 2743
rect 26282 2729 26296 2743
rect 7250 2705 7264 2719
rect 26402 2705 26416 2719
rect 7346 2681 7360 2695
rect 16370 2681 16384 2695
rect 23978 2681 23992 2695
rect 25610 2681 25624 2695
rect 7370 2657 7384 2671
rect 13682 2657 13696 2671
rect 13730 2657 13744 2671
rect 21146 2657 21160 2671
rect 21194 2657 21208 2671
rect 22898 2657 22912 2671
rect 7682 2633 7696 2647
rect 7706 2633 7720 2647
rect 7754 2633 7768 2647
rect 9674 2633 9688 2647
rect 12818 2633 12832 2647
rect 20810 2633 20824 2647
rect 24170 2633 24184 2647
rect 24866 2633 24880 2647
rect 7730 2609 7744 2623
rect 8618 2609 8632 2623
rect 8930 2609 8944 2623
rect 10106 2609 10120 2623
rect 10202 2609 10216 2623
rect 26858 2609 26872 2623
rect 7874 2585 7888 2599
rect 10010 2585 10024 2599
rect 11546 2585 11560 2599
rect 12770 2585 12784 2599
rect 19490 2585 19504 2599
rect 20162 2585 20176 2599
rect 24170 2585 24184 2599
rect 24458 2585 24472 2599
rect 8042 2561 8056 2575
rect 8138 2561 8152 2575
rect 8426 2561 8440 2575
rect 9482 2561 9496 2575
rect 10922 2561 10936 2575
rect 13874 2561 13888 2575
rect 22730 2561 22744 2575
rect 27434 2561 27448 2575
rect 8474 2537 8488 2551
rect 14738 2537 14752 2551
rect 8522 2513 8536 2527
rect 21170 2513 21184 2527
rect 24626 2513 24640 2527
rect 8570 2489 8584 2503
rect 8594 2489 8608 2503
rect 8954 2489 8968 2503
rect 17474 2489 17488 2503
rect 9050 2465 9064 2479
rect 12002 2465 12016 2479
rect 12122 2465 12136 2479
rect 26042 2465 26056 2479
rect 9338 2441 9352 2455
rect 11066 2441 11080 2455
rect 23690 2441 23704 2455
rect 9506 2417 9520 2431
rect 9554 2417 9568 2431
rect 9626 2417 9640 2431
rect 22442 2417 22456 2431
rect 9578 2393 9592 2407
rect 19106 2393 19120 2407
rect 20258 2393 20272 2407
rect 9698 2369 9712 2383
rect 15146 2369 15160 2383
rect 9794 2345 9808 2359
rect 20234 2345 20248 2359
rect 25226 2345 25240 2359
rect 25778 2345 25792 2359
rect 9818 2321 9832 2335
rect 11498 2321 11512 2335
rect 11930 2321 11944 2335
rect 12362 2321 12376 2335
rect 14522 2321 14536 2335
rect 16562 2321 16576 2335
rect 22346 2321 22360 2335
rect 24194 2321 24208 2335
rect 26114 2321 26128 2335
rect 10034 2297 10048 2311
rect 23738 2297 23752 2311
rect 10034 2273 10048 2287
rect 13922 2273 13936 2287
rect 17114 2273 17128 2287
rect 10058 2249 10072 2263
rect 10130 2249 10144 2263
rect 10202 2249 10216 2263
rect 10802 2249 10816 2263
rect 12170 2249 12184 2263
rect 25826 2249 25840 2263
rect 10082 2225 10096 2239
rect 22274 2225 22288 2239
rect 10442 2201 10456 2215
rect 18842 2201 18856 2215
rect 21770 2201 21784 2215
rect 10706 2177 10720 2191
rect 10730 2177 10744 2191
rect 10802 2177 10816 2191
rect 12050 2177 12064 2191
rect 14642 2177 14656 2191
rect 14738 2177 14752 2191
rect 22178 2177 22192 2191
rect 10922 2153 10936 2167
rect 11114 2153 11128 2167
rect 23810 2153 23824 2167
rect 10994 2129 11008 2143
rect 12962 2129 12976 2143
rect 13058 2129 13072 2143
rect 20546 2129 20560 2143
rect 22178 2129 22192 2143
rect 22778 2129 22792 2143
rect 11042 2105 11056 2119
rect 11090 2105 11104 2119
rect 11162 2105 11176 2119
rect 11978 2105 11992 2119
rect 12050 2105 12064 2119
rect 19394 2105 19408 2119
rect 11066 2081 11080 2095
rect 27506 2081 27520 2095
rect 11162 2057 11176 2071
rect 21698 2057 21712 2071
rect 11426 2033 11440 2047
rect 13250 2033 13264 2047
rect 13442 2033 13456 2047
rect 22106 2033 22120 2047
rect 11546 2009 11560 2023
rect 16034 2009 16048 2023
rect 20354 2009 20368 2023
rect 11594 1985 11608 1999
rect 24506 1985 24520 1999
rect 26522 1985 26536 1999
rect 11882 1961 11896 1975
rect 15314 1961 15328 1975
rect 15890 1961 15904 1975
rect 17114 1961 17128 1975
rect 21482 1961 21496 1975
rect 11954 1937 11968 1951
rect 12194 1937 12208 1951
rect 12290 1937 12304 1951
rect 24698 1937 24712 1951
rect 12194 1913 12208 1927
rect 12386 1913 12400 1927
rect 12602 1913 12616 1927
rect 23306 1913 23320 1927
rect 12410 1889 12424 1903
rect 25970 1889 25984 1903
rect 12746 1865 12760 1879
rect 12794 1865 12808 1879
rect 12866 1865 12880 1879
rect 16778 1865 16792 1879
rect 23762 1865 23776 1879
rect 12986 1841 13000 1855
rect 15362 1841 15376 1855
rect 16538 1841 16552 1855
rect 18842 1841 18856 1855
rect 27266 1841 27280 1855
rect 13154 1817 13168 1831
rect 22130 1817 22144 1831
rect 27626 1817 27640 1831
rect 27963 1817 27977 1831
rect 13682 1793 13696 1807
rect 13790 1793 13804 1807
rect 14306 1793 14320 1807
rect 14618 1793 14632 1807
rect 15146 1793 15160 1807
rect 21674 1793 21688 1807
rect 27602 1793 27616 1807
rect 27963 1793 27977 1807
rect 14474 1769 14488 1783
rect 14822 1769 14836 1783
rect 15890 1769 15904 1783
rect 21722 1769 21736 1783
rect 22778 1769 22792 1783
rect 26930 1769 26944 1783
rect 27578 1769 27592 1783
rect 27963 1769 27977 1783
rect 14522 1745 14536 1759
rect 25322 1745 25336 1759
rect 27554 1745 27568 1759
rect 27963 1745 27977 1759
rect 19394 1721 19408 1735
rect 27074 1721 27088 1735
rect 27530 1721 27544 1735
rect 27963 1721 27977 1735
rect 14042 888 14056 902
rect 14618 888 14632 902
rect 16610 888 16624 902
rect 24554 888 24568 902
rect 13970 864 13984 878
rect 20762 864 20776 878
rect 22370 864 22384 878
rect 22850 864 22864 878
rect 23810 864 23824 878
rect 24626 864 24640 878
rect 27026 864 27040 878
rect 13778 840 13792 854
rect 18050 840 18064 854
rect 13466 816 13480 830
rect 14066 816 14080 830
rect 15170 816 15184 830
rect 22874 816 22888 830
rect 13370 792 13384 806
rect 19034 792 19048 806
rect 13202 768 13216 782
rect 23546 768 23560 782
rect 12458 744 12472 758
rect 15938 744 15952 758
rect 16466 744 16480 758
rect 22130 744 22144 758
rect 12146 720 12160 734
rect 26810 720 26824 734
rect 11258 696 11272 710
rect 22826 696 22840 710
rect 10370 672 10384 686
rect 11354 672 11368 686
rect 11810 672 11824 686
rect 14690 672 14704 686
rect 14810 672 14824 686
rect 22586 672 22600 686
rect 10346 648 10360 662
rect 11138 648 11152 662
rect 16346 648 16360 662
rect 27050 648 27064 662
rect 10226 624 10240 638
rect 12650 624 12664 638
rect 12698 624 12712 638
rect 14090 624 14104 638
rect 14138 624 14152 638
rect 25970 624 25984 638
rect 10106 600 10120 614
rect 17810 600 17824 614
rect 22154 600 22168 614
rect 23642 600 23656 614
rect 10082 576 10096 590
rect 15698 576 15712 590
rect 16418 576 16432 590
rect 25730 576 25744 590
rect 8810 552 8824 566
rect 11666 552 11680 566
rect 11714 552 11728 566
rect 24506 552 24520 566
rect 8786 528 8800 542
rect 20786 528 20800 542
rect 21674 528 21688 542
rect 24986 528 25000 542
rect 8426 504 8440 518
rect 19298 504 19312 518
rect 20450 504 20464 518
rect 26762 504 26776 518
rect 8282 480 8296 494
rect 24938 480 24952 494
rect 8138 456 8152 470
rect 16874 456 16888 470
rect 17402 456 17416 470
rect 20018 456 20032 470
rect 22226 456 22240 470
rect 23282 456 23296 470
rect 24482 456 24496 470
rect 25010 456 25024 470
rect 25130 456 25144 470
rect 7778 432 7792 446
rect 15218 432 15232 446
rect 17762 432 17776 446
rect 22250 432 22264 446
rect 7418 408 7432 422
rect 16562 408 16576 422
rect 7154 384 7168 398
rect 10754 384 10768 398
rect 11210 384 11224 398
rect 20690 384 20704 398
rect 7034 360 7048 374
rect 12506 360 12520 374
rect 12554 360 12568 374
rect 18410 360 18424 374
rect 6266 336 6280 350
rect 13826 336 13840 350
rect 20402 336 20416 350
rect 27002 336 27016 350
rect 5018 312 5032 326
rect 5066 312 5080 326
rect 5570 312 5584 326
rect 18986 312 19000 326
rect 4778 288 4792 302
rect 10514 288 10528 302
rect 13346 288 13360 302
rect 14186 288 14200 302
rect 20546 288 20560 302
rect 22754 288 22768 302
rect 26978 288 26992 302
rect 4490 264 4504 278
rect 22394 264 22408 278
rect 4346 240 4360 254
rect 6578 240 6592 254
rect 6842 240 6856 254
rect 24530 240 24544 254
rect 4274 216 4288 230
rect 23426 216 23440 230
rect 4226 192 4240 206
rect 19250 192 19264 206
rect 3986 168 4000 182
rect 5162 168 5176 182
rect 5210 168 5224 182
rect 6338 168 6352 182
rect 6506 168 6520 182
rect 21650 168 21664 182
rect 3602 144 3616 158
rect 13538 144 13552 158
rect 24314 144 24328 158
rect 27963 144 27977 158
rect 2882 120 2896 134
rect 4034 120 4048 134
rect 9842 120 9856 134
rect 9938 120 9952 134
rect 19058 120 19072 134
rect 2834 96 2848 110
rect 14930 96 14944 110
rect 27050 96 27064 110
rect 27963 96 27977 110
rect 70 72 84 86
rect 1778 72 1792 86
rect 2714 72 2728 86
rect 14834 72 14848 86
rect 27026 72 27040 86
rect 27963 72 27977 86
rect 70 48 84 62
rect 1730 48 1744 62
rect 2474 48 2488 62
rect 11690 48 11704 62
rect 14210 48 14224 62
rect 18602 48 18616 62
rect 27963 48 27977 62
rect 70 24 84 38
rect 16130 24 16144 38
rect 27002 24 27016 38
rect 27963 24 27977 38
rect 70 0 84 14
rect 26954 0 26968 14
rect 26978 0 26992 14
rect 27963 0 27977 14
<< metal2 >>
rect 0 8867 70 8879
rect 0 8843 70 8855
rect 0 8819 70 8831
rect 123 8616 323 9034
rect 339 8616 351 9034
rect 363 8616 375 9034
rect 387 8616 399 9034
rect 411 8616 423 9034
rect 2391 8928 2403 9034
rect 3951 8952 3963 9034
rect 3952 8938 3970 8952
rect 2392 8914 2410 8928
rect 2043 8616 2055 8890
rect 2211 8616 2223 8794
rect 2379 8616 2391 8914
rect 3243 8616 3255 8914
rect 3675 8616 3687 8770
rect 3939 8616 3951 8938
rect 4131 8616 4143 8938
rect 6171 8760 6183 9034
rect 7275 8616 7287 8962
rect 7707 8736 7719 9034
rect 9243 8712 9255 9034
rect 9291 8616 9303 8674
rect 9891 8616 9903 8986
rect 10779 8664 10791 9034
rect 12315 8832 12327 9034
rect 11211 8616 11223 8818
rect 11715 8616 11727 8650
rect 12363 8616 12375 8650
rect 13347 8616 13359 8794
rect 13851 8640 13863 9034
rect 15387 8640 15399 9034
rect 16047 9024 16059 9034
rect 16048 9010 16066 9024
rect 14835 8616 14847 8626
rect 16035 8616 16047 9010
rect 16935 9000 16947 9034
rect 18459 8976 18471 9034
rect 17139 8616 17151 8746
rect 17283 8616 17295 8818
rect 17523 8616 17535 8818
rect 18699 8616 18711 8794
rect 19983 8760 19995 9034
rect 19179 8616 19191 8698
rect 19227 8616 19239 8746
rect 20259 8616 20271 8842
rect 22743 8760 22755 9034
rect 23031 8952 23043 9034
rect 24555 8904 24567 9034
rect 22744 8746 22762 8760
rect 21099 8616 21111 8626
rect 22731 8616 22743 8746
rect 22779 8616 22791 8866
rect 26079 8832 26091 9034
rect 23355 8616 23367 8722
rect 25827 8616 25839 8746
rect 27507 8616 27519 8818
rect 27531 8640 27543 8770
rect 27555 8712 27567 8914
rect 27579 8784 27591 8794
rect 27579 8736 27591 8746
rect 27603 8688 27615 8746
rect 27627 8688 27639 8818
rect 27651 8616 27851 9034
rect 27977 8771 28047 8783
rect 27977 8747 28047 8759
rect 27977 8723 28047 8735
rect 27977 8699 28047 8711
rect 27977 8675 28047 8687
rect 27977 8651 28047 8663
rect 27977 8627 28047 8639
rect 0 4218 70 4230
rect 0 4194 70 4206
rect 0 4170 70 4182
rect 0 4146 70 4158
rect 123 1711 323 7817
rect 339 1711 351 7817
rect 363 1711 375 7817
rect 387 1711 399 7817
rect 411 1711 423 7817
rect 1611 4255 1623 7817
rect 1659 4327 1671 7817
rect 1731 4351 1743 7817
rect 1755 4375 1767 7817
rect 1803 4423 1815 7817
rect 1851 4447 1863 7817
rect 1611 1711 1623 4121
rect 1635 1711 1647 4265
rect 1659 1711 1671 4289
rect 1683 1711 1695 4217
rect 1731 1711 1743 4217
rect 1779 1711 1791 4385
rect 1875 4111 1887 7817
rect 1899 4495 1911 7817
rect 1923 4519 1935 7817
rect 1971 4543 1983 7817
rect 1995 4567 2007 7817
rect 1899 1711 1911 4457
rect 2091 4087 2103 7817
rect 2115 4591 2127 7817
rect 2139 4615 2151 7817
rect 2187 4639 2199 7817
rect 2235 4663 2247 7817
rect 2283 4687 2295 7817
rect 2307 4711 2319 7817
rect 2331 4735 2343 7817
rect 2259 1711 2271 4049
rect 2307 1711 2319 4025
rect 2379 4015 2391 7817
rect 2427 4759 2439 7817
rect 2451 4783 2463 7817
rect 2451 1711 2463 4697
rect 2475 3991 2487 7817
rect 2523 4807 2535 7817
rect 2547 4231 2559 7817
rect 2571 4447 2583 7817
rect 2619 4447 2631 7817
rect 2667 4831 2679 7817
rect 2739 4855 2751 7817
rect 2499 1711 2511 3953
rect 2547 1711 2559 3929
rect 2571 1711 2583 3905
rect 2619 1711 2631 4217
rect 2667 1711 2679 3881
rect 2763 3871 2775 7817
rect 2787 4879 2799 7817
rect 2787 1711 2799 3833
rect 2811 1711 2823 3809
rect 2835 3799 2847 7817
rect 2859 3775 2871 7817
rect 2907 4903 2919 7817
rect 2955 4951 2967 7817
rect 3003 4975 3015 7817
rect 2907 1711 2919 3737
rect 2931 1711 2943 4913
rect 3051 1711 3063 4985
rect 3075 4255 3087 7817
rect 3099 5023 3111 7817
rect 3147 5047 3159 7817
rect 3195 3727 3207 7817
rect 3219 5071 3231 7817
rect 3291 4255 3303 7817
rect 3315 5095 3327 7817
rect 3339 3703 3351 7817
rect 3387 5119 3399 7817
rect 3411 5143 3423 7817
rect 3459 4135 3471 7817
rect 3507 5167 3519 7817
rect 3531 5191 3543 7817
rect 3579 5215 3591 7817
rect 3627 5239 3639 7817
rect 3411 1711 3423 3665
rect 3459 1711 3471 3737
rect 3603 1711 3615 4361
rect 3651 1711 3663 3641
rect 3723 1711 3735 5249
rect 3747 4039 3759 7817
rect 3771 5311 3783 7817
rect 3795 5335 3807 7817
rect 3843 5383 3855 7817
rect 3867 5431 3879 7817
rect 3747 1711 3759 3617
rect 3771 1711 3783 5273
rect 3819 1711 3831 3593
rect 3843 1711 3855 5345
rect 3867 1711 3879 5393
rect 3891 3583 3903 7817
rect 3939 5455 3951 7817
rect 3987 5479 3999 7817
rect 4011 5503 4023 7817
rect 4035 5527 4047 7817
rect 4083 5575 4095 7817
rect 4203 5599 4215 7817
rect 3915 1711 3927 4961
rect 3939 1711 3951 3593
rect 3963 1711 3975 3809
rect 4083 1711 4095 5537
rect 4227 5383 4239 7817
rect 4155 1711 4167 3545
rect 4179 1711 4191 5009
rect 4251 4303 4263 7817
rect 4299 3535 4311 7817
rect 4323 4303 4335 7817
rect 4347 5623 4359 7817
rect 4371 5647 4383 7817
rect 4419 5671 4431 7817
rect 4203 1711 4215 3521
rect 4299 1711 4311 3497
rect 4395 1711 4407 3809
rect 4419 1711 4431 4337
rect 4443 4231 4455 7817
rect 4443 1711 4455 3473
rect 4467 3463 4479 7817
rect 4515 5695 4527 7817
rect 4539 4711 4551 7817
rect 4563 5719 4575 7817
rect 4611 5767 4623 7817
rect 4515 1711 4527 3425
rect 4539 1711 4551 3401
rect 4563 1711 4575 3377
rect 4587 1711 4599 5729
rect 4659 3559 4671 7817
rect 4731 5791 4743 7817
rect 4755 5815 4767 7817
rect 4779 5839 4791 7817
rect 4827 4831 4839 7817
rect 4851 5863 4863 7817
rect 4875 5887 4887 7817
rect 4923 5911 4935 7817
rect 4947 5839 4959 7817
rect 4971 5935 4983 7817
rect 5019 5959 5031 7817
rect 5043 5863 5055 7817
rect 5067 5983 5079 7817
rect 4635 1711 4647 3353
rect 4659 1711 4671 3329
rect 4683 1711 4695 3641
rect 4707 1711 4719 3305
rect 4755 1711 4767 3281
rect 4803 1711 4815 3257
rect 4851 1711 4863 3233
rect 4875 1711 4887 3209
rect 4923 1711 4935 3185
rect 4971 1711 4983 4697
rect 4995 1711 5007 4049
rect 5115 3655 5127 7817
rect 5139 4351 5151 7817
rect 5163 3223 5175 7817
rect 5211 3271 5223 7817
rect 5259 6031 5271 7817
rect 5331 6079 5343 7817
rect 5355 6127 5367 7817
rect 5403 6151 5415 7817
rect 5451 6223 5463 7817
rect 5475 6247 5487 7817
rect 5499 6271 5511 7817
rect 5547 6319 5559 7817
rect 5091 1711 5103 3161
rect 5115 1711 5127 3137
rect 5187 1711 5199 3113
rect 5259 1711 5271 5993
rect 5283 1711 5295 3689
rect 5307 1711 5319 6041
rect 5331 1711 5343 3689
rect 5355 1711 5367 6089
rect 5403 1711 5415 3089
rect 5427 1711 5439 6161
rect 5451 1711 5463 6185
rect 5499 1711 5511 4577
rect 5523 1711 5535 3065
rect 5547 1711 5559 6281
rect 5571 5767 5583 7817
rect 5619 3079 5631 7817
rect 5667 3055 5679 7817
rect 5691 4303 5703 7817
rect 5739 5167 5751 7817
rect 5787 4255 5799 7817
rect 5811 3679 5823 7817
rect 5835 5167 5847 7817
rect 5883 5527 5895 7817
rect 5907 6343 5919 7817
rect 5955 6367 5967 7817
rect 5691 1711 5703 3017
rect 6003 3007 6015 7817
rect 6027 2983 6039 7817
rect 6051 6391 6063 7817
rect 6075 3031 6087 7817
rect 6123 5287 6135 7817
rect 6147 3031 6159 7817
rect 6171 5287 6183 7817
rect 6195 6415 6207 7817
rect 6051 1711 6063 2945
rect 6099 1711 6111 2921
rect 6219 2911 6231 7817
rect 6267 6439 6279 7817
rect 6291 6463 6303 7817
rect 6339 6487 6351 7817
rect 6291 1711 6303 5465
rect 6363 1711 6375 6497
rect 6387 3151 6399 7817
rect 6411 6535 6423 7817
rect 6435 6559 6447 7817
rect 6483 6583 6495 7817
rect 6507 6607 6519 7817
rect 6435 1711 6447 6329
rect 6531 3463 6543 7817
rect 6555 5359 6567 7817
rect 6459 1711 6471 3137
rect 6483 1711 6495 3449
rect 6555 1711 6567 5057
rect 6603 4807 6615 7817
rect 6627 4399 6639 7817
rect 6651 6631 6663 7817
rect 6603 1711 6615 2873
rect 6627 1711 6639 2849
rect 6651 1711 6663 5441
rect 6675 2863 6687 5825
rect 6699 5359 6711 7817
rect 6723 5455 6735 7817
rect 6699 1711 6711 4217
rect 6723 1711 6735 3281
rect 6747 1711 6759 4385
rect 6771 2863 6783 7817
rect 6819 3607 6831 7817
rect 6843 5503 6855 7817
rect 6867 3127 6879 7817
rect 6915 6511 6927 7817
rect 6939 6655 6951 7817
rect 6963 6511 6975 7817
rect 7011 6679 7023 7817
rect 7035 6703 7047 7817
rect 7059 6751 7071 7817
rect 6795 1711 6807 2825
rect 6819 1711 6831 2801
rect 6891 1711 6903 2777
rect 6939 1711 6951 3329
rect 7011 1711 7023 4817
rect 7035 2935 7047 6665
rect 7059 1711 7071 6713
rect 7107 5743 7119 7817
rect 7131 6679 7143 7817
rect 7179 5743 7191 7817
rect 7107 1711 7119 3617
rect 7131 1711 7143 4217
rect 7227 3319 7239 7817
rect 7251 6775 7263 7817
rect 7323 6799 7335 7817
rect 7347 6823 7359 7817
rect 7371 6847 7383 7817
rect 7203 1711 7215 2753
rect 7227 1711 7239 2729
rect 7251 1711 7263 2705
rect 7299 1711 7311 5369
rect 7323 1711 7335 5585
rect 7395 5335 7407 7817
rect 7419 6871 7431 7817
rect 7467 5335 7479 7817
rect 7491 6895 7503 7817
rect 7539 6919 7551 7817
rect 7587 6943 7599 7817
rect 7347 1711 7359 2681
rect 7371 1711 7383 2657
rect 7443 1711 7455 4409
rect 7467 1711 7479 3785
rect 7515 1711 7527 3785
rect 7539 1711 7551 2825
rect 7587 1711 7599 6929
rect 7611 3631 7623 7817
rect 7635 6967 7647 7817
rect 7635 1711 7647 5369
rect 7683 5311 7695 7817
rect 7659 1711 7671 4025
rect 7707 2647 7719 6305
rect 7731 5455 7743 7817
rect 7803 5383 7815 7817
rect 7827 5455 7839 7817
rect 7851 6991 7863 7817
rect 7683 1711 7695 2633
rect 7731 1711 7743 2609
rect 7755 1711 7767 2633
rect 7803 1711 7815 3137
rect 7827 1711 7839 4625
rect 7851 2743 7863 5441
rect 7899 3847 7911 7817
rect 7923 5455 7935 7817
rect 7947 7015 7959 7817
rect 7995 5479 8007 7817
rect 7875 1711 7887 2585
rect 7923 1711 7935 5081
rect 7947 3679 7959 5441
rect 7995 1711 8007 5441
rect 8019 3919 8031 7817
rect 8043 4447 8055 7817
rect 8091 6871 8103 7817
rect 8067 5455 8079 6329
rect 8115 5455 8127 7817
rect 8163 6871 8175 7817
rect 8043 1711 8055 2561
rect 8115 1711 8127 5369
rect 8139 2575 8151 6233
rect 8163 1711 8175 3977
rect 8187 1711 8199 6809
rect 8211 4855 8223 7817
rect 8235 6823 8247 7817
rect 8259 7039 8271 7817
rect 8235 1711 8247 3977
rect 8259 1711 8271 4697
rect 8283 3415 8295 6857
rect 8307 4183 8319 7817
rect 8355 6871 8367 7817
rect 8331 1711 8343 3593
rect 8355 1711 8367 4169
rect 8379 1711 8391 3401
rect 8427 2575 8439 7817
rect 8451 7063 8463 7817
rect 8475 5479 8487 7817
rect 8499 7087 8511 7817
rect 8523 7111 8535 7817
rect 8571 5383 8583 7817
rect 8595 7135 8607 7817
rect 8451 1711 8463 5081
rect 8475 1711 8487 2537
rect 8523 1711 8535 2513
rect 8595 2503 8607 5777
rect 8619 2623 8631 7817
rect 8667 4783 8679 7817
rect 8715 7159 8727 7817
rect 8571 1711 8583 2489
rect 8643 1711 8655 2801
rect 8667 1711 8679 3281
rect 8715 1711 8727 4289
rect 8739 3295 8751 7145
rect 8787 6895 8799 7817
rect 8835 7159 8847 7817
rect 8907 3583 8919 7817
rect 8763 1711 8775 3569
rect 8931 3535 8943 7817
rect 8931 1711 8943 2609
rect 8955 2503 8967 7817
rect 9003 7183 9015 7817
rect 9027 5815 9039 7817
rect 9051 2479 9063 7817
rect 9099 4543 9111 7817
rect 9123 4039 9135 7817
rect 9147 7207 9159 7817
rect 9195 7231 9207 7817
rect 9219 4447 9231 7817
rect 9243 6919 9255 7817
rect 9267 7255 9279 7817
rect 9339 4783 9351 7817
rect 9363 7087 9375 7817
rect 9387 5863 9399 7817
rect 9411 6919 9423 7817
rect 9435 7279 9447 7817
rect 9483 5095 9495 7817
rect 9507 3679 9519 7817
rect 9531 3991 9543 7817
rect 9339 1711 9351 2441
rect 9483 1711 9495 2561
rect 9507 1711 9519 2417
rect 9531 1711 9543 3929
rect 9555 2431 9567 5849
rect 9579 2839 9591 7817
rect 9603 3991 9615 7817
rect 9579 1711 9591 2393
rect 9603 1711 9615 3161
rect 9627 2431 9639 7817
rect 9651 1711 9663 6113
rect 9675 2647 9687 7817
rect 9699 3559 9711 7817
rect 9747 7327 9759 7817
rect 9795 7351 9807 7817
rect 9699 1711 9711 2369
rect 9723 1711 9735 6113
rect 9747 1711 9759 7289
rect 9819 4375 9831 7817
rect 9843 7375 9855 7817
rect 9891 7303 9903 7817
rect 9795 1711 9807 2345
rect 9819 1711 9831 2321
rect 9891 1711 9903 3593
rect 9915 1711 9927 7385
rect 9939 7303 9951 7817
rect 9963 7423 9975 7817
rect 9987 7447 9999 7817
rect 9987 1711 9999 5777
rect 10011 1711 10023 2585
rect 10035 2311 10047 7817
rect 10035 1711 10047 2273
rect 10059 2263 10071 7817
rect 10083 2239 10095 7817
rect 10107 2623 10119 7817
rect 10155 4423 10167 7817
rect 10131 1711 10143 2249
rect 10179 1711 10191 7433
rect 10203 2623 10215 7817
rect 10275 3895 10287 7817
rect 10299 4567 10311 7817
rect 10323 7447 10335 7817
rect 10203 1711 10215 2249
rect 10275 1711 10287 3545
rect 10299 1711 10311 4025
rect 10323 1711 10335 6209
rect 10347 1711 10359 7337
rect 10371 3463 10383 7817
rect 10419 5959 10431 7817
rect 10419 1711 10431 4817
rect 10443 1711 10455 2201
rect 10467 1711 10479 4817
rect 10491 2839 10503 7817
rect 10515 4039 10527 7817
rect 10539 5359 10551 7817
rect 10587 7471 10599 7817
rect 10563 1711 10575 5849
rect 10611 5503 10623 7817
rect 10635 6295 10647 7817
rect 10635 1711 10647 5801
rect 10659 1711 10671 4697
rect 10683 3751 10695 7817
rect 10707 4711 10719 7817
rect 10731 2191 10743 5441
rect 10707 1711 10719 2177
rect 10779 1711 10791 6977
rect 10803 2263 10815 7817
rect 10875 7063 10887 7817
rect 10899 5455 10911 7817
rect 10803 1711 10815 2177
rect 10851 1711 10863 3617
rect 10875 1711 10887 4409
rect 10923 2575 10935 7817
rect 10947 6295 10959 7817
rect 10995 7495 11007 7817
rect 11019 7159 11031 7817
rect 10923 1711 10935 2153
rect 10971 1711 10983 7145
rect 11043 5095 11055 7817
rect 11067 7519 11079 7817
rect 10995 1711 11007 2129
rect 11019 1711 11031 5057
rect 11067 2455 11079 7145
rect 11091 2119 11103 7241
rect 11115 7159 11127 7817
rect 11139 3175 11151 7817
rect 11043 1711 11055 2105
rect 11067 1711 11079 2081
rect 11115 1711 11127 2153
rect 11163 2119 11175 7817
rect 11211 7543 11223 7817
rect 11259 3823 11271 7817
rect 11283 7543 11295 7817
rect 11307 7471 11319 7817
rect 11163 1711 11175 2057
rect 11331 1711 11343 5561
rect 11355 2743 11367 7817
rect 11403 7567 11415 7817
rect 11475 7591 11487 7817
rect 11379 1711 11391 7457
rect 11427 1711 11439 2033
rect 11475 1711 11487 5801
rect 11499 2335 11511 7817
rect 11523 3703 11535 7817
rect 11571 7615 11583 7817
rect 11547 2599 11559 7577
rect 11595 4063 11607 7817
rect 11547 1711 11559 2009
rect 11571 1711 11583 3809
rect 11619 3679 11631 7601
rect 11643 5191 11655 7817
rect 11691 7591 11703 7817
rect 11595 1711 11607 1985
rect 11643 1711 11655 2825
rect 11691 1711 11703 5609
rect 11715 5191 11727 7817
rect 11763 7615 11775 7817
rect 11811 7639 11823 7817
rect 11835 6439 11847 7817
rect 11859 7663 11871 7817
rect 11883 5863 11895 7817
rect 11907 4687 11919 7817
rect 11763 1711 11775 4625
rect 11787 1711 11799 3233
rect 11859 1711 11871 4625
rect 11883 1711 11895 1961
rect 11907 1711 11919 4097
rect 11931 2335 11943 7649
rect 11955 3103 11967 7817
rect 11979 4231 11991 7817
rect 12003 7663 12015 7817
rect 11955 1711 11967 1937
rect 11979 1711 11991 2105
rect 12003 1711 12015 2465
rect 12027 1711 12039 4673
rect 12051 2191 12063 7817
rect 12075 6943 12087 7817
rect 12099 4111 12111 7817
rect 12147 3703 12159 7817
rect 12171 3823 12183 7817
rect 12219 7063 12231 7817
rect 12267 7663 12279 7817
rect 12291 6271 12303 7817
rect 12051 1711 12063 2105
rect 12099 1711 12111 3689
rect 12123 1711 12135 2465
rect 12171 1711 12183 2249
rect 12195 1951 12207 6257
rect 12315 5263 12327 7817
rect 12363 5263 12375 7817
rect 12195 1711 12207 1913
rect 12243 1711 12255 3593
rect 12267 1711 12279 2729
rect 12291 1711 12303 1937
rect 12339 1711 12351 3377
rect 12363 1711 12375 2321
rect 12387 1927 12399 5249
rect 12411 3487 12423 7817
rect 12435 4303 12447 7817
rect 12459 4375 12471 7817
rect 12483 6847 12495 7817
rect 12531 4399 12543 7817
rect 12555 5263 12567 7817
rect 12579 6847 12591 7817
rect 12627 4711 12639 7817
rect 12651 3943 12663 7817
rect 12411 1711 12423 1889
rect 12483 1711 12495 3929
rect 12675 3391 12687 7817
rect 12723 7663 12735 7817
rect 12747 3535 12759 7817
rect 12771 7687 12783 7817
rect 12579 1711 12591 3281
rect 12603 1711 12615 1913
rect 12675 1711 12687 2825
rect 12747 1711 12759 1865
rect 12771 1711 12783 2585
rect 12795 1879 12807 3785
rect 12819 3295 12831 7817
rect 12843 6919 12855 7817
rect 12867 7639 12879 7817
rect 12915 7711 12927 7817
rect 12939 7735 12951 7817
rect 12819 1711 12831 2633
rect 12867 1711 12879 1865
rect 12915 1711 12927 6665
rect 12963 2143 12975 7817
rect 13011 7759 13023 7817
rect 13035 7783 13047 7817
rect 12987 1711 12999 1841
rect 13011 1711 13023 6737
rect 13083 5599 13095 7817
rect 13131 7807 13143 7817
rect 13035 1711 13047 4961
rect 13059 1711 13071 2129
rect 13107 1711 13119 3281
rect 13131 1711 13143 5849
rect 13155 3535 13167 7817
rect 13179 5263 13191 7817
rect 13203 3799 13215 7745
rect 13227 3799 13239 7817
rect 13251 2047 13263 7817
rect 13275 4399 13287 7769
rect 13299 3103 13311 7817
rect 13155 1711 13167 1817
rect 13323 1711 13335 5441
rect 13347 2743 13359 7793
rect 13419 1711 13431 4241
rect 13467 3535 13479 7817
rect 13491 6919 13503 7817
rect 13515 6439 13527 7817
rect 13563 7351 13575 7817
rect 13611 3823 13623 7817
rect 13443 1711 13455 2033
rect 13515 1711 13527 3353
rect 13587 1711 13599 3089
rect 13635 1711 13647 6929
rect 13659 1711 13671 3545
rect 13683 2671 13695 7817
rect 13707 4111 13719 7817
rect 13731 4831 13743 7817
rect 13755 7759 13767 7817
rect 13779 7591 13791 7817
rect 13827 7279 13839 7817
rect 13851 7567 13863 7817
rect 13683 1711 13695 1793
rect 13731 1711 13743 2657
rect 13755 1711 13767 6953
rect 13791 1807 13803 6257
rect 13827 1711 13839 6905
rect 13899 3151 13911 7817
rect 13875 1711 13887 2561
rect 13923 2287 13935 7745
rect 13947 6367 13959 7817
rect 13971 4831 13983 7817
rect 13947 1711 13959 3641
rect 13971 1711 13983 4769
rect 13995 1711 14007 5417
rect 14019 5239 14031 7817
rect 14067 6991 14079 7817
rect 14115 6175 14127 7817
rect 14115 1711 14127 5345
rect 14187 3103 14199 7817
rect 14211 4231 14223 7817
rect 14235 6343 14247 7817
rect 14259 4111 14271 6449
rect 14283 5383 14295 7817
rect 14235 1711 14247 4097
rect 14283 1711 14295 3137
rect 14307 2815 14319 7817
rect 14307 1711 14319 1793
rect 14331 1711 14343 7409
rect 14355 7303 14367 7817
rect 14379 1711 14391 4697
rect 14403 3943 14415 7817
rect 14427 4783 14439 7817
rect 14403 1711 14415 3665
rect 14427 1711 14439 3785
rect 14451 3151 14463 7673
rect 14475 2743 14487 7817
rect 14475 1711 14487 1769
rect 14499 1711 14511 2825
rect 14523 2335 14535 7817
rect 14547 4711 14559 7817
rect 14523 1711 14535 1745
rect 14571 1711 14583 4769
rect 14595 4255 14607 7817
rect 14595 1711 14607 3665
rect 14619 1807 14631 7265
rect 14643 2191 14655 7817
rect 14667 3679 14679 7817
rect 14691 4975 14703 7817
rect 14667 1711 14679 3137
rect 14715 1711 14727 7025
rect 14739 2551 14751 7817
rect 14763 7111 14775 7817
rect 14787 5263 14799 7817
rect 14811 4135 14823 7817
rect 14883 4351 14895 7817
rect 14931 4759 14943 7817
rect 14739 1711 14751 2177
rect 14787 1711 14799 4097
rect 14823 1783 14835 3569
rect 14859 1711 14871 4121
rect 14883 1711 14895 4193
rect 14955 1711 14967 6305
rect 14979 1711 14991 4073
rect 15003 3343 15015 7817
rect 15027 3103 15039 7817
rect 15051 5575 15063 7817
rect 15075 4207 15087 7049
rect 15099 5431 15111 7817
rect 15027 1711 15039 2777
rect 15051 1711 15063 4193
rect 15099 1711 15111 5177
rect 15123 3343 15135 7817
rect 15147 2383 15159 7817
rect 15195 5191 15207 7817
rect 15219 7711 15231 7817
rect 15243 5623 15255 7817
rect 15267 5575 15279 7817
rect 15315 1975 15327 7817
rect 15339 6175 15351 7817
rect 15147 1711 15159 1793
rect 15339 1711 15351 5921
rect 15363 1855 15375 7817
rect 15387 2959 15399 6161
rect 15483 4519 15495 7817
rect 15843 6703 15855 7817
rect 15747 1711 15759 4505
rect 15891 1975 15903 7817
rect 15891 1711 15903 1769
rect 15915 1711 15927 4193
rect 15987 1711 15999 7241
rect 16035 5935 16047 7817
rect 16155 6103 16167 7817
rect 16035 1711 16047 2009
rect 16107 1711 16119 4793
rect 16155 1711 16167 2993
rect 16203 1711 16215 6449
rect 16251 1711 16263 6641
rect 16323 1711 16335 5489
rect 16371 1711 16383 2681
rect 16443 1711 16455 5801
rect 16515 5383 16527 7817
rect 16515 1711 16527 4073
rect 16563 2335 16575 7817
rect 16587 4087 16599 6737
rect 16707 4207 16719 7817
rect 16755 6535 16767 7817
rect 16827 4951 16839 7817
rect 16539 1711 16551 1841
rect 16659 1711 16671 4073
rect 16731 1711 16743 4289
rect 16755 1711 16767 3905
rect 16779 1711 16791 1865
rect 16827 1711 16839 3953
rect 16851 3223 16863 7817
rect 16875 7375 16887 7817
rect 16899 3991 16911 7817
rect 16947 7303 16959 7817
rect 16971 5815 16983 7817
rect 16995 6007 17007 7817
rect 17043 6007 17055 7817
rect 17067 6103 17079 7817
rect 16947 1711 16959 5369
rect 17091 5287 17103 7817
rect 16971 1711 16983 3665
rect 17019 1711 17031 5009
rect 17067 1711 17079 4433
rect 17091 1711 17103 3329
rect 17115 2287 17127 7817
rect 17115 1711 17127 1961
rect 17139 1711 17151 6113
rect 17187 5479 17199 7817
rect 17211 6487 17223 7817
rect 17235 6535 17247 7817
rect 17163 1711 17175 4433
rect 17211 1711 17223 2993
rect 17235 1711 17247 6425
rect 17259 3343 17271 6281
rect 17283 4447 17295 7817
rect 17283 1711 17295 2945
rect 17307 2791 17319 6521
rect 17331 3199 17343 7817
rect 17355 7351 17367 7817
rect 17379 6175 17391 7817
rect 17427 6271 17439 7817
rect 17451 6295 17463 7817
rect 17475 2503 17487 7817
rect 17499 7207 17511 7817
rect 17571 6943 17583 7817
rect 17595 4783 17607 7817
rect 17643 2767 17655 7817
rect 17691 5239 17703 7817
rect 17715 7255 17727 7817
rect 17739 5239 17751 7817
rect 17787 5023 17799 7817
rect 17811 3559 17823 7817
rect 17835 4135 17847 7817
rect 17883 3295 17895 7817
rect 17907 4039 17919 7817
rect 17931 7087 17943 7817
rect 17955 7039 17967 7817
rect 17955 1711 17967 7001
rect 18003 6343 18015 7817
rect 17979 1711 17991 5153
rect 18027 4711 18039 7817
rect 18003 1711 18015 3881
rect 18051 3439 18063 7817
rect 18075 1711 18087 7649
rect 18099 3127 18111 7817
rect 18147 7711 18159 7817
rect 18123 2791 18135 5273
rect 18099 1711 18111 2777
rect 18147 1711 18159 5345
rect 18195 1711 18207 4553
rect 18267 1711 18279 7313
rect 18291 6367 18303 7817
rect 18291 1711 18303 5489
rect 18315 1711 18327 6401
rect 18363 1711 18375 7217
rect 18483 1711 18495 7409
rect 18531 1711 18543 4553
rect 18651 1711 18663 3905
rect 18723 1711 18735 4433
rect 18771 1711 18783 4121
rect 18843 2215 18855 7817
rect 18867 3919 18879 7817
rect 18915 6535 18927 7817
rect 18843 1711 18855 1841
rect 18867 1711 18879 2873
rect 18891 1711 18903 6497
rect 18915 1711 18927 6401
rect 18963 4543 18975 7817
rect 18987 5095 18999 7817
rect 19011 6415 19023 7817
rect 18939 1711 18951 3881
rect 19011 1711 19023 5561
rect 19059 5047 19071 7817
rect 19083 1711 19095 5321
rect 19107 2407 19119 7817
rect 19131 1711 19143 4577
rect 19179 3895 19191 7817
rect 19155 1711 19167 3617
rect 19203 1711 19215 6209
rect 19227 4135 19239 7817
rect 19275 7735 19287 7817
rect 19299 6223 19311 7817
rect 19323 7351 19335 7817
rect 19347 6775 19359 7817
rect 19275 1711 19287 4313
rect 19347 1711 19359 6017
rect 19371 1711 19383 3521
rect 19395 2119 19407 7817
rect 19443 4279 19455 7817
rect 19395 1711 19407 1721
rect 19443 1711 19455 2825
rect 19467 1711 19479 4049
rect 19515 3271 19527 7817
rect 19539 7039 19551 7817
rect 19563 6463 19575 7817
rect 19587 5695 19599 7817
rect 19635 7231 19647 7817
rect 19491 1711 19503 2585
rect 19611 1711 19623 6857
rect 19659 5887 19671 7817
rect 19683 5407 19695 7817
rect 19707 4807 19719 7817
rect 19755 4399 19767 7817
rect 19803 7735 19815 7817
rect 19875 7711 19887 7817
rect 19899 6247 19911 7817
rect 19923 5071 19935 7817
rect 19971 3751 19983 7817
rect 19995 3175 20007 7817
rect 20019 5095 20031 7817
rect 20067 4855 20079 7817
rect 20091 5287 20103 7817
rect 20115 6391 20127 7817
rect 20163 3391 20175 7817
rect 20187 5335 20199 7817
rect 20211 5215 20223 7817
rect 20235 5095 20247 7817
rect 20163 1711 20175 2585
rect 20187 1711 20199 4697
rect 20259 2407 20271 5321
rect 20235 1711 20247 2345
rect 20283 1711 20295 7697
rect 20307 5095 20319 7817
rect 20331 7351 20343 7817
rect 20307 1711 20319 2729
rect 20331 1711 20343 3017
rect 20355 2023 20367 5081
rect 20379 4855 20391 7817
rect 20427 6175 20439 7817
rect 20451 5095 20463 7817
rect 20475 4903 20487 7817
rect 20499 6175 20511 7817
rect 20523 7759 20535 7817
rect 20379 1711 20391 4289
rect 20499 1711 20511 5945
rect 20523 1711 20535 7697
rect 20547 2143 20559 6161
rect 20571 2959 20583 7817
rect 20595 5863 20607 7817
rect 20619 7231 20631 7817
rect 20571 1711 20583 2777
rect 20619 1711 20631 6473
rect 20643 1711 20655 6521
rect 20667 4375 20679 7817
rect 20691 3247 20703 7817
rect 20715 4351 20727 7817
rect 20739 5095 20751 7817
rect 20763 5431 20775 7745
rect 20787 4423 20799 7817
rect 20739 1711 20751 3977
rect 20811 2647 20823 7817
rect 20835 5503 20847 7817
rect 20859 7759 20871 7817
rect 20835 1711 20847 4217
rect 20859 1711 20871 7697
rect 20907 5647 20919 7817
rect 20931 5719 20943 7817
rect 20883 1711 20895 4409
rect 20907 1711 20919 4385
rect 20955 4087 20967 7817
rect 20979 6559 20991 7817
rect 21003 5095 21015 7817
rect 21051 6127 21063 7817
rect 20955 1711 20967 2873
rect 20979 1711 20991 4409
rect 21003 1711 21015 5057
rect 21087 4423 21099 7601
rect 21027 1711 21039 4001
rect 21075 1711 21087 4217
rect 21123 1711 21135 7121
rect 21147 2671 21159 7745
rect 21171 2527 21183 7817
rect 21195 2839 21207 7817
rect 21243 4831 21255 7817
rect 21195 1711 21207 2657
rect 21219 1711 21231 4049
rect 21267 1711 21279 6065
rect 21291 5167 21303 7817
rect 21339 4543 21351 7817
rect 21375 4423 21387 4937
rect 21411 4615 21423 7817
rect 21315 1711 21327 3209
rect 21339 1711 21351 4409
rect 21363 1711 21375 3689
rect 21435 3415 21447 7817
rect 21411 1711 21423 2993
rect 21459 1711 21471 3593
rect 21483 1975 21495 7817
rect 21531 6247 21543 7817
rect 21531 1711 21543 6209
rect 21555 4111 21567 7817
rect 21579 7159 21591 7817
rect 21627 7351 21639 7817
rect 21555 1711 21567 3545
rect 21579 1711 21591 6257
rect 21627 1711 21639 7289
rect 21651 4231 21663 7817
rect 21675 1807 21687 7817
rect 21699 2071 21711 7337
rect 21723 5791 21735 7817
rect 21747 2839 21759 7817
rect 21771 4687 21783 7817
rect 21819 4063 21831 7817
rect 21843 3175 21855 7817
rect 21867 4903 21879 7817
rect 21723 1711 21735 1769
rect 21771 1711 21783 2201
rect 21843 1711 21855 2729
rect 21867 1711 21879 3905
rect 21891 1711 21903 5753
rect 21915 2767 21927 7817
rect 21939 6847 21951 7817
rect 21939 1711 21951 3929
rect 21963 3511 21975 7817
rect 21963 1711 21975 3281
rect 21987 1711 21999 6569
rect 22011 5071 22023 7817
rect 22035 5215 22047 7817
rect 22059 5191 22071 7817
rect 22035 1711 22047 4841
rect 22059 1711 22071 4673
rect 22083 1711 22095 4481
rect 22107 2047 22119 4889
rect 22131 1831 22143 5201
rect 22179 2191 22191 7817
rect 22179 1711 22191 2129
rect 22275 1711 22287 2225
rect 22323 1711 22335 3641
rect 22347 1711 22359 2321
rect 22443 1711 22455 2417
rect 22467 1711 22479 7073
rect 22491 1711 22503 3041
rect 22539 1711 22551 7169
rect 22587 3247 22599 7817
rect 22731 7471 22743 7817
rect 22563 1711 22575 3161
rect 22635 1711 22647 4241
rect 22659 1711 22671 4025
rect 22683 1711 22695 4097
rect 22731 1711 22743 2561
rect 22779 2143 22791 7817
rect 22827 5047 22839 7817
rect 22851 4855 22863 7817
rect 22899 2671 22911 7817
rect 22947 4903 22959 7817
rect 22971 5863 22983 7817
rect 22995 4207 23007 7817
rect 23043 5527 23055 7817
rect 23091 5455 23103 7817
rect 22779 1711 22791 1769
rect 22923 1711 22935 3209
rect 22947 1711 22959 3809
rect 22971 1711 22983 3761
rect 23019 1711 23031 4625
rect 23043 1711 23055 2921
rect 23067 1711 23079 2969
rect 23115 1711 23127 3737
rect 23139 1711 23151 7529
rect 23163 5503 23175 7817
rect 23211 4903 23223 7817
rect 23283 6727 23295 7817
rect 23187 1711 23199 4841
rect 23235 1711 23247 6665
rect 23259 1711 23271 5849
rect 23307 1927 23319 7817
rect 23331 4855 23343 7817
rect 23403 7711 23415 7817
rect 23331 1711 23343 4025
rect 23355 1711 23367 3617
rect 23379 1711 23391 5585
rect 23403 1711 23415 3809
rect 23427 3559 23439 7817
rect 23451 6103 23463 7817
rect 23475 1711 23487 7649
rect 23499 6391 23511 7817
rect 23523 7663 23535 7817
rect 23499 1711 23511 6209
rect 23535 3535 23547 4889
rect 23571 3847 23583 7817
rect 23619 5623 23631 7817
rect 23643 5503 23655 7817
rect 23691 7087 23703 7817
rect 23523 1711 23535 3089
rect 23595 1711 23607 4817
rect 23619 1711 23631 4025
rect 23655 2791 23667 4841
rect 23691 1711 23703 2441
rect 23715 1711 23727 6113
rect 23739 4735 23751 7817
rect 23739 1711 23751 2297
rect 23763 1879 23775 7817
rect 23787 7495 23799 7817
rect 23787 1711 23799 3593
rect 23811 2167 23823 6377
rect 23835 3799 23847 7817
rect 23859 5527 23871 7817
rect 23859 1711 23871 5465
rect 23883 3175 23895 5513
rect 23907 4591 23919 7817
rect 23955 6631 23967 7817
rect 23907 1711 23919 4529
rect 23931 1711 23943 5369
rect 23979 4663 23991 7817
rect 24003 4879 24015 7817
rect 24027 6367 24039 7817
rect 23955 1711 23967 4577
rect 23979 1711 23991 2681
rect 24003 1711 24015 4721
rect 24051 1711 24063 2897
rect 24075 2839 24087 7817
rect 24099 5503 24111 7817
rect 24123 6343 24135 7817
rect 24147 4543 24159 7721
rect 24075 1711 24087 2777
rect 24123 1711 24135 3713
rect 24171 2647 24183 7817
rect 24171 1711 24183 2585
rect 24195 2335 24207 7817
rect 24219 7207 24231 7817
rect 24219 1711 24231 7169
rect 24243 2791 24255 4817
rect 24267 3679 24279 7817
rect 24291 4831 24303 7817
rect 24315 5815 24327 7817
rect 24363 5383 24375 7817
rect 24387 5503 24399 7817
rect 24291 1711 24303 4745
rect 24339 1711 24351 4937
rect 24387 1711 24399 2945
rect 24411 1711 24423 6017
rect 24435 3631 24447 7817
rect 24435 1711 24447 3593
rect 24459 2599 24471 4961
rect 24483 4519 24495 7817
rect 24507 1999 24519 7817
rect 24531 5911 24543 7817
rect 24543 4567 24555 4817
rect 24579 4255 24591 7817
rect 24603 4831 24615 7817
rect 24603 1711 24615 4217
rect 24627 2527 24639 7817
rect 24675 7687 24687 7817
rect 24651 3007 24663 7193
rect 24675 1711 24687 7649
rect 24699 1951 24711 7817
rect 24723 1711 24735 4793
rect 24747 2887 24759 7817
rect 24795 6151 24807 7817
rect 24771 1711 24783 5249
rect 24807 3751 24819 4817
rect 24843 4471 24855 7817
rect 24843 1711 24855 3833
rect 24867 1711 24879 2633
rect 24891 1711 24903 7241
rect 24915 3847 24927 7817
rect 24939 4591 24951 7817
rect 24963 6295 24975 7817
rect 24963 1711 24975 4745
rect 24987 4399 24999 7673
rect 25011 5551 25023 7817
rect 25035 3751 25047 7817
rect 25059 6127 25071 7817
rect 25083 4759 25095 6401
rect 25107 3487 25119 7817
rect 25155 3367 25167 7817
rect 25227 2359 25239 7817
rect 25251 3679 25263 7817
rect 25275 6055 25287 7817
rect 25323 1759 25335 7817
rect 25347 7447 25359 7817
rect 25371 6271 25383 7817
rect 25395 4159 25407 7817
rect 25443 4591 25455 7817
rect 25467 3079 25479 7817
rect 25491 4831 25503 7817
rect 25515 4447 25527 7817
rect 25563 5167 25575 7817
rect 25491 1711 25503 2801
rect 25539 1711 25551 4697
rect 25587 2839 25599 7817
rect 25635 5119 25647 7817
rect 25683 6439 25695 7817
rect 25707 6655 25719 7817
rect 25731 6607 25743 7817
rect 25779 5743 25791 7817
rect 25611 2695 25623 4817
rect 25683 1711 25695 4961
rect 25707 1711 25719 5153
rect 25803 4831 25815 7817
rect 25779 1711 25791 2345
rect 25803 1711 25815 3737
rect 25827 2263 25839 4817
rect 25851 1711 25863 5129
rect 25875 4831 25887 7817
rect 25899 5839 25911 7817
rect 25923 6895 25935 7817
rect 25971 1903 25983 7817
rect 25995 2863 26007 7817
rect 26043 2479 26055 7817
rect 26091 3967 26103 7817
rect 26115 2335 26127 7817
rect 26139 6799 26151 7817
rect 26187 3919 26199 7817
rect 26211 3823 26223 7817
rect 26235 5311 26247 7817
rect 26283 2743 26295 7817
rect 26307 5023 26319 7817
rect 26331 3535 26343 7817
rect 26355 6247 26367 7817
rect 26331 1711 26343 3161
rect 26379 1711 26391 2825
rect 26403 2719 26415 7817
rect 26427 4735 26439 7817
rect 26475 6007 26487 7817
rect 26523 3079 26535 7817
rect 26547 3679 26559 7817
rect 26523 1711 26535 1985
rect 26547 1711 26559 3305
rect 26571 1711 26583 6113
rect 26595 3583 26607 7817
rect 26643 6319 26655 7817
rect 26619 3559 26631 5921
rect 26691 4783 26703 7817
rect 26763 7639 26775 7817
rect 26715 4759 26727 7313
rect 26787 6439 26799 7817
rect 26811 5863 26823 7817
rect 26595 1711 26607 3545
rect 26643 1711 26655 4745
rect 26667 1711 26679 3617
rect 26691 1711 26703 4721
rect 26739 1711 26751 5081
rect 26835 4183 26847 7817
rect 26883 5983 26895 7817
rect 26907 5695 26919 7817
rect 26859 1711 26871 2609
rect 26883 1711 26895 5489
rect 26907 1711 26919 5657
rect 26931 1783 26943 7817
rect 26955 7399 26967 7817
rect 26955 1711 26967 4769
rect 26979 4735 26991 4817
rect 27003 3919 27015 7817
rect 27027 6919 27039 7817
rect 27051 3463 27063 7817
rect 27099 7519 27111 7817
rect 27075 1735 27087 5681
rect 27123 4927 27135 7817
rect 27147 4999 27159 7817
rect 27195 3607 27207 7817
rect 27219 6199 27231 7817
rect 27267 1855 27279 7817
rect 27315 4807 27327 7817
rect 27339 4783 27351 7817
rect 27363 3151 27375 7817
rect 27411 3103 27423 7817
rect 27435 2575 27447 7817
rect 27459 5071 27471 7817
rect 27507 2095 27519 7817
rect 27531 1735 27543 4337
rect 27555 1759 27567 5489
rect 27579 1783 27591 5273
rect 27603 1807 27615 4673
rect 27627 1831 27639 6809
rect 27651 1711 27851 7817
rect 27977 5226 28047 5238
rect 27977 3858 28047 3870
rect 27977 1818 28047 1830
rect 27977 1794 28047 1806
rect 27977 1770 28047 1782
rect 27977 1746 28047 1758
rect 27977 1722 28047 1734
rect 0 73 70 85
rect 0 49 70 61
rect 0 25 70 37
rect 0 1 70 13
rect 123 0 323 912
rect 339 0 351 912
rect 363 0 375 912
rect 387 0 399 912
rect 411 0 423 912
rect 1731 62 1743 912
rect 1779 86 1791 912
rect 2475 62 2487 912
rect 2715 86 2727 912
rect 2835 110 2847 912
rect 2883 134 2895 912
rect 3603 158 3615 912
rect 3987 182 3999 912
rect 4035 134 4047 912
rect 4227 206 4239 912
rect 4275 230 4287 912
rect 4347 254 4359 912
rect 4491 278 4503 912
rect 4779 302 4791 912
rect 5019 326 5031 912
rect 5067 326 5079 912
rect 5163 182 5175 912
rect 5211 182 5223 912
rect 5571 326 5583 912
rect 6267 350 6279 912
rect 6339 182 6351 912
rect 6507 182 6519 912
rect 6579 254 6591 912
rect 6843 254 6855 912
rect 7035 374 7047 912
rect 7155 398 7167 912
rect 7419 422 7431 912
rect 7779 446 7791 912
rect 8139 470 8151 912
rect 8283 494 8295 912
rect 8427 518 8439 912
rect 8787 542 8799 912
rect 8811 566 8823 912
rect 9843 134 9855 912
rect 9939 134 9951 912
rect 10083 590 10095 912
rect 10107 614 10119 912
rect 10227 638 10239 912
rect 10347 662 10359 912
rect 10371 686 10383 912
rect 10515 302 10527 912
rect 10755 398 10767 912
rect 11139 662 11151 912
rect 11211 398 11223 912
rect 11259 710 11271 912
rect 11355 686 11367 912
rect 11667 566 11679 912
rect 11691 62 11703 912
rect 11715 566 11727 912
rect 11811 686 11823 912
rect 12147 734 12159 912
rect 12459 758 12471 912
rect 12507 374 12519 912
rect 12555 374 12567 912
rect 12651 638 12663 912
rect 12699 638 12711 912
rect 13203 782 13215 912
rect 13347 302 13359 912
rect 13371 806 13383 912
rect 13467 830 13479 912
rect 13539 158 13551 912
rect 13779 854 13791 912
rect 13827 350 13839 912
rect 13971 878 13983 912
rect 14043 902 14055 912
rect 14067 830 14079 912
rect 14091 638 14103 912
rect 14139 638 14151 912
rect 14187 302 14199 912
rect 14211 62 14223 912
rect 14619 902 14631 912
rect 14691 686 14703 912
rect 14811 686 14823 912
rect 14835 86 14847 912
rect 14931 110 14943 912
rect 15171 830 15183 912
rect 15219 446 15231 912
rect 15699 590 15711 912
rect 15939 758 15951 912
rect 16131 38 16143 912
rect 16347 662 16359 912
rect 16419 590 16431 912
rect 16467 758 16479 912
rect 16563 422 16575 912
rect 16611 902 16623 912
rect 16875 470 16887 912
rect 17403 470 17415 912
rect 17763 446 17775 912
rect 17811 614 17823 912
rect 18051 854 18063 912
rect 18411 374 18423 912
rect 18603 62 18615 912
rect 18987 326 18999 912
rect 19035 806 19047 912
rect 19059 134 19071 912
rect 19251 206 19263 912
rect 19299 518 19311 912
rect 20019 470 20031 912
rect 20403 350 20415 912
rect 20451 518 20463 912
rect 20547 302 20559 912
rect 20691 398 20703 912
rect 20763 878 20775 912
rect 20787 542 20799 912
rect 21651 182 21663 912
rect 21675 542 21687 912
rect 22131 758 22143 912
rect 22155 614 22167 912
rect 22227 470 22239 912
rect 22251 446 22263 912
rect 22371 878 22383 912
rect 22395 278 22407 912
rect 22587 686 22599 912
rect 22755 302 22767 912
rect 22827 710 22839 912
rect 22851 878 22863 912
rect 22875 830 22887 912
rect 23283 470 23295 912
rect 23427 230 23439 912
rect 23547 782 23559 912
rect 23643 614 23655 912
rect 23811 878 23823 912
rect 24315 158 24327 912
rect 24483 470 24495 912
rect 24507 566 24519 912
rect 24531 254 24543 912
rect 24555 902 24567 912
rect 24627 878 24639 912
rect 24939 494 24951 912
rect 24987 542 24999 912
rect 25011 470 25023 912
rect 25131 470 25143 912
rect 25731 590 25743 912
rect 25971 638 25983 912
rect 26763 518 26775 912
rect 26811 734 26823 912
rect 26955 14 26967 912
rect 26979 14 26991 288
rect 27003 38 27015 336
rect 27027 86 27039 864
rect 27051 110 27063 648
rect 27651 0 27851 912
rect 27977 145 28047 157
rect 27977 97 28047 109
rect 27977 73 28047 85
rect 27977 49 28047 61
rect 27977 25 28047 37
rect 27977 1 28047 13
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7817
box 0 0 1464 799
use inv g8364
timestamp 1386238110
transform 1 0 1587 0 1 7817
box 0 0 120 799
use nor2 g8043
timestamp 1386235306
transform 1 0 1707 0 1 7817
box 0 0 120 799
use nand3 g8291
timestamp 1386234893
transform 1 0 1827 0 1 7817
box 0 0 120 799
use and2 g8112
timestamp 1386234845
transform 1 0 1947 0 1 7817
box 0 0 120 799
use nand2 g8060
timestamp 1386234792
transform 1 0 2067 0 1 7817
box 0 0 96 799
use nand2 g8182
timestamp 1386234792
transform 1 0 2163 0 1 7817
box 0 0 96 799
use nand2 g8369
timestamp 1386234792
transform 1 0 2259 0 1 7817
box 0 0 96 799
use rowcrosser PcWe
timestamp 1386086759
transform 1 0 2355 0 1 7817
box 0 0 48 799
use nand2 g8066
timestamp 1386234792
transform 1 0 2403 0 1 7817
box 0 0 96 799
use nand2 g8169
timestamp 1386234792
transform 1 0 2499 0 1 7817
box 0 0 96 799
use inv g8107
timestamp 1386238110
transform 1 0 2595 0 1 7817
box 0 0 120 799
use nand2 g8229
timestamp 1386234792
transform 1 0 2715 0 1 7817
box 0 0 96 799
use and2 g8370
timestamp 1386234845
transform 1 0 2811 0 1 7817
box 0 0 120 799
use inv g8313
timestamp 1386238110
transform 1 0 2931 0 1 7817
box 0 0 120 799
use nor2 g8039
timestamp 1386235306
transform 1 0 3051 0 1 7817
box 0 0 120 799
use nand2 g8344
timestamp 1386234792
transform 1 0 3171 0 1 7817
box 0 0 96 799
use nand2 g8222
timestamp 1386234792
transform 1 0 3267 0 1 7817
box 0 0 96 799
use nor2 g8098
timestamp 1386235306
transform 1 0 3363 0 1 7817
box 0 0 120 799
use nor2 g8102
timestamp 1386235306
transform 1 0 3483 0 1 7817
box 0 0 120 799
use inv g8314
timestamp 1386238110
transform 1 0 3603 0 1 7817
box 0 0 120 799
use nand2 g8327
timestamp 1386234792
transform 1 0 3723 0 1 7817
box 0 0 96 799
use nand2 g8187
timestamp 1386234792
transform 1 0 3819 0 1 7817
box 0 0 96 799
use rowcrosser nWait
timestamp 1386086759
transform 1 0 3915 0 1 7817
box 0 0 48 799
use nand2 g8135
timestamp 1386234792
transform 1 0 3963 0 1 7817
box 0 0 96 799
use inv g8171
timestamp 1386238110
transform 1 0 4059 0 1 7817
box 0 0 120 799
use nand2 g8295
timestamp 1386234792
transform 1 0 4179 0 1 7817
box 0 0 96 799
use nand3 g8287
timestamp 1386234893
transform 1 0 4275 0 1 7817
box 0 0 120 799
use nand2 g8154
timestamp 1386234792
transform 1 0 4395 0 1 7817
box 0 0 96 799
use nand2 g8261
timestamp 1386234792
transform 1 0 4491 0 1 7817
box 0 0 96 799
use inv g8276
timestamp 1386238110
transform 1 0 4587 0 1 7817
box 0 0 120 799
use nand2 g8130
timestamp 1386234792
transform 1 0 4707 0 1 7817
box 0 0 96 799
use nand2 g8082
timestamp 1386234792
transform 1 0 4803 0 1 7817
box 0 0 96 799
use nand2 g8318
timestamp 1386234792
transform 1 0 4899 0 1 7817
box 0 0 96 799
use nand2 g8377
timestamp 1386234792
transform 1 0 4995 0 1 7817
box 0 0 96 799
use nand2 g8390
timestamp 1386234792
transform 1 0 5091 0 1 7817
box 0 0 96 799
use inv g8168
timestamp 1386238110
transform 1 0 5187 0 1 7817
box 0 0 120 799
use nor2 g8238
timestamp 1386235306
transform 1 0 5307 0 1 7817
box 0 0 120 799
use nand2 g8225
timestamp 1386234792
transform 1 0 5427 0 1 7817
box 0 0 96 799
use nor2 g8143
timestamp 1386235306
transform 1 0 5523 0 1 7817
box 0 0 120 799
use and2 g8333
timestamp 1386234845
transform 1 0 5643 0 1 7817
box 0 0 120 799
use nand2 g8149
timestamp 1386234792
transform 1 0 5763 0 1 7817
box 0 0 96 799
use nor2 g8042
timestamp 1386235306
transform 1 0 5859 0 1 7817
box 0 0 120 799
use nand3 g8069
timestamp 1386234893
transform 1 0 5979 0 1 7817
box 0 0 120 799
use nand4 g8338
timestamp 1386234936
transform 1 0 6099 0 1 7817
box 0 0 144 799
use nor2 g8280
timestamp 1386235306
transform 1 0 6243 0 1 7817
box 0 0 120 799
use nand2 g8249
timestamp 1386234792
transform 1 0 6363 0 1 7817
box 0 0 96 799
use nand3 g8064
timestamp 1386234893
transform 1 0 6459 0 1 7817
box 0 0 120 799
use nand2 g8310
timestamp 1386234792
transform 1 0 6579 0 1 7817
box 0 0 96 799
use nor2 g8235
timestamp 1386235306
transform 1 0 6675 0 1 7817
box 0 0 120 799
use nand2 g8058
timestamp 1386234792
transform 1 0 6795 0 1 7817
box 0 0 96 799
use nand2 g8362
timestamp 1386234792
transform 1 0 6891 0 1 7817
box 0 0 96 799
use nand2 g8055
timestamp 1386234792
transform 1 0 6987 0 1 7817
box 0 0 96 799
use nor2 g8088
timestamp 1386235306
transform 1 0 7083 0 1 7817
box 0 0 120 799
use nand2 g8214
timestamp 1386234792
transform 1 0 7203 0 1 7817
box 0 0 96 799
use nand4 g8056
timestamp 1386234936
transform 1 0 7299 0 1 7817
box 0 0 144 799
use nor2 g8281
timestamp 1386235306
transform 1 0 7443 0 1 7817
box 0 0 120 799
use nand2 g8366
timestamp 1386234792
transform 1 0 7563 0 1 7817
box 0 0 96 799
use inv g8269
timestamp 1386238110
transform 1 0 7659 0 1 7817
box 0 0 120 799
use nand2 g8183
timestamp 1386234792
transform 1 0 7779 0 1 7817
box 0 0 96 799
use nand2 g8170
timestamp 1386234792
transform 1 0 7875 0 1 7817
box 0 0 96 799
use nand2 g8124
timestamp 1386234792
transform 1 0 7971 0 1 7817
box 0 0 96 799
use nor2 g8106
timestamp 1386235306
transform 1 0 8067 0 1 7817
box 0 0 120 799
use nand2 g8414
timestamp 1386234792
transform 1 0 8187 0 1 7817
box 0 0 96 799
use inv g8119
timestamp 1386238110
transform 1 0 8283 0 1 7817
box 0 0 120 799
use nand4 g8275
timestamp 1386234936
transform 1 0 8403 0 1 7817
box 0 0 144 799
use nand2 g8418
timestamp 1386234792
transform 1 0 8547 0 1 7817
box 0 0 96 799
use inv g8146
timestamp 1386238110
transform 1 0 8643 0 1 7817
box 0 0 120 799
use inv g8127
timestamp 1386238110
transform 1 0 8763 0 1 7817
box 0 0 120 799
use nand2 g8155
timestamp 1386234792
transform 1 0 8883 0 1 7817
box 0 0 96 799
use nand2 g8290
timestamp 1386234792
transform 1 0 8979 0 1 7817
box 0 0 96 799
use nand2 g8033
timestamp 1386234792
transform 1 0 9075 0 1 7817
box 0 0 96 799
use nand4 g8252
timestamp 1386234936
transform 1 0 9171 0 1 7817
box 0 0 144 799
use nand4 g8334
timestamp 1386234936
transform 1 0 9315 0 1 7817
box 0 0 144 799
use nand2 g8244
timestamp 1386234792
transform 1 0 9459 0 1 7817
box 0 0 96 799
use nand2 g8240
timestamp 1386234792
transform 1 0 9555 0 1 7817
box 0 0 96 799
use and2 g8407
timestamp 1386234845
transform 1 0 9651 0 1 7817
box 0 0 120 799
use nand2 g8139
timestamp 1386234792
transform 1 0 9771 0 1 7817
box 0 0 96 799
use rowcrosser g8048
timestamp 1386086759
transform 1 0 9867 0 1 7817
box 0 0 48 799
use nand2 g8118
timestamp 1386234792
transform 1 0 9915 0 1 7817
box 0 0 96 799
use nand3 g8363
timestamp 1386234893
transform 1 0 10011 0 1 7817
box 0 0 120 799
use inv g8111
timestamp 1386238110
transform 1 0 10131 0 1 7817
box 0 0 120 799
use nand2 g8381
timestamp 1386234792
transform 1 0 10251 0 1 7817
box 0 0 96 799
use inv g8403
timestamp 1386238110
transform 1 0 10347 0 1 7817
box 0 0 120 799
use nand2 g8347
timestamp 1386234792
transform 1 0 10467 0 1 7817
box 0 0 96 799
use nand2 g8357
timestamp 1386234792
transform 1 0 10563 0 1 7817
box 0 0 96 799
use xor2 g8120
timestamp 1386237344
transform 1 0 10659 0 1 7817
box 0 0 192 799
use nand3 g8091
timestamp 1386234893
transform 1 0 10851 0 1 7817
box 0 0 120 799
use nand3 g8134
timestamp 1386234893
transform 1 0 10971 0 1 7817
box 0 0 120 799
use nand2 g8386
timestamp 1386234792
transform 1 0 11091 0 1 7817
box 0 0 96 799
use rowcrosser AluEn
timestamp 1386086759
transform 1 0 11187 0 1 7817
box 0 0 48 799
use nand2 g8320
timestamp 1386234792
transform 1 0 11235 0 1 7817
box 0 0 96 799
use inv g8354
timestamp 1386238110
transform 1 0 11331 0 1 7817
box 0 0 120 799
use nand2 g8374
timestamp 1386234792
transform 1 0 11451 0 1 7817
box 0 0 96 799
use and2 g8050
timestamp 1386234845
transform 1 0 11547 0 1 7817
box 0 0 120 799
use nor2 g8218
timestamp 1386235306
transform 1 0 11667 0 1 7817
box 0 0 120 799
use nand4 g8284
timestamp 1386234936
transform 1 0 11787 0 1 7817
box 0 0 144 799
use nand2 g8198
timestamp 1386234792
transform 1 0 11931 0 1 7817
box 0 0 96 799
use nand2 g8272
timestamp 1386234792
transform 1 0 12027 0 1 7817
box 0 0 96 799
use and2 g8199
timestamp 1386234845
transform 1 0 12123 0 1 7817
box 0 0 120 799
use nand2 g8306
timestamp 1386234792
transform 1 0 12243 0 1 7817
box 0 0 96 799
use rowcrosser RwSel_91_1_93_
timestamp 1386086759
transform 1 0 12339 0 1 7817
box 0 0 48 799
use nand3 g8221
timestamp 1386234893
transform 1 0 12387 0 1 7817
box 0 0 120 799
use nand2 g8319
timestamp 1386234792
transform 1 0 12507 0 1 7817
box 0 0 96 799
use nand2 g8220
timestamp 1386234792
transform 1 0 12603 0 1 7817
box 0 0 96 799
use nand2 g8392
timestamp 1386234792
transform 1 0 12699 0 1 7817
box 0 0 96 799
use nand2 g8194
timestamp 1386234792
transform 1 0 12795 0 1 7817
box 0 0 96 799
use nand2 g8230
timestamp 1386234792
transform 1 0 12891 0 1 7817
box 0 0 96 799
use nor2 g8271
timestamp 1386235306
transform 1 0 12987 0 1 7817
box 0 0 120 799
use nand2 g8340
timestamp 1386234792
transform 1 0 13107 0 1 7817
box 0 0 96 799
use nor2 rm_assigns_buf_StatusReg_1
timestamp 1386235306
transform 1 0 13203 0 1 7817
box 0 0 120 799
use buffer g8399
timestamp 1386236986
transform 1 0 13323 0 1 7817
box 0 0 120 799
use nand2 g8421
timestamp 1386234792
transform 1 0 13443 0 1 7817
box 0 0 96 799
use inv g8074
timestamp 1386238110
transform 1 0 13539 0 1 7817
box 0 0 120 799
use nand4 g8209
timestamp 1386234936
transform 1 0 13659 0 1 7817
box 0 0 144 799
use and2 g8103
timestamp 1386234845
transform 1 0 13803 0 1 7817
box 0 0 120 799
use nor2 g8268
timestamp 1386235306
transform 1 0 13923 0 1 7817
box 0 0 120 799
use inv g8283
timestamp 1386238110
transform 1 0 14043 0 1 7817
box 0 0 120 799
use nand2 g8411
timestamp 1386234792
transform 1 0 14163 0 1 7817
box 0 0 96 799
use nor2 g8321
timestamp 1386235306
transform 1 0 14259 0 1 7817
box 0 0 120 799
use nor2 g8379
timestamp 1386235306
transform 1 0 14379 0 1 7817
box 0 0 120 799
use nor2 g8180
timestamp 1386235306
transform 1 0 14499 0 1 7817
box 0 0 120 799
use nand2 g8052
timestamp 1386234792
transform 1 0 14619 0 1 7817
box 0 0 96 799
use nand4 g8417
timestamp 1386234936
transform 1 0 14715 0 1 7817
box 0 0 144 799
use inv g8136
timestamp 1386238110
transform 1 0 14859 0 1 7817
box 0 0 120 799
use nand2 g8110
timestamp 1386234792
transform 1 0 14979 0 1 7817
box 0 0 96 799
use nand2 g8153
timestamp 1386234792
transform 1 0 15075 0 1 7817
box 0 0 96 799
use nand3 g8361
timestamp 1386234893
transform 1 0 15171 0 1 7817
box 0 0 120 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 15291 0 1 7817
box 0 0 96 799
use scandtype stateSub_reg_91_2_93_
timestamp 1386241841
transform 1 0 15387 0 1 7817
box 0 0 624 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 16011 0 1 7817
box 0 0 48 799
use scandtype g8372
timestamp 1386241841
transform 1 0 16059 0 1 7817
box 0 0 624 799
use inv g8294
timestamp 1386238110
transform 1 0 16683 0 1 7817
box 0 0 120 799
use nand3 g8099
timestamp 1386234893
transform 1 0 16803 0 1 7817
box 0 0 120 799
use nand2 g8057
timestamp 1386234792
transform 1 0 16923 0 1 7817
box 0 0 96 799
use nand4 g8190
timestamp 1386234936
transform 1 0 17019 0 1 7817
box 0 0 144 799
use nand2 g8304
timestamp 1386234792
transform 1 0 17163 0 1 7817
box 0 0 96 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 17259 0 1 7817
box 0 0 48 799
use nand2 g8092
timestamp 1386234792
transform 1 0 17307 0 1 7817
box 0 0 96 799
use nand4 g8277
timestamp 1386234936
transform 1 0 17403 0 1 7817
box 0 0 144 799
use and2 g8081
timestamp 1386234845
transform 1 0 17547 0 1 7817
box 0 0 120 799
use nand2 g8243
timestamp 1386234792
transform 1 0 17667 0 1 7817
box 0 0 96 799
use nand2 g8296
timestamp 1386234792
transform 1 0 17763 0 1 7817
box 0 0 96 799
use nand3 g8348
timestamp 1386234893
transform 1 0 17859 0 1 7817
box 0 0 120 799
use nand2 g8234
timestamp 1386234792
transform 1 0 17979 0 1 7817
box 0 0 96 799
use inv StatusReg_reg_91_1_93_
timestamp 1386238110
transform 1 0 18075 0 1 7817
box 0 0 120 799
use scandtype g8324
timestamp 1386241841
transform 1 0 18195 0 1 7817
box 0 0 624 799
use and2 g8293
timestamp 1386234845
transform 1 0 18819 0 1 7817
box 0 0 120 799
use nand2 g8312
timestamp 1386234792
transform 1 0 18939 0 1 7817
box 0 0 96 799
use inv g8213
timestamp 1386238110
transform 1 0 19035 0 1 7817
box 0 0 120 799
use rowcrosser ALE
timestamp 1386086759
transform 1 0 19155 0 1 7817
box 0 0 48 799
use rowcrosser LrWe
timestamp 1386086759
transform 1 0 19203 0 1 7817
box 0 0 48 799
use nand3 g8096
timestamp 1386234893
transform 1 0 19251 0 1 7817
box 0 0 120 799
use inv g8212
timestamp 1386238110
transform 1 0 19371 0 1 7817
box 0 0 120 799
use nand3 g8084
timestamp 1386234893
transform 1 0 19491 0 1 7817
box 0 0 120 799
use nand3 g8265
timestamp 1386234893
transform 1 0 19611 0 1 7817
box 0 0 120 799
use inv g8200
timestamp 1386238110
transform 1 0 19731 0 1 7817
box 0 0 120 799
use nand2 g8400
timestamp 1386234792
transform 1 0 19851 0 1 7817
box 0 0 96 799
use nand2 g8108
timestamp 1386234792
transform 1 0 19947 0 1 7817
box 0 0 96 799
use nand2 g8049
timestamp 1386234792
transform 1 0 20043 0 1 7817
box 0 0 96 799
use nand4 g8144
timestamp 1386234936
transform 1 0 20139 0 1 7817
box 0 0 144 799
use and2 g8159
timestamp 1386234845
transform 1 0 20283 0 1 7817
box 0 0 120 799
use nand4 g8177
timestamp 1386234936
transform 1 0 20403 0 1 7817
box 0 0 144 799
use nand2 g8356
timestamp 1386234792
transform 1 0 20547 0 1 7817
box 0 0 96 799
use nand3 g8251
timestamp 1386234893
transform 1 0 20643 0 1 7817
box 0 0 120 799
use nand3 g8036
timestamp 1386234893
transform 1 0 20763 0 1 7817
box 0 0 120 799
use nand4 g8226
timestamp 1386234936
transform 1 0 20883 0 1 7817
box 0 0 144 799
use inv g8264
timestamp 1386238110
transform 1 0 21027 0 1 7817
box 0 0 120 799
use nor2 g8332
timestamp 1386235306
transform 1 0 21147 0 1 7817
box 0 0 120 799
use inv g8089
timestamp 1386238110
transform 1 0 21267 0 1 7817
box 0 0 120 799
use and2 g8206
timestamp 1386234845
transform 1 0 21387 0 1 7817
box 0 0 120 799
use nand2 g8237
timestamp 1386234792
transform 1 0 21507 0 1 7817
box 0 0 96 799
use nand2 g8278
timestamp 1386234792
transform 1 0 21603 0 1 7817
box 0 0 96 799
use nand2 g8376
timestamp 1386234792
transform 1 0 21699 0 1 7817
box 0 0 96 799
use nand2 g8181
timestamp 1386234792
transform 1 0 21795 0 1 7817
box 0 0 96 799
use nand2 g8216
timestamp 1386234792
transform 1 0 21891 0 1 7817
box 0 0 96 799
use nand2 StatusReg_reg_91_0_93_
timestamp 1386234792
transform 1 0 21987 0 1 7817
box 0 0 96 799
use scandtype g8253
timestamp 1386241841
transform 1 0 22083 0 1 7817
box 0 0 624 799
use rowcrosser AluWe
timestamp 1386086759
transform 1 0 22707 0 1 7817
box 0 0 48 799
use rowcrosser Rs1Sel_91_0_93_
timestamp 1386086759
transform 1 0 22755 0 1 7817
box 0 0 48 799
use nor2 g8373
timestamp 1386235306
transform 1 0 22803 0 1 7817
box 0 0 120 799
use nand2 g8186
timestamp 1386234792
transform 1 0 22923 0 1 7817
box 0 0 96 799
use inv g8427
timestamp 1386238110
transform 1 0 23019 0 1 7817
box 0 0 120 799
use inv g8090
timestamp 1386238110
transform 1 0 23139 0 1 7817
box 0 0 120 799
use nand3 g8195
timestamp 1386234893
transform 1 0 23259 0 1 7817
box 0 0 120 799
use nand2 g8223
timestamp 1386234792
transform 1 0 23379 0 1 7817
box 0 0 96 799
use and2 g8410
timestamp 1386234845
transform 1 0 23475 0 1 7817
box 0 0 120 799
use and2 g8133
timestamp 1386234845
transform 1 0 23595 0 1 7817
box 0 0 120 799
use nand2 g8341
timestamp 1386234792
transform 1 0 23715 0 1 7817
box 0 0 96 799
use nor2 g8041
timestamp 1386235306
transform 1 0 23811 0 1 7817
box 0 0 120 799
use nand3 g8406
timestamp 1386234893
transform 1 0 23931 0 1 7817
box 0 0 120 799
use nand2 g8289
timestamp 1386234792
transform 1 0 24051 0 1 7817
box 0 0 96 799
use nand2 g8128
timestamp 1386234792
transform 1 0 24147 0 1 7817
box 0 0 96 799
use nand2 g8397
timestamp 1386234792
transform 1 0 24243 0 1 7817
box 0 0 96 799
use and2 g8100
timestamp 1386234845
transform 1 0 24339 0 1 7817
box 0 0 120 799
use nand2 g8350
timestamp 1386234792
transform 1 0 24459 0 1 7817
box 0 0 96 799
use nand2 g8117
timestamp 1386234792
transform 1 0 24555 0 1 7817
box 0 0 96 799
use and2 g8167
timestamp 1386234845
transform 1 0 24651 0 1 7817
box 0 0 120 799
use inv g8191
timestamp 1386238110
transform 1 0 24771 0 1 7817
box 0 0 120 799
use nand2 g8227
timestamp 1386234792
transform 1 0 24891 0 1 7817
box 0 0 96 799
use nand2 g8387
timestamp 1386234792
transform 1 0 24987 0 1 7817
box 0 0 96 799
use inv g8270
timestamp 1386238110
transform 1 0 25083 0 1 7817
box 0 0 120 799
use nand2 g8073
timestamp 1386234792
transform 1 0 25203 0 1 7817
box 0 0 96 799
use nand3 g8163
timestamp 1386234893
transform 1 0 25299 0 1 7817
box 0 0 120 799
use nand3 g8273
timestamp 1386234893
transform 1 0 25419 0 1 7817
box 0 0 120 799
use nor2 g8337
timestamp 1386235306
transform 1 0 25539 0 1 7817
box 0 0 120 799
use nand2 g8051
timestamp 1386234792
transform 1 0 25659 0 1 7817
box 0 0 96 799
use nand2 g8147
timestamp 1386234792
transform 1 0 25755 0 1 7817
box 0 0 96 799
use nand2 g8217
timestamp 1386234792
transform 1 0 25851 0 1 7817
box 0 0 96 799
use nor2 g8353
timestamp 1386235306
transform 1 0 25947 0 1 7817
box 0 0 120 799
use nand2 g8367
timestamp 1386234792
transform 1 0 26067 0 1 7817
box 0 0 96 799
use nand2 g8248
timestamp 1386234792
transform 1 0 26163 0 1 7817
box 0 0 96 799
use nand3 g8114
timestamp 1386234893
transform 1 0 26259 0 1 7817
box 0 0 120 799
use and2 g8174
timestamp 1386234845
transform 1 0 26379 0 1 7817
box 0 0 120 799
use and2 g8393
timestamp 1386234845
transform 1 0 26499 0 1 7817
box 0 0 120 799
use inv g8305
timestamp 1386238110
transform 1 0 26619 0 1 7817
box 0 0 120 799
use nand3 g8241
timestamp 1386234893
transform 1 0 26739 0 1 7817
box 0 0 120 799
use nand3 g8382
timestamp 1386234893
transform 1 0 26859 0 1 7817
box 0 0 120 799
use nand2 g8067
timestamp 1386234792
transform 1 0 26979 0 1 7817
box 0 0 96 799
use nand2 g8158
timestamp 1386234792
transform 1 0 27075 0 1 7817
box 0 0 96 799
use and2 g8063
timestamp 1386234845
transform 1 0 27171 0 1 7817
box 0 0 120 799
use nand2 g8257
timestamp 1386234792
transform 1 0 27291 0 1 7817
box 0 0 96 799
use nand2 PcSel_91_1_93_
timestamp 1386234792
transform 1 0 27387 0 1 7817
box 0 0 96 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 27483 0 1 7817
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27531 0 1 7817
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 912
box 0 0 1464 799
use nand3 stateSub_reg_91_0_93_
timestamp 1386234893
transform 1 0 1587 0 1 912
box 0 0 120 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 1707 0 1 912
box 0 0 48 799
use rowcrosser Flags_91_3_93_
timestamp 1386086759
transform 1 0 1755 0 1 912
box 0 0 48 799
use scandtype g8409
timestamp 1386241841
transform 1 0 1803 0 1 912
box 0 0 624 799
use nand2 g8352
timestamp 1386234792
transform 1 0 2427 0 1 912
box 0 0 96 799
use nor2 g8150
timestamp 1386235306
transform 1 0 2523 0 1 912
box 0 0 120 799
use inv g8178
timestamp 1386238110
transform 1 0 2643 0 1 912
box 0 0 120 799
use nand2 g8250
timestamp 1386234792
transform 1 0 2763 0 1 912
box 0 0 96 799
use nand2 state_reg_91_1_93_
timestamp 1386234792
transform 1 0 2859 0 1 912
box 0 0 96 799
use scandtype g8416
timestamp 1386241841
transform 1 0 2955 0 1 912
box 0 0 624 799
use inv g8148
timestamp 1386238110
transform 1 0 3579 0 1 912
box 0 0 120 799
use nand2 g8196
timestamp 1386234792
transform 1 0 3699 0 1 912
box 0 0 96 799
use nand2 g8211
timestamp 1386234792
transform 1 0 3795 0 1 912
box 0 0 96 799
use nand3 g8300
timestamp 1386234893
transform 1 0 3891 0 1 912
box 0 0 120 799
use inv g8175
timestamp 1386238110
transform 1 0 4011 0 1 912
box 0 0 120 799
use nand3 g8078
timestamp 1386234893
transform 1 0 4131 0 1 912
box 0 0 120 799
use and2 g8388
timestamp 1386234845
transform 1 0 4251 0 1 912
box 0 0 120 799
use nand2 g8093
timestamp 1386234792
transform 1 0 4371 0 1 912
box 0 0 96 799
use nand4 g8104
timestamp 1386234936
transform 1 0 4467 0 1 912
box 0 0 144 799
use nand3 g8391
timestamp 1386234893
transform 1 0 4611 0 1 912
box 0 0 120 799
use nand2 g8307
timestamp 1386234792
transform 1 0 4731 0 1 912
box 0 0 96 799
use nor2 g8389
timestamp 1386235306
transform 1 0 4827 0 1 912
box 0 0 120 799
use nand2 g8335
timestamp 1386234792
transform 1 0 4947 0 1 912
box 0 0 96 799
use nand2 g8160
timestamp 1386234792
transform 1 0 5043 0 1 912
box 0 0 96 799
use nand2 g8076
timestamp 1386234792
transform 1 0 5139 0 1 912
box 0 0 96 799
use nand4 g8224
timestamp 1386234936
transform 1 0 5235 0 1 912
box 0 0 144 799
use nand2 g8161
timestamp 1386234792
transform 1 0 5379 0 1 912
box 0 0 96 799
use nand3 StatusReg_reg_91_2_93_
timestamp 1386234893
transform 1 0 5475 0 1 912
box 0 0 120 799
use scandtype g8094
timestamp 1386241841
transform 1 0 5595 0 1 912
box 0 0 624 799
use mux2 g8121
timestamp 1386235218
transform 1 0 6219 0 1 912
box 0 0 192 799
use nand3 g8037
timestamp 1386234893
transform 1 0 6411 0 1 912
box 0 0 120 799
use nand4 g8266
timestamp 1386234936
transform 1 0 6531 0 1 912
box 0 0 144 799
use nand2 g8401
timestamp 1386234792
transform 1 0 6675 0 1 912
box 0 0 96 799
use nand2 g8189
timestamp 1386234792
transform 1 0 6771 0 1 912
box 0 0 96 799
use inv g8125
timestamp 1386238110
transform 1 0 6867 0 1 912
box 0 0 120 799
use nand2 g8297
timestamp 1386234792
transform 1 0 6987 0 1 912
box 0 0 96 799
use nand2 g8232
timestamp 1386234792
transform 1 0 7083 0 1 912
box 0 0 96 799
use nand2 g8152
timestamp 1386234792
transform 1 0 7179 0 1 912
box 0 0 96 799
use nand3 g8303
timestamp 1386234893
transform 1 0 7275 0 1 912
box 0 0 120 799
use nand2 g8328
timestamp 1386234792
transform 1 0 7395 0 1 912
box 0 0 96 799
use nor2 g8394
timestamp 1386235306
transform 1 0 7491 0 1 912
box 0 0 120 799
use nand2 g8080
timestamp 1386234792
transform 1 0 7611 0 1 912
box 0 0 96 799
use nand4 g8395
timestamp 1386234936
transform 1 0 7707 0 1 912
box 0 0 144 799
use inv g8282
timestamp 1386238110
transform 1 0 7851 0 1 912
box 0 0 120 799
use inv g8267
timestamp 1386238110
transform 1 0 7971 0 1 912
box 0 0 120 799
use nand3 g8274
timestamp 1386234893
transform 1 0 8091 0 1 912
box 0 0 120 799
use nand2 g8236
timestamp 1386234792
transform 1 0 8211 0 1 912
box 0 0 96 799
use nand2 g8101
timestamp 1386234792
transform 1 0 8307 0 1 912
box 0 0 96 799
use nand2 g8349
timestamp 1386234792
transform 1 0 8403 0 1 912
box 0 0 96 799
use inv g8412
timestamp 1386238110
transform 1 0 8499 0 1 912
box 0 0 120 799
use nor2 g8185
timestamp 1386235306
transform 1 0 8619 0 1 912
box 0 0 120 799
use nand2 IntReq_reg
timestamp 1386234792
transform 1 0 8739 0 1 912
box 0 0 96 799
use scandtype g8365
timestamp 1386241841
transform 1 0 8835 0 1 912
box 0 0 624 799
use nand2 g8255
timestamp 1386234792
transform 1 0 9459 0 1 912
box 0 0 96 799
use and2 g8086
timestamp 1386234845
transform 1 0 9555 0 1 912
box 0 0 120 799
use nand2 g8301
timestamp 1386234792
transform 1 0 9675 0 1 912
box 0 0 96 799
use nand2 g8192
timestamp 1386234792
transform 1 0 9771 0 1 912
box 0 0 96 799
use nand2 g8292
timestamp 1386234792
transform 1 0 9867 0 1 912
box 0 0 96 799
use nand2 g8254
timestamp 1386234792
transform 1 0 9963 0 1 912
box 0 0 96 799
use nand2 g8116
timestamp 1386234792
transform 1 0 10059 0 1 912
box 0 0 96 799
use nand2 g8166
timestamp 1386234792
transform 1 0 10155 0 1 912
box 0 0 96 799
use nand4 g8145
timestamp 1386234936
transform 1 0 10251 0 1 912
box 0 0 144 799
use nand2 g8426
timestamp 1386234792
transform 1 0 10395 0 1 912
box 0 0 96 799
use inv g8315
timestamp 1386238110
transform 1 0 10491 0 1 912
box 0 0 120 799
use nor2 g8228
timestamp 1386235306
transform 1 0 10611 0 1 912
box 0 0 120 799
use nand2 g8342
timestamp 1386234792
transform 1 0 10731 0 1 912
box 0 0 96 799
use and2 g8072
timestamp 1386234845
transform 1 0 10827 0 1 912
box 0 0 120 799
use nand4 g8279
timestamp 1386234936
transform 1 0 10947 0 1 912
box 0 0 144 799
use nand2 g8259
timestamp 1386234792
transform 1 0 11091 0 1 912
box 0 0 96 799
use inv g8105
timestamp 1386238110
transform 1 0 11187 0 1 912
box 0 0 120 799
use nand2 g8375
timestamp 1386234792
transform 1 0 11307 0 1 912
box 0 0 96 799
use inv g8129
timestamp 1386238110
transform 1 0 11403 0 1 912
box 0 0 120 799
use nand2 g8122
timestamp 1386234792
transform 1 0 11523 0 1 912
box 0 0 96 799
use nand3 g8059
timestamp 1386234893
transform 1 0 11619 0 1 912
box 0 0 120 799
use nand2 g8062
timestamp 1386234792
transform 1 0 11739 0 1 912
box 0 0 96 799
use nand2 g8097
timestamp 1386234792
transform 1 0 11835 0 1 912
box 0 0 96 799
use nand4 g8025
timestamp 1386234936
transform 1 0 11931 0 1 912
box 0 0 144 799
use nand4 g8247
timestamp 1386234936
transform 1 0 12075 0 1 912
box 0 0 144 799
use nand2 g8263
timestamp 1386234792
transform 1 0 12219 0 1 912
box 0 0 96 799
use nor2 g8256
timestamp 1386235306
transform 1 0 12315 0 1 912
box 0 0 120 799
use nand2 g8131
timestamp 1386234792
transform 1 0 12435 0 1 912
box 0 0 96 799
use nand2 g8087
timestamp 1386234792
transform 1 0 12531 0 1 912
box 0 0 96 799
use nand2 g8345
timestamp 1386234792
transform 1 0 12627 0 1 912
box 0 0 96 799
use nor2 g8322
timestamp 1386235306
transform 1 0 12723 0 1 912
box 0 0 120 799
use inv g8286
timestamp 1386238110
transform 1 0 12843 0 1 912
box 0 0 120 799
use nand3 g8368
timestamp 1386234893
transform 1 0 12963 0 1 912
box 0 0 120 799
use nand2 g8201
timestamp 1386234792
transform 1 0 13083 0 1 912
box 0 0 96 799
use inv g8137
timestamp 1386238110
transform 1 0 13179 0 1 912
box 0 0 120 799
use nand2 g8331
timestamp 1386234792
transform 1 0 13299 0 1 912
box 0 0 96 799
use nand2 g8336
timestamp 1386234792
transform 1 0 13395 0 1 912
box 0 0 96 799
use and2 g8242
timestamp 1386234845
transform 1 0 13491 0 1 912
box 0 0 120 799
use nand2 g8207
timestamp 1386234792
transform 1 0 13611 0 1 912
box 0 0 96 799
use nand2 g8423
timestamp 1386234792
transform 1 0 13707 0 1 912
box 0 0 96 799
use inv g8383
timestamp 1386238110
transform 1 0 13803 0 1 912
box 0 0 120 799
use nand2 g8044
timestamp 1386234792
transform 1 0 13923 0 1 912
box 0 0 96 799
use nand4 g8405
timestamp 1386234936
transform 1 0 14019 0 1 912
box 0 0 144 799
use nand2 g8173
timestamp 1386234792
transform 1 0 14163 0 1 912
box 0 0 96 799
use nand2 g8398
timestamp 1386234792
transform 1 0 14259 0 1 912
box 0 0 96 799
use nand2 g8157
timestamp 1386234792
transform 1 0 14355 0 1 912
box 0 0 96 799
use nand2 g8325
timestamp 1386234792
transform 1 0 14451 0 1 912
box 0 0 96 799
use nand2 g8040
timestamp 1386234792
transform 1 0 14547 0 1 912
box 0 0 96 799
use nand3 g8068
timestamp 1386234893
transform 1 0 14643 0 1 912
box 0 0 120 799
use nand4 g8140
timestamp 1386234936
transform 1 0 14763 0 1 912
box 0 0 144 799
use nand2 g8141
timestamp 1386234792
transform 1 0 14907 0 1 912
box 0 0 96 799
use nor2 g8210
timestamp 1386235306
transform 1 0 15003 0 1 912
box 0 0 120 799
use and2 InISR_reg
timestamp 1386234845
transform 1 0 15123 0 1 912
box 0 0 120 799
use scandtype g8317
timestamp 1386241841
transform 1 0 15243 0 1 912
box 0 0 624 799
use nand2 g8203
timestamp 1386234792
transform 1 0 15867 0 1 912
box 0 0 96 799
use inv g8065
timestamp 1386238110
transform 1 0 15963 0 1 912
box 0 0 120 799
use nand2 g8404
timestamp 1386234792
transform 1 0 16083 0 1 912
box 0 0 96 799
use inv g8413
timestamp 1386238110
transform 1 0 16179 0 1 912
box 0 0 120 799
use nand2 g8113
timestamp 1386234792
transform 1 0 16299 0 1 912
box 0 0 96 799
use nand2 g8358
timestamp 1386234792
transform 1 0 16395 0 1 912
box 0 0 96 799
use nand2 g8070
timestamp 1386234792
transform 1 0 16491 0 1 912
box 0 0 96 799
use inv g8323
timestamp 1386238110
transform 1 0 16587 0 1 912
box 0 0 120 799
use nand2 g8408
timestamp 1386234792
transform 1 0 16707 0 1 912
box 0 0 96 799
use inv g8380
timestamp 1386238110
transform 1 0 16803 0 1 912
box 0 0 120 799
use and2 g8038
timestamp 1386234845
transform 1 0 16923 0 1 912
box 0 0 120 799
use nand4 g8233
timestamp 1386234936
transform 1 0 17043 0 1 912
box 0 0 144 799
use nor2 IRQ2_reg
timestamp 1386235306
transform 1 0 17187 0 1 912
box 0 0 120 799
use scandtype g8151
timestamp 1386241841
transform 1 0 17307 0 1 912
box 0 0 624 799
use nand2 g8138
timestamp 1386234792
transform 1 0 17931 0 1 912
box 0 0 96 799
use nand2 g8402
timestamp 1386234792
transform 1 0 18027 0 1 912
box 0 0 96 799
use inv g8188
timestamp 1386238110
transform 1 0 18123 0 1 912
box 0 0 120 799
use nand2 g8176
timestamp 1386234792
transform 1 0 18243 0 1 912
box 0 0 96 799
use inv g8172
timestamp 1386238110
transform 1 0 18339 0 1 912
box 0 0 120 799
use inv g8422
timestamp 1386238110
transform 1 0 18459 0 1 912
box 0 0 120 799
use inv g8162
timestamp 1386238110
transform 1 0 18579 0 1 912
box 0 0 120 799
use inv g8031
timestamp 1386238110
transform 1 0 18699 0 1 912
box 0 0 120 799
use nand4 g8095
timestamp 1386234936
transform 1 0 18819 0 1 912
box 0 0 144 799
use nand4 g8299
timestamp 1386234936
transform 1 0 18963 0 1 912
box 0 0 144 799
use and2 g8126
timestamp 1386234845
transform 1 0 19107 0 1 912
box 0 0 120 799
use nand2 g8326
timestamp 1386234792
transform 1 0 19227 0 1 912
box 0 0 96 799
use nand2 g8396
timestamp 1386234792
transform 1 0 19323 0 1 912
box 0 0 96 799
use nand2 IRQ1_reg
timestamp 1386234792
transform 1 0 19419 0 1 912
box 0 0 96 799
use scandtype g8329
timestamp 1386241841
transform 1 0 19515 0 1 912
box 0 0 624 799
use nor2 g8205
timestamp 1386235306
transform 1 0 20139 0 1 912
box 0 0 120 799
use nand2 g8339
timestamp 1386234792
transform 1 0 20259 0 1 912
box 0 0 96 799
use and2 g8164
timestamp 1386234845
transform 1 0 20355 0 1 912
box 0 0 120 799
use nand3 g8260
timestamp 1386234893
transform 1 0 20475 0 1 912
box 0 0 120 799
use nor2 g8245
timestamp 1386235306
transform 1 0 20595 0 1 912
box 0 0 120 799
use nand2 g8165
timestamp 1386234792
transform 1 0 20715 0 1 912
box 0 0 96 799
use nand3 g8034
timestamp 1386234893
transform 1 0 20811 0 1 912
box 0 0 120 799
use nand3 g8351
timestamp 1386234893
transform 1 0 20931 0 1 912
box 0 0 120 799
use inv g8215
timestamp 1386238110
transform 1 0 21051 0 1 912
box 0 0 120 799
use nor2 g8343
timestamp 1386235306
transform 1 0 21171 0 1 912
box 0 0 120 799
use nand2 g8288
timestamp 1386234792
transform 1 0 21291 0 1 912
box 0 0 96 799
use inv g8239
timestamp 1386238110
transform 1 0 21387 0 1 912
box 0 0 120 799
use nand2 g8079
timestamp 1386234792
transform 1 0 21507 0 1 912
box 0 0 96 799
use nand2 g8384
timestamp 1386234792
transform 1 0 21603 0 1 912
box 0 0 96 799
use inv g8262
timestamp 1386238110
transform 1 0 21699 0 1 912
box 0 0 120 799
use nand2 g8311
timestamp 1386234792
transform 1 0 21819 0 1 912
box 0 0 96 799
use nand2 g8109
timestamp 1386234792
transform 1 0 21915 0 1 912
box 0 0 96 799
use nand2 g8085
timestamp 1386234792
transform 1 0 22011 0 1 912
box 0 0 96 799
use nand2 g8298
timestamp 1386234792
transform 1 0 22107 0 1 912
box 0 0 96 799
use nand2 g8346
timestamp 1386234792
transform 1 0 22203 0 1 912
box 0 0 96 799
use nand3 g8184
timestamp 1386234893
transform 1 0 22299 0 1 912
box 0 0 120 799
use nand2 g8132
timestamp 1386234792
transform 1 0 22419 0 1 912
box 0 0 96 799
use nand2 g8355
timestamp 1386234792
transform 1 0 22515 0 1 912
box 0 0 96 799
use nand2 g8385
timestamp 1386234792
transform 1 0 22611 0 1 912
box 0 0 96 799
use nand2 g8219
timestamp 1386234792
transform 1 0 22707 0 1 912
box 0 0 96 799
use nand2 g8330
timestamp 1386234792
transform 1 0 22803 0 1 912
box 0 0 96 799
use nand2 g8061
timestamp 1386234792
transform 1 0 22899 0 1 912
box 0 0 96 799
use nand2 g8360
timestamp 1386234792
transform 1 0 22995 0 1 912
box 0 0 96 799
use nor2 g8258
timestamp 1386235306
transform 1 0 23091 0 1 912
box 0 0 120 799
use nand2 g8115
timestamp 1386234792
transform 1 0 23211 0 1 912
box 0 0 96 799
use nand4 g8202
timestamp 1386234936
transform 1 0 23307 0 1 912
box 0 0 144 799
use nand3 g8246
timestamp 1386234893
transform 1 0 23451 0 1 912
box 0 0 120 799
use nand2 g8208
timestamp 1386234792
transform 1 0 23571 0 1 912
box 0 0 96 799
use nand2 g8231
timestamp 1386234792
transform 1 0 23667 0 1 912
box 0 0 96 799
use and2 g8156
timestamp 1386234845
transform 1 0 23763 0 1 912
box 0 0 120 799
use nand4 g8047
timestamp 1386234936
transform 1 0 23883 0 1 912
box 0 0 144 799
use nor2 g8179
timestamp 1386235306
transform 1 0 24027 0 1 912
box 0 0 120 799
use inv g8371
timestamp 1386238110
transform 1 0 24147 0 1 912
box 0 0 120 799
use nand2 g8193
timestamp 1386234792
transform 1 0 24267 0 1 912
box 0 0 96 799
use nand2 g8071
timestamp 1386234792
transform 1 0 24363 0 1 912
box 0 0 96 799
use nand3 g8285
timestamp 1386234893
transform 1 0 24459 0 1 912
box 0 0 120 799
use and2 g8083
timestamp 1386234845
transform 1 0 24579 0 1 912
box 0 0 120 799
use inv g8204
timestamp 1386238110
transform 1 0 24699 0 1 912
box 0 0 120 799
use nand2 g8053
timestamp 1386234792
transform 1 0 24819 0 1 912
box 0 0 96 799
use nand3 state_reg_91_0_93_
timestamp 1386234893
transform 1 0 24915 0 1 912
box 0 0 120 799
use scandtype g8142
timestamp 1386241841
transform 1 0 25035 0 1 912
box 0 0 624 799
use nand2 g8302
timestamp 1386234792
transform 1 0 25659 0 1 912
box 0 0 96 799
use and2 stateSub_reg_91_1_93_
timestamp 1386234845
transform 1 0 25755 0 1 912
box 0 0 120 799
use scandtype g8075
timestamp 1386241841
transform 1 0 25875 0 1 912
box 0 0 624 799
use nand3 g8197
timestamp 1386234893
transform 1 0 26499 0 1 912
box 0 0 120 799
use nand2 g8032
timestamp 1386234792
transform 1 0 26619 0 1 912
box 0 0 96 799
use nor2 g8316
timestamp 1386235306
transform 1 0 26715 0 1 912
box 0 0 120 799
use nand2 Flags_91_0_93_
timestamp 1386234792
transform 1 0 26835 0 1 912
box 0 0 96 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 26931 0 1 912
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27531 0 1 912
box 0 0 320 799
<< labels >>
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 411 9034 423 9034 5 nReset
rlabel metal2 387 9034 399 9034 5 Clock
rlabel metal2 363 9034 375 9034 5 Test
rlabel metal2 339 9034 351 9034 5 SDO
rlabel metal2 123 9034 323 9034 5 Vdd!
rlabel metal2 0 8819 0 8831 4 nWait
rlabel metal2 0 8843 0 8855 4 nME
rlabel metal2 0 8867 0 8879 4 ALE
rlabel metal2 0 4146 0 4158 4 ENB
rlabel metal2 0 4170 0 4182 4 nIRQ
rlabel metal2 0 4194 0 4206 4 nWE
rlabel metal2 0 4218 0 4230 4 nOE
rlabel metal2 0 1 0 13 2 Flags[0]
rlabel metal2 0 25 0 37 2 Flags[2]
rlabel metal2 0 49 0 61 2 Flags[3]
rlabel metal2 0 73 0 85 2 Flags[1]
rlabel metal2 27651 0 27851 0 1 GND!
rlabel metal2 28047 1 28047 13 8 OpcodeCondIn[5]
rlabel metal2 28047 25 28047 37 8 OpcodeCondIn[4]
rlabel metal2 28047 49 28047 61 8 OpcodeCondIn[6]
rlabel metal2 28047 73 28047 85 8 OpcodeCondIn[7]
rlabel metal2 28047 97 28047 109 8 OpcodeCondIn[2]
rlabel metal2 28047 145 28047 157 8 OpcodeCondIn[0]
rlabel metal2 28047 3858 28047 3870 6 SysBus[1]
rlabel metal2 28047 5226 28047 5238 6 AluOR[1]
rlabel metal2 28047 1722 28047 1734 6 OpcodeCondIn[1]
rlabel metal2 28047 1746 28047 1758 6 OpcodeCondIn[3]
rlabel metal2 28047 1770 28047 1782 6 SysBus[2]
rlabel metal2 28047 1794 28047 1806 6 SysBus[3]
rlabel metal2 28047 1818 28047 1830 6 SysBus[0]
rlabel metal2 27651 9034 27850 9034 5 GND!
rlabel metal2 28047 8627 28047 8639 6 AluOR[0]
rlabel metal2 28047 8651 28047 8663 6 Rs1Sel[0]
rlabel metal2 28047 8675 28047 8687 6 RwSel[1]
rlabel metal2 28047 8699 28047 8711 6 Rs1Sel[1]
rlabel metal2 28047 8723 28047 8735 6 RwSel[0]
rlabel metal2 28047 8747 28047 8759 6 RegWe
rlabel metal2 28047 8771 28047 8783 6 CFlag
rlabel metal2 2391 9034 2403 9034 4 AluEn
rlabel metal2 3951 9034 3963 9034 4 AluWe
rlabel metal2 6171 9034 6183 9034 4 Op2Sel[1]
rlabel metal2 7707 9034 7719 9034 4 Op2Sel[0]
rlabel metal2 9243 9034 9255 9034 4 ImmSel
rlabel metal2 10779 9034 10791 9034 4 Op1Sel
rlabel metal2 12315 9034 12327 9034 4 PcWe
rlabel metal2 13851 9034 13863 9034 4 PcEn
rlabel metal2 15387 9034 15399 9034 6 PcSel[2]
rlabel metal2 16047 9034 16059 9034 6 PcSel[1]
rlabel metal2 16935 9034 16947 9034 6 PcSel[0]
rlabel metal2 18459 9034 18471 9034 6 LrEn
rlabel metal2 19983 9034 19995 9034 6 WdSel
rlabel metal2 22743 9034 22755 9034 6 LrWe
rlabel metal2 23031 9034 23043 9034 6 LrSel
rlabel metal2 24555 9034 24567 9034 6 IrWe
rlabel metal2 26079 9034 26091 9034 6 MemEn
rlabel m2contact 1737 55 1737 55 2 Flags[3]
rlabel m2contact 1785 79 1785 79 2 Flags[1]
rlabel m2contact 2481 55 2481 55 2 OpcodeCondIn[6]
rlabel m2contact 2721 79 2721 79 2 n_283
rlabel m2contact 2841 103 2841 103 2 n_216
rlabel m2contact 2889 127 2889 127 2 n_120
rlabel m2contact 3609 151 3609 151 2 OpcodeCondIn[0]
rlabel m2contact 3993 175 3993 175 2 n_192
rlabel m2contact 4041 127 4041 127 2 n_120
rlabel m2contact 4233 199 4233 199 2 n_187
rlabel m2contact 4281 223 4281 223 2 n_238
rlabel m2contact 4353 247 4353 247 2 n_291
rlabel m2contact 4497 271 4497 271 2 n_9
rlabel m2contact 4785 295 4785 295 2 OpcodeCondIn[5]
rlabel m2contact 5025 319 5025 319 2 n_16
rlabel m2contact 5073 319 5073 319 2 n_16
rlabel m2contact 5169 175 5169 175 2 n_192
rlabel m2contact 5217 175 5217 175 2 n_249
rlabel m2contact 5577 319 5577 319 2 n_228
rlabel m2contact 6273 343 6273 343 2 OpcodeCondIn[4]
rlabel m2contact 6345 175 6345 175 2 n_249
rlabel m2contact 6513 175 6513 175 2 n_204
rlabel m2contact 6585 247 6585 247 2 n_291
rlabel m2contact 6849 247 6849 247 2 n_8
rlabel m2contact 7041 367 7041 367 2 n_113
rlabel m2contact 7161 391 7161 391 2 n_93
rlabel m2contact 7425 415 7425 415 2 n_48
rlabel m2contact 7785 439 7785 439 2 n_270
rlabel m2contact 8145 463 8145 463 2 n_14
rlabel m2contact 8289 487 8289 487 2 n_125
rlabel m2contact 8433 511 8433 511 2 n_235
rlabel m2contact 8793 535 8793 535 2 n_145
rlabel m2contact 8817 559 8817 559 2 n_183
rlabel m2contact 9849 127 9849 127 2 n_120
rlabel m2contact 9945 127 9945 127 2 n_211
rlabel m2contact 10089 583 10089 583 2 n_505
rlabel m2contact 10113 607 10113 607 2 IRQ2
rlabel m2contact 10233 631 10233 631 2 n_302
rlabel m2contact 10353 655 10353 655 2 OpcodeCondIn[2]
rlabel m2contact 10377 679 10377 679 2 n_223
rlabel m2contact 10521 295 10521 295 2 OpcodeCondIn[5]
rlabel m2contact 10761 391 10761 391 2 n_93
rlabel m2contact 11145 655 11145 655 2 OpcodeCondIn[2]
rlabel m2contact 11217 391 11217 391 2 n_134
rlabel m2contact 11265 703 11265 703 2 n_150
rlabel m2contact 11361 679 11361 679 2 n_223
rlabel m2contact 11673 559 11673 559 2 n_183
rlabel m2contact 11697 55 11697 55 2 OpcodeCondIn[6]
rlabel m2contact 11721 559 11721 559 2 n_260
rlabel m2contact 11817 679 11817 679 2 n_361
rlabel m2contact 12153 727 12153 727 2 n_393
rlabel m2contact 12465 751 12465 751 2 n_37
rlabel m2contact 12513 367 12513 367 2 n_113
rlabel m2contact 12561 367 12561 367 2 n_244
rlabel m2contact 12657 631 12657 631 2 n_302
rlabel m2contact 12705 631 12705 631 2 n_332
rlabel m2contact 13209 775 13209 775 2 n_181
rlabel m2contact 13353 295 13353 295 2 OpcodeCondIn[5]
rlabel m2contact 13377 799 13377 799 4 n_298
rlabel m2contact 13473 823 13473 823 4 n_44
rlabel m2contact 13545 151 13545 151 2 OpcodeCondIn[0]
rlabel m2contact 13785 847 13785 847 4 n_167
rlabel m2contact 13833 343 13833 343 2 OpcodeCondIn[4]
rlabel m2contact 13977 871 13977 871 4 OpcodeCondIn[7]
rlabel m2contact 14049 895 14049 895 4 n_66
rlabel m2contact 14073 823 14073 823 4 n_44
rlabel m2contact 14097 631 14097 631 2 n_332
rlabel m2contact 14145 631 14145 631 2 n_376
rlabel m2contact 14193 295 14193 295 2 OpcodeCondIn[5]
rlabel m2contact 14217 55 14217 55 2 OpcodeCondIn[6]
rlabel m2contact 14625 895 14625 895 6 n_66
rlabel m2contact 14697 679 14697 679 8 n_361
rlabel m2contact 14817 679 14817 679 8 n_288
rlabel m2contact 14841 79 14841 79 8 n_283
rlabel m2contact 14937 103 14937 103 8 n_216
rlabel m2contact 15177 823 15177 823 6 n_201
rlabel m2contact 15225 439 15225 439 8 n_270
rlabel m2contact 15705 583 15705 583 8 n_505
rlabel m2contact 15945 751 15945 751 8 n_37
rlabel m2contact 16137 31 16137 31 8 Flags[2]
rlabel m2contact 16353 655 16353 655 8 OpcodeCondIn[2]
rlabel m2contact 16425 583 16425 583 8 n_254
rlabel m2contact 16473 751 16473 751 8 n_303
rlabel m2contact 16569 415 16569 415 8 n_48
rlabel m2contact 16617 895 16617 895 6 n_314
rlabel m2contact 16881 463 16881 463 8 n_14
rlabel m2contact 17409 463 17409 463 8 IRQ1
rlabel m2contact 17769 439 17769 439 8 n_504
rlabel m2contact 17817 607 17817 607 8 IRQ2
rlabel m2contact 18057 847 18057 847 6 n_167
rlabel m2contact 18417 367 18417 367 8 n_244
rlabel m2contact 18609 55 18609 55 8 OpcodeCondIn[6]
rlabel m2contact 18993 319 18993 319 8 n_228
rlabel m2contact 19041 799 19041 799 6 n_298
rlabel m2contact 19065 127 19065 127 8 n_211
rlabel m2contact 19257 199 19257 199 8 n_187
rlabel m2contact 19305 511 19305 511 8 n_235
rlabel m2contact 20025 463 20025 463 8 IRQ1
rlabel m2contact 20409 343 20409 343 8 OpcodeCondIn[4]
rlabel m2contact 20457 511 20457 511 8 n_57
rlabel m2contact 20553 295 20553 295 8 OpcodeCondIn[5]
rlabel m2contact 20697 391 20697 391 8 n_134
rlabel m2contact 20769 871 20769 871 6 OpcodeCondIn[7]
rlabel m2contact 20793 535 20793 535 8 n_145
rlabel m2contact 21657 175 21657 175 8 n_204
rlabel m2contact 21681 535 21681 535 8 n_258
rlabel m2contact 22137 751 22137 751 8 n_303
rlabel m2contact 22161 607 22161 607 8 n_143
rlabel m2contact 22233 463 22233 463 8 IRQ1
rlabel m2contact 22257 439 22257 439 8 n_504
rlabel m2contact 22377 871 22377 871 6 OpcodeCondIn[7]
rlabel m2contact 22401 271 22401 271 8 n_9
rlabel m2contact 22593 679 22593 679 8 n_288
rlabel m2contact 22761 295 22761 295 8 OpcodeCondIn[5]
rlabel m2contact 22833 703 22833 703 8 n_150
rlabel m2contact 22857 871 22857 871 6 OpcodeCondIn[7]
rlabel m2contact 22881 823 22881 823 6 n_201
rlabel m2contact 23289 463 23289 463 8 n_136
rlabel m2contact 23433 223 23433 223 8 n_238
rlabel m2contact 23553 775 23553 775 8 n_181
rlabel m2contact 23649 607 23649 607 8 n_143
rlabel m2contact 23817 871 23817 871 6 OpcodeCondIn[7]
rlabel m2contact 24321 151 24321 151 8 OpcodeCondIn[0]
rlabel m2contact 24489 463 24489 463 8 n_136
rlabel m2contact 24513 559 24513 559 8 n_260
rlabel m2contact 24537 247 24537 247 8 n_8
rlabel m2contact 24561 895 24561 895 6 n_314
rlabel m2contact 24633 871 24633 871 6 OpcodeCondIn[7]
rlabel m2contact 24945 487 24945 487 8 n_125
rlabel m2contact 24993 535 24993 535 8 n_258
rlabel m2contact 25017 463 25017 463 8 n_310
rlabel m2contact 25137 463 25137 463 8 n_310
rlabel m2contact 25737 583 25737 583 8 n_254
rlabel m2contact 25977 631 25977 631 8 n_376
rlabel m2contact 26769 511 26769 511 8 n_57
rlabel m2contact 26817 727 26817 727 8 n_393
rlabel m2contact 26961 7 26961 7 8 Flags[0]
rlabel m2contact 26985 7 26985 7 8 OpcodeCondIn[5]
rlabel m2contact 26985 295 26985 295 8 OpcodeCondIn[5]
rlabel m2contact 27009 31 27009 31 8 OpcodeCondIn[4]
rlabel m2contact 27009 343 27009 343 8 OpcodeCondIn[4]
rlabel m2contact 27033 79 27033 79 8 OpcodeCondIn[7]
rlabel m2contact 27033 871 27033 871 6 OpcodeCondIn[7]
rlabel m2contact 27057 103 27057 103 8 OpcodeCondIn[2]
rlabel m2contact 27057 655 27057 655 8 OpcodeCondIn[2]
rlabel m2contact 1617 4248 1617 4248 4 n_43
rlabel m2contact 1617 4128 1617 4128 4 n_384
rlabel m2contact 1641 4272 1641 4272 4 n_343
rlabel m2contact 1665 4296 1665 4296 4 n_220
rlabel m2contact 1665 4320 1665 4320 4 n_18
rlabel m2contact 1689 4224 1689 4224 4 nOE
rlabel m2contact 1737 4224 1737 4224 4 Flags[3]
rlabel m2contact 1737 4344 1737 4344 4 OpcodeCondIn[1]
rlabel m2contact 1761 4368 1761 4368 4 OpcodeCondIn[0]
rlabel m2contact 1785 4392 1785 4392 4 Flags[1]
rlabel m2contact 1809 4416 1809 4416 4 n_140
rlabel m2contact 1857 4440 1857 4440 4 n_377
rlabel m2contact 1881 4104 1881 4104 4 n_357
rlabel m2contact 1905 4464 1905 4464 4 n_247
rlabel m2contact 1905 4488 1905 4488 4 n_320
rlabel m2contact 1929 4512 1929 4512 4 n_391
rlabel m2contact 1977 4536 1977 4536 4 n_95
rlabel m2contact 2001 4560 2001 4560 4 n_118
rlabel m2contact 2097 4080 2097 4080 4 n_255
rlabel m2contact 2121 4584 2121 4584 4 n_227
rlabel m2contact 2145 4608 2145 4608 4 n_304
rlabel m2contact 2193 4632 2193 4632 4 n_359
rlabel m2contact 2241 4656 2241 4656 4 n_360
rlabel m2contact 2265 4056 2265 4056 4 n_19
rlabel m2contact 2289 4680 2289 4680 4 n_87
rlabel m2contact 2313 4032 2313 4032 4 stateSub[0]
rlabel m2contact 2313 4704 2313 4704 4 state[0]
rlabel m2contact 2337 4728 2337 4728 4 n_149
rlabel m2contact 2385 4008 2385 4008 4 AluEn
rlabel m2contact 2433 4752 2433 4752 4 n_11
rlabel m2contact 2457 4704 2457 4704 4 state[0]
rlabel m2contact 2457 4776 2457 4776 4 OpcodeCondIn[7]
rlabel m2contact 2481 3984 2481 3984 4 n_21
rlabel m2contact 2505 3960 2505 3960 4 n_13
rlabel m2contact 2529 4800 2529 4800 4 n_379
rlabel m2contact 2553 4224 2553 4224 4 Flags[3]
rlabel m2contact 2553 3936 2553 3936 4 n_49
rlabel m2contact 2577 4440 2577 4440 4 n_377
rlabel m2contact 2577 3912 2577 3912 4 n_112
rlabel m2contact 2625 4224 2625 4224 4 n_153
rlabel m2contact 2625 4440 2625 4440 4 n_373
rlabel m2contact 2673 3888 2673 3888 4 n_282
rlabel m2contact 2673 4824 2673 4824 4 n_299
rlabel m2contact 2745 4848 2745 4848 4 n_322
rlabel m2contact 2769 3864 2769 3864 4 SysBus[1]
rlabel m2contact 2793 3840 2793 3840 4 n_213
rlabel m2contact 2793 4872 2793 4872 4 n_323
rlabel m2contact 2817 3816 2817 3816 4 n_237
rlabel m2contact 2841 3792 2841 3792 4 n_117
rlabel m2contact 2865 3768 2865 3768 4 n_34
rlabel m2contact 2913 3744 2913 3744 4 state[1]
rlabel m2contact 2913 4896 2913 4896 4 n_158
rlabel m2contact 2937 4920 2937 4920 4 n_151
rlabel m2contact 2961 4944 2961 4944 4 n_53
rlabel m2contact 3009 4968 3009 4968 4 n_98
rlabel m2contact 3057 4992 3057 4992 4 n_292
rlabel m2contact 3081 4248 3081 4248 4 n_43
rlabel m2contact 3105 5016 3105 5016 4 n_172
rlabel m2contact 3153 5040 3153 5040 4 n_74
rlabel m2contact 3201 3720 3201 3720 4 n_363
rlabel m2contact 3225 5064 3225 5064 4 n_382
rlabel m2contact 3297 4248 3297 4248 4 n_43
rlabel m2contact 3321 5088 3321 5088 4 n_232
rlabel m2contact 3345 3696 3345 3696 4 n_89
rlabel m2contact 3393 5112 3393 5112 4 n_83
rlabel m2contact 3417 3672 3417 3672 4 n_218
rlabel m2contact 3417 5136 3417 5136 4 n_91
rlabel m2contact 3465 4128 3465 4128 4 n_384
rlabel m2contact 3465 3744 3465 3744 4 state[1]
rlabel m2contact 3513 5160 3513 5160 4 n_234
rlabel m2contact 3537 5184 3537 5184 4 n_20
rlabel m2contact 3585 5208 3585 5208 4 n_273
rlabel m2contact 3609 4368 3609 4368 4 OpcodeCondIn[0]
rlabel m2contact 3633 5232 3633 5232 4 n_341
rlabel m2contact 3657 3648 3657 3648 4 n_12
rlabel m2contact 3729 5256 3729 5256 4 n_239
rlabel m2contact 3753 4032 3753 4032 4 stateSub[0]
rlabel m2contact 3753 3624 3753 3624 4 n_240
rlabel m2contact 3777 5280 3777 5280 4 n_285
rlabel m2contact 3777 5304 3777 5304 4 n_31
rlabel m2contact 3801 5328 3801 5328 4 n_39
rlabel m2contact 3825 3600 3825 3600 4 n_191
rlabel m2contact 3849 5352 3849 5352 4 n_142
rlabel m2contact 3849 5376 3849 5376 4 n_219
rlabel m2contact 3873 5400 3873 5400 4 n_182
rlabel m2contact 3873 5424 3873 5424 4 n_7
rlabel m2contact 3897 3576 3897 3576 4 n_35
rlabel m2contact 3921 4968 3921 4968 4 n_98
rlabel m2contact 3945 3600 3945 3600 4 n_191
rlabel m2contact 3945 5448 3945 5448 4 AluWe
rlabel m2contact 3969 3816 3969 3816 4 n_237
rlabel m2contact 3993 5472 3993 5472 4 n_261
rlabel m2contact 4017 5496 4017 5496 4 OpcodeCondIn[3]
rlabel m2contact 4041 5520 4041 5520 4 n_269
rlabel m2contact 4089 5544 4089 5544 4 n_121
rlabel m2contact 4089 5568 4089 5568 4 n_311
rlabel m2contact 4161 3552 4161 3552 4 n_222
rlabel m2contact 4185 5016 4185 5016 4 n_172
rlabel m2contact 4209 3528 4209 3528 4 n_186
rlabel m2contact 4209 5592 4209 5592 4 n_230
rlabel m2contact 4233 5376 4233 5376 4 n_219
rlabel m2contact 4257 4296 4257 4296 4 n_220
rlabel m2contact 4305 3528 4305 3528 4 n_186
rlabel m2contact 4305 3504 4305 3504 4 n_215
rlabel m2contact 4329 4296 4329 4296 4 n_81
rlabel m2contact 4353 5616 4353 5616 4 OpcodeCondIn[6]
rlabel m2contact 4377 5640 4377 5640 4 n_82
rlabel m2contact 4401 3816 4401 3816 4 n_237
rlabel m2contact 4425 4344 4425 4344 4 OpcodeCondIn[1]
rlabel m2contact 4425 5664 4425 5664 4 n_38
rlabel m2contact 4449 4224 4449 4224 4 n_153
rlabel m2contact 4449 3480 4449 3480 4 n_27
rlabel m2contact 4473 3456 4473 3456 4 n_97
rlabel m2contact 4521 5688 4521 5688 4 n_148
rlabel m2contact 4521 3432 4521 3432 4 n_25
rlabel m2contact 4545 4704 4545 4704 4 state[0]
rlabel m2contact 4545 3408 4545 3408 4 n_199
rlabel m2contact 4569 5712 4569 5712 4 n_168
rlabel m2contact 4569 3384 4569 3384 4 n_280
rlabel m2contact 4593 5736 4593 5736 4 n_281
rlabel m2contact 4617 5760 4617 5760 4 n_130
rlabel m2contact 4641 3360 4641 3360 4 n_70
rlabel m2contact 4665 3552 4665 3552 4 n_222
rlabel m2contact 4665 3336 4665 3336 4 n_306
rlabel m2contact 4689 3648 4689 3648 4 n_12
rlabel m2contact 4713 3312 4713 3312 4 n_352
rlabel m2contact 4737 5784 4737 5784 4 n_106
rlabel m2contact 4761 3288 4761 3288 4 n_110
rlabel m2contact 4761 5808 4761 5808 4 n_276
rlabel m2contact 4785 5832 4785 5832 4 n_346
rlabel m2contact 4809 3264 4809 3264 4 n_26
rlabel m2contact 4833 4824 4833 4824 4 n_299
rlabel m2contact 4857 3240 4857 3240 4 StatusReg[0]
rlabel m2contact 4857 5856 4857 5856 4 n_217
rlabel m2contact 4881 5880 4881 5880 4 n_300
rlabel m2contact 4881 3216 4881 3216 4 n_54
rlabel m2contact 4929 5904 4929 5904 4 n_327
rlabel m2contact 4929 3192 4929 3192 4 n_41
rlabel m2contact 4953 5832 4953 5832 4 n_346
rlabel m2contact 4977 4704 4977 4704 4 state[0]
rlabel m2contact 4977 5928 4977 5928 4 n_347
rlabel m2contact 5001 4056 5001 4056 4 n_19
rlabel m2contact 5025 5952 5025 5952 4 n_71
rlabel m2contact 5049 5856 5049 5856 4 n_217
rlabel m2contact 5073 5976 5073 5976 4 n_72
rlabel m2contact 5097 3168 5097 3168 4 n_193
rlabel m2contact 5121 3648 5121 3648 4 n_12
rlabel m2contact 5121 3144 5121 3144 4 n_61
rlabel m2contact 5145 4344 5145 4344 4 OpcodeCondIn[1]
rlabel m2contact 5169 3216 5169 3216 4 n_54
rlabel m2contact 5193 3120 5193 3120 4 n_198
rlabel m2contact 5217 3264 5217 3264 4 n_26
rlabel m2contact 5265 6000 5265 6000 4 n_328
rlabel m2contact 5265 6024 5265 6024 4 n_63
rlabel m2contact 5289 3696 5289 3696 4 n_89
rlabel m2contact 5313 6048 5313 6048 4 n_109
rlabel m2contact 5337 3696 5337 3696 4 n_365
rlabel m2contact 5337 6072 5337 6072 4 n_163
rlabel m2contact 5361 6096 5361 6096 4 n_366
rlabel m2contact 5361 6120 5361 6120 4 n_139
rlabel m2contact 5409 6144 5409 6144 4 n_221
rlabel m2contact 5409 3096 5409 3096 4 n_100
rlabel m2contact 5433 6168 5433 6168 4 n_128
rlabel m2contact 5457 6192 5457 6192 4 n_177
rlabel m2contact 5457 6216 5457 6216 4 n_196
rlabel m2contact 5481 6240 5481 6240 4 n_195
rlabel m2contact 5505 4584 5505 4584 4 n_227
rlabel m2contact 5505 6264 5505 6264 4 n_197
rlabel m2contact 5529 3072 5529 3072 4 n_225
rlabel m2contact 5553 6288 5553 6288 4 n_51
rlabel m2contact 5553 6312 5553 6312 4 n_159
rlabel m2contact 5577 5760 5577 5760 4 n_130
rlabel m2contact 5625 3072 5625 3072 4 n_225
rlabel m2contact 5673 3048 5673 3048 4 n_185
rlabel m2contact 5697 4296 5697 4296 4 n_81
rlabel m2contact 5697 3024 5697 3024 4 n_392
rlabel m2contact 5745 5160 5745 5160 4 n_234
rlabel m2contact 5793 4248 5793 4248 4 n_43
rlabel m2contact 5817 3672 5817 3672 4 n_218
rlabel m2contact 5841 5160 5841 5160 4 n_253
rlabel m2contact 5889 5520 5889 5520 4 n_269
rlabel m2contact 5913 6336 5913 6336 4 n_203
rlabel m2contact 5961 6360 5961 6360 4 n_284
rlabel m2contact 6009 3000 6009 3000 4 n_378
rlabel m2contact 6033 2976 6033 2976 4 n_358
rlabel m2contact 6057 6384 6057 6384 4 n_321
rlabel m2contact 6057 2952 6057 2952 4 n_506
rlabel m2contact 6081 3024 6081 3024 4 n_392
rlabel m2contact 6105 2928 6105 2928 4 StatusReg[2]
rlabel m2contact 6129 5280 6129 5280 4 n_285
rlabel m2contact 6153 3024 6153 3024 4 n_264
rlabel m2contact 6177 5280 6177 5280 4 n_316
rlabel m2contact 6201 6408 6201 6408 4 n_339
rlabel m2contact 6225 2904 6225 2904 4 n_340
rlabel m2contact 6273 6432 6273 6432 4 n_86
rlabel m2contact 6297 5472 6297 5472 4 n_261
rlabel m2contact 6297 6456 6297 6456 4 n_58
rlabel m2contact 6345 6480 6345 6480 4 n_132
rlabel m2contact 6369 6504 6369 6504 4 n_309
rlabel m2contact 6393 3144 6393 3144 4 n_61
rlabel m2contact 6417 6528 6417 6528 4 n_30
rlabel m2contact 6441 6336 6441 6336 4 n_203
rlabel m2contact 6441 6552 6441 6552 4 n_103
rlabel m2contact 6465 3144 6465 3144 4 n_202
rlabel m2contact 6489 3456 6489 3456 4 n_97
rlabel m2contact 6489 6576 6489 6576 4 n_40
rlabel m2contact 6513 6600 6513 6600 4 n_60
rlabel m2contact 6537 3456 6537 3456 4 n_28
rlabel m2contact 6561 5064 6561 5064 4 n_382
rlabel m2contact 6561 5352 6561 5352 4 n_142
rlabel m2contact 6609 4800 6609 4800 4 n_379
rlabel m2contact 6609 2880 6609 2880 4 n_386
rlabel m2contact 6633 4392 6633 4392 4 Flags[1]
rlabel m2contact 6633 2856 6633 2856 4 n_346
rlabel m2contact 6657 5448 6657 5448 4 AluWe
rlabel m2contact 6657 6624 6657 6624 4 n_380
rlabel m2contact 6681 2856 6681 2856 4 n_346
rlabel m2contact 6681 5832 6681 5832 4 n_346
rlabel m2contact 6705 4224 6705 4224 4 n_153
rlabel m2contact 6705 5352 6705 5352 4 n_75
rlabel m2contact 6729 3288 6729 3288 4 n_110
rlabel m2contact 6729 5448 6729 5448 4 n_32
rlabel m2contact 6753 4392 6753 4392 4 n_157
rlabel m2contact 6777 2856 6777 2856 4 n_76
rlabel m2contact 6801 2832 6801 2832 4 stateSub[1]
rlabel m2contact 6825 3600 6825 3600 4 n_191
rlabel m2contact 6825 2808 6825 2808 4 n_10
rlabel m2contact 6849 5496 6849 5496 4 OpcodeCondIn[3]
rlabel m2contact 6873 3120 6873 3120 4 n_198
rlabel m2contact 6897 2784 6897 2784 4 n_268
rlabel m2contact 6921 6504 6921 6504 4 n_309
rlabel m2contact 6945 3336 6945 3336 4 n_306
rlabel m2contact 6945 6648 6945 6648 4 n_59
rlabel m2contact 6969 6504 6969 6504 4 n_362
rlabel m2contact 7017 4824 7017 4824 4 n_299
rlabel m2contact 7017 6672 7017 6672 4 StatusReg[2]
rlabel m2contact 7041 2928 7041 2928 4 StatusReg[2]
rlabel m2contact 7041 6672 7041 6672 4 StatusReg[2]
rlabel m2contact 7041 6696 7041 6696 4 n_507
rlabel m2contact 7065 6720 7065 6720 4 n_301
rlabel m2contact 7065 6744 7065 6744 4 n_47
rlabel m2contact 7113 3624 7113 3624 4 n_240
rlabel m2contact 7113 5736 7113 5736 4 n_281
rlabel m2contact 7137 4224 7137 4224 4 n_153
rlabel m2contact 7137 6672 7137 6672 4 n_135
rlabel m2contact 7185 5736 7185 5736 4 n_308
rlabel m2contact 7209 2760 7209 2760 4 n_155
rlabel m2contact 7233 3312 7233 3312 4 n_352
rlabel m2contact 7233 2736 7233 2736 4 n_170
rlabel m2contact 7257 6768 7257 6768 4 n_188
rlabel m2contact 7257 2712 7257 2712 4 n_156
rlabel m2contact 7305 5376 7305 5376 4 n_219
rlabel m2contact 7329 5592 7329 5592 4 n_230
rlabel m2contact 7329 6792 7329 6792 4 n_33
rlabel m2contact 7353 2688 7353 2688 4 n_224
rlabel m2contact 7353 6816 7353 6816 4 n_85
rlabel m2contact 7377 6840 7377 6840 4 n_78
rlabel m2contact 7377 2664 7377 2664 4 n_231
rlabel m2contact 7401 5328 7401 5328 4 n_39
rlabel m2contact 7425 6864 7425 6864 4 n_164
rlabel m2contact 7449 4416 7449 4416 4 n_140
rlabel m2contact 7473 3792 7473 3792 4 n_117
rlabel m2contact 7473 5328 7473 5328 4 n_344
rlabel m2contact 7497 6888 7497 6888 4 n_294
rlabel m2contact 7521 3792 7521 3792 4 n_56
rlabel m2contact 7545 2832 7545 2832 4 stateSub[1]
rlabel m2contact 7545 6912 7545 6912 4 n_370
rlabel m2contact 7593 6936 7593 6936 4 n_174
rlabel m2contact 7617 3624 7617 3624 4 n_240
rlabel m2contact 7641 5376 7641 5376 4 n_219
rlabel m2contact 7641 6960 7641 6960 4 n_102
rlabel m2contact 7665 4032 7665 4032 4 stateSub[0]
rlabel m2contact 7689 5304 7689 5304 4 n_31
rlabel m2contact 7689 2640 7689 2640 4 n_159
rlabel m2contact 7713 2640 7713 2640 4 n_159
rlabel m2contact 7713 6312 7713 6312 4 n_159
rlabel m2contact 7737 5448 7737 5448 4 n_32
rlabel m2contact 7737 2616 7737 2616 4 n_124
rlabel m2contact 7761 2640 7761 2640 4 n_205
rlabel m2contact 7809 5376 7809 5376 4 n_219
rlabel m2contact 7809 3144 7809 3144 4 n_202
rlabel m2contact 7833 4632 7833 4632 4 n_359
rlabel m2contact 7833 5448 7833 5448 4 n_170
rlabel m2contact 7857 2736 7857 2736 4 n_170
rlabel m2contact 7857 5448 7857 5448 4 n_170
rlabel m2contact 7857 6984 7857 6984 4 n_126
rlabel m2contact 7881 2592 7881 2592 4 n_52
rlabel m2contact 7905 3840 7905 3840 4 n_213
rlabel m2contact 7929 5088 7929 5088 4 n_232
rlabel m2contact 7929 5448 7929 5448 4 n_218
rlabel m2contact 7953 3672 7953 3672 4 n_218
rlabel m2contact 7953 5448 7953 5448 4 n_218
rlabel m2contact 7953 7008 7953 7008 4 n_214
rlabel m2contact 8001 5472 8001 5472 4 n_261
rlabel m2contact 8001 5448 8001 5448 4 n_203
rlabel m2contact 8025 3912 8025 3912 4 n_112
rlabel m2contact 8049 4440 8049 4440 4 n_373
rlabel m2contact 8049 2568 8049 2568 4 n_195
rlabel m2contact 8073 5448 8073 5448 4 n_203
rlabel m2contact 8073 6336 8073 6336 4 n_203
rlabel m2contact 8097 6864 8097 6864 4 n_164
rlabel m2contact 8121 5376 8121 5376 4 n_219
rlabel m2contact 8121 5448 8121 5448 4 n_73
rlabel m2contact 8145 2568 8145 2568 4 n_195
rlabel m2contact 8145 6240 8145 6240 4 n_195
rlabel m2contact 8169 3984 8169 3984 4 n_21
rlabel m2contact 8169 6864 8169 6864 4 n_199
rlabel m2contact 8193 6816 8193 6816 4 n_85
rlabel m2contact 8217 4848 8217 4848 4 n_322
rlabel m2contact 8241 6816 8241 6816 4 SysBus[0]
rlabel m2contact 8241 3984 8241 3984 4 n_62
rlabel m2contact 8265 4704 8265 4704 4 state[0]
rlabel m2contact 8265 7032 8265 7032 4 n_324
rlabel m2contact 8289 3408 8289 3408 4 n_199
rlabel m2contact 8289 6864 8289 6864 4 n_199
rlabel m2contact 8313 4176 8313 4176 4 nIRQ
rlabel m2contact 8337 3600 8337 3600 4 n_191
rlabel m2contact 8361 4176 8361 4176 4 n_80
rlabel m2contact 8361 6864 8361 6864 4 n_3
rlabel m2contact 8385 3408 8385 3408 4 n_176
rlabel m2contact 8433 2568 8433 2568 4 n_262
rlabel m2contact 8457 5088 8457 5088 4 n_232
rlabel m2contact 8457 7056 8457 7056 4 n_287
rlabel m2contact 8481 5472 8481 5472 4 n_261
rlabel m2contact 8481 2544 8481 2544 4 n_293
rlabel m2contact 8505 7080 8505 7080 4 n_184
rlabel m2contact 8529 7104 8529 7104 4 n_263
rlabel m2contact 8529 2520 8529 2520 4 n_50
rlabel m2contact 8577 5376 8577 5376 4 n_219
rlabel m2contact 8577 2496 8577 2496 4 n_106
rlabel m2contact 8601 2496 8601 2496 4 n_106
rlabel m2contact 8601 5784 8601 5784 4 n_106
rlabel m2contact 8601 7128 8601 7128 4 n_88
rlabel m2contact 8625 2616 8625 2616 4 n_124
rlabel m2contact 8649 2808 8649 2808 4 n_10
rlabel m2contact 8673 4776 8673 4776 4 OpcodeCondIn[7]
rlabel m2contact 8673 3288 8673 3288 4 n_110
rlabel m2contact 8721 4296 8721 4296 4 n_81
rlabel m2contact 8721 7152 8721 7152 4 n_110
rlabel m2contact 8745 3288 8745 3288 4 n_110
rlabel m2contact 8745 7152 8745 7152 4 n_110
rlabel m2contact 8769 3576 8769 3576 4 n_35
rlabel m2contact 8793 6888 8793 6888 4 n_294
rlabel m2contact 8841 7152 8841 7152 4 n_295
rlabel m2contact 8913 3576 8913 3576 4 n_251
rlabel m2contact 8937 3528 8937 3528 4 n_186
rlabel m2contact 8937 2616 8937 2616 4 n_271
rlabel m2contact 8961 2496 8961 2496 4 n_259
rlabel m2contact 9009 7176 9009 7176 4 n_277
rlabel m2contact 9033 5808 9033 5808 4 n_276
rlabel m2contact 9057 2472 9057 2472 4 n_278
rlabel m2contact 9105 4536 9105 4536 4 n_95
rlabel m2contact 9129 4032 9129 4032 4 stateSub[0]
rlabel m2contact 9153 7200 9153 7200 4 n_96
rlabel m2contact 9201 7224 9201 7224 4 n_345
rlabel m2contact 9225 4440 9225 4440 4 n_373
rlabel m2contact 9249 6912 9249 6912 4 n_370
rlabel m2contact 9273 7248 9273 7248 4 n_355
rlabel m2contact 9345 4776 9345 4776 4 OpcodeCondIn[7]
rlabel m2contact 9345 2448 9345 2448 4 IntReq
rlabel m2contact 9369 7080 9369 7080 4 n_184
rlabel m2contact 9393 5856 9393 5856 4 n_217
rlabel m2contact 9417 6912 9417 6912 4 OpcodeCondIn[4]
rlabel m2contact 9441 7272 9441 7272 4 n_147
rlabel m2contact 9489 5088 9489 5088 4 n_232
rlabel m2contact 9489 2568 9489 2568 4 n_262
rlabel m2contact 9513 3672 9513 3672 4 n_218
rlabel m2contact 9513 2424 9513 2424 4 n_217
rlabel m2contact 9537 3936 9537 3936 4 n_49
rlabel m2contact 9537 3984 9537 3984 4 n_62
rlabel m2contact 9561 2424 9561 2424 4 n_217
rlabel m2contact 9561 5856 9561 5856 4 n_217
rlabel m2contact 9585 2832 9585 2832 4 stateSub[1]
rlabel m2contact 9585 2400 9585 2400 4 n_138
rlabel m2contact 9609 3168 9609 3168 4 n_193
rlabel m2contact 9609 3984 9609 3984 4 n_144
rlabel m2contact 9633 2424 9633 2424 4 n_146
rlabel m2contact 9657 6120 9657 6120 4 n_139
rlabel m2contact 9681 2640 9681 2640 4 n_205
rlabel m2contact 9705 3552 9705 3552 4 n_222
rlabel m2contact 9705 2376 9705 2376 4 n_307
rlabel m2contact 9729 6120 9729 6120 4 n_367
rlabel m2contact 9753 7296 9753 7296 4 PcSel[0]
rlabel m2contact 9753 7320 9753 7320 4 n_241
rlabel m2contact 9801 7344 9801 7344 4 OpcodeCondIn[2]
rlabel m2contact 9801 2352 9801 2352 4 n_92
rlabel m2contact 9825 4368 9825 4368 4 OpcodeCondIn[0]
rlabel m2contact 9825 2328 9825 2328 4 stateSub[2]
rlabel m2contact 9849 7368 9849 7368 4 n_6
rlabel m2contact 9897 3600 9897 3600 4 n_191
rlabel m2contact 9897 7296 9897 7296 4 PcSel[0]
rlabel m2contact 9921 7392 9921 7392 4 n_152
rlabel m2contact 9945 7296 9945 7296 4 n_257
rlabel m2contact 9969 7416 9969 7416 4 n_245
rlabel m2contact 9993 5784 9993 5784 4 n_106
rlabel m2contact 9993 7440 9993 7440 4 n_256
rlabel m2contact 10017 2592 10017 2592 4 n_52
rlabel m2contact 10041 2304 10041 2304 4 n_236
rlabel m2contact 10041 2280 10041 2280 4 n_315
rlabel m2contact 10065 2256 10065 2256 4 n_114
rlabel m2contact 10089 2232 10089 2232 4 n_122
rlabel m2contact 10113 2616 10113 2616 4 n_271
rlabel m2contact 10137 2256 10137 2256 4 n_114
rlabel m2contact 10161 4416 10161 4416 4 n_140
rlabel m2contact 10185 7440 10185 7440 4 n_256
rlabel m2contact 10209 2616 10209 2616 4 n_23
rlabel m2contact 10209 2256 10209 2256 4 n_349
rlabel m2contact 10281 3888 10281 3888 4 n_282
rlabel m2contact 10281 3552 10281 3552 4 n_222
rlabel m2contact 10305 4560 10305 4560 4 n_118
rlabel m2contact 10305 4032 10305 4032 4 stateSub[0]
rlabel m2contact 10329 6216 10329 6216 4 n_196
rlabel m2contact 10329 7440 10329 7440 4 n_305
rlabel m2contact 10353 7344 10353 7344 4 OpcodeCondIn[2]
rlabel m2contact 10377 3456 10377 3456 4 n_28
rlabel m2contact 10425 4824 10425 4824 4 n_299
rlabel m2contact 10425 5952 10425 5952 4 n_71
rlabel m2contact 10449 2208 10449 2208 4 n_67
rlabel m2contact 10473 4824 10473 4824 4 n_296
rlabel m2contact 10497 2832 10497 2832 4 stateSub[1]
rlabel m2contact 10521 4032 10521 4032 4 stateSub[0]
rlabel m2contact 10545 5352 10545 5352 4 n_75
rlabel m2contact 10569 5856 10569 5856 4 n_217
rlabel m2contact 10593 7464 10593 7464 4 n_17
rlabel m2contact 10617 5496 10617 5496 4 OpcodeCondIn[3]
rlabel m2contact 10641 5808 10641 5808 4 n_276
rlabel m2contact 10641 6288 10641 6288 4 n_51
rlabel m2contact 10665 4704 10665 4704 4 state[0]
rlabel m2contact 10689 3744 10689 3744 4 state[1]
rlabel m2contact 10713 4704 10713 4704 4 state[0]
rlabel m2contact 10713 2184 10713 2184 4 n_73
rlabel m2contact 10737 2184 10737 2184 4 n_73
rlabel m2contact 10737 5448 10737 5448 4 n_73
rlabel m2contact 10785 6984 10785 6984 4 n_126
rlabel m2contact 10809 2256 10809 2256 4 n_349
rlabel m2contact 10809 2184 10809 2184 4 n_207
rlabel m2contact 10857 3624 10857 3624 4 n_240
rlabel m2contact 10881 4416 10881 4416 4 n_140
rlabel m2contact 10881 7056 10881 7056 4 n_287
rlabel m2contact 10905 5448 10905 5448 4 n_297
rlabel m2contact 10929 2568 10929 2568 4 n_262
rlabel m2contact 10929 2160 10929 2160 4 n_104
rlabel m2contact 10953 6288 10953 6288 4 n_313
rlabel m2contact 10977 7152 10977 7152 4 n_295
rlabel m2contact 11001 7488 11001 7488 4 n_169
rlabel m2contact 11001 2136 11001 2136 4 n_267
rlabel m2contact 11025 5064 11025 5064 4 n_382
rlabel m2contact 11025 7152 11025 7152 4 IntReq
rlabel m2contact 11049 5088 11049 5088 4 n_232
rlabel m2contact 11049 2112 11049 2112 4 n_355
rlabel m2contact 11073 2448 11073 2448 4 IntReq
rlabel m2contact 11073 7152 11073 7152 4 IntReq
rlabel m2contact 11073 7512 11073 7512 4 n_233
rlabel m2contact 11073 2088 11073 2088 4 RwSel[1]
rlabel m2contact 11097 2112 11097 2112 4 n_355
rlabel m2contact 11097 7248 11097 7248 4 n_355
rlabel m2contact 11121 2160 11121 2160 4 n_104
rlabel m2contact 11121 7152 11121 7152 4 n_166
rlabel m2contact 11145 3168 11145 3168 4 n_193
rlabel m2contact 11169 2112 11169 2112 4 n_194
rlabel m2contact 11169 2064 11169 2064 4 n_105
rlabel m2contact 11217 7536 11217 7536 4 nWait
rlabel m2contact 11265 3816 11265 3816 4 n_237
rlabel m2contact 11289 7536 11289 7536 4 nWait
rlabel m2contact 11313 7464 11313 7464 4 n_17
rlabel m2contact 11337 5568 11337 5568 4 n_311
rlabel m2contact 11361 2736 11361 2736 4 n_170
rlabel m2contact 11385 7464 11385 7464 4 LrWe
rlabel m2contact 11409 7560 11409 7560 4 n_84
rlabel m2contact 11433 2040 11433 2040 4 n_42
rlabel m2contact 11481 5808 11481 5808 4 n_276
rlabel m2contact 11481 7584 11481 7584 4 n_52
rlabel m2contact 11505 2328 11505 2328 4 stateSub[2]
rlabel m2contact 11529 3696 11529 3696 4 n_365
rlabel m2contact 11553 2592 11553 2592 4 n_52
rlabel m2contact 11553 7584 11553 7584 4 n_52
rlabel m2contact 11553 2016 11553 2016 4 n_286
rlabel m2contact 11577 3816 11577 3816 4 n_237
rlabel m2contact 11577 7608 11577 7608 4 n_218
rlabel m2contact 11601 4056 11601 4056 4 n_19
rlabel m2contact 11601 1992 11601 1992 4 n_326
rlabel m2contact 11625 3672 11625 3672 4 n_218
rlabel m2contact 11625 7608 11625 7608 4 n_218
rlabel m2contact 11649 5184 11649 5184 4 n_20
rlabel m2contact 11649 2832 11649 2832 4 stateSub[1]
rlabel m2contact 11697 5616 11697 5616 4 OpcodeCondIn[6]
rlabel m2contact 11697 7584 11697 7584 4 n_348
rlabel m2contact 11721 5184 11721 5184 4 Op1Sel
rlabel m2contact 11769 4632 11769 4632 4 n_359
rlabel m2contact 11769 7608 11769 7608 4 n_372
rlabel m2contact 11793 3240 11793 3240 4 StatusReg[0]
rlabel m2contact 11817 7632 11817 7632 4 n_79
rlabel m2contact 11841 6432 11841 6432 4 n_86
rlabel m2contact 11865 4632 11865 4632 4 n_359
rlabel m2contact 11865 7656 11865 7656 4 stateSub[2]
rlabel m2contact 11889 5856 11889 5856 4 n_217
rlabel m2contact 11889 1968 11889 1968 4 StatusReg[3]
rlabel m2contact 11913 4104 11913 4104 4 n_357
rlabel m2contact 11913 4680 11913 4680 4 n_87
rlabel m2contact 11937 2328 11937 2328 4 stateSub[2]
rlabel m2contact 11937 7656 11937 7656 4 stateSub[2]
rlabel m2contact 11961 3096 11961 3096 4 n_100
rlabel m2contact 11961 1944 11961 1944 4 n_197
rlabel m2contact 11985 4224 11985 4224 4 n_153
rlabel m2contact 11985 2112 11985 2112 4 n_194
rlabel m2contact 12009 2472 12009 2472 4 n_278
rlabel m2contact 12009 7656 12009 7656 4 n_101
rlabel m2contact 12033 4680 12033 4680 4 n_107
rlabel m2contact 12057 2184 12057 2184 4 n_207
rlabel m2contact 12057 2112 12057 2112 4 n_330
rlabel m2contact 12081 6936 12081 6936 4 n_174
rlabel m2contact 12105 3696 12105 3696 4 n_365
rlabel m2contact 12105 4104 12105 4104 4 n_208
rlabel m2contact 12129 2472 12129 2472 4 n_162
rlabel m2contact 12153 3696 12153 3696 4 n_55
rlabel m2contact 12177 3816 12177 3816 4 n_237
rlabel m2contact 12177 2256 12177 2256 4 n_349
rlabel m2contact 12201 1944 12201 1944 4 n_197
rlabel m2contact 12201 6264 12201 6264 4 n_197
rlabel m2contact 12201 1920 12201 1920 4 Rs1Sel[0]
rlabel m2contact 12225 7056 12225 7056 4 n_287
rlabel m2contact 12249 3600 12249 3600 4 n_191
rlabel m2contact 12273 2736 12273 2736 4 n_170
rlabel m2contact 12273 7656 12273 7656 4 n_101
rlabel m2contact 12297 6264 12297 6264 4 n_175
rlabel m2contact 12297 1944 12297 1944 4 n_171
rlabel m2contact 12321 5256 12321 5256 4 n_239
rlabel m2contact 12345 3384 12345 3384 4 n_280
rlabel m2contact 12369 2328 12369 2328 4 stateSub[2]
rlabel m2contact 12369 5256 12369 5256 4 Rs1Sel[0]
rlabel m2contact 12393 1920 12393 1920 4 Rs1Sel[0]
rlabel m2contact 12393 5256 12393 5256 4 Rs1Sel[0]
rlabel m2contact 12417 3480 12417 3480 4 n_27
rlabel m2contact 12417 1896 12417 1896 4 n_111
rlabel m2contact 12441 4296 12441 4296 4 n_81
rlabel m2contact 12465 4368 12465 4368 4 OpcodeCondIn[0]
rlabel m2contact 12489 3936 12489 3936 4 n_49
rlabel m2contact 12489 6840 12489 6840 4 n_78
rlabel m2contact 12537 4392 12537 4392 4 n_157
rlabel m2contact 12561 5256 12561 5256 4 n_108
rlabel m2contact 12585 3288 12585 3288 4 n_110
rlabel m2contact 12585 6840 12585 6840 4 n_160
rlabel m2contact 12609 1920 12609 1920 4 n_289
rlabel m2contact 12633 4704 12633 4704 4 state[0]
rlabel m2contact 12657 3936 12657 3936 4 n_49
rlabel m2contact 12681 3384 12681 3384 4 n_280
rlabel m2contact 12681 2832 12681 2832 4 stateSub[1]
rlabel m2contact 12729 7656 12729 7656 4 n_180
rlabel m2contact 12753 3528 12753 3528 4 n_186
rlabel m2contact 12753 1872 12753 1872 4 n_56
rlabel m2contact 12777 2592 12777 2592 4 n_52
rlabel m2contact 12777 7680 12777 7680 4 n_161
rlabel m2contact 12801 1872 12801 1872 4 n_56
rlabel m2contact 12801 3792 12801 3792 4 n_56
rlabel m2contact 12825 3288 12825 3288 4 n_110
rlabel m2contact 12825 2640 12825 2640 4 n_205
rlabel m2contact 12849 6912 12849 6912 4 OpcodeCondIn[4]
rlabel m2contact 12873 7632 12873 7632 4 n_79
rlabel m2contact 12873 1872 12873 1872 4 n_69
rlabel m2contact 12921 6672 12921 6672 4 n_135
rlabel m2contact 12921 7704 12921 7704 4 n_274
rlabel m2contact 12945 7728 12945 7728 4 n_189
rlabel m2contact 12969 2136 12969 2136 4 n_267
rlabel m2contact 12993 1848 12993 1848 4 n_46
rlabel m2contact 13017 6744 13017 6744 4 n_47
rlabel m2contact 13017 7752 13017 7752 4 n_56
rlabel m2contact 13041 4968 13041 4968 4 n_98
rlabel m2contact 13041 7776 13041 7776 4 n_157
rlabel m2contact 13065 2136 13065 2136 4 n_99
rlabel m2contact 13089 5592 13089 5592 4 n_230
rlabel m2contact 13113 3288 13113 3288 4 n_110
rlabel m2contact 13137 5856 13137 5856 4 n_217
rlabel m2contact 13137 7800 13137 7800 4 n_170
rlabel m2contact 13161 3528 13161 3528 4 n_186
rlabel m2contact 13161 1824 13161 1824 4 n_22
rlabel m2contact 13185 5256 13185 5256 4 n_108
rlabel m2contact 13209 3792 13209 3792 4 n_56
rlabel m2contact 13209 7752 13209 7752 4 n_56
rlabel m2contact 13233 3792 13233 3792 4 n_56
rlabel m2contact 13257 2040 13257 2040 4 n_42
rlabel m2contact 13281 4392 13281 4392 4 n_157
rlabel m2contact 13281 7776 13281 7776 4 n_157
rlabel m2contact 13305 3096 13305 3096 4 n_100
rlabel m2contact 13329 5448 13329 5448 4 n_297
rlabel m2contact 13353 2736 13353 2736 4 n_170
rlabel m2contact 13353 7800 13353 7800 4 n_170
rlabel m2contact 13425 4248 13425 4248 4 n_43
rlabel m2contact 13449 2040 13449 2040 4 n_42
rlabel m2contact 13473 3528 13473 3528 4 n_186
rlabel m2contact 13497 6912 13497 6912 4 OpcodeCondIn[4]
rlabel m2contact 13521 3360 13521 3360 4 n_70
rlabel m2contact 13521 6432 13521 6432 4 n_86
rlabel m2contact 13569 7344 13569 7344 4 OpcodeCondIn[2]
rlabel m2contact 13593 3096 13593 3096 4 n_179
rlabel m2contact 13617 3816 13617 3816 4 n_237
rlabel m2contact 13641 6936 13641 6936 4 n_174
rlabel m2contact 13665 3552 13665 3552 4 n_222
rlabel m2contact 13689 2664 13689 2664 4 n_231
rlabel m2contact 13689 1800 13689 1800 4 n_175
rlabel m2contact 13713 4104 13713 4104 4 n_208
rlabel m2contact 13737 4824 13737 4824 4 n_296
rlabel m2contact 13737 2664 13737 2664 4 n_141
rlabel m2contact 13761 6960 13761 6960 4 n_102
rlabel m2contact 13761 7752 13761 7752 4 n_315
rlabel m2contact 13785 7584 13785 7584 4 n_348
rlabel m2contact 13797 1800 13797 1800 4 n_175
rlabel m2contact 13797 6264 13797 6264 4 n_175
rlabel m2contact 13833 6912 13833 6912 4 OpcodeCondIn[4]
rlabel m2contact 13833 7272 13833 7272 4 n_147
rlabel m2contact 13857 7560 13857 7560 4 n_84
rlabel m2contact 13881 2568 13881 2568 4 n_262
rlabel m2contact 13905 3144 13905 3144 4 n_202
rlabel m2contact 13929 2280 13929 2280 4 n_315
rlabel m2contact 13929 7752 13929 7752 4 n_315
rlabel m2contact 13953 3648 13953 3648 4 n_12
rlabel m2contact 13953 6360 13953 6360 4 n_284
rlabel m2contact 13977 4776 13977 4776 4 OpcodeCondIn[7]
rlabel m2contact 13977 4824 13977 4824 4 n_325
rlabel m2contact 14001 5424 14001 5424 4 n_7
rlabel m2contact 14025 5232 14025 5232 4 n_341
rlabel m2contact 14073 6984 14073 6984 4 n_126
rlabel m2contact 14121 6168 14121 6168 4 n_128
rlabel m2contact 14121 5352 14121 5352 4 n_75
rlabel m2contact 14193 3096 14193 3096 4 n_179
rlabel m2contact 14217 4224 14217 4224 4 n_153
rlabel m2contact 14241 6336 14241 6336 6 n_203
rlabel m2contact 14241 4104 14241 4104 6 n_58
rlabel m2contact 14265 4104 14265 4104 6 n_58
rlabel m2contact 14265 6456 14265 6456 6 n_58
rlabel m2contact 14289 5376 14289 5376 6 n_219
rlabel m2contact 14289 3144 14289 3144 6 n_161
rlabel m2contact 14313 2808 14313 2808 6 n_10
rlabel m2contact 14313 1800 14313 1800 6 n_147
rlabel m2contact 14337 7416 14337 7416 6 n_245
rlabel m2contact 14361 7296 14361 7296 6 n_257
rlabel m2contact 14385 4704 14385 4704 6 state[0]
rlabel m2contact 14409 3936 14409 3936 6 n_49
rlabel m2contact 14409 3672 14409 3672 6 n_218
rlabel m2contact 14433 4776 14433 4776 6 OpcodeCondIn[7]
rlabel m2contact 14433 3792 14433 3792 6 n_56
rlabel m2contact 14457 3144 14457 3144 6 n_161
rlabel m2contact 14457 7680 14457 7680 6 n_161
rlabel m2contact 14481 2736 14481 2736 6 n_170
rlabel m2contact 14481 1776 14481 1776 6 n_251
rlabel m2contact 14505 2832 14505 2832 6 stateSub[1]
rlabel m2contact 14529 2328 14529 2328 6 stateSub[2]
rlabel m2contact 14529 1752 14529 1752 6 n_252
rlabel m2contact 14553 4704 14553 4704 6 state[0]
rlabel m2contact 14577 4776 14577 4776 6 n_65
rlabel m2contact 14601 4248 14601 4248 6 n_43
rlabel m2contact 14601 3672 14601 3672 6 n_218
rlabel m2contact 14625 1800 14625 1800 6 n_147
rlabel m2contact 14625 7272 14625 7272 6 n_147
rlabel m2contact 14649 2184 14649 2184 6 n_207
rlabel m2contact 14673 3672 14673 3672 6 n_218
rlabel m2contact 14673 3144 14673 3144 6 n_381
rlabel m2contact 14697 4968 14697 4968 6 n_243
rlabel m2contact 14721 7032 14721 7032 6 n_324
rlabel m2contact 14745 2544 14745 2544 6 n_293
rlabel m2contact 14745 2184 14745 2184 6 n_389
rlabel m2contact 14769 7104 14769 7104 6 n_263
rlabel m2contact 14793 5256 14793 5256 6 n_364
rlabel m2contact 14793 4104 14793 4104 6 n_165
rlabel m2contact 14817 4128 14817 4128 6 n_384
rlabel m2contact 14829 1776 14829 1776 6 n_251
rlabel m2contact 14829 3576 14829 3576 6 n_251
rlabel m2contact 14865 4128 14865 4128 6 n_173
rlabel m2contact 14889 4200 14889 4200 6 nWE
rlabel m2contact 14889 4344 14889 4344 6 OpcodeCondIn[1]
rlabel m2contact 14937 4752 14937 4752 6 n_11
rlabel m2contact 14961 6312 14961 6312 6 n_159
rlabel m2contact 14985 4080 14985 4080 6 n_255
rlabel m2contact 15009 3336 15009 3336 6 n_306
rlabel m2contact 15033 2784 15033 2784 6 n_268
rlabel m2contact 15033 3096 15033 3096 6 n_179
rlabel m2contact 15057 5568 15057 5568 6 n_311
rlabel m2contact 15057 4200 15057 4200 6 n_287
rlabel m2contact 15081 4200 15081 4200 6 n_287
rlabel m2contact 15081 7056 15081 7056 6 n_287
rlabel m2contact 15105 5184 15105 5184 6 Op1Sel
rlabel m2contact 15105 5424 15105 5424 6 n_229
rlabel m2contact 15129 3336 15129 3336 6 n_306
rlabel m2contact 15153 2376 15153 2376 6 n_307
rlabel m2contact 15153 1800 15153 1800 6 n_154
rlabel m2contact 15201 5184 15201 5184 6 n_178
rlabel m2contact 15225 7704 15225 7704 6 n_274
rlabel m2contact 15249 5616 15249 5616 6 OpcodeCondIn[6]
rlabel m2contact 15273 5568 15273 5568 6 n_279
rlabel m2contact 15321 1968 15321 1968 6 StatusReg[3]
rlabel m2contact 15345 5928 15345 5928 6 n_347
rlabel m2contact 15345 6168 15345 6168 6 n_506
rlabel m2contact 15369 1848 15369 1848 6 n_46
rlabel m2contact 15393 2952 15393 2952 6 n_506
rlabel m2contact 15393 6168 15393 6168 6 n_506
rlabel m2contact 15489 4512 15489 4512 6 n_391
rlabel m2contact 15753 4512 15753 4512 6 InISR
rlabel m2contact 15849 6696 15849 6696 6 n_507
rlabel m2contact 15897 1968 15897 1968 6 StatusReg[3]
rlabel m2contact 15897 1776 15897 1776 6 n_36
rlabel m2contact 15921 4200 15921 4200 6 n_29
rlabel m2contact 15993 7248 15993 7248 6 n_355
rlabel m2contact 16041 2016 16041 2016 6 n_286
rlabel m2contact 16041 5928 16041 5928 6 PcSel[1]
rlabel m2contact 16113 4800 16113 4800 6 n_379
rlabel m2contact 16161 6096 16161 6096 6 n_366
rlabel m2contact 16161 3000 16161 3000 6 n_378
rlabel m2contact 16209 6456 16209 6456 6 n_58
rlabel m2contact 16257 6648 16257 6648 6 n_59
rlabel m2contact 16329 5496 16329 5496 6 OpcodeCondIn[3]
rlabel m2contact 16377 2688 16377 2688 6 n_224
rlabel m2contact 16449 5808 16449 5808 6 n_276
rlabel m2contact 16521 5376 16521 5376 6 n_219
rlabel m2contact 16521 4080 16521 4080 6 n_47
rlabel m2contact 16545 1848 16545 1848 6 n_46
rlabel m2contact 16569 2328 16569 2328 6 stateSub[2]
rlabel m2contact 16593 4080 16593 4080 6 n_47
rlabel m2contact 16593 6744 16593 6744 6 n_47
rlabel m2contact 16665 4080 16665 4080 6 n_333
rlabel m2contact 16713 4200 16713 4200 6 n_29
rlabel m2contact 16737 4296 16737 4296 6 n_81
rlabel m2contact 16761 3912 16761 3912 6 n_112
rlabel m2contact 16761 6528 16761 6528 6 n_30
rlabel m2contact 16785 1872 16785 1872 6 n_69
rlabel m2contact 16833 3960 16833 3960 6 n_13
rlabel m2contact 16833 4944 16833 4944 6 n_53
rlabel m2contact 16857 3216 16857 3216 6 n_54
rlabel m2contact 16881 7368 16881 7368 6 n_6
rlabel m2contact 16905 3984 16905 3984 6 n_144
rlabel m2contact 16953 5376 16953 5376 6 n_219
rlabel m2contact 16953 7296 16953 7296 6 n_257
rlabel m2contact 16977 3672 16977 3672 6 n_218
rlabel m2contact 16977 5808 16977 5808 6 n_290
rlabel m2contact 17001 6000 17001 6000 6 n_328
rlabel m2contact 17025 5016 17025 5016 6 n_172
rlabel m2contact 17049 6000 17049 6000 6 n_265
rlabel m2contact 17073 4440 17073 4440 6 n_373
rlabel m2contact 17073 6096 17073 6096 6 n_266
rlabel m2contact 17097 5280 17097 5280 6 n_316
rlabel m2contact 17097 3336 17097 3336 6 n_313
rlabel m2contact 17121 2280 17121 2280 6 n_315
rlabel m2contact 17121 1968 17121 1968 6 n_331
rlabel m2contact 17145 6120 17145 6120 6 n_367
rlabel m2contact 17169 4440 17169 4440 6 PcWe
rlabel m2contact 17193 5472 17193 5472 6 n_261
rlabel m2contact 17217 6480 17217 6480 6 n_132
rlabel m2contact 17217 3000 17217 3000 6 n_123
rlabel m2contact 17241 6432 17241 6432 6 n_86
rlabel m2contact 17241 6528 17241 6528 6 n_268
rlabel m2contact 17265 3336 17265 3336 6 n_313
rlabel m2contact 17265 6288 17265 6288 6 n_313
rlabel m2contact 17289 4440 17289 4440 6 PcWe
rlabel m2contact 17289 2952 17289 2952 6 n_209
rlabel m2contact 17313 2784 17313 2784 6 n_268
rlabel m2contact 17313 6528 17313 6528 6 n_268
rlabel m2contact 17337 3192 17337 3192 6 n_41
rlabel m2contact 17361 7344 17361 7344 6 OpcodeCondIn[2]
rlabel m2contact 17385 6168 17385 6168 6 n_90
rlabel m2contact 17433 6264 17433 6264 6 n_318
rlabel m2contact 17457 6288 17457 6288 6 n_212
rlabel m2contact 17481 2496 17481 2496 6 n_259
rlabel m2contact 17505 7200 17505 7200 6 n_96
rlabel m2contact 17577 6936 17577 6936 6 n_174
rlabel m2contact 17601 4776 17601 4776 6 n_65
rlabel m2contact 17649 2760 17649 2760 6 n_155
rlabel m2contact 17697 5232 17697 5232 6 n_341
rlabel m2contact 17721 7248 17721 7248 6 n_355
rlabel m2contact 17745 5232 17745 5232 6 AluOR[1]
rlabel m2contact 17793 5016 17793 5016 6 n_172
rlabel m2contact 17817 3552 17817 3552 6 n_222
rlabel m2contact 17841 4128 17841 4128 6 n_173
rlabel m2contact 17889 3288 17889 3288 6 n_110
rlabel m2contact 17913 4032 17913 4032 6 stateSub[0]
rlabel m2contact 17937 7080 17937 7080 6 n_184
rlabel m2contact 17961 7008 17961 7008 6 n_214
rlabel m2contact 17961 7032 17961 7032 6 n_45
rlabel m2contact 17985 5160 17985 5160 6 n_253
rlabel m2contact 18009 3888 18009 3888 6 n_282
rlabel m2contact 18009 6336 18009 6336 6 n_4
rlabel m2contact 18033 4704 18033 4704 6 state[0]
rlabel m2contact 18057 3432 18057 3432 6 n_25
rlabel m2contact 18081 7656 18081 7656 6 n_180
rlabel m2contact 18105 3120 18105 3120 6 n_198
rlabel m2contact 18105 2784 18105 2784 6 n_316
rlabel m2contact 18129 2784 18129 2784 6 n_316
rlabel m2contact 18129 5280 18129 5280 6 n_316
rlabel m2contact 18153 5352 18153 5352 6 n_75
rlabel m2contact 18153 7704 18153 7704 6 n_274
rlabel m2contact 18201 4560 18201 4560 6 n_118
rlabel m2contact 18273 7320 18273 7320 6 n_241
rlabel m2contact 18297 5496 18297 5496 6 OpcodeCondIn[3]
rlabel m2contact 18297 6360 18297 6360 6 n_388
rlabel m2contact 18321 6408 18321 6408 6 n_339
rlabel m2contact 18369 7224 18369 7224 6 n_345
rlabel m2contact 18489 7416 18489 7416 6 n_245
rlabel m2contact 18537 4560 18537 4560 6 n_246
rlabel m2contact 18657 3912 18657 3912 6 n_112
rlabel m2contact 18729 4440 18729 4440 6 n_226
rlabel m2contact 18777 4128 18777 4128 6 WdSel
rlabel m2contact 18849 2208 18849 2208 6 n_67
rlabel m2contact 18849 1848 18849 1848 6 n_250
rlabel m2contact 18873 3912 18873 3912 6 n_112
rlabel m2contact 18873 2880 18873 2880 6 n_386
rlabel m2contact 18897 6504 18897 6504 6 n_362
rlabel m2contact 18921 6408 18921 6408 6 n_339
rlabel m2contact 18921 6528 18921 6528 6 n_68
rlabel m2contact 18945 3888 18945 3888 6 ImmSel
rlabel m2contact 18969 4536 18969 4536 6 n_95
rlabel m2contact 18993 5088 18993 5088 6 n_232
rlabel m2contact 19017 5568 19017 5568 6 n_279
rlabel m2contact 19017 6408 19017 6408 6 n_94
rlabel m2contact 19065 5040 19065 5040 6 n_74
rlabel m2contact 19089 5328 19089 5328 6 n_344
rlabel m2contact 19113 2400 19113 2400 6 n_138
rlabel m2contact 19137 4584 19137 4584 6 n_227
rlabel m2contact 19161 3624 19161 3624 6 n_240
rlabel m2contact 19185 3888 19185 3888 6 ImmSel
rlabel m2contact 19209 6216 19209 6216 6 n_196
rlabel m2contact 19233 4128 19233 4128 6 WdSel
rlabel m2contact 19281 4320 19281 4320 6 n_18
rlabel m2contact 19281 7728 19281 7728 6 n_189
rlabel m2contact 19305 6216 19305 6216 6 n_196
rlabel m2contact 19329 7344 19329 7344 6 OpcodeCondIn[2]
rlabel m2contact 19353 6024 19353 6024 6 n_63
rlabel m2contact 19353 6768 19353 6768 6 n_188
rlabel m2contact 19377 3528 19377 3528 6 n_186
rlabel m2contact 19401 2112 19401 2112 6 n_330
rlabel m2contact 19401 1728 19401 1728 6 n_64
rlabel m2contact 19449 4272 19449 4272 6 n_343
rlabel m2contact 19449 2832 19449 2832 6 stateSub[1]
rlabel m2contact 19473 4056 19473 4056 6 n_19
rlabel m2contact 19497 2592 19497 2592 6 n_52
rlabel m2contact 19521 3264 19521 3264 6 n_26
rlabel m2contact 19545 7032 19545 7032 6 n_45
rlabel m2contact 19569 6456 19569 6456 6 n_58
rlabel m2contact 19593 5688 19593 5688 6 n_148
rlabel m2contact 19617 6864 19617 6864 6 n_3
rlabel m2contact 19641 7224 19641 7224 6 n_345
rlabel m2contact 19665 5880 19665 5880 6 n_300
rlabel m2contact 19689 5400 19689 5400 6 n_182
rlabel m2contact 19713 4800 19713 4800 6 n_379
rlabel m2contact 19761 4392 19761 4392 6 n_157
rlabel m2contact 19809 7728 19809 7728 6 n_189
rlabel m2contact 19881 7704 19881 7704 6 n_274
rlabel m2contact 19905 6240 19905 6240 6 n_195
rlabel m2contact 19929 5064 19929 5064 6 n_382
rlabel m2contact 19977 3744 19977 3744 6 state[1]
rlabel m2contact 20001 3168 20001 3168 6 n_193
rlabel m2contact 20025 5088 20025 5088 6 n_15
rlabel m2contact 20073 4848 20073 4848 6 n_322
rlabel m2contact 20097 5280 20097 5280 6 SysBus[2]
rlabel m2contact 20121 6384 20121 6384 6 n_321
rlabel m2contact 20169 3384 20169 3384 6 n_280
rlabel m2contact 20169 2592 20169 2592 6 n_52
rlabel m2contact 20193 4704 20193 4704 6 state[0]
rlabel m2contact 20193 5328 20193 5328 6 n_138
rlabel m2contact 20217 5208 20217 5208 6 n_273
rlabel m2contact 20241 2352 20241 2352 6 n_92
rlabel m2contact 20241 5088 20241 5088 6 n_15
rlabel m2contact 20265 2400 20265 2400 6 n_138
rlabel m2contact 20265 5328 20265 5328 6 n_138
rlabel m2contact 20289 7704 20289 7704 6 n_274
rlabel m2contact 20313 2736 20313 2736 6 n_170
rlabel m2contact 20313 5088 20313 5088 6 n_286
rlabel m2contact 20337 3024 20337 3024 6 n_264
rlabel m2contact 20337 7344 20337 7344 6 OpcodeCondIn[2]
rlabel m2contact 20361 2016 20361 2016 6 n_286
rlabel m2contact 20361 5088 20361 5088 6 n_286
rlabel m2contact 20385 4848 20385 4848 6 n_322
rlabel m2contact 20385 4296 20385 4296 6 n_81
rlabel m2contact 20433 6168 20433 6168 6 n_90
rlabel m2contact 20457 5088 20457 5088 6 n_24
rlabel m2contact 20481 4896 20481 4896 6 n_158
rlabel m2contact 20505 5952 20505 5952 6 n_71
rlabel m2contact 20505 6168 20505 6168 6 n_99
rlabel m2contact 20529 7704 20529 7704 6 n_274
rlabel m2contact 20529 7752 20529 7752 6 n_229
rlabel m2contact 20553 2136 20553 2136 6 n_99
rlabel m2contact 20553 6168 20553 6168 6 n_99
rlabel m2contact 20577 2952 20577 2952 6 n_209
rlabel m2contact 20577 2784 20577 2784 6 n_275
rlabel m2contact 20601 5856 20601 5856 6 n_217
rlabel m2contact 20625 6480 20625 6480 6 n_132
rlabel m2contact 20625 7224 20625 7224 6 n_345
rlabel m2contact 20649 6528 20649 6528 6 n_68
rlabel m2contact 20673 4368 20673 4368 6 OpcodeCondIn[0]
rlabel m2contact 20697 3240 20697 3240 6 StatusReg[0]
rlabel m2contact 20721 4344 20721 4344 6 OpcodeCondIn[1]
rlabel m2contact 20745 3984 20745 3984 6 n_144
rlabel m2contact 20745 5088 20745 5088 6 n_24
rlabel m2contact 20769 5424 20769 5424 6 n_229
rlabel m2contact 20769 7752 20769 7752 6 n_229
rlabel m2contact 20793 4416 20793 4416 6 n_140
rlabel m2contact 20817 2640 20817 2640 6 n_205
rlabel m2contact 20841 4224 20841 4224 6 n_153
rlabel m2contact 20841 5496 20841 5496 6 OpcodeCondIn[3]
rlabel m2contact 20865 7704 20865 7704 6 n_274
rlabel m2contact 20865 7752 20865 7752 6 n_141
rlabel m2contact 20889 4416 20889 4416 6 n_140
rlabel m2contact 20913 5640 20913 5640 6 n_82
rlabel m2contact 20913 4392 20913 4392 6 n_272
rlabel m2contact 20937 5712 20937 5712 6 n_168
rlabel m2contact 20961 2880 20961 2880 6 n_386
rlabel m2contact 20961 4080 20961 4080 6 n_333
rlabel m2contact 20985 6552 20985 6552 6 n_103
rlabel m2contact 20985 4416 20985 4416 6 n_372
rlabel m2contact 21009 5064 21009 5064 6 n_382
rlabel m2contact 21009 5088 21009 5088 6 n_375
rlabel m2contact 21033 4008 21033 4008 6 AluEn
rlabel m2contact 21057 6120 21057 6120 6 n_367
rlabel m2contact 21081 4224 21081 4224 6 n_153
rlabel m2contact 21093 4416 21093 4416 6 n_372
rlabel m2contact 21093 7608 21093 7608 6 n_372
rlabel m2contact 21129 7128 21129 7128 6 n_88
rlabel m2contact 21153 2664 21153 2664 6 n_141
rlabel m2contact 21153 7752 21153 7752 6 n_141
rlabel m2contact 21177 2520 21177 2520 6 n_50
rlabel m2contact 21201 2832 21201 2832 6 stateSub[1]
rlabel m2contact 21201 2664 21201 2664 6 n_115
rlabel m2contact 21225 4056 21225 4056 6 n_19
rlabel m2contact 21249 4824 21249 4824 6 n_325
rlabel m2contact 21273 6072 21273 6072 6 n_163
rlabel m2contact 21297 5160 21297 5160 6 n_253
rlabel m2contact 21321 3216 21321 3216 6 n_54
rlabel m2contact 21345 4536 21345 4536 6 n_95
rlabel m2contact 21345 4416 21345 4416 6 n_53
rlabel m2contact 21369 3696 21369 3696 6 n_55
rlabel m2contact 21381 4416 21381 4416 6 n_53
rlabel m2contact 21381 4944 21381 4944 6 n_53
rlabel m2contact 21417 4608 21417 4608 6 n_304
rlabel m2contact 21417 3000 21417 3000 6 n_123
rlabel m2contact 21441 3408 21441 3408 6 n_176
rlabel m2contact 21465 3600 21465 3600 6 n_191
rlabel m2contact 21489 1968 21489 1968 6 n_331
rlabel m2contact 21537 6216 21537 6216 6 n_196
rlabel m2contact 21537 6240 21537 6240 6 n_116
rlabel m2contact 21561 3552 21561 3552 6 n_222
rlabel m2contact 21561 4104 21561 4104 6 n_165
rlabel m2contact 21585 7152 21585 7152 6 n_166
rlabel m2contact 21585 6264 21585 6264 6 n_318
rlabel m2contact 21633 7296 21633 7296 6 n_257
rlabel m2contact 21633 7344 21633 7344 6 n_105
rlabel m2contact 21657 4224 21657 4224 6 n_153
rlabel m2contact 21681 1800 21681 1800 6 n_154
rlabel m2contact 21705 2064 21705 2064 6 n_105
rlabel m2contact 21705 7344 21705 7344 6 n_105
rlabel m2contact 21729 5784 21729 5784 6 n_106
rlabel m2contact 21729 1776 21729 1776 6 n_36
rlabel m2contact 21753 2832 21753 2832 6 stateSub[1]
rlabel m2contact 21777 2208 21777 2208 6 n_67
rlabel m2contact 21777 4680 21777 4680 6 n_107
rlabel m2contact 21825 4056 21825 4056 6 n_19
rlabel m2contact 21849 3168 21849 3168 6 n_193
rlabel m2contact 21849 2736 21849 2736 6 n_170
rlabel m2contact 21873 3912 21873 3912 6 n_112
rlabel m2contact 21873 4896 21873 4896 6 n_42
rlabel m2contact 21897 5760 21897 5760 6 n_130
rlabel m2contact 21921 2760 21921 2760 6 n_155
rlabel m2contact 21945 3936 21945 3936 6 n_49
rlabel m2contact 21945 6840 21945 6840 6 n_160
rlabel m2contact 21969 3504 21969 3504 6 n_215
rlabel m2contact 21969 3288 21969 3288 6 n_110
rlabel m2contact 21993 6576 21993 6576 6 n_40
rlabel m2contact 22017 5064 22017 5064 6 n_137
rlabel m2contact 22041 4848 22041 4848 6 n_322
rlabel m2contact 22041 5208 22041 5208 6 n_22
rlabel m2contact 22065 5184 22065 5184 6 n_178
rlabel m2contact 22065 4680 22065 4680 6 SysBus[3]
rlabel m2contact 22089 4488 22089 4488 6 n_320
rlabel m2contact 22113 2040 22113 2040 6 n_42
rlabel m2contact 22113 4896 22113 4896 6 n_42
rlabel m2contact 22137 1824 22137 1824 6 n_22
rlabel m2contact 22137 5208 22137 5208 6 n_22
rlabel m2contact 22185 2184 22185 2184 6 n_389
rlabel m2contact 22185 2136 22185 2136 6 ALE
rlabel m2contact 22281 2232 22281 2232 6 n_122
rlabel m2contact 22329 3648 22329 3648 6 n_12
rlabel m2contact 22353 2328 22353 2328 6 stateSub[2]
rlabel m2contact 22449 2424 22449 2424 6 n_146
rlabel m2contact 22473 7080 22473 7080 6 n_184
rlabel m2contact 22497 3048 22497 3048 6 n_185
rlabel m2contact 22545 7176 22545 7176 6 n_277
rlabel m2contact 22569 3168 22569 3168 6 n_193
rlabel m2contact 22593 3240 22593 3240 6 StatusReg[0]
rlabel m2contact 22641 4248 22641 4248 6 n_43
rlabel m2contact 22665 4032 22665 4032 6 stateSub[0]
rlabel m2contact 22689 4104 22689 4104 6 n_165
rlabel m2contact 22737 2568 22737 2568 6 n_262
rlabel m2contact 22737 7464 22737 7464 6 LrWe
rlabel m2contact 22785 1776 22785 1776 6 n_36
rlabel m2contact 22785 2136 22785 2136 6 ALE
rlabel m2contact 22833 5040 22833 5040 6 n_74
rlabel m2contact 22857 4848 22857 4848 6 n_5
rlabel m2contact 22905 2664 22905 2664 6 n_115
rlabel m2contact 22929 3216 22929 3216 6 n_54
rlabel m2contact 22953 3816 22953 3816 6 n_237
rlabel m2contact 22953 4896 22953 4896 6 n_186
rlabel m2contact 22977 3768 22977 3768 6 n_34
rlabel m2contact 22977 5856 22977 5856 6 n_217
rlabel m2contact 23001 4200 23001 4200 6 n_29
rlabel m2contact 23025 4632 23025 4632 6 n_359
rlabel m2contact 23049 5520 23049 5520 6 n_269
rlabel m2contact 23049 2928 23049 2928 6 StatusReg[2]
rlabel m2contact 23073 2976 23073 2976 6 n_358
rlabel m2contact 23097 5448 23097 5448 6 n_297
rlabel m2contact 23121 3744 23121 3744 6 state[1]
rlabel m2contact 23145 7536 23145 7536 6 nWait
rlabel m2contact 23169 5496 23169 5496 6 OpcodeCondIn[3]
rlabel m2contact 23193 4848 23193 4848 6 n_5
rlabel m2contact 23217 4896 23217 4896 6 n_186
rlabel m2contact 23241 6672 23241 6672 6 n_135
rlabel m2contact 23265 5856 23265 5856 6 n_217
rlabel m2contact 23289 6720 23289 6720 6 n_301
rlabel m2contact 23313 1920 23313 1920 6 n_289
rlabel m2contact 23337 4032 23337 4032 6 stateSub[0]
rlabel m2contact 23337 4848 23337 4848 6 n_275
rlabel m2contact 23361 3624 23361 3624 6 n_240
rlabel m2contact 23385 5592 23385 5592 6 n_230
rlabel m2contact 23409 3816 23409 3816 6 n_237
rlabel m2contact 23409 7704 23409 7704 6 n_274
rlabel m2contact 23433 3552 23433 3552 6 n_222
rlabel m2contact 23457 6096 23457 6096 6 n_266
rlabel m2contact 23481 7656 23481 7656 6 n_180
rlabel m2contact 23505 6216 23505 6216 6 n_196
rlabel m2contact 23505 6384 23505 6384 6 n_104
rlabel m2contact 23529 7656 23529 7656 6 n_180
rlabel m2contact 23529 3096 23529 3096 6 n_179
rlabel m2contact 23541 3528 23541 3528 6 n_186
rlabel m2contact 23541 4896 23541 4896 6 n_186
rlabel m2contact 23577 3840 23577 3840 6 n_213
rlabel m2contact 23601 4824 23601 4824 6 n_325
rlabel m2contact 23625 4032 23625 4032 6 stateSub[0]
rlabel m2contact 23625 5616 23625 5616 6 OpcodeCondIn[6]
rlabel m2contact 23649 5496 23649 5496 6 OpcodeCondIn[3]
rlabel m2contact 23661 2784 23661 2784 6 n_275
rlabel m2contact 23661 4848 23661 4848 6 n_275
rlabel m2contact 23697 7080 23697 7080 6 n_184
rlabel m2contact 23697 2448 23697 2448 6 IntReq
rlabel m2contact 23721 6120 23721 6120 6 n_367
rlabel m2contact 23745 4728 23745 4728 6 n_149
rlabel m2contact 23745 2304 23745 2304 6 n_236
rlabel m2contact 23769 1872 23769 1872 6 n_69
rlabel m2contact 23793 3600 23793 3600 6 n_191
rlabel m2contact 23793 7488 23793 7488 6 n_169
rlabel m2contact 23817 2160 23817 2160 6 n_104
rlabel m2contact 23817 6384 23817 6384 6 n_104
rlabel m2contact 23841 3792 23841 3792 6 n_56
rlabel m2contact 23865 5472 23865 5472 6 n_261
rlabel m2contact 23865 5520 23865 5520 6 n_193
rlabel m2contact 23889 3168 23889 3168 6 n_193
rlabel m2contact 23889 5520 23889 5520 6 n_193
rlabel m2contact 23913 4584 23913 4584 6 n_227
rlabel m2contact 23913 4536 23913 4536 6 n_189
rlabel m2contact 23937 5376 23937 5376 6 n_219
rlabel m2contact 23961 4584 23961 4584 6 n_227
rlabel m2contact 23961 6624 23961 6624 6 n_380
rlabel m2contact 23985 4656 23985 4656 6 n_360
rlabel m2contact 23985 2688 23985 2688 6 n_224
rlabel m2contact 24009 4872 24009 4872 6 n_323
rlabel m2contact 24009 4728 24009 4728 6 n_190
rlabel m2contact 24033 6360 24033 6360 6 n_388
rlabel m2contact 24057 2904 24057 2904 6 n_340
rlabel m2contact 24081 2832 24081 2832 6 stateSub[1]
rlabel m2contact 24081 2784 24081 2784 6 n_325
rlabel m2contact 24105 5496 24105 5496 6 OpcodeCondIn[3]
rlabel m2contact 24129 3720 24129 3720 6 n_363
rlabel m2contact 24129 6336 24129 6336 6 n_4
rlabel m2contact 24153 4536 24153 4536 6 n_189
rlabel m2contact 24153 7728 24153 7728 6 n_189
rlabel m2contact 24177 2640 24177 2640 6 n_205
rlabel m2contact 24177 2592 24177 2592 6 n_243
rlabel m2contact 24201 2328 24201 2328 6 stateSub[2]
rlabel m2contact 24225 7176 24225 7176 6 n_277
rlabel m2contact 24225 7200 24225 7200 6 n_123
rlabel m2contact 24249 2784 24249 2784 6 n_325
rlabel m2contact 24249 4824 24249 4824 6 n_325
rlabel m2contact 24273 3672 24273 3672 6 n_218
rlabel m2contact 24297 4752 24297 4752 6 n_11
rlabel m2contact 24297 4824 24297 4824 6 n_246
rlabel m2contact 24321 5808 24321 5808 6 n_290
rlabel m2contact 24345 4944 24345 4944 6 n_53
rlabel m2contact 24369 5376 24369 5376 6 n_219
rlabel m2contact 24393 5496 24393 5496 6 OpcodeCondIn[3]
rlabel m2contact 24393 2952 24393 2952 6 n_209
rlabel m2contact 24417 6024 24417 6024 6 n_63
rlabel m2contact 24441 3624 24441 3624 6 n_240
rlabel m2contact 24441 3600 24441 3600 6 n_210
rlabel m2contact 24465 2592 24465 2592 6 n_243
rlabel m2contact 24465 4968 24465 4968 6 n_243
rlabel m2contact 24489 4512 24489 4512 6 InISR
rlabel m2contact 24513 1992 24513 1992 6 n_326
rlabel m2contact 24537 5904 24537 5904 6 n_327
rlabel m2contact 24549 4560 24549 4560 6 n_246
rlabel m2contact 24549 4824 24549 4824 6 n_246
rlabel m2contact 24585 4248 24585 4248 6 n_43
rlabel m2contact 24609 4224 24609 4224 6 n_153
rlabel m2contact 24609 4824 24609 4824 6 state[1]
rlabel m2contact 24633 2520 24633 2520 6 n_50
rlabel m2contact 24657 3000 24657 3000 6 n_123
rlabel m2contact 24657 7200 24657 7200 6 n_123
rlabel m2contact 24681 7656 24681 7656 6 n_180
rlabel m2contact 24681 7680 24681 7680 6 n_272
rlabel m2contact 24705 1944 24705 1944 6 n_171
rlabel m2contact 24729 4800 24729 4800 6 n_379
rlabel m2contact 24753 2880 24753 2880 6 n_386
rlabel m2contact 24777 5256 24777 5256 6 n_364
rlabel m2contact 24801 6144 24801 6144 6 n_221
rlabel m2contact 24813 3744 24813 3744 6 state[1]
rlabel m2contact 24813 4824 24813 4824 6 state[1]
rlabel m2contact 24849 4464 24849 4464 6 n_247
rlabel m2contact 24849 3840 24849 3840 6 n_213
rlabel m2contact 24873 2640 24873 2640 6 n_205
rlabel m2contact 24897 7248 24897 7248 6 n_355
rlabel m2contact 24921 3840 24921 3840 6 n_213
rlabel m2contact 24945 4584 24945 4584 6 n_227
rlabel m2contact 24969 6288 24969 6288 6 n_212
rlabel m2contact 24969 4752 24969 4752 6 n_94
rlabel m2contact 24993 4392 24993 4392 6 n_272
rlabel m2contact 24993 7680 24993 7680 6 n_272
rlabel m2contact 25017 5544 25017 5544 6 n_121
rlabel m2contact 25041 3744 25041 3744 6 state[1]
rlabel m2contact 25065 6120 25065 6120 6 n_367
rlabel m2contact 25089 4752 25089 4752 6 n_94
rlabel m2contact 25089 6408 25089 6408 6 n_94
rlabel m2contact 25113 3480 25113 3480 6 n_27
rlabel m2contact 25161 3360 25161 3360 6 n_70
rlabel m2contact 25233 2352 25233 2352 6 n_92
rlabel m2contact 25257 3672 25257 3672 6 n_218
rlabel m2contact 25281 6048 25281 6048 6 n_109
rlabel m2contact 25329 1752 25329 1752 6 n_252
rlabel m2contact 25353 7440 25353 7440 6 n_305
rlabel m2contact 25377 6264 25377 6264 6 n_318
rlabel m2contact 25401 4152 25401 4152 6 ENB
rlabel m2contact 25449 4584 25449 4584 6 n_227
rlabel m2contact 25473 3072 25473 3072 6 n_225
rlabel m2contact 25497 2808 25497 2808 6 n_10
rlabel m2contact 25497 4824 25497 4824 6 n_224
rlabel m2contact 25521 4440 25521 4440 6 n_226
rlabel m2contact 25545 4704 25545 4704 6 state[0]
rlabel m2contact 25569 5160 25569 5160 6 n_253
rlabel m2contact 25593 2832 25593 2832 6 stateSub[1]
rlabel m2contact 25617 2688 25617 2688 6 n_224
rlabel m2contact 25617 4824 25617 4824 6 n_224
rlabel m2contact 25641 5112 25641 5112 6 n_83
rlabel m2contact 25689 6432 25689 6432 6 n_86
rlabel m2contact 25689 4968 25689 4968 6 n_243
rlabel m2contact 25713 5160 25713 5160 6 n_253
rlabel m2contact 25713 6648 25713 6648 6 n_59
rlabel m2contact 25737 6600 25737 6600 6 n_60
rlabel m2contact 25785 5736 25785 5736 6 n_308
rlabel m2contact 25785 2352 25785 2352 6 n_92
rlabel m2contact 25809 3744 25809 3744 6 state[1]
rlabel m2contact 25809 4824 25809 4824 6 n_349
rlabel m2contact 25833 2256 25833 2256 6 n_349
rlabel m2contact 25833 4824 25833 4824 6 n_349
rlabel m2contact 25857 5136 25857 5136 6 n_91
rlabel m2contact 25881 4824 25881 4824 6 n_242
rlabel m2contact 25905 5832 25905 5832 6 n_346
rlabel m2contact 25929 6888 25929 6888 6 n_294
rlabel m2contact 25977 1896 25977 1896 6 n_111
rlabel m2contact 26001 2856 26001 2856 6 n_76
rlabel m2contact 26049 2472 26049 2472 6 n_162
rlabel m2contact 26097 3960 26097 3960 6 n_13
rlabel m2contact 26121 2328 26121 2328 6 stateSub[2]
rlabel m2contact 26145 6792 26145 6792 6 n_33
rlabel m2contact 26193 3912 26193 3912 6 n_112
rlabel m2contact 26217 3816 26217 3816 6 n_237
rlabel m2contact 26241 5304 26241 5304 6 n_31
rlabel m2contact 26289 2736 26289 2736 6 n_170
rlabel m2contact 26313 5016 26313 5016 6 n_172
rlabel m2contact 26337 3528 26337 3528 6 n_186
rlabel m2contact 26337 3168 26337 3168 6 n_193
rlabel m2contact 26361 6240 26361 6240 6 n_116
rlabel m2contact 26385 2832 26385 2832 6 stateSub[1]
rlabel m2contact 26409 2712 26409 2712 6 n_156
rlabel m2contact 26433 4728 26433 4728 6 n_190
rlabel m2contact 26481 6000 26481 6000 6 n_265
rlabel m2contact 26529 3072 26529 3072 6 n_225
rlabel m2contact 26529 1992 26529 1992 6 n_326
rlabel m2contact 26553 3672 26553 3672 6 n_218
rlabel m2contact 26553 3312 26553 3312 6 n_352
rlabel m2contact 26577 6120 26577 6120 6 n_367
rlabel m2contact 26601 3576 26601 3576 6 n_251
rlabel m2contact 26601 3552 26601 3552 6 PcSel[1]
rlabel m2contact 26625 3552 26625 3552 6 PcSel[1]
rlabel m2contact 26625 5928 26625 5928 6 PcSel[1]
rlabel m2contact 26649 6312 26649 6312 6 n_159
rlabel m2contact 26649 4752 26649 4752 6 n_241
rlabel m2contact 26673 3624 26673 3624 6 n_240
rlabel m2contact 26697 4776 26697 4776 6 n_65
rlabel m2contact 26697 4728 26697 4728 6 n_242
rlabel m2contact 26721 4752 26721 4752 6 n_241
rlabel m2contact 26721 7320 26721 7320 6 n_241
rlabel m2contact 26745 5088 26745 5088 6 n_375
rlabel m2contact 26769 7632 26769 7632 6 n_79
rlabel m2contact 26793 6432 26793 6432 6 n_86
rlabel m2contact 26817 5856 26817 5856 6 n_217
rlabel m2contact 26841 4176 26841 4176 6 n_80
rlabel m2contact 26865 2616 26865 2616 6 n_23
rlabel m2contact 26889 5496 26889 5496 6 OpcodeCondIn[3]
rlabel m2contact 26889 5976 26889 5976 6 n_72
rlabel m2contact 26913 5664 26913 5664 6 n_38
rlabel m2contact 26913 5688 26913 5688 6 n_64
rlabel m2contact 26937 1776 26937 1776 6 n_36
rlabel m2contact 26961 7392 26961 7392 6 n_152
rlabel m2contact 26961 4776 26961 4776 6 Flags[0]
rlabel m2contact 26985 4728 26985 4728 6 n_242
rlabel m2contact 26985 4824 26985 4824 6 n_242
rlabel m2contact 27009 3912 27009 3912 6 n_112
rlabel m2contact 27033 6912 27033 6912 6 OpcodeCondIn[4]
rlabel m2contact 27057 3456 27057 3456 6 n_28
rlabel m2contact 27081 1728 27081 1728 6 n_64
rlabel m2contact 27081 5688 27081 5688 6 n_64
rlabel m2contact 27105 7512 27105 7512 6 n_233
rlabel m2contact 27129 4920 27129 4920 6 n_151
rlabel m2contact 27153 4992 27153 4992 6 n_292
rlabel m2contact 27201 3600 27201 3600 6 n_210
rlabel m2contact 27225 6192 27225 6192 6 n_177
rlabel m2contact 27273 1848 27273 1848 6 n_250
rlabel m2contact 27321 4800 27321 4800 6 n_379
rlabel m2contact 27345 4776 27345 4776 6 Flags[0]
rlabel m2contact 27369 3144 27369 3144 6 n_381
rlabel m2contact 27417 3096 27417 3096 6 n_179
rlabel m2contact 27441 2568 27441 2568 6 n_262
rlabel m2contact 27465 5064 27465 5064 6 n_137
rlabel m2contact 27513 2088 27513 2088 6 RwSel[1]
rlabel m2contact 27537 1728 27537 1728 6 OpcodeCondIn[1]
rlabel m2contact 27537 4344 27537 4344 6 OpcodeCondIn[1]
rlabel m2contact 27561 1752 27561 1752 6 OpcodeCondIn[3]
rlabel m2contact 27561 5496 27561 5496 6 OpcodeCondIn[3]
rlabel m2contact 27585 1776 27585 1776 6 SysBus[2]
rlabel m2contact 27585 5280 27585 5280 6 SysBus[2]
rlabel m2contact 27609 1800 27609 1800 6 SysBus[3]
rlabel m2contact 27609 4680 27609 4680 6 SysBus[3]
rlabel m2contact 27633 1824 27633 1824 6 SysBus[0]
rlabel m2contact 27633 6816 27633 6816 6 SysBus[0]
rlabel m2contact 2049 8897 2049 8897 4 IrWe
rlabel m2contact 2217 8801 2217 8801 4 CFlag
rlabel m2contact 2385 8921 2385 8921 4 AluEn
rlabel metal2 2403 8921 2403 8921 4 AluEn
rlabel m2contact 3249 8921 3249 8921 4 Rs1Sel[1]
rlabel m2contact 3681 8777 3681 8777 4 AluOR[0]
rlabel m2contact 3945 8945 3945 8945 4 AluWe
rlabel metal2 3963 8945 3963 8945 4 AluWe
rlabel m2contact 4137 8945 4137 8945 4 LrSel
rlabel m2contact 6177 8753 6177 8753 4 Op2Sel[1]
rlabel m2contact 7281 8969 7281 8969 4 LrEn
rlabel m2contact 7713 8729 7713 8729 4 Op2Sel[0]
rlabel m2contact 9249 8705 9249 8705 4 ImmSel
rlabel m2contact 9297 8681 9297 8681 4 RegWe
rlabel m2contact 9897 8993 9897 8993 4 PcSel[0]
rlabel m2contact 10785 8657 10785 8657 4 Op1Sel
rlabel m2contact 11217 8825 11217 8825 4 nWait
rlabel m2contact 11721 8657 11721 8657 4 Op1Sel
rlabel m2contact 12321 8825 12321 8825 4 PcWe
rlabel m2contact 12369 8657 12369 8657 4 Rs1Sel[0]
rlabel m2contact 13353 8801 13353 8801 4 CFlag
rlabel m2contact 13857 8633 13857 8633 4 PcEn
rlabel m2contact 14841 8633 14841 8633 6 PcEn
rlabel m2contact 15393 8633 15393 8633 6 PcSel[2]
rlabel m2contact 16041 9017 16041 9017 6 PcSel[1]
rlabel metal2 16059 9017 16059 9017 6 PcSel[1]
rlabel m2contact 16941 8993 16941 8993 6 PcSel[0]
rlabel m2contact 17145 8753 17145 8753 6 Op2Sel[1]
rlabel m2contact 17289 8825 17289 8825 6 PcWe
rlabel m2contact 17529 8825 17529 8825 6 MemEn
rlabel m2contact 18465 8969 18465 8969 6 LrEn
rlabel m2contact 18705 8801 18705 8801 6 CFlag
rlabel m2contact 19185 8705 19185 8705 6 ImmSel
rlabel m2contact 19233 8753 19233 8753 6 WdSel
rlabel m2contact 19989 8753 19989 8753 6 WdSel
rlabel m2contact 20265 8849 20265 8849 6 nME
rlabel m2contact 21105 8633 21105 8633 6 PcSel[2]
rlabel m2contact 22737 8753 22737 8753 6 LrWe
rlabel metal2 22755 8753 22755 8753 6 LrWe
rlabel m2contact 22785 8873 22785 8873 6 ALE
rlabel m2contact 23037 8945 23037 8945 6 LrSel
rlabel m2contact 23361 8729 23361 8729 6 Op2Sel[0]
rlabel m2contact 24561 8897 24561 8897 6 IrWe
rlabel m2contact 25833 8753 25833 8753 6 RwSel[0]
rlabel m2contact 26085 8825 26085 8825 6 MemEn
rlabel m2contact 27513 8825 27513 8825 6 RwSel[1]
rlabel m2contact 27537 8633 27537 8633 6 AluOR[0]
rlabel m2contact 27537 8777 27537 8777 6 AluOR[0]
rlabel m2contact 27561 8705 27561 8705 6 Rs1Sel[1]
rlabel m2contact 27561 8921 27561 8921 6 Rs1Sel[1]
rlabel m2contact 27585 8729 27585 8729 6 RwSel[0]
rlabel m2contact 27585 8753 27585 8753 6 RwSel[0]
rlabel m2contact 27585 8777 27585 8777 6 CFlag
rlabel m2contact 27585 8801 27585 8801 6 CFlag
rlabel m2contact 27609 8681 27609 8681 6 RegWe
rlabel m2contact 27609 8753 27609 8753 6 RegWe
rlabel m2contact 27633 8681 27633 8681 6 RwSel[1]
rlabel m2contact 27633 8825 27633 8825 6 RwSel[1]
<< end >>
