../../Design/Implementation/verilog/behavioural/opcodes.svh