../../../Design/Implementation/verilog/behavioural/io_serial.sv