magic
tech c035u
timestamp 1398682356
<< metal1 >>
rect -28 17559 0 17569
rect -28 17536 0 17546
rect -28 17498 0 17523
rect -28 16853 0 16878
rect -28 16830 0 16840
rect -28 16807 0 16817
rect -28 16784 0 16794
rect -28 16761 0 16771
rect -28 16694 0 16704
rect 1008 16672 1030 16682
rect -28 16448 0 16458
rect -28 16425 0 16435
rect -28 16387 0 16412
rect -28 15742 0 15767
rect -28 15719 0 15729
rect -28 15696 0 15706
rect -28 15673 0 15683
rect -28 15650 0 15660
rect -28 15583 0 15593
rect 1008 15561 1030 15571
rect -28 15337 0 15347
rect -28 15314 0 15324
rect -28 15276 0 15301
rect -28 14631 0 14656
rect -28 14608 0 14618
rect -28 14585 0 14595
rect -28 14562 0 14572
rect -28 14539 0 14549
rect -28 14472 0 14482
rect 1008 14450 1030 14460
rect -28 14226 0 14236
rect -28 14203 0 14213
rect -28 14165 0 14190
rect -28 13520 0 13545
rect -28 13497 0 13507
rect -28 13474 0 13484
rect -28 13451 0 13461
rect -28 13428 0 13438
rect -28 13361 0 13371
rect 1008 13339 1030 13349
rect -28 13115 0 13125
rect -28 13092 0 13102
rect -28 13054 0 13079
rect -28 12409 0 12434
rect -28 12386 0 12396
rect -28 12363 0 12373
rect -28 12340 0 12350
rect -28 12317 0 12327
rect -28 12250 0 12260
rect 1008 12228 1030 12238
rect -28 12004 0 12014
rect -28 11981 0 11991
rect -28 11943 0 11968
rect -28 11298 0 11323
rect -28 11275 0 11285
rect -28 11252 0 11262
rect -28 11229 0 11239
rect -28 11206 0 11216
rect -28 11139 0 11149
rect 1008 11117 1030 11127
rect -28 10893 0 10903
rect -28 10870 0 10880
rect -28 10832 0 10857
rect -28 10187 0 10212
rect -28 10164 0 10174
rect -28 10141 0 10151
rect -28 10118 0 10128
rect -28 10095 0 10105
rect -28 10028 0 10038
rect 1008 10006 1030 10016
rect -28 9782 0 9792
rect -28 9759 0 9769
rect -28 9721 0 9746
rect -28 9076 0 9101
rect -28 9053 0 9063
rect -28 9030 0 9040
rect -28 9007 0 9017
rect -28 8984 0 8994
rect -28 8917 0 8927
rect 1008 8895 1030 8905
rect -28 8671 0 8681
rect -28 8648 0 8658
rect -28 8610 0 8635
rect -28 7965 0 7990
rect -28 7942 0 7952
rect -28 7919 0 7929
rect -28 7896 0 7906
rect -28 7873 0 7883
rect -28 7806 0 7816
rect 1008 7784 1030 7794
rect -28 7560 0 7570
rect -28 7537 0 7547
rect -28 7499 0 7524
rect -28 6854 0 6879
rect -28 6831 0 6841
rect -28 6808 0 6818
rect -28 6785 0 6795
rect -28 6762 0 6772
rect -28 6695 0 6705
rect 1008 6673 1030 6683
rect -28 6449 0 6459
rect -28 6426 0 6436
rect -28 6388 0 6413
rect -28 5743 0 5768
rect -28 5720 0 5730
rect -28 5697 0 5707
rect -28 5674 0 5684
rect -28 5651 0 5661
rect -28 5584 0 5594
rect 1008 5562 1030 5572
rect -28 5338 0 5348
rect -28 5315 0 5325
rect -28 5277 0 5302
rect -28 4632 0 4657
rect -28 4609 0 4619
rect -28 4586 0 4596
rect -28 4563 0 4573
rect -28 4540 0 4550
rect -28 4473 0 4483
rect 1008 4451 1030 4461
rect -28 4227 0 4237
rect -28 4204 0 4214
rect -28 4166 0 4191
rect -28 3521 0 3546
rect -28 3498 0 3508
rect -28 3475 0 3485
rect -28 3452 0 3462
rect -28 3429 0 3439
rect -28 3362 0 3372
rect 1008 3340 1030 3350
rect -28 3116 0 3126
rect -28 3093 0 3103
rect -28 3055 0 3080
rect -28 2410 0 2435
rect -28 2387 0 2397
rect -28 2364 0 2374
rect -28 2341 0 2351
rect -28 2318 0 2328
rect -28 2251 0 2261
rect 1008 2229 1030 2239
rect -28 2005 0 2015
rect -28 1982 0 1992
rect -28 1944 0 1969
rect -28 1299 0 1324
rect -28 1276 0 1286
rect -28 1253 0 1263
rect -28 1230 0 1240
rect -28 1207 0 1217
rect -28 1140 0 1150
rect 1008 1118 1030 1128
rect -28 894 0 904
rect -28 871 0 881
rect -28 833 0 858
rect -28 188 0 213
rect -28 165 0 175
rect -28 142 0 152
rect -28 119 0 129
rect -28 96 0 106
rect -28 29 0 39
rect 1008 7 1030 17
<< metal2 >>
rect 72 17776 84 17807
rect 864 17776 876 17807
use IrAA IrAA_0
array 0 0 1008 0 7 1111
timestamp 1397224710
transform 1 0 0 0 1 8888
box 0 0 1008 1111
use IrBA IrBA_0
array 0 0 1008 0 2 1111
timestamp 1397224710
transform 1 0 0 0 1 5555
box 0 0 1008 1111
use IrBB IrBB_0
array 0 0 1008 0 4 1111
timestamp 1397224710
transform 1 0 0 0 1 0
box 0 0 1008 1111
<< labels >>
rlabel metal1 -28 165 -28 175 3 Clock
rlabel metal1 -28 1276 -28 1286 3 Clock
rlabel metal1 -28 2387 -28 2397 3 Clock
rlabel metal1 -28 3498 -28 3508 3 Clock
rlabel metal1 -28 4609 -28 4619 3 Clock
rlabel metal1 -28 5720 -28 5730 3 Clock
rlabel metal1 -28 6831 -28 6841 3 Clock
rlabel metal1 -28 7942 -28 7952 3 Clock
rlabel metal1 -28 9053 -28 9063 3 Clock
rlabel metal1 -28 10164 -28 10174 3 Clock
rlabel metal1 -28 11275 -28 11285 3 Clock
rlabel metal1 -28 12386 -28 12396 3 Clock
rlabel metal1 -28 13497 -28 13507 3 Clock
rlabel metal1 -28 14608 -28 14618 3 Clock
rlabel metal1 -28 15719 -28 15729 3 Clock
rlabel metal1 -28 16830 -28 16840 3 Clock
rlabel metal1 -28 119 -28 129 2 nReset
rlabel metal1 -28 1230 -28 1240 2 nReset
rlabel metal1 -28 2341 -28 2351 2 nReset
rlabel metal1 -28 3452 -28 3462 2 nReset
rlabel metal1 -28 4563 -28 4573 2 nReset
rlabel metal1 -28 5674 -28 5684 2 nReset
rlabel metal1 -28 6785 -28 6795 2 nReset
rlabel metal1 -28 7896 -28 7906 2 nReset
rlabel metal1 -28 9007 -28 9017 2 nReset
rlabel metal1 -28 10118 -28 10128 2 nReset
rlabel metal1 -28 11229 -28 11239 2 nReset
rlabel metal1 -28 12340 -28 12350 2 nReset
rlabel metal1 -28 13451 -28 13461 2 nReset
rlabel metal1 -28 14562 -28 14572 2 nReset
rlabel metal1 -28 15673 -28 15683 2 nReset
rlabel metal1 -28 16784 -28 16794 2 nReset
rlabel metal1 -28 142 -28 152 3 Test
rlabel metal1 -28 1253 -28 1263 3 Test
rlabel metal1 -28 2364 -28 2374 3 Test
rlabel metal1 -28 3475 -28 3485 3 Test
rlabel metal1 -28 4586 -28 4596 3 Test
rlabel metal1 -28 5697 -28 5707 3 Test
rlabel metal1 -28 6808 -28 6818 3 Test
rlabel metal1 -28 7919 -28 7929 3 Test
rlabel metal1 -28 9030 -28 9040 3 Test
rlabel metal1 -28 10141 -28 10151 3 Test
rlabel metal1 -28 11252 -28 11262 3 Test
rlabel metal1 -28 12363 -28 12373 3 Test
rlabel metal1 -28 13474 -28 13484 3 Test
rlabel metal1 -28 14585 -28 14595 3 Test
rlabel metal1 -28 15696 -28 15706 3 Test
rlabel metal1 -28 16807 -28 16817 3 Test
rlabel metal1 -28 188 -28 213 3 GND!
rlabel metal1 -28 1299 -28 1324 3 GND!
rlabel metal1 -28 2410 -28 2435 3 GND!
rlabel metal1 -28 3521 -28 3546 3 GND!
rlabel metal1 -28 4632 -28 4657 3 GND!
rlabel metal1 -28 5743 -28 5768 3 GND!
rlabel metal1 -28 6854 -28 6879 3 GND!
rlabel metal1 -28 7965 -28 7990 3 GND!
rlabel metal1 -28 9076 -28 9101 3 GND!
rlabel metal1 -28 10187 -28 10212 3 GND!
rlabel metal1 -28 11298 -28 11323 3 GND!
rlabel metal1 -28 12409 -28 12434 3 GND!
rlabel metal1 -28 13520 -28 13545 3 GND!
rlabel metal1 -28 14631 -28 14656 3 GND!
rlabel metal1 -28 15742 -28 15767 3 GND!
rlabel metal1 -28 16853 -28 16878 3 GND!
rlabel metal1 -28 833 -28 858 3 Vdd!
rlabel metal1 -28 1944 -28 1969 3 Vdd!
rlabel metal1 -28 3055 -28 3080 3 Vdd!
rlabel metal1 -28 4166 -28 4191 3 Vdd!
rlabel metal1 -28 5277 -28 5302 3 Vdd!
rlabel metal1 -28 6388 -28 6413 3 Vdd!
rlabel metal1 -28 7499 -28 7524 3 Vdd!
rlabel metal1 -28 8610 -28 8635 3 Vdd!
rlabel metal1 -28 9721 -28 9746 3 Vdd!
rlabel metal1 -28 10832 -28 10857 3 Vdd!
rlabel metal1 -28 11943 -28 11968 3 Vdd!
rlabel metal1 -28 13054 -28 13079 3 Vdd!
rlabel metal1 -28 14165 -28 14190 3 Vdd!
rlabel metal1 -28 15276 -28 15301 3 Vdd!
rlabel metal1 -28 16387 -28 16412 3 Vdd!
rlabel metal1 -28 17498 -28 17523 3 Vdd!
rlabel metal1 -28 871 -28 881 3 SDI
rlabel metal1 -28 1982 -28 1992 3 SDI
rlabel metal1 -28 3093 -28 3103 3 SDI
rlabel metal1 -28 4204 -28 4214 3 SDI
rlabel metal1 -28 5315 -28 5325 3 SDI
rlabel metal1 -28 6426 -28 6436 3 SDI
rlabel metal1 -28 7537 -28 7547 3 SDI
rlabel metal1 -28 8648 -28 8658 3 SDI
rlabel metal1 -28 9759 -28 9769 3 SDI
rlabel metal1 -28 10870 -28 10880 3 SDI
rlabel metal1 -28 11981 -28 11991 3 SDI
rlabel metal1 -28 13092 -28 13102 3 SDI
rlabel metal1 -28 14203 -28 14213 3 SDI
rlabel metal1 -28 15314 -28 15324 3 SDI
rlabel metal1 -28 16425 -28 16435 3 SDI
rlabel metal1 -28 17536 -28 17546 3 SDI
rlabel metal1 -28 894 -28 904 3 ScanReturn
rlabel metal1 -28 2005 -28 2015 3 ScanReturn
rlabel metal1 -28 3116 -28 3126 3 ScanReturn
rlabel metal1 -28 4227 -28 4237 3 ScanReturn
rlabel metal1 -28 5338 -28 5348 3 ScanReturn
rlabel metal1 -28 6449 -28 6459 3 ScanReturn
rlabel metal1 -28 7560 -28 7570 3 ScanReturn
rlabel metal1 -28 8671 -28 8681 3 ScanReturn
rlabel metal1 -28 9782 -28 9792 3 ScanReturn
rlabel metal1 -28 10893 -28 10903 3 ScanReturn
rlabel metal1 -28 12004 -28 12014 3 ScanReturn
rlabel metal1 -28 13115 -28 13125 3 ScanReturn
rlabel metal1 -28 14226 -28 14236 3 ScanReturn
rlabel metal1 -28 15337 -28 15347 3 ScanReturn
rlabel metal1 -28 16448 -28 16458 3 ScanReturn
rlabel metal1 -28 17559 -28 17569 3 ScanReturn
rlabel metal1 1030 7 1030 17 7 Imm[0]
rlabel metal1 1030 1118 1030 1128 7 Imm[1]
rlabel metal1 1030 2229 1030 2239 7 Imm[2]
rlabel metal1 1030 3340 1030 3350 7 Imm[3]
rlabel metal1 1030 4451 1030 4461 7 Imm[4]
rlabel metal1 1030 5562 1030 5572 7 Imm[5]
rlabel metal1 1030 6673 1030 6683 7 Imm[6]
rlabel metal1 1030 7784 1030 7794 7 Imm[7]
rlabel metal1 1030 8895 1030 8905 7 Imm[8]
rlabel metal1 1030 10006 1030 10016 7 Imm[9]
rlabel metal1 1030 11117 1030 11127 7 Imm[10]
rlabel metal1 1030 12228 1030 12238 7 Imm[11]
rlabel metal1 1030 13339 1030 13349 7 Imm[12]
rlabel metal1 1030 14450 1030 14460 7 Imm[13]
rlabel metal1 1030 15561 1030 15571 7 Imm[14]
rlabel metal1 1030 16672 1030 16682 7 Imm[15]
rlabel metal1 -28 29 -28 39 3 SysBus[0]
rlabel metal1 -28 1140 -28 1150 3 SysBus[1]
rlabel metal1 -28 2251 -28 2261 3 SysBus[2]
rlabel metal1 -28 3362 -28 3372 3 SysBus[3]
rlabel metal1 -28 4473 -28 4483 3 SysBus[4]
rlabel metal1 -28 5584 -28 5594 3 SysBus[5]
rlabel metal1 -28 6695 -28 6705 3 SysBus[6]
rlabel metal1 -28 7806 -28 7816 3 SysBus[7]
rlabel metal1 -28 8917 -28 8927 3 SysBus[8]
rlabel metal1 -28 10028 -28 10038 3 SysBus[9]
rlabel metal1 -28 11139 -28 11149 3 SysBus[10]
rlabel metal1 -28 12250 -28 12260 3 SysBus[11]
rlabel metal1 -28 13361 -28 13371 3 SysBus[12]
rlabel metal1 -28 14472 -28 14482 3 SysBus[13]
rlabel metal1 -28 15583 -28 15593 3 SysBus[14]
rlabel metal1 -28 16694 -28 16704 3 SysBus[15]
rlabel metal1 -28 96 -28 106 3 Ir[0]
rlabel metal1 -28 1207 -28 1217 3 Ir[1]
rlabel metal1 -28 2318 -28 2328 3 Ir[2]
rlabel metal1 -28 3429 -28 3439 3 Ir[3]
rlabel metal1 -28 4540 -28 4550 3 Ir[4]
rlabel metal1 -28 5651 -28 5661 3 Ir[5]
rlabel metal1 -28 6762 -28 6772 3 Ir[6]
rlabel metal1 -28 7873 -28 7883 3 Ir[7]
rlabel metal1 -28 8984 -28 8994 3 Ir[8]
rlabel metal1 -28 10095 -28 10105 3 Ir[9]
rlabel metal1 -28 11206 -28 11216 3 Ir[10]
rlabel metal1 -28 12317 -28 12327 3 Ir[11]
rlabel metal1 -28 13428 -28 13438 3 Ir[12]
rlabel metal1 -28 14539 -28 14549 3 Ir[13]
rlabel metal1 -28 15650 -28 15660 3 Ir[14]
rlabel metal1 -28 16761 -28 16771 3 Ir[15]
rlabel metal2 864 17807 876 17807 5 ImmSel
rlabel metal2 72 17807 84 17807 5 IrWe
<< end >>
