magic
tech c035u
timestamp 1394303457
<< metal1 >>
rect 4050 1062 5500 1072
rect 5514 1062 14837 1072
rect 0 155 1469 165
rect 0 95 1492 105
rect 1506 95 5380 105
rect 5394 95 5548 105
rect 5562 95 14841 105
rect 2442 73 14841 83
rect 5106 51 14841 61
rect 14586 29 14841 39
rect 14802 7 14841 17
<< m2contact >>
rect 4036 1060 4050 1074
rect 5500 1060 5514 1074
rect 1492 93 1506 107
rect 5380 93 5394 107
rect 5548 93 5562 107
rect 2428 71 2442 85
rect 5092 49 5106 63
rect 14572 27 14586 41
rect 14788 5 14802 19
<< metal2 >>
rect 5 970 205 1079
rect 221 970 233 1079
rect 245 970 257 1079
rect 269 970 281 1079
rect 293 970 305 1079
rect 1541 1050 1553 1079
rect 2213 1050 2225 1079
rect 2261 1050 2273 1079
rect 2333 1050 2345 1079
rect 2693 1050 2705 1079
rect 2837 1050 2849 1079
rect 3053 1050 3065 1079
rect 3797 1050 3809 1079
rect 3965 1050 3977 1079
rect 4037 1050 4049 1060
rect 4349 1050 4361 1079
rect 4565 1050 4577 1079
rect 5309 1050 5321 1079
rect 5477 970 5489 1079
rect 5501 970 5513 1060
rect 5573 1050 5657 1062
rect 5693 1050 5705 1079
rect 6437 1050 6449 1079
rect 6653 1050 6665 1079
rect 6845 1050 6857 1079
rect 7589 1050 7601 1079
rect 7805 1050 7817 1079
rect 5573 970 5585 1050
rect 7997 1049 8009 1079
rect 8741 1050 8753 1079
rect 8957 1050 8969 1079
rect 9149 1050 9161 1079
rect 9893 1050 9905 1079
rect 10109 1050 10121 1079
rect 10301 1050 10313 1079
rect 11045 1050 11057 1079
rect 11261 1050 11273 1079
rect 11453 1050 11465 1079
rect 12197 1050 12209 1079
rect 12413 1050 12425 1079
rect 12605 1050 12617 1079
rect 13349 1050 13361 1079
rect 13565 1050 13577 1079
rect 13757 1049 13769 1079
rect 14501 1050 14513 1079
rect 14717 1049 14729 1079
rect 5 0 205 171
rect 221 0 233 171
rect 245 0 257 171
rect 269 0 281 171
rect 293 0 305 171
rect 1493 107 1505 111
rect 1541 0 1553 113
rect 2213 0 2225 112
rect 2261 0 2273 111
rect 2333 0 2345 111
rect 2429 85 2441 111
rect 2693 0 2705 111
rect 2837 0 2849 111
rect 3053 0 3065 111
rect 3797 0 3809 111
rect 3965 0 3977 114
rect 4349 0 4361 113
rect 4565 0 4577 113
rect 5093 63 5105 111
rect 5309 0 5321 111
rect 5381 107 5393 111
rect 5477 0 5489 171
rect 5549 107 5561 171
rect 5693 0 5705 122
rect 6437 0 6449 111
rect 6653 0 6665 111
rect 6845 0 6857 111
rect 7589 0 7601 111
rect 7805 0 7817 111
rect 7997 0 8009 111
rect 8741 0 8753 111
rect 8957 0 8969 111
rect 9149 0 9161 111
rect 9893 0 9905 111
rect 10109 0 10121 111
rect 10301 0 10313 111
rect 11045 0 11057 111
rect 11261 0 11273 111
rect 11453 0 11465 111
rect 12197 0 12209 112
rect 12413 0 12425 111
rect 12605 0 12617 112
rect 13349 0 13361 111
rect 13565 0 13577 111
rect 13757 0 13769 111
rect 14501 0 14513 111
rect 14573 41 14585 111
rect 14717 0 14729 111
rect 14789 19 14801 112
use leftbuf  leftbuf_0
timestamp 1386242881
transform 1 0 5 0 1 171
box 0 0 1464 799
use IrAA  IrAA_0
timestamp 1394294731
transform 1 0 1469 0 1 111
box 0 0 1008 939
use Pc_slice  Pc_slice_0
timestamp 1394294966
transform 1 0 2477 0 1 111
box 0 0 2952 939
use mux2  mux2_0
timestamp 1386235218
transform 1 0 5429 0 1 171
box 0 0 192 799
use regBlock_slice  regBlock_slice_0
timestamp 1394295027
transform 1 0 5621 0 1 111
box 0 0 9216 939
<< labels >>
rlabel metal1 5573 100 5573 100 1 SysBus
rlabel metal1 14835 1067 14835 1067 6 AluOut
rlabel metal1 14830 34 14830 34 1 Rd1
rlabel metal1 14832 11 14832 11 1 Rd2
rlabel metal2 5 0 205 0 1 Vdd!
rlabel metal2 221 0 233 0 1 SDI
rlabel metal2 245 0 257 0 1 Test
rlabel metal2 269 0 281 0 1 Clock
rlabel metal2 293 0 305 0 1 nReset
rlabel metal2 2333 0 2345 0 1 ImmSel
rlabel metal2 2261 0 2273 0 1 Ext1
rlabel metal2 2213 0 2225 0 1 Ext0
rlabel metal2 2693 0 2705 0 1 PcIncCin
rlabel metal2 2837 0 2849 0 1 LrSel
rlabel metal2 3053 0 3065 0 1 LrWe
rlabel metal2 3797 0 3809 0 1 LrEn
rlabel metal2 3965 0 3977 0 1 PcSel[0]
rlabel metal2 4349 0 4361 0 1 PcSel[1]
rlabel metal2 4565 0 4577 0 1 PcWe
rlabel metal2 5309 0 5321 0 1 PcEn
rlabel metal2 5477 0 5489 0 1 WdSel
rlabel metal2 5693 0 5705 0 1 Rq[0]
rlabel metal2 6437 0 6449 0 1 Rs1[0]
rlabel metal2 6653 0 6665 0 1 Ps2[0]
rlabel metal2 6845 0 6857 0 1 Rw[1]
rlabel metal2 7589 0 7601 0 1 Rs1[1]
rlabel metal2 7805 0 7817 0 1 Rs2[1]
rlabel metal2 7997 0 8009 0 1 Rw[2]
rlabel metal2 8741 0 8753 0 1 Rs1[2]
rlabel metal2 8957 0 8969 0 1 Rs2[2]
rlabel metal2 9149 0 9161 0 1 Rw[3]
rlabel metal2 9893 0 9905 0 1 Rs1[3]
rlabel metal2 10109 0 10121 0 1 Rs2[3]
rlabel metal2 10301 0 10313 0 1 Rw[4]
rlabel metal2 11045 0 11057 0 1 Rs1[4]
rlabel metal2 11261 0 11273 0 1 Rs2[4]
rlabel metal2 11453 0 11465 0 1 Rw[5]
rlabel metal2 12197 0 12209 0 1 Rs1[5]
rlabel metal2 12413 0 12425 0 1 Rs2[5]
rlabel metal2 12605 0 12617 0 1 Rw[6]
rlabel metal2 13349 0 13361 0 1 Rs1[6]
rlabel metal2 13565 0 13577 0 1 Rs2[6]
rlabel metal2 13757 0 13769 0 1 Rw[7]
rlabel metal2 14501 0 14513 0 1 Rs1[7]
rlabel metal2 14717 0 14729 0 1 Rs2[7]
rlabel metal2 1541 0 1553 0 1 IrWe
rlabel metal1 14829 100 14829 100 1 SysBus
rlabel metal1 14830 78 14830 78 1 Imm
rlabel metal1 14831 56 14831 56 1 Pc
rlabel metal2 14717 1079 14729 1079 5 Rs2[7]
rlabel metal2 14501 1079 14513 1079 5 Rs1[7]
rlabel metal2 13757 1079 13769 1079 5 Rw[7]
rlabel metal2 13565 1079 13577 1079 5 Rs2[6]
rlabel metal2 13349 1079 13361 1079 5 Rs1[6]
rlabel metal2 12605 1079 12617 1079 5 Rw[6]
rlabel metal2 12197 1079 12209 1079 5 Rs1[5]
rlabel metal2 12413 1079 12425 1079 5 Rs2[5]
rlabel metal2 11453 1079 11465 1079 5 Rw[5]
rlabel metal2 11261 1079 11273 1079 5 Rs2[4]
rlabel metal2 11045 1079 11057 1079 5 Rs1[4]
rlabel metal2 10301 1079 10313 1079 5 Rw[4]
rlabel metal2 10109 1079 10121 1079 5 Rs2[3]
rlabel metal2 9893 1079 9905 1079 5 Rs1[3]
rlabel metal2 9149 1079 9161 1079 5 Rw[3]
rlabel metal2 8957 1079 8969 1079 5 Rs2[2]
rlabel metal2 8741 1079 8753 1079 5 Rs1[2]
rlabel metal2 7997 1079 8009 1079 5 Rw[2]
rlabel metal2 7805 1079 7817 1079 5 Rs2[1]
rlabel metal2 7589 1079 7601 1079 5 Rs1[1]
rlabel metal2 6845 1079 6857 1079 5 Rw[1]
rlabel metal2 6653 1079 6665 1079 5 Rs2[0]
rlabel metal2 6437 1079 6449 1079 5 Rs1[0]
rlabel metal2 5693 1079 5705 1079 5 Rw[0]
rlabel metal2 5477 1079 5489 1079 5 WdSel
rlabel metal2 5309 1079 5321 1079 5 PcEn
rlabel metal2 4565 1079 4577 1079 5 PcWe
rlabel metal2 4349 1079 4361 1079 5 PcSel[1]
rlabel metal2 3965 1079 3977 1079 5 PcSel[0]
rlabel metal2 3797 1079 3809 1079 5 LrEn
rlabel metal2 3053 1079 3065 1079 5 LrWe
rlabel metal2 2837 1079 2849 1079 5 LrSel
rlabel metal2 2693 1079 2705 1079 5 PcIncCout
rlabel metal2 2333 1079 2345 1079 5 ImmSel
rlabel metal2 2261 1079 2273 1079 5 Ext1
rlabel metal2 2213 1079 2225 1079 5 Ext0
rlabel metal2 1541 1079 1553 1079 5 IrWe
rlabel metal2 5 1079 205 1079 5 Vdd!
rlabel metal2 221 1079 233 1079 5 SDO
rlabel metal2 245 1079 257 1079 5 Test
rlabel metal2 269 1079 281 1079 5 Clock
rlabel metal2 293 1079 305 1079 5 nReset
rlabel metal1 0 95 0 105 3 SysBus
rlabel metal1 0 155 0 165 3 Ir
<< end >>
