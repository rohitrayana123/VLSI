magic
tech c035u
timestamp 1394566734
<< nwell >>
rect 1464 941 3240 1339
rect 15048 941 15432 1339
rect 23034 941 23856 1339
<< pwell >>
rect 1464 540 3240 941
rect 15048 547 15432 941
rect 23034 540 23856 941
<< pohmic >>
rect 1464 616 1470 626
rect 3234 616 3240 626
rect 15048 616 15054 626
rect 15426 616 15432 626
rect 23034 616 23040 626
rect 23850 616 23856 626
<< nohmic >>
rect 1464 1276 1470 1286
rect 3234 1276 3240 1286
rect 15048 1276 15054 1286
rect 15426 1276 15432 1286
rect 23034 1276 23040 1286
rect 23850 1276 23856 1286
<< psubstratetap >>
rect 1470 616 3234 632
rect 15054 616 15426 632
rect 23040 616 23850 632
<< nsubstratetap >>
rect 1470 1270 3234 1286
rect 15054 1270 15426 1286
rect 23040 1270 23850 1286
<< metal1 >>
rect 3637 1734 6167 1744
rect 4069 1712 6143 1722
rect 4501 1690 6119 1700
rect 4933 1667 5903 1677
rect 5365 1646 5879 1656
rect 5797 1624 5855 1634
rect 4189 1520 5519 1530
rect 4237 1498 5471 1508
rect 3805 1476 5039 1486
rect 3757 1454 5087 1464
rect 3372 1432 4607 1442
rect 3325 1410 4655 1420
rect 3301 1388 3719 1398
rect 3733 1388 4151 1398
rect 4597 1388 5015 1398
rect 5029 1388 5447 1398
rect 3541 1366 3959 1376
rect 3973 1366 4391 1376
rect 4837 1366 5255 1376
rect 5269 1366 5687 1376
rect 3397 1344 3551 1354
rect 3829 1344 3983 1354
rect 4261 1344 4415 1354
rect 4693 1344 4847 1354
rect 5125 1344 5279 1354
rect 5557 1344 5711 1354
rect 1464 1322 3240 1332
rect 15048 1322 15432 1332
rect 23034 1322 23856 1332
rect 1464 1299 3240 1309
rect 15048 1299 15432 1309
rect 23034 1299 23856 1309
rect 1464 1270 1470 1286
rect 3234 1270 3240 1286
rect 1464 1261 3240 1270
rect 15048 1270 15054 1286
rect 15426 1270 15432 1286
rect 15048 1261 15432 1270
rect 23034 1270 23040 1286
rect 23850 1270 23856 1286
rect 23034 1261 23856 1270
rect 1464 632 3240 641
rect 1464 616 1470 632
rect 3234 616 3240 632
rect 15048 632 15432 641
rect 15048 616 15054 632
rect 15426 616 15432 632
rect 23034 632 23856 641
rect 23034 616 23040 632
rect 23850 616 23856 632
rect 1464 593 3240 603
rect 15048 593 15432 603
rect 1464 570 3240 580
rect 15048 570 15432 580
rect 1464 547 3240 557
rect 15048 547 15432 557
rect 20869 28 20903 38
rect 20917 28 20951 38
rect 20965 28 20999 38
rect 21013 28 21047 38
rect 21061 28 21095 38
rect 21109 28 21143 38
rect 21157 28 21191 38
rect 21205 28 21503 38
rect 21517 28 21551 38
rect 21565 28 21599 38
rect 21613 28 21647 38
rect 21661 28 21959 38
rect 21973 28 22007 38
rect 22021 28 22319 38
rect 22333 28 23976 38
<< m2contact >>
rect 3623 1732 3637 1746
rect 6167 1732 6181 1746
rect 4055 1710 4069 1724
rect 6143 1710 6157 1724
rect 4487 1688 4501 1702
rect 6119 1688 6133 1702
rect 4919 1665 4933 1679
rect 5903 1665 5917 1679
rect 5351 1643 5365 1657
rect 5879 1643 5893 1657
rect 5783 1622 5797 1636
rect 5855 1621 5869 1635
rect 4175 1518 4189 1532
rect 5519 1518 5533 1532
rect 4223 1496 4237 1510
rect 5471 1496 5485 1510
rect 3791 1474 3805 1488
rect 5039 1474 5053 1488
rect 3743 1452 3757 1466
rect 5087 1452 5101 1466
rect 3358 1430 3372 1444
rect 4607 1430 4621 1444
rect 3311 1408 3325 1422
rect 4655 1408 4669 1422
rect 3287 1386 3301 1400
rect 3719 1386 3733 1400
rect 4151 1386 4165 1400
rect 4583 1386 4597 1400
rect 5015 1386 5029 1400
rect 5447 1386 5461 1400
rect 3527 1364 3541 1378
rect 3959 1364 3973 1378
rect 4391 1364 4405 1378
rect 4823 1364 4837 1378
rect 5255 1364 5269 1378
rect 5687 1364 5701 1378
rect 3383 1342 3397 1356
rect 3551 1342 3565 1356
rect 3815 1342 3829 1356
rect 3983 1342 3997 1356
rect 4247 1342 4261 1356
rect 4415 1342 4429 1356
rect 4679 1342 4693 1356
rect 4847 1342 4861 1356
rect 5111 1342 5125 1356
rect 5279 1342 5293 1356
rect 5543 1342 5557 1356
rect 5711 1342 5725 1356
rect 20855 26 20869 40
rect 20903 26 20917 40
rect 20951 26 20965 40
rect 20999 26 21013 40
rect 21047 26 21061 40
rect 21095 26 21109 40
rect 21143 26 21157 40
rect 21191 26 21205 40
rect 21503 25 21517 39
rect 21551 25 21565 39
rect 21599 25 21613 39
rect 21647 25 21661 39
rect 21959 26 21973 40
rect 22007 26 22021 40
rect 22319 26 22333 40
rect 23976 26 23990 40
<< metal2 >>
rect 0 1339 200 1795
rect 216 1339 228 1795
rect 240 1339 252 1795
rect 264 1339 276 1795
rect 288 1339 300 1795
rect 3288 1400 3300 1795
rect 3312 1422 3324 1795
rect 3360 1444 3372 1795
rect 3288 1339 3300 1386
rect 3312 1339 3324 1408
rect 3360 1339 3372 1430
rect 3528 1378 3540 1795
rect 3384 1339 3396 1342
rect 3528 1339 3540 1364
rect 3552 1339 3564 1342
rect 3624 1339 3636 1732
rect 3744 1466 3756 1795
rect 3792 1488 3804 1795
rect 3720 1339 3732 1386
rect 3744 1339 3756 1452
rect 3792 1339 3804 1474
rect 3816 1339 3828 1342
rect 3960 1339 3972 1364
rect 3984 1339 3996 1342
rect 4056 1339 4068 1710
rect 4176 1532 4188 1795
rect 4152 1339 4164 1386
rect 4176 1339 4188 1518
rect 4224 1510 4236 1795
rect 4224 1339 4236 1496
rect 4248 1339 4260 1342
rect 4392 1339 4404 1364
rect 4416 1339 4428 1342
rect 4488 1339 4500 1688
rect 4584 1400 4596 1795
rect 4584 1339 4596 1386
rect 4608 1339 4620 1430
rect 4656 1339 4668 1408
rect 4824 1378 4836 1795
rect 4680 1339 4692 1342
rect 4824 1339 4836 1364
rect 4848 1339 4860 1342
rect 4920 1339 4932 1665
rect 5016 1339 5028 1386
rect 5040 1339 5052 1474
rect 5088 1339 5100 1452
rect 5112 1339 5124 1342
rect 5256 1339 5268 1364
rect 5280 1339 5292 1342
rect 5352 1339 5364 1643
rect 5448 1339 5460 1386
rect 5472 1339 5484 1496
rect 5520 1339 5532 1518
rect 5544 1339 5556 1342
rect 5688 1339 5700 1364
rect 5712 1339 5724 1342
rect 5784 1339 5796 1622
rect 5856 1618 5868 1621
rect 5880 1618 5892 1643
rect 5904 1618 5916 1665
rect 5954 1618 5966 1795
rect 6120 1618 6132 1688
rect 6144 1618 6156 1710
rect 6168 1618 6180 1732
rect 6264 1618 6276 1795
rect 6288 1618 6300 1795
rect 6312 1618 6324 1795
rect 15624 1624 15636 1795
rect 15744 1624 15756 1795
rect 15864 1624 15876 1795
rect 15984 1624 15996 1795
rect 16104 1624 16116 1795
rect 17280 1624 17292 1795
rect 17712 1624 17724 1795
rect 17904 1624 17916 1795
rect 17976 1624 17988 1795
rect 18072 1624 18084 1795
rect 21744 1624 21756 1795
rect 21960 1624 21972 1795
rect 22080 1624 22092 1795
rect 22200 1624 22212 1795
rect 22584 1624 22596 1795
rect 23976 1339 24176 1795
rect 0 0 200 540
rect 216 0 228 540
rect 240 0 252 540
rect 264 0 276 540
rect 288 0 300 540
rect 3456 530 3468 540
rect 3600 530 3612 540
rect 3456 518 3612 530
rect 3888 530 3900 540
rect 4032 530 4044 540
rect 3888 518 4044 530
rect 4320 530 4332 540
rect 4464 530 4476 540
rect 4320 518 4476 530
rect 4752 530 4764 540
rect 4896 530 4908 540
rect 4752 518 4908 530
rect 5184 530 5196 540
rect 5328 530 5340 540
rect 5184 518 5340 530
rect 5616 530 5628 540
rect 5760 530 5772 540
rect 5616 518 5772 530
rect 15504 0 15516 165
rect 15768 0 15780 165
rect 15936 0 15948 165
rect 16104 0 16116 165
rect 16128 0 16140 165
rect 16200 0 16212 165
rect 16416 0 16428 165
rect 16560 0 16572 165
rect 16896 0 16908 165
rect 17256 0 17268 165
rect 17664 0 17676 165
rect 18000 0 18012 165
rect 18312 0 18324 165
rect 18648 0 18660 165
rect 18768 0 18780 165
rect 18816 0 18828 165
rect 18984 0 18996 165
rect 20784 0 20796 165
rect 20809 0 20821 165
rect 20856 0 20868 26
rect 20904 0 20916 26
rect 20952 0 20964 26
rect 21000 0 21012 26
rect 21048 0 21060 26
rect 21096 0 21108 26
rect 21144 0 21156 26
rect 21168 0 21180 165
rect 21192 0 21204 26
rect 21432 0 21444 165
rect 21504 0 21516 25
rect 21552 0 21564 25
rect 21600 0 21612 25
rect 21648 0 21660 25
rect 21888 0 21900 165
rect 21960 0 21972 26
rect 22008 0 22020 26
rect 22248 0 22260 165
rect 22320 0 22332 26
rect 22608 0 22620 165
rect 22776 0 22788 165
rect 23016 73 23028 165
rect 23016 61 23748 73
rect 23736 0 23748 61
rect 23976 40 24176 540
rect 23990 26 24176 40
rect 23976 0 24176 26
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 0 0 1 540
box 0 0 1464 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 3240 0 1 540
box 0 0 192 799
use tiehigh tiehigh_3
timestamp 1386086759
transform 1 0 3432 0 1 540
box 0 0 48 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 3480 0 1 540
box 0 0 192 799
use mux2 mux2_8
timestamp 1386235218
transform 1 0 3672 0 1 540
box 0 0 192 799
use tiehigh tiehigh_4
timestamp 1386086759
transform 1 0 3864 0 1 540
box 0 0 48 799
use mux2 mux2_9
timestamp 1386235218
transform 1 0 3912 0 1 540
box 0 0 192 799
use mux2 mux2_10
timestamp 1386235218
transform 1 0 4104 0 1 540
box 0 0 192 799
use tiehigh tiehigh_5
timestamp 1386086759
transform 1 0 4296 0 1 540
box 0 0 48 799
use mux2 mux2_11
timestamp 1386235218
transform 1 0 4344 0 1 540
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4536 0 1 540
box 0 0 192 799
use tiehigh tiehigh_2
timestamp 1386086759
transform 1 0 4728 0 1 540
box 0 0 48 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 4776 0 1 540
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 4968 0 1 540
box 0 0 192 799
use tiehigh tiehigh_1
timestamp 1386086759
transform 1 0 5160 0 1 540
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 5208 0 1 540
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 5400 0 1 540
box 0 0 192 799
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 5592 0 1 540
box 0 0 48 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 5640 0 1 540
box 0 0 192 799
use regBlock_decoder regBlock_decoder_0
timestamp 1394493274
transform 1 0 5832 0 1 0
box 0 0 9216 1618
use ALUDecoder ALUDecoder_0
timestamp 1394559852
transform 1 0 15432 0 1 165
box 0 0 7602 1459
use rightend rightend_0
timestamp 1386235834
transform 1 0 23856 0 1 540
box 0 0 320 799
<< labels >>
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 240 1795 252 1795 1 Test
rlabel metal2 264 1795 276 1795 1 Clock
rlabel metal2 288 1795 300 1795 1 nReset
rlabel metal2 0 1795 200 1795 5 Vdd!
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 15624 1795 15636 1795 5 Ir[15]
rlabel metal2 15744 1795 15756 1795 5 Ir[14]
rlabel metal2 15864 1795 15876 1795 5 Ir[13]
rlabel metal2 15984 1795 15996 1795 5 Ir[12]
rlabel metal2 16104 1795 16116 1795 5 Ir[11]
rlabel metal2 17280 1795 17292 1795 5 CFlag
rlabel metal2 17712 1795 17724 1795 5 Flags[2]
rlabel metal2 17904 1795 17916 1795 5 Flags[1]
rlabel metal2 18072 1795 18084 1795 5 Flagss[0]
rlabel metal2 22200 1795 22212 1795 5 Ir[0]
rlabel metal2 22080 1795 22092 1795 5 Ir[1]
rlabel metal2 21960 1795 21972 1795 5 Ir[2]
rlabel metal2 21744 1795 21756 1795 5 Ir[3]
rlabel metal2 22584 1795 22596 1795 5 AluEn
rlabel metal2 22776 0 22788 0 1 LLI
rlabel metal2 22608 0 22620 0 1 ShOut
rlabel metal2 21888 0 21900 0 1 Sh2
rlabel metal2 20809 0 20821 0 1 ShR
rlabel metal2 22248 0 22260 0 1 Sh1
rlabel metal2 21432 0 21444 0 1 Sh4
rlabel metal2 20784 0 20796 0 1 Sh8
rlabel metal2 15504 0 15516 0 1 ZeroA
rlabel metal2 16200 0 16212 0 1 N
rlabel metal2 18648 0 18660 0 1 NOR
rlabel metal2 18816 0 18828 0 1 ShB
rlabel metal2 18768 0 18780 0 1 ASign
rlabel metal2 18984 0 18996 0 1 ShL
rlabel metal2 18000 0 18012 0 1 NOT
rlabel metal2 17664 0 17676 0 1 XOR
rlabel metal2 17256 0 17268 0 1 OR
rlabel metal2 16896 0 16908 0 1 AND
rlabel metal2 16560 0 16572 0 1 FAOut
rlabel metal2 16416 0 16428 0 1 nZ
rlabel metal2 16128 0 16140 0 1 COut
rlabel metal2 16104 0 16116 0 1 LastCIn
rlabel metal2 15936 0 15948 0 1 CIn_slice
rlabel metal2 15768 0 15780 0 1 SUB
rlabel metal2 18312 0 18324 0 1 NAND
rlabel metal2 21168 0 21180 0 1 ShInBit
rlabel metal2 4824 1795 4836 1795 5 RwSel[1]
rlabel metal2 4176 1795 4188 1795 5 Ir[8]
rlabel metal2 4224 1795 4236 1795 5 Ir[5]
rlabel metal2 3792 1795 3804 1795 5 Ir[6]
rlabel metal2 3744 1795 3756 1795 5 Ir[9]
rlabel metal2 3360 1795 3372 1795 5 Ir[7]
rlabel metal2 3312 1795 3324 1795 5 Ir[10]
rlabel metal2 3528 1795 3540 1795 5 Rs1Sel[1]
rlabel metal2 3288 1795 3300 1795 5 Rs1Sel[0]
rlabel metal2 5954 1795 5966 1795 5 RegWe
rlabel metal2 6312 1795 6324 1795 5 Ir[4]
rlabel metal2 6288 1795 6300 1795 5 Ir[3]
rlabel metal2 6264 1795 6276 1795 5 Ir[2]
rlabel metal2 17976 1795 17988 1795 5 Flags[3]
rlabel metal2 4584 1795 4596 1795 5 RwSel[0]
rlabel metal2 23976 1795 24176 1795 1 GND!
rlabel metal2 23736 0 23748 0 1 OutEn
rlabel metal2 21144 0 21156 0 5 Sh8G_R
rlabel metal2 21096 0 21108 0 5 Sh8F_R
rlabel metal2 21048 0 21060 0 5 Sh8E_R
rlabel metal2 21000 0 21012 0 5 Sh8D_R
rlabel metal2 20856 0 20868 0 5 Sh8A_R
rlabel metal2 20904 0 20916 0 5 Sh8B_R
rlabel metal2 20952 0 20964 0 5 Sh8C_R
rlabel metal2 21192 0 21204 0 5 Sh8H_R
rlabel metal2 21552 0 21564 0 5 Sh4A_R
rlabel metal2 21600 0 21612 0 5 Sh4B_R
rlabel metal2 21648 0 21660 0 5 Sh4C_R
rlabel metal2 21504 0 21516 0 5 Sh4Z_R
rlabel metal2 21960 0 21972 0 5 Sh2A_R
rlabel metal2 22008 0 22020 0 5 Sh2B_R
rlabel metal2 23978 0 24176 0 1 GND!
rlabel metal2 22320 0 22332 0 1 Sh1_R_In
rlabel metal2 216 1795 228 1795 5 SDO
<< end >>
