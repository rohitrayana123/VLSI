magic
tech c035u
timestamp 1398806367
<< nwell >>
rect 7104 665 7656 1063
<< pwell >>
rect 7104 264 7656 665
<< pohmic >>
rect 7104 340 7110 350
rect 7648 340 7656 350
<< nohmic >>
rect 7104 1000 7110 1010
rect 7648 1000 7656 1010
<< psubstratetap >>
rect 7136 604 7152 620
rect 7223 604 7239 620
rect 7310 604 7326 620
rect 7397 604 7413 620
rect 7484 604 7500 620
rect 7571 604 7587 620
rect 7110 340 7648 356
<< nsubstratetap >>
rect 7110 994 7648 1010
<< metal1 >>
rect 2005 1222 2159 1232
rect 2845 1222 2975 1232
rect 2989 1222 3119 1232
rect 3133 1222 3263 1232
rect 3277 1222 4271 1232
rect 4285 1222 4286 1232
rect 1909 1200 2063 1210
rect 2197 1200 2375 1210
rect 2413 1200 2471 1210
rect 3421 1200 3551 1210
rect 3565 1200 3695 1210
rect 3709 1200 4151 1210
rect 4165 1200 4583 1210
rect 6013 1201 6167 1211
rect 6675 1200 6709 1210
rect 7055 1200 7089 1210
rect 0 1178 623 1188
rect 709 1178 743 1188
rect 973 1178 1247 1188
rect 1573 1178 1607 1188
rect 1789 1178 2039 1188
rect 2101 1178 2231 1188
rect 2293 1178 2447 1188
rect 2701 1178 3911 1188
rect 4045 1178 4319 1188
rect 4333 1178 4439 1188
rect 4981 1178 5015 1188
rect 5653 1178 5687 1188
rect 5893 1178 5927 1188
rect 6109 1179 6143 1189
rect 6675 1176 6685 1200
rect 6709 1178 7055 1188
rect 7079 1176 7089 1200
rect 0 1156 503 1166
rect 517 1156 1871 1166
rect 1885 1156 1967 1166
rect 1981 1156 2735 1166
rect 2749 1156 2879 1166
rect 2893 1156 3311 1166
rect 3325 1156 3455 1166
rect 3469 1156 3743 1166
rect 3757 1156 4487 1166
rect 4501 1156 4775 1166
rect 4789 1156 5471 1166
rect 5485 1156 6935 1166
rect 0 1134 383 1144
rect 397 1134 1511 1144
rect 1525 1134 2255 1144
rect 2269 1134 2568 1144
rect 2582 1134 2855 1144
rect 2869 1134 2999 1144
rect 3013 1134 3719 1144
rect 3733 1134 4343 1144
rect 4357 1134 4463 1144
rect 4477 1134 4607 1144
rect 4621 1134 4751 1144
rect 4837 1134 5039 1144
rect 5101 1134 5135 1144
rect 5509 1134 5711 1144
rect 5749 1134 6047 1144
rect 6061 1134 6239 1144
rect 6253 1134 6359 1144
rect 6373 1134 6479 1144
rect 6829 1134 7031 1144
rect 0 1112 263 1122
rect 277 1112 1847 1122
rect 1861 1112 4007 1122
rect 4021 1112 4127 1122
rect 4141 1112 5447 1122
rect 5461 1112 5591 1122
rect 5605 1112 6767 1122
rect 6781 1112 6911 1122
rect 0 1090 143 1100
rect 157 1090 1487 1100
rect 1501 1090 1703 1100
rect 1717 1090 2351 1100
rect 2365 1090 3863 1100
rect 3877 1090 3983 1100
rect 3997 1090 4727 1100
rect 4741 1090 5423 1100
rect 5437 1090 5567 1100
rect 5581 1090 5807 1100
rect 5821 1090 6623 1100
rect 6637 1090 6887 1100
rect 0 1068 23 1078
rect 37 1068 1631 1078
rect 1645 1068 2543 1078
rect 2557 1068 3839 1078
rect 3853 1068 3959 1078
rect 3973 1068 4079 1078
rect 4093 1068 4199 1078
rect 4213 1068 5399 1078
rect 5413 1068 5543 1078
rect 5557 1068 6599 1078
rect 6613 1068 6743 1078
rect 6757 1068 6863 1078
rect 6973 1068 7007 1078
rect 7104 1046 7656 1056
rect 7104 1023 7656 1033
rect 7104 994 7110 1010
rect 7648 994 7656 1010
rect 7104 985 7656 994
rect 7136 365 7152 604
rect 7223 365 7239 604
rect 7310 365 7326 604
rect 7397 365 7413 604
rect 7484 365 7500 604
rect 7571 365 7587 604
rect 7104 356 7656 365
rect 7104 340 7110 356
rect 7648 340 7656 356
rect 7104 317 7656 327
rect 7104 294 7656 304
rect 7104 271 7656 281
rect 51 237 61 261
rect 85 249 1823 259
rect 1837 249 2327 259
rect 2341 249 5159 259
rect 5173 249 5783 259
rect 51 227 85 237
rect 205 227 4103 237
rect 4117 227 4223 237
rect 4237 227 4871 237
rect 5222 227 5279 237
rect 5365 227 5663 237
rect 325 205 1727 215
rect 1741 205 1943 215
rect 1957 205 2135 215
rect 2149 205 2591 215
rect 2605 205 3887 215
rect 3901 205 4247 215
rect 4261 205 5183 215
rect 5197 205 5831 215
rect 5845 205 6671 215
rect 445 183 2711 193
rect 2725 183 3143 193
rect 3157 183 3287 193
rect 3301 183 3431 193
rect 3445 183 3575 193
rect 3589 183 4895 193
rect 4909 183 5615 193
rect 5629 183 5951 193
rect 5965 183 6647 193
rect 6661 183 6791 193
rect 565 161 1535 171
rect 1549 161 1751 171
rect 1765 161 3023 171
rect 3037 161 3167 171
rect 3181 161 3599 171
rect 3613 161 4631 171
rect 4645 161 4919 171
rect 4933 161 5975 171
rect 349 139 767 149
rect 781 139 1127 149
rect 1141 139 2495 149
rect 3197 137 3215 147
rect 3277 139 3647 149
rect 4549 139 5303 149
rect 6565 139 6815 149
rect 661 117 2639 127
rect 3229 112 3263 122
rect 3321 117 3359 127
rect 3397 117 5208 127
rect 5365 117 6191 127
rect 7340 117 7377 127
rect 517 95 863 105
rect 997 95 1367 105
rect 1477 95 2927 105
rect 3349 93 3383 103
rect 3445 95 3791 105
rect 4693 95 7343 105
rect 7367 93 7377 117
rect 709 73 1151 83
rect 1837 73 3071 83
rect 3397 69 3431 79
rect 4405 73 5376 83
rect 6013 73 6311 83
rect 6445 69 6455 79
rect 685 51 935 61
rect 1141 51 1655 61
rect 2245 51 3183 61
rect 3565 51 5231 61
rect 51 29 85 39
rect 51 5 61 29
rect 781 29 1319 39
rect 2581 29 3307 39
rect 85 7 2783 17
rect 2893 7 3503 17
rect 5437 7 5471 17
rect 5485 7 5519 17
rect 5533 7 5567 17
rect 5581 7 5615 17
rect 5629 7 5663 17
rect 5677 7 5711 17
rect 5725 7 5759 17
rect 5773 7 6071 17
rect 6085 7 6119 17
rect 6133 7 6167 17
rect 6181 7 6215 17
rect 6229 7 6527 17
rect 6541 7 6575 17
rect 6589 7 6887 17
<< m2contact >>
rect 1991 1220 2005 1234
rect 2159 1220 2173 1234
rect 2831 1220 2845 1234
rect 2975 1220 2989 1234
rect 3119 1220 3133 1234
rect 3263 1220 3277 1234
rect 4271 1220 4285 1234
rect 1895 1198 1909 1212
rect 2063 1198 2077 1212
rect 2183 1198 2197 1212
rect 2375 1198 2389 1212
rect 2399 1198 2413 1212
rect 2471 1198 2485 1212
rect 3407 1198 3421 1212
rect 3551 1198 3565 1212
rect 3695 1198 3709 1212
rect 4151 1198 4165 1212
rect 4583 1198 4597 1212
rect 5999 1199 6013 1213
rect 6167 1199 6181 1213
rect 623 1176 637 1190
rect 695 1176 709 1190
rect 743 1176 757 1190
rect 959 1176 973 1190
rect 1247 1176 1261 1190
rect 1559 1176 1573 1190
rect 1607 1176 1621 1190
rect 1775 1176 1789 1190
rect 2039 1176 2053 1190
rect 2087 1177 2101 1191
rect 2231 1176 2245 1190
rect 2279 1176 2293 1190
rect 2447 1176 2461 1190
rect 2687 1176 2701 1190
rect 3911 1176 3925 1190
rect 4031 1176 4045 1190
rect 4319 1176 4333 1190
rect 4439 1176 4453 1190
rect 4967 1176 4981 1190
rect 5015 1176 5029 1190
rect 5639 1176 5653 1190
rect 5687 1176 5701 1190
rect 5879 1176 5893 1190
rect 5927 1176 5941 1190
rect 6095 1176 6109 1190
rect 6143 1176 6157 1190
rect 6695 1176 6709 1190
rect 7055 1176 7069 1190
rect 503 1154 517 1168
rect 1871 1154 1885 1168
rect 1967 1154 1981 1168
rect 2735 1154 2749 1168
rect 2879 1154 2893 1168
rect 3311 1154 3325 1168
rect 3455 1154 3469 1168
rect 3743 1154 3757 1168
rect 4487 1155 4501 1169
rect 4775 1153 4789 1167
rect 5471 1154 5485 1168
rect 6935 1154 6949 1168
rect 383 1132 397 1146
rect 1511 1132 1525 1146
rect 2255 1132 2269 1146
rect 2568 1132 2582 1146
rect 2855 1132 2869 1146
rect 2999 1132 3013 1146
rect 3719 1132 3733 1146
rect 4343 1132 4357 1146
rect 4463 1132 4477 1146
rect 4607 1132 4621 1146
rect 4751 1132 4765 1146
rect 4823 1132 4837 1146
rect 5039 1132 5053 1146
rect 5087 1132 5101 1146
rect 5135 1132 5149 1146
rect 5495 1132 5509 1146
rect 5711 1132 5725 1146
rect 5735 1132 5749 1146
rect 6047 1132 6061 1146
rect 6239 1132 6253 1146
rect 6359 1132 6373 1146
rect 6479 1132 6493 1146
rect 6815 1132 6829 1146
rect 7031 1132 7045 1146
rect 263 1110 277 1124
rect 1847 1110 1861 1124
rect 4007 1110 4021 1124
rect 4127 1110 4141 1124
rect 5447 1110 5461 1124
rect 5591 1110 5605 1124
rect 6767 1110 6781 1124
rect 6911 1110 6925 1124
rect 143 1088 157 1102
rect 1487 1088 1501 1102
rect 1703 1088 1717 1102
rect 2351 1088 2365 1102
rect 3863 1088 3877 1102
rect 3983 1088 3997 1102
rect 4727 1088 4741 1102
rect 5423 1088 5437 1102
rect 5567 1088 5581 1102
rect 5807 1088 5821 1102
rect 6623 1088 6637 1102
rect 6887 1088 6901 1102
rect 23 1066 37 1080
rect 1631 1066 1645 1080
rect 2543 1066 2557 1080
rect 3839 1066 3853 1080
rect 3959 1066 3973 1080
rect 4079 1066 4093 1080
rect 4199 1066 4213 1080
rect 5399 1066 5413 1080
rect 5543 1066 5557 1080
rect 6599 1066 6613 1080
rect 6743 1066 6757 1080
rect 6863 1066 6877 1080
rect 6959 1066 6973 1080
rect 7007 1066 7021 1080
rect 71 247 85 261
rect 1823 247 1837 261
rect 2327 247 2341 261
rect 5159 247 5173 261
rect 5783 247 5797 261
rect 191 225 205 239
rect 4103 225 4117 239
rect 4223 225 4237 239
rect 4871 225 4885 239
rect 5208 225 5222 239
rect 5279 225 5293 239
rect 5351 225 5365 239
rect 5663 225 5677 239
rect 311 203 325 217
rect 1727 203 1741 217
rect 1943 203 1957 217
rect 2135 203 2149 217
rect 2591 203 2605 217
rect 3887 203 3901 217
rect 4247 203 4261 217
rect 5183 204 5197 218
rect 5831 203 5845 217
rect 6671 203 6685 217
rect 431 181 445 195
rect 2711 181 2725 195
rect 3143 181 3157 195
rect 3287 181 3301 195
rect 3431 181 3445 195
rect 3575 181 3589 195
rect 4895 181 4909 195
rect 5615 181 5629 195
rect 5951 181 5965 195
rect 6647 181 6661 195
rect 6791 181 6805 195
rect 551 159 565 173
rect 1535 159 1549 173
rect 1751 159 1765 173
rect 3023 158 3037 172
rect 3167 159 3181 173
rect 3599 159 3613 173
rect 4631 159 4645 173
rect 4919 159 4933 173
rect 5975 159 5989 173
rect 335 137 349 151
rect 767 137 781 151
rect 1127 137 1141 151
rect 2495 137 2509 151
rect 3183 135 3197 149
rect 3215 134 3229 148
rect 3263 137 3277 151
rect 3647 137 3661 151
rect 4535 137 4549 151
rect 5303 137 5317 151
rect 6551 137 6565 151
rect 6815 137 6829 151
rect 647 115 661 129
rect 2639 115 2653 129
rect 3215 110 3229 124
rect 3263 110 3277 124
rect 3307 115 3321 129
rect 3359 115 3373 129
rect 3383 115 3397 129
rect 5208 115 5222 129
rect 5351 115 5365 129
rect 6191 115 6205 129
rect 503 93 517 107
rect 863 93 877 107
rect 983 93 997 107
rect 1367 93 1381 107
rect 1463 93 1477 107
rect 2927 93 2941 107
rect 3335 91 3349 105
rect 3383 91 3397 105
rect 3431 93 3445 107
rect 3791 93 3805 107
rect 4679 93 4693 107
rect 7343 93 7357 107
rect 695 71 709 85
rect 1151 71 1165 85
rect 1823 71 1837 85
rect 3071 72 3085 86
rect 3383 67 3397 81
rect 3431 67 3445 81
rect 4391 71 4405 85
rect 5376 71 5390 85
rect 5999 71 6013 85
rect 6311 71 6325 85
rect 6431 67 6445 81
rect 6455 67 6469 81
rect 671 49 685 63
rect 935 49 949 63
rect 1127 49 1141 63
rect 1655 49 1669 63
rect 2231 49 2245 63
rect 3183 49 3197 63
rect 3551 49 3565 63
rect 5231 49 5245 63
rect 767 27 781 41
rect 1319 27 1333 41
rect 2567 27 2581 41
rect 3307 27 3321 41
rect 71 5 85 19
rect 2783 5 2797 19
rect 2879 5 2893 19
rect 3503 5 3517 19
rect 5423 5 5437 19
rect 5471 5 5485 19
rect 5519 5 5533 19
rect 5567 5 5581 19
rect 5615 5 5629 19
rect 5663 5 5677 19
rect 5711 5 5725 19
rect 5759 5 5773 19
rect 6071 5 6085 19
rect 6119 5 6133 19
rect 6167 5 6181 19
rect 6215 5 6229 19
rect 6527 5 6541 19
rect 6575 5 6589 19
rect 6887 5 6901 19
<< metal2 >>
rect 24 1063 36 1066
rect 144 1063 156 1088
rect 264 1063 276 1110
rect 384 1063 396 1132
rect 504 1063 516 1154
rect 624 1063 636 1176
rect 696 1063 708 1176
rect 744 1063 756 1176
rect 960 1063 972 1176
rect 1056 1063 1068 1239
rect 1248 1190 1260 1239
rect 1248 1063 1260 1176
rect 1320 1063 1332 1239
rect 1416 1063 1428 1239
rect 1488 1063 1500 1088
rect 1512 1063 1524 1132
rect 1560 1063 1572 1176
rect 1608 1063 1620 1176
rect 1632 1063 1644 1066
rect 1704 1063 1716 1088
rect 1776 1063 1788 1176
rect 1848 1063 1860 1110
rect 1872 1063 1884 1154
rect 1896 1063 1908 1198
rect 1968 1063 1980 1154
rect 1992 1063 2004 1220
rect 2040 1063 2052 1176
rect 2064 1063 2076 1198
rect 2088 1063 2100 1177
rect 2160 1063 2172 1220
rect 2184 1063 2196 1198
rect 2232 1063 2244 1176
rect 2256 1063 2268 1132
rect 2280 1063 2292 1176
rect 2352 1063 2364 1088
rect 2376 1063 2388 1198
rect 2400 1063 2412 1198
rect 2448 1063 2460 1176
rect 2472 1063 2484 1198
rect 2544 1063 2556 1066
rect 2568 1063 2580 1132
rect 2688 1063 2700 1176
rect 2736 1063 2748 1154
rect 2832 1063 2844 1220
rect 2856 1063 2868 1132
rect 2880 1063 2892 1154
rect 2976 1063 2988 1220
rect 3000 1063 3012 1132
rect 3120 1063 3132 1220
rect 3264 1063 3276 1220
rect 3312 1063 3324 1154
rect 3408 1063 3420 1198
rect 3456 1063 3468 1154
rect 3552 1063 3564 1198
rect 3696 1063 3708 1198
rect 3720 1063 3732 1132
rect 3744 1063 3756 1154
rect 3840 1063 3852 1066
rect 3864 1063 3876 1088
rect 3912 1063 3924 1176
rect 3960 1063 3972 1066
rect 3984 1063 3996 1088
rect 4008 1063 4020 1110
rect 4032 1063 4044 1176
rect 4080 1063 4092 1066
rect 4128 1063 4140 1110
rect 4152 1063 4164 1198
rect 4200 1063 4212 1066
rect 4272 1063 4284 1220
rect 4320 1063 4332 1176
rect 4344 1063 4356 1132
rect 4440 1063 4452 1176
rect 4464 1063 4476 1132
rect 4488 1063 4500 1155
rect 4584 1063 4596 1198
rect 4608 1063 4620 1132
rect 4728 1063 4740 1088
rect 4752 1063 4764 1132
rect 4776 1063 4788 1153
rect 4824 1063 4836 1132
rect 4968 1063 4980 1176
rect 5016 1063 5028 1176
rect 5040 1063 5052 1132
rect 5088 1063 5100 1132
rect 5136 1063 5148 1132
rect 5400 1063 5412 1066
rect 5424 1063 5436 1088
rect 5448 1063 5460 1110
rect 5472 1063 5484 1154
rect 5496 1063 5508 1132
rect 5544 1063 5556 1066
rect 5568 1063 5580 1088
rect 5592 1063 5604 1110
rect 5640 1063 5652 1176
rect 5688 1063 5700 1176
rect 5712 1063 5724 1132
rect 5736 1063 5748 1132
rect 5808 1063 5820 1088
rect 5880 1063 5892 1176
rect 5928 1063 5940 1176
rect 6000 1063 6012 1199
rect 6048 1063 6060 1132
rect 6072 1063 6084 1239
rect 6096 1063 6108 1176
rect 6144 1063 6156 1176
rect 6168 1063 6180 1199
rect 6240 1063 6252 1132
rect 6264 1063 6276 1239
rect 6360 1063 6372 1132
rect 6384 1063 6396 1239
rect 6480 1063 6492 1132
rect 6504 1063 6516 1239
rect 6600 1063 6612 1066
rect 6624 1063 6636 1088
rect 6696 1063 6708 1176
rect 6744 1063 6756 1066
rect 6768 1063 6780 1110
rect 6816 1063 6828 1132
rect 6864 1063 6876 1066
rect 6888 1063 6900 1088
rect 6912 1063 6924 1110
rect 6936 1063 6948 1154
rect 6960 1063 6972 1066
rect 7008 1063 7020 1066
rect 7032 1063 7044 1132
rect 7056 1063 7068 1176
rect 72 261 84 264
rect 192 239 204 264
rect 312 217 324 264
rect 432 195 444 264
rect 552 173 564 264
rect 72 0 84 5
rect 336 0 348 137
rect 648 129 660 264
rect 768 151 780 264
rect 864 107 876 264
rect 504 0 516 93
rect 672 0 684 49
rect 696 0 708 71
rect 936 63 948 264
rect 1128 151 1140 264
rect 768 0 780 27
rect 984 0 996 93
rect 1152 85 1164 264
rect 1128 0 1140 49
rect 1320 41 1332 264
rect 1368 107 1380 264
rect 1536 173 1548 264
rect 1464 0 1476 93
rect 1656 63 1668 264
rect 1728 217 1740 264
rect 1752 173 1764 264
rect 1824 261 1836 264
rect 1944 217 1956 264
rect 2136 217 2148 264
rect 2328 261 2340 264
rect 2496 151 2508 264
rect 2592 217 2604 264
rect 2640 129 2652 264
rect 2712 195 2724 264
rect 1824 0 1836 71
rect 2232 0 2244 49
rect 2568 0 2580 27
rect 2784 19 2796 264
rect 2928 107 2940 264
rect 3024 172 3036 264
rect 3072 86 3084 264
rect 3144 195 3156 264
rect 3168 173 3180 264
rect 3216 148 3228 264
rect 3288 195 3300 264
rect 3184 63 3196 135
rect 3264 124 3276 137
rect 3360 129 3372 264
rect 3432 195 3444 264
rect 2880 0 2892 5
rect 3216 0 3228 110
rect 3308 41 3320 115
rect 3384 105 3396 115
rect 3336 0 3348 91
rect 3432 81 3444 93
rect 3384 0 3396 67
rect 3504 19 3516 264
rect 3576 195 3588 264
rect 3600 173 3612 264
rect 3648 151 3660 264
rect 3792 107 3804 264
rect 3888 217 3900 264
rect 4104 239 4116 264
rect 4224 239 4236 264
rect 4248 217 4260 264
rect 4392 85 4404 264
rect 4536 151 4548 264
rect 4632 173 4644 264
rect 4680 107 4692 264
rect 4872 239 4884 264
rect 4896 195 4908 264
rect 4920 173 4932 264
rect 5160 261 5172 264
rect 5184 218 5196 264
rect 5209 129 5221 225
rect 5232 63 5244 264
rect 5280 239 5292 264
rect 5304 151 5316 264
rect 5352 239 5364 264
rect 5616 195 5628 264
rect 5784 261 5796 264
rect 3552 0 3564 49
rect 5352 0 5364 115
rect 5377 0 5389 71
rect 5664 19 5676 225
rect 5832 217 5844 264
rect 5952 195 5964 264
rect 5976 173 5988 264
rect 6192 129 6204 264
rect 6312 85 6324 264
rect 6432 81 6444 264
rect 6552 151 6564 264
rect 6648 195 6660 264
rect 6672 217 6684 264
rect 6792 195 6804 264
rect 7080 256 7092 264
rect 7080 244 7188 256
rect 5424 0 5436 5
rect 5472 0 5484 5
rect 5520 0 5532 5
rect 5568 0 5580 5
rect 5616 0 5628 5
rect 5664 0 5676 5
rect 5712 0 5724 5
rect 5760 0 5772 5
rect 6000 0 6012 71
rect 6072 0 6084 5
rect 6120 0 6132 5
rect 6168 0 6180 5
rect 6216 0 6228 5
rect 6456 0 6468 67
rect 6528 0 6540 5
rect 6576 0 6588 5
rect 6816 0 6828 137
rect 6888 0 6900 5
rect 7176 0 7188 244
rect 7344 0 7356 93
use inv inv_0
timestamp 1386238110
transform 1 0 0 0 1 264
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 120 0 1 264
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 240 0 1 264
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 360 0 1 264
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 480 0 1 264
box 0 0 120 799
use and2 and2_4
timestamp 1386234845
transform 1 0 600 0 1 264
box 0 0 120 799
use xor2 xor2_3
timestamp 1396952988
transform 1 0 720 0 1 264
box 0 0 192 799
use xor2 xor2_4
timestamp 1396952988
transform 1 0 912 0 1 264
box 0 0 192 799
use xor2 xor2_5
timestamp 1396952988
transform 1 0 1104 0 1 264
box 0 0 192 799
use rowcrosser rowcrosser_1
timestamp 1397224710
transform 1 0 1296 0 1 264
box 0 0 48 799
use inv inv_6
timestamp 1386238110
transform 1 0 1344 0 1 264
box 0 0 120 799
use nand3 nand3_3
timestamp 1396952988
transform 1 0 1464 0 1 264
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 1584 0 1 264
box 0 0 96 799
use nand3 nand3_0
timestamp 1396952988
transform 1 0 1680 0 1 264
box 0 0 120 799
use nand3 nand3_1
timestamp 1396952988
transform 1 0 1800 0 1 264
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 1920 0 1 264
box 0 0 96 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 2016 0 1 264
box 0 0 96 799
use nand2 nand2_16
timestamp 1386234792
transform 1 0 2112 0 1 264
box 0 0 96 799
use nand2 nand2_17
timestamp 1386234792
transform 1 0 2208 0 1 264
box 0 0 96 799
use nand3 nand3_2
timestamp 1396952988
transform 1 0 2304 0 1 264
box 0 0 120 799
use nand2 nand2_18
timestamp 1386234792
transform 1 0 2424 0 1 264
box 0 0 96 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 2520 0 1 264
box 0 0 144 799
use nor3 nor3_6
timestamp 1386235396
transform 1 0 2664 0 1 264
box 0 0 144 799
use nor3 nor3_7
timestamp 1386235396
transform 1 0 2808 0 1 264
box 0 0 144 799
use nor3 nor3_8
timestamp 1386235396
transform 1 0 2952 0 1 264
box 0 0 144 799
use nor3 nor3_9
timestamp 1386235396
transform 1 0 3096 0 1 264
box 0 0 144 799
use nor3 nor3_10
timestamp 1386235396
transform 1 0 3240 0 1 264
box 0 0 144 799
use nor3 nor3_11
timestamp 1386235396
transform 1 0 3384 0 1 264
box 0 0 144 799
use nor3 nor3_12
timestamp 1386235396
transform 1 0 3528 0 1 264
box 0 0 144 799
use nor3 nor3_13
timestamp 1386235396
transform 1 0 3672 0 1 264
box 0 0 144 799
use nand3 nand3_4
timestamp 1396952988
transform 1 0 3816 0 1 264
box 0 0 120 799
use nand3 nand3_5
timestamp 1396952988
transform 1 0 3936 0 1 264
box 0 0 120 799
use nand3 nand3_6
timestamp 1396952988
transform 1 0 4056 0 1 264
box 0 0 120 799
use nand3 nand3_7
timestamp 1396952988
transform 1 0 4176 0 1 264
box 0 0 120 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 4296 0 1 264
box 0 0 120 799
use nor3 nor3_15
timestamp 1386235396
transform 1 0 4416 0 1 264
box 0 0 144 799
use nor3 nor3_16
timestamp 1386235396
transform 1 0 4560 0 1 264
box 0 0 144 799
use nor3 nor3_2
timestamp 1386235396
transform 1 0 4704 0 1 264
box 0 0 144 799
use nor3 nor3_3
timestamp 1386235396
transform 1 0 4848 0 1 264
box 0 0 144 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 4992 0 1 264
box 0 0 120 799
use nor3 nor3_4
timestamp 1386235396
transform 1 0 5112 0 1 264
box 0 0 144 799
use and2 and2_3
timestamp 1386234845
transform 1 0 5256 0 1 264
box 0 0 120 799
use nand4 nand4_2
timestamp 1386234936
transform 1 0 5376 0 1 264
box 0 0 144 799
use nand4 nand4_3
timestamp 1386234936
transform 1 0 5520 0 1 264
box 0 0 144 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 5664 0 1 264
box 0 0 96 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 5760 0 1 264
box 0 0 144 799
use nand3 nand3_9
timestamp 1396952988
transform 1 0 5904 0 1 264
box 0 0 120 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 6024 0 1 264
box 0 0 96 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 6120 0 1 264
box 0 0 96 799
use and2 and2_0
timestamp 1386234845
transform 1 0 6216 0 1 264
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 6336 0 1 264
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 6456 0 1 264
box 0 0 120 799
use nand4 nand4_4
timestamp 1386234936
transform 1 0 6576 0 1 264
box 0 0 144 799
use nand3 nand3_10
timestamp 1396952988
transform 1 0 6720 0 1 264
box 0 0 120 799
use nand4 nand4_5
timestamp 1386234936
transform 1 0 6840 0 1 264
box 0 0 144 799
use nand3 nand3_11
timestamp 1396952988
transform 1 0 6984 0 1 264
box 0 0 120 799
<< labels >>
rlabel metal2 6264 1239 6276 1239 5 imm4[2]
rlabel metal2 6384 1239 6396 1239 5 imm4[1]
rlabel metal2 6504 1239 6516 1239 5 imm4[0]
rlabel metal2 6072 1239 6084 1239 5 imm4[3]
rlabel metal2 1248 1239 1260 1239 5 C
rlabel metal2 1056 1239 1068 1239 5 V
rlabel metal2 1320 1239 1332 1239 5 N
rlabel metal2 1416 1239 1428 1239 5 Z
rlabel m2contact 3917 1183 3917 1183 1 ABnC
rlabel m2contact 4277 1225 4277 1225 1 AnBnC
rlabel m2contact 4156 1203 4156 1203 1 AnBC
rlabel m2contact 4037 1180 4037 1180 1 ABC
rlabel metal1 5250 143 5250 143 1 ShSign
rlabel metal1 336 211 336 211 1 nC
rlabel metal1 104 253 104 253 1 nA
rlabel metal1 210 231 210 231 1 nB
rlabel metal1 459 186 459 186 1 nD
rlabel metal1 579 164 579 164 1 nE
rlabel metal1 668 123 668 123 1 UseC
rlabel metal2 72 0 84 0 1 ZeroA
rlabel metal2 336 0 348 0 1 SUB
rlabel metal2 504 0 516 0 1 CIn_slice
rlabel metal2 672 0 684 0 1 LastCIn
rlabel metal2 696 0 708 0 1 COut
rlabel metal2 984 0 996 0 1 nZ
rlabel metal2 768 0 780 0 1 N
rlabel metal2 1128 0 1140 0 1 FAOut
rlabel metal2 1464 0 1476 0 1 AND
rlabel metal2 1824 0 1836 0 1 OR
rlabel metal2 2232 0 2244 0 1 XOR
rlabel metal2 2568 0 2580 0 1 NOT
rlabel metal2 2880 0 2892 0 1 NAND
rlabel metal2 3216 0 3228 0 1 NOR
rlabel metal2 3336 0 3348 0 1 ASign
rlabel metal2 3384 0 3396 0 1 ShB
rlabel metal2 3552 0 3564 0 1 ShL
rlabel metal2 5352 0 5364 0 1 Sh8
rlabel metal2 5377 0 5389 0 1 ShR
rlabel metal2 6000 0 6012 0 1 Sh4
rlabel metal2 6456 0 6468 0 1 Sh2
rlabel metal2 6816 0 6828 0 1 Sh1
rlabel metal2 7176 0 7188 0 1 ShOut
rlabel metal2 7344 0 7356 0 1 LLI
rlabel metal1 7656 317 7656 327 7 Clock
rlabel metal1 7656 1046 7656 1056 1 ScanReturn
rlabel metal1 7656 1023 7656 1033 1 Scan
rlabel metal1 7656 340 7656 365 7 GND!
rlabel metal1 7656 985 7656 1010 7 Vdd!
rlabel metal1 0 1068 0 1078 3 OpCode[4]
rlabel metal1 0 1090 0 1100 3 OpCode[3]
rlabel metal1 0 1112 0 1122 3 OpCode[2]
rlabel metal1 0 1134 0 1144 3 OpCode[1]
rlabel metal1 0 1156 0 1166 3 OpCode[0]
rlabel metal1 0 1178 0 1188 3 Cin
rlabel metal2 6072 0 6084 0 1 ShiftIn
rlabel metal2 6120 0 6132 0 1 ShiftIn
rlabel metal2 6168 0 6180 0 1 ShiftIn
rlabel metal2 6216 0 6228 0 1 ShiftIn
rlabel metal2 6528 0 6540 0 1 ShiftIn
rlabel metal2 6576 0 6588 0 1 ShiftIn
rlabel metal2 6888 0 6900 0 1 ShiftIn
rlabel metal1 7656 294 7656 304 7 Test
rlabel metal1 7656 271 7656 281 7 nReset
rlabel metal2 5424 0 5436 0 1 ShiftIn
rlabel metal2 5472 0 5484 0 1 ShiftIn
rlabel metal2 5520 0 5532 0 1 ShiftIn
rlabel metal2 5568 0 5580 0 1 ShiftIn
rlabel metal2 5616 0 5628 0 1 ShiftIn
rlabel metal2 5664 0 5676 0 1 ShiftIn
rlabel metal2 5712 0 5724 0 1 ShiftIn
rlabel metal2 5760 0 5772 0 1 ShiftIn
<< end >>
