magic
tech c035u
timestamp 1397224710
<< metal1 >>
rect 14 19475 14361 19485
rect 37 19451 14554 19461
rect 60 19427 14746 19437
rect 14938 19425 14972 19435
rect 83 19403 14938 19413
rect 14962 19401 14972 19425
rect 15130 19402 15164 19412
rect 106 19379 15130 19389
rect 15154 19377 15164 19402
rect 129 19355 3945 19365
rect 152 19331 4377 19341
rect 175 19307 4761 19317
rect 198 19283 3993 19293
rect 221 19259 4425 19269
rect 244 19235 4809 19245
rect 267 19211 6949 19221
rect 22138 19209 22171 19219
rect 290 19187 6925 19197
rect 6939 19187 22137 19197
rect 22161 19185 22171 19209
rect 313 19163 6901 19173
rect 6915 19163 22329 19173
rect 336 19139 22449 19149
rect 22569 19137 22603 19147
rect 359 19115 22569 19125
rect 22593 19113 22603 19137
rect 2879 17675 2890 17685
rect 14 16788 365 16798
rect 25391 16787 25408 16797
rect 2842 16721 2890 16731
rect 25391 16721 25408 16731
rect 2842 16699 2890 16709
rect 2879 16564 2890 16574
rect 37 15677 365 15687
rect 25391 15676 25408 15686
rect 2842 15610 2890 15620
rect 25391 15610 25408 15620
rect 2842 15588 2890 15598
rect 2879 15453 2890 15463
rect 60 14566 365 14576
rect 25391 14565 25408 14575
rect 2842 14499 2890 14509
rect 25391 14499 25408 14509
rect 2842 14477 2890 14487
rect 2879 14342 2890 14352
rect 83 13455 365 13465
rect 25391 13454 25408 13464
rect 2842 13388 2890 13398
rect 25391 13388 25408 13398
rect 2842 13366 2890 13376
rect 2879 13231 2890 13241
rect 106 12344 365 12354
rect 25391 12343 25408 12353
rect 2842 12277 2890 12287
rect 25391 12277 25408 12287
rect 2842 12255 2890 12265
rect 2879 12120 2890 12130
rect 95 11255 131 11265
rect 95 11231 105 11255
rect 129 11233 365 11243
rect 25391 11232 25408 11242
rect 2842 11166 2890 11176
rect 25391 11166 25408 11176
rect 2842 11144 2890 11154
rect 2879 11009 2890 11019
rect 118 10144 152 10154
rect 118 10120 128 10144
rect 152 10122 365 10132
rect 25391 10121 25408 10131
rect 2842 10055 2890 10065
rect 25391 10055 25408 10065
rect 2842 10033 2890 10043
rect 2879 9898 2890 9908
rect 141 9033 175 9043
rect 141 9009 151 9033
rect 175 9011 365 9021
rect 25391 9010 25408 9020
rect 2842 8944 2890 8954
rect 25391 8944 25408 8954
rect 2842 8922 2890 8932
rect 2879 8787 2890 8797
rect 164 7922 198 7932
rect 164 7898 174 7922
rect 198 7900 365 7910
rect 25391 7899 25408 7909
rect 2842 7833 2890 7843
rect 25391 7833 25408 7843
rect 2842 7811 2890 7821
rect 2879 7676 2890 7686
rect 187 6811 221 6821
rect 187 6787 197 6811
rect 221 6789 365 6799
rect 25391 6788 25408 6798
rect 2842 6722 2890 6732
rect 25391 6722 25408 6732
rect 2842 6700 2890 6710
rect 2879 6565 2890 6575
rect 210 5700 244 5710
rect 210 5676 220 5700
rect 244 5678 365 5688
rect 25391 5677 25408 5687
rect 2842 5611 2890 5621
rect 25391 5611 25408 5621
rect 2842 5589 2890 5599
rect 2879 5454 2890 5464
rect 233 4589 267 4599
rect 233 4565 243 4589
rect 267 4567 365 4577
rect 25391 4566 25408 4576
rect 2842 4500 2890 4510
rect 25391 4500 25408 4510
rect 2842 4478 2890 4488
rect 2879 4343 2890 4353
rect 256 3478 290 3488
rect 256 3454 266 3478
rect 290 3456 365 3466
rect 25391 3455 25408 3465
rect 2842 3389 2890 3399
rect 25391 3389 25408 3399
rect 2842 3367 2890 3377
rect 2879 3232 2890 3242
rect 279 2367 313 2377
rect 279 2343 289 2367
rect 313 2345 365 2355
rect 25391 2344 25408 2354
rect 2842 2278 2890 2288
rect 25391 2278 25408 2288
rect 2842 2256 2890 2266
rect 2879 2121 2890 2131
rect 302 1256 335 1266
rect 302 1232 312 1256
rect 336 1234 365 1244
rect 25391 1233 25408 1243
rect 2842 1167 2890 1177
rect 25391 1167 25408 1177
rect 2842 1145 2890 1155
rect 2879 1010 2890 1020
rect 325 145 359 155
rect 325 121 335 145
rect 359 123 365 133
rect 25391 122 25408 132
rect 2842 56 2890 66
rect 25391 56 25408 66
rect 2842 34 2890 44
rect 570 8 3105 18
rect 17063 7 19713 17
rect 19727 7 19760 17
rect 19774 7 19809 17
rect 19823 7 19857 17
rect 19871 7 19905 17
rect 19919 7 19953 17
rect 19967 7 20001 17
rect 20015 7 20049 17
rect 20063 7 20361 17
rect 20375 7 20409 17
rect 20423 7 20456 17
rect 20470 7 20505 17
rect 20519 7 20817 17
rect 20831 7 20865 17
rect 20879 7 21249 17
rect 21263 7 25186 17
<< m2contact >>
rect 0 19473 14 19487
rect 14361 19474 14375 19488
rect 23 19449 37 19463
rect 14554 19449 14568 19463
rect 46 19425 60 19439
rect 14746 19425 14760 19439
rect 69 19401 83 19415
rect 14938 19401 14952 19415
rect 92 19377 106 19391
rect 15130 19377 15144 19392
rect 115 19353 129 19367
rect 3945 19353 3959 19367
rect 138 19329 152 19343
rect 4377 19329 4391 19343
rect 161 19305 175 19319
rect 4761 19305 4775 19319
rect 184 19281 198 19295
rect 3993 19281 4007 19295
rect 207 19257 221 19271
rect 4425 19257 4439 19271
rect 230 19233 244 19247
rect 4809 19233 4823 19247
rect 253 19209 267 19223
rect 6949 19209 6963 19223
rect 276 19185 290 19199
rect 6925 19185 6939 19199
rect 22137 19185 22151 19199
rect 299 19161 313 19175
rect 6901 19161 6915 19175
rect 22329 19160 22343 19174
rect 322 19137 336 19151
rect 22449 19137 22463 19151
rect 345 19113 359 19127
rect 22569 19113 22583 19127
rect 2865 17673 2879 17687
rect 0 16786 14 16800
rect 2865 16562 2879 16576
rect 23 15675 37 15689
rect 2865 15451 2879 15465
rect 46 14564 60 14578
rect 2865 14340 2879 14354
rect 69 13453 83 13467
rect 2865 13229 2879 13243
rect 92 12342 106 12356
rect 2865 12118 2879 12132
rect 115 11231 129 11245
rect 2865 11007 2879 11021
rect 138 10120 152 10134
rect 2865 9896 2879 9910
rect 161 9009 175 9023
rect 2865 8785 2879 8799
rect 184 7898 198 7912
rect 2865 7674 2879 7688
rect 207 6787 221 6801
rect 2865 6563 2879 6577
rect 230 5676 244 5690
rect 2865 5452 2879 5466
rect 253 4565 267 4579
rect 2865 4341 2879 4355
rect 276 3454 290 3468
rect 2865 3230 2879 3244
rect 299 2343 313 2357
rect 2865 2119 2879 2133
rect 322 1232 336 1246
rect 2865 1008 2879 1022
rect 345 121 359 135
rect 556 6 570 20
rect 3105 5 3119 19
rect 17049 5 17063 19
rect 19713 5 19727 19
rect 19760 5 19774 19
rect 19809 5 19823 19
rect 19857 5 19871 19
rect 19905 5 19919 19
rect 19953 5 19967 19
rect 20001 5 20015 19
rect 20049 5 20063 19
rect 20361 5 20375 19
rect 20409 5 20423 19
rect 20456 5 20470 19
rect 20505 5 20519 19
rect 20817 5 20831 19
rect 20865 5 20879 19
rect 21249 5 21263 19
rect 25186 5 25200 19
<< metal2 >>
rect 1 16800 13 19473
rect 1 0 13 16786
rect 24 15689 36 19449
rect 24 0 36 15675
rect 47 14578 59 19425
rect 47 0 59 14564
rect 70 13467 82 19401
rect 70 0 82 13453
rect 93 12356 105 19377
rect 93 0 105 12342
rect 116 11245 128 19353
rect 116 0 128 11231
rect 139 10134 151 19329
rect 139 0 151 10120
rect 162 9023 174 19305
rect 162 0 174 9009
rect 185 7912 197 19281
rect 185 0 197 7898
rect 208 6801 220 19257
rect 208 0 220 6787
rect 231 5690 243 19233
rect 231 0 243 5676
rect 254 4579 266 19209
rect 254 0 266 4565
rect 277 3468 289 19185
rect 277 0 289 3454
rect 300 2357 312 19161
rect 300 0 312 2343
rect 323 1246 335 19137
rect 323 0 335 1232
rect 346 135 358 19113
rect 370 19105 570 19490
rect 586 19105 598 19490
rect 610 19105 622 19490
rect 634 19105 646 19490
rect 658 19105 670 19490
rect 3922 19105 3934 19490
rect 3946 19105 3958 19353
rect 3994 19105 4006 19281
rect 4162 19105 4174 19490
rect 4378 19105 4390 19329
rect 4426 19105 4438 19257
rect 4762 19105 4774 19305
rect 4810 19105 4822 19233
rect 5122 19105 5134 19490
rect 5314 19105 5326 19490
rect 6348 19105 6360 19490
rect 6902 19105 6914 19161
rect 6926 19105 6938 19185
rect 6950 19105 6962 19209
rect 14339 19105 14351 19490
rect 14363 19105 14375 19474
rect 14555 19105 14567 19449
rect 14603 19105 14615 19490
rect 14747 19105 14759 19425
rect 14939 19105 14951 19401
rect 15131 19105 15143 19377
rect 15323 19105 15335 19490
rect 17122 19105 17134 19490
rect 17314 19105 17326 19490
rect 17386 19105 17398 19490
rect 17482 19105 17494 19490
rect 22138 19105 22150 19185
rect 22330 19105 22342 19160
rect 22450 19105 22462 19137
rect 22570 19105 22582 19113
rect 25186 19105 25386 19490
rect 2866 17603 2878 17673
rect 2866 16492 2878 16562
rect 2866 15381 2878 15451
rect 2866 14270 2878 14340
rect 2866 13159 2878 13229
rect 2866 12048 2878 12118
rect 2866 10937 2878 11007
rect 2866 9826 2878 9896
rect 2866 8715 2878 8785
rect 2866 7604 2878 7674
rect 2866 6493 2878 6563
rect 2866 5382 2878 5452
rect 2866 4271 2878 4341
rect 2866 3160 2878 3230
rect 2866 2049 2878 2119
rect 2866 938 2878 1008
rect 346 0 358 121
rect 370 20 570 27
rect 370 6 556 20
rect 370 0 570 6
rect 586 0 598 27
rect 610 0 622 27
rect 634 0 646 27
rect 658 0 670 27
rect 1906 0 1918 27
rect 2698 0 2710 27
rect 3106 19 3118 27
rect 3250 0 3262 27
rect 3466 0 3478 27
rect 4210 0 4222 27
rect 4378 0 4390 27
rect 4762 0 4774 27
rect 4954 0 4966 27
rect 5170 0 5182 27
rect 5914 0 5926 27
rect 6082 0 6094 27
rect 15490 0 15502 27
rect 15682 0 15694 27
rect 15922 0 15934 27
rect 16570 21 16582 27
rect 16762 21 16774 27
rect 16570 9 16774 21
rect 17050 19 17062 27
rect 19714 19 19726 27
rect 19762 19 19774 27
rect 19810 19 19822 27
rect 19858 19 19870 27
rect 19906 19 19918 27
rect 19954 19 19966 27
rect 20002 19 20014 27
rect 20050 19 20062 27
rect 20362 19 20374 27
rect 20410 19 20422 27
rect 20458 19 20470 27
rect 20506 19 20518 27
rect 20818 19 20830 27
rect 20866 19 20878 27
rect 21250 19 21262 27
rect 23626 0 23638 27
rect 24370 0 24382 27
rect 24586 0 24598 27
rect 24730 0 24742 27
rect 24778 0 24790 27
rect 24826 0 24838 27
rect 24874 0 24886 27
rect 24946 0 24958 27
rect 25186 19 25386 27
rect 25200 5 25386 19
rect 25186 0 25386 5
use slice17 slice17_0
timestamp 1397224710
transform 1 0 370 0 1 17803
box 0 0 25016 1302
use leftbuf_slice leftbuf_slice_0
array 0 0 1469 0 15 1111
timestamp 1396389552
transform 1 0 365 0 1 27
box 0 0 1469 1111
use IrAA IrAA_0
array 0 0 1008 0 7 1111
timestamp 1397224710
transform 1 0 1834 0 1 8915
box 0 0 1008 1111
use tielow tielow_0
timestamp 1386086605
transform 1 0 2842 0 1 16804
box 0 0 48 799
use tielow tielow_1
timestamp 1386086605
transform 1 0 2842 0 1 15693
box 0 0 48 799
use tielow tielow_2
timestamp 1386086605
transform 1 0 2842 0 1 14582
box 0 0 48 799
use tielow tielow_3
timestamp 1386086605
transform 1 0 2842 0 1 13471
box 0 0 48 799
use tielow tielow_4
timestamp 1386086605
transform 1 0 2842 0 1 12360
box 0 0 48 799
use tielow tielow_5
timestamp 1386086605
transform 1 0 2842 0 1 11249
box 0 0 48 799
use tielow tielow_6
timestamp 1386086605
transform 1 0 2842 0 1 10138
box 0 0 48 799
use tielow tielow_7
timestamp 1386086605
transform 1 0 2842 0 1 9027
box 0 0 48 799
use IrBA IrBA_0
array 0 0 1008 0 2 1111
timestamp 1397224710
transform 1 0 1834 0 1 5582
box 0 0 1008 1111
use tielow tielow_8
timestamp 1386086605
transform 1 0 2842 0 1 7916
box 0 0 48 799
use tielow tielow_9
timestamp 1386086605
transform 1 0 2842 0 1 6805
box 0 0 48 799
use tielow tielow_10
timestamp 1386086605
transform 1 0 2842 0 1 5694
box 0 0 48 799
use IrBB IrBB_0
array 0 0 1008 0 4 1111
timestamp 1397224710
transform 1 0 1834 0 1 27
box 0 0 1008 1111
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 2842 0 1 4583
box 0 0 48 799
use tielow tielow_12
timestamp 1386086605
transform 1 0 2842 0 1 3472
box 0 0 48 799
use tielow tielow_13
timestamp 1386086605
transform 1 0 2842 0 1 2361
box 0 0 48 799
use tielow tielow_14
timestamp 1386086605
transform 1 0 2842 0 1 1250
box 0 0 48 799
use tielow tielow_15
timestamp 1386086605
transform 1 0 2842 0 1 139
box 0 0 48 799
use Datapath_slice Datapath_slice_0
array 0 0 20472 0 15 1111
timestamp 1397224710
transform 1 0 2890 0 1 27
box 0 0 20472 1111
use LLIcell_U LLIcell_U_0
array 0 0 192 0 7 1111
timestamp 1396390011
transform 1 0 23362 0 1 8915
box 0 0 192 1111
use LLIcell_L LLIcell_L_0
array 0 0 192 0 7 1111
timestamp 1396390031
transform 1 0 23362 0 1 27
box 0 0 192 1111
use Datapath_end_high Datapath_end_high_0
array 0 0 1837 0 11 1111
timestamp 1397220089
transform 1 0 23554 0 1 4471
box 0 0 1837 1111
use Datapath_end_low Datapath_end_low_0
array 0 0 1837 0 3 1111
timestamp 1397224710
transform 1 0 23554 0 1 27
box 0 0 1837 1111
<< labels >>
rlabel metal2 1 0 13 0 1 Ir[15]
rlabel metal2 24 0 36 0 1 Ir[14]
rlabel metal2 47 0 59 0 1 Ir[13]
rlabel metal2 70 0 82 0 1 Ir[12]
rlabel metal2 93 0 105 0 1 Ir[11]
rlabel metal2 116 0 128 0 1 Ir[10]
rlabel metal2 139 0 151 0 1 Ir[9]
rlabel metal2 162 0 174 0 1 Ir[8]
rlabel metal2 185 0 197 0 1 Ir[7]
rlabel metal2 208 0 220 0 1 Ir[6]
rlabel metal2 231 0 243 0 1 Ir[5]
rlabel metal2 254 0 266 0 1 Ir[4]
rlabel metal2 277 0 289 0 1 Ir[3]
rlabel metal2 300 0 312 0 1 Ir[2]
rlabel metal2 323 0 335 0 1 Ir[1]
rlabel metal2 346 0 358 0 1 Ir[0]
rlabel metal2 658 0 670 0 1 nReset
rlabel metal2 634 0 646 0 1 Clock
rlabel metal2 610 0 622 0 1 Test
rlabel metal2 586 0 598 0 1 SDI
rlabel metal2 370 0 570 0 1 Vdd!
rlabel metal2 24586 0 24598 0 1 MemEn
rlabel metal2 24946 0 24958 0 1 StatusRegEn
rlabel metal2 24730 0 24742 0 1 StatusReg[3]
rlabel metal2 24778 0 24790 0 1 StatusReg[2]
rlabel metal2 24826 0 24838 0 1 StatusReg[1]
rlabel metal2 24874 0 24886 0 1 StatusReg[0]
rlabel metal2 25186 0 25386 0 1 GND!
rlabel metal2 4210 0 4222 0 1 LrEn
rlabel metal2 4378 0 4390 0 1 PcSel[0]
rlabel metal2 4762 0 4774 0 1 PcSel[1]
rlabel metal2 23626 0 23638 0 1 AluWe
rlabel metal2 24370 0 24382 0 1 AluEn
rlabel metal2 5170 0 5182 0 1 PcWe
rlabel metal2 4954 0 4966 0 1 PcSel[2]
rlabel metal2 5914 0 5926 0 1 PcEn
rlabel metal2 6082 0 6094 0 1 WdSel
rlabel metal2 15490 0 15502 0 1 Op1Sel
rlabel metal2 15682 0 15694 0 1 Op2Sel[0]
rlabel metal2 15922 0 15934 0 1 Op2Sel[1]
rlabel metal2 1906 0 1918 0 1 IrWe
rlabel metal2 2698 0 2710 0 1 ImmSel
rlabel metal2 3466 0 3478 0 1 LrWe
rlabel metal2 3250 0 3262 0 1 LrSel
rlabel metal1 25408 56 25408 66 7 DataOut[0]
rlabel metal1 25408 1167 25408 1177 7 DataOut[1]
rlabel metal1 25408 2278 25408 2288 7 DataOut[2]
rlabel metal1 25408 3389 25408 3399 7 DataOut[3]
rlabel metal1 25408 4500 25408 4510 7 DataOut[4]
rlabel metal1 25408 5611 25408 5621 7 DataOut[5]
rlabel metal1 25408 6722 25408 6732 7 DataOut[6]
rlabel metal1 25408 7833 25408 7843 7 DataOut[7]
rlabel metal1 25408 8944 25408 8954 7 DataOut[8]
rlabel metal1 25408 10055 25408 10065 7 DataOut[9]
rlabel metal1 25408 11166 25408 11176 7 DataOut[10]
rlabel metal1 25408 12277 25408 12287 7 DataOut[11]
rlabel metal1 25408 13388 25408 13398 7 DataOut[12]
rlabel metal1 25408 14499 25408 14509 7 DataOut[13]
rlabel metal1 25408 15610 25408 15620 7 DataOut[14]
rlabel metal1 25408 16721 25408 16731 7 DataOut[15]
rlabel metal2 6 19178 6 19178 1 Ir[15]
rlabel metal2 30 19177 30 19177 1 Ir[14]
rlabel metal2 53 19177 53 19177 1 Ir[13]
rlabel metal2 76 19178 76 19178 1 Ir[12]
rlabel metal2 99 19178 99 19178 1 Ir[11]
rlabel metal2 122 19177 122 19177 1 Ir[10]
rlabel metal2 145 19178 145 19178 1 Ir[9]
rlabel metal2 168 19178 168 19178 1 Ir[8]
rlabel metal2 191 19180 191 19180 1 Ir[7]
rlabel metal2 214 19181 214 19181 1 Ir[6]
rlabel metal2 237 19182 237 19182 1 Ir[5]
rlabel metal2 260 19183 260 19183 1 Ir[4]
rlabel metal2 283 19182 283 19182 1 Ir[3]
rlabel metal2 586 19490 598 19490 5 SDO
rlabel metal2 370 19490 570 19490 5 Vdd!
rlabel metal2 658 19490 670 19490 1 nReset
rlabel metal2 634 19490 646 19490 1 Clock
rlabel metal2 610 19490 622 19490 1 Test
rlabel metal2 25186 19490 25386 19490 1 GND!
rlabel metal1 25408 122 25408 132 7 DataIn[0]
rlabel metal1 25408 1233 25408 1243 7 DataIn[1]
rlabel metal1 25408 2344 25408 2354 7 DataIn[2]
rlabel metal1 25408 3455 25408 3465 7 DataIn[3]
rlabel metal1 25408 4566 25408 4576 7 DataIn[4]
rlabel metal1 25408 5677 25408 5687 7 DataIn[5]
rlabel metal1 25408 6788 25408 6798 7 DataIn[6]
rlabel metal1 25408 7899 25408 7909 7 DataIn[7]
rlabel metal1 25408 9010 25408 9020 7 DataIn[8]
rlabel metal1 25408 10121 25408 10131 7 DataIn[9]
rlabel metal1 25408 11232 25408 11242 7 DataIn[10]
rlabel metal1 25408 12343 25408 12353 7 DataIn[11]
rlabel metal1 25408 13454 25408 13464 7 DataIn[12]
rlabel metal1 25408 14565 25408 14575 7 DataIn[13]
rlabel metal1 25408 15676 25408 15686 7 DataIn[14]
rlabel metal1 25408 16787 25408 16797 7 DataIn[15]
rlabel metal2 22144 19180 22144 19180 1 Ir[3]
rlabel metal2 22335 19155 22335 19155 1 Ir[2]
rlabel metal2 22455 19130 22455 19130 1 Ir[1]
rlabel metal2 22576 19108 22576 19108 1 Ir[0]
rlabel metal2 17482 19490 17494 19490 5 Flags[0]
rlabel metal2 17386 19490 17398 19490 5 Flags[3]
rlabel metal2 17314 19490 17326 19490 5 Flags[1]
rlabel metal2 17122 19490 17134 19490 5 Flags[2]
rlabel metal2 15323 19490 15335 19490 5 CFlag
rlabel metal2 14339 19490 14351 19490 5 AluOR[1]
rlabel metal2 14603 19490 14615 19490 5 AluOR[0]
rlabel metal2 14368 19467 14368 19467 1 Ir[15]
rlabel metal2 14559 19442 14559 19442 1 Ir[14]
rlabel metal2 15137 19370 15137 19370 1 Ir[11]
rlabel metal2 14945 19395 14945 19395 1 Ir[12]
rlabel metal2 14752 19419 14752 19419 1 Ir[13]
rlabel metal2 6906 19153 6906 19153 1 Ir[2]
rlabel metal2 6932 19177 6932 19177 1 Ir[3]
rlabel metal2 6955 19201 6955 19201 1 Ir[4]
rlabel metal2 6348 19490 6360 19490 5 RegWe
rlabel metal2 4000 19273 4000 19273 1 Ir[7]
rlabel metal2 3951 19346 3951 19346 1 Ir[10]
rlabel metal2 4432 19250 4432 19250 1 Ir[6]
rlabel metal2 4383 19321 4383 19321 1 Ir[9]
rlabel metal2 4767 19298 4767 19298 1 Ir[8]
rlabel metal2 4817 19227 4817 19227 1 Ir[5]
rlabel metal2 3922 19490 3934 19490 5 Rs1Sel[0]
rlabel metal2 4162 19490 4174 19490 5 Rs1Sel[1]
rlabel metal2 5122 19490 5134 19490 5 RwSel[0]
rlabel metal2 5314 19490 5326 19490 5 RwSel[1]
<< end >>
