magic
tech c035u
timestamp 1397223953
<< nwell >>
rect 264 506 508 904
rect 1396 506 2105 904
rect 3521 506 4156 904
rect 4948 506 5113 904
<< pwell >>
rect 264 105 508 506
rect 1396 105 2105 506
rect 3521 105 4156 506
rect 4948 105 5113 506
<< pohmic >>
rect 264 181 266 191
rect 504 181 508 191
rect 1396 181 1398 191
rect 2103 181 2105 191
rect 3521 181 3523 191
rect 4154 181 4156 191
rect 4948 181 4950 191
rect 5111 181 5113 191
<< nohmic >>
rect 264 841 265 851
rect 504 841 508 851
rect 1396 841 1398 851
rect 2103 841 2105 851
rect 3521 841 3523 851
rect 4154 841 4156 851
rect 4948 841 4950 851
rect 5111 841 5113 851
<< psubstratetap >>
rect 290 457 306 473
rect 347 457 363 473
rect 404 457 420 473
rect 461 457 477 473
rect 1430 457 1446 473
rect 1487 457 1503 473
rect 1544 457 1560 473
rect 1601 457 1617 473
rect 1658 457 1674 473
rect 1715 457 1731 473
rect 1772 457 1788 473
rect 1829 457 1845 473
rect 1886 457 1902 473
rect 1943 457 1959 473
rect 2000 457 2016 473
rect 2057 457 2073 473
rect 3539 457 3555 473
rect 3596 457 3612 473
rect 3653 457 3669 473
rect 3710 457 3726 473
rect 3767 457 3783 473
rect 3824 457 3840 473
rect 3881 457 3897 473
rect 3938 457 3954 473
rect 3995 457 4011 473
rect 4052 457 4068 473
rect 4109 457 4125 473
rect 4964 457 4980 473
rect 5021 457 5037 473
rect 5078 457 5094 473
rect 266 181 504 197
rect 1398 181 2103 197
rect 3523 181 4154 197
rect 4950 181 5111 197
<< nsubstratetap >>
rect 265 835 504 851
rect 1398 835 2103 851
rect 3523 835 4154 851
rect 4950 835 5111 851
<< metal1 >>
rect 135 1112 191 1124
rect 205 1112 1083 1124
rect 1097 1112 2632 1124
rect 2646 1112 3448 1124
rect 3462 1112 4875 1124
rect 4889 1112 5856 1124
rect 5870 1112 6624 1124
rect 6638 1112 7416 1124
rect 0 1090 71 1100
rect 85 1090 843 1100
rect 857 1090 2392 1100
rect 2406 1090 3328 1100
rect 3342 1090 4755 1100
rect 4769 1090 5640 1100
rect 5654 1090 6408 1100
rect 6422 1090 7296 1100
rect 0 1068 47 1078
rect 61 1068 819 1078
rect 833 1068 2512 1078
rect 2526 1068 3232 1078
rect 3246 1068 4635 1078
rect 4649 1068 5736 1078
rect 5750 1068 6384 1078
rect 6398 1068 7176 1078
rect 0 1045 23 1055
rect 37 1045 963 1055
rect 977 1045 2368 1055
rect 2382 1045 3208 1055
rect 3222 1045 4611 1055
rect 4625 1045 5616 1055
rect 5630 1045 6504 1055
rect 6518 1045 7152 1055
rect 8126 1046 8304 1056
rect 8318 1046 8496 1056
rect 8510 1046 8688 1056
rect 8702 1046 8880 1056
rect 8894 1046 9072 1056
rect 737 1022 2152 1032
rect 2166 1022 2992 1032
rect 3006 1022 4515 1032
rect 4529 1022 5520 1032
rect 5534 1022 6192 1032
rect 6206 1022 6960 1032
rect 6974 1022 7896 1032
rect 8054 1020 8568 1030
rect 8582 1020 8952 1030
rect 8966 1020 9144 1030
rect 9182 1019 9217 1029
rect 713 1000 2128 1010
rect 2142 1000 3112 1010
rect 3126 1000 4419 1010
rect 4433 1000 5400 1010
rect 5414 1000 6288 1010
rect 6302 1000 6936 1010
rect 6950 1000 7776 1010
rect 8990 997 9217 1007
rect 689 977 2272 987
rect 2286 977 2968 987
rect 2982 977 4395 987
rect 4409 977 5376 987
rect 5390 977 6168 987
rect 6182 977 7056 987
rect 7070 977 7752 987
rect 8006 976 8184 986
rect 8198 976 8760 986
rect 8798 975 9217 985
rect 0 954 579 964
rect 593 954 1203 964
rect 1217 954 2752 964
rect 2766 954 4299 964
rect 4313 954 5280 964
rect 5294 954 5976 964
rect 5990 954 6744 964
rect 6758 954 7656 964
rect 8606 953 9217 963
rect 0 932 555 942
rect 569 932 1179 942
rect 1193 932 2872 942
rect 2886 932 4203 942
rect 4217 932 5160 942
rect 5174 932 6072 942
rect 6086 932 6720 942
rect 6734 932 7536 942
rect 8414 931 9217 941
rect 0 909 531 919
rect 545 909 1323 919
rect 1337 909 2728 919
rect 2742 909 4179 919
rect 4193 909 5136 919
rect 5150 909 5952 919
rect 5966 909 6840 919
rect 6854 909 7512 919
rect 8222 909 9217 919
rect 264 887 508 897
rect 1396 887 2105 897
rect 3521 887 4156 897
rect 4948 887 5113 897
rect 264 864 508 874
rect 1396 864 2105 874
rect 3521 864 4156 874
rect 4948 864 5113 874
rect 264 835 265 851
rect 504 835 508 851
rect 264 826 508 835
rect 1396 835 1398 851
rect 2103 835 2105 851
rect 1396 826 2105 835
rect 3521 835 3523 851
rect 4154 835 4156 851
rect 3521 826 4156 835
rect 4948 835 4950 851
rect 5111 835 5113 851
rect 4948 826 5113 835
rect 290 206 306 457
rect 347 206 363 457
rect 404 206 420 457
rect 461 206 477 457
rect 1430 206 1446 457
rect 1487 206 1503 457
rect 1544 206 1560 457
rect 1601 206 1617 457
rect 1658 206 1674 457
rect 1715 206 1731 457
rect 1772 206 1788 457
rect 1829 206 1845 457
rect 1886 206 1902 457
rect 1943 206 1959 457
rect 2000 206 2016 457
rect 2057 206 2073 457
rect 3539 206 3555 457
rect 3596 206 3612 457
rect 3653 206 3669 457
rect 3710 206 3726 457
rect 3767 206 3783 457
rect 3824 206 3840 457
rect 3881 206 3897 457
rect 3938 206 3954 457
rect 3995 206 4011 457
rect 4052 206 4068 457
rect 4109 206 4125 457
rect 4964 206 4980 457
rect 5021 206 5037 457
rect 5078 206 5094 457
rect 264 197 508 206
rect 264 181 266 197
rect 504 181 508 197
rect 1396 197 2105 206
rect 1396 181 1398 197
rect 2103 181 2105 197
rect 3521 197 4156 206
rect 3521 181 3523 197
rect 4154 181 4156 197
rect 4948 197 5113 206
rect 4948 181 4950 197
rect 5111 181 5113 197
rect 264 158 508 168
rect 1396 158 2105 168
rect 3521 158 4156 168
rect 4948 158 5113 168
rect 264 135 508 145
rect 1396 135 2105 145
rect 3521 135 4156 145
rect 4948 135 5113 145
rect 264 112 508 122
rect 1396 112 2105 122
rect 3521 112 4156 122
rect 4948 112 5113 122
<< m2contact >>
rect 121 1112 135 1126
rect 191 1111 205 1125
rect 1083 1111 1097 1125
rect 2632 1111 2646 1125
rect 3448 1111 3462 1125
rect 4875 1111 4889 1125
rect 5856 1111 5870 1125
rect 6624 1111 6638 1125
rect 7416 1111 7430 1125
rect 71 1088 85 1102
rect 843 1088 857 1102
rect 2392 1088 2406 1102
rect 3328 1088 3342 1102
rect 4755 1088 4769 1102
rect 5640 1088 5654 1102
rect 6408 1088 6422 1102
rect 7296 1088 7310 1102
rect 47 1066 61 1080
rect 819 1066 833 1080
rect 2512 1066 2526 1080
rect 3232 1066 3246 1080
rect 4635 1066 4649 1080
rect 5736 1066 5750 1080
rect 6384 1066 6398 1080
rect 7176 1066 7190 1080
rect 23 1043 37 1057
rect 963 1043 977 1057
rect 2368 1043 2382 1057
rect 3208 1043 3222 1057
rect 4611 1043 4625 1057
rect 5616 1043 5630 1057
rect 6504 1043 6518 1057
rect 7152 1043 7166 1057
rect 8112 1043 8126 1057
rect 8304 1044 8318 1058
rect 8496 1044 8510 1058
rect 8688 1045 8702 1059
rect 8880 1044 8894 1058
rect 9072 1044 9086 1058
rect 723 1020 737 1034
rect 2152 1020 2166 1034
rect 2992 1020 3006 1034
rect 4515 1020 4529 1034
rect 5520 1020 5534 1034
rect 6192 1020 6206 1034
rect 6960 1020 6974 1034
rect 7896 1020 7910 1034
rect 8040 1018 8054 1032
rect 8568 1018 8582 1032
rect 8952 1018 8966 1032
rect 9144 1018 9158 1032
rect 9168 1017 9182 1031
rect 699 998 713 1012
rect 2128 998 2142 1012
rect 3112 998 3126 1012
rect 4419 998 4433 1012
rect 5400 998 5414 1012
rect 6288 998 6302 1012
rect 6936 998 6950 1012
rect 7776 998 7790 1012
rect 8976 995 8990 1009
rect 675 975 689 989
rect 2272 975 2286 989
rect 2968 975 2982 989
rect 4395 975 4409 989
rect 5376 975 5390 989
rect 6168 975 6182 989
rect 7056 975 7070 989
rect 7752 975 7766 989
rect 7992 974 8006 988
rect 8184 974 8198 988
rect 8760 974 8774 988
rect 8784 973 8798 987
rect 579 952 593 966
rect 1203 952 1217 966
rect 2752 952 2766 966
rect 4299 952 4313 966
rect 5280 952 5294 966
rect 5976 952 5990 966
rect 6744 952 6758 966
rect 7656 952 7670 966
rect 8592 951 8606 965
rect 555 930 569 944
rect 1179 930 1193 944
rect 2872 930 2886 944
rect 4203 930 4217 944
rect 5160 930 5174 944
rect 6072 930 6086 944
rect 6720 930 6734 944
rect 7536 930 7550 944
rect 8400 929 8414 943
rect 531 907 545 921
rect 1323 907 1337 921
rect 2728 907 2742 921
rect 4179 907 4193 921
rect 5136 907 5150 921
rect 5952 907 5966 921
rect 6840 907 6854 921
rect 7512 907 7526 921
rect 8208 907 8222 921
<< metal2 >>
rect 122 1126 134 1131
rect 24 904 36 1043
rect 48 904 60 1066
rect 72 904 84 1088
rect 192 904 204 1111
rect 676 989 688 1131
rect 700 1012 712 1131
rect 724 1034 736 1131
rect 532 904 544 907
rect 556 904 568 930
rect 580 904 592 952
rect 676 904 688 975
rect 700 904 712 998
rect 724 904 736 1020
rect 820 904 832 1066
rect 844 904 856 1088
rect 964 904 976 1043
rect 1084 904 1096 1111
rect 1180 904 1192 930
rect 1204 904 1216 952
rect 1324 904 1336 907
rect 2129 904 2141 998
rect 2153 904 2165 1020
rect 2273 904 2285 975
rect 2369 904 2381 1043
rect 2393 904 2405 1088
rect 2513 904 2525 1066
rect 2633 904 2645 1111
rect 2729 904 2741 907
rect 2753 904 2765 952
rect 2873 904 2885 930
rect 2969 904 2981 975
rect 2993 904 3005 1020
rect 3113 904 3125 998
rect 3209 904 3221 1043
rect 3233 904 3245 1066
rect 3329 904 3341 1088
rect 3449 904 3461 1111
rect 4180 904 4192 907
rect 4204 904 4216 930
rect 4300 904 4312 952
rect 4396 904 4408 975
rect 4420 904 4432 998
rect 4516 904 4528 1020
rect 4612 904 4624 1043
rect 4636 904 4648 1066
rect 4756 904 4768 1088
rect 4876 904 4888 1111
rect 5137 904 5149 907
rect 5161 904 5173 930
rect 5281 904 5293 952
rect 5377 904 5389 975
rect 5401 904 5413 998
rect 5521 904 5533 1020
rect 5617 904 5629 1043
rect 5641 904 5653 1088
rect 5737 904 5749 1066
rect 5857 904 5869 1111
rect 5953 904 5965 907
rect 5977 904 5989 952
rect 6073 904 6085 930
rect 6169 904 6181 975
rect 6193 904 6205 1020
rect 6289 904 6301 998
rect 6385 904 6397 1066
rect 6409 904 6421 1088
rect 6505 904 6517 1043
rect 6625 904 6637 1111
rect 6721 904 6733 930
rect 6745 904 6757 952
rect 6841 904 6853 907
rect 6937 904 6949 998
rect 6961 904 6973 1020
rect 7057 904 7069 975
rect 7153 904 7165 1043
rect 7177 904 7189 1066
rect 7297 904 7309 1088
rect 7417 904 7429 1111
rect 8113 1057 8125 1131
rect 7513 904 7525 907
rect 7537 904 7549 930
rect 7657 904 7669 952
rect 7753 904 7765 975
rect 7777 904 7789 998
rect 7897 904 7909 1020
rect 7993 904 8005 974
rect 8041 904 8053 1018
rect 8113 904 8125 1043
rect 8137 904 8149 1131
rect 8185 904 8197 974
rect 8209 904 8221 907
rect 8305 904 8317 1044
rect 8329 904 8341 1131
rect 8377 904 8389 1131
rect 8401 904 8413 929
rect 8497 904 8509 1044
rect 8521 904 8533 1131
rect 8569 904 8581 1018
rect 8593 904 8605 951
rect 8689 904 8701 1045
rect 8713 904 8725 1131
rect 8761 904 8773 974
rect 8785 904 8797 973
rect 8881 904 8893 1044
rect 8905 904 8917 1131
rect 8953 904 8965 1018
rect 8977 904 8989 995
rect 9073 904 9085 1044
rect 9097 904 9109 1131
rect 9145 904 9157 1018
rect 9169 904 9181 1017
rect 120 93 180 105
rect 240 83 252 105
rect 72 71 252 83
rect 72 0 84 71
rect 628 61 640 105
rect 772 83 784 105
rect 892 93 952 105
rect 1012 93 1072 105
rect 1132 95 1144 105
rect 1132 83 1236 95
rect 1252 93 1312 105
rect 1372 93 1980 105
rect 2201 93 2261 105
rect 772 71 1044 83
rect 628 49 828 61
rect 816 0 828 49
rect 1032 0 1044 71
rect 1224 0 1236 83
rect 1968 0 1980 93
rect 2321 83 2333 105
rect 2441 93 2501 105
rect 2561 93 2621 105
rect 2681 83 2693 105
rect 2801 93 2861 105
rect 2184 71 2333 83
rect 2376 71 2693 83
rect 2921 83 2933 105
rect 3041 93 3101 105
rect 3161 83 3173 105
rect 3257 93 3317 105
rect 3377 93 3437 105
rect 3497 93 3540 105
rect 4228 93 4288 105
rect 2921 71 3132 83
rect 3161 71 3348 83
rect 2184 0 2196 71
rect 2376 0 2388 71
rect 3120 0 3132 71
rect 3336 0 3348 71
rect 3528 0 3540 93
rect 4348 83 4360 105
rect 4444 93 4504 105
rect 4564 83 4576 105
rect 4684 93 4744 105
rect 4804 93 4864 105
rect 4924 83 4936 105
rect 5209 93 5269 105
rect 5329 95 5341 105
rect 5329 83 5436 95
rect 5449 93 5509 105
rect 5569 95 5581 105
rect 5569 83 5652 95
rect 5665 93 5725 105
rect 5785 93 5845 105
rect 5905 83 5917 105
rect 6001 93 6061 105
rect 4272 71 4360 83
rect 4488 71 4576 83
rect 4680 71 4936 83
rect 4272 0 4284 71
rect 4488 0 4500 71
rect 4680 0 4692 71
rect 5424 0 5436 83
rect 5640 0 5652 83
rect 5832 71 5917 83
rect 5832 0 5844 71
rect 6121 61 6133 105
rect 6217 93 6277 105
rect 6337 83 6349 105
rect 6433 93 6493 105
rect 6553 93 6613 105
rect 6673 83 6685 105
rect 6769 93 6829 105
rect 6889 83 6901 105
rect 6985 93 7045 105
rect 6337 71 6663 83
rect 6673 71 6871 83
rect 6889 71 7088 83
rect 6651 61 6663 71
rect 6859 61 6871 71
rect 6121 49 6588 61
rect 6651 49 6804 61
rect 6859 49 6996 61
rect 6576 0 6588 49
rect 6792 0 6804 49
rect 6984 0 6996 49
rect 7076 17 7088 71
rect 7105 39 7117 105
rect 7225 93 7285 105
rect 7345 93 7405 105
rect 7465 61 7477 105
rect 7585 93 7645 105
rect 7705 83 7717 105
rect 7825 93 7885 105
rect 7945 95 7957 105
rect 7945 83 9108 95
rect 7705 73 7931 83
rect 7705 71 8892 73
rect 7919 61 8892 71
rect 7465 51 7907 61
rect 7465 49 8148 51
rect 7895 39 8148 49
rect 7105 29 7883 39
rect 7105 27 7956 29
rect 7871 17 7956 27
rect 7076 5 7740 17
rect 7728 0 7740 5
rect 7944 0 7956 17
rect 8136 0 8148 39
rect 8880 0 8892 61
rect 9096 0 9108 83
use nor3 nor3_2
timestamp 1386235396
transform 1 0 0 0 1 105
box 0 0 144 799
use and2 and2_10
timestamp 1386234845
transform 1 0 144 0 1 105
box 0 0 120 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 508 0 1 105
box 0 0 144 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 652 0 1 105
box 0 0 144 799
use nor2 nor2_12
timestamp 1386235306
transform 1 0 796 0 1 105
box 0 0 120 799
use and2 and2_11
timestamp 1386234845
transform 1 0 916 0 1 105
box 0 0 120 799
use and2 and2_12
timestamp 1386234845
transform 1 0 1036 0 1 105
box 0 0 120 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 1156 0 1 105
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 1276 0 1 105
box 0 0 120 799
use nor2 nor2_6
timestamp 1386235306
transform 1 0 2105 0 1 105
box 0 0 120 799
use and2 and2_5
timestamp 1386234845
transform 1 0 2225 0 1 105
box 0 0 120 799
use nor2 nor2_13
timestamp 1386235306
transform 1 0 2345 0 1 105
box 0 0 120 799
use and2 and2_13
timestamp 1386234845
transform 1 0 2465 0 1 105
box 0 0 120 799
use and2 and2_14
timestamp 1386234845
transform 1 0 2585 0 1 105
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 2705 0 1 105
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 2825 0 1 105
box 0 0 120 799
use nor2 nor2_7
timestamp 1386235306
transform 1 0 2945 0 1 105
box 0 0 120 799
use and2 and2_6
timestamp 1386234845
transform 1 0 3065 0 1 105
box 0 0 120 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 3185 0 1 105
box 0 0 96 799
use nor2 nor2_14
timestamp 1386235306
transform 1 0 3281 0 1 105
box 0 0 120 799
use and2 and2_15
timestamp 1386234845
transform 1 0 3401 0 1 105
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 4156 0 1 105
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 4252 0 1 105
box 0 0 120 799
use nand2 nand2_3
timestamp 1386234792
transform 1 0 4372 0 1 105
box 0 0 96 799
use nor2 nor2_8
timestamp 1386235306
transform 1 0 4468 0 1 105
box 0 0 120 799
use nor2 nor2_15
timestamp 1386235306
transform 1 0 4588 0 1 105
box 0 0 120 799
use and2 and2_16
timestamp 1386234845
transform 1 0 4708 0 1 105
box 0 0 120 799
use and2 and2_17
timestamp 1386234845
transform 1 0 4828 0 1 105
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 5113 0 1 105
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 5233 0 1 105
box 0 0 120 799
use nor2 nor2_9
timestamp 1386235306
transform 1 0 5353 0 1 105
box 0 0 120 799
use and2 and2_7
timestamp 1386234845
transform 1 0 5473 0 1 105
box 0 0 120 799
use nand2 nand2_7
timestamp 1386234792
transform 1 0 5593 0 1 105
box 0 0 96 799
use nor2 nor2_16
timestamp 1386235306
transform 1 0 5689 0 1 105
box 0 0 120 799
use and2 and2_18
timestamp 1386234845
transform 1 0 5809 0 1 105
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 5929 0 1 105
box 0 0 96 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 6025 0 1 105
box 0 0 120 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 6145 0 1 105
box 0 0 96 799
use nor2 nor2_10
timestamp 1386235306
transform 1 0 6241 0 1 105
box 0 0 120 799
use nand2 nand2_8
timestamp 1386234792
transform 1 0 6361 0 1 105
box 0 0 96 799
use nor2 nor2_17
timestamp 1386235306
transform 1 0 6457 0 1 105
box 0 0 120 799
use and2 and2_19
timestamp 1386234845
transform 1 0 6577 0 1 105
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 6697 0 1 105
box 0 0 96 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 6793 0 1 105
box 0 0 120 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 6913 0 1 105
box 0 0 96 799
use nor2 nor2_11
timestamp 1386235306
transform 1 0 7009 0 1 105
box 0 0 120 799
use and2 and2_20
timestamp 1386234845
transform 1 0 7129 0 1 105
box 0 0 120 799
use and2 and2_21
timestamp 1386234845
transform 1 0 7249 0 1 105
box 0 0 120 799
use and2 and2_22
timestamp 1386234845
transform 1 0 7369 0 1 105
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 7489 0 1 105
box 0 0 120 799
use and2 and2_4
timestamp 1386234845
transform 1 0 7609 0 1 105
box 0 0 120 799
use and2 and2_8
timestamp 1386234845
transform 1 0 7729 0 1 105
box 0 0 120 799
use and2 and2_9
timestamp 1386234845
transform 1 0 7849 0 1 105
box 0 0 120 799
use tielow tielow_0
timestamp 1386086605
transform 1 0 7969 0 1 105
box 0 0 48 799
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 8017 0 1 105
box 0 0 48 799
use mux2 mux2_0
array 0 4 192 0 0 799
timestamp 1386235218
transform 1 0 8065 0 1 105
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 9025 0 1 105
box 0 0 192 799
<< labels >>
rlabel metal2 724 1131 736 1131 5 Rs2In[2]
rlabel metal2 700 1131 712 1131 5 Rs2In[1]
rlabel metal2 676 1131 688 1131 5 Rs2In[0]
rlabel metal2 122 1131 134 1131 5 We
rlabel metal2 8329 1131 8341 1131 5 Ir[14]
rlabel metal2 8521 1131 8533 1131 5 Ir[13]
rlabel metal2 8713 1131 8725 1131 5 Ir[12]
rlabel metal2 8905 1131 8917 1131 5 Ir[11]
rlabel metal2 8137 1131 8149 1131 5 Ir[15]
rlabel metal2 8377 1131 8389 1131 1 AluOR[0]
rlabel metal2 8113 1131 8125 1131 1 AluOR[1]
rlabel metal2 9097 1131 9109 1131 5 Cin
rlabel metal2 72 0 84 0 1 Rw[0]
rlabel metal2 816 0 828 0 1 Rs1[0]
rlabel metal2 1032 0 1044 0 1 Rs2[0]
rlabel metal2 2184 0 2196 0 1 Rs2[1]
rlabel metal2 2376 0 2388 0 1 Rw[2]
rlabel metal2 3120 0 3132 0 1 Rs1[2]
rlabel metal2 3336 0 3348 0 1 Rs2[2]
rlabel metal2 3528 0 3540 0 1 Rw[3]
rlabel metal2 4272 0 4284 0 1 Rs1[3]
rlabel metal2 5424 0 5436 0 1 Rs1[4]
rlabel metal2 5640 0 5652 0 1 Rs2[4]
rlabel metal2 5832 0 5844 0 1 Rw[5]
rlabel metal2 6576 0 6588 0 1 Rs1[5]
rlabel metal2 6792 0 6804 0 1 Rs2[5]
rlabel metal2 6984 0 6996 0 1 Rw[6]
rlabel metal2 7728 0 7740 0 1 Rs1[6]
rlabel metal2 7944 0 7956 0 1 Rs2[6]
rlabel metal2 8136 0 8148 0 1 Rw[7]
rlabel metal2 8880 0 8892 0 1 Rs1[7]
rlabel metal2 9096 0 9108 0 1 Rs2[7]
rlabel metal2 1224 0 1236 0 1 Rw[1]
rlabel metal2 1968 0 1980 0 1 Rs1[1]
rlabel metal2 4488 0 4500 0 1 Rs2[3]
rlabel metal2 4680 0 4692 0 1 Rw[4]
rlabel metal1 0 1045 0 1055 3 RwIn[0]
rlabel metal1 0 1068 0 1078 3 RwIn[1]
rlabel metal1 0 1090 0 1100 3 RwIn[2]
rlabel metal1 0 909 0 919 3 Rs1In[0]
rlabel metal1 0 932 0 942 3 Rs1In[1]
rlabel metal1 0 954 0 964 3 Rs1In[2]
rlabel metal1 9217 909 9217 919 7 AluOp[0]
rlabel metal1 9217 931 9217 941 7 AluOp[1]
rlabel metal1 9217 953 9217 963 7 AluOp[2]
rlabel metal1 9217 975 9217 985 7 AluOp[3]
rlabel metal1 9217 997 9217 1007 7 AluOp[4]
rlabel metal1 9217 1019 9217 1029 7 AluBin
<< end >>
