magic
tech c035u
timestamp 1395936165
<< nwell >>
rect 27435 46019 57587 46064
rect 27435 13033 27480 46019
rect 57542 13033 57587 46019
rect 27435 12988 57587 13033
<< nohmic >>
rect 27440 46027 57582 46059
rect 27440 13025 27472 46027
rect 57550 13025 57582 46027
rect 27440 12993 57582 13025
<< metal1 >>
rect 28368 45994 28378 46038
rect 28416 45994 28426 46038
rect 28368 45984 28426 45994
rect 27461 45096 27514 45106
rect 27504 45085 27514 45096
rect 28368 45085 28378 45984
rect 28464 45085 28474 46038
rect 31800 46021 31810 46038
rect 31848 45994 31858 46038
rect 35328 46021 35338 46038
rect 29952 45984 31858 45994
rect 29952 45970 29962 45984
rect 35376 45994 35386 46038
rect 38856 45994 38866 46038
rect 38904 46021 38914 46038
rect 39048 46021 39058 46038
rect 45912 45994 45922 46038
rect 45960 46021 45970 46038
rect 46104 46021 46114 46038
rect 49416 45994 49426 46038
rect 49464 46021 49474 46038
rect 49608 46021 49618 46038
rect 52944 45994 52954 46038
rect 31885 45984 35386 45994
rect 35400 45984 52978 45994
rect 29928 45960 29962 45970
rect 29928 45949 29938 45960
rect 35400 45970 35410 45984
rect 52968 45973 52978 45984
rect 52992 45973 53002 46038
rect 53136 46021 53146 46038
rect 53016 45984 55546 45994
rect 53016 45973 53026 45984
rect 55536 45973 55546 45984
rect 29989 45960 35410 45970
rect 38917 45960 52943 45970
rect 53040 45960 55522 45970
rect 29952 45936 31799 45946
rect 29952 45922 29962 45936
rect 31813 45936 35327 45946
rect 53040 45946 53050 45960
rect 45973 45936 53050 45946
rect 53064 45936 55487 45946
rect 29904 45912 29962 45922
rect 30000 45912 31871 45922
rect 29904 45058 29914 45912
rect 30000 45898 30010 45912
rect 29952 45888 30010 45898
rect 27461 45048 29914 45058
rect 27504 40642 27514 45023
rect 27528 40669 27538 45048
rect 28368 44266 28378 45023
rect 28464 44293 28474 45023
rect 29928 44293 29938 45887
rect 29952 44293 29962 45888
rect 29976 44293 29986 45863
rect 35328 44461 35338 45935
rect 39048 44581 39058 45935
rect 53064 45922 53074 45936
rect 55512 45946 55522 45960
rect 55512 45936 55570 45946
rect 46117 45912 53074 45922
rect 55309 45912 55522 45922
rect 55512 45901 55522 45912
rect 55560 45901 55570 45936
rect 52981 45888 55474 45898
rect 49464 44581 49474 45887
rect 49608 44581 49618 45887
rect 52944 45874 52954 45887
rect 52944 45864 53015 45874
rect 55464 45874 55474 45888
rect 55464 45864 55594 45874
rect 53136 45850 53146 45863
rect 53136 45840 55474 45850
rect 52992 44578 53002 45839
rect 55296 44581 55306 45815
rect 55464 44581 55474 45840
rect 55488 44581 55498 45839
rect 55512 44581 55522 45839
rect 52992 44568 53015 44578
rect 55536 44578 55546 45839
rect 55560 44605 55570 45839
rect 55584 45298 55594 45864
rect 55584 45288 57561 45298
rect 57504 45277 57514 45288
rect 57480 45240 57561 45250
rect 57480 45157 57490 45240
rect 57504 45130 57514 45215
rect 57456 45120 57514 45130
rect 55536 44568 55583 44578
rect 36576 44544 55607 44554
rect 36576 44461 36586 44544
rect 53005 44520 55343 44530
rect 55477 44520 55642 44530
rect 39048 44461 39058 44519
rect 47557 44496 55535 44506
rect 55632 44506 55642 44520
rect 55632 44496 55690 44506
rect 47352 44472 55655 44482
rect 47352 44461 47362 44472
rect 55680 44482 55690 44496
rect 55680 44472 55714 44482
rect 47725 44448 55679 44458
rect 55704 44458 55714 44472
rect 55704 44448 55786 44458
rect 55776 44437 55786 44448
rect 34152 44424 55751 44434
rect 28368 44256 30010 44266
rect 27504 40632 27562 40642
rect 27461 40608 27514 40618
rect 27504 40597 27514 40608
rect 27528 40570 27538 40607
rect 27461 40560 27538 40570
rect 27504 36181 27514 40535
rect 27528 36178 27538 40560
rect 27552 36205 27562 40632
rect 27528 36168 27586 36178
rect 27461 36144 27538 36154
rect 27528 36133 27538 36144
rect 27576 36106 27586 36168
rect 27461 36096 27586 36106
rect 27504 31765 27514 36071
rect 27528 31762 27538 36071
rect 27552 31789 27562 36071
rect 27528 31752 27586 31762
rect 27461 31728 27538 31738
rect 27504 27373 27514 31703
rect 27528 27373 27538 31728
rect 27552 27373 27562 31727
rect 27576 27370 27586 31752
rect 27576 27360 27610 27370
rect 27461 27336 27586 27346
rect 27504 22909 27514 27311
rect 27528 22906 27538 27311
rect 27552 22933 27562 27311
rect 27576 23458 27586 27336
rect 27600 23506 27610 27360
rect 28464 23533 28474 44231
rect 29976 44218 29986 44231
rect 29904 44208 29986 44218
rect 29904 44194 29914 44208
rect 29880 44184 29914 44194
rect 30000 44194 30010 44256
rect 30000 44184 30479 44194
rect 29880 23533 29890 44184
rect 29904 44160 30610 44170
rect 29904 23533 29914 44160
rect 30600 44149 30610 44160
rect 34152 44149 34162 44424
rect 35544 44400 55463 44410
rect 35328 44269 35338 44399
rect 35544 44365 35554 44400
rect 55501 44400 55799 44410
rect 44832 44376 55487 44386
rect 44832 44365 44842 44376
rect 55573 44376 55823 44386
rect 45565 44352 55559 44362
rect 55597 44352 55858 44362
rect 35352 44328 55738 44338
rect 35352 44269 35362 44328
rect 44568 44304 55714 44314
rect 35544 44269 35554 44303
rect 36576 44269 36586 44303
rect 39048 44269 39058 44303
rect 44568 44269 44578 44304
rect 55704 44293 55714 44304
rect 55728 44293 55738 44328
rect 55752 44293 55762 44327
rect 55776 44293 55786 44327
rect 47616 44280 55631 44290
rect 47616 44269 47626 44280
rect 55800 44290 55810 44327
rect 55848 44317 55858 44352
rect 55800 44280 55882 44290
rect 55872 44269 55882 44280
rect 49621 44256 52991 44266
rect 53029 44256 55810 44266
rect 55800 44245 55810 44256
rect 34392 44232 55583 44242
rect 34392 44149 34402 44232
rect 55824 44242 55834 44255
rect 55824 44232 55895 44242
rect 39061 44208 55919 44218
rect 35328 44170 35338 44207
rect 49477 44184 55330 44194
rect 35328 44160 55295 44170
rect 55320 44170 55330 44184
rect 55357 44184 55823 44194
rect 55861 44184 55954 44194
rect 55320 44160 55858 44170
rect 55296 44149 55306 44159
rect 29928 23533 29938 44135
rect 29952 23533 29962 44135
rect 55464 41365 55474 44135
rect 55488 41365 55498 44135
rect 55512 41365 55522 44135
rect 55536 41365 55546 44135
rect 55560 41365 55570 44135
rect 55584 41365 55594 44135
rect 55608 41365 55618 44135
rect 55632 41365 55642 44135
rect 55656 41365 55666 44135
rect 55680 41365 55690 44135
rect 55704 41365 55714 44135
rect 55728 41365 55738 44135
rect 55752 41365 55762 44135
rect 55776 41365 55786 44135
rect 55800 41365 55810 44135
rect 55824 41365 55834 44135
rect 55848 41365 55858 44160
rect 55872 41365 55882 44159
rect 55896 41365 55906 44159
rect 55920 41365 55930 44159
rect 55417 41338 55450 41346
rect 55944 41338 55954 44184
rect 55417 41336 55954 41338
rect 55440 41328 55954 41336
rect 55417 41270 55450 41280
rect 55440 41266 55450 41270
rect 55920 41266 55930 41303
rect 55440 41256 55930 41266
rect 55464 40189 55474 41231
rect 55488 40189 55498 41231
rect 55512 40189 55522 41231
rect 55536 40189 55546 41231
rect 55560 40189 55570 41231
rect 55584 40189 55594 41231
rect 55608 40189 55618 41231
rect 55632 40189 55642 41231
rect 55656 40189 55666 41231
rect 55680 40189 55690 41231
rect 55704 40189 55714 41231
rect 55728 40189 55738 41231
rect 55752 40189 55762 41231
rect 55776 40189 55786 41231
rect 55800 40189 55810 41231
rect 55824 40189 55834 41231
rect 55848 40189 55858 41231
rect 55872 40189 55882 41231
rect 55417 40162 55450 40170
rect 55896 40162 55906 41231
rect 57456 40837 57466 45120
rect 57504 45096 57561 45106
rect 57480 40861 57490 45095
rect 57504 40861 57514 45096
rect 57469 40824 57561 40834
rect 57432 40800 57503 40810
rect 57432 40693 57442 40800
rect 57504 40776 57561 40786
rect 57456 40693 57466 40775
rect 57480 40666 57490 40775
rect 57504 40669 57514 40776
rect 55417 40160 55906 40162
rect 55440 40152 55906 40160
rect 57408 40656 57490 40666
rect 55417 40094 55450 40104
rect 55440 40090 55450 40094
rect 55872 40090 55882 40127
rect 55440 40080 55882 40090
rect 55464 39013 55474 40055
rect 55488 39013 55498 40055
rect 55512 39013 55522 40055
rect 55536 39013 55546 40055
rect 55560 39013 55570 40055
rect 55584 39013 55594 40055
rect 55608 39013 55618 40055
rect 55632 39013 55642 40055
rect 55656 39013 55666 40055
rect 55680 39013 55690 40055
rect 55704 39013 55714 40055
rect 55728 39013 55738 40055
rect 55752 39013 55762 40055
rect 55776 39013 55786 40055
rect 55800 39013 55810 40055
rect 55824 39013 55834 40055
rect 55417 38986 55450 38994
rect 55848 38986 55858 40055
rect 55417 38984 55858 38986
rect 55440 38976 55858 38984
rect 55417 38918 55450 38928
rect 55440 38914 55450 38918
rect 55824 38914 55834 38951
rect 55440 38904 55834 38914
rect 55464 37837 55474 38879
rect 55488 37837 55498 38879
rect 55512 37837 55522 38879
rect 55536 37837 55546 38879
rect 55560 37837 55570 38879
rect 55584 37837 55594 38879
rect 55608 37837 55618 38879
rect 55632 37837 55642 38879
rect 55656 37837 55666 38879
rect 55680 37837 55690 38879
rect 55704 37837 55714 38879
rect 55728 37837 55738 38879
rect 55752 37837 55762 38879
rect 55776 37837 55786 38879
rect 55417 37810 55450 37818
rect 55800 37810 55810 38879
rect 55417 37808 55810 37810
rect 55440 37800 55810 37808
rect 55417 37742 55450 37752
rect 55440 37738 55450 37742
rect 55776 37738 55786 37775
rect 55440 37728 55786 37738
rect 55464 36661 55474 37703
rect 55488 36661 55498 37703
rect 55512 36661 55522 37703
rect 55536 36661 55546 37703
rect 55560 36661 55570 37703
rect 55584 36661 55594 37703
rect 55608 36661 55618 37703
rect 55632 36661 55642 37703
rect 55656 36661 55666 37703
rect 55680 36661 55690 37703
rect 55704 36661 55714 37703
rect 55728 36661 55738 37703
rect 55752 36661 55762 37703
rect 55417 36634 55450 36642
rect 57408 36634 57418 40656
rect 57480 40632 57561 40642
rect 55417 36632 57418 36634
rect 55440 36624 57418 36632
rect 55417 36566 55450 36576
rect 55440 36562 55450 36566
rect 57432 36562 57442 40631
rect 55440 36552 57442 36562
rect 55464 35485 55474 36527
rect 55488 35485 55498 36527
rect 55512 35485 55522 36527
rect 55536 35485 55546 36527
rect 55560 35485 55570 36527
rect 55584 35485 55594 36527
rect 55608 35485 55618 36527
rect 55632 35485 55642 36527
rect 55656 35485 55666 36527
rect 55680 35485 55690 36527
rect 55704 35485 55714 36527
rect 55728 35485 55738 36527
rect 55752 35485 55762 36527
rect 57456 36370 57466 40631
rect 57480 36397 57490 40632
rect 57504 36397 57514 40607
rect 57456 36360 57561 36370
rect 57456 36336 57479 36346
rect 57456 36229 57466 36336
rect 57480 36312 57561 36322
rect 57480 36229 57490 36312
rect 57504 36202 57514 36287
rect 57432 36192 57514 36202
rect 55417 35458 55450 35466
rect 57432 35458 57442 36192
rect 57504 36168 57561 36178
rect 55417 35456 57442 35458
rect 55440 35448 57442 35456
rect 55417 35390 55450 35400
rect 55440 35386 55450 35390
rect 57456 35386 57466 36167
rect 55440 35376 57466 35386
rect 55464 34309 55474 35351
rect 55488 34309 55498 35351
rect 55512 34309 55522 35351
rect 55536 34309 55546 35351
rect 55560 34309 55570 35351
rect 55584 34309 55594 35351
rect 55608 34309 55618 35351
rect 55632 34309 55642 35351
rect 55656 34309 55666 35351
rect 55680 34309 55690 35351
rect 55704 34309 55714 35351
rect 55728 34309 55738 35351
rect 55752 34309 55762 35351
rect 55417 34282 55450 34290
rect 57480 34282 57490 36167
rect 55417 34280 57490 34282
rect 55440 34272 57490 34280
rect 55417 34214 55450 34224
rect 55440 34210 55450 34214
rect 57504 34210 57514 36168
rect 55440 34200 57514 34210
rect 55464 33133 55474 34175
rect 55488 33133 55498 34175
rect 55512 33133 55522 34175
rect 55536 33133 55546 34175
rect 55560 33133 55570 34175
rect 55584 33133 55594 34175
rect 55608 33133 55618 34175
rect 55632 33133 55642 34175
rect 55656 33133 55666 34175
rect 55680 33133 55690 34175
rect 55704 33133 55714 34175
rect 55728 33133 55738 34175
rect 55752 33130 55762 34175
rect 55752 33120 55786 33130
rect 55417 33106 55450 33114
rect 55417 33104 55762 33106
rect 55440 33096 55762 33104
rect 55752 33085 55762 33096
rect 55776 33085 55786 33120
rect 55608 33058 55618 33071
rect 55608 33048 55810 33058
rect 55417 33038 55450 33048
rect 55440 33034 55450 33038
rect 55440 33024 55618 33034
rect 55464 31957 55474 32999
rect 55488 31954 55498 32999
rect 55512 31981 55522 32999
rect 55536 31981 55546 32999
rect 55560 31981 55570 32999
rect 55584 31981 55594 32999
rect 55608 31981 55618 33024
rect 55632 31981 55642 33023
rect 55656 31981 55666 33023
rect 55680 31981 55690 33023
rect 55704 31981 55714 33023
rect 55728 31981 55738 33023
rect 55752 31981 55762 33023
rect 55776 31981 55786 33023
rect 55800 31981 55810 33048
rect 55488 31944 55834 31954
rect 55417 31930 55450 31938
rect 55417 31928 55498 31930
rect 55440 31920 55498 31928
rect 55488 31885 55498 31920
rect 55417 31862 55450 31872
rect 55512 31882 55522 31919
rect 55824 31909 55834 31944
rect 55512 31872 55858 31882
rect 55440 31858 55450 31862
rect 55440 31848 55522 31858
rect 55464 30778 55474 31823
rect 55488 30805 55498 31823
rect 55512 30805 55522 31848
rect 55536 30805 55546 31847
rect 55560 30805 55570 31847
rect 55584 30805 55594 31847
rect 55608 30805 55618 31847
rect 55632 30805 55642 31847
rect 55656 30805 55666 31847
rect 55680 30805 55690 31847
rect 55704 30805 55714 31847
rect 55728 30805 55738 31847
rect 55752 30805 55762 31847
rect 55776 30805 55786 31847
rect 55800 30805 55810 31847
rect 55824 30805 55834 31847
rect 55848 31762 55858 31872
rect 55848 31752 57527 31762
rect 55464 30768 55858 30778
rect 55417 30754 55450 30762
rect 55417 30752 55474 30754
rect 55440 30744 55474 30752
rect 55464 30709 55474 30744
rect 55488 30709 55498 30743
rect 55512 30709 55522 30743
rect 55536 30709 55546 30743
rect 55560 30709 55570 30743
rect 55584 30709 55594 30743
rect 55608 30709 55618 30743
rect 55632 30709 55642 30743
rect 55656 30709 55666 30743
rect 55680 30709 55690 30743
rect 55704 30709 55714 30743
rect 55417 30686 55450 30696
rect 55728 30706 55738 30743
rect 55848 30733 55858 30768
rect 55728 30696 55882 30706
rect 55440 30682 55450 30686
rect 55440 30672 55738 30682
rect 55464 29605 55474 30647
rect 55488 29605 55498 30647
rect 55512 29605 55522 30647
rect 55536 29602 55546 30647
rect 55560 29629 55570 30647
rect 55584 29629 55594 30647
rect 55608 29629 55618 30647
rect 55632 29629 55642 30647
rect 55656 29629 55666 30647
rect 55680 29629 55690 30647
rect 55704 29629 55714 30647
rect 55728 29629 55738 30672
rect 55752 29629 55762 30671
rect 55776 29629 55786 30671
rect 55800 29629 55810 30671
rect 55824 29629 55834 30671
rect 55848 29629 55858 30671
rect 55872 29629 55882 30696
rect 55536 29592 55906 29602
rect 55417 29578 55450 29586
rect 55417 29576 55546 29578
rect 55440 29568 55546 29576
rect 55536 29533 55546 29568
rect 55560 29533 55570 29567
rect 55584 29533 55594 29567
rect 55608 29533 55618 29567
rect 55417 29510 55450 29520
rect 55632 29530 55642 29567
rect 55896 29557 55906 29592
rect 55632 29520 55930 29530
rect 55440 29506 55450 29510
rect 55440 29496 55642 29506
rect 55464 28429 55474 29471
rect 55488 28429 55498 29471
rect 55512 28429 55522 29471
rect 55536 28429 55546 29471
rect 55560 28429 55570 29471
rect 55584 28429 55594 29471
rect 55608 28429 55618 29471
rect 55632 28429 55642 29496
rect 55656 28429 55666 29495
rect 55680 28426 55690 29495
rect 55704 28453 55714 29495
rect 55728 28453 55738 29495
rect 55752 28453 55762 29495
rect 55776 28453 55786 29495
rect 55800 28453 55810 29495
rect 55824 28453 55834 29495
rect 55848 28453 55858 29495
rect 55872 28453 55882 29495
rect 55896 28453 55906 29495
rect 55920 28453 55930 29520
rect 55680 28416 55954 28426
rect 55417 28402 55450 28410
rect 55417 28400 55690 28402
rect 55440 28392 55690 28400
rect 55680 28381 55690 28392
rect 55944 28381 55954 28416
rect 55584 28354 55594 28367
rect 55584 28344 55978 28354
rect 55417 28334 55450 28344
rect 55440 28330 55450 28334
rect 55440 28320 55594 28330
rect 55464 27253 55474 28295
rect 55488 27253 55498 28295
rect 55512 27253 55522 28295
rect 55536 27253 55546 28295
rect 55560 27253 55570 28295
rect 55584 27253 55594 28320
rect 55608 27253 55618 28319
rect 55632 27253 55642 28319
rect 55656 27253 55666 28319
rect 55680 27253 55690 28319
rect 55704 27253 55714 28319
rect 55728 27253 55738 28319
rect 55752 27253 55762 28319
rect 55776 27253 55786 28319
rect 55800 27253 55810 28319
rect 55824 27253 55834 28319
rect 55848 27250 55858 28319
rect 55872 27277 55882 28319
rect 55896 27277 55906 28319
rect 55920 27277 55930 28319
rect 55944 27277 55954 28319
rect 55968 27277 55978 28344
rect 55848 27240 56002 27250
rect 55417 27226 55450 27234
rect 55417 27224 55858 27226
rect 55440 27216 55858 27224
rect 55848 27205 55858 27216
rect 55992 27205 56002 27240
rect 55584 27178 55594 27191
rect 55584 27168 56026 27178
rect 55417 27158 55450 27168
rect 55440 27154 55450 27158
rect 55440 27144 55594 27154
rect 55464 26077 55474 27119
rect 55488 26077 55498 27119
rect 55512 26077 55522 27119
rect 55536 26077 55546 27119
rect 55560 26074 55570 27119
rect 55584 26101 55594 27144
rect 55608 26101 55618 27143
rect 55632 26101 55642 27143
rect 55656 26101 55666 27143
rect 55680 26101 55690 27143
rect 55704 26101 55714 27143
rect 55728 26101 55738 27143
rect 55752 26101 55762 27143
rect 55776 26101 55786 27143
rect 55800 26101 55810 27143
rect 55824 26101 55834 27143
rect 55848 26101 55858 27143
rect 55872 26101 55882 27143
rect 55896 26101 55906 27143
rect 55920 26101 55930 27143
rect 55944 26101 55954 27143
rect 55968 26101 55978 27143
rect 55992 26101 56002 27143
rect 56016 26101 56026 27168
rect 55560 26064 56050 26074
rect 55417 26050 55450 26058
rect 55417 26048 55570 26050
rect 55440 26040 55570 26048
rect 55560 26029 55570 26040
rect 56040 26029 56050 26064
rect 55536 26002 55546 26015
rect 55536 25992 56074 26002
rect 55417 25982 55450 25992
rect 55440 25978 55450 25982
rect 55440 25968 55546 25978
rect 55464 24901 55474 25943
rect 55488 24901 55498 25943
rect 55512 24901 55522 25943
rect 55536 24901 55546 25968
rect 55560 24901 55570 25967
rect 55584 24901 55594 25967
rect 55608 24901 55618 25967
rect 55632 24901 55642 25967
rect 55656 24901 55666 25967
rect 55680 24901 55690 25967
rect 55704 24898 55714 25967
rect 55728 24925 55738 25967
rect 55752 24925 55762 25967
rect 55776 24925 55786 25967
rect 55800 24925 55810 25967
rect 55824 24925 55834 25967
rect 55848 24925 55858 25967
rect 55872 24925 55882 25967
rect 55896 24925 55906 25967
rect 55920 24925 55930 25967
rect 55944 24925 55954 25967
rect 55968 24925 55978 25967
rect 55992 24925 56002 25967
rect 56016 24925 56026 25967
rect 56040 24925 56050 25967
rect 56064 24925 56074 25992
rect 55704 24888 56098 24898
rect 55417 24874 55450 24882
rect 55417 24872 55714 24874
rect 55440 24864 55714 24872
rect 55704 24829 55714 24864
rect 55728 24829 55738 24863
rect 55752 24829 55762 24863
rect 55776 24829 55786 24863
rect 55800 24829 55810 24863
rect 55824 24829 55834 24863
rect 55848 24829 55858 24863
rect 55872 24829 55882 24863
rect 55896 24829 55906 24863
rect 55920 24829 55930 24863
rect 55944 24829 55954 24863
rect 55968 24829 55978 24863
rect 55992 24829 56002 24863
rect 55417 24806 55450 24816
rect 56016 24826 56026 24863
rect 56088 24853 56098 24888
rect 56016 24816 56122 24826
rect 55440 24802 55450 24806
rect 55440 24792 56026 24802
rect 55464 23725 55474 24767
rect 55488 23725 55498 24767
rect 55512 23725 55522 24767
rect 55536 23722 55546 24767
rect 55560 23749 55570 24767
rect 55584 23749 55594 24767
rect 55608 23749 55618 24767
rect 55632 23749 55642 24767
rect 55656 23749 55666 24767
rect 55680 23749 55690 24767
rect 55704 23749 55714 24767
rect 55728 23749 55738 24767
rect 55752 23749 55762 24767
rect 55776 23749 55786 24767
rect 55800 23749 55810 24767
rect 55824 23749 55834 24767
rect 55848 23749 55858 24767
rect 55872 23749 55882 24767
rect 55896 23749 55906 24767
rect 55920 23749 55930 24767
rect 55944 23749 55954 24767
rect 55968 23749 55978 24767
rect 55992 23749 56002 24767
rect 56016 23749 56026 24792
rect 56040 23749 56050 24791
rect 56064 23749 56074 24791
rect 56088 23749 56098 24791
rect 56112 23749 56122 24816
rect 55536 23712 56146 23722
rect 55417 23698 55450 23706
rect 55417 23696 55546 23698
rect 55440 23688 55546 23696
rect 55536 23653 55546 23688
rect 55560 23653 55570 23687
rect 55584 23653 55594 23687
rect 55608 23653 55618 23687
rect 55632 23653 55642 23687
rect 55656 23653 55666 23687
rect 55680 23653 55690 23687
rect 55704 23653 55714 23687
rect 55417 23630 55450 23640
rect 55728 23650 55738 23687
rect 56136 23677 56146 23712
rect 55728 23640 56170 23650
rect 55440 23626 55450 23630
rect 55440 23616 55738 23626
rect 55464 23533 55474 23591
rect 55488 23533 55498 23591
rect 55512 23533 55522 23591
rect 55536 23533 55546 23591
rect 55560 23533 55570 23591
rect 55584 23533 55594 23591
rect 55608 23533 55618 23591
rect 55632 23533 55642 23591
rect 55656 23533 55666 23591
rect 55680 23533 55690 23591
rect 55704 23533 55714 23591
rect 55728 23533 55738 23616
rect 55752 23533 55762 23615
rect 55776 23533 55786 23615
rect 55800 23533 55810 23615
rect 55824 23533 55834 23615
rect 55848 23533 55858 23615
rect 55872 23533 55882 23615
rect 55896 23533 55906 23615
rect 55920 23533 55930 23615
rect 55944 23533 55954 23615
rect 55968 23533 55978 23615
rect 55992 23533 56002 23615
rect 56016 23533 56026 23615
rect 56040 23533 56050 23615
rect 56064 23533 56074 23615
rect 56088 23533 56098 23615
rect 56112 23533 56122 23615
rect 56136 23533 56146 23615
rect 56160 23533 56170 23640
rect 30480 23506 30490 23519
rect 27600 23496 29986 23506
rect 29976 23485 29986 23496
rect 30200 23496 30490 23506
rect 30200 23485 30210 23496
rect 30667 23506 30677 23519
rect 30517 23496 30677 23506
rect 30229 23472 30594 23482
rect 30229 23458 30239 23472
rect 30620 23458 30630 23471
rect 27576 23448 30239 23458
rect 30312 23448 30630 23458
rect 27528 22896 27586 22906
rect 27461 22872 27538 22882
rect 27504 18445 27514 22847
rect 27528 22618 27538 22872
rect 27552 22642 27562 22871
rect 27576 22666 27586 22896
rect 28464 22693 28474 23423
rect 29880 22762 29890 23423
rect 29869 22752 29890 22762
rect 29904 22738 29914 23423
rect 29845 22728 29914 22738
rect 29928 22714 29938 23423
rect 29797 22704 29938 22714
rect 29952 22690 29962 23423
rect 29976 22693 29986 23423
rect 29749 22680 29962 22690
rect 30010 22690 30020 23423
rect 30033 22714 30043 23389
rect 30056 22738 30066 23423
rect 30079 22762 30089 23389
rect 30102 22786 30112 23423
rect 30125 22810 30135 23389
rect 30148 22834 30158 23423
rect 30171 22858 30181 23389
rect 30201 22885 30211 23423
rect 30312 22861 30322 23448
rect 30644 23434 30654 23471
rect 30336 23424 30654 23434
rect 30336 22861 30346 23424
rect 30360 23400 30503 23410
rect 30360 22861 30370 23400
rect 30171 22848 30240 22858
rect 30148 22824 30383 22834
rect 30125 22800 30407 22810
rect 31944 22810 31954 23519
rect 32136 22834 32146 23519
rect 32136 22824 32351 22834
rect 32928 22834 32938 23519
rect 32928 22824 33167 22834
rect 33480 22834 33490 23519
rect 33696 22858 33706 23519
rect 33696 22848 34007 22858
rect 33480 22824 34031 22834
rect 34440 22834 34450 23519
rect 34608 22858 34618 23519
rect 34992 22882 35002 23519
rect 35184 22906 35194 23519
rect 35184 22896 35207 22906
rect 35400 22906 35410 23519
rect 35400 22896 35639 22906
rect 36144 22906 36154 23519
rect 36312 22930 36322 23519
rect 36312 22920 37247 22930
rect 36144 22896 37967 22906
rect 34992 22872 38447 22882
rect 34608 22848 39335 22858
rect 34440 22824 40223 22834
rect 31944 22800 38423 22810
rect 38461 22800 41338 22810
rect 30102 22776 33983 22786
rect 34045 22776 41303 22786
rect 41328 22786 41338 22800
rect 41328 22776 42143 22786
rect 30079 22752 35183 22762
rect 35221 22752 42167 22762
rect 30056 22728 35615 22738
rect 35653 22728 42983 22738
rect 30033 22704 37223 22714
rect 37261 22704 44567 22714
rect 30010 22680 37943 22690
rect 37981 22680 44605 22690
rect 27576 22656 28391 22666
rect 28405 22656 30167 22666
rect 30181 22656 30199 22666
rect 30254 22656 32327 22666
rect 32365 22656 39311 22666
rect 39349 22656 42959 22666
rect 42997 22656 45383 22666
rect 45720 22666 45730 23519
rect 45912 22690 45922 23519
rect 46152 22714 46162 23519
rect 53856 23506 53866 23519
rect 50976 23496 53866 23506
rect 46152 22704 46199 22714
rect 45912 22680 47663 22690
rect 45720 22656 48572 22666
rect 27552 22632 29879 22642
rect 29989 22632 30284 22642
rect 30421 22632 33959 22642
rect 34021 22632 42119 22642
rect 42157 22632 44543 22642
rect 44581 22632 46175 22642
rect 46213 22632 48634 22642
rect 30312 22618 30322 22631
rect 27528 22608 30322 22618
rect 30312 22597 30322 22608
rect 30336 22597 30346 22631
rect 30360 22597 30370 22631
rect 30384 22618 30394 22631
rect 30384 22608 33154 22618
rect 33144 22597 33154 22608
rect 33181 22608 40210 22618
rect 40200 22597 40210 22608
rect 40237 22608 42154 22618
rect 42144 22597 42154 22608
rect 42181 22608 44587 22618
rect 44577 22597 44587 22608
rect 44619 22608 47650 22618
rect 47640 22597 47650 22608
rect 48624 22618 48634 22632
rect 47677 22608 48607 22618
rect 48624 22608 49402 22618
rect 48597 22597 48607 22608
rect 49392 22597 49402 22608
rect 50976 22597 50986 23496
rect 54792 23506 54802 23519
rect 53893 23496 54802 23506
rect 54888 23506 54898 23519
rect 54829 23496 54898 23506
rect 51672 23472 54599 23482
rect 51672 22597 51682 23472
rect 54637 23472 54743 23482
rect 54781 23472 54839 23482
rect 51816 23448 54815 23458
rect 51816 22597 51826 23448
rect 52608 23424 54767 23434
rect 52608 22597 52618 23424
rect 53424 23400 53879 23410
rect 53424 22597 53434 23400
rect 54216 23400 54623 23410
rect 54216 22597 54226 23400
rect 54960 22618 54970 23519
rect 55296 23506 55306 23519
rect 55296 23496 56194 23506
rect 55464 22618 55474 23471
rect 55488 22642 55498 23471
rect 55512 22666 55522 23471
rect 55536 22690 55546 23471
rect 55560 22714 55570 23471
rect 55584 22738 55594 23471
rect 55608 22762 55618 23471
rect 55632 22786 55642 23471
rect 55656 22810 55666 23471
rect 55680 22834 55690 23471
rect 55704 22858 55714 23471
rect 55728 22882 55738 23471
rect 55752 22906 55762 23471
rect 55776 22930 55786 23471
rect 55800 22954 55810 23471
rect 55824 22978 55834 23471
rect 55848 23002 55858 23471
rect 55872 23026 55882 23471
rect 55896 23050 55906 23471
rect 55920 23074 55930 23471
rect 55944 23098 55954 23471
rect 55968 23122 55978 23471
rect 55992 23146 56002 23471
rect 56016 23170 56026 23471
rect 56040 23194 56050 23471
rect 56064 23218 56074 23471
rect 56088 23242 56098 23471
rect 56112 23266 56122 23471
rect 56136 23290 56146 23471
rect 56160 23314 56170 23471
rect 56184 23341 56194 23496
rect 56160 23304 56519 23314
rect 56136 23280 56543 23290
rect 56112 23256 56567 23266
rect 56088 23232 56591 23242
rect 56064 23208 56615 23218
rect 56040 23184 56639 23194
rect 56016 23160 56663 23170
rect 55992 23136 56687 23146
rect 55968 23112 56711 23122
rect 55944 23088 56735 23098
rect 55920 23064 56759 23074
rect 55896 23040 56783 23050
rect 55872 23016 56807 23026
rect 55848 22992 56831 23002
rect 55824 22968 56855 22978
rect 55800 22944 56879 22954
rect 57504 22944 57561 22954
rect 57504 22933 57514 22944
rect 55776 22920 56903 22930
rect 55752 22896 57561 22906
rect 55728 22872 56927 22882
rect 55704 22848 56951 22858
rect 55680 22824 56975 22834
rect 55656 22800 56999 22810
rect 57504 22789 57514 22871
rect 55632 22776 57023 22786
rect 55608 22752 57561 22762
rect 55584 22728 57047 22738
rect 55560 22704 57071 22714
rect 57504 22714 57514 22727
rect 57109 22704 57514 22714
rect 55536 22680 57143 22690
rect 55512 22656 57407 22666
rect 55488 22632 57455 22642
rect 54960 22608 55042 22618
rect 55464 22608 57514 22618
rect 55032 22597 55042 22608
rect 27461 18408 27538 18418
rect 27504 14578 27514 18383
rect 27528 14605 27538 18408
rect 28392 14584 28402 22583
rect 28464 18178 28474 22583
rect 29736 22394 29746 22583
rect 29784 22429 29794 22583
rect 29832 22429 29842 22583
rect 29856 22429 29866 22583
rect 29880 22429 29890 22583
rect 29736 22384 29903 22394
rect 56520 22374 56530 22583
rect 56544 22374 56554 22583
rect 56568 22374 56578 22583
rect 56592 22374 56602 22583
rect 56616 22374 56626 22583
rect 29797 22360 29903 22370
rect 56640 22347 56650 22583
rect 56664 22350 56674 22583
rect 56688 22350 56698 22583
rect 56712 22350 56722 22583
rect 56736 22350 56746 22583
rect 56509 22337 56650 22347
rect 29832 18205 29842 22335
rect 29856 18205 29866 22335
rect 29880 18205 29890 22335
rect 56760 22323 56770 22583
rect 56784 22326 56794 22583
rect 56808 22326 56818 22583
rect 56832 22326 56842 22583
rect 56856 22326 56866 22583
rect 56880 22326 56890 22583
rect 56904 22326 56914 22583
rect 56928 22326 56938 22583
rect 56952 22326 56962 22583
rect 56976 22326 56986 22583
rect 56509 22313 56770 22323
rect 57000 22299 57010 22583
rect 56509 22289 57010 22299
rect 56509 22265 56783 22275
rect 56509 22241 56735 22251
rect 56520 18829 56530 22216
rect 56544 18829 56554 22216
rect 56568 18829 56578 22216
rect 56592 18829 56602 22216
rect 56616 18829 56626 22216
rect 56664 18829 56674 22216
rect 56688 18829 56698 22216
rect 56712 18829 56722 22216
rect 56808 18829 56818 22264
rect 56832 18829 56842 22264
rect 56856 18829 56866 22264
rect 56880 18829 56890 22264
rect 56904 18802 56914 22264
rect 56509 18792 56914 18802
rect 28464 18168 29903 18178
rect 29832 14584 29842 18143
rect 29856 14584 29866 18143
rect 56520 17413 56530 18767
rect 56544 17413 56554 18767
rect 56568 17413 56578 18767
rect 56592 17413 56602 18767
rect 56616 17413 56626 18767
rect 56664 17413 56674 18767
rect 56688 17413 56698 18767
rect 56712 17386 56722 18767
rect 56509 17376 56722 17386
rect 56520 17149 56530 17351
rect 56544 17149 56554 17351
rect 56568 17149 56578 17351
rect 56592 17149 56602 17351
rect 56616 17149 56626 17351
rect 56664 17149 56674 17351
rect 56688 17149 56698 17351
rect 56808 17122 56818 18767
rect 56509 17112 56818 17122
rect 56520 16813 56530 17087
rect 56544 16813 56554 17087
rect 56568 16813 56578 17087
rect 56592 16813 56602 17087
rect 56616 16813 56626 17087
rect 56664 16813 56674 17087
rect 56688 16786 56698 17087
rect 56509 16776 56698 16786
rect 56520 15013 56530 16751
rect 56544 15013 56554 16751
rect 56568 15013 56578 16751
rect 56592 15013 56602 16751
rect 56616 15013 56626 16751
rect 56664 15013 56674 16751
rect 56832 15013 56842 18767
rect 56856 15013 56866 18767
rect 56880 14986 56890 18767
rect 56509 14976 56890 14986
rect 56520 14605 56530 14951
rect 56544 14605 56554 14951
rect 56568 14605 56578 14951
rect 56592 14698 56602 14951
rect 56616 14725 56626 14951
rect 56664 14725 56674 14951
rect 56592 14688 56735 14698
rect 56832 14674 56842 14951
rect 56856 14677 56866 14951
rect 56928 14677 56938 22264
rect 56688 14664 56842 14674
rect 56616 14629 56626 14663
rect 56688 14626 56698 14664
rect 56952 14650 56962 22264
rect 56976 14653 56986 22264
rect 57024 14653 57034 22583
rect 56712 14640 56962 14650
rect 56712 14629 56722 14640
rect 56640 14616 56698 14626
rect 56640 14602 56650 14616
rect 57048 14626 57058 22583
rect 56773 14616 57058 14626
rect 56605 14592 56650 14602
rect 56701 14592 56975 14602
rect 27504 14568 27562 14578
rect 27552 14560 27562 14568
rect 56653 14568 56927 14578
rect 27504 14544 27527 14554
rect 27504 14434 27514 14544
rect 27552 14550 29903 14560
rect 56509 14554 56542 14560
rect 57024 14557 57034 14591
rect 56509 14550 56855 14554
rect 56520 14544 56855 14550
rect 29880 14526 29903 14536
rect 28392 14461 28402 14519
rect 29832 14461 29842 14519
rect 29856 14461 29866 14519
rect 29880 14461 29890 14526
rect 56492 14530 56503 14537
rect 56492 14520 56735 14530
rect 57072 14530 57082 22583
rect 57096 18466 57106 22583
rect 57144 18493 57154 22583
rect 57408 18493 57418 22583
rect 57456 18493 57466 22583
rect 57504 18493 57514 22608
rect 57096 18456 57561 18466
rect 57480 18445 57490 18456
rect 57144 14533 57154 18431
rect 57408 18274 57418 18431
rect 57456 18418 57466 18431
rect 57456 18408 57561 18418
rect 57480 18301 57490 18383
rect 57504 18301 57514 18383
rect 57408 18264 57561 18274
rect 56797 14520 57082 14530
rect 57480 14506 57490 18239
rect 56509 14496 57490 14506
rect 56736 14482 56746 14496
rect 56736 14472 56807 14482
rect 56869 14472 57143 14482
rect 30333 14434 30343 14447
rect 27504 14424 30343 14434
rect 29808 14400 29831 14410
rect 28392 13957 28402 14399
rect 29808 14338 29818 14400
rect 29917 14400 30284 14410
rect 30357 14410 30367 14447
rect 56640 14434 56650 14471
rect 56664 14437 56674 14471
rect 56688 14437 56698 14471
rect 56712 14437 56722 14471
rect 56736 14448 57023 14458
rect 56736 14437 56746 14448
rect 30312 14400 30367 14410
rect 31872 14424 56650 14434
rect 30312 14386 30322 14400
rect 29832 14376 30322 14386
rect 29832 14365 29842 14376
rect 29904 14338 29914 14351
rect 29808 14328 29914 14338
rect 29832 13930 29842 14303
rect 27461 13920 29842 13930
rect 28392 13117 28402 13895
rect 29856 13117 29866 14303
rect 29880 13090 29890 14303
rect 31872 13093 31882 14424
rect 56832 14424 56855 14434
rect 32016 14400 37607 14410
rect 32016 13093 32026 14400
rect 56832 14410 56842 14424
rect 37621 14400 56842 14410
rect 35376 14376 56663 14386
rect 35376 13093 35386 14376
rect 35520 14352 43727 14362
rect 35520 13093 35530 14352
rect 56712 14362 56722 14375
rect 43741 14352 56722 14362
rect 38904 14328 56543 14338
rect 38904 13093 38914 14328
rect 56736 14338 56746 14375
rect 56760 14341 56770 14375
rect 56653 14328 56746 14338
rect 39048 14304 49703 14314
rect 39048 13093 39058 14304
rect 56784 14314 56794 14375
rect 49717 14304 56794 14314
rect 45960 14280 56759 14290
rect 45960 13093 45970 14280
rect 56808 14290 56818 14375
rect 56784 14280 56818 14290
rect 46104 14256 49847 14266
rect 46104 13093 46114 14256
rect 49861 14256 56591 14266
rect 56677 14256 56687 14266
rect 56784 14266 56794 14280
rect 56712 14256 56794 14266
rect 49488 14232 56567 14242
rect 49488 13093 49498 14232
rect 56712 14242 56722 14256
rect 56605 14232 56722 14242
rect 49632 14208 56663 14218
rect 49632 13093 49642 14208
rect 53016 14184 56639 14194
rect 53016 13093 53026 14184
rect 53160 14160 56615 14170
rect 53160 13093 53170 14160
rect 53208 14136 56591 14146
rect 28368 13080 29890 13090
rect 28368 13066 28378 13080
rect 28344 13056 28378 13066
rect 28344 13014 28354 13056
rect 28405 13056 28450 13066
rect 28392 13014 28402 13055
rect 28440 13014 28450 13056
rect 53208 13066 53218 14136
rect 56520 13810 56530 14111
rect 56808 14002 56818 14280
rect 57504 14029 57514 18239
rect 56808 13992 57561 14002
rect 57504 13954 57514 13967
rect 57504 13944 57561 13954
rect 56520 13800 57561 13810
rect 29869 13056 53218 13066
rect 31872 13014 31882 13031
rect 32016 13014 32026 13031
rect 32064 13014 32074 13056
rect 35376 13014 35386 13031
rect 35520 13014 35530 13031
rect 35568 13014 35578 13056
rect 38904 13014 38914 13031
rect 39048 13014 39058 13031
rect 39096 13014 39106 13056
rect 45960 13014 45970 13031
rect 46104 13014 46114 13031
rect 46152 13014 46162 13056
rect 49488 13014 49498 13031
rect 49632 13014 49642 13031
rect 49680 13014 49690 13056
rect 53016 13014 53026 13031
rect 53160 13014 53170 13031
rect 53208 13014 53218 13056
<< m2contact >>
rect 31799 46007 31813 46021
rect 35327 46007 35341 46021
rect 31871 45983 31885 45997
rect 38903 46007 38917 46021
rect 39047 46007 39061 46021
rect 45959 46007 45973 46021
rect 46103 46007 46117 46021
rect 49463 46007 49477 46021
rect 49607 46007 49621 46021
rect 29975 45959 29989 45973
rect 53135 46007 53149 46021
rect 38903 45959 38917 45973
rect 52943 45959 52957 45973
rect 52967 45959 52981 45973
rect 52991 45959 53005 45973
rect 53015 45959 53029 45973
rect 29927 45935 29941 45949
rect 31799 45935 31813 45949
rect 35327 45935 35341 45949
rect 39047 45935 39061 45949
rect 45959 45935 45973 45949
rect 27503 45071 27517 45085
rect 28367 45071 28381 45085
rect 28463 45071 28477 45085
rect 29927 45887 29941 45901
rect 31871 45911 31885 45925
rect 27503 45023 27517 45037
rect 28367 45023 28381 45037
rect 28463 45023 28477 45037
rect 29975 45863 29989 45877
rect 46103 45911 46117 45925
rect 55487 45935 55501 45949
rect 55535 45959 55549 45973
rect 55295 45911 55309 45925
rect 49463 45887 49477 45901
rect 49607 45887 49621 45901
rect 52943 45887 52957 45901
rect 52967 45887 52981 45901
rect 53015 45863 53029 45877
rect 53135 45863 53149 45877
rect 55511 45887 55525 45901
rect 55559 45887 55573 45901
rect 52991 45839 53005 45853
rect 39047 44567 39061 44581
rect 49463 44567 49477 44581
rect 49607 44567 49621 44581
rect 55295 45815 55309 45829
rect 55487 45839 55501 45853
rect 55511 45839 55525 45853
rect 55535 45839 55549 45853
rect 55559 45839 55573 45853
rect 53015 44567 53029 44581
rect 55295 44567 55309 44581
rect 55463 44567 55477 44581
rect 55487 44567 55501 44581
rect 55511 44567 55525 44581
rect 57503 45263 57517 45277
rect 57503 45215 57517 45229
rect 57479 45143 57493 45157
rect 55559 44591 55573 44605
rect 55583 44567 55597 44581
rect 55607 44543 55621 44557
rect 39047 44519 39061 44533
rect 52991 44519 53005 44533
rect 55343 44519 55357 44533
rect 55463 44519 55477 44533
rect 47543 44495 47557 44509
rect 55535 44495 55549 44509
rect 55655 44471 55669 44485
rect 35327 44447 35341 44461
rect 36575 44447 36589 44461
rect 39047 44447 39061 44461
rect 47351 44447 47365 44461
rect 47711 44447 47725 44461
rect 55679 44447 55693 44461
rect 28463 44279 28477 44293
rect 29927 44279 29941 44293
rect 29951 44279 29965 44293
rect 29975 44279 29989 44293
rect 28463 44231 28477 44245
rect 29975 44231 29989 44245
rect 27527 40655 27541 40669
rect 27527 40607 27541 40621
rect 27503 40583 27517 40597
rect 27503 40535 27517 40549
rect 27503 36167 27517 36181
rect 27551 36191 27565 36205
rect 27527 36119 27541 36133
rect 27503 36071 27517 36085
rect 27527 36071 27541 36085
rect 27551 36071 27565 36085
rect 27503 31751 27517 31765
rect 27551 31775 27565 31789
rect 27503 31703 27517 31717
rect 27551 31727 27565 31741
rect 27503 27359 27517 27373
rect 27527 27359 27541 27373
rect 27551 27359 27565 27373
rect 27503 27311 27517 27325
rect 27527 27311 27541 27325
rect 27551 27311 27565 27325
rect 27503 22895 27517 22909
rect 30479 44183 30493 44197
rect 55751 44423 55765 44437
rect 55775 44423 55789 44437
rect 35327 44399 35341 44413
rect 55463 44399 55477 44413
rect 55487 44399 55501 44413
rect 55799 44399 55813 44413
rect 55487 44375 55501 44389
rect 55559 44375 55573 44389
rect 55823 44375 55837 44389
rect 35543 44351 35557 44365
rect 44831 44351 44845 44365
rect 45551 44351 45565 44365
rect 55559 44351 55573 44365
rect 55583 44351 55597 44365
rect 35543 44303 35557 44317
rect 36575 44303 36589 44317
rect 39047 44303 39061 44317
rect 55751 44327 55765 44341
rect 55775 44327 55789 44341
rect 55799 44327 55813 44341
rect 55631 44279 55645 44293
rect 55703 44279 55717 44293
rect 55727 44279 55741 44293
rect 55751 44279 55765 44293
rect 55775 44279 55789 44293
rect 55847 44303 55861 44317
rect 35327 44255 35341 44269
rect 35351 44255 35365 44269
rect 35543 44255 35557 44269
rect 36575 44255 36589 44269
rect 39047 44255 39061 44269
rect 44567 44255 44581 44269
rect 47615 44255 47629 44269
rect 49607 44255 49621 44269
rect 52991 44255 53005 44269
rect 53015 44255 53029 44269
rect 55823 44255 55837 44269
rect 55871 44255 55885 44269
rect 55583 44231 55597 44245
rect 55799 44231 55813 44245
rect 55895 44231 55909 44245
rect 35327 44207 35341 44221
rect 39047 44207 39061 44221
rect 55919 44207 55933 44221
rect 49463 44183 49477 44197
rect 55295 44159 55309 44173
rect 55343 44183 55357 44197
rect 55823 44183 55837 44197
rect 55847 44183 55861 44197
rect 29927 44135 29941 44149
rect 29951 44135 29965 44149
rect 30599 44135 30613 44149
rect 34151 44135 34165 44149
rect 34391 44135 34405 44149
rect 55295 44135 55309 44149
rect 55463 44135 55477 44149
rect 55487 44135 55501 44149
rect 55511 44135 55525 44149
rect 55535 44135 55549 44149
rect 55559 44135 55573 44149
rect 55583 44135 55597 44149
rect 55607 44135 55621 44149
rect 55631 44135 55645 44149
rect 55655 44135 55669 44149
rect 55679 44135 55693 44149
rect 55703 44135 55717 44149
rect 55727 44135 55741 44149
rect 55751 44135 55765 44149
rect 55775 44135 55789 44149
rect 55799 44135 55813 44149
rect 55823 44135 55837 44149
rect 55871 44159 55885 44173
rect 55895 44159 55909 44173
rect 55919 44159 55933 44173
rect 55463 41351 55477 41365
rect 55487 41351 55501 41365
rect 55511 41351 55525 41365
rect 55535 41351 55549 41365
rect 55559 41351 55573 41365
rect 55583 41351 55597 41365
rect 55607 41351 55621 41365
rect 55631 41351 55645 41365
rect 55655 41351 55669 41365
rect 55679 41351 55693 41365
rect 55703 41351 55717 41365
rect 55727 41351 55741 41365
rect 55751 41351 55765 41365
rect 55775 41351 55789 41365
rect 55799 41351 55813 41365
rect 55823 41351 55837 41365
rect 55847 41351 55861 41365
rect 55871 41351 55885 41365
rect 55895 41351 55909 41365
rect 55919 41351 55933 41365
rect 55919 41303 55933 41317
rect 55463 41231 55477 41245
rect 55487 41231 55501 41245
rect 55511 41231 55525 41245
rect 55535 41231 55549 41245
rect 55559 41231 55573 41245
rect 55583 41231 55597 41245
rect 55607 41231 55621 41245
rect 55631 41231 55645 41245
rect 55655 41231 55669 41245
rect 55679 41231 55693 41245
rect 55703 41231 55717 41245
rect 55727 41231 55741 41245
rect 55751 41231 55765 41245
rect 55775 41231 55789 41245
rect 55799 41231 55813 41245
rect 55823 41231 55837 41245
rect 55847 41231 55861 41245
rect 55871 41231 55885 41245
rect 55895 41231 55909 41245
rect 55463 40175 55477 40189
rect 55487 40175 55501 40189
rect 55511 40175 55525 40189
rect 55535 40175 55549 40189
rect 55559 40175 55573 40189
rect 55583 40175 55597 40189
rect 55607 40175 55621 40189
rect 55631 40175 55645 40189
rect 55655 40175 55669 40189
rect 55679 40175 55693 40189
rect 55703 40175 55717 40189
rect 55727 40175 55741 40189
rect 55751 40175 55765 40189
rect 55775 40175 55789 40189
rect 55799 40175 55813 40189
rect 55823 40175 55837 40189
rect 55847 40175 55861 40189
rect 55871 40175 55885 40189
rect 57479 45095 57493 45109
rect 57479 40847 57493 40861
rect 57503 40847 57517 40861
rect 57455 40823 57469 40837
rect 57503 40799 57517 40813
rect 57455 40775 57469 40789
rect 57479 40775 57493 40789
rect 57431 40679 57445 40693
rect 57455 40679 57469 40693
rect 55871 40127 55885 40141
rect 55463 40055 55477 40069
rect 55487 40055 55501 40069
rect 55511 40055 55525 40069
rect 55535 40055 55549 40069
rect 55559 40055 55573 40069
rect 55583 40055 55597 40069
rect 55607 40055 55621 40069
rect 55631 40055 55645 40069
rect 55655 40055 55669 40069
rect 55679 40055 55693 40069
rect 55703 40055 55717 40069
rect 55727 40055 55741 40069
rect 55751 40055 55765 40069
rect 55775 40055 55789 40069
rect 55799 40055 55813 40069
rect 55823 40055 55837 40069
rect 55847 40055 55861 40069
rect 55463 38999 55477 39013
rect 55487 38999 55501 39013
rect 55511 38999 55525 39013
rect 55535 38999 55549 39013
rect 55559 38999 55573 39013
rect 55583 38999 55597 39013
rect 55607 38999 55621 39013
rect 55631 38999 55645 39013
rect 55655 38999 55669 39013
rect 55679 38999 55693 39013
rect 55703 38999 55717 39013
rect 55727 38999 55741 39013
rect 55751 38999 55765 39013
rect 55775 38999 55789 39013
rect 55799 38999 55813 39013
rect 55823 38999 55837 39013
rect 55823 38951 55837 38965
rect 55463 38879 55477 38893
rect 55487 38879 55501 38893
rect 55511 38879 55525 38893
rect 55535 38879 55549 38893
rect 55559 38879 55573 38893
rect 55583 38879 55597 38893
rect 55607 38879 55621 38893
rect 55631 38879 55645 38893
rect 55655 38879 55669 38893
rect 55679 38879 55693 38893
rect 55703 38879 55717 38893
rect 55727 38879 55741 38893
rect 55751 38879 55765 38893
rect 55775 38879 55789 38893
rect 55799 38879 55813 38893
rect 55463 37823 55477 37837
rect 55487 37823 55501 37837
rect 55511 37823 55525 37837
rect 55535 37823 55549 37837
rect 55559 37823 55573 37837
rect 55583 37823 55597 37837
rect 55607 37823 55621 37837
rect 55631 37823 55645 37837
rect 55655 37823 55669 37837
rect 55679 37823 55693 37837
rect 55703 37823 55717 37837
rect 55727 37823 55741 37837
rect 55751 37823 55765 37837
rect 55775 37823 55789 37837
rect 55775 37775 55789 37789
rect 55463 37703 55477 37717
rect 55487 37703 55501 37717
rect 55511 37703 55525 37717
rect 55535 37703 55549 37717
rect 55559 37703 55573 37717
rect 55583 37703 55597 37717
rect 55607 37703 55621 37717
rect 55631 37703 55645 37717
rect 55655 37703 55669 37717
rect 55679 37703 55693 37717
rect 55703 37703 55717 37717
rect 55727 37703 55741 37717
rect 55751 37703 55765 37717
rect 55463 36647 55477 36661
rect 55487 36647 55501 36661
rect 55511 36647 55525 36661
rect 55535 36647 55549 36661
rect 55559 36647 55573 36661
rect 55583 36647 55597 36661
rect 55607 36647 55621 36661
rect 55631 36647 55645 36661
rect 55655 36647 55669 36661
rect 55679 36647 55693 36661
rect 55703 36647 55717 36661
rect 55727 36647 55741 36661
rect 55751 36647 55765 36661
rect 57503 40655 57517 40669
rect 57431 40631 57445 40645
rect 57455 40631 57469 40645
rect 55463 36527 55477 36541
rect 55487 36527 55501 36541
rect 55511 36527 55525 36541
rect 55535 36527 55549 36541
rect 55559 36527 55573 36541
rect 55583 36527 55597 36541
rect 55607 36527 55621 36541
rect 55631 36527 55645 36541
rect 55655 36527 55669 36541
rect 55679 36527 55693 36541
rect 55703 36527 55717 36541
rect 55727 36527 55741 36541
rect 55751 36527 55765 36541
rect 57503 40607 57517 40621
rect 57479 36383 57493 36397
rect 57503 36383 57517 36397
rect 57479 36335 57493 36349
rect 57503 36287 57517 36301
rect 57455 36215 57469 36229
rect 57479 36215 57493 36229
rect 55463 35471 55477 35485
rect 55487 35471 55501 35485
rect 55511 35471 55525 35485
rect 55535 35471 55549 35485
rect 55559 35471 55573 35485
rect 55583 35471 55597 35485
rect 55607 35471 55621 35485
rect 55631 35471 55645 35485
rect 55655 35471 55669 35485
rect 55679 35471 55693 35485
rect 55703 35471 55717 35485
rect 55727 35471 55741 35485
rect 55751 35471 55765 35485
rect 57455 36167 57469 36181
rect 57479 36167 57493 36181
rect 55463 35351 55477 35365
rect 55487 35351 55501 35365
rect 55511 35351 55525 35365
rect 55535 35351 55549 35365
rect 55559 35351 55573 35365
rect 55583 35351 55597 35365
rect 55607 35351 55621 35365
rect 55631 35351 55645 35365
rect 55655 35351 55669 35365
rect 55679 35351 55693 35365
rect 55703 35351 55717 35365
rect 55727 35351 55741 35365
rect 55751 35351 55765 35365
rect 55463 34295 55477 34309
rect 55487 34295 55501 34309
rect 55511 34295 55525 34309
rect 55535 34295 55549 34309
rect 55559 34295 55573 34309
rect 55583 34295 55597 34309
rect 55607 34295 55621 34309
rect 55631 34295 55645 34309
rect 55655 34295 55669 34309
rect 55679 34295 55693 34309
rect 55703 34295 55717 34309
rect 55727 34295 55741 34309
rect 55751 34295 55765 34309
rect 55463 34175 55477 34189
rect 55487 34175 55501 34189
rect 55511 34175 55525 34189
rect 55535 34175 55549 34189
rect 55559 34175 55573 34189
rect 55583 34175 55597 34189
rect 55607 34175 55621 34189
rect 55631 34175 55645 34189
rect 55655 34175 55669 34189
rect 55679 34175 55693 34189
rect 55703 34175 55717 34189
rect 55727 34175 55741 34189
rect 55751 34175 55765 34189
rect 55463 33119 55477 33133
rect 55487 33119 55501 33133
rect 55511 33119 55525 33133
rect 55535 33119 55549 33133
rect 55559 33119 55573 33133
rect 55583 33119 55597 33133
rect 55607 33119 55621 33133
rect 55631 33119 55645 33133
rect 55655 33119 55669 33133
rect 55679 33119 55693 33133
rect 55703 33119 55717 33133
rect 55727 33119 55741 33133
rect 55607 33071 55621 33085
rect 55751 33071 55765 33085
rect 55775 33071 55789 33085
rect 55463 32999 55477 33013
rect 55487 32999 55501 33013
rect 55511 32999 55525 33013
rect 55535 32999 55549 33013
rect 55559 32999 55573 33013
rect 55583 32999 55597 33013
rect 55463 31943 55477 31957
rect 55631 33023 55645 33037
rect 55655 33023 55669 33037
rect 55679 33023 55693 33037
rect 55703 33023 55717 33037
rect 55727 33023 55741 33037
rect 55751 33023 55765 33037
rect 55775 33023 55789 33037
rect 55511 31967 55525 31981
rect 55535 31967 55549 31981
rect 55559 31967 55573 31981
rect 55583 31967 55597 31981
rect 55607 31967 55621 31981
rect 55631 31967 55645 31981
rect 55655 31967 55669 31981
rect 55679 31967 55693 31981
rect 55703 31967 55717 31981
rect 55727 31967 55741 31981
rect 55751 31967 55765 31981
rect 55775 31967 55789 31981
rect 55799 31967 55813 31981
rect 55511 31919 55525 31933
rect 55487 31871 55501 31885
rect 55823 31895 55837 31909
rect 55463 31823 55477 31837
rect 55487 31823 55501 31837
rect 55535 31847 55549 31861
rect 55559 31847 55573 31861
rect 55583 31847 55597 31861
rect 55607 31847 55621 31861
rect 55631 31847 55645 31861
rect 55655 31847 55669 31861
rect 55679 31847 55693 31861
rect 55703 31847 55717 31861
rect 55727 31847 55741 31861
rect 55751 31847 55765 31861
rect 55775 31847 55789 31861
rect 55799 31847 55813 31861
rect 55823 31847 55837 31861
rect 57527 31751 57541 31765
rect 55487 30791 55501 30805
rect 55511 30791 55525 30805
rect 55535 30791 55549 30805
rect 55559 30791 55573 30805
rect 55583 30791 55597 30805
rect 55607 30791 55621 30805
rect 55631 30791 55645 30805
rect 55655 30791 55669 30805
rect 55679 30791 55693 30805
rect 55703 30791 55717 30805
rect 55727 30791 55741 30805
rect 55751 30791 55765 30805
rect 55775 30791 55789 30805
rect 55799 30791 55813 30805
rect 55823 30791 55837 30805
rect 55487 30743 55501 30757
rect 55511 30743 55525 30757
rect 55535 30743 55549 30757
rect 55559 30743 55573 30757
rect 55583 30743 55597 30757
rect 55607 30743 55621 30757
rect 55631 30743 55645 30757
rect 55655 30743 55669 30757
rect 55679 30743 55693 30757
rect 55703 30743 55717 30757
rect 55727 30743 55741 30757
rect 55463 30695 55477 30709
rect 55487 30695 55501 30709
rect 55511 30695 55525 30709
rect 55535 30695 55549 30709
rect 55559 30695 55573 30709
rect 55583 30695 55597 30709
rect 55607 30695 55621 30709
rect 55631 30695 55645 30709
rect 55655 30695 55669 30709
rect 55679 30695 55693 30709
rect 55703 30695 55717 30709
rect 55847 30719 55861 30733
rect 55463 30647 55477 30661
rect 55487 30647 55501 30661
rect 55511 30647 55525 30661
rect 55535 30647 55549 30661
rect 55559 30647 55573 30661
rect 55583 30647 55597 30661
rect 55607 30647 55621 30661
rect 55631 30647 55645 30661
rect 55655 30647 55669 30661
rect 55679 30647 55693 30661
rect 55703 30647 55717 30661
rect 55463 29591 55477 29605
rect 55487 29591 55501 29605
rect 55511 29591 55525 29605
rect 55751 30671 55765 30685
rect 55775 30671 55789 30685
rect 55799 30671 55813 30685
rect 55823 30671 55837 30685
rect 55847 30671 55861 30685
rect 55559 29615 55573 29629
rect 55583 29615 55597 29629
rect 55607 29615 55621 29629
rect 55631 29615 55645 29629
rect 55655 29615 55669 29629
rect 55679 29615 55693 29629
rect 55703 29615 55717 29629
rect 55727 29615 55741 29629
rect 55751 29615 55765 29629
rect 55775 29615 55789 29629
rect 55799 29615 55813 29629
rect 55823 29615 55837 29629
rect 55847 29615 55861 29629
rect 55871 29615 55885 29629
rect 55559 29567 55573 29581
rect 55583 29567 55597 29581
rect 55607 29567 55621 29581
rect 55631 29567 55645 29581
rect 55535 29519 55549 29533
rect 55559 29519 55573 29533
rect 55583 29519 55597 29533
rect 55607 29519 55621 29533
rect 55895 29543 55909 29557
rect 55463 29471 55477 29485
rect 55487 29471 55501 29485
rect 55511 29471 55525 29485
rect 55535 29471 55549 29485
rect 55559 29471 55573 29485
rect 55583 29471 55597 29485
rect 55607 29471 55621 29485
rect 55655 29495 55669 29509
rect 55679 29495 55693 29509
rect 55703 29495 55717 29509
rect 55727 29495 55741 29509
rect 55751 29495 55765 29509
rect 55775 29495 55789 29509
rect 55799 29495 55813 29509
rect 55823 29495 55837 29509
rect 55847 29495 55861 29509
rect 55871 29495 55885 29509
rect 55895 29495 55909 29509
rect 55463 28415 55477 28429
rect 55487 28415 55501 28429
rect 55511 28415 55525 28429
rect 55535 28415 55549 28429
rect 55559 28415 55573 28429
rect 55583 28415 55597 28429
rect 55607 28415 55621 28429
rect 55631 28415 55645 28429
rect 55655 28415 55669 28429
rect 55703 28439 55717 28453
rect 55727 28439 55741 28453
rect 55751 28439 55765 28453
rect 55775 28439 55789 28453
rect 55799 28439 55813 28453
rect 55823 28439 55837 28453
rect 55847 28439 55861 28453
rect 55871 28439 55885 28453
rect 55895 28439 55909 28453
rect 55919 28439 55933 28453
rect 55583 28367 55597 28381
rect 55679 28367 55693 28381
rect 55943 28367 55957 28381
rect 55463 28295 55477 28309
rect 55487 28295 55501 28309
rect 55511 28295 55525 28309
rect 55535 28295 55549 28309
rect 55559 28295 55573 28309
rect 55607 28319 55621 28333
rect 55631 28319 55645 28333
rect 55655 28319 55669 28333
rect 55679 28319 55693 28333
rect 55703 28319 55717 28333
rect 55727 28319 55741 28333
rect 55751 28319 55765 28333
rect 55775 28319 55789 28333
rect 55799 28319 55813 28333
rect 55823 28319 55837 28333
rect 55847 28319 55861 28333
rect 55871 28319 55885 28333
rect 55895 28319 55909 28333
rect 55919 28319 55933 28333
rect 55943 28319 55957 28333
rect 55463 27239 55477 27253
rect 55487 27239 55501 27253
rect 55511 27239 55525 27253
rect 55535 27239 55549 27253
rect 55559 27239 55573 27253
rect 55583 27239 55597 27253
rect 55607 27239 55621 27253
rect 55631 27239 55645 27253
rect 55655 27239 55669 27253
rect 55679 27239 55693 27253
rect 55703 27239 55717 27253
rect 55727 27239 55741 27253
rect 55751 27239 55765 27253
rect 55775 27239 55789 27253
rect 55799 27239 55813 27253
rect 55823 27239 55837 27253
rect 55871 27263 55885 27277
rect 55895 27263 55909 27277
rect 55919 27263 55933 27277
rect 55943 27263 55957 27277
rect 55967 27263 55981 27277
rect 55583 27191 55597 27205
rect 55847 27191 55861 27205
rect 55991 27191 56005 27205
rect 55463 27119 55477 27133
rect 55487 27119 55501 27133
rect 55511 27119 55525 27133
rect 55535 27119 55549 27133
rect 55559 27119 55573 27133
rect 55463 26063 55477 26077
rect 55487 26063 55501 26077
rect 55511 26063 55525 26077
rect 55535 26063 55549 26077
rect 55607 27143 55621 27157
rect 55631 27143 55645 27157
rect 55655 27143 55669 27157
rect 55679 27143 55693 27157
rect 55703 27143 55717 27157
rect 55727 27143 55741 27157
rect 55751 27143 55765 27157
rect 55775 27143 55789 27157
rect 55799 27143 55813 27157
rect 55823 27143 55837 27157
rect 55847 27143 55861 27157
rect 55871 27143 55885 27157
rect 55895 27143 55909 27157
rect 55919 27143 55933 27157
rect 55943 27143 55957 27157
rect 55967 27143 55981 27157
rect 55991 27143 56005 27157
rect 55583 26087 55597 26101
rect 55607 26087 55621 26101
rect 55631 26087 55645 26101
rect 55655 26087 55669 26101
rect 55679 26087 55693 26101
rect 55703 26087 55717 26101
rect 55727 26087 55741 26101
rect 55751 26087 55765 26101
rect 55775 26087 55789 26101
rect 55799 26087 55813 26101
rect 55823 26087 55837 26101
rect 55847 26087 55861 26101
rect 55871 26087 55885 26101
rect 55895 26087 55909 26101
rect 55919 26087 55933 26101
rect 55943 26087 55957 26101
rect 55967 26087 55981 26101
rect 55991 26087 56005 26101
rect 56015 26087 56029 26101
rect 55535 26015 55549 26029
rect 55559 26015 55573 26029
rect 56039 26015 56053 26029
rect 55463 25943 55477 25957
rect 55487 25943 55501 25957
rect 55511 25943 55525 25957
rect 55559 25967 55573 25981
rect 55583 25967 55597 25981
rect 55607 25967 55621 25981
rect 55631 25967 55645 25981
rect 55655 25967 55669 25981
rect 55679 25967 55693 25981
rect 55703 25967 55717 25981
rect 55727 25967 55741 25981
rect 55751 25967 55765 25981
rect 55775 25967 55789 25981
rect 55799 25967 55813 25981
rect 55823 25967 55837 25981
rect 55847 25967 55861 25981
rect 55871 25967 55885 25981
rect 55895 25967 55909 25981
rect 55919 25967 55933 25981
rect 55943 25967 55957 25981
rect 55967 25967 55981 25981
rect 55991 25967 56005 25981
rect 56015 25967 56029 25981
rect 56039 25967 56053 25981
rect 55463 24887 55477 24901
rect 55487 24887 55501 24901
rect 55511 24887 55525 24901
rect 55535 24887 55549 24901
rect 55559 24887 55573 24901
rect 55583 24887 55597 24901
rect 55607 24887 55621 24901
rect 55631 24887 55645 24901
rect 55655 24887 55669 24901
rect 55679 24887 55693 24901
rect 55727 24911 55741 24925
rect 55751 24911 55765 24925
rect 55775 24911 55789 24925
rect 55799 24911 55813 24925
rect 55823 24911 55837 24925
rect 55847 24911 55861 24925
rect 55871 24911 55885 24925
rect 55895 24911 55909 24925
rect 55919 24911 55933 24925
rect 55943 24911 55957 24925
rect 55967 24911 55981 24925
rect 55991 24911 56005 24925
rect 56015 24911 56029 24925
rect 56039 24911 56053 24925
rect 56063 24911 56077 24925
rect 55727 24863 55741 24877
rect 55751 24863 55765 24877
rect 55775 24863 55789 24877
rect 55799 24863 55813 24877
rect 55823 24863 55837 24877
rect 55847 24863 55861 24877
rect 55871 24863 55885 24877
rect 55895 24863 55909 24877
rect 55919 24863 55933 24877
rect 55943 24863 55957 24877
rect 55967 24863 55981 24877
rect 55991 24863 56005 24877
rect 56015 24863 56029 24877
rect 55703 24815 55717 24829
rect 55727 24815 55741 24829
rect 55751 24815 55765 24829
rect 55775 24815 55789 24829
rect 55799 24815 55813 24829
rect 55823 24815 55837 24829
rect 55847 24815 55861 24829
rect 55871 24815 55885 24829
rect 55895 24815 55909 24829
rect 55919 24815 55933 24829
rect 55943 24815 55957 24829
rect 55967 24815 55981 24829
rect 55991 24815 56005 24829
rect 56087 24839 56101 24853
rect 55463 24767 55477 24781
rect 55487 24767 55501 24781
rect 55511 24767 55525 24781
rect 55535 24767 55549 24781
rect 55559 24767 55573 24781
rect 55583 24767 55597 24781
rect 55607 24767 55621 24781
rect 55631 24767 55645 24781
rect 55655 24767 55669 24781
rect 55679 24767 55693 24781
rect 55703 24767 55717 24781
rect 55727 24767 55741 24781
rect 55751 24767 55765 24781
rect 55775 24767 55789 24781
rect 55799 24767 55813 24781
rect 55823 24767 55837 24781
rect 55847 24767 55861 24781
rect 55871 24767 55885 24781
rect 55895 24767 55909 24781
rect 55919 24767 55933 24781
rect 55943 24767 55957 24781
rect 55967 24767 55981 24781
rect 55991 24767 56005 24781
rect 55463 23711 55477 23725
rect 55487 23711 55501 23725
rect 55511 23711 55525 23725
rect 56039 24791 56053 24805
rect 56063 24791 56077 24805
rect 56087 24791 56101 24805
rect 55559 23735 55573 23749
rect 55583 23735 55597 23749
rect 55607 23735 55621 23749
rect 55631 23735 55645 23749
rect 55655 23735 55669 23749
rect 55679 23735 55693 23749
rect 55703 23735 55717 23749
rect 55727 23735 55741 23749
rect 55751 23735 55765 23749
rect 55775 23735 55789 23749
rect 55799 23735 55813 23749
rect 55823 23735 55837 23749
rect 55847 23735 55861 23749
rect 55871 23735 55885 23749
rect 55895 23735 55909 23749
rect 55919 23735 55933 23749
rect 55943 23735 55957 23749
rect 55967 23735 55981 23749
rect 55991 23735 56005 23749
rect 56015 23735 56029 23749
rect 56039 23735 56053 23749
rect 56063 23735 56077 23749
rect 56087 23735 56101 23749
rect 56111 23735 56125 23749
rect 55559 23687 55573 23701
rect 55583 23687 55597 23701
rect 55607 23687 55621 23701
rect 55631 23687 55645 23701
rect 55655 23687 55669 23701
rect 55679 23687 55693 23701
rect 55703 23687 55717 23701
rect 55727 23687 55741 23701
rect 55535 23639 55549 23653
rect 55559 23639 55573 23653
rect 55583 23639 55597 23653
rect 55607 23639 55621 23653
rect 55631 23639 55645 23653
rect 55655 23639 55669 23653
rect 55679 23639 55693 23653
rect 55703 23639 55717 23653
rect 56135 23663 56149 23677
rect 55463 23591 55477 23605
rect 55487 23591 55501 23605
rect 55511 23591 55525 23605
rect 55535 23591 55549 23605
rect 55559 23591 55573 23605
rect 55583 23591 55597 23605
rect 55607 23591 55621 23605
rect 55631 23591 55645 23605
rect 55655 23591 55669 23605
rect 55679 23591 55693 23605
rect 55703 23591 55717 23605
rect 55751 23615 55765 23629
rect 55775 23615 55789 23629
rect 55799 23615 55813 23629
rect 55823 23615 55837 23629
rect 55847 23615 55861 23629
rect 55871 23615 55885 23629
rect 55895 23615 55909 23629
rect 55919 23615 55933 23629
rect 55943 23615 55957 23629
rect 55967 23615 55981 23629
rect 55991 23615 56005 23629
rect 56015 23615 56029 23629
rect 56039 23615 56053 23629
rect 56063 23615 56077 23629
rect 56087 23615 56101 23629
rect 56111 23615 56125 23629
rect 56135 23615 56149 23629
rect 28463 23519 28477 23533
rect 29879 23519 29893 23533
rect 29903 23519 29917 23533
rect 29927 23519 29941 23533
rect 29951 23519 29965 23533
rect 30479 23519 30493 23533
rect 30666 23519 30680 23533
rect 31943 23519 31957 23533
rect 32135 23519 32149 23533
rect 32927 23519 32941 23533
rect 33479 23519 33493 23533
rect 33695 23519 33709 23533
rect 34439 23519 34453 23533
rect 34607 23519 34621 23533
rect 34991 23519 35005 23533
rect 35183 23519 35197 23533
rect 35399 23519 35413 23533
rect 36143 23519 36157 23533
rect 36311 23519 36325 23533
rect 45719 23519 45733 23533
rect 45911 23519 45925 23533
rect 46151 23519 46165 23533
rect 53855 23519 53869 23533
rect 54791 23519 54805 23533
rect 54887 23519 54901 23533
rect 54959 23519 54973 23533
rect 55295 23519 55309 23533
rect 55463 23519 55477 23533
rect 55487 23519 55501 23533
rect 55511 23519 55525 23533
rect 55535 23519 55549 23533
rect 55559 23519 55573 23533
rect 55583 23519 55597 23533
rect 55607 23519 55621 23533
rect 55631 23519 55645 23533
rect 55655 23519 55669 23533
rect 55679 23519 55693 23533
rect 55703 23519 55717 23533
rect 55727 23519 55741 23533
rect 55751 23519 55765 23533
rect 55775 23519 55789 23533
rect 55799 23519 55813 23533
rect 55823 23519 55837 23533
rect 55847 23519 55861 23533
rect 55871 23519 55885 23533
rect 55895 23519 55909 23533
rect 55919 23519 55933 23533
rect 55943 23519 55957 23533
rect 55967 23519 55981 23533
rect 55991 23519 56005 23533
rect 56015 23519 56029 23533
rect 56039 23519 56053 23533
rect 56063 23519 56077 23533
rect 56087 23519 56101 23533
rect 56111 23519 56125 23533
rect 56135 23519 56149 23533
rect 56159 23519 56173 23533
rect 30503 23495 30517 23509
rect 29975 23471 29989 23485
rect 30199 23471 30213 23485
rect 30594 23471 30608 23485
rect 30618 23471 30632 23485
rect 30642 23471 30656 23485
rect 28463 23423 28477 23437
rect 29879 23423 29893 23437
rect 29903 23423 29917 23437
rect 29927 23423 29941 23437
rect 29951 23423 29965 23437
rect 29975 23423 29989 23437
rect 30009 23423 30023 23437
rect 30055 23423 30069 23437
rect 30101 23423 30115 23437
rect 30147 23423 30161 23437
rect 30199 23423 30213 23437
rect 27551 22919 27565 22933
rect 27503 22847 27517 22861
rect 27551 22871 27565 22885
rect 29855 22751 29869 22765
rect 29831 22727 29845 22741
rect 29783 22703 29797 22717
rect 28463 22679 28477 22693
rect 29735 22679 29749 22693
rect 29975 22679 29989 22693
rect 30032 23389 30046 23403
rect 30078 23389 30092 23403
rect 30124 23389 30138 23403
rect 30170 23389 30184 23403
rect 30199 22871 30213 22885
rect 30503 23399 30517 23413
rect 30240 22847 30254 22861
rect 30311 22847 30325 22861
rect 30335 22847 30349 22861
rect 30359 22847 30373 22861
rect 30383 22823 30397 22837
rect 30407 22799 30421 22813
rect 32351 22823 32365 22837
rect 33167 22823 33181 22837
rect 34007 22847 34021 22861
rect 34031 22823 34045 22837
rect 35207 22895 35221 22909
rect 35639 22895 35653 22909
rect 37247 22919 37261 22933
rect 37967 22895 37981 22909
rect 38447 22871 38461 22885
rect 39335 22847 39349 22861
rect 40223 22823 40237 22837
rect 38423 22799 38437 22813
rect 38447 22799 38461 22813
rect 33983 22775 33997 22789
rect 34031 22775 34045 22789
rect 41303 22775 41317 22789
rect 42143 22775 42157 22789
rect 35183 22751 35197 22765
rect 35207 22751 35221 22765
rect 42167 22751 42181 22765
rect 35615 22727 35629 22741
rect 35639 22727 35653 22741
rect 42983 22727 42997 22741
rect 37223 22703 37237 22717
rect 37247 22703 37261 22717
rect 44567 22703 44581 22717
rect 37943 22679 37957 22693
rect 37967 22679 37981 22693
rect 44605 22679 44619 22693
rect 28391 22655 28405 22669
rect 30167 22655 30181 22669
rect 30199 22655 30213 22669
rect 30240 22655 30254 22669
rect 32327 22655 32341 22669
rect 32351 22655 32365 22669
rect 39311 22655 39325 22669
rect 39335 22655 39349 22669
rect 42959 22655 42973 22669
rect 42983 22655 42997 22669
rect 45383 22655 45397 22669
rect 46199 22703 46213 22717
rect 47663 22679 47677 22693
rect 48572 22655 48586 22669
rect 29879 22631 29893 22645
rect 29975 22631 29989 22645
rect 30284 22631 30298 22645
rect 30311 22631 30325 22645
rect 30335 22631 30349 22645
rect 30359 22631 30373 22645
rect 30383 22631 30397 22645
rect 30407 22631 30421 22645
rect 33959 22631 33973 22645
rect 34007 22631 34021 22645
rect 42119 22631 42133 22645
rect 42143 22631 42157 22645
rect 44543 22631 44557 22645
rect 44567 22631 44581 22645
rect 46175 22631 46189 22645
rect 46199 22631 46213 22645
rect 33167 22607 33181 22621
rect 40223 22607 40237 22621
rect 42167 22607 42181 22621
rect 44605 22607 44619 22621
rect 47663 22607 47677 22621
rect 53879 23495 53893 23509
rect 54815 23495 54829 23509
rect 54599 23471 54613 23485
rect 54623 23471 54637 23485
rect 54743 23471 54757 23485
rect 54767 23471 54781 23485
rect 54839 23471 54853 23485
rect 54815 23447 54829 23461
rect 54767 23423 54781 23437
rect 53879 23399 53893 23413
rect 54623 23399 54637 23413
rect 55463 23471 55477 23485
rect 55487 23471 55501 23485
rect 55511 23471 55525 23485
rect 55535 23471 55549 23485
rect 55559 23471 55573 23485
rect 55583 23471 55597 23485
rect 55607 23471 55621 23485
rect 55631 23471 55645 23485
rect 55655 23471 55669 23485
rect 55679 23471 55693 23485
rect 55703 23471 55717 23485
rect 55727 23471 55741 23485
rect 55751 23471 55765 23485
rect 55775 23471 55789 23485
rect 55799 23471 55813 23485
rect 55823 23471 55837 23485
rect 55847 23471 55861 23485
rect 55871 23471 55885 23485
rect 55895 23471 55909 23485
rect 55919 23471 55933 23485
rect 55943 23471 55957 23485
rect 55967 23471 55981 23485
rect 55991 23471 56005 23485
rect 56015 23471 56029 23485
rect 56039 23471 56053 23485
rect 56063 23471 56077 23485
rect 56087 23471 56101 23485
rect 56111 23471 56125 23485
rect 56135 23471 56149 23485
rect 56159 23471 56173 23485
rect 56183 23327 56197 23341
rect 56519 23303 56533 23317
rect 56543 23279 56557 23293
rect 56567 23255 56581 23269
rect 56591 23231 56605 23245
rect 56615 23207 56629 23221
rect 56639 23183 56653 23197
rect 56663 23159 56677 23173
rect 56687 23135 56701 23149
rect 56711 23111 56725 23125
rect 56735 23087 56749 23101
rect 56759 23063 56773 23077
rect 56783 23039 56797 23053
rect 56807 23015 56821 23029
rect 56831 22991 56845 23005
rect 56855 22967 56869 22981
rect 56879 22943 56893 22957
rect 56903 22919 56917 22933
rect 57503 22919 57517 22933
rect 56927 22871 56941 22885
rect 57503 22871 57517 22885
rect 56951 22847 56965 22861
rect 56975 22823 56989 22837
rect 56999 22799 57013 22813
rect 57023 22775 57037 22789
rect 57503 22775 57517 22789
rect 57047 22727 57061 22741
rect 57503 22727 57517 22741
rect 57071 22703 57085 22717
rect 57095 22703 57109 22717
rect 57143 22679 57157 22693
rect 57407 22655 57421 22669
rect 57455 22631 57469 22645
rect 28391 22583 28405 22597
rect 28463 22583 28477 22597
rect 29735 22583 29749 22597
rect 29783 22583 29797 22597
rect 29831 22583 29845 22597
rect 29855 22583 29869 22597
rect 29879 22583 29893 22597
rect 30309 22583 30323 22597
rect 30333 22583 30347 22597
rect 30357 22583 30371 22597
rect 33143 22583 33157 22597
rect 40199 22583 40213 22597
rect 42143 22583 42157 22597
rect 44576 22583 44590 22597
rect 47639 22583 47653 22597
rect 48596 22583 48610 22597
rect 49391 22583 49405 22597
rect 50975 22583 50989 22597
rect 51671 22583 51685 22597
rect 51815 22583 51829 22597
rect 52607 22583 52621 22597
rect 53423 22583 53437 22597
rect 54215 22583 54229 22597
rect 55031 22583 55045 22597
rect 56519 22583 56533 22597
rect 56543 22583 56557 22597
rect 56567 22583 56581 22597
rect 56591 22583 56605 22597
rect 56615 22583 56629 22597
rect 56639 22583 56653 22597
rect 56663 22583 56677 22597
rect 56687 22583 56701 22597
rect 56711 22583 56725 22597
rect 56735 22583 56749 22597
rect 56759 22583 56773 22597
rect 56783 22583 56797 22597
rect 56807 22583 56821 22597
rect 56831 22583 56845 22597
rect 56855 22583 56869 22597
rect 56879 22583 56893 22597
rect 56903 22583 56917 22597
rect 56927 22583 56941 22597
rect 56951 22583 56965 22597
rect 56975 22583 56989 22597
rect 56999 22583 57013 22597
rect 57023 22583 57037 22597
rect 57047 22583 57061 22597
rect 57071 22583 57085 22597
rect 57095 22583 57109 22597
rect 57143 22583 57157 22597
rect 57407 22583 57421 22597
rect 57455 22583 57469 22597
rect 27503 18431 27517 18445
rect 27503 18383 27517 18397
rect 27527 14591 27541 14605
rect 29783 22415 29797 22429
rect 29831 22415 29845 22429
rect 29855 22415 29869 22429
rect 29879 22415 29893 22429
rect 29903 22383 29917 22397
rect 29783 22359 29797 22373
rect 29903 22359 29917 22373
rect 56519 22360 56533 22374
rect 56543 22360 56557 22374
rect 56567 22360 56581 22374
rect 56591 22360 56605 22374
rect 56615 22360 56629 22374
rect 29831 22335 29845 22349
rect 29855 22335 29869 22349
rect 29879 22335 29893 22349
rect 56495 22336 56509 22350
rect 56663 22336 56677 22350
rect 56687 22336 56701 22350
rect 56711 22336 56725 22350
rect 56735 22336 56749 22350
rect 56495 22312 56509 22326
rect 56783 22312 56797 22326
rect 56807 22312 56821 22326
rect 56831 22312 56845 22326
rect 56855 22312 56869 22326
rect 56879 22312 56893 22326
rect 56903 22312 56917 22326
rect 56927 22312 56941 22326
rect 56951 22312 56965 22326
rect 56975 22312 56989 22326
rect 56495 22288 56509 22302
rect 56495 22264 56509 22278
rect 56783 22264 56797 22278
rect 56807 22264 56821 22278
rect 56831 22264 56845 22278
rect 56855 22264 56869 22278
rect 56879 22264 56893 22278
rect 56903 22264 56917 22278
rect 56927 22264 56941 22278
rect 56951 22264 56965 22278
rect 56975 22264 56989 22278
rect 56495 22240 56509 22254
rect 56735 22240 56749 22254
rect 56519 22216 56533 22230
rect 56543 22216 56557 22230
rect 56567 22216 56581 22230
rect 56591 22216 56605 22230
rect 56615 22216 56629 22230
rect 56663 22216 56677 22230
rect 56687 22216 56701 22230
rect 56711 22216 56725 22230
rect 56519 18815 56533 18829
rect 56543 18815 56557 18829
rect 56567 18815 56581 18829
rect 56591 18815 56605 18829
rect 56615 18815 56629 18829
rect 56663 18815 56677 18829
rect 56687 18815 56701 18829
rect 56711 18815 56725 18829
rect 56807 18815 56821 18829
rect 56831 18815 56845 18829
rect 56855 18815 56869 18829
rect 56879 18815 56893 18829
rect 56495 18791 56509 18805
rect 56519 18767 56533 18781
rect 56543 18767 56557 18781
rect 56567 18767 56581 18781
rect 56591 18767 56605 18781
rect 56615 18767 56629 18781
rect 56663 18767 56677 18781
rect 56687 18767 56701 18781
rect 56711 18767 56725 18781
rect 56807 18767 56821 18781
rect 56831 18767 56845 18781
rect 56855 18767 56869 18781
rect 56879 18767 56893 18781
rect 29831 18191 29845 18205
rect 29855 18191 29869 18205
rect 29879 18191 29893 18205
rect 29903 18167 29917 18181
rect 29831 18143 29845 18157
rect 29855 18143 29869 18157
rect 29879 18143 29893 18157
rect 56519 17399 56533 17413
rect 56543 17399 56557 17413
rect 56567 17399 56581 17413
rect 56591 17399 56605 17413
rect 56615 17399 56629 17413
rect 56663 17399 56677 17413
rect 56687 17399 56701 17413
rect 56495 17375 56509 17389
rect 56519 17351 56533 17365
rect 56543 17351 56557 17365
rect 56567 17351 56581 17365
rect 56591 17351 56605 17365
rect 56615 17351 56629 17365
rect 56663 17351 56677 17365
rect 56687 17351 56701 17365
rect 56519 17135 56533 17149
rect 56543 17135 56557 17149
rect 56567 17135 56581 17149
rect 56591 17135 56605 17149
rect 56615 17135 56629 17149
rect 56663 17135 56677 17149
rect 56687 17135 56701 17149
rect 56495 17111 56509 17125
rect 56519 17087 56533 17101
rect 56543 17087 56557 17101
rect 56567 17087 56581 17101
rect 56591 17087 56605 17101
rect 56615 17087 56629 17101
rect 56663 17087 56677 17101
rect 56687 17087 56701 17101
rect 56519 16799 56533 16813
rect 56543 16799 56557 16813
rect 56567 16799 56581 16813
rect 56591 16799 56605 16813
rect 56615 16799 56629 16813
rect 56663 16799 56677 16813
rect 56495 16775 56509 16789
rect 56519 16751 56533 16765
rect 56543 16751 56557 16765
rect 56567 16751 56581 16765
rect 56591 16751 56605 16765
rect 56615 16751 56629 16765
rect 56663 16751 56677 16765
rect 56519 14999 56533 15013
rect 56543 14999 56557 15013
rect 56567 14999 56581 15013
rect 56591 14999 56605 15013
rect 56615 14999 56629 15013
rect 56663 14999 56677 15013
rect 56831 14999 56845 15013
rect 56855 14999 56869 15013
rect 56495 14975 56509 14989
rect 56519 14951 56533 14965
rect 56543 14951 56557 14965
rect 56567 14951 56581 14965
rect 56591 14951 56605 14965
rect 56615 14951 56629 14965
rect 56663 14951 56677 14965
rect 56831 14951 56845 14965
rect 56855 14951 56869 14965
rect 56615 14711 56629 14725
rect 56663 14711 56677 14725
rect 56735 14687 56749 14701
rect 56615 14663 56629 14677
rect 56615 14615 56629 14629
rect 56855 14663 56869 14677
rect 56927 14663 56941 14677
rect 56975 14639 56989 14653
rect 57023 14639 57037 14653
rect 56519 14591 56533 14605
rect 56543 14591 56557 14605
rect 56567 14591 56581 14605
rect 56591 14591 56605 14605
rect 56711 14615 56725 14629
rect 56759 14615 56773 14629
rect 56687 14591 56701 14605
rect 56975 14591 56989 14605
rect 57023 14591 57037 14605
rect 28391 14570 28405 14584
rect 29831 14570 29845 14584
rect 29855 14570 29869 14584
rect 56639 14567 56653 14581
rect 56927 14567 56941 14581
rect 27527 14543 27541 14557
rect 29903 14549 29917 14563
rect 56495 14549 56509 14563
rect 56855 14543 56869 14557
rect 57023 14543 57037 14557
rect 28391 14519 28405 14533
rect 29831 14519 29845 14533
rect 29855 14519 29869 14533
rect 29903 14525 29917 14539
rect 56478 14525 56492 14539
rect 56735 14519 56749 14533
rect 56783 14519 56797 14533
rect 57143 18479 57157 18493
rect 57407 18479 57421 18493
rect 57455 18479 57469 18493
rect 57503 18479 57517 18493
rect 57143 18431 57157 18445
rect 57407 18431 57421 18445
rect 57455 18431 57469 18445
rect 57479 18431 57493 18445
rect 57479 18383 57493 18397
rect 57503 18383 57517 18397
rect 57479 18287 57493 18301
rect 57503 18287 57517 18301
rect 57479 18239 57493 18253
rect 57503 18239 57517 18253
rect 57143 14519 57157 14533
rect 56495 14495 56509 14509
rect 56639 14471 56653 14485
rect 56663 14471 56677 14485
rect 56687 14471 56701 14485
rect 56711 14471 56725 14485
rect 56807 14471 56821 14485
rect 56855 14471 56869 14485
rect 57143 14471 57157 14485
rect 28391 14447 28405 14461
rect 29831 14447 29845 14461
rect 29855 14447 29869 14461
rect 29879 14447 29893 14461
rect 30332 14447 30346 14461
rect 30356 14447 30370 14461
rect 28391 14399 28405 14413
rect 29831 14399 29845 14413
rect 29903 14399 29917 14413
rect 30284 14399 30298 14413
rect 57023 14447 57037 14461
rect 29831 14351 29845 14365
rect 29903 14351 29917 14365
rect 29831 14303 29845 14317
rect 29855 14303 29869 14317
rect 29879 14303 29893 14317
rect 28391 13943 28405 13957
rect 28391 13895 28405 13909
rect 28391 13103 28405 13117
rect 29855 13103 29869 13117
rect 56663 14423 56677 14437
rect 56687 14423 56701 14437
rect 56711 14423 56725 14437
rect 56735 14423 56749 14437
rect 37607 14399 37621 14413
rect 56855 14423 56869 14437
rect 56663 14375 56677 14389
rect 56711 14375 56725 14389
rect 56735 14375 56749 14389
rect 56759 14375 56773 14389
rect 56783 14375 56797 14389
rect 56807 14375 56821 14389
rect 43727 14351 43741 14365
rect 56543 14327 56557 14341
rect 56639 14327 56653 14341
rect 56759 14327 56773 14341
rect 49703 14303 49717 14317
rect 56759 14279 56773 14293
rect 49847 14255 49861 14269
rect 56591 14255 56605 14269
rect 56663 14255 56677 14269
rect 56687 14255 56701 14269
rect 56567 14231 56581 14245
rect 56591 14231 56605 14245
rect 56663 14207 56677 14221
rect 56639 14183 56653 14197
rect 56615 14159 56629 14173
rect 31871 13079 31885 13093
rect 32015 13079 32029 13093
rect 35375 13079 35389 13093
rect 35519 13079 35533 13093
rect 38903 13079 38917 13093
rect 39047 13079 39061 13093
rect 45959 13079 45973 13093
rect 46103 13079 46117 13093
rect 49487 13079 49501 13093
rect 49631 13079 49645 13093
rect 53015 13079 53029 13093
rect 53159 13079 53173 13093
rect 28391 13055 28405 13069
rect 29855 13055 29869 13069
rect 56591 14135 56605 14149
rect 56519 14111 56533 14125
rect 57503 14015 57517 14029
rect 57503 13967 57517 13981
rect 31871 13031 31885 13045
rect 32015 13031 32029 13045
rect 35375 13031 35389 13045
rect 35519 13031 35533 13045
rect 38903 13031 38917 13045
rect 39047 13031 39061 13045
rect 45959 13031 45973 13045
rect 46103 13031 46117 13045
rect 49487 13031 49501 13045
rect 49631 13031 49645 13045
rect 53015 13031 53029 13045
rect 53159 13031 53173 13045
<< metal2 >>
rect 29928 45901 29940 45935
rect 29976 45877 29988 45959
rect 31800 45949 31812 46007
rect 31872 45925 31884 45983
rect 35328 45949 35340 46007
rect 38904 45973 38916 46007
rect 39048 45949 39060 46007
rect 45960 45949 45972 46007
rect 46104 45925 46116 46007
rect 49464 45901 49476 46007
rect 49608 45901 49620 46007
rect 52944 45901 52956 45959
rect 52968 45901 52980 45959
rect 52992 45853 53004 45959
rect 53016 45877 53028 45959
rect 53136 45877 53148 46007
rect 55296 45829 55308 45911
rect 55488 45853 55500 45935
rect 55512 45853 55524 45887
rect 55536 45853 55548 45959
rect 55560 45853 55572 45887
rect 57504 45229 57516 45263
rect 57480 45109 57492 45143
rect 27504 45037 27516 45071
rect 28368 45037 28380 45071
rect 28464 45037 28476 45071
rect 39048 44533 39060 44567
rect 35328 44413 35340 44447
rect 35544 44317 35556 44351
rect 36576 44317 36588 44447
rect 39048 44317 39060 44447
rect 28464 44245 28476 44279
rect 29928 44149 29940 44279
rect 29952 44149 29964 44279
rect 29976 44245 29988 44279
rect 35328 44221 35340 44255
rect 30480 44124 30492 44183
rect 30595 44135 30599 44149
rect 34147 44135 34151 44149
rect 34387 44135 34391 44149
rect 35352 44148 35364 44255
rect 35544 44148 35556 44255
rect 36576 44148 36588 44255
rect 39048 44221 39060 44255
rect 44568 44148 44580 44255
rect 44832 44148 44844 44351
rect 45552 44148 45564 44351
rect 47352 44148 47364 44447
rect 47544 44148 47556 44495
rect 47616 44148 47628 44255
rect 47712 44148 47724 44447
rect 49464 44197 49476 44567
rect 49608 44269 49620 44567
rect 52992 44269 53004 44519
rect 53016 44269 53028 44567
rect 55296 44173 55308 44567
rect 55464 44533 55476 44567
rect 55344 44197 55356 44519
rect 55488 44413 55500 44567
rect 55464 44149 55476 44399
rect 55488 44149 55500 44375
rect 55512 44149 55524 44567
rect 55536 44149 55548 44495
rect 55560 44389 55572 44591
rect 55584 44365 55596 44567
rect 55560 44149 55572 44351
rect 55584 44149 55596 44231
rect 55608 44149 55620 44543
rect 55632 44149 55644 44279
rect 55656 44149 55668 44471
rect 55680 44149 55692 44447
rect 55752 44341 55764 44423
rect 55776 44341 55788 44423
rect 55800 44341 55812 44399
rect 55704 44149 55716 44279
rect 55728 44149 55740 44279
rect 55752 44149 55764 44279
rect 55776 44149 55788 44279
rect 55824 44269 55836 44375
rect 55800 44149 55812 44231
rect 55848 44197 55860 44303
rect 55824 44149 55836 44183
rect 55872 44173 55884 44255
rect 55896 44173 55908 44231
rect 55920 44173 55932 44207
rect 35347 44136 35364 44148
rect 35539 44136 35556 44148
rect 36573 44136 36588 44148
rect 44564 44136 44580 44148
rect 44828 44136 44844 44148
rect 45548 44136 45564 44148
rect 47347 44136 47364 44148
rect 47539 44136 47556 44148
rect 47611 44136 47628 44148
rect 47707 44136 47724 44148
rect 30595 44124 30607 44135
rect 34147 44124 34159 44135
rect 34387 44124 34399 44135
rect 35347 44124 35359 44136
rect 35539 44124 35551 44136
rect 36573 44124 36585 44136
rect 44564 44124 44576 44136
rect 44828 44124 44840 44136
rect 45548 44124 45560 44136
rect 47347 44124 47359 44136
rect 47539 44124 47551 44136
rect 47611 44124 47623 44136
rect 47707 44124 47719 44136
rect 55296 44124 55308 44135
rect 55464 41245 55476 41351
rect 55488 41245 55500 41351
rect 55512 41245 55524 41351
rect 55536 41245 55548 41351
rect 55560 41245 55572 41351
rect 55584 41245 55596 41351
rect 55608 41245 55620 41351
rect 55632 41245 55644 41351
rect 55656 41245 55668 41351
rect 55680 41245 55692 41351
rect 55704 41245 55716 41351
rect 55728 41245 55740 41351
rect 55752 41245 55764 41351
rect 55776 41245 55788 41351
rect 55800 41245 55812 41351
rect 55824 41245 55836 41351
rect 55848 41245 55860 41351
rect 55872 41245 55884 41351
rect 55896 41245 55908 41351
rect 55920 41317 55932 41351
rect 57456 40789 57468 40823
rect 57480 40789 57492 40847
rect 57504 40813 57516 40847
rect 27528 40621 27540 40655
rect 57432 40645 57444 40679
rect 57456 40645 57468 40679
rect 57504 40621 57516 40655
rect 27504 40549 27516 40583
rect 55464 40069 55476 40175
rect 55488 40069 55500 40175
rect 55512 40069 55524 40175
rect 55536 40069 55548 40175
rect 55560 40069 55572 40175
rect 55584 40069 55596 40175
rect 55608 40069 55620 40175
rect 55632 40069 55644 40175
rect 55656 40069 55668 40175
rect 55680 40069 55692 40175
rect 55704 40069 55716 40175
rect 55728 40069 55740 40175
rect 55752 40069 55764 40175
rect 55776 40069 55788 40175
rect 55800 40069 55812 40175
rect 55824 40069 55836 40175
rect 55848 40069 55860 40175
rect 55872 40141 55884 40175
rect 55464 38893 55476 38999
rect 55488 38893 55500 38999
rect 55512 38893 55524 38999
rect 55536 38893 55548 38999
rect 55560 38893 55572 38999
rect 55584 38893 55596 38999
rect 55608 38893 55620 38999
rect 55632 38893 55644 38999
rect 55656 38893 55668 38999
rect 55680 38893 55692 38999
rect 55704 38893 55716 38999
rect 55728 38893 55740 38999
rect 55752 38893 55764 38999
rect 55776 38893 55788 38999
rect 55800 38893 55812 38999
rect 55824 38965 55836 38999
rect 55464 37717 55476 37823
rect 55488 37717 55500 37823
rect 55512 37717 55524 37823
rect 55536 37717 55548 37823
rect 55560 37717 55572 37823
rect 55584 37717 55596 37823
rect 55608 37717 55620 37823
rect 55632 37717 55644 37823
rect 55656 37717 55668 37823
rect 55680 37717 55692 37823
rect 55704 37717 55716 37823
rect 55728 37717 55740 37823
rect 55752 37717 55764 37823
rect 55776 37789 55788 37823
rect 55464 36541 55476 36647
rect 55488 36541 55500 36647
rect 55512 36541 55524 36647
rect 55536 36541 55548 36647
rect 55560 36541 55572 36647
rect 55584 36541 55596 36647
rect 55608 36541 55620 36647
rect 55632 36541 55644 36647
rect 55656 36541 55668 36647
rect 55680 36541 55692 36647
rect 55704 36541 55716 36647
rect 55728 36541 55740 36647
rect 55752 36541 55764 36647
rect 57480 36349 57492 36383
rect 57504 36301 57516 36383
rect 27504 36085 27516 36167
rect 27528 36085 27540 36119
rect 27552 36085 27564 36191
rect 57456 36181 57468 36215
rect 57480 36181 57492 36215
rect 55464 35365 55476 35471
rect 55488 35365 55500 35471
rect 55512 35365 55524 35471
rect 55536 35365 55548 35471
rect 55560 35365 55572 35471
rect 55584 35365 55596 35471
rect 55608 35365 55620 35471
rect 55632 35365 55644 35471
rect 55656 35365 55668 35471
rect 55680 35365 55692 35471
rect 55704 35365 55716 35471
rect 55728 35365 55740 35471
rect 55752 35365 55764 35471
rect 55464 34189 55476 34295
rect 55488 34189 55500 34295
rect 55512 34189 55524 34295
rect 55536 34189 55548 34295
rect 55560 34189 55572 34295
rect 55584 34189 55596 34295
rect 55608 34189 55620 34295
rect 55632 34189 55644 34295
rect 55656 34189 55668 34295
rect 55680 34189 55692 34295
rect 55704 34189 55716 34295
rect 55728 34189 55740 34295
rect 55752 34189 55764 34295
rect 55464 33013 55476 33119
rect 55488 33013 55500 33119
rect 55512 33013 55524 33119
rect 55536 33013 55548 33119
rect 55560 33013 55572 33119
rect 55584 33013 55596 33119
rect 55608 33085 55620 33119
rect 55632 33037 55644 33119
rect 55656 33037 55668 33119
rect 55680 33037 55692 33119
rect 55704 33037 55716 33119
rect 55728 33037 55740 33119
rect 55752 33037 55764 33071
rect 55776 33037 55788 33071
rect 55464 31837 55476 31943
rect 55512 31933 55524 31967
rect 55488 31837 55500 31871
rect 55536 31861 55548 31967
rect 55560 31861 55572 31967
rect 55584 31861 55596 31967
rect 55608 31861 55620 31967
rect 55632 31861 55644 31967
rect 55656 31861 55668 31967
rect 55680 31861 55692 31967
rect 55704 31861 55716 31967
rect 55728 31861 55740 31967
rect 55752 31861 55764 31967
rect 55776 31861 55788 31967
rect 55800 31861 55812 31967
rect 55824 31861 55836 31895
rect 27504 31717 27516 31751
rect 27552 31741 27564 31775
rect 57541 31752 57561 31764
rect 55488 30757 55500 30791
rect 55512 30757 55524 30791
rect 55536 30757 55548 30791
rect 55560 30757 55572 30791
rect 55584 30757 55596 30791
rect 55608 30757 55620 30791
rect 55632 30757 55644 30791
rect 55656 30757 55668 30791
rect 55680 30757 55692 30791
rect 55704 30757 55716 30791
rect 55728 30757 55740 30791
rect 55464 30661 55476 30695
rect 55488 30661 55500 30695
rect 55512 30661 55524 30695
rect 55536 30661 55548 30695
rect 55560 30661 55572 30695
rect 55584 30661 55596 30695
rect 55608 30661 55620 30695
rect 55632 30661 55644 30695
rect 55656 30661 55668 30695
rect 55680 30661 55692 30695
rect 55704 30661 55716 30695
rect 55752 30685 55764 30791
rect 55776 30685 55788 30791
rect 55800 30685 55812 30791
rect 55824 30685 55836 30791
rect 55848 30685 55860 30719
rect 55464 29485 55476 29591
rect 55488 29485 55500 29591
rect 55512 29485 55524 29591
rect 55560 29581 55572 29615
rect 55584 29581 55596 29615
rect 55608 29581 55620 29615
rect 55632 29581 55644 29615
rect 55536 29485 55548 29519
rect 55560 29485 55572 29519
rect 55584 29485 55596 29519
rect 55608 29485 55620 29519
rect 55656 29509 55668 29615
rect 55680 29509 55692 29615
rect 55704 29509 55716 29615
rect 55728 29509 55740 29615
rect 55752 29509 55764 29615
rect 55776 29509 55788 29615
rect 55800 29509 55812 29615
rect 55824 29509 55836 29615
rect 55848 29509 55860 29615
rect 55872 29509 55884 29615
rect 55896 29509 55908 29543
rect 55464 28309 55476 28415
rect 55488 28309 55500 28415
rect 55512 28309 55524 28415
rect 55536 28309 55548 28415
rect 55560 28309 55572 28415
rect 55584 28381 55596 28415
rect 55608 28333 55620 28415
rect 55632 28333 55644 28415
rect 55656 28333 55668 28415
rect 55680 28333 55692 28367
rect 55704 28333 55716 28439
rect 55728 28333 55740 28439
rect 55752 28333 55764 28439
rect 55776 28333 55788 28439
rect 55800 28333 55812 28439
rect 55824 28333 55836 28439
rect 55848 28333 55860 28439
rect 55872 28333 55884 28439
rect 55896 28333 55908 28439
rect 55920 28333 55932 28439
rect 55944 28333 55956 28367
rect 27504 27325 27516 27359
rect 27528 27325 27540 27359
rect 27552 27325 27564 27359
rect 55464 27133 55476 27239
rect 55488 27133 55500 27239
rect 55512 27133 55524 27239
rect 55536 27133 55548 27239
rect 55560 27133 55572 27239
rect 55584 27205 55596 27239
rect 55608 27157 55620 27239
rect 55632 27157 55644 27239
rect 55656 27157 55668 27239
rect 55680 27157 55692 27239
rect 55704 27157 55716 27239
rect 55728 27157 55740 27239
rect 55752 27157 55764 27239
rect 55776 27157 55788 27239
rect 55800 27157 55812 27239
rect 55824 27157 55836 27239
rect 55848 27157 55860 27191
rect 55872 27157 55884 27263
rect 55896 27157 55908 27263
rect 55920 27157 55932 27263
rect 55944 27157 55956 27263
rect 55968 27157 55980 27263
rect 55992 27157 56004 27191
rect 55464 25957 55476 26063
rect 55488 25957 55500 26063
rect 55512 25957 55524 26063
rect 55536 26029 55548 26063
rect 55560 25981 55572 26015
rect 55584 25981 55596 26087
rect 55608 25981 55620 26087
rect 55632 25981 55644 26087
rect 55656 25981 55668 26087
rect 55680 25981 55692 26087
rect 55704 25981 55716 26087
rect 55728 25981 55740 26087
rect 55752 25981 55764 26087
rect 55776 25981 55788 26087
rect 55800 25981 55812 26087
rect 55824 25981 55836 26087
rect 55848 25981 55860 26087
rect 55872 25981 55884 26087
rect 55896 25981 55908 26087
rect 55920 25981 55932 26087
rect 55944 25981 55956 26087
rect 55968 25981 55980 26087
rect 55992 25981 56004 26087
rect 56016 25981 56028 26087
rect 56040 25981 56052 26015
rect 55464 24781 55476 24887
rect 55488 24781 55500 24887
rect 55512 24781 55524 24887
rect 55536 24781 55548 24887
rect 55560 24781 55572 24887
rect 55584 24781 55596 24887
rect 55608 24781 55620 24887
rect 55632 24781 55644 24887
rect 55656 24781 55668 24887
rect 55680 24781 55692 24887
rect 55728 24877 55740 24911
rect 55752 24877 55764 24911
rect 55776 24877 55788 24911
rect 55800 24877 55812 24911
rect 55824 24877 55836 24911
rect 55848 24877 55860 24911
rect 55872 24877 55884 24911
rect 55896 24877 55908 24911
rect 55920 24877 55932 24911
rect 55944 24877 55956 24911
rect 55968 24877 55980 24911
rect 55992 24877 56004 24911
rect 56016 24877 56028 24911
rect 55704 24781 55716 24815
rect 55728 24781 55740 24815
rect 55752 24781 55764 24815
rect 55776 24781 55788 24815
rect 55800 24781 55812 24815
rect 55824 24781 55836 24815
rect 55848 24781 55860 24815
rect 55872 24781 55884 24815
rect 55896 24781 55908 24815
rect 55920 24781 55932 24815
rect 55944 24781 55956 24815
rect 55968 24781 55980 24815
rect 55992 24781 56004 24815
rect 56040 24805 56052 24911
rect 56064 24805 56076 24911
rect 56088 24805 56100 24839
rect 55464 23605 55476 23711
rect 55488 23605 55500 23711
rect 55512 23605 55524 23711
rect 55560 23701 55572 23735
rect 55584 23701 55596 23735
rect 55608 23701 55620 23735
rect 55632 23701 55644 23735
rect 55656 23701 55668 23735
rect 55680 23701 55692 23735
rect 55704 23701 55716 23735
rect 55728 23701 55740 23735
rect 55536 23605 55548 23639
rect 55560 23605 55572 23639
rect 55584 23605 55596 23639
rect 55608 23605 55620 23639
rect 55632 23605 55644 23639
rect 55656 23605 55668 23639
rect 55680 23605 55692 23639
rect 55704 23605 55716 23639
rect 55752 23629 55764 23735
rect 55776 23629 55788 23735
rect 55800 23629 55812 23735
rect 55824 23629 55836 23735
rect 55848 23629 55860 23735
rect 55872 23629 55884 23735
rect 55896 23629 55908 23735
rect 55920 23629 55932 23735
rect 55944 23629 55956 23735
rect 55968 23629 55980 23735
rect 55992 23629 56004 23735
rect 56016 23629 56028 23735
rect 56040 23629 56052 23735
rect 56064 23629 56076 23735
rect 56088 23629 56100 23735
rect 56112 23629 56124 23735
rect 56136 23629 56148 23663
rect 28464 23437 28476 23519
rect 29880 23437 29892 23519
rect 29904 23437 29916 23519
rect 29928 23437 29940 23519
rect 29952 23437 29964 23519
rect 29976 23437 29988 23471
rect 30010 23437 30022 23552
rect 30033 23403 30045 23552
rect 30056 23437 30068 23552
rect 30079 23403 30091 23552
rect 30102 23437 30114 23552
rect 30125 23403 30137 23552
rect 30148 23437 30160 23552
rect 30171 23403 30183 23552
rect 30480 23533 30492 23552
rect 30200 23437 30212 23471
rect 30504 23413 30516 23495
rect 30595 23485 30607 23552
rect 30619 23485 30631 23552
rect 30643 23485 30655 23552
rect 30667 23533 30679 23552
rect 31939 23533 31951 23552
rect 32131 23533 32143 23552
rect 32923 23533 32935 23552
rect 33475 23533 33487 23552
rect 33691 23533 33703 23552
rect 34435 23533 34447 23552
rect 34603 23533 34615 23552
rect 34987 23533 34999 23552
rect 35179 23533 35191 23552
rect 35395 23533 35407 23552
rect 36139 23533 36151 23552
rect 36307 23533 36319 23552
rect 45715 23533 45727 23552
rect 45907 23533 45919 23552
rect 46147 23533 46159 23552
rect 53851 23533 53863 23552
rect 31939 23519 31943 23533
rect 32131 23519 32135 23533
rect 32923 23519 32927 23533
rect 33475 23519 33479 23533
rect 33691 23519 33695 23533
rect 34435 23519 34439 23533
rect 34603 23519 34607 23533
rect 34987 23519 34991 23533
rect 35179 23519 35183 23533
rect 35395 23519 35399 23533
rect 36139 23519 36143 23533
rect 36307 23519 36311 23533
rect 45715 23519 45719 23533
rect 45907 23519 45911 23533
rect 46147 23519 46151 23533
rect 53851 23519 53855 23533
rect 54595 23532 54607 23552
rect 54739 23532 54751 23552
rect 54787 23533 54799 23552
rect 54595 23520 54612 23532
rect 54739 23520 54756 23532
rect 53880 23413 53892 23495
rect 54600 23485 54612 23520
rect 54744 23485 54756 23520
rect 54787 23519 54791 23533
rect 54835 23532 54847 23552
rect 54883 23533 54895 23552
rect 54955 23533 54967 23552
rect 55296 23533 55308 23552
rect 54835 23520 54852 23532
rect 54624 23413 54636 23471
rect 54768 23437 54780 23471
rect 54816 23461 54828 23495
rect 54840 23485 54852 23520
rect 54883 23519 54887 23533
rect 54955 23519 54959 23533
rect 55464 23485 55476 23519
rect 55488 23485 55500 23519
rect 55512 23485 55524 23519
rect 55536 23485 55548 23519
rect 55560 23485 55572 23519
rect 55584 23485 55596 23519
rect 55608 23485 55620 23519
rect 55632 23485 55644 23519
rect 55656 23485 55668 23519
rect 55680 23485 55692 23519
rect 55704 23485 55716 23519
rect 55728 23485 55740 23519
rect 55752 23485 55764 23519
rect 55776 23485 55788 23519
rect 55800 23485 55812 23519
rect 55824 23485 55836 23519
rect 55848 23485 55860 23519
rect 55872 23485 55884 23519
rect 55896 23485 55908 23519
rect 55920 23485 55932 23519
rect 55944 23485 55956 23519
rect 55968 23485 55980 23519
rect 55992 23485 56004 23519
rect 56016 23485 56028 23519
rect 56040 23485 56052 23519
rect 56064 23485 56076 23519
rect 56088 23485 56100 23519
rect 56112 23485 56124 23519
rect 56136 23485 56148 23519
rect 56160 23485 56172 23519
rect 27504 22861 27516 22895
rect 27552 22885 27564 22919
rect 28392 22597 28404 22655
rect 28464 22597 28476 22679
rect 29736 22597 29748 22679
rect 29784 22597 29796 22703
rect 29832 22597 29844 22727
rect 29856 22597 29868 22751
rect 29976 22645 29988 22679
rect 30200 22669 30212 22871
rect 30241 22669 30253 22847
rect 29880 22597 29892 22631
rect 30168 22551 30180 22655
rect 30312 22645 30324 22847
rect 30336 22645 30348 22847
rect 30360 22645 30372 22847
rect 30384 22645 30396 22823
rect 30408 22645 30420 22799
rect 32352 22669 32364 22823
rect 30285 22551 30297 22631
rect 32328 22596 32340 22655
rect 33168 22621 33180 22823
rect 32325 22584 32340 22596
rect 30309 22551 30321 22583
rect 30333 22551 30345 22583
rect 30357 22551 30369 22583
rect 32325 22551 32337 22584
rect 33141 22583 33143 22597
rect 33960 22596 33972 22631
rect 33957 22584 33972 22596
rect 33984 22596 33996 22775
rect 34008 22645 34020 22847
rect 34032 22789 34044 22823
rect 35208 22765 35220 22895
rect 35184 22596 35196 22751
rect 35640 22741 35652 22895
rect 35616 22596 35628 22727
rect 37248 22717 37260 22919
rect 37224 22596 37236 22703
rect 37968 22693 37980 22895
rect 38448 22813 38460 22871
rect 33984 22584 34005 22596
rect 35184 22584 35205 22596
rect 35616 22584 35637 22596
rect 33141 22551 33153 22583
rect 33957 22551 33969 22584
rect 33993 22551 34005 22584
rect 35193 22551 35205 22584
rect 35625 22551 35637 22584
rect 37221 22584 37236 22596
rect 37944 22596 37956 22679
rect 38424 22596 38436 22799
rect 39336 22669 39348 22847
rect 39312 22596 39324 22655
rect 40224 22621 40236 22823
rect 37944 22584 37965 22596
rect 38424 22584 38445 22596
rect 39312 22584 39333 22596
rect 37221 22551 37233 22584
rect 37953 22551 37965 22584
rect 38433 22551 38445 22584
rect 39321 22551 39333 22584
rect 40213 22583 40221 22597
rect 41304 22596 41316 22775
rect 42144 22645 42156 22775
rect 42120 22596 42132 22631
rect 42168 22621 42180 22751
rect 42984 22669 42996 22727
rect 40209 22551 40221 22583
rect 41301 22584 41316 22596
rect 42117 22584 42132 22596
rect 41301 22551 41313 22584
rect 42117 22551 42129 22584
rect 42157 22583 42165 22597
rect 42960 22596 42972 22655
rect 44568 22645 44580 22703
rect 44544 22596 44556 22631
rect 44606 22621 44618 22679
rect 42960 22584 42981 22596
rect 44544 22584 44565 22596
rect 42153 22551 42165 22583
rect 42969 22551 42981 22584
rect 44553 22551 44565 22584
rect 45384 22596 45396 22655
rect 46200 22645 46212 22703
rect 45381 22584 45396 22596
rect 46176 22596 46188 22631
rect 47664 22621 47676 22679
rect 46176 22584 46197 22596
rect 44577 22551 44589 22583
rect 45381 22551 45393 22584
rect 46185 22551 46197 22584
rect 47653 22583 47661 22597
rect 47649 22551 47661 22583
rect 48573 22551 48585 22655
rect 49405 22583 49413 22597
rect 50989 22583 50997 22597
rect 51685 22583 51693 22597
rect 48597 22551 48609 22583
rect 49401 22551 49413 22583
rect 50985 22551 50997 22583
rect 51681 22551 51693 22583
rect 51813 22583 51815 22597
rect 52621 22583 52629 22597
rect 51813 22551 51825 22583
rect 52617 22551 52629 22583
rect 53421 22583 53423 22597
rect 54229 22583 54237 22597
rect 53421 22551 53433 22583
rect 54225 22551 54237 22583
rect 55029 22583 55031 22597
rect 55029 22551 55041 22583
rect 56184 22551 56196 23327
rect 56520 22597 56532 23303
rect 56544 22597 56556 23279
rect 56568 22597 56580 23255
rect 56592 22597 56604 23231
rect 56616 22597 56628 23207
rect 56640 22597 56652 23183
rect 56664 22597 56676 23159
rect 56688 22597 56700 23135
rect 56712 22597 56724 23111
rect 56736 22597 56748 23087
rect 56760 22597 56772 23063
rect 56784 22597 56796 23039
rect 56808 22597 56820 23015
rect 56832 22597 56844 22991
rect 56856 22597 56868 22967
rect 56880 22597 56892 22943
rect 56904 22597 56916 22919
rect 57504 22885 57516 22919
rect 56928 22597 56940 22871
rect 56952 22597 56964 22847
rect 56976 22597 56988 22823
rect 57000 22597 57012 22799
rect 57024 22597 57036 22775
rect 57504 22741 57516 22775
rect 57048 22597 57060 22727
rect 57072 22597 57084 22703
rect 57096 22597 57108 22703
rect 57144 22597 57156 22679
rect 57408 22597 57420 22655
rect 57456 22597 57468 22631
rect 29784 22373 29796 22415
rect 29832 22349 29844 22415
rect 29856 22349 29868 22415
rect 29880 22349 29892 22415
rect 29917 22384 29946 22396
rect 29917 22360 29946 22372
rect 56467 22336 56495 22348
rect 56467 22312 56495 22324
rect 56467 22288 56495 22300
rect 56467 22264 56495 22276
rect 56467 22240 56495 22252
rect 56520 22230 56532 22360
rect 56544 22230 56556 22360
rect 56568 22230 56580 22360
rect 56592 22230 56604 22360
rect 56616 22230 56628 22360
rect 56664 22230 56676 22336
rect 56688 22230 56700 22336
rect 56712 22230 56724 22336
rect 56736 22254 56748 22336
rect 56784 22278 56796 22312
rect 56808 22278 56820 22312
rect 56832 22278 56844 22312
rect 56856 22278 56868 22312
rect 56880 22278 56892 22312
rect 56904 22278 56916 22312
rect 56928 22278 56940 22312
rect 56952 22278 56964 22312
rect 56976 22278 56988 22312
rect 56467 18791 56495 18803
rect 56520 18781 56532 18815
rect 56544 18781 56556 18815
rect 56568 18781 56580 18815
rect 56592 18781 56604 18815
rect 56616 18781 56628 18815
rect 56664 18781 56676 18815
rect 56688 18781 56700 18815
rect 56712 18781 56724 18815
rect 56808 18781 56820 18815
rect 56832 18781 56844 18815
rect 56856 18781 56868 18815
rect 56880 18781 56892 18815
rect 57144 18445 57156 18479
rect 57408 18445 57420 18479
rect 57456 18445 57468 18479
rect 27504 18397 27516 18431
rect 57480 18397 57492 18431
rect 57504 18397 57516 18479
rect 57480 18253 57492 18287
rect 57504 18253 57516 18287
rect 29832 18157 29844 18191
rect 29856 18157 29868 18191
rect 29880 18157 29892 18191
rect 29917 18167 29946 18179
rect 29893 18155 29916 18156
rect 29893 18144 29946 18155
rect 29904 18143 29946 18144
rect 56467 17375 56495 17387
rect 56520 17365 56532 17399
rect 56544 17365 56556 17399
rect 56568 17365 56580 17399
rect 56592 17365 56604 17399
rect 56616 17365 56628 17399
rect 56664 17365 56676 17399
rect 56688 17365 56700 17399
rect 56467 17111 56495 17123
rect 56520 17101 56532 17135
rect 56544 17101 56556 17135
rect 56568 17101 56580 17135
rect 56592 17101 56604 17135
rect 56616 17101 56628 17135
rect 56664 17101 56676 17135
rect 56688 17101 56700 17135
rect 56467 16775 56495 16787
rect 56520 16765 56532 16799
rect 56544 16765 56556 16799
rect 56568 16765 56580 16799
rect 56592 16765 56604 16799
rect 56616 16765 56628 16799
rect 56664 16765 56676 16799
rect 56467 14989 56509 14994
rect 56467 14982 56495 14989
rect 56520 14965 56532 14999
rect 56544 14965 56556 14999
rect 56568 14965 56580 14999
rect 56592 14965 56604 14999
rect 56616 14965 56628 14999
rect 56664 14965 56676 14999
rect 56832 14965 56844 14999
rect 56856 14965 56868 14999
rect 56616 14677 56628 14711
rect 27528 14557 27540 14591
rect 28392 14533 28404 14570
rect 29832 14533 29844 14570
rect 29856 14533 29868 14570
rect 29917 14550 29946 14562
rect 56467 14550 56495 14562
rect 29917 14526 29946 14538
rect 56467 14526 56478 14538
rect 56467 14509 56507 14514
rect 56467 14502 56495 14509
rect 28392 14413 28404 14447
rect 29832 14413 29844 14447
rect 29832 14317 29844 14351
rect 29856 14317 29868 14447
rect 29880 14317 29892 14447
rect 30285 14413 30297 14491
rect 30333 14461 30345 14491
rect 30357 14461 30369 14491
rect 37617 14460 37629 14491
rect 37608 14448 37629 14460
rect 43725 14460 43737 14491
rect 49713 14460 49725 14491
rect 43725 14448 43740 14460
rect 37608 14413 37620 14448
rect 29904 14365 29916 14399
rect 43728 14365 43740 14448
rect 49704 14448 49725 14460
rect 49845 14460 49857 14491
rect 49845 14448 49860 14460
rect 49704 14317 49716 14448
rect 49848 14269 49860 14448
rect 56520 14125 56532 14591
rect 56544 14341 56556 14591
rect 56568 14245 56580 14591
rect 56592 14269 56604 14591
rect 56592 14149 56604 14231
rect 56616 14173 56628 14615
rect 56640 14485 56652 14567
rect 56664 14485 56676 14711
rect 56688 14485 56700 14591
rect 56712 14485 56724 14615
rect 56736 14533 56748 14687
rect 56664 14389 56676 14423
rect 56640 14197 56652 14327
rect 56688 14269 56700 14423
rect 56712 14389 56724 14423
rect 56736 14389 56748 14423
rect 56760 14389 56772 14615
rect 56856 14557 56868 14663
rect 56928 14581 56940 14663
rect 56976 14605 56988 14639
rect 57024 14605 57036 14639
rect 56784 14389 56796 14519
rect 56808 14389 56820 14471
rect 56856 14437 56868 14471
rect 57024 14461 57036 14543
rect 57144 14485 57156 14519
rect 56760 14293 56772 14327
rect 56664 14221 56676 14255
rect 57504 13981 57516 14015
rect 28392 13909 28404 13943
rect 28392 13069 28404 13103
rect 29856 13069 29868 13103
rect 31872 13045 31884 13079
rect 32016 13045 32028 13079
rect 35376 13045 35388 13079
rect 35520 13045 35532 13079
rect 38904 13045 38916 13079
rect 39048 13045 39060 13079
rect 45960 13045 45972 13079
rect 46104 13045 46116 13079
rect 49488 13045 49500 13079
rect 49632 13045 49644 13079
rect 53016 13045 53028 13079
rect 53160 13045 53172 13079
<< metal4 >>
rect 27627 50850 29187 52410
rect 31153 50850 32713 52410
rect 34679 50850 36239 52410
rect 38205 50850 39765 52410
rect 41731 50850 43291 52410
rect 45257 50850 46817 52410
rect 48783 50850 50343 52410
rect 52309 50850 53869 52410
rect 55835 50850 57395 52410
rect 21089 44398 22649 45958
rect 62373 44398 63933 45958
rect 21089 39926 22649 41486
rect 62373 39926 63933 41486
rect 21089 35454 22649 37014
rect 62373 35454 63933 37014
rect 21089 30982 22649 32542
rect 62373 30982 63933 32542
rect 21089 26510 22649 28070
rect 62373 26510 63933 28070
rect 21089 22038 22649 23598
rect 62373 22038 63933 23598
rect 21089 17566 22649 19126
rect 62373 17566 63933 19126
rect 21089 13094 22649 14654
rect 62373 13094 63933 14654
rect 27627 6642 29187 8202
rect 31153 6642 32713 8202
rect 34679 6642 36239 8202
rect 38205 6642 39765 8202
rect 41731 6642 43291 8202
rect 45257 6642 46817 8202
rect 48783 6642 50343 8202
rect 52309 6642 53869 8202
rect 55835 6642 57395 8202
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 21011 -1 0 52488
box 0 0 6450 6450
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 27547 1 0 46038
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 29267 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 29353 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 29439 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 29525 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 29611 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 29697 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 29783 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 29869 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 29955 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 30041 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 30127 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 30213 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 30299 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 30385 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 30471 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 30557 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 30643 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 30729 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 30815 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 30901 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 0 -1 30987 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 0 -1 31073 1 0 46038
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 32793 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 0 -1 32879 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 0 -1 32965 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 0 -1 33051 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 0 -1 33137 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 0 -1 33223 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 0 -1 33309 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 0 -1 33395 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 0 -1 33481 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 0 -1 33567 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 0 -1 33653 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 0 -1 33739 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 0 -1 33825 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 0 -1 33911 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 33997 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 34083 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 34169 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 34255 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 34341 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 34427 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 34513 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 34599 1 0 46038
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 36319 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 36405 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 36491 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 36577 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 36663 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 36749 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 36835 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 36921 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 37007 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 37093 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 37179 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 37265 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 37351 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 37437 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 37523 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 37609 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 37695 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 37781 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 37867 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 37953 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 38039 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 38125 1 0 46038
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 39845 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 39931 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 40017 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 40103 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 40189 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 40275 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 40361 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 40447 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 40533 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 40619 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 40705 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 40791 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 40877 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 40963 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 41049 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 41135 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 41221 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 41307 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 41393 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 41479 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 41565 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 41651 1 0 46038
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 43371 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 43457 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 43543 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 43629 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 43715 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 0 -1 43801 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 0 -1 43887 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 0 -1 43973 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 0 -1 44059 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 0 -1 44145 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 0 -1 44231 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 0 -1 44317 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 0 -1 44403 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 0 -1 44489 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 0 -1 44575 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 0 -1 44661 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 0 -1 44747 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 0 -1 44833 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 0 -1 44919 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 0 -1 45005 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 0 -1 45091 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 0 -1 45177 1 0 46038
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 46897 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 0 -1 46983 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 0 -1 47069 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 0 -1 47155 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 0 -1 47241 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 0 -1 47327 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 0 -1 47413 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 0 -1 47499 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 0 -1 47585 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 0 -1 47671 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 0 -1 47757 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 0 -1 47843 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 0 -1 47929 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 0 -1 48015 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 0 -1 48101 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 0 -1 48187 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 0 -1 48273 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 0 -1 48359 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 0 -1 48445 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 0 -1 48531 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 0 -1 48617 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 0 -1 48703 1 0 46038
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 50423 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 0 -1 50509 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 0 -1 50595 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 0 -1 50681 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 0 -1 50767 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 0 -1 50853 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 0 -1 50939 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 0 -1 51025 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 0 -1 51111 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 0 -1 51197 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 0 -1 51283 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 0 -1 51369 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 0 -1 51455 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 0 -1 51541 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 0 -1 51627 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 0 -1 51713 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 0 -1 51799 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 0 -1 51885 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 0 -1 51971 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 0 -1 52057 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 0 -1 52143 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 0 -1 52229 1 0 46038
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 53949 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 0 -1 54035 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 0 -1 54121 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 0 -1 54207 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 0 -1 54293 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 0 -1 54379 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 0 -1 54465 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 0 -1 54551 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 0 -1 54637 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 0 -1 54723 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 0 -1 54809 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 0 -1 54895 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 0 -1 54981 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 0 -1 55067 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 0 -1 55153 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 0 -1 55239 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 0 -1 55325 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 0 -1 55411 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 0 -1 55497 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 0 -1 55583 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 0 -1 55669 1 0 46038
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 0 -1 55755 1 0 46038
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 57475 1 0 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 0 -1 57561 1 0 46038
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 64011 0 -1 52488
box 0 0 6450 6450
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 27461 0 -1 46038
box 0 0 6450 1720
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform -1 0 27461 0 -1 44318
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform -1 0 27461 0 -1 44232
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform -1 0 27461 0 -1 44146
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 57561 0 1 44318
box 0 0 6450 1720
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 57561 0 1 44232
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 57561 0 1 44146
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform -1 0 27461 0 -1 44060
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform -1 0 27461 0 -1 43974
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform -1 0 27461 0 -1 43888
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform -1 0 27461 0 -1 43802
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform -1 0 27461 0 -1 43716
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform -1 0 27461 0 -1 43630
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform -1 0 27461 0 -1 43544
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform -1 0 27461 0 -1 43458
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform -1 0 27461 0 -1 43372
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform -1 0 27461 0 -1 43286
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform -1 0 27461 0 -1 43200
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform -1 0 27461 0 -1 43114
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform -1 0 27461 0 -1 43028
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform -1 0 27461 0 -1 42942
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform -1 0 27461 0 -1 42856
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform -1 0 27461 0 -1 42770
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform -1 0 27461 0 -1 42684
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform -1 0 27461 0 -1 42598
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform -1 0 27461 0 -1 42512
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform -1 0 27461 0 -1 42426
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform -1 0 27461 0 -1 42340
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform -1 0 27461 0 -1 42254
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform -1 0 27461 0 -1 42168
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform -1 0 27461 0 -1 42082
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform -1 0 27461 0 -1 41996
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform -1 0 27461 0 -1 41910
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform -1 0 27461 0 -1 41824
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform -1 0 27461 0 -1 41738
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform -1 0 27461 0 -1 41652
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 27461 0 -1 41566
box 0 0 6450 1720
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform -1 0 27461 0 -1 39846
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform -1 0 27461 0 -1 39760
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform -1 0 27461 0 -1 39674
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform -1 0 27461 0 -1 39588
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform -1 0 27461 0 -1 39502
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform -1 0 27461 0 -1 39416
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform -1 0 27461 0 -1 39330
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform -1 0 27461 0 -1 39244
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform -1 0 27461 0 -1 39158
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform -1 0 27461 0 -1 39072
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform -1 0 27461 0 -1 38986
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform -1 0 27461 0 -1 38900
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform -1 0 27461 0 -1 38814
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform -1 0 27461 0 -1 38728
box 0 0 6450 86
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform -1 0 27461 0 -1 38642
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform -1 0 27461 0 -1 38556
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform -1 0 27461 0 -1 38470
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform -1 0 27461 0 -1 38384
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform -1 0 27461 0 -1 38298
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform -1 0 27461 0 -1 38212
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform -1 0 27461 0 -1 38126
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform -1 0 27461 0 -1 38040
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform -1 0 27461 0 -1 37954
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform -1 0 27461 0 -1 37868
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform -1 0 27461 0 -1 37782
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform -1 0 27461 0 -1 37696
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform -1 0 27461 0 -1 37610
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform -1 0 27461 0 -1 37524
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform -1 0 27461 0 -1 37438
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform -1 0 27461 0 -1 37352
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform -1 0 27461 0 -1 37266
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform -1 0 27461 0 -1 37180
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 27461 0 -1 37094
box 0 0 6450 1720
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform -1 0 27461 0 -1 35374
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform -1 0 27461 0 -1 35288
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform -1 0 27461 0 -1 35202
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform -1 0 27461 0 -1 35116
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform -1 0 27461 0 -1 35030
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform -1 0 27461 0 -1 34944
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform -1 0 27461 0 -1 34858
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform -1 0 27461 0 -1 34772
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform -1 0 27461 0 -1 34686
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform -1 0 27461 0 -1 34600
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform -1 0 27461 0 -1 34514
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform -1 0 27461 0 -1 34428
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform -1 0 27461 0 -1 34342
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform -1 0 27461 0 -1 34256
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform -1 0 27461 0 -1 34170
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform -1 0 27461 0 -1 34084
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform -1 0 27461 0 -1 33998
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform -1 0 27461 0 -1 33912
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform -1 0 27461 0 -1 33826
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform -1 0 27461 0 -1 33740
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform -1 0 27461 0 -1 33654
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform -1 0 27461 0 -1 33568
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform -1 0 27461 0 -1 33482
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform -1 0 27461 0 -1 33396
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform -1 0 27461 0 -1 33310
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform -1 0 27461 0 -1 33224
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform -1 0 27461 0 -1 33138
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform -1 0 27461 0 -1 33052
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform -1 0 27461 0 -1 32966
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform -1 0 27461 0 -1 32880
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform -1 0 27461 0 -1 32794
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform -1 0 27461 0 -1 32708
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 27461 0 -1 32622
box 0 0 6450 1720
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform -1 0 27461 0 -1 30902
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform -1 0 27461 0 -1 30816
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform -1 0 27461 0 -1 30730
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform -1 0 27461 0 -1 30644
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform -1 0 27461 0 -1 30558
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform -1 0 27461 0 -1 30472
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform -1 0 27461 0 -1 30386
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform -1 0 27461 0 -1 30300
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform -1 0 27461 0 -1 30214
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform -1 0 27461 0 -1 30128
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform -1 0 27461 0 -1 30042
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform -1 0 27461 0 -1 29956
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform -1 0 27461 0 -1 29870
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform -1 0 27461 0 -1 29784
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform -1 0 27461 0 -1 29698
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform -1 0 27461 0 -1 29612
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform -1 0 27461 0 -1 29526
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform -1 0 27461 0 -1 29440
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform -1 0 27461 0 -1 29354
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform -1 0 27461 0 -1 29268
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform -1 0 27461 0 -1 29182
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform -1 0 27461 0 -1 29096
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform -1 0 27461 0 -1 29010
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform -1 0 27461 0 -1 28924
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform -1 0 27461 0 -1 28838
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform -1 0 27461 0 -1 28752
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform -1 0 27461 0 -1 28666
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform -1 0 27461 0 -1 28580
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform -1 0 27461 0 -1 28494
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform -1 0 27461 0 -1 28408
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform -1 0 27461 0 -1 28322
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform -1 0 27461 0 -1 28236
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 27461 0 -1 28150
box 0 0 6450 1720
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform -1 0 27461 0 -1 26430
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform -1 0 27461 0 -1 26344
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform -1 0 27461 0 -1 26258
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform -1 0 27461 0 -1 26172
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform -1 0 27461 0 -1 26086
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform -1 0 27461 0 -1 26000
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform -1 0 27461 0 -1 25914
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform -1 0 27461 0 -1 25828
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform -1 0 27461 0 -1 25742
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform -1 0 27461 0 -1 25656
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform -1 0 27461 0 -1 25570
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 27461 0 -1 25484
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 27461 0 -1 25398
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 27461 0 -1 25312
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 27461 0 -1 25226
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 27461 0 -1 25140
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 27461 0 -1 25054
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 27461 0 -1 24968
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 27461 0 -1 24882
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 27461 0 -1 24796
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 27461 0 -1 24710
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 27461 0 -1 24624
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 27461 0 -1 24538
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 27461 0 -1 24452
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 27461 0 -1 24366
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 27461 0 -1 24280
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform -1 0 27461 0 -1 24194
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform -1 0 27461 0 -1 24108
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform -1 0 27461 0 -1 24022
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform -1 0 27461 0 -1 23936
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform -1 0 27461 0 -1 23850
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform -1 0 27461 0 -1 23764
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 27461 0 -1 23678
box 0 0 6450 1720
use datapath datapath_0
timestamp 1395690245
transform 1 0 30009 0 1 23552
box 0 0 25408 20572
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 57561 0 1 44060
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 57561 0 1 43974
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 57561 0 1 43888
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 57561 0 1 43802
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 57561 0 1 43716
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 57561 0 1 43630
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 57561 0 1 43544
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 57561 0 1 43458
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 57561 0 1 43372
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 57561 0 1 43286
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 57561 0 1 43200
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 57561 0 1 43114
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 57561 0 1 43028
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 57561 0 1 42942
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 57561 0 1 42856
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 57561 0 1 42770
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 57561 0 1 42684
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 57561 0 1 42598
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 57561 0 1 42512
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 57561 0 1 42426
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 57561 0 1 42340
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 57561 0 1 42254
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 57561 0 1 42168
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 57561 0 1 42082
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 57561 0 1 41996
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 57561 0 1 41910
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 57561 0 1 41824
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 57561 0 1 41738
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 57561 0 1 41652
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 57561 0 1 41566
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 57561 0 1 39846
box 0 0 6450 1720
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 57561 0 1 39760
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 57561 0 1 39674
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 57561 0 1 39588
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 57561 0 1 39502
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 57561 0 1 39416
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 57561 0 1 39330
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 57561 0 1 39244
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 57561 0 1 39158
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 57561 0 1 39072
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 57561 0 1 38986
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 57561 0 1 38900
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 57561 0 1 38814
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 57561 0 1 38728
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 57561 0 1 38642
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 57561 0 1 38556
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 57561 0 1 38470
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 57561 0 1 38384
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 57561 0 1 38298
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 57561 0 1 38212
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 57561 0 1 38126
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 57561 0 1 38040
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 57561 0 1 37954
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 57561 0 1 37868
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 57561 0 1 37782
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 57561 0 1 37696
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 57561 0 1 37610
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 57561 0 1 37524
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 57561 0 1 37438
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 57561 0 1 37352
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 57561 0 1 37266
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 57561 0 1 37180
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 57561 0 1 37094
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 57561 0 1 35374
box 0 0 6450 1720
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 57561 0 1 35288
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 57561 0 1 35202
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 57561 0 1 35116
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 57561 0 1 35030
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 57561 0 1 34944
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 57561 0 1 34858
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 57561 0 1 34772
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 57561 0 1 34686
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 57561 0 1 34600
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 57561 0 1 34514
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 57561 0 1 34428
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 57561 0 1 34342
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 57561 0 1 34256
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 57561 0 1 34170
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 57561 0 1 34084
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 57561 0 1 33998
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 57561 0 1 33912
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 57561 0 1 33826
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 57561 0 1 33740
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 57561 0 1 33654
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 57561 0 1 33568
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 57561 0 1 33482
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 57561 0 1 33396
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 57561 0 1 33310
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 57561 0 1 33224
box 0 0 6450 86
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 57561 0 1 33138
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 57561 0 1 33052
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 57561 0 1 32966
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 57561 0 1 32880
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 57561 0 1 32794
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 57561 0 1 32708
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 57561 0 1 32622
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 57561 0 1 30902
box 0 0 6450 1720
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 57561 0 1 30816
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 57561 0 1 30730
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 57561 0 1 30644
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 57561 0 1 30558
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 57561 0 1 30472
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 57561 0 1 30386
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 57561 0 1 30300
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 57561 0 1 30214
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 57561 0 1 30128
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 57561 0 1 30042
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 57561 0 1 29956
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 57561 0 1 29870
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 57561 0 1 29784
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 57561 0 1 29698
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 57561 0 1 29612
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 57561 0 1 29526
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 57561 0 1 29440
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 57561 0 1 29354
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 57561 0 1 29268
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 57561 0 1 29182
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 57561 0 1 29096
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 57561 0 1 29010
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 57561 0 1 28924
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 57561 0 1 28838
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 57561 0 1 28752
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 57561 0 1 28666
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 57561 0 1 28580
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 57561 0 1 28494
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 57561 0 1 28408
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 57561 0 1 28322
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 57561 0 1 28236
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 57561 0 1 28150
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 57561 0 1 26430
box 0 0 6450 1720
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 57561 0 1 26344
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 57561 0 1 26258
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 57561 0 1 26172
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 57561 0 1 26086
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 57561 0 1 26000
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 57561 0 1 25914
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 57561 0 1 25828
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 57561 0 1 25742
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 57561 0 1 25656
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 57561 0 1 25570
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 57561 0 1 25484
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 57561 0 1 25398
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 57561 0 1 25312
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 57561 0 1 25226
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 57561 0 1 25140
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 57561 0 1 25054
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 57561 0 1 24968
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 57561 0 1 24882
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 57561 0 1 24796
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 57561 0 1 24710
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 57561 0 1 24624
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 57561 0 1 24538
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 57561 0 1 24452
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 57561 0 1 24366
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 57561 0 1 24280
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 57561 0 1 24194
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 57561 0 1 24108
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 57561 0 1 24022
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 57561 0 1 23936
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 57561 0 1 23850
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 57561 0 1 23764
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 57561 0 1 23678
box 0 0 6450 86
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform -1 0 27461 0 -1 21958
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform -1 0 27461 0 -1 21872
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform -1 0 27461 0 -1 21786
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform -1 0 27461 0 -1 21700
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform -1 0 27461 0 -1 21614
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform -1 0 27461 0 -1 21528
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform -1 0 27461 0 -1 21442
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform -1 0 27461 0 -1 21356
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform -1 0 27461 0 -1 21270
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform -1 0 27461 0 -1 21184
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform -1 0 27461 0 -1 21098
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform -1 0 27461 0 -1 21012
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform -1 0 27461 0 -1 20926
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform -1 0 27461 0 -1 20840
box 0 0 6450 86
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform -1 0 27461 0 -1 20754
box 0 0 6450 86
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform -1 0 27461 0 -1 20668
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform -1 0 27461 0 -1 20582
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform -1 0 27461 0 -1 20496
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform -1 0 27461 0 -1 20410
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform -1 0 27461 0 -1 20324
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform -1 0 27461 0 -1 20238
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform -1 0 27461 0 -1 20152
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform -1 0 27461 0 -1 20066
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform -1 0 27461 0 -1 19980
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform -1 0 27461 0 -1 19894
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform -1 0 27461 0 -1 19808
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform -1 0 27461 0 -1 19722
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform -1 0 27461 0 -1 19636
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform -1 0 27461 0 -1 19550
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform -1 0 27461 0 -1 19464
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform -1 0 27461 0 -1 19378
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform -1 0 27461 0 -1 19292
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 27461 0 -1 19206
box 0 0 6450 1720
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform -1 0 27461 0 -1 17486
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform -1 0 27461 0 -1 17400
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform -1 0 27461 0 -1 17314
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform -1 0 27461 0 -1 17228
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform -1 0 27461 0 -1 17142
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform -1 0 27461 0 -1 17056
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform -1 0 27461 0 -1 16970
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform -1 0 27461 0 -1 16884
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform -1 0 27461 0 -1 16798
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform -1 0 27461 0 -1 16712
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform -1 0 27461 0 -1 16626
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform -1 0 27461 0 -1 16540
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform -1 0 27461 0 -1 16454
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform -1 0 27461 0 -1 16368
box 0 0 6450 86
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform -1 0 27461 0 -1 16282
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform -1 0 27461 0 -1 16196
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform -1 0 27461 0 -1 16110
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform -1 0 27461 0 -1 16024
box 0 0 6450 86
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform -1 0 27461 0 -1 15938
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform -1 0 27461 0 -1 15852
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform -1 0 27461 0 -1 15766
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform -1 0 27461 0 -1 15680
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform -1 0 27461 0 -1 15594
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform -1 0 27461 0 -1 15508
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform -1 0 27461 0 -1 15422
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform -1 0 27461 0 -1 15336
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform -1 0 27461 0 -1 15250
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform -1 0 27461 0 -1 15164
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform -1 0 27461 0 -1 15078
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform -1 0 27461 0 -1 14992
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform -1 0 27461 0 -1 14906
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform -1 0 27461 0 -1 14820
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 27461 0 -1 14734
box 0 0 6450 1720
use control control_0
timestamp 1395929462
transform 1 0 29946 0 1 14491
box 0 0 26521 8060
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 57561 0 1 21958
box 0 0 6450 1720
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 57561 0 1 21872
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 57561 0 1 21786
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 57561 0 1 21700
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 57561 0 1 21614
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 57561 0 1 21528
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 57561 0 1 21442
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 1 0 57561 0 1 21356
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 1 0 57561 0 1 21270
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 1 0 57561 0 1 21184
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 1 0 57561 0 1 21098
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 1 0 57561 0 1 21012
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 1 0 57561 0 1 20926
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 1 0 57561 0 1 20840
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 1 0 57561 0 1 20754
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 1 0 57561 0 1 20668
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 1 0 57561 0 1 20582
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 1 0 57561 0 1 20496
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 1 0 57561 0 1 20410
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 1 0 57561 0 1 20324
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 1 0 57561 0 1 20238
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 1 0 57561 0 1 20152
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 1 0 57561 0 1 20066
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 1 0 57561 0 1 19980
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 1 0 57561 0 1 19894
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 1 0 57561 0 1 19808
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 1 0 57561 0 1 19722
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 1 0 57561 0 1 19636
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 1 0 57561 0 1 19550
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 1 0 57561 0 1 19464
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 1 0 57561 0 1 19378
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 1 0 57561 0 1 19292
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 1 0 57561 0 1 19206
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 57561 0 1 17486
box 0 0 6450 1720
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 1 0 57561 0 1 17400
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 1 0 57561 0 1 17314
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 1 0 57561 0 1 17228
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 1 0 57561 0 1 17142
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 1 0 57561 0 1 17056
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 1 0 57561 0 1 16970
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 1 0 57561 0 1 16884
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 1 0 57561 0 1 16798
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 1 0 57561 0 1 16712
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 1 0 57561 0 1 16626
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 1 0 57561 0 1 16540
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 1 0 57561 0 1 16454
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 1 0 57561 0 1 16368
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 1 0 57561 0 1 16282
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 1 0 57561 0 1 16196
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 1 0 57561 0 1 16110
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 1 0 57561 0 1 16024
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 1 0 57561 0 1 15938
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 1 0 57561 0 1 15852
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 1 0 57561 0 1 15766
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 1 0 57561 0 1 15680
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 1 0 57561 0 1 15594
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 1 0 57561 0 1 15508
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 1 0 57561 0 1 15422
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 1 0 57561 0 1 15336
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 1 0 57561 0 1 15250
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 1 0 57561 0 1 15164
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 1 0 57561 0 1 15078
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 1 0 57561 0 1 14992
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 1 0 57561 0 1 14906
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 1 0 57561 0 1 14820
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 1 0 57561 0 1 14734
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 57561 0 1 13014
box 0 0 6450 1720
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 21011 0 1 6564
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 27461 -1 0 13014
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 27547 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 29267 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 29353 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 29439 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 29525 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 29611 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 29697 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 29783 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 29869 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 29955 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 30041 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 30127 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 30213 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 30299 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 30385 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 30471 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 30557 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 30643 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 30729 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 30815 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 30901 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 30987 -1 0 13014
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 31073 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 32793 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 32879 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 32965 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 33051 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 33137 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 33223 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 33309 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 33395 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 33481 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 33567 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 33653 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 33739 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 33825 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 33911 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 33997 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 34083 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 34169 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 34255 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 34341 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 34427 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 34513 -1 0 13014
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 34599 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 36319 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 36405 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 36491 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 36577 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 36663 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 36749 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 36835 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 36921 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 37007 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 37093 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 37179 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 37265 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 37351 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 37437 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 37523 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 37609 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 37695 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 37781 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 37867 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 37953 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 38039 -1 0 13014
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 38125 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 39845 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 39931 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 40017 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 40103 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 40189 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 40275 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 40361 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 40447 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 40533 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 40619 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 40705 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 40791 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 40877 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 40963 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 41049 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 41135 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 41221 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 41307 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 41393 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 41479 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 41565 -1 0 13014
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 41651 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 43371 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 43457 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 43543 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 43629 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 43715 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 43801 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 43887 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 43973 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 44059 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 44145 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 44231 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 44317 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 44403 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 44489 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 44575 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 44661 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 44747 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 44833 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 44919 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 45005 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 45091 -1 0 13014
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 45177 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 46897 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 46983 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 47069 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 47155 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 47241 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 47327 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 47413 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 47499 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 47585 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 47671 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 47757 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 47843 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 47929 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 48015 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 48101 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 48187 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 48273 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 48359 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 48445 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 48531 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 48617 -1 0 13014
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 48703 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 50423 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 50509 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 50595 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 50681 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 50767 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 50853 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 50939 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 51025 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 51111 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 51197 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 51283 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 51369 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 51455 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 51541 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 51627 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 51713 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 51799 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 51885 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 51971 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 52057 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 52143 -1 0 13014
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 52229 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 53949 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 54035 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 54121 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 54207 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 54293 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 54379 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 54465 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 54551 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 54637 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 54723 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 54809 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 54895 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 54981 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 55067 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 55153 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 55239 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 55325 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 55411 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 55497 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 55583 -1 0 13014
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 55669 -1 0 13014
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 55755 -1 0 13014
box 0 0 6450 1720
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 57475 -1 0 13014
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 64011 1 0 6564
box 0 0 6450 6450
<< labels >>
rlabel metal4 27627 6642 29187 8202 0 nIRQ
rlabel metal4 31153 6642 32713 8202 0 Data[0]
rlabel metal4 34679 6642 36239 8202 0 Data[1]
rlabel metal4 38205 6642 39765 8202 0 Data[2]
rlabel metal4 41731 6642 43291 8202 0 vdde!
rlabel metal4 45257 6642 46817 8202 0 Data[3]
rlabel metal4 48783 6642 50343 8202 0 Data[4]
rlabel metal4 52309 6642 53869 8202 0 Data[5]
rlabel metal4 55835 6642 57395 8202 0 gnde!
rlabel metal4 62373 13094 63933 14654 0 Data[6]
rlabel metal4 62373 17566 63933 19126 0 Data[7]
rlabel metal4 62373 22038 63933 23598 0 Data[8]
rlabel metal4 62373 26510 63933 28070 0 gnde!
rlabel metal4 62373 30982 63933 32542 0 GND!
rlabel metal4 62373 35454 63933 37014 0 Data[9]
rlabel metal4 62373 39926 63933 41486 0 Data[10]
rlabel metal4 62373 44398 63933 45958 0 Data[11]
rlabel metal4 55835 50850 57395 52410 0 vdde!
rlabel metal4 52309 50850 53869 52410 0 Data[12]
rlabel metal4 48783 50850 50343 52410 0 Data[13]
rlabel metal4 45257 50850 46817 52410 0 Data[14]
rlabel metal4 41731 50850 43291 52410 0 gnde!
rlabel metal4 38205 50850 39765 52410 0 Data[15]
rlabel metal4 34679 50850 36239 52410 0 ALE
rlabel metal4 31153 50850 32713 52410 0 nME
rlabel metal4 27627 50850 29187 52410 0 nWait
rlabel metal4 21089 44398 22649 45958 0 nOE
rlabel metal4 21089 39926 22649 41486 0 RnW
rlabel metal4 21089 35454 22649 37014 0 SDO
rlabel metal4 21089 30982 22649 32542 0 Vdd!
rlabel metal4 21089 26510 22649 28070 0 SDI
rlabel metal4 21089 22038 22649 23598 0 Test
rlabel metal4 21089 17566 22649 19126 0 Clock
rlabel metal4 21089 13094 22649 14654 0 nReset
<< end >>
