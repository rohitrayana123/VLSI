magic
tech c035u
timestamp 1398680265
<< pohmic >>
rect 0 16160 37 16170
<< metal1 >>
rect 0 17069 37 17079
rect 0 17047 37 17057
rect 0 17024 37 17034
rect 0 16933 37 16943
rect 0 16911 37 16921
rect 0 16888 37 16898
rect 0 16866 37 16876
rect 0 16843 37 16853
rect 0 16805 37 16830
rect 0 16160 37 16185
rect 0 16137 37 16147
rect 0 16114 37 16124
rect 0 16091 37 16101
rect 0 15901 60 15911
rect 9253 15877 9289 15887
rect 9253 15855 9289 15865
rect 0 15806 37 15816
rect 0 15783 37 15793
rect 0 15745 37 15770
rect 0 15100 37 15125
rect 0 15077 37 15087
rect 0 15054 37 15064
rect 0 15031 37 15041
rect 0 14901 60 14911
rect 9253 14877 9289 14887
rect 9253 14855 9289 14865
rect 0 14806 37 14816
rect 0 14783 37 14793
rect 0 14745 37 14770
rect 0 14100 37 14125
rect 0 14077 37 14087
rect 0 14054 37 14064
rect 0 14031 37 14041
rect 0 13901 60 13911
rect 9253 13877 9289 13887
rect 9253 13855 9289 13865
rect 0 13806 37 13816
rect 0 13783 37 13793
rect 0 13745 37 13770
rect 0 13100 37 13125
rect 0 13077 37 13087
rect 0 13054 37 13064
rect 0 13031 37 13041
rect 0 12901 60 12911
rect 9253 12877 9289 12887
rect 9253 12855 9289 12865
rect 0 12806 37 12816
rect 0 12783 37 12793
rect 0 12745 37 12770
rect 0 12100 37 12125
rect 0 12077 37 12087
rect 0 12054 37 12064
rect 0 12031 37 12041
rect 0 11901 60 11911
rect 9253 11877 9289 11887
rect 9253 11855 9289 11865
rect 0 11806 37 11816
rect 0 11783 37 11793
rect 0 11745 37 11770
rect 0 11100 37 11125
rect 0 11077 37 11087
rect 0 11054 37 11064
rect 0 11031 37 11041
rect 0 10901 60 10911
rect 9253 10877 9289 10887
rect 9253 10855 9289 10865
rect 0 10806 37 10816
rect 0 10783 37 10793
rect 0 10745 37 10770
rect 0 10100 37 10125
rect 0 10077 37 10087
rect 0 10054 37 10064
rect 0 10031 37 10041
rect 0 9901 60 9911
rect 9253 9877 9289 9887
rect 9253 9855 9289 9865
rect 0 9806 37 9816
rect 0 9783 37 9793
rect 0 9745 37 9770
rect 0 9100 37 9125
rect 0 9077 37 9087
rect 0 9054 37 9064
rect 0 9031 37 9041
rect 0 8901 60 8911
rect 9253 8877 9289 8887
rect 9253 8855 9289 8865
rect 0 8806 37 8816
rect 0 8783 37 8793
rect 0 8745 37 8770
rect 0 8100 37 8125
rect 0 8077 37 8087
rect 0 8054 37 8064
rect 0 8031 37 8041
rect 0 7901 60 7911
rect 9253 7877 9289 7887
rect 9253 7855 9289 7865
rect 0 7806 37 7816
rect 0 7783 37 7793
rect 0 7745 37 7770
rect 0 7100 37 7125
rect 0 7077 37 7087
rect 0 7054 37 7064
rect 0 7031 37 7041
rect 0 6901 60 6911
rect 9253 6877 9289 6887
rect 9253 6855 9289 6865
rect 0 6806 37 6816
rect 0 6783 37 6793
rect 0 6745 37 6770
rect 0 6100 37 6125
rect 0 6077 37 6087
rect 0 6054 37 6064
rect 0 6031 37 6041
rect 0 5901 60 5911
rect 9253 5877 9289 5887
rect 9253 5855 9289 5865
rect 0 5806 37 5816
rect 0 5783 37 5793
rect 0 5745 37 5770
rect 0 5100 37 5125
rect 0 5077 37 5087
rect 0 5054 37 5064
rect 0 5031 37 5041
rect 0 4901 60 4911
rect 9253 4877 9289 4887
rect 9253 4855 9289 4865
rect 0 4806 37 4816
rect 0 4783 37 4793
rect 0 4745 37 4770
rect 0 4100 37 4125
rect 0 4077 37 4087
rect 0 4054 37 4064
rect 0 4031 37 4041
rect 0 3901 60 3911
rect 9253 3877 9289 3887
rect 9253 3855 9289 3865
rect 0 3806 37 3816
rect 0 3783 37 3793
rect 0 3745 37 3770
rect 0 3100 37 3125
rect 0 3077 37 3087
rect 0 3054 37 3064
rect 0 3031 37 3041
rect 0 2901 60 2911
rect 9253 2877 9289 2887
rect 9253 2855 9289 2865
rect 0 2806 37 2816
rect 0 2783 37 2793
rect 0 2745 37 2770
rect 0 2100 37 2125
rect 0 2077 37 2087
rect 0 2054 37 2064
rect 0 2031 37 2041
rect 0 1901 60 1911
rect 9253 1877 9289 1887
rect 9253 1855 9289 1865
rect 0 1806 37 1816
rect 0 1783 37 1793
rect 0 1745 37 1770
rect 0 1100 37 1125
rect 0 1077 37 1087
rect 0 1054 37 1064
rect 0 1031 37 1041
rect 0 901 60 911
rect 9253 877 9289 887
rect 9253 855 9289 865
rect 0 806 37 816
rect 0 783 37 793
rect 0 745 37 770
rect 0 100 37 125
rect 0 77 37 87
rect 0 54 37 64
rect 0 31 37 41
<< m2contact >>
rect 60 15901 74 15915
rect 60 14901 74 14915
rect 60 13901 74 13915
rect 60 12901 74 12915
rect 60 11901 74 11915
rect 60 10901 74 10915
rect 60 9901 74 9915
rect 60 8901 74 8915
rect 60 7901 74 7915
rect 60 6901 74 6915
rect 60 5901 74 5915
rect 60 4901 74 4915
rect 60 3901 74 3915
rect 60 2901 74 2915
rect 60 1901 74 1915
rect 60 901 74 915
<< metal2 >>
rect 159 17110 171 17130
rect 713 17110 725 17130
rect 737 17110 749 17130
rect 761 17110 773 17130
rect 61 15894 73 15901
rect 109 15894 121 15979
rect 853 15894 865 15979
rect 1069 15894 1081 15979
rect 1261 15894 1273 15979
rect 2005 15894 2017 15979
rect 2221 15894 2233 15979
rect 2413 15894 2425 15979
rect 3157 15894 3169 15979
rect 3373 15894 3385 15979
rect 3565 15894 3577 15979
rect 4309 15894 4321 15979
rect 4525 15894 4537 15979
rect 4717 15894 4729 15979
rect 5461 15894 5473 15979
rect 5677 15894 5689 15979
rect 5869 15894 5881 15979
rect 6613 15894 6625 15979
rect 6829 15894 6841 15979
rect 7021 15894 7033 15979
rect 7765 15894 7777 15979
rect 7981 15894 7993 15979
rect 8173 15894 8185 15979
rect 8917 15894 8929 15979
rect 9133 15894 9145 15979
rect 61 14894 73 14901
rect 109 14894 121 15000
rect 853 14894 865 15000
rect 1069 14894 1081 15000
rect 1261 14894 1273 15000
rect 2005 14894 2017 15000
rect 2221 14894 2233 15000
rect 2413 14894 2425 15000
rect 3157 14894 3169 15000
rect 3373 14894 3385 15000
rect 3565 14894 3577 15000
rect 4309 14894 4321 15000
rect 4525 14894 4537 15000
rect 4717 14894 4729 15000
rect 5461 14894 5473 15000
rect 5677 14894 5689 15000
rect 5869 14894 5881 15000
rect 6613 14894 6625 15000
rect 6829 14894 6841 15000
rect 7021 14894 7033 15000
rect 7765 14894 7777 15000
rect 7981 14894 7993 15000
rect 8173 14894 8185 15000
rect 8917 14894 8929 15000
rect 9133 14894 9145 15000
rect 61 13894 73 13901
rect 109 13894 121 14000
rect 853 13894 865 14000
rect 1069 13894 1081 14000
rect 1261 13894 1273 14000
rect 2005 13894 2017 14000
rect 2221 13894 2233 14000
rect 2413 13894 2425 14000
rect 3157 13894 3169 14000
rect 3373 13894 3385 14000
rect 3565 13894 3577 14000
rect 4309 13894 4321 14000
rect 4525 13894 4537 14000
rect 4717 13894 4729 14000
rect 5461 13894 5473 14000
rect 5677 13894 5689 14000
rect 5869 13894 5881 14000
rect 6613 13894 6625 14000
rect 6829 13894 6841 14000
rect 7021 13894 7033 14000
rect 7765 13894 7777 14000
rect 7981 13894 7993 14000
rect 8173 13894 8185 14000
rect 8917 13894 8929 14000
rect 9133 13894 9145 14000
rect 61 12894 73 12901
rect 109 12894 121 13000
rect 853 12894 865 13000
rect 1069 12894 1081 13000
rect 1261 12894 1273 13000
rect 2005 12894 2017 13000
rect 2221 12894 2233 13000
rect 2413 12894 2425 13000
rect 3157 12894 3169 13000
rect 3373 12894 3385 13000
rect 3565 12894 3577 13000
rect 4309 12894 4321 13000
rect 4525 12894 4537 13000
rect 4717 12894 4729 13000
rect 5461 12894 5473 13000
rect 5677 12894 5689 13000
rect 5869 12894 5881 13000
rect 6613 12894 6625 13000
rect 6829 12894 6841 13000
rect 7021 12894 7033 13000
rect 7765 12894 7777 13000
rect 7981 12894 7993 13000
rect 8173 12894 8185 13000
rect 8917 12894 8929 13000
rect 9133 12894 9145 13000
rect 61 11894 73 11901
rect 109 11894 121 12000
rect 853 11894 865 12000
rect 1069 11894 1081 12000
rect 1261 11894 1273 12000
rect 2005 11894 2017 12000
rect 2221 11894 2233 12000
rect 2413 11894 2425 12000
rect 3157 11894 3169 12000
rect 3373 11894 3385 12000
rect 3565 11894 3577 12000
rect 4309 11894 4321 12000
rect 4525 11894 4537 12000
rect 4717 11894 4729 12000
rect 5461 11894 5473 12000
rect 5677 11894 5689 12000
rect 5869 11894 5881 12000
rect 6613 11894 6625 12000
rect 6829 11894 6841 12000
rect 7021 11894 7033 12000
rect 7765 11894 7777 12000
rect 7981 11894 7993 12000
rect 8173 11894 8185 12000
rect 8917 11894 8929 12000
rect 9133 11894 9145 12000
rect 61 10894 73 10901
rect 109 10894 121 11000
rect 853 10894 865 11000
rect 1069 10894 1081 11000
rect 1261 10894 1273 11000
rect 2005 10894 2017 11000
rect 2221 10894 2233 11000
rect 2413 10894 2425 11000
rect 3157 10894 3169 11000
rect 3373 10894 3385 11000
rect 3565 10894 3577 11000
rect 4309 10894 4321 11000
rect 4525 10894 4537 11000
rect 4717 10894 4729 11000
rect 5461 10894 5473 11000
rect 5677 10894 5689 11000
rect 5869 10894 5881 11000
rect 6613 10894 6625 11000
rect 6829 10894 6841 11000
rect 7021 10894 7033 11000
rect 7765 10894 7777 11000
rect 7981 10894 7993 11000
rect 8173 10894 8185 11000
rect 8917 10894 8929 11000
rect 9133 10894 9145 11000
rect 61 9894 73 9901
rect 109 9894 121 10000
rect 853 9894 865 10000
rect 1069 9894 1081 10000
rect 1261 9894 1273 10000
rect 2005 9894 2017 10000
rect 2221 9894 2233 10000
rect 2413 9894 2425 10000
rect 3157 9894 3169 10000
rect 3373 9894 3385 10000
rect 3565 9894 3577 10000
rect 4309 9894 4321 10000
rect 4525 9894 4537 10000
rect 4717 9894 4729 10000
rect 5461 9894 5473 10000
rect 5677 9894 5689 10000
rect 5869 9894 5881 10000
rect 6613 9894 6625 10000
rect 6829 9894 6841 10000
rect 7021 9894 7033 10000
rect 7765 9894 7777 10000
rect 7981 9894 7993 10000
rect 8173 9894 8185 10000
rect 8917 9894 8929 10000
rect 9133 9894 9145 10000
rect 61 8894 73 8901
rect 109 8894 121 9000
rect 853 8894 865 9000
rect 1069 8894 1081 9000
rect 1261 8894 1273 9000
rect 2005 8894 2017 9000
rect 2221 8894 2233 9000
rect 2413 8894 2425 9000
rect 3157 8894 3169 9000
rect 3373 8894 3385 9000
rect 3565 8894 3577 9000
rect 4309 8894 4321 9000
rect 4525 8894 4537 9000
rect 4717 8894 4729 9000
rect 5461 8894 5473 9000
rect 5677 8894 5689 9000
rect 5869 8894 5881 9000
rect 6613 8894 6625 9000
rect 6829 8894 6841 9000
rect 7021 8894 7033 9000
rect 7765 8894 7777 9000
rect 7981 8894 7993 9000
rect 8173 8894 8185 9000
rect 8917 8894 8929 9000
rect 9133 8894 9145 9000
rect 61 7894 73 7901
rect 109 7894 121 8000
rect 853 7894 865 8000
rect 1069 7894 1081 8000
rect 1261 7894 1273 8000
rect 2005 7894 2017 8000
rect 2221 7894 2233 8000
rect 2413 7894 2425 8000
rect 3157 7894 3169 8000
rect 3373 7894 3385 8000
rect 3565 7894 3577 8000
rect 4309 7894 4321 8000
rect 4525 7894 4537 8000
rect 4717 7894 4729 8000
rect 5461 7894 5473 8000
rect 5677 7894 5689 8000
rect 5869 7894 5881 8000
rect 6613 7894 6625 8000
rect 6829 7894 6841 8000
rect 7021 7894 7033 8000
rect 7765 7894 7777 8000
rect 7981 7894 7993 8000
rect 8173 7894 8185 8000
rect 8917 7894 8929 8000
rect 9133 7894 9145 8000
rect 61 6894 73 6901
rect 109 6894 121 7000
rect 853 6894 865 7000
rect 1069 6894 1081 7000
rect 1261 6894 1273 7000
rect 2005 6894 2017 7000
rect 2221 6894 2233 7000
rect 2413 6894 2425 7000
rect 3157 6894 3169 7000
rect 3373 6894 3385 7000
rect 3565 6894 3577 7000
rect 4309 6894 4321 7000
rect 4525 6894 4537 7000
rect 4717 6894 4729 7000
rect 5461 6894 5473 7000
rect 5677 6894 5689 7000
rect 5869 6894 5881 7000
rect 6613 6894 6625 7000
rect 6829 6894 6841 7000
rect 7021 6894 7033 7000
rect 7765 6894 7777 7000
rect 7981 6894 7993 7000
rect 8173 6894 8185 7000
rect 8917 6894 8929 7000
rect 9133 6894 9145 7000
rect 61 5894 73 5901
rect 109 5894 121 6000
rect 853 5894 865 6000
rect 1069 5894 1081 6000
rect 1261 5894 1273 6000
rect 2005 5894 2017 6000
rect 2221 5894 2233 6000
rect 2413 5894 2425 6000
rect 3157 5894 3169 6000
rect 3373 5894 3385 6000
rect 3565 5894 3577 6000
rect 4309 5894 4321 6000
rect 4525 5894 4537 6000
rect 4717 5894 4729 6000
rect 5461 5894 5473 6000
rect 5677 5894 5689 6000
rect 5869 5894 5881 6000
rect 6613 5894 6625 6000
rect 6829 5894 6841 6000
rect 7021 5894 7033 6000
rect 7765 5894 7777 6000
rect 7981 5894 7993 6000
rect 8173 5894 8185 6000
rect 8917 5894 8929 6000
rect 9133 5894 9145 6000
rect 61 4894 73 4901
rect 109 4894 121 5000
rect 853 4894 865 5000
rect 1069 4894 1081 5000
rect 1261 4894 1273 5000
rect 2005 4894 2017 5000
rect 2221 4894 2233 5000
rect 2413 4894 2425 5000
rect 3157 4894 3169 5000
rect 3373 4894 3385 5000
rect 3565 4894 3577 5000
rect 4309 4894 4321 5000
rect 4525 4894 4537 5000
rect 4717 4894 4729 5000
rect 5461 4894 5473 5000
rect 5677 4894 5689 5000
rect 5869 4894 5881 5000
rect 6613 4894 6625 5000
rect 6829 4894 6841 5000
rect 7021 4894 7033 5000
rect 7765 4894 7777 5000
rect 7981 4894 7993 5000
rect 8173 4894 8185 5000
rect 8917 4894 8929 5000
rect 9133 4894 9145 5000
rect 61 3894 73 3901
rect 109 3894 121 4000
rect 853 3894 865 4000
rect 1069 3894 1081 4000
rect 1261 3894 1273 4000
rect 2005 3894 2017 4000
rect 2221 3894 2233 4000
rect 2413 3894 2425 4000
rect 3157 3894 3169 4000
rect 3373 3894 3385 4000
rect 3565 3894 3577 4000
rect 4309 3894 4321 4000
rect 4525 3894 4537 4000
rect 4717 3894 4729 4000
rect 5461 3894 5473 4000
rect 5677 3894 5689 4000
rect 5869 3894 5881 4000
rect 6613 3894 6625 4000
rect 6829 3894 6841 4000
rect 7021 3894 7033 4000
rect 7765 3894 7777 4000
rect 7981 3894 7993 4000
rect 8173 3894 8185 4000
rect 8917 3894 8929 4000
rect 9133 3894 9145 4000
rect 61 2894 73 2901
rect 109 2894 121 3000
rect 853 2894 865 3000
rect 1069 2894 1081 3000
rect 1261 2894 1273 3000
rect 2005 2894 2017 3000
rect 2221 2894 2233 3000
rect 2413 2894 2425 3000
rect 3157 2894 3169 3000
rect 3373 2894 3385 3000
rect 3565 2894 3577 3000
rect 4309 2894 4321 3000
rect 4525 2894 4537 3000
rect 4717 2894 4729 3000
rect 5461 2894 5473 3000
rect 5677 2894 5689 3000
rect 5869 2894 5881 3000
rect 6613 2894 6625 3000
rect 6829 2894 6841 3000
rect 7021 2894 7033 3000
rect 7765 2894 7777 3000
rect 7981 2894 7993 3000
rect 8173 2894 8185 3000
rect 8917 2894 8929 3000
rect 9133 2894 9145 3000
rect 61 1894 73 1901
rect 109 1894 121 2000
rect 853 1894 865 2000
rect 1069 1894 1081 2000
rect 1261 1894 1273 2000
rect 2005 1894 2017 2000
rect 2221 1894 2233 2000
rect 2413 1894 2425 2000
rect 3157 1894 3169 2000
rect 3373 1894 3385 2000
rect 3565 1894 3577 2000
rect 4309 1894 4321 2000
rect 4525 1894 4537 2000
rect 4717 1894 4729 2000
rect 5461 1894 5473 2000
rect 5677 1894 5689 2000
rect 5869 1894 5881 2000
rect 6613 1894 6625 2000
rect 6829 1894 6841 2000
rect 7021 1894 7033 2000
rect 7765 1894 7777 2000
rect 7981 1894 7993 2000
rect 8173 1894 8185 2000
rect 8917 1894 8929 2000
rect 9133 1894 9145 2000
rect 61 894 73 901
rect 109 894 121 1000
rect 853 894 865 1000
rect 1069 894 1081 1000
rect 1261 894 1273 1000
rect 2005 894 2017 1000
rect 2221 894 2233 1000
rect 2413 894 2425 1000
rect 3157 894 3169 1000
rect 3373 894 3385 1000
rect 3565 894 3577 1000
rect 4309 894 4321 1000
rect 4525 894 4537 1000
rect 4717 894 4729 1000
rect 5461 894 5473 1000
rect 5677 894 5689 1000
rect 5869 894 5881 1000
rect 6613 894 6625 1000
rect 6829 894 6841 1000
rect 7021 894 7033 1000
rect 7765 894 7777 1000
rect 7981 894 7993 1000
rect 8173 894 8185 1000
rect 8917 894 8929 1000
rect 9133 894 9145 1000
use regBlock_decoder regBlock_decoder_0
timestamp 1397223953
transform 1 0 37 0 1 15979
box 0 0 9217 1131
use regBlock_slice regBlock_slice_0
array 0 0 80 0 15 1000
timestamp 1396393625
transform 1 0 37 0 1 -21
box 0 21 9216 915
<< labels >>
rlabel metal1 0 31 0 41 3 nReset
rlabel metal1 0 1031 0 1041 3 nReset
rlabel metal1 0 2031 0 2041 3 nReset
rlabel metal1 0 3031 0 3041 3 nReset
rlabel metal1 0 4031 0 4041 3 nReset
rlabel metal1 0 5031 0 5041 3 nReset
rlabel metal1 0 6031 0 6041 3 nReset
rlabel metal1 0 7031 0 7041 3 nReset
rlabel metal1 0 8031 0 8041 3 nReset
rlabel metal1 0 9031 0 9041 3 nReset
rlabel metal1 0 10031 0 10041 3 nReset
rlabel metal1 0 11031 0 11041 3 nReset
rlabel metal1 0 12031 0 12041 3 nReset
rlabel metal1 0 13031 0 13041 3 nReset
rlabel metal1 0 14031 0 14041 3 nReset
rlabel metal1 0 15031 0 15041 3 nReset
rlabel metal1 0 54 0 64 3 Test
rlabel metal1 0 1054 0 1064 3 Test
rlabel metal1 0 2054 0 2064 3 Test
rlabel metal1 0 3054 0 3064 3 Test
rlabel metal1 0 4054 0 4064 3 Test
rlabel metal1 0 5054 0 5064 3 Test
rlabel metal1 0 6054 0 6064 3 Test
rlabel metal1 0 7054 0 7064 3 Test
rlabel metal1 0 8054 0 8064 3 Test
rlabel metal1 0 9054 0 9064 3 Test
rlabel metal1 0 10054 0 10064 3 Test
rlabel metal1 0 11054 0 11064 3 Test
rlabel metal1 0 12054 0 12064 3 Test
rlabel metal1 0 13054 0 13064 3 Test
rlabel metal1 0 14054 0 14064 3 Test
rlabel metal1 0 15054 0 15064 3 Test
rlabel metal1 0 77 0 87 3 Clock
rlabel metal1 0 1077 0 1087 3 Clock
rlabel metal1 0 2077 0 2087 3 Clock
rlabel metal1 0 3077 0 3087 3 Clock
rlabel metal1 0 4077 0 4087 3 Clock
rlabel metal1 0 5077 0 5087 3 Clock
rlabel metal1 0 6077 0 6087 3 Clock
rlabel metal1 0 7077 0 7087 3 Clock
rlabel metal1 0 8077 0 8087 3 Clock
rlabel metal1 0 9077 0 9087 3 Clock
rlabel metal1 0 10077 0 10087 3 Clock
rlabel metal1 0 11077 0 11087 3 Clock
rlabel metal1 0 12077 0 12087 3 Clock
rlabel metal1 0 13077 0 13087 3 Clock
rlabel metal1 0 14077 0 14087 3 Clock
rlabel metal1 0 15077 0 15087 3 Clock
rlabel metal1 0 100 0 125 3 GND!
rlabel metal1 0 1100 0 1125 3 GND!
rlabel metal1 0 2100 0 2125 3 GND!
rlabel metal1 0 3100 0 3125 3 GND!
rlabel metal1 0 4100 0 4125 3 GND!
rlabel metal1 0 5100 0 5125 3 GND!
rlabel metal1 0 6100 0 6125 3 GND!
rlabel metal1 0 7100 0 7125 3 GND!
rlabel metal1 0 8100 0 8125 3 GND!
rlabel metal1 0 9100 0 9125 3 GND!
rlabel metal1 0 10100 0 10125 3 GND!
rlabel metal1 0 11100 0 11125 3 GND!
rlabel metal1 0 12100 0 12125 3 GND!
rlabel metal1 0 13100 0 13125 3 GND!
rlabel metal1 0 14100 0 14125 3 GND!
rlabel metal1 0 15100 0 15125 3 GND!
rlabel metal1 0 745 0 770 3 Vdd!
rlabel metal1 0 1745 0 1770 3 Vdd!
rlabel metal1 0 2745 0 2770 3 Vdd!
rlabel metal1 0 3745 0 3770 3 Vdd!
rlabel metal1 0 4745 0 4770 3 Vdd!
rlabel metal1 0 5745 0 5770 3 Vdd!
rlabel metal1 0 6745 0 6770 3 Vdd!
rlabel metal1 0 7745 0 7770 3 Vdd!
rlabel metal1 0 8745 0 8770 3 Vdd!
rlabel metal1 0 9745 0 9770 3 Vdd!
rlabel metal1 0 10745 0 10770 3 Vdd!
rlabel metal1 0 11745 0 11770 3 Vdd!
rlabel metal1 0 12745 0 12770 3 Vdd!
rlabel metal1 0 13745 0 13770 3 Vdd!
rlabel metal1 0 14745 0 14770 3 Vdd!
rlabel metal1 0 15745 0 15770 3 Vdd!
rlabel metal1 0 783 0 793 3 SDI
rlabel metal1 0 1783 0 1793 3 SDI
rlabel metal1 0 2783 0 2793 3 SDI
rlabel metal1 0 3783 0 3793 3 SDI
rlabel metal1 0 4783 0 4793 3 SDI
rlabel metal1 0 5783 0 5793 3 SDI
rlabel metal1 0 6783 0 6793 3 SDI
rlabel metal1 0 7783 0 7793 3 SDI
rlabel metal1 0 8783 0 8793 3 SDI
rlabel metal1 0 9783 0 9793 3 SDI
rlabel metal1 0 10783 0 10793 3 SDI
rlabel metal1 0 11783 0 11793 3 SDI
rlabel metal1 0 12783 0 12793 3 SDI
rlabel metal1 0 13783 0 13793 3 SDI
rlabel metal1 0 14783 0 14793 3 SDI
rlabel metal1 0 15783 0 15793 3 SDI
rlabel metal1 0 806 0 816 3 ScanReturn
rlabel metal1 0 1806 0 1816 3 ScanReturn
rlabel metal1 0 2806 0 2816 3 ScanReturn
rlabel metal1 0 3806 0 3816 3 ScanReturn
rlabel metal1 0 4806 0 4816 3 ScanReturn
rlabel metal1 0 5806 0 5816 3 ScanReturn
rlabel metal1 0 6806 0 6816 3 ScanReturn
rlabel metal1 0 7806 0 7816 3 ScanReturn
rlabel metal1 0 8806 0 8816 3 ScanReturn
rlabel metal1 0 9806 0 9816 3 ScanReturn
rlabel metal1 0 10806 0 10816 3 ScanReturn
rlabel metal1 0 11806 0 11816 3 ScanReturn
rlabel metal1 0 12806 0 12816 3 ScanReturn
rlabel metal1 0 13806 0 13816 3 ScanReturn
rlabel metal1 0 14806 0 14816 3 ScanReturn
rlabel metal1 0 15806 0 15816 3 ScanReturn
rlabel metal1 0 901 0 911 3 WData[0]
rlabel metal1 0 1901 0 1911 3 WData[1]
rlabel metal1 0 2901 0 2911 3 WData[2]
rlabel metal1 0 3901 0 3911 3 WData[3]
rlabel metal1 0 4901 0 4911 3 WData[4]
rlabel metal1 0 5901 0 5911 3 WData[5]
rlabel metal1 0 6901 0 6911 3 WData[6]
rlabel metal1 0 7901 0 7911 3 WData[7]
rlabel metal1 0 8901 0 8911 3 WData[8]
rlabel metal1 0 9901 0 9911 3 WData[9]
rlabel metal1 0 10901 0 10911 3 WData[10]
rlabel metal1 0 11901 0 11911 3 WData[11]
rlabel metal1 0 12901 0 12911 3 WData[12]
rlabel metal1 0 13901 0 13911 3 WData[13]
rlabel metal1 0 14901 0 14911 3 WData[14]
rlabel metal1 0 15901 0 15911 3 WData[15]
rlabel metal1 9289 855 9289 865 7 Rd2[0]
rlabel metal1 9289 1855 9289 1865 7 Rd2[1]
rlabel metal1 9289 2855 9289 2865 7 Rd2[2]
rlabel metal1 9289 3855 9289 3865 7 Rd2[3]
rlabel metal1 9289 4855 9289 4865 7 Rd2[4]
rlabel metal1 9289 5855 9289 5865 7 Rd2[5]
rlabel metal1 9289 6855 9289 6865 7 Rd2[6]
rlabel metal1 9289 7855 9289 7865 7 Rd2[7]
rlabel metal1 9289 8855 9289 8865 7 Rd2[8]
rlabel metal1 9289 9855 9289 9865 7 Rd2[9]
rlabel metal1 9289 10855 9289 10865 7 Rd2[10]
rlabel metal1 9289 11855 9289 11865 7 Rd2[11]
rlabel metal1 9289 12855 9289 12865 7 Rd2[12]
rlabel metal1 9289 13855 9289 13865 7 Rd2[13]
rlabel metal1 9289 14855 9289 14865 7 Rd2[14]
rlabel metal1 9289 15855 9289 15865 7 Rd2[15]
rlabel metal1 9289 877 9289 887 7 Rd1[0]
rlabel metal1 9289 1877 9289 1887 7 Rd1[1]
rlabel metal1 9289 2877 9289 2887 7 Rd1[2]
rlabel metal1 9289 3877 9289 3887 7 Rd1[3]
rlabel metal1 9289 4877 9289 4887 7 Rd1[4]
rlabel metal1 9289 5877 9289 5887 7 Rd1[5]
rlabel metal1 9289 6877 9289 6887 7 Rd1[6]
rlabel metal1 9289 7877 9289 7887 7 Rd1[7]
rlabel metal1 9289 8877 9289 8887 7 Rd1[8]
rlabel metal1 9289 9877 9289 9887 7 Rd1[9]
rlabel metal1 9289 10877 9289 10887 7 Rd1[10]
rlabel metal1 9289 11877 9289 11887 7 Rd1[11]
rlabel metal1 9289 12877 9289 12887 7 Rd1[12]
rlabel metal1 9289 13877 9289 13887 7 Rd1[13]
rlabel metal1 9289 14877 9289 14887 7 Rd1[14]
rlabel metal1 9289 15877 9289 15887 7 Rd1[15]
rlabel metal1 0 16888 0 16898 3 Rs1[0]
rlabel metal1 0 16911 0 16921 3 Rs1[1]
rlabel metal1 0 16933 0 16943 3 Rs1[2]
rlabel metal1 0 17024 0 17034 3 Rw[0]
rlabel metal1 0 17047 0 17057 3 Rw[1]
rlabel metal1 0 17069 0 17079 3 Rw[2]
rlabel metal2 159 17130 171 17130 5 We
rlabel metal2 713 17130 725 17130 5 Rs2[0]
rlabel metal2 737 17130 749 17130 5 Rs2[1]
rlabel metal2 761 17130 773 17130 5 Rs2[2]
rlabel metal1 0 16091 0 16101 3 nReset
rlabel metal1 0 16114 0 16124 3 Test
rlabel metal1 0 16137 0 16147 3 Clock
rlabel metal1 0 16160 0 16185 3 GND!
rlabel metal1 0 16843 0 16853 3 Scan
rlabel metal1 0 16866 0 16876 3 ScanReturn
rlabel metal1 0 16805 0 16830 3 Vdd!
<< end >>
