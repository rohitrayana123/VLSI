../../../../c035u/Datapath/datapath.sv