magic
tech c035u
timestamp 1396965088
<< nwell >>
rect 25803 1395 26450 1793
<< pwell >>
rect 25803 994 26450 1395
<< pohmic >>
rect 25803 1070 25808 1080
rect 26443 1070 26450 1080
<< nohmic >>
rect 25803 1730 25808 1740
rect 26443 1730 26450 1740
<< psubstratetap >>
rect 25808 1070 26443 1086
<< nsubstratetap >>
rect 25808 1724 26443 1740
<< metal1 >>
rect 6808 8564 6826 8578
rect 9028 8566 19130 8576
rect 22156 8566 24866 8576
rect 5320 8542 16454 8552
rect 21340 8542 24338 8552
rect 5056 8518 13190 8528
rect 18892 8518 23210 8528
rect 23788 8518 26186 8528
rect 2320 8492 2338 8506
rect 3232 8494 4298 8504
rect 4888 8494 10610 8504
rect 13168 8494 13946 8504
rect 15628 8494 18962 8504
rect 19708 8494 25466 8504
rect 84 8470 10922 8480
rect 11200 8468 11218 8482
rect 12496 8470 23798 8480
rect 84 8446 10370 8456
rect 10432 8444 10450 8458
rect 16240 8444 16258 8458
rect 16960 8446 17270 8456
rect 18544 8446 26546 8456
rect 4060 8422 6458 8432
rect 6784 8422 7394 8432
rect 9256 8422 11534 8432
rect 20296 8420 20314 8434
rect 21328 8422 24614 8432
rect 26392 8422 26450 8432
rect 26488 8422 26869 8432
rect 4072 8398 5738 8408
rect 6400 8398 14006 8408
rect 21472 8398 26474 8408
rect 26512 8398 26869 8408
rect 5716 8374 8714 8384
rect 9520 8372 9538 8386
rect 21736 8374 25430 8384
rect 26440 8374 26498 8384
rect 26536 8374 26869 8384
rect 5728 8350 14690 8360
rect 14704 8350 22166 8360
rect 22180 8350 25154 8360
rect 26464 8350 26869 8360
rect 22696 8326 26522 8336
rect 26560 8326 26869 8336
rect 13744 7493 17306 7503
rect 13672 7469 14450 7479
rect 13096 7445 16850 7455
rect 16864 7445 19898 7455
rect 19912 7445 26282 7455
rect 12976 7421 14642 7431
rect 12952 7397 24314 7407
rect 12448 7373 12506 7383
rect 12904 7373 16610 7383
rect 12016 7349 22394 7359
rect 22408 7349 23570 7359
rect 23584 7349 25874 7359
rect 11992 7325 13490 7335
rect 13504 7325 14546 7335
rect 20176 7325 20858 7335
rect 11512 7301 12698 7311
rect 12760 7301 24026 7311
rect 11464 7277 20378 7287
rect 11368 7253 19970 7263
rect 19984 7253 22922 7263
rect 11296 7229 20162 7239
rect 10936 7205 10946 7215
rect 11008 7205 26330 7215
rect 10840 7181 22514 7191
rect 10264 7157 10346 7167
rect 10504 7157 13634 7167
rect 13648 7157 16538 7167
rect 16552 7157 21170 7167
rect 21184 7157 21938 7167
rect 21952 7157 24050 7167
rect 24064 7157 25586 7167
rect 10072 7133 11618 7143
rect 11632 7133 15026 7143
rect 10000 7109 22130 7119
rect 9952 7085 14066 7095
rect 14848 7085 14942 7095
rect 9928 7061 21746 7071
rect 9592 7037 13730 7047
rect 13744 7037 18986 7047
rect 19000 7037 22994 7047
rect 23008 7037 24146 7047
rect 9400 7013 11090 7023
rect 11104 7013 14834 7023
rect 9328 6989 9386 6999
rect 9520 6989 10058 6999
rect 10120 6989 21962 6999
rect 21976 6989 23642 6999
rect 8992 6965 14618 6975
rect 8992 6941 16322 6951
rect 21736 6941 22214 6951
rect 8920 6917 23546 6927
rect 8632 6893 21722 6903
rect 8440 6869 20642 6879
rect 8248 6845 23834 6855
rect 8080 6821 14474 6831
rect 14488 6821 14858 6831
rect 14872 6821 22850 6831
rect 7912 6797 12602 6807
rect 12688 6797 16466 6807
rect 7864 6773 9482 6783
rect 9496 6773 9578 6783
rect 9592 6773 19178 6783
rect 24976 6773 25034 6783
rect 25120 6773 25394 6783
rect 7696 6749 7730 6759
rect 7816 6749 9194 6759
rect 9208 6749 9626 6759
rect 9784 6749 25106 6759
rect 7672 6725 25442 6735
rect 7600 6701 24962 6711
rect 7600 6677 22898 6687
rect 7288 6653 15794 6663
rect 7264 6629 18218 6639
rect 20128 6629 20306 6639
rect 7144 6605 18770 6615
rect 18784 6605 23738 6615
rect 7096 6581 7106 6591
rect 7192 6581 22730 6591
rect 7072 6557 9434 6567
rect 9448 6557 12746 6567
rect 12856 6557 20114 6567
rect 7048 6533 10490 6543
rect 10504 6533 13154 6543
rect 13168 6533 14570 6543
rect 14584 6533 18170 6543
rect 18184 6533 22538 6543
rect 7024 6509 9674 6519
rect 9688 6509 10202 6519
rect 10216 6509 18890 6519
rect 18904 6509 21338 6519
rect 7000 6485 23858 6495
rect 6976 6461 10778 6471
rect 10792 6461 16010 6471
rect 16696 6461 25706 6471
rect 6904 6437 13346 6447
rect 13624 6437 13922 6447
rect 16672 6437 16730 6447
rect 20080 6437 24350 6447
rect 6712 6413 12314 6423
rect 12328 6413 15626 6423
rect 16432 6413 21554 6423
rect 6688 6389 9098 6399
rect 9112 6389 13322 6399
rect 13552 6389 14234 6399
rect 16192 6389 26474 6399
rect 6664 6365 9122 6375
rect 9136 6365 25202 6375
rect 6496 6341 8858 6351
rect 8920 6341 12074 6351
rect 12160 6341 16826 6351
rect 17008 6341 17066 6351
rect 18640 6341 23018 6351
rect 6376 6317 6386 6327
rect 6448 6317 20066 6327
rect 20536 6317 21026 6327
rect 21280 6317 25778 6327
rect 6352 6293 12482 6303
rect 12496 6293 13898 6303
rect 16168 6293 22634 6303
rect 22648 6293 23354 6303
rect 6304 6269 13706 6279
rect 13816 6269 22418 6279
rect 6232 6245 26210 6255
rect 6208 6221 7370 6231
rect 7432 6221 17378 6231
rect 17392 6221 21266 6231
rect 6064 6197 6074 6207
rect 6160 6197 9362 6207
rect 9376 6197 12794 6207
rect 12808 6197 18698 6207
rect 18712 6197 21794 6207
rect 21808 6197 22274 6207
rect 22288 6197 23474 6207
rect 25360 6197 25634 6207
rect 5968 6173 11474 6183
rect 11584 6173 14942 6183
rect 14956 6173 16274 6183
rect 16288 6173 18626 6183
rect 18640 6173 24506 6183
rect 24520 6173 25346 6183
rect 5800 6149 20522 6159
rect 20536 6149 20690 6159
rect 5752 6125 6554 6135
rect 6616 6125 14282 6135
rect 16144 6125 19082 6135
rect 20368 6125 20822 6135
rect 21688 6125 22034 6135
rect 24808 6125 24866 6135
rect 5704 6101 11282 6111
rect 11296 6101 21674 6111
rect 21688 6101 23582 6111
rect 23596 6101 26162 6111
rect 5608 6077 7658 6087
rect 7672 6077 13250 6087
rect 13264 6077 14306 6087
rect 14320 6077 18842 6087
rect 18856 6077 22970 6087
rect 22984 6077 24794 6087
rect 24808 6077 25850 6087
rect 5488 6053 8498 6063
rect 8512 6053 10322 6063
rect 10336 6053 13562 6063
rect 13576 6053 15674 6063
rect 15688 6053 17954 6063
rect 17968 6053 20354 6063
rect 20368 6053 22850 6063
rect 5440 6029 20090 6039
rect 5392 6005 11330 6015
rect 11344 6005 12554 6015
rect 12568 6005 15122 6015
rect 15136 6005 15410 6015
rect 15424 6005 17522 6015
rect 17536 6005 20738 6015
rect 20752 6005 25970 6015
rect 5248 5981 19226 5991
rect 5224 5957 6194 5967
rect 6256 5957 17474 5967
rect 17920 5957 17930 5967
rect 5104 5933 20210 5943
rect 5056 5909 5066 5919
rect 5128 5909 13814 5919
rect 14896 5909 14942 5919
rect 15016 5909 20306 5919
rect 5008 5885 19586 5895
rect 20464 5885 21002 5895
rect 4960 5861 5210 5871
rect 5224 5861 11018 5871
rect 11080 5861 11210 5871
rect 11272 5861 20474 5871
rect 24232 5861 24326 5871
rect 4936 5837 23234 5847
rect 23248 5837 24218 5847
rect 4816 5813 7418 5823
rect 7432 5813 8234 5823
rect 8248 5813 9410 5823
rect 9424 5813 10106 5823
rect 10120 5813 13058 5823
rect 13072 5813 16298 5823
rect 16312 5813 20450 5823
rect 4768 5789 18506 5799
rect 18520 5789 26042 5799
rect 4720 5765 20666 5775
rect 4672 5741 5330 5751
rect 5344 5741 11066 5751
rect 11152 5741 19154 5751
rect 19168 5741 22490 5751
rect 4672 5717 8594 5727
rect 8680 5717 20906 5727
rect 4576 5693 8282 5703
rect 8296 5693 9290 5703
rect 9304 5693 13514 5703
rect 13528 5693 14186 5703
rect 14200 5693 14786 5703
rect 14800 5693 19922 5703
rect 19936 5693 22058 5703
rect 22072 5693 22778 5703
rect 22792 5693 25514 5703
rect 4528 5669 16034 5679
rect 16096 5669 23402 5679
rect 4504 5645 23090 5655
rect 4456 5621 8642 5631
rect 8800 5621 16466 5631
rect 16528 5621 24722 5631
rect 4432 5597 18458 5607
rect 18928 5597 18962 5607
rect 20800 5597 26066 5607
rect 4336 5573 21242 5583
rect 21472 5573 21650 5583
rect 4240 5549 13226 5559
rect 13408 5549 15362 5559
rect 15376 5549 17762 5559
rect 17776 5549 19682 5559
rect 19696 5549 20786 5559
rect 20800 5549 20822 5559
rect 20836 5549 21458 5559
rect 21472 5549 21602 5559
rect 21616 5549 24170 5559
rect 4216 5525 12866 5535
rect 12880 5525 14342 5535
rect 14356 5525 14402 5535
rect 14416 5525 17738 5535
rect 17752 5525 23498 5535
rect 4192 5501 7706 5511
rect 7768 5501 12434 5511
rect 12448 5501 14498 5511
rect 14512 5501 17210 5511
rect 17224 5501 24458 5511
rect 25312 5501 25490 5511
rect 4168 5477 18914 5487
rect 18928 5477 25298 5487
rect 4120 5453 6338 5463
rect 6352 5453 6962 5463
rect 6976 5453 7778 5463
rect 7792 5453 8546 5463
rect 8560 5453 10922 5463
rect 10936 5453 18722 5463
rect 19048 5453 19058 5463
rect 19144 5453 19322 5463
rect 19864 5453 20306 5463
rect 4096 5429 22322 5439
rect 4048 5405 15434 5415
rect 15856 5405 20138 5415
rect 4048 5381 21506 5391
rect 4024 5357 23306 5367
rect 3976 5333 9818 5343
rect 9832 5333 20954 5343
rect 22696 5333 23102 5343
rect 3928 5309 12026 5319
rect 12112 5309 18122 5319
rect 18304 5309 22994 5319
rect 3904 5285 11570 5295
rect 11632 5285 23450 5295
rect 3832 5261 9698 5271
rect 9760 5261 20402 5271
rect 20776 5261 21098 5271
rect 22264 5261 22826 5271
rect 25624 5261 25946 5271
rect 3808 5237 25610 5247
rect 3712 5213 4538 5223
rect 4552 5213 7898 5223
rect 7912 5213 13082 5223
rect 13096 5213 17138 5223
rect 17152 5213 22682 5223
rect 22696 5213 25994 5223
rect 3616 5189 22250 5199
rect 22264 5189 24938 5199
rect 3616 5165 5258 5175
rect 5320 5165 17690 5175
rect 17704 5165 24266 5175
rect 24280 5165 24842 5175
rect 3568 5141 5618 5151
rect 5632 5141 6410 5151
rect 6424 5141 18578 5151
rect 19024 5141 24098 5151
rect 3472 5117 12386 5127
rect 12544 5117 14426 5127
rect 14440 5117 25634 5127
rect 3448 5093 13754 5103
rect 13768 5093 21290 5103
rect 3184 5069 25370 5079
rect 3160 5045 11498 5055
rect 11512 5045 17906 5055
rect 17920 5045 25562 5055
rect 3136 5021 23882 5031
rect 3088 4997 13778 5007
rect 14176 4997 19982 5007
rect 20344 4997 24170 5007
rect 3064 4973 6362 4983
rect 6376 4973 6842 4983
rect 6856 4973 8858 4983
rect 8872 4973 18386 4983
rect 18400 4973 19706 4983
rect 19720 4973 21818 4983
rect 3040 4949 4610 4959
rect 4624 4949 4730 4959
rect 4744 4949 5546 4959
rect 5560 4949 6050 4959
rect 6136 4949 24194 4959
rect 3016 4925 7922 4935
rect 7936 4925 19850 4935
rect 19864 4925 22298 4935
rect 22312 4925 23066 4935
rect 23080 4925 23762 4935
rect 2896 4901 3650 4911
rect 3664 4901 6506 4911
rect 6520 4901 12818 4911
rect 12832 4901 25274 4911
rect 2896 4877 16706 4887
rect 16912 4877 23954 4887
rect 2824 4853 10226 4863
rect 10240 4853 19826 4863
rect 20248 4853 20978 4863
rect 2776 4829 9938 4839
rect 9952 4829 12986 4839
rect 13120 4829 19562 4839
rect 20056 4829 20834 4839
rect 2752 4805 10802 4815
rect 10888 4805 26869 4815
rect 2704 4781 3290 4791
rect 3304 4781 3674 4791
rect 3688 4781 4466 4791
rect 4480 4781 5186 4791
rect 5200 4781 7682 4791
rect 7696 4781 7874 4791
rect 7888 4781 7970 4791
rect 7984 4781 8618 4791
rect 8632 4781 13418 4791
rect 13432 4781 15506 4791
rect 15520 4781 20546 4791
rect 20560 4781 23258 4791
rect 23272 4781 25274 4791
rect 2680 4757 25010 4767
rect 25096 4757 25322 4767
rect 2632 4733 10250 4743
rect 10552 4733 12458 4743
rect 12472 4733 23042 4743
rect 23296 4733 23318 4743
rect 23680 4733 25730 4743
rect 2608 4709 5354 4719
rect 5368 4709 10130 4719
rect 10144 4709 11162 4719
rect 11176 4709 20594 4719
rect 20608 4709 22586 4719
rect 22600 4709 22874 4719
rect 22888 4709 23522 4719
rect 23536 4709 23834 4719
rect 25072 4709 25226 4719
rect 2584 4685 3266 4695
rect 3328 4685 19130 4695
rect 19144 4685 26018 4695
rect 2560 4661 13130 4671
rect 13288 4661 14210 4671
rect 14272 4661 19346 4671
rect 19648 4661 24326 4671
rect 25000 4661 25130 4671
rect 25216 4661 25442 4671
rect 25792 4661 26378 4671
rect 2536 4637 8954 4647
rect 9040 4637 25490 4647
rect 2488 4613 11234 4623
rect 11248 4613 17186 4623
rect 17200 4613 19706 4623
rect 21064 4613 22214 4623
rect 22576 4613 24002 4623
rect 24280 4613 24350 4623
rect 25024 4613 25466 4623
rect 2440 4589 3938 4599
rect 4000 4589 14666 4599
rect 14752 4589 24818 4599
rect 25384 4589 25850 4599
rect 2416 4565 2906 4575
rect 2920 4565 4274 4575
rect 4288 4565 9914 4575
rect 9928 4565 10898 4575
rect 10912 4565 14042 4575
rect 14056 4565 22658 4575
rect 22888 4565 23546 4575
rect 2392 4541 7946 4551
rect 7960 4541 22514 4551
rect 2344 4517 3338 4527
rect 3352 4517 19802 4527
rect 22072 4517 22538 4527
rect 2320 4493 3578 4503
rect 3592 4493 6026 4503
rect 6040 4493 7754 4503
rect 7768 4493 10706 4503
rect 10720 4493 12674 4503
rect 12688 4493 13874 4503
rect 13888 4493 14282 4503
rect 14296 4493 14882 4503
rect 14896 4493 15722 4503
rect 15736 4493 16682 4503
rect 16696 4493 19538 4503
rect 19552 4493 21530 4503
rect 21544 4493 22010 4503
rect 22024 4493 22082 4503
rect 22096 4493 26306 4503
rect 2296 4469 4394 4479
rect 4408 4469 7154 4479
rect 7168 4469 7466 4479
rect 7480 4469 8306 4479
rect 8320 4469 20810 4479
rect 20824 4469 21770 4479
rect 21784 4469 23282 4479
rect 2296 4445 19610 4455
rect 21544 4445 21746 4455
rect 22024 4445 23102 4455
rect 2224 4421 2978 4431
rect 2992 4421 3242 4431
rect 3256 4421 3890 4431
rect 3904 4421 4634 4431
rect 4648 4421 9314 4431
rect 9328 4421 13298 4431
rect 13312 4421 17882 4431
rect 17896 4421 19946 4431
rect 19960 4421 20762 4431
rect 2176 4397 13274 4407
rect 13288 4397 14162 4407
rect 14176 4397 19490 4407
rect 19504 4397 22706 4407
rect 2128 4373 19418 4383
rect 19552 4373 19898 4383
rect 2104 4349 2234 4359
rect 2248 4349 2354 4359
rect 2368 4349 5930 4359
rect 5944 4349 6602 4359
rect 6616 4349 9458 4359
rect 9472 4349 10274 4359
rect 10288 4349 12362 4359
rect 12376 4349 12914 4359
rect 12928 4349 13178 4359
rect 13192 4349 16922 4359
rect 16936 4349 17978 4359
rect 17992 4349 20498 4359
rect 20512 4349 25082 4359
rect 2080 4325 19874 4335
rect 2032 4301 6530 4311
rect 6592 4301 18314 4311
rect 18712 4301 21074 4311
rect 21088 4301 21650 4311
rect 1984 4277 3554 4287
rect 3568 4277 4610 4287
rect 4624 4277 5162 4287
rect 5176 4277 7322 4287
rect 7336 4277 10562 4287
rect 10648 4277 23066 4287
rect 1936 4253 9794 4263
rect 9904 4253 21914 4263
rect 1888 4229 4370 4239
rect 4384 4229 9098 4239
rect 9112 4229 16994 4239
rect 17272 4229 23138 4239
rect 1840 4205 10466 4215
rect 10480 4205 18050 4215
rect 18064 4205 25754 4215
rect 1792 4181 5042 4191
rect 5056 4181 6770 4191
rect 6784 4181 15386 4191
rect 15400 4181 15578 4191
rect 15592 4181 24602 4191
rect 1768 4157 3482 4167
rect 3496 4157 10682 4167
rect 10696 4157 15554 4167
rect 15664 4157 17858 4167
rect 18760 4157 19322 4167
rect 1720 4133 9218 4143
rect 9304 4133 11378 4143
rect 11392 4133 15746 4143
rect 15760 4133 17114 4143
rect 17128 4133 19250 4143
rect 19264 4133 21866 4143
rect 21880 4133 22154 4143
rect 22168 4133 25250 4143
rect 1696 4109 2258 4119
rect 2272 4109 4058 4119
rect 4072 4109 8738 4119
rect 8752 4109 13586 4119
rect 13600 4109 18074 4119
rect 18088 4109 19754 4119
rect 19768 4109 21890 4119
rect 21904 4109 25802 4119
rect 1672 4085 7082 4095
rect 7096 4085 9218 4095
rect 9232 4085 11690 4095
rect 11704 4085 21122 4095
rect 21136 4085 21482 4095
rect 21904 4085 22490 4095
rect 1648 4061 7058 4071
rect 7072 4061 8066 4071
rect 8080 4061 8186 4071
rect 8200 4061 8378 4071
rect 8392 4061 11402 4071
rect 11416 4061 11522 4071
rect 11536 4061 11666 4071
rect 11680 4061 12194 4071
rect 12208 4061 20330 4071
rect 20344 4061 25898 4071
rect 1624 4037 1898 4047
rect 1912 4037 4586 4047
rect 4600 4037 8402 4047
rect 8416 4037 12650 4047
rect 12664 4037 18194 4047
rect 18208 4037 21386 4047
rect 84 4013 10010 4023
rect 10024 4013 13658 4023
rect 13672 4013 17090 4023
rect 17104 4013 21506 4023
rect 84 3989 25418 3999
rect 1696 3965 19466 3975
rect 19768 3965 20210 3975
rect 2008 3941 26450 3951
rect 2056 3917 4826 3927
rect 4840 3917 5498 3927
rect 5512 3917 12578 3927
rect 12592 3917 13946 3927
rect 13960 3917 14090 3927
rect 14104 3917 15602 3927
rect 15616 3917 18818 3927
rect 18832 3917 21602 3927
rect 21616 3917 26090 3927
rect 2512 3893 23090 3903
rect 2608 3869 10970 3879
rect 10984 3869 16802 3879
rect 16912 3869 19274 3879
rect 19288 3869 19778 3879
rect 2632 3845 4874 3855
rect 4888 3845 19202 3855
rect 19216 3845 24242 3855
rect 2704 3821 13538 3831
rect 13552 3821 19658 3831
rect 2728 3797 4202 3807
rect 4264 3797 22466 3807
rect 2944 3773 20042 3783
rect 3232 3749 13898 3759
rect 14056 3749 14342 3759
rect 14536 3749 18962 3759
rect 19024 3749 19346 3759
rect 19360 3749 22106 3759
rect 22120 3749 22442 3759
rect 22456 3749 24386 3759
rect 3256 3725 3290 3735
rect 3400 3725 16754 3735
rect 16768 3725 22346 3735
rect 3304 3701 5402 3711
rect 5416 3701 7202 3711
rect 7216 3701 7730 3711
rect 7744 3701 11546 3711
rect 11560 3701 14210 3711
rect 14224 3701 17858 3711
rect 17872 3701 20882 3711
rect 20896 3701 22610 3711
rect 22624 3701 22946 3711
rect 22960 3701 25658 3711
rect 3448 3677 5090 3687
rect 5104 3677 6098 3687
rect 6112 3677 6794 3687
rect 6808 3677 15410 3687
rect 15424 3677 24626 3687
rect 3520 3653 19370 3663
rect 19480 3653 19682 3663
rect 22624 3653 23234 3663
rect 3688 3629 9530 3639
rect 9544 3629 18410 3639
rect 18424 3629 20618 3639
rect 22960 3629 23582 3639
rect 3736 3605 24050 3615
rect 3784 3581 19082 3591
rect 19216 3581 20858 3591
rect 3808 3557 8522 3567
rect 8536 3557 18818 3567
rect 18832 3557 25058 3567
rect 3856 3533 25706 3543
rect 3928 3509 4298 3519
rect 4312 3509 6074 3519
rect 6088 3509 8210 3519
rect 8224 3509 10346 3519
rect 10360 3509 11906 3519
rect 11920 3509 13202 3519
rect 13216 3509 15314 3519
rect 15328 3509 17330 3519
rect 17344 3509 22466 3519
rect 22480 3509 24074 3519
rect 3952 3485 21098 3495
rect 24088 3485 24098 3495
rect 4120 3461 8138 3471
rect 8152 3461 21986 3471
rect 22000 3461 22754 3471
rect 22768 3461 23186 3471
rect 23200 3461 24986 3471
rect 25000 3461 25754 3471
rect 4312 3437 6914 3447
rect 6928 3437 7298 3447
rect 7312 3437 11594 3447
rect 11608 3437 13010 3447
rect 13024 3437 20930 3447
rect 20944 3437 24530 3447
rect 24544 3437 24746 3447
rect 24760 3437 25250 3447
rect 25264 3437 25682 3447
rect 4336 3413 8714 3423
rect 8728 3413 10178 3423
rect 10192 3413 13970 3423
rect 13984 3413 14906 3423
rect 14920 3413 15890 3423
rect 15904 3413 17018 3423
rect 17032 3413 17354 3423
rect 17368 3413 21794 3423
rect 21808 3413 22274 3423
rect 22288 3413 25130 3423
rect 25696 3413 26042 3423
rect 4408 3389 6242 3399
rect 6256 3389 14330 3399
rect 14344 3389 17426 3399
rect 17440 3389 18266 3399
rect 18856 3389 18890 3399
rect 22768 3389 23474 3399
rect 4504 3365 6458 3375
rect 6472 3365 15530 3375
rect 15544 3365 19274 3375
rect 4720 3341 11930 3351
rect 11944 3341 19514 3351
rect 4768 3317 7778 3327
rect 7792 3317 8258 3327
rect 8272 3317 13346 3327
rect 13360 3317 26258 3327
rect 4840 3293 6386 3303
rect 6400 3293 9962 3303
rect 9976 3293 14942 3303
rect 14956 3293 18938 3303
rect 4888 3269 5066 3279
rect 5152 3269 22202 3279
rect 4960 3245 9386 3255
rect 9400 3245 11882 3255
rect 11896 3245 12770 3255
rect 12784 3245 15626 3255
rect 15640 3245 15938 3255
rect 15952 3245 19034 3255
rect 4984 3221 7802 3231
rect 7816 3221 9746 3231
rect 9760 3221 10610 3231
rect 10624 3221 11810 3231
rect 11824 3221 13370 3231
rect 13384 3221 14810 3231
rect 14824 3221 15818 3231
rect 15832 3221 16778 3231
rect 16792 3221 20258 3231
rect 20272 3221 23318 3231
rect 5008 3197 11210 3207
rect 11224 3197 14114 3207
rect 14704 3197 23210 3207
rect 5080 3173 21314 3183
rect 21328 3173 21698 3183
rect 23224 3173 26426 3183
rect 5176 3149 5210 3159
rect 5272 3149 7106 3159
rect 7240 3149 7994 3159
rect 8104 3149 12626 3159
rect 12640 3149 15698 3159
rect 15712 3149 23378 3159
rect 23392 3149 25154 3159
rect 5224 3125 20834 3135
rect 5296 3101 8786 3111
rect 8848 3101 26114 3111
rect 5368 3077 10418 3087
rect 10624 3077 14450 3087
rect 15112 3077 18866 3087
rect 18880 3077 20186 3087
rect 5488 3053 6266 3063
rect 6328 3053 21194 3063
rect 5656 3029 23258 3039
rect 5848 3005 9986 3015
rect 10048 3005 23786 3015
rect 5848 2981 25178 2991
rect 5896 2957 12938 2967
rect 12952 2957 26186 2967
rect 5920 2933 8018 2943
rect 8128 2933 17834 2943
rect 17848 2933 21026 2943
rect 21040 2933 21626 2943
rect 21640 2933 23786 2943
rect 23800 2933 25178 2943
rect 6136 2909 13994 2919
rect 14008 2909 16586 2919
rect 16600 2909 22826 2919
rect 22840 2909 23162 2919
rect 6472 2885 11114 2895
rect 11128 2885 14138 2895
rect 14152 2885 15482 2895
rect 15496 2885 16706 2895
rect 16720 2885 16874 2895
rect 16888 2885 24914 2895
rect 6592 2861 8474 2871
rect 8488 2861 25922 2871
rect 6736 2837 16754 2847
rect 16816 2837 16826 2847
rect 17584 2837 25034 2847
rect 6880 2813 6938 2823
rect 6952 2813 14234 2823
rect 14248 2813 15698 2823
rect 15712 2813 19730 2823
rect 19744 2813 25538 2823
rect 7120 2789 8090 2799
rect 8104 2789 10154 2799
rect 10168 2789 10298 2799
rect 10312 2789 11714 2799
rect 11728 2789 16658 2799
rect 16672 2789 20234 2799
rect 23176 2789 23642 2799
rect 7144 2765 9002 2775
rect 9064 2765 23618 2775
rect 7240 2741 16634 2751
rect 16792 2741 25826 2751
rect 7288 2717 9554 2727
rect 9568 2717 9866 2727
rect 9880 2717 19922 2727
rect 19936 2717 20474 2727
rect 20488 2717 20906 2727
rect 20920 2717 21578 2727
rect 21592 2717 22034 2727
rect 22048 2717 25226 2727
rect 7336 2693 19394 2703
rect 19744 2693 19982 2703
rect 20200 2693 20282 2703
rect 7360 2669 7490 2679
rect 7552 2669 9842 2679
rect 9904 2669 13466 2679
rect 13576 2669 14306 2679
rect 15160 2669 20018 2679
rect 20032 2669 24098 2679
rect 7384 2645 7706 2655
rect 7720 2645 25322 2655
rect 7888 2621 7922 2631
rect 8008 2621 8330 2631
rect 8344 2621 23042 2631
rect 7936 2597 20714 2607
rect 8200 2573 8234 2583
rect 8296 2573 12338 2583
rect 12352 2573 24122 2583
rect 8344 2549 17066 2559
rect 17632 2549 21842 2559
rect 24136 2549 24146 2559
rect 8392 2525 10586 2535
rect 10600 2525 14930 2535
rect 15208 2525 22178 2535
rect 8536 2501 15770 2511
rect 15784 2501 18362 2511
rect 18376 2501 22370 2511
rect 8680 2477 20306 2487
rect 20728 2477 21074 2487
rect 22384 2477 23018 2487
rect 8848 2453 9146 2463
rect 9352 2453 11786 2463
rect 11848 2453 14594 2463
rect 15256 2453 16226 2463
rect 16528 2453 16946 2463
rect 17800 2453 19442 2463
rect 9184 2429 18002 2439
rect 18016 2429 19298 2439
rect 9448 2405 9482 2415
rect 9616 2405 12578 2415
rect 12712 2405 20426 2415
rect 9664 2381 13994 2391
rect 14080 2381 14378 2391
rect 14392 2381 14546 2391
rect 15568 2381 16442 2391
rect 16576 2381 25946 2391
rect 9688 2357 11186 2367
rect 11248 2357 16730 2367
rect 18952 2357 18986 2367
rect 9808 2333 9914 2343
rect 10192 2333 10322 2343
rect 10672 2333 10850 2343
rect 10864 2333 20570 2343
rect 20584 2333 23426 2343
rect 10312 2309 10370 2319
rect 10720 2309 19058 2319
rect 10744 2285 15290 2295
rect 10816 2261 24554 2271
rect 10840 2237 10946 2247
rect 11008 2237 13850 2247
rect 13864 2237 24938 2247
rect 10888 2213 11450 2223
rect 11464 2213 14018 2223
rect 11032 2189 18482 2199
rect 18496 2189 22802 2199
rect 22816 2189 24290 2199
rect 24304 2189 24866 2199
rect 11104 2165 26426 2175
rect 11152 2141 12194 2151
rect 12208 2141 23930 2151
rect 11200 2117 20978 2127
rect 11224 2093 16298 2103
rect 16312 2093 23978 2103
rect 11320 2069 12506 2079
rect 12520 2069 17714 2079
rect 23992 2069 24098 2079
rect 11344 2045 13682 2055
rect 13792 2045 14474 2055
rect 11560 2021 17042 2031
rect 17056 2021 20378 2031
rect 11752 1997 16442 2007
rect 12256 1973 13442 1983
rect 12352 1949 13034 1959
rect 13120 1949 16370 1959
rect 12568 1925 12602 1935
rect 12808 1925 21002 1935
rect 12856 1901 17930 1911
rect 12904 1877 16394 1887
rect 13000 1853 13322 1863
rect 13408 1853 24410 1863
rect 26440 1853 26869 1863
rect 13192 1829 13754 1839
rect 26488 1829 26869 1839
rect 13216 1805 13814 1815
rect 26464 1805 26869 1815
rect 25803 1776 26450 1786
rect 25803 1753 26450 1763
rect 25803 1724 25808 1740
rect 26443 1724 26450 1740
rect 25803 1715 26450 1724
rect 25803 1086 26450 1095
rect 25803 1070 25808 1086
rect 26443 1070 26450 1086
rect 25803 1047 26450 1057
rect 25803 1024 26450 1034
rect 25803 1001 26450 1011
rect 16600 972 18866 982
rect 15904 948 18434 958
rect 15352 924 17546 934
rect 13864 900 23306 910
rect 11056 876 25490 886
rect 10960 852 25562 862
rect 10792 828 14114 838
rect 14488 828 16850 838
rect 16960 828 22898 838
rect 10456 804 15218 814
rect 15232 804 19298 814
rect 10408 780 22178 790
rect 10384 756 20282 766
rect 9496 732 20666 742
rect 9064 708 17642 718
rect 17656 708 22802 718
rect 9016 684 23426 694
rect 8968 660 20618 670
rect 8752 636 19970 646
rect 8728 612 25394 622
rect 8656 588 17138 598
rect 17464 586 17482 600
rect 18976 588 19946 598
rect 8176 564 19634 574
rect 7840 540 20018 550
rect 7624 516 24386 526
rect 7576 492 8210 502
rect 8584 492 21002 502
rect 23008 490 23026 504
rect 7552 468 12386 478
rect 13048 468 22298 478
rect 7192 444 18578 454
rect 18592 444 21626 454
rect 6712 420 19418 430
rect 6664 396 6722 406
rect 7048 396 21818 406
rect 6184 372 8426 382
rect 8440 372 11402 382
rect 13312 372 24146 382
rect 6088 348 23138 358
rect 5296 324 6770 334
rect 6832 324 13466 334
rect 13480 324 20834 334
rect 5128 300 16826 310
rect 3856 276 14978 286
rect 15064 276 25442 286
rect 3736 252 6026 262
rect 6040 252 21146 262
rect 2656 228 20570 238
rect 2584 204 22394 214
rect 2392 180 3986 190
rect 4144 180 11666 190
rect 13600 180 24002 190
rect 2344 156 4346 166
rect 4432 154 4450 168
rect 4648 156 25610 166
rect 84 132 12602 142
rect 13696 132 21770 142
rect 84 108 2426 118
rect 2488 108 18026 118
rect 6280 84 7814 94
rect 8128 84 9554 94
rect 10360 84 14210 94
rect 15016 84 17042 94
rect 25576 84 26869 94
rect 7504 60 25562 70
rect 25600 60 26869 70
rect 10600 36 25586 46
rect 25624 36 26869 46
rect 11320 12 26869 22
<< m2contact >>
rect 6794 8564 6808 8578
rect 9014 8564 9028 8578
rect 19130 8564 19144 8578
rect 22142 8564 22156 8578
rect 24866 8564 24880 8578
rect 5306 8540 5320 8554
rect 16454 8540 16468 8554
rect 21326 8540 21340 8554
rect 24338 8540 24352 8554
rect 5042 8516 5056 8530
rect 13190 8516 13204 8530
rect 18878 8516 18892 8530
rect 23210 8516 23224 8530
rect 23774 8516 23788 8530
rect 26186 8516 26200 8530
rect 2306 8492 2320 8506
rect 3218 8492 3232 8506
rect 4298 8492 4312 8506
rect 4874 8492 4888 8506
rect 10610 8492 10624 8506
rect 13154 8492 13168 8506
rect 13946 8492 13960 8506
rect 15614 8492 15628 8506
rect 18962 8492 18976 8506
rect 19694 8492 19708 8506
rect 25466 8492 25480 8506
rect 70 8468 84 8482
rect 10922 8468 10936 8482
rect 11186 8468 11200 8482
rect 12482 8468 12496 8482
rect 23798 8468 23812 8482
rect 70 8444 84 8458
rect 10370 8444 10384 8458
rect 10418 8444 10432 8458
rect 16226 8444 16240 8458
rect 16946 8444 16960 8458
rect 17270 8444 17284 8458
rect 18530 8444 18544 8458
rect 26546 8444 26560 8458
rect 4046 8420 4060 8434
rect 6458 8420 6472 8434
rect 6770 8420 6784 8434
rect 7394 8420 7408 8434
rect 9242 8420 9256 8434
rect 11534 8420 11548 8434
rect 20282 8420 20296 8434
rect 21314 8420 21328 8434
rect 24614 8420 24628 8434
rect 26378 8420 26392 8434
rect 26450 8420 26464 8434
rect 26474 8420 26488 8434
rect 26869 8420 26883 8434
rect 4058 8396 4072 8410
rect 5738 8396 5752 8410
rect 6386 8396 6400 8410
rect 14006 8396 14020 8410
rect 21458 8396 21472 8410
rect 26474 8396 26488 8410
rect 26498 8396 26512 8410
rect 26869 8396 26883 8410
rect 5702 8372 5716 8386
rect 8714 8372 8728 8386
rect 9506 8372 9520 8386
rect 21722 8372 21736 8386
rect 25430 8372 25444 8386
rect 26426 8372 26440 8386
rect 26498 8372 26512 8386
rect 26522 8372 26536 8386
rect 26869 8372 26883 8386
rect 5714 8348 5728 8362
rect 14690 8348 14704 8362
rect 22166 8348 22180 8362
rect 25154 8348 25168 8362
rect 26450 8348 26464 8362
rect 26869 8348 26883 8362
rect 22682 8324 22696 8338
rect 26522 8324 26536 8338
rect 26546 8324 26560 8338
rect 26869 8324 26883 8338
rect 13730 7491 13744 7505
rect 17306 7491 17320 7505
rect 13658 7467 13672 7481
rect 14450 7467 14464 7481
rect 13082 7443 13096 7457
rect 16850 7443 16864 7457
rect 19898 7443 19912 7457
rect 26282 7443 26296 7457
rect 12962 7419 12976 7433
rect 14642 7419 14656 7433
rect 12938 7395 12952 7409
rect 24314 7395 24328 7409
rect 12434 7371 12448 7385
rect 12506 7371 12520 7385
rect 12890 7371 12904 7385
rect 16610 7371 16624 7385
rect 12002 7347 12016 7361
rect 22394 7347 22408 7361
rect 23570 7347 23584 7361
rect 25874 7347 25888 7361
rect 11978 7323 11992 7337
rect 13490 7323 13504 7337
rect 14546 7323 14560 7337
rect 20162 7323 20176 7337
rect 20858 7323 20872 7337
rect 11498 7299 11512 7313
rect 12698 7299 12712 7313
rect 12746 7299 12760 7313
rect 24026 7299 24040 7313
rect 11450 7275 11464 7289
rect 20378 7275 20392 7289
rect 11354 7251 11368 7265
rect 19970 7251 19984 7265
rect 22922 7251 22936 7265
rect 11282 7227 11296 7241
rect 20162 7227 20176 7241
rect 10922 7203 10936 7217
rect 10946 7203 10960 7217
rect 10994 7203 11008 7217
rect 26330 7203 26344 7217
rect 10826 7179 10840 7193
rect 22514 7179 22528 7193
rect 10250 7155 10264 7169
rect 10346 7155 10360 7169
rect 10490 7155 10504 7169
rect 13634 7155 13648 7169
rect 16538 7155 16552 7169
rect 21170 7155 21184 7169
rect 21938 7155 21952 7169
rect 24050 7155 24064 7169
rect 25586 7155 25600 7169
rect 10058 7131 10072 7145
rect 11618 7131 11632 7145
rect 15026 7131 15040 7145
rect 9986 7107 10000 7121
rect 22130 7107 22144 7121
rect 9938 7083 9952 7097
rect 14066 7083 14080 7097
rect 14834 7083 14848 7097
rect 14942 7083 14956 7097
rect 9914 7059 9928 7073
rect 21746 7059 21760 7073
rect 9578 7035 9592 7049
rect 13730 7035 13744 7049
rect 18986 7035 19000 7049
rect 22994 7035 23008 7049
rect 24146 7035 24160 7049
rect 9386 7011 9400 7025
rect 11090 7011 11104 7025
rect 14834 7011 14848 7025
rect 9314 6987 9328 7001
rect 9386 6987 9400 7001
rect 9506 6987 9520 7001
rect 10058 6987 10072 7001
rect 10106 6987 10120 7001
rect 21962 6987 21976 7001
rect 23642 6987 23656 7001
rect 8978 6963 8992 6977
rect 14618 6963 14632 6977
rect 8978 6939 8992 6953
rect 16322 6939 16336 6953
rect 21722 6939 21736 6953
rect 22214 6939 22228 6953
rect 8906 6915 8920 6929
rect 23546 6915 23560 6929
rect 8618 6891 8632 6905
rect 21722 6891 21736 6905
rect 8426 6867 8440 6881
rect 20642 6867 20656 6881
rect 8234 6843 8248 6857
rect 23834 6843 23848 6857
rect 8066 6819 8080 6833
rect 14474 6819 14488 6833
rect 14858 6819 14872 6833
rect 22850 6819 22864 6833
rect 7898 6795 7912 6809
rect 12602 6795 12616 6809
rect 12674 6795 12688 6809
rect 16466 6795 16480 6809
rect 7850 6771 7864 6785
rect 9482 6771 9496 6785
rect 9578 6771 9592 6785
rect 19178 6771 19192 6785
rect 24962 6771 24976 6785
rect 25034 6771 25048 6785
rect 25106 6771 25120 6785
rect 25394 6771 25408 6785
rect 7682 6747 7696 6761
rect 7730 6747 7744 6761
rect 7802 6747 7816 6761
rect 9194 6747 9208 6761
rect 9626 6747 9640 6761
rect 9770 6747 9784 6761
rect 25106 6747 25120 6761
rect 7658 6723 7672 6737
rect 25442 6723 25456 6737
rect 7586 6699 7600 6713
rect 24962 6699 24976 6713
rect 7586 6675 7600 6689
rect 22898 6675 22912 6689
rect 7274 6651 7288 6665
rect 15794 6651 15808 6665
rect 7250 6627 7264 6641
rect 18218 6627 18232 6641
rect 20114 6627 20128 6641
rect 20306 6627 20320 6641
rect 7130 6603 7144 6617
rect 18770 6603 18784 6617
rect 23738 6603 23752 6617
rect 7082 6579 7096 6593
rect 7106 6579 7120 6593
rect 7178 6579 7192 6593
rect 22730 6579 22744 6593
rect 7058 6555 7072 6569
rect 9434 6555 9448 6569
rect 12746 6555 12760 6569
rect 12842 6555 12856 6569
rect 20114 6555 20128 6569
rect 7034 6531 7048 6545
rect 10490 6531 10504 6545
rect 13154 6531 13168 6545
rect 14570 6531 14584 6545
rect 18170 6531 18184 6545
rect 22538 6531 22552 6545
rect 7010 6507 7024 6521
rect 9674 6507 9688 6521
rect 10202 6507 10216 6521
rect 18890 6507 18904 6521
rect 21338 6507 21352 6521
rect 6986 6483 7000 6497
rect 23858 6483 23872 6497
rect 6962 6459 6976 6473
rect 10778 6459 10792 6473
rect 16010 6459 16024 6473
rect 16682 6459 16696 6473
rect 25706 6459 25720 6473
rect 6890 6435 6904 6449
rect 13346 6435 13360 6449
rect 13610 6435 13624 6449
rect 13922 6435 13936 6449
rect 16658 6435 16672 6449
rect 16730 6435 16744 6449
rect 20066 6435 20080 6449
rect 24350 6435 24364 6449
rect 6698 6411 6712 6425
rect 12314 6411 12328 6425
rect 15626 6411 15640 6425
rect 16418 6411 16432 6425
rect 21554 6411 21568 6425
rect 6674 6387 6688 6401
rect 9098 6387 9112 6401
rect 13322 6387 13336 6401
rect 13538 6387 13552 6401
rect 14234 6387 14248 6401
rect 16178 6387 16192 6401
rect 26474 6387 26488 6401
rect 6650 6363 6664 6377
rect 9122 6363 9136 6377
rect 25202 6363 25216 6377
rect 6482 6339 6496 6353
rect 8858 6339 8872 6353
rect 8906 6339 8920 6353
rect 12074 6339 12088 6353
rect 12146 6339 12160 6353
rect 16826 6339 16840 6353
rect 16994 6339 17008 6353
rect 17066 6339 17080 6353
rect 18626 6339 18640 6353
rect 23018 6339 23032 6353
rect 6362 6315 6376 6329
rect 6386 6315 6400 6329
rect 6434 6315 6448 6329
rect 20066 6315 20080 6329
rect 20522 6315 20536 6329
rect 21026 6315 21040 6329
rect 21266 6315 21280 6329
rect 25778 6315 25792 6329
rect 6338 6291 6352 6305
rect 12482 6291 12496 6305
rect 13898 6291 13912 6305
rect 16154 6291 16168 6305
rect 22634 6291 22648 6305
rect 23354 6291 23368 6305
rect 6290 6267 6304 6281
rect 13706 6267 13720 6281
rect 13802 6267 13816 6281
rect 22418 6267 22432 6281
rect 6218 6243 6232 6257
rect 26210 6243 26224 6257
rect 6194 6219 6208 6233
rect 7370 6219 7384 6233
rect 7418 6219 7432 6233
rect 17378 6219 17392 6233
rect 21266 6219 21280 6233
rect 6050 6195 6064 6209
rect 6074 6195 6088 6209
rect 6146 6195 6160 6209
rect 9362 6195 9376 6209
rect 12794 6195 12808 6209
rect 18698 6195 18712 6209
rect 21794 6195 21808 6209
rect 22274 6195 22288 6209
rect 23474 6195 23488 6209
rect 25346 6195 25360 6209
rect 25634 6195 25648 6209
rect 5954 6171 5968 6185
rect 11474 6171 11488 6185
rect 11570 6171 11584 6185
rect 14942 6171 14956 6185
rect 16274 6171 16288 6185
rect 18626 6171 18640 6185
rect 24506 6171 24520 6185
rect 25346 6171 25360 6185
rect 5786 6147 5800 6161
rect 20522 6147 20536 6161
rect 20690 6147 20704 6161
rect 5738 6123 5752 6137
rect 6554 6123 6568 6137
rect 6602 6123 6616 6137
rect 14282 6123 14296 6137
rect 16130 6123 16144 6137
rect 19082 6123 19096 6137
rect 20354 6123 20368 6137
rect 20822 6123 20836 6137
rect 21674 6123 21688 6137
rect 22034 6123 22048 6137
rect 24794 6123 24808 6137
rect 24866 6123 24880 6137
rect 5690 6099 5704 6113
rect 11282 6099 11296 6113
rect 21674 6099 21688 6113
rect 23582 6099 23596 6113
rect 26162 6099 26176 6113
rect 5594 6075 5608 6089
rect 7658 6075 7672 6089
rect 13250 6075 13264 6089
rect 14306 6075 14320 6089
rect 18842 6075 18856 6089
rect 22970 6075 22984 6089
rect 24794 6075 24808 6089
rect 25850 6075 25864 6089
rect 5474 6051 5488 6065
rect 8498 6051 8512 6065
rect 10322 6051 10336 6065
rect 13562 6051 13576 6065
rect 15674 6051 15688 6065
rect 17954 6051 17968 6065
rect 20354 6051 20368 6065
rect 22850 6051 22864 6065
rect 5426 6027 5440 6041
rect 20090 6027 20104 6041
rect 5378 6003 5392 6017
rect 11330 6003 11344 6017
rect 12554 6003 12568 6017
rect 15122 6003 15136 6017
rect 15410 6003 15424 6017
rect 17522 6003 17536 6017
rect 20738 6003 20752 6017
rect 25970 6003 25984 6017
rect 5234 5979 5248 5993
rect 19226 5979 19240 5993
rect 5210 5955 5224 5969
rect 6194 5955 6208 5969
rect 6242 5955 6256 5969
rect 17474 5955 17488 5969
rect 17906 5955 17920 5969
rect 17930 5955 17944 5969
rect 5090 5931 5104 5945
rect 20210 5931 20224 5945
rect 5042 5907 5056 5921
rect 5066 5907 5080 5921
rect 5114 5907 5128 5921
rect 13814 5907 13828 5921
rect 14882 5907 14896 5921
rect 14942 5907 14956 5921
rect 15002 5907 15016 5921
rect 20306 5907 20320 5921
rect 4994 5883 5008 5897
rect 19586 5883 19600 5897
rect 20450 5883 20464 5897
rect 21002 5883 21016 5897
rect 4946 5859 4960 5873
rect 5210 5859 5224 5873
rect 11018 5859 11032 5873
rect 11066 5859 11080 5873
rect 11210 5859 11224 5873
rect 11258 5859 11272 5873
rect 20474 5859 20488 5873
rect 24218 5859 24232 5873
rect 24326 5859 24340 5873
rect 4922 5835 4936 5849
rect 23234 5835 23248 5849
rect 24218 5835 24232 5849
rect 4802 5811 4816 5825
rect 7418 5811 7432 5825
rect 8234 5811 8248 5825
rect 9410 5811 9424 5825
rect 10106 5811 10120 5825
rect 13058 5811 13072 5825
rect 16298 5811 16312 5825
rect 20450 5811 20464 5825
rect 4754 5787 4768 5801
rect 18506 5787 18520 5801
rect 26042 5787 26056 5801
rect 4706 5763 4720 5777
rect 20666 5763 20680 5777
rect 4658 5739 4672 5753
rect 5330 5739 5344 5753
rect 11066 5739 11080 5753
rect 11138 5739 11152 5753
rect 19154 5739 19168 5753
rect 22490 5739 22504 5753
rect 4658 5715 4672 5729
rect 8594 5715 8608 5729
rect 8666 5715 8680 5729
rect 20906 5715 20920 5729
rect 4562 5691 4576 5705
rect 8282 5691 8296 5705
rect 9290 5691 9304 5705
rect 13514 5691 13528 5705
rect 14186 5691 14200 5705
rect 14786 5691 14800 5705
rect 19922 5691 19936 5705
rect 22058 5691 22072 5705
rect 22778 5691 22792 5705
rect 25514 5691 25528 5705
rect 4514 5667 4528 5681
rect 16034 5667 16048 5681
rect 16082 5667 16096 5681
rect 23402 5667 23416 5681
rect 4490 5643 4504 5657
rect 23090 5643 23104 5657
rect 4442 5619 4456 5633
rect 8642 5619 8656 5633
rect 8786 5619 8800 5633
rect 16466 5619 16480 5633
rect 16514 5619 16528 5633
rect 24722 5619 24736 5633
rect 4418 5595 4432 5609
rect 18458 5595 18472 5609
rect 18914 5595 18928 5609
rect 18962 5595 18976 5609
rect 20786 5595 20800 5609
rect 26066 5595 26080 5609
rect 4322 5571 4336 5585
rect 21242 5571 21256 5585
rect 21458 5571 21472 5585
rect 21650 5571 21664 5585
rect 4226 5547 4240 5561
rect 13226 5547 13240 5561
rect 13394 5547 13408 5561
rect 15362 5547 15376 5561
rect 17762 5547 17776 5561
rect 19682 5547 19696 5561
rect 20786 5547 20800 5561
rect 20822 5547 20836 5561
rect 21458 5547 21472 5561
rect 21602 5547 21616 5561
rect 24170 5547 24184 5561
rect 4202 5523 4216 5537
rect 12866 5523 12880 5537
rect 14342 5523 14356 5537
rect 14402 5523 14416 5537
rect 17738 5523 17752 5537
rect 23498 5523 23512 5537
rect 4178 5499 4192 5513
rect 7706 5499 7720 5513
rect 7754 5499 7768 5513
rect 12434 5499 12448 5513
rect 14498 5499 14512 5513
rect 17210 5499 17224 5513
rect 24458 5499 24472 5513
rect 25298 5499 25312 5513
rect 25490 5499 25504 5513
rect 4154 5475 4168 5489
rect 18914 5475 18928 5489
rect 25298 5475 25312 5489
rect 4106 5451 4120 5465
rect 6338 5451 6352 5465
rect 6962 5451 6976 5465
rect 7778 5451 7792 5465
rect 8546 5451 8560 5465
rect 10922 5451 10936 5465
rect 18722 5451 18736 5465
rect 19034 5451 19048 5465
rect 19058 5451 19072 5465
rect 19130 5451 19144 5465
rect 19322 5451 19336 5465
rect 19850 5451 19864 5465
rect 20306 5451 20320 5465
rect 4082 5427 4096 5441
rect 22322 5427 22336 5441
rect 4034 5403 4048 5417
rect 15434 5403 15448 5417
rect 15842 5403 15856 5417
rect 20138 5403 20152 5417
rect 4034 5379 4048 5393
rect 21506 5379 21520 5393
rect 4010 5355 4024 5369
rect 23306 5355 23320 5369
rect 3962 5331 3976 5345
rect 9818 5331 9832 5345
rect 20954 5331 20968 5345
rect 22682 5331 22696 5345
rect 23102 5331 23116 5345
rect 3914 5307 3928 5321
rect 12026 5307 12040 5321
rect 12098 5307 12112 5321
rect 18122 5307 18136 5321
rect 18290 5307 18304 5321
rect 22994 5307 23008 5321
rect 3890 5283 3904 5297
rect 11570 5283 11584 5297
rect 11618 5283 11632 5297
rect 23450 5283 23464 5297
rect 3818 5259 3832 5273
rect 9698 5259 9712 5273
rect 9746 5259 9760 5273
rect 20402 5259 20416 5273
rect 20762 5259 20776 5273
rect 21098 5259 21112 5273
rect 22250 5259 22264 5273
rect 22826 5259 22840 5273
rect 25610 5259 25624 5273
rect 25946 5259 25960 5273
rect 3794 5235 3808 5249
rect 25610 5235 25624 5249
rect 3698 5211 3712 5225
rect 4538 5211 4552 5225
rect 7898 5211 7912 5225
rect 13082 5211 13096 5225
rect 17138 5211 17152 5225
rect 22682 5211 22696 5225
rect 25994 5211 26008 5225
rect 3602 5187 3616 5201
rect 22250 5187 22264 5201
rect 24938 5187 24952 5201
rect 3602 5163 3616 5177
rect 5258 5163 5272 5177
rect 5306 5163 5320 5177
rect 17690 5163 17704 5177
rect 24266 5163 24280 5177
rect 24842 5163 24856 5177
rect 3554 5139 3568 5153
rect 5618 5139 5632 5153
rect 6410 5139 6424 5153
rect 18578 5139 18592 5153
rect 19010 5139 19024 5153
rect 24098 5139 24112 5153
rect 3458 5115 3472 5129
rect 12386 5115 12400 5129
rect 12530 5115 12544 5129
rect 14426 5115 14440 5129
rect 25634 5115 25648 5129
rect 3434 5091 3448 5105
rect 13754 5091 13768 5105
rect 21290 5091 21304 5105
rect 3170 5067 3184 5081
rect 25370 5067 25384 5081
rect 3146 5043 3160 5057
rect 11498 5043 11512 5057
rect 17906 5043 17920 5057
rect 25562 5043 25576 5057
rect 3122 5019 3136 5033
rect 23882 5019 23896 5033
rect 3074 4995 3088 5009
rect 13778 4995 13792 5009
rect 14162 4995 14176 5009
rect 19982 4995 19996 5009
rect 20330 4995 20344 5009
rect 24170 4995 24184 5009
rect 3050 4971 3064 4985
rect 6362 4971 6376 4985
rect 6842 4971 6856 4985
rect 8858 4971 8872 4985
rect 18386 4971 18400 4985
rect 19706 4971 19720 4985
rect 21818 4971 21832 4985
rect 3026 4947 3040 4961
rect 4610 4947 4624 4961
rect 4730 4947 4744 4961
rect 5546 4947 5560 4961
rect 6050 4947 6064 4961
rect 6122 4947 6136 4961
rect 24194 4947 24208 4961
rect 3002 4923 3016 4937
rect 7922 4923 7936 4937
rect 19850 4923 19864 4937
rect 22298 4923 22312 4937
rect 23066 4923 23080 4937
rect 23762 4923 23776 4937
rect 2882 4899 2896 4913
rect 3650 4899 3664 4913
rect 6506 4899 6520 4913
rect 12818 4899 12832 4913
rect 25274 4899 25288 4913
rect 2882 4875 2896 4889
rect 16706 4875 16720 4889
rect 16898 4875 16912 4889
rect 23954 4875 23968 4889
rect 2810 4851 2824 4865
rect 10226 4851 10240 4865
rect 19826 4851 19840 4865
rect 20234 4851 20248 4865
rect 20978 4851 20992 4865
rect 2762 4827 2776 4841
rect 9938 4827 9952 4841
rect 12986 4827 13000 4841
rect 13106 4827 13120 4841
rect 19562 4827 19576 4841
rect 20042 4827 20056 4841
rect 20834 4827 20848 4841
rect 2738 4803 2752 4817
rect 10802 4803 10816 4817
rect 10874 4803 10888 4817
rect 26869 4803 26883 4817
rect 2690 4779 2704 4793
rect 3290 4779 3304 4793
rect 3674 4779 3688 4793
rect 4466 4779 4480 4793
rect 5186 4779 5200 4793
rect 7682 4779 7696 4793
rect 7874 4779 7888 4793
rect 7970 4779 7984 4793
rect 8618 4779 8632 4793
rect 13418 4779 13432 4793
rect 15506 4779 15520 4793
rect 20546 4779 20560 4793
rect 23258 4779 23272 4793
rect 25274 4779 25288 4793
rect 2666 4755 2680 4769
rect 25010 4755 25024 4769
rect 25082 4755 25096 4769
rect 25322 4755 25336 4769
rect 2618 4731 2632 4745
rect 10250 4731 10264 4745
rect 10538 4731 10552 4745
rect 12458 4731 12472 4745
rect 23042 4731 23056 4745
rect 23282 4731 23296 4745
rect 23318 4731 23332 4745
rect 23666 4731 23680 4745
rect 25730 4731 25744 4745
rect 2594 4707 2608 4721
rect 5354 4707 5368 4721
rect 10130 4707 10144 4721
rect 11162 4707 11176 4721
rect 20594 4707 20608 4721
rect 22586 4707 22600 4721
rect 22874 4707 22888 4721
rect 23522 4707 23536 4721
rect 23834 4707 23848 4721
rect 25058 4707 25072 4721
rect 25226 4707 25240 4721
rect 2570 4683 2584 4697
rect 3266 4683 3280 4697
rect 3314 4683 3328 4697
rect 19130 4683 19144 4697
rect 26018 4683 26032 4697
rect 2546 4659 2560 4673
rect 13130 4659 13144 4673
rect 13274 4659 13288 4673
rect 14210 4659 14224 4673
rect 14258 4659 14272 4673
rect 19346 4659 19360 4673
rect 19634 4659 19648 4673
rect 24326 4659 24340 4673
rect 24986 4659 25000 4673
rect 25130 4659 25144 4673
rect 25202 4659 25216 4673
rect 25442 4659 25456 4673
rect 25778 4659 25792 4673
rect 26378 4659 26392 4673
rect 2522 4635 2536 4649
rect 8954 4635 8968 4649
rect 9026 4635 9040 4649
rect 25490 4635 25504 4649
rect 2474 4611 2488 4625
rect 11234 4611 11248 4625
rect 17186 4611 17200 4625
rect 19706 4611 19720 4625
rect 21050 4611 21064 4625
rect 22214 4611 22228 4625
rect 22562 4611 22576 4625
rect 24002 4611 24016 4625
rect 24266 4611 24280 4625
rect 24350 4611 24364 4625
rect 25010 4611 25024 4625
rect 25466 4611 25480 4625
rect 2426 4587 2440 4601
rect 3938 4587 3952 4601
rect 3986 4587 4000 4601
rect 14666 4587 14680 4601
rect 14738 4587 14752 4601
rect 24818 4587 24832 4601
rect 25370 4587 25384 4601
rect 25850 4587 25864 4601
rect 2402 4563 2416 4577
rect 2906 4563 2920 4577
rect 4274 4563 4288 4577
rect 9914 4563 9928 4577
rect 10898 4563 10912 4577
rect 14042 4563 14056 4577
rect 22658 4563 22672 4577
rect 22874 4563 22888 4577
rect 23546 4563 23560 4577
rect 2378 4539 2392 4553
rect 7946 4539 7960 4553
rect 22514 4539 22528 4553
rect 2330 4515 2344 4529
rect 3338 4515 3352 4529
rect 19802 4515 19816 4529
rect 22058 4515 22072 4529
rect 22538 4515 22552 4529
rect 2306 4491 2320 4505
rect 3578 4491 3592 4505
rect 6026 4491 6040 4505
rect 7754 4491 7768 4505
rect 10706 4491 10720 4505
rect 12674 4491 12688 4505
rect 13874 4491 13888 4505
rect 14282 4491 14296 4505
rect 14882 4491 14896 4505
rect 15722 4491 15736 4505
rect 16682 4491 16696 4505
rect 19538 4491 19552 4505
rect 21530 4491 21544 4505
rect 22010 4491 22024 4505
rect 22082 4491 22096 4505
rect 26306 4491 26320 4505
rect 2282 4467 2296 4481
rect 4394 4467 4408 4481
rect 7154 4467 7168 4481
rect 7466 4467 7480 4481
rect 8306 4467 8320 4481
rect 20810 4467 20824 4481
rect 21770 4467 21784 4481
rect 23282 4467 23296 4481
rect 2282 4443 2296 4457
rect 19610 4443 19624 4457
rect 21530 4443 21544 4457
rect 21746 4443 21760 4457
rect 22010 4443 22024 4457
rect 23102 4443 23116 4457
rect 2210 4419 2224 4433
rect 2978 4419 2992 4433
rect 3242 4419 3256 4433
rect 3890 4419 3904 4433
rect 4634 4419 4648 4433
rect 9314 4419 9328 4433
rect 13298 4419 13312 4433
rect 17882 4419 17896 4433
rect 19946 4419 19960 4433
rect 20762 4419 20776 4433
rect 2162 4395 2176 4409
rect 13274 4395 13288 4409
rect 14162 4395 14176 4409
rect 19490 4395 19504 4409
rect 22706 4395 22720 4409
rect 2114 4371 2128 4385
rect 19418 4371 19432 4385
rect 19538 4371 19552 4385
rect 19898 4371 19912 4385
rect 2090 4347 2104 4361
rect 2234 4347 2248 4361
rect 2354 4347 2368 4361
rect 5930 4347 5944 4361
rect 6602 4347 6616 4361
rect 9458 4347 9472 4361
rect 10274 4347 10288 4361
rect 12362 4347 12376 4361
rect 12914 4347 12928 4361
rect 13178 4347 13192 4361
rect 16922 4347 16936 4361
rect 17978 4347 17992 4361
rect 20498 4347 20512 4361
rect 25082 4347 25096 4361
rect 2066 4323 2080 4337
rect 19874 4323 19888 4337
rect 2018 4299 2032 4313
rect 6530 4299 6544 4313
rect 6578 4299 6592 4313
rect 18314 4299 18328 4313
rect 18698 4299 18712 4313
rect 21074 4299 21088 4313
rect 21650 4299 21664 4313
rect 1970 4275 1984 4289
rect 3554 4275 3568 4289
rect 4610 4275 4624 4289
rect 5162 4275 5176 4289
rect 7322 4275 7336 4289
rect 10562 4275 10576 4289
rect 10634 4275 10648 4289
rect 23066 4275 23080 4289
rect 1922 4251 1936 4265
rect 9794 4251 9808 4265
rect 9890 4251 9904 4265
rect 21914 4251 21928 4265
rect 1874 4227 1888 4241
rect 4370 4227 4384 4241
rect 9098 4227 9112 4241
rect 16994 4227 17008 4241
rect 17258 4227 17272 4241
rect 23138 4227 23152 4241
rect 1826 4203 1840 4217
rect 10466 4203 10480 4217
rect 18050 4203 18064 4217
rect 25754 4203 25768 4217
rect 1778 4179 1792 4193
rect 5042 4179 5056 4193
rect 6770 4179 6784 4193
rect 15386 4179 15400 4193
rect 15578 4179 15592 4193
rect 24602 4179 24616 4193
rect 1754 4155 1768 4169
rect 3482 4155 3496 4169
rect 10682 4155 10696 4169
rect 15554 4155 15568 4169
rect 15650 4155 15664 4169
rect 17858 4155 17872 4169
rect 18746 4155 18760 4169
rect 19322 4155 19336 4169
rect 1706 4131 1720 4145
rect 9218 4131 9232 4145
rect 9290 4131 9304 4145
rect 11378 4131 11392 4145
rect 15746 4131 15760 4145
rect 17114 4131 17128 4145
rect 19250 4131 19264 4145
rect 21866 4131 21880 4145
rect 22154 4131 22168 4145
rect 25250 4131 25264 4145
rect 1682 4107 1696 4121
rect 2258 4107 2272 4121
rect 4058 4107 4072 4121
rect 8738 4107 8752 4121
rect 13586 4107 13600 4121
rect 18074 4107 18088 4121
rect 19754 4107 19768 4121
rect 21890 4107 21904 4121
rect 25802 4107 25816 4121
rect 1658 4083 1672 4097
rect 7082 4083 7096 4097
rect 9218 4083 9232 4097
rect 11690 4083 11704 4097
rect 21122 4083 21136 4097
rect 21482 4083 21496 4097
rect 21890 4083 21904 4097
rect 22490 4083 22504 4097
rect 1634 4059 1648 4073
rect 7058 4059 7072 4073
rect 8066 4059 8080 4073
rect 8186 4059 8200 4073
rect 8378 4059 8392 4073
rect 11402 4059 11416 4073
rect 11522 4059 11536 4073
rect 11666 4059 11680 4073
rect 12194 4059 12208 4073
rect 20330 4059 20344 4073
rect 25898 4059 25912 4073
rect 1610 4035 1624 4049
rect 1898 4035 1912 4049
rect 4586 4035 4600 4049
rect 8402 4035 8416 4049
rect 12650 4035 12664 4049
rect 18194 4035 18208 4049
rect 21386 4035 21400 4049
rect 70 4011 84 4025
rect 10010 4011 10024 4025
rect 13658 4011 13672 4025
rect 17090 4011 17104 4025
rect 21506 4011 21520 4025
rect 70 3987 84 4001
rect 25418 3987 25432 4001
rect 1682 3963 1696 3977
rect 19466 3963 19480 3977
rect 19754 3963 19768 3977
rect 20210 3963 20224 3977
rect 1994 3939 2008 3953
rect 26450 3939 26464 3953
rect 2042 3915 2056 3929
rect 4826 3915 4840 3929
rect 5498 3915 5512 3929
rect 12578 3915 12592 3929
rect 13946 3915 13960 3929
rect 14090 3915 14104 3929
rect 15602 3915 15616 3929
rect 18818 3915 18832 3929
rect 21602 3915 21616 3929
rect 26090 3915 26104 3929
rect 2498 3891 2512 3905
rect 23090 3891 23104 3905
rect 2594 3867 2608 3881
rect 10970 3867 10984 3881
rect 16802 3867 16816 3881
rect 16898 3867 16912 3881
rect 19274 3867 19288 3881
rect 19778 3867 19792 3881
rect 2618 3843 2632 3857
rect 4874 3843 4888 3857
rect 19202 3843 19216 3857
rect 24242 3843 24256 3857
rect 2690 3819 2704 3833
rect 13538 3819 13552 3833
rect 19658 3819 19672 3833
rect 2714 3795 2728 3809
rect 4202 3795 4216 3809
rect 4250 3795 4264 3809
rect 22466 3795 22480 3809
rect 2930 3771 2944 3785
rect 20042 3771 20056 3785
rect 3218 3747 3232 3761
rect 13898 3747 13912 3761
rect 14042 3747 14056 3761
rect 14342 3747 14356 3761
rect 14522 3747 14536 3761
rect 18962 3747 18976 3761
rect 19010 3747 19024 3761
rect 19346 3747 19360 3761
rect 22106 3747 22120 3761
rect 22442 3747 22456 3761
rect 24386 3747 24400 3761
rect 3242 3723 3256 3737
rect 3290 3723 3304 3737
rect 3386 3723 3400 3737
rect 16754 3723 16768 3737
rect 22346 3723 22360 3737
rect 3290 3699 3304 3713
rect 5402 3699 5416 3713
rect 7202 3699 7216 3713
rect 7730 3699 7744 3713
rect 11546 3699 11560 3713
rect 14210 3699 14224 3713
rect 17858 3699 17872 3713
rect 20882 3699 20896 3713
rect 22610 3699 22624 3713
rect 22946 3699 22960 3713
rect 25658 3699 25672 3713
rect 3434 3675 3448 3689
rect 5090 3675 5104 3689
rect 6098 3675 6112 3689
rect 6794 3675 6808 3689
rect 15410 3675 15424 3689
rect 24626 3675 24640 3689
rect 3506 3651 3520 3665
rect 19370 3651 19384 3665
rect 19466 3651 19480 3665
rect 19682 3651 19696 3665
rect 22610 3651 22624 3665
rect 23234 3651 23248 3665
rect 3674 3627 3688 3641
rect 9530 3627 9544 3641
rect 18410 3627 18424 3641
rect 20618 3627 20632 3641
rect 22946 3627 22960 3641
rect 23582 3627 23596 3641
rect 3722 3603 3736 3617
rect 24050 3603 24064 3617
rect 3770 3579 3784 3593
rect 19082 3579 19096 3593
rect 19202 3579 19216 3593
rect 20858 3579 20872 3593
rect 3794 3555 3808 3569
rect 8522 3555 8536 3569
rect 18818 3555 18832 3569
rect 25058 3555 25072 3569
rect 3842 3531 3856 3545
rect 25706 3531 25720 3545
rect 3914 3507 3928 3521
rect 4298 3507 4312 3521
rect 6074 3507 6088 3521
rect 8210 3507 8224 3521
rect 10346 3507 10360 3521
rect 11906 3507 11920 3521
rect 13202 3507 13216 3521
rect 15314 3507 15328 3521
rect 17330 3507 17344 3521
rect 22466 3507 22480 3521
rect 24074 3507 24088 3521
rect 3938 3483 3952 3497
rect 21098 3483 21112 3497
rect 24074 3483 24088 3497
rect 24098 3483 24112 3497
rect 4106 3459 4120 3473
rect 8138 3459 8152 3473
rect 21986 3459 22000 3473
rect 22754 3459 22768 3473
rect 23186 3459 23200 3473
rect 24986 3459 25000 3473
rect 25754 3459 25768 3473
rect 4298 3435 4312 3449
rect 6914 3435 6928 3449
rect 7298 3435 7312 3449
rect 11594 3435 11608 3449
rect 13010 3435 13024 3449
rect 20930 3435 20944 3449
rect 24530 3435 24544 3449
rect 24746 3435 24760 3449
rect 25250 3435 25264 3449
rect 25682 3435 25696 3449
rect 4322 3411 4336 3425
rect 8714 3411 8728 3425
rect 10178 3411 10192 3425
rect 13970 3411 13984 3425
rect 14906 3411 14920 3425
rect 15890 3411 15904 3425
rect 17018 3411 17032 3425
rect 17354 3411 17368 3425
rect 21794 3411 21808 3425
rect 22274 3411 22288 3425
rect 25130 3411 25144 3425
rect 25682 3411 25696 3425
rect 26042 3411 26056 3425
rect 4394 3387 4408 3401
rect 6242 3387 6256 3401
rect 14330 3387 14344 3401
rect 17426 3387 17440 3401
rect 18266 3387 18280 3401
rect 18842 3387 18856 3401
rect 18890 3387 18904 3401
rect 22754 3387 22768 3401
rect 23474 3387 23488 3401
rect 4490 3363 4504 3377
rect 6458 3363 6472 3377
rect 15530 3363 15544 3377
rect 19274 3363 19288 3377
rect 4706 3339 4720 3353
rect 11930 3339 11944 3353
rect 19514 3339 19528 3353
rect 4754 3315 4768 3329
rect 7778 3315 7792 3329
rect 8258 3315 8272 3329
rect 13346 3315 13360 3329
rect 26258 3315 26272 3329
rect 4826 3291 4840 3305
rect 6386 3291 6400 3305
rect 9962 3291 9976 3305
rect 14942 3291 14956 3305
rect 18938 3291 18952 3305
rect 4874 3267 4888 3281
rect 5066 3267 5080 3281
rect 5138 3267 5152 3281
rect 22202 3267 22216 3281
rect 4946 3243 4960 3257
rect 9386 3243 9400 3257
rect 11882 3243 11896 3257
rect 12770 3243 12784 3257
rect 15626 3243 15640 3257
rect 15938 3243 15952 3257
rect 19034 3243 19048 3257
rect 4970 3219 4984 3233
rect 7802 3219 7816 3233
rect 9746 3219 9760 3233
rect 10610 3219 10624 3233
rect 11810 3219 11824 3233
rect 13370 3219 13384 3233
rect 14810 3219 14824 3233
rect 15818 3219 15832 3233
rect 16778 3219 16792 3233
rect 20258 3219 20272 3233
rect 23318 3219 23332 3233
rect 4994 3195 5008 3209
rect 11210 3195 11224 3209
rect 14114 3195 14128 3209
rect 14690 3195 14704 3209
rect 23210 3195 23224 3209
rect 5066 3171 5080 3185
rect 21314 3171 21328 3185
rect 21698 3171 21712 3185
rect 23210 3171 23224 3185
rect 26426 3171 26440 3185
rect 5162 3147 5176 3161
rect 5210 3147 5224 3161
rect 5258 3147 5272 3161
rect 7106 3147 7120 3161
rect 7226 3147 7240 3161
rect 7994 3147 8008 3161
rect 8090 3147 8104 3161
rect 12626 3147 12640 3161
rect 15698 3147 15712 3161
rect 23378 3147 23392 3161
rect 25154 3147 25168 3161
rect 5210 3123 5224 3137
rect 20834 3123 20848 3137
rect 5282 3099 5296 3113
rect 8786 3099 8800 3113
rect 8834 3099 8848 3113
rect 26114 3099 26128 3113
rect 5354 3075 5368 3089
rect 10418 3075 10432 3089
rect 10610 3075 10624 3089
rect 14450 3075 14464 3089
rect 15098 3075 15112 3089
rect 18866 3075 18880 3089
rect 20186 3075 20200 3089
rect 5474 3051 5488 3065
rect 6266 3051 6280 3065
rect 6314 3051 6328 3065
rect 21194 3051 21208 3065
rect 5642 3027 5656 3041
rect 23258 3027 23272 3041
rect 5834 3003 5848 3017
rect 9986 3003 10000 3017
rect 10034 3003 10048 3017
rect 23786 3003 23800 3017
rect 5834 2979 5848 2993
rect 25178 2979 25192 2993
rect 5882 2955 5896 2969
rect 12938 2955 12952 2969
rect 26186 2955 26200 2969
rect 5906 2931 5920 2945
rect 8018 2931 8032 2945
rect 8114 2931 8128 2945
rect 17834 2931 17848 2945
rect 21026 2931 21040 2945
rect 21626 2931 21640 2945
rect 23786 2931 23800 2945
rect 25178 2931 25192 2945
rect 6122 2907 6136 2921
rect 13994 2907 14008 2921
rect 16586 2907 16600 2921
rect 22826 2907 22840 2921
rect 23162 2907 23176 2921
rect 6458 2883 6472 2897
rect 11114 2883 11128 2897
rect 14138 2883 14152 2897
rect 15482 2883 15496 2897
rect 16706 2883 16720 2897
rect 16874 2883 16888 2897
rect 24914 2883 24928 2897
rect 6578 2859 6592 2873
rect 8474 2859 8488 2873
rect 25922 2859 25936 2873
rect 6722 2835 6736 2849
rect 16754 2835 16768 2849
rect 16802 2835 16816 2849
rect 16826 2835 16840 2849
rect 17570 2835 17584 2849
rect 25034 2835 25048 2849
rect 6866 2811 6880 2825
rect 6938 2811 6952 2825
rect 14234 2811 14248 2825
rect 15698 2811 15712 2825
rect 19730 2811 19744 2825
rect 25538 2811 25552 2825
rect 7106 2787 7120 2801
rect 8090 2787 8104 2801
rect 10154 2787 10168 2801
rect 10298 2787 10312 2801
rect 11714 2787 11728 2801
rect 16658 2787 16672 2801
rect 20234 2787 20248 2801
rect 23162 2787 23176 2801
rect 23642 2787 23656 2801
rect 7130 2763 7144 2777
rect 9002 2763 9016 2777
rect 9050 2763 9064 2777
rect 23618 2763 23632 2777
rect 7226 2739 7240 2753
rect 16634 2739 16648 2753
rect 16778 2739 16792 2753
rect 25826 2739 25840 2753
rect 7274 2715 7288 2729
rect 9554 2715 9568 2729
rect 9866 2715 9880 2729
rect 19922 2715 19936 2729
rect 20474 2715 20488 2729
rect 20906 2715 20920 2729
rect 21578 2715 21592 2729
rect 22034 2715 22048 2729
rect 25226 2715 25240 2729
rect 7322 2691 7336 2705
rect 19394 2691 19408 2705
rect 19730 2691 19744 2705
rect 19982 2691 19996 2705
rect 20186 2691 20200 2705
rect 20282 2691 20296 2705
rect 7346 2667 7360 2681
rect 7490 2667 7504 2681
rect 7538 2667 7552 2681
rect 9842 2667 9856 2681
rect 9890 2667 9904 2681
rect 13466 2667 13480 2681
rect 13562 2667 13576 2681
rect 14306 2667 14320 2681
rect 15146 2667 15160 2681
rect 20018 2667 20032 2681
rect 24098 2667 24112 2681
rect 7370 2643 7384 2657
rect 7706 2643 7720 2657
rect 25322 2643 25336 2657
rect 7874 2619 7888 2633
rect 7922 2619 7936 2633
rect 7994 2619 8008 2633
rect 8330 2619 8344 2633
rect 23042 2619 23056 2633
rect 7922 2595 7936 2609
rect 20714 2595 20728 2609
rect 8186 2571 8200 2585
rect 8234 2571 8248 2585
rect 8282 2571 8296 2585
rect 12338 2571 12352 2585
rect 24122 2571 24136 2585
rect 8330 2547 8344 2561
rect 17066 2547 17080 2561
rect 17618 2547 17632 2561
rect 21842 2547 21856 2561
rect 24122 2547 24136 2561
rect 24146 2547 24160 2561
rect 8378 2523 8392 2537
rect 10586 2523 10600 2537
rect 14930 2523 14944 2537
rect 15194 2523 15208 2537
rect 22178 2523 22192 2537
rect 8522 2499 8536 2513
rect 15770 2499 15784 2513
rect 18362 2499 18376 2513
rect 22370 2499 22384 2513
rect 8666 2475 8680 2489
rect 20306 2475 20320 2489
rect 20714 2475 20728 2489
rect 21074 2475 21088 2489
rect 22370 2475 22384 2489
rect 23018 2475 23032 2489
rect 8834 2451 8848 2465
rect 9146 2451 9160 2465
rect 9338 2451 9352 2465
rect 11786 2451 11800 2465
rect 11834 2451 11848 2465
rect 14594 2451 14608 2465
rect 15242 2451 15256 2465
rect 16226 2451 16240 2465
rect 16514 2451 16528 2465
rect 16946 2451 16960 2465
rect 17786 2451 17800 2465
rect 19442 2451 19456 2465
rect 9170 2427 9184 2441
rect 18002 2427 18016 2441
rect 19298 2427 19312 2441
rect 9434 2403 9448 2417
rect 9482 2403 9496 2417
rect 9602 2403 9616 2417
rect 12578 2403 12592 2417
rect 12698 2403 12712 2417
rect 20426 2403 20440 2417
rect 9650 2379 9664 2393
rect 13994 2379 14008 2393
rect 14066 2379 14080 2393
rect 14378 2379 14392 2393
rect 14546 2379 14560 2393
rect 15554 2379 15568 2393
rect 16442 2379 16456 2393
rect 16562 2379 16576 2393
rect 25946 2379 25960 2393
rect 9674 2355 9688 2369
rect 11186 2355 11200 2369
rect 11234 2355 11248 2369
rect 16730 2355 16744 2369
rect 18938 2355 18952 2369
rect 18986 2355 19000 2369
rect 9794 2331 9808 2345
rect 9914 2331 9928 2345
rect 10178 2331 10192 2345
rect 10322 2331 10336 2345
rect 10658 2331 10672 2345
rect 10850 2331 10864 2345
rect 20570 2331 20584 2345
rect 23426 2331 23440 2345
rect 10298 2307 10312 2321
rect 10370 2307 10384 2321
rect 10706 2307 10720 2321
rect 19058 2307 19072 2321
rect 10730 2283 10744 2297
rect 15290 2283 15304 2297
rect 10802 2259 10816 2273
rect 24554 2259 24568 2273
rect 10826 2235 10840 2249
rect 10946 2235 10960 2249
rect 10994 2235 11008 2249
rect 13850 2235 13864 2249
rect 24938 2235 24952 2249
rect 10874 2211 10888 2225
rect 11450 2211 11464 2225
rect 14018 2211 14032 2225
rect 11018 2187 11032 2201
rect 18482 2187 18496 2201
rect 22802 2187 22816 2201
rect 24290 2187 24304 2201
rect 24866 2187 24880 2201
rect 11090 2163 11104 2177
rect 26426 2163 26440 2177
rect 11138 2139 11152 2153
rect 12194 2139 12208 2153
rect 23930 2139 23944 2153
rect 11186 2115 11200 2129
rect 20978 2115 20992 2129
rect 11210 2091 11224 2105
rect 16298 2091 16312 2105
rect 23978 2091 23992 2105
rect 11306 2067 11320 2081
rect 12506 2067 12520 2081
rect 17714 2067 17728 2081
rect 23978 2067 23992 2081
rect 24098 2067 24112 2081
rect 11330 2043 11344 2057
rect 13682 2043 13696 2057
rect 13778 2043 13792 2057
rect 14474 2043 14488 2057
rect 11546 2019 11560 2033
rect 17042 2019 17056 2033
rect 20378 2019 20392 2033
rect 11738 1995 11752 2009
rect 16442 1995 16456 2009
rect 12242 1971 12256 1985
rect 13442 1971 13456 1985
rect 12338 1947 12352 1961
rect 13034 1947 13048 1961
rect 13106 1947 13120 1961
rect 16370 1947 16384 1961
rect 12554 1923 12568 1937
rect 12602 1923 12616 1937
rect 12794 1923 12808 1937
rect 21002 1923 21016 1937
rect 12842 1899 12856 1913
rect 17930 1899 17944 1913
rect 12890 1875 12904 1889
rect 16394 1875 16408 1889
rect 12986 1851 13000 1865
rect 13322 1851 13336 1865
rect 13394 1851 13408 1865
rect 24410 1851 24424 1865
rect 26426 1851 26440 1865
rect 26869 1851 26883 1865
rect 13178 1827 13192 1841
rect 13754 1827 13768 1841
rect 26474 1827 26488 1841
rect 26869 1827 26883 1841
rect 13202 1803 13216 1817
rect 13814 1803 13828 1817
rect 26450 1803 26464 1817
rect 26869 1803 26883 1817
rect 16586 970 16600 984
rect 18866 970 18880 984
rect 15890 946 15904 960
rect 18434 946 18448 960
rect 15338 922 15352 936
rect 17546 922 17560 936
rect 13850 898 13864 912
rect 23306 898 23320 912
rect 11042 874 11056 888
rect 25490 874 25504 888
rect 10946 850 10960 864
rect 25562 850 25576 864
rect 10778 826 10792 840
rect 14114 826 14128 840
rect 14474 826 14488 840
rect 16850 826 16864 840
rect 16946 826 16960 840
rect 22898 826 22912 840
rect 10442 802 10456 816
rect 15218 802 15232 816
rect 19298 802 19312 816
rect 10394 778 10408 792
rect 22178 778 22192 792
rect 10370 754 10384 768
rect 20282 754 20296 768
rect 9482 730 9496 744
rect 20666 730 20680 744
rect 9050 706 9064 720
rect 17642 706 17656 720
rect 22802 706 22816 720
rect 9002 682 9016 696
rect 23426 682 23440 696
rect 8954 658 8968 672
rect 20618 658 20632 672
rect 8738 634 8752 648
rect 19970 634 19984 648
rect 8714 610 8728 624
rect 25394 610 25408 624
rect 8642 586 8656 600
rect 17138 586 17152 600
rect 17450 586 17464 600
rect 18962 586 18976 600
rect 19946 586 19960 600
rect 8162 562 8176 576
rect 19634 562 19648 576
rect 7826 538 7840 552
rect 20018 538 20032 552
rect 7610 514 7624 528
rect 24386 514 24400 528
rect 7562 490 7576 504
rect 8210 490 8224 504
rect 8570 490 8584 504
rect 21002 490 21016 504
rect 22994 490 23008 504
rect 7538 466 7552 480
rect 12386 466 12400 480
rect 13034 466 13048 480
rect 22298 466 22312 480
rect 7178 442 7192 456
rect 18578 442 18592 456
rect 21626 442 21640 456
rect 6698 418 6712 432
rect 19418 418 19432 432
rect 6650 394 6664 408
rect 6722 394 6736 408
rect 7034 394 7048 408
rect 21818 394 21832 408
rect 6170 370 6184 384
rect 8426 370 8440 384
rect 11402 370 11416 384
rect 13298 370 13312 384
rect 24146 370 24160 384
rect 6074 346 6088 360
rect 23138 346 23152 360
rect 5282 322 5296 336
rect 6770 322 6784 336
rect 6818 322 6832 336
rect 13466 322 13480 336
rect 20834 322 20848 336
rect 5114 298 5128 312
rect 16826 298 16840 312
rect 3842 274 3856 288
rect 14978 274 14992 288
rect 15050 274 15064 288
rect 25442 274 25456 288
rect 3722 250 3736 264
rect 6026 250 6040 264
rect 21146 250 21160 264
rect 2642 226 2656 240
rect 20570 226 20584 240
rect 2570 202 2584 216
rect 22394 202 22408 216
rect 2378 178 2392 192
rect 3986 178 4000 192
rect 4130 178 4144 192
rect 11666 178 11680 192
rect 13586 178 13600 192
rect 24002 178 24016 192
rect 2330 154 2344 168
rect 4346 154 4360 168
rect 4418 154 4432 168
rect 4634 154 4648 168
rect 25610 154 25624 168
rect 70 130 84 144
rect 12602 130 12616 144
rect 13682 130 13696 144
rect 21770 130 21784 144
rect 70 106 84 120
rect 2426 106 2440 120
rect 2474 106 2488 120
rect 18026 106 18040 120
rect 6266 82 6280 96
rect 7814 82 7828 96
rect 8114 82 8128 96
rect 9554 82 9568 96
rect 10346 82 10360 96
rect 14210 82 14224 96
rect 15002 82 15016 96
rect 17042 82 17056 96
rect 25562 82 25576 96
rect 26869 82 26883 96
rect 7490 58 7504 72
rect 25562 58 25576 72
rect 25586 58 25600 72
rect 26869 58 26883 72
rect 10586 34 10600 48
rect 25586 34 25600 48
rect 25610 34 25624 48
rect 26869 34 26883 48
rect 11306 10 11320 24
rect 26869 10 26883 24
<< metal2 >>
rect 0 8469 70 8481
rect 0 8445 70 8457
rect 123 8314 323 8588
rect 339 8314 351 8588
rect 363 8314 375 8588
rect 387 8314 399 8588
rect 411 8314 423 8588
rect 2319 8506 2331 8588
rect 3219 8506 3231 8588
rect 2320 8492 2338 8506
rect 2307 8314 2319 8492
rect 4047 8434 4059 8588
rect 4875 8506 4887 8588
rect 4059 8314 4071 8396
rect 4299 8314 4311 8492
rect 5043 8314 5055 8516
rect 5307 8314 5319 8540
rect 5703 8386 5715 8588
rect 5739 8410 5751 8588
rect 6807 8578 6819 8588
rect 6808 8564 6826 8578
rect 5715 8314 5727 8348
rect 6387 8314 6399 8396
rect 6459 8314 6471 8420
rect 6771 8314 6783 8420
rect 6795 8314 6807 8564
rect 7395 8434 7407 8588
rect 9015 8578 9027 8588
rect 8715 8314 8727 8372
rect 9243 8314 9255 8420
rect 9519 8386 9531 8588
rect 10431 8458 10443 8588
rect 10432 8444 10450 8458
rect 9520 8372 9538 8386
rect 9507 8314 9519 8372
rect 10371 8314 10383 8444
rect 10419 8314 10431 8444
rect 10611 8314 10623 8492
rect 11199 8482 11211 8588
rect 11200 8468 11218 8482
rect 10923 8314 10935 8468
rect 11187 8314 11199 8468
rect 11535 8434 11547 8588
rect 13155 8506 13167 8588
rect 13191 8530 13203 8588
rect 12483 8314 12495 8468
rect 13947 8314 13959 8492
rect 14007 8410 14019 8588
rect 15615 8506 15627 8588
rect 16239 8458 16251 8588
rect 16455 8554 16467 8588
rect 17271 8458 17283 8588
rect 18879 8530 18891 8588
rect 16240 8444 16258 8458
rect 14691 8314 14703 8348
rect 16227 8314 16239 8444
rect 16947 8314 16959 8444
rect 18531 8314 18543 8444
rect 18963 8314 18975 8492
rect 19131 8314 19143 8564
rect 19695 8506 19707 8588
rect 20295 8434 20307 8588
rect 21327 8554 21339 8588
rect 22143 8578 22155 8588
rect 20296 8420 20314 8434
rect 20283 8314 20295 8420
rect 21315 8314 21327 8420
rect 21459 8314 21471 8396
rect 21723 8314 21735 8372
rect 22167 8362 22179 8588
rect 23775 8530 23787 8588
rect 22683 8314 22695 8324
rect 23211 8314 23223 8516
rect 23799 8482 23811 8588
rect 24339 8314 24351 8540
rect 24615 8434 24627 8588
rect 24867 8314 24879 8564
rect 25431 8386 25443 8588
rect 25155 8314 25167 8348
rect 25467 8314 25479 8492
rect 26187 8314 26199 8516
rect 26379 8314 26391 8420
rect 26427 8314 26439 8372
rect 26451 8362 26463 8420
rect 26475 8410 26487 8420
rect 26499 8386 26511 8396
rect 26523 8338 26535 8372
rect 26547 8338 26559 8444
rect 26571 8314 26771 8588
rect 26883 8421 26953 8433
rect 26883 8397 26953 8409
rect 26883 8373 26953 8385
rect 26883 8349 26953 8361
rect 26883 8325 26953 8337
rect 0 4012 70 4024
rect 0 3988 70 4000
rect 123 1793 323 7515
rect 339 1793 351 7515
rect 363 1793 375 7515
rect 387 1793 399 7515
rect 411 1793 423 7515
rect 1611 4049 1623 7515
rect 1635 4073 1647 7515
rect 1659 4097 1671 7515
rect 1683 4121 1695 7515
rect 1707 4145 1719 7515
rect 1755 4169 1767 7515
rect 1779 4193 1791 7515
rect 1827 4217 1839 7515
rect 1875 4241 1887 7515
rect 1899 4049 1911 7515
rect 1923 4265 1935 7515
rect 1971 4289 1983 7515
rect 1683 1793 1695 3963
rect 1995 3953 2007 7515
rect 2019 4313 2031 7515
rect 2067 4337 2079 7515
rect 2091 4361 2103 7515
rect 2115 4385 2127 7515
rect 2163 4409 2175 7515
rect 2211 4433 2223 7515
rect 2283 4481 2295 7515
rect 2307 4505 2319 7515
rect 2331 4529 2343 7515
rect 2379 4553 2391 7515
rect 2403 4577 2415 7515
rect 2427 4601 2439 7515
rect 2475 4625 2487 7515
rect 2043 1793 2055 3915
rect 2091 1793 2103 4347
rect 2235 1793 2247 4347
rect 2259 1793 2271 4107
rect 2283 1793 2295 4443
rect 2355 1793 2367 4347
rect 2499 3905 2511 7515
rect 2523 4649 2535 7515
rect 2571 4697 2583 7515
rect 2595 4721 2607 7515
rect 2619 4745 2631 7515
rect 2667 4769 2679 7515
rect 2691 4793 2703 7515
rect 2547 1793 2559 4659
rect 2595 1793 2607 3867
rect 2619 1793 2631 3843
rect 2691 1793 2703 3819
rect 2715 3809 2727 7515
rect 2763 4841 2775 7515
rect 2811 4865 2823 7515
rect 2883 4913 2895 7515
rect 2739 1793 2751 4803
rect 2883 1793 2895 4875
rect 2907 4577 2919 7515
rect 2931 3785 2943 7515
rect 2979 4433 2991 7515
rect 3003 4937 3015 7515
rect 3027 4961 3039 7515
rect 3051 4985 3063 7515
rect 3075 5009 3087 7515
rect 3123 5033 3135 7515
rect 3147 5057 3159 7515
rect 3171 5081 3183 7515
rect 3219 3761 3231 7515
rect 3243 4433 3255 7515
rect 3267 4697 3279 7515
rect 3291 3737 3303 4779
rect 3315 4697 3327 7515
rect 3339 4529 3351 7515
rect 3387 3737 3399 7515
rect 3435 5105 3447 7515
rect 3459 5129 3471 7515
rect 3243 1793 3255 3723
rect 3291 1793 3303 3699
rect 3435 1793 3447 3675
rect 3483 1793 3495 4155
rect 3507 3665 3519 7515
rect 3555 5153 3567 7515
rect 3579 4505 3591 7515
rect 3603 5201 3615 7515
rect 3555 1793 3567 4275
rect 3603 1793 3615 5163
rect 3651 4913 3663 7515
rect 3675 4793 3687 7515
rect 3699 5225 3711 7515
rect 3675 1793 3687 3627
rect 3723 3617 3735 7515
rect 3771 3593 3783 7515
rect 3795 5249 3807 7515
rect 3795 1793 3807 3555
rect 3819 1793 3831 5259
rect 3843 3545 3855 7515
rect 3891 5297 3903 7515
rect 3915 5321 3927 7515
rect 3939 4601 3951 7515
rect 3963 5345 3975 7515
rect 3987 4601 3999 7515
rect 4035 5417 4047 7515
rect 3891 1793 3903 4419
rect 3915 1793 3927 3507
rect 3939 1793 3951 3483
rect 4011 1793 4023 5355
rect 4035 1793 4047 5379
rect 4059 4121 4071 7515
rect 4107 5465 4119 7515
rect 4155 5489 4167 7515
rect 4203 5537 4215 7515
rect 4083 1793 4095 5427
rect 4107 1793 4119 3459
rect 4179 1793 4191 5499
rect 4203 1793 4215 3795
rect 4227 1793 4239 5547
rect 4275 4577 4287 7515
rect 4251 1793 4263 3795
rect 4299 3521 4311 7515
rect 4323 5585 4335 7515
rect 4371 4241 4383 7515
rect 4395 4481 4407 7515
rect 4419 5609 4431 7515
rect 4299 1793 4311 3435
rect 4323 1793 4335 3411
rect 4395 1793 4407 3387
rect 4443 1793 4455 5619
rect 4467 4793 4479 7515
rect 4491 5657 4503 7515
rect 4515 5681 4527 7515
rect 4563 5705 4575 7515
rect 4491 1793 4503 3363
rect 4539 1793 4551 5211
rect 4587 4049 4599 7515
rect 4611 4961 4623 7515
rect 4635 4433 4647 7515
rect 4659 5753 4671 7515
rect 4707 5777 4719 7515
rect 4611 1793 4623 4275
rect 4659 1793 4671 5715
rect 4731 4961 4743 7515
rect 4755 5801 4767 7515
rect 4803 5825 4815 7515
rect 4827 3929 4839 7515
rect 4875 3857 4887 7515
rect 4923 5849 4935 7515
rect 4947 5873 4959 7515
rect 4995 5897 5007 7515
rect 5043 5921 5055 7515
rect 5091 5945 5103 7515
rect 5115 5921 5127 7515
rect 4707 1793 4719 3339
rect 4755 1793 4767 3315
rect 4827 1793 4839 3291
rect 4875 1793 4887 3267
rect 4947 1793 4959 3243
rect 4971 1793 4983 3219
rect 4995 1793 5007 3195
rect 5043 1793 5055 4179
rect 5067 3281 5079 5907
rect 5067 1793 5079 3171
rect 5091 1793 5103 3675
rect 5139 3281 5151 7515
rect 5163 4289 5175 7515
rect 5211 5969 5223 7515
rect 5235 5993 5247 7515
rect 5163 1793 5175 3147
rect 5187 1793 5199 4779
rect 5211 3161 5223 5859
rect 5259 5177 5271 7515
rect 5211 1793 5223 3123
rect 5259 1793 5271 3147
rect 5283 3113 5295 7515
rect 5307 1793 5319 5163
rect 5331 1793 5343 5739
rect 5355 4721 5367 7515
rect 5379 6017 5391 7515
rect 5403 3713 5415 7515
rect 5427 6041 5439 7515
rect 5475 6065 5487 7515
rect 5499 3929 5511 7515
rect 5547 4961 5559 7515
rect 5595 6089 5607 7515
rect 5619 5153 5631 7515
rect 5355 1793 5367 3075
rect 5475 1793 5487 3051
rect 5643 3041 5655 7515
rect 5691 6113 5703 7515
rect 5739 6137 5751 7515
rect 5787 6161 5799 7515
rect 5835 3017 5847 7515
rect 5835 1793 5847 2979
rect 5883 1793 5895 2955
rect 5907 2945 5919 7515
rect 5931 4361 5943 7515
rect 5955 6185 5967 7515
rect 6027 4505 6039 7515
rect 6051 6209 6063 7515
rect 6051 1793 6063 4947
rect 6075 3521 6087 6195
rect 6099 3689 6111 7515
rect 6123 4961 6135 7515
rect 6195 6233 6207 7515
rect 6219 6257 6231 7515
rect 6123 1793 6135 2907
rect 6147 1793 6159 6195
rect 6243 5969 6255 7515
rect 6195 1793 6207 5955
rect 6243 1793 6255 3387
rect 6267 3065 6279 7515
rect 6291 1793 6303 6267
rect 6315 3065 6327 7515
rect 6339 6305 6351 7515
rect 6363 6329 6375 7515
rect 6435 6329 6447 7515
rect 6339 1793 6351 5451
rect 6363 1793 6375 4971
rect 6387 3305 6399 6315
rect 6411 1793 6423 5139
rect 6459 3377 6471 7515
rect 6483 6353 6495 7515
rect 6459 1793 6471 2883
rect 6507 1793 6519 4899
rect 6531 4313 6543 7515
rect 6555 6137 6567 7515
rect 6579 4313 6591 7515
rect 6603 6137 6615 7515
rect 6651 6377 6663 7515
rect 6675 6401 6687 7515
rect 6699 6425 6711 7515
rect 6579 1793 6591 2859
rect 6603 1793 6615 4347
rect 6723 2849 6735 7515
rect 6771 4193 6783 7515
rect 6795 3689 6807 7515
rect 6843 4985 6855 7515
rect 6891 6449 6903 7515
rect 6915 3449 6927 7515
rect 6963 6473 6975 7515
rect 7011 6521 7023 7515
rect 7035 6545 7047 7515
rect 7059 6569 7071 7515
rect 7083 6593 7095 7515
rect 7131 6617 7143 7515
rect 6867 1793 6879 2811
rect 6939 1793 6951 2811
rect 6963 1793 6975 5451
rect 6987 1793 6999 6483
rect 7059 1793 7071 4059
rect 7083 1793 7095 4083
rect 7107 3161 7119 6579
rect 7155 4481 7167 7515
rect 7179 6593 7191 7515
rect 7107 1793 7119 2787
rect 7131 1793 7143 2763
rect 7203 1793 7215 3699
rect 7227 3161 7239 7515
rect 7251 6641 7263 7515
rect 7275 6665 7287 7515
rect 7323 4289 7335 7515
rect 7227 1793 7239 2739
rect 7275 1793 7287 2715
rect 7299 1793 7311 3435
rect 7323 1793 7335 2691
rect 7347 2681 7359 7515
rect 7371 6233 7383 7515
rect 7419 6233 7431 7515
rect 7371 1793 7383 2643
rect 7419 1793 7431 5811
rect 7467 4481 7479 7515
rect 7539 2681 7551 7515
rect 7587 6713 7599 7515
rect 7659 6737 7671 7515
rect 7683 6761 7695 7515
rect 7491 1793 7503 2667
rect 7587 1793 7599 6675
rect 7659 1793 7671 6075
rect 7707 5513 7719 7515
rect 7683 1793 7695 4779
rect 7731 3713 7743 6747
rect 7755 5513 7767 7515
rect 7779 5465 7791 7515
rect 7803 6761 7815 7515
rect 7851 6785 7863 7515
rect 7875 4793 7887 7515
rect 7899 6809 7911 7515
rect 7707 1793 7719 2643
rect 7755 1793 7767 4491
rect 7779 1793 7791 3315
rect 7803 1793 7815 3219
rect 7875 1793 7887 2619
rect 7899 1793 7911 5211
rect 7923 2633 7935 4923
rect 7947 4553 7959 7515
rect 7923 1793 7935 2595
rect 7971 1793 7983 4779
rect 7995 3161 8007 7515
rect 8067 6833 8079 7515
rect 7995 1793 8007 2619
rect 8019 1793 8031 2931
rect 8067 1793 8079 4059
rect 8091 3161 8103 7515
rect 8115 2945 8127 7515
rect 8139 3473 8151 7515
rect 8187 4073 8199 7515
rect 8211 3521 8223 7515
rect 8235 6857 8247 7515
rect 8091 1793 8103 2787
rect 8235 2585 8247 5811
rect 8283 5705 8295 7515
rect 8307 4481 8319 7515
rect 8187 1793 8199 2571
rect 8259 1793 8271 3315
rect 8331 2633 8343 7515
rect 8379 4073 8391 7515
rect 8403 4049 8415 7515
rect 8427 6881 8439 7515
rect 8475 2873 8487 7515
rect 8283 1793 8295 2571
rect 8331 1793 8343 2547
rect 8379 1793 8391 2523
rect 8499 1793 8511 6051
rect 8523 3569 8535 7515
rect 8595 5729 8607 7515
rect 8619 6905 8631 7515
rect 8643 5633 8655 7515
rect 8667 5729 8679 7515
rect 8523 1793 8535 2499
rect 8547 1793 8559 5451
rect 8619 1793 8631 4779
rect 8715 3425 8727 7515
rect 8739 4121 8751 7515
rect 8787 5633 8799 7515
rect 8835 3113 8847 7515
rect 8859 6353 8871 7515
rect 8907 6929 8919 7515
rect 8667 1793 8679 2475
rect 8787 1793 8799 3099
rect 8835 1793 8847 2451
rect 8859 1793 8871 4971
rect 8907 1793 8919 6339
rect 8955 4649 8967 7515
rect 8979 6977 8991 7515
rect 8979 1793 8991 6939
rect 9003 2777 9015 7515
rect 9027 4649 9039 7515
rect 9051 2777 9063 7515
rect 9099 6401 9111 7515
rect 9123 6377 9135 7515
rect 9099 1793 9111 4227
rect 9147 2465 9159 7515
rect 9195 6761 9207 7515
rect 9219 4145 9231 7515
rect 9291 5705 9303 7515
rect 9315 7001 9327 7515
rect 9171 1793 9183 2427
rect 9219 1793 9231 4083
rect 9291 1793 9303 4131
rect 9315 1793 9327 4419
rect 9339 2465 9351 7515
rect 9387 7025 9399 7515
rect 9363 1793 9375 6195
rect 9387 3257 9399 6987
rect 9435 6569 9447 7515
rect 9507 7001 9519 7515
rect 9411 1793 9423 5811
rect 9435 1793 9447 2403
rect 9459 1793 9471 4347
rect 9483 2417 9495 6771
rect 9531 1793 9543 3627
rect 9555 2729 9567 7515
rect 9579 7049 9591 7515
rect 9579 1793 9591 6771
rect 9603 2417 9615 7515
rect 9627 1793 9639 6747
rect 9651 2393 9663 7515
rect 9675 6521 9687 7515
rect 9699 5273 9711 7515
rect 9747 5273 9759 7515
rect 9771 6761 9783 7515
rect 9795 4265 9807 7515
rect 9819 5345 9831 7515
rect 9675 1793 9687 2355
rect 9747 1793 9759 3219
rect 9843 2681 9855 7515
rect 9891 4265 9903 7515
rect 9915 7073 9927 7515
rect 9939 7097 9951 7515
rect 9795 1793 9807 2331
rect 9867 1793 9879 2715
rect 9891 1793 9903 2667
rect 9915 2345 9927 4563
rect 9939 1793 9951 4827
rect 9963 3305 9975 7515
rect 9987 7121 9999 7515
rect 9987 1793 9999 3003
rect 10011 1793 10023 4011
rect 10035 3017 10047 7515
rect 10059 7145 10071 7515
rect 10107 7001 10119 7515
rect 10059 1793 10071 6987
rect 10107 1793 10119 5811
rect 10131 1793 10143 4707
rect 10155 2801 10167 7515
rect 10179 3425 10191 7515
rect 10203 6521 10215 7515
rect 10251 7169 10263 7515
rect 10179 1793 10191 2331
rect 10227 1793 10239 4851
rect 10251 1793 10263 4731
rect 10275 1793 10287 4347
rect 10299 2801 10311 7515
rect 10323 2345 10335 6051
rect 10347 3521 10359 7155
rect 10371 2321 10383 7515
rect 10419 3089 10431 7515
rect 10467 4217 10479 7515
rect 10491 7169 10503 7515
rect 10299 1793 10311 2307
rect 10491 1793 10503 6531
rect 10539 4745 10551 7515
rect 10563 1793 10575 4275
rect 10587 2537 10599 7515
rect 10611 3233 10623 7515
rect 10635 4289 10647 7515
rect 10683 4169 10695 7515
rect 10707 4505 10719 7515
rect 10611 1793 10623 3075
rect 10659 1793 10671 2331
rect 10707 1793 10719 2307
rect 10731 2297 10743 7515
rect 10779 6473 10791 7515
rect 10803 4817 10815 7515
rect 10827 7193 10839 7515
rect 10851 2345 10863 7515
rect 10875 4817 10887 7515
rect 10923 7217 10935 7515
rect 10803 1793 10815 2259
rect 10827 1793 10839 2235
rect 10875 1793 10887 2211
rect 10899 1793 10911 4563
rect 10923 1793 10935 5451
rect 10947 2249 10959 7203
rect 10971 3881 10983 7515
rect 10995 7217 11007 7515
rect 11019 5873 11031 7515
rect 11067 5873 11079 7515
rect 11091 7025 11103 7515
rect 10995 1793 11007 2235
rect 11019 1793 11031 2187
rect 11067 1793 11079 5739
rect 11115 2897 11127 7515
rect 11139 5753 11151 7515
rect 11091 1793 11103 2163
rect 11139 1793 11151 2139
rect 11163 1793 11175 4707
rect 11187 2369 11199 7515
rect 11211 3209 11223 5859
rect 11235 4625 11247 7515
rect 11259 5873 11271 7515
rect 11283 7241 11295 7515
rect 11187 1793 11199 2115
rect 11211 1793 11223 2091
rect 11235 1793 11247 2355
rect 11283 1793 11295 6099
rect 11331 6017 11343 7515
rect 11355 7265 11367 7515
rect 11307 1793 11319 2067
rect 11331 1793 11343 2043
rect 11379 1793 11391 4131
rect 11403 4073 11415 7515
rect 11451 7289 11463 7515
rect 11475 6185 11487 7515
rect 11499 7313 11511 7515
rect 11451 1793 11463 2211
rect 11499 1793 11511 5043
rect 11523 1793 11535 4059
rect 11547 3713 11559 7515
rect 11571 6185 11583 7515
rect 11547 1793 11559 2019
rect 11571 1793 11583 5283
rect 11595 3449 11607 7515
rect 11619 7145 11631 7515
rect 11619 1793 11631 5283
rect 11667 4073 11679 7515
rect 11691 4097 11703 7515
rect 11715 2801 11727 7515
rect 11739 2009 11751 7515
rect 11787 2465 11799 7515
rect 11811 3233 11823 7515
rect 11835 2465 11847 7515
rect 11883 3257 11895 7515
rect 11907 3521 11919 7515
rect 11931 3353 11943 7515
rect 11979 7337 11991 7515
rect 12003 7361 12015 7515
rect 12027 5321 12039 7515
rect 12075 6353 12087 7515
rect 12099 5321 12111 7515
rect 12147 6353 12159 7515
rect 12195 4073 12207 7515
rect 12195 1793 12207 2139
rect 12243 1985 12255 7515
rect 12315 6425 12327 7515
rect 12339 2585 12351 7515
rect 12387 5129 12399 7515
rect 12435 7385 12447 7515
rect 12339 1793 12351 1947
rect 12363 1793 12375 4347
rect 12435 1793 12447 5499
rect 12459 1793 12471 4731
rect 12483 1793 12495 6291
rect 12507 2081 12519 7371
rect 12555 6017 12567 7515
rect 12531 1793 12543 5115
rect 12579 3929 12591 7515
rect 12555 1793 12567 1923
rect 12579 1793 12591 2403
rect 12603 1937 12615 6795
rect 12627 3161 12639 7515
rect 12675 6809 12687 7515
rect 12699 7313 12711 7515
rect 12747 7313 12759 7515
rect 12651 1793 12663 4035
rect 12675 1793 12687 4491
rect 12699 1793 12711 2403
rect 12747 1793 12759 6555
rect 12795 6209 12807 7515
rect 12819 4913 12831 7515
rect 12843 6569 12855 7515
rect 12891 7385 12903 7515
rect 12771 1793 12783 3243
rect 12795 1793 12807 1923
rect 12843 1793 12855 1899
rect 12867 1793 12879 5523
rect 12915 4361 12927 7515
rect 12939 7409 12951 7515
rect 12891 1793 12903 1875
rect 12939 1793 12951 2955
rect 12963 1793 12975 7419
rect 12987 4841 12999 7515
rect 13011 3449 13023 7515
rect 13035 1961 13047 7515
rect 13083 7457 13095 7515
rect 12987 1793 12999 1851
rect 13059 1793 13071 5811
rect 13083 1793 13095 5211
rect 13107 4841 13119 7515
rect 13131 4673 13143 7515
rect 13107 1793 13119 1947
rect 13155 1793 13167 6531
rect 13179 4361 13191 7515
rect 13203 3521 13215 7515
rect 13227 5561 13239 7515
rect 13179 1793 13191 1827
rect 13203 1793 13215 1803
rect 13251 1793 13263 6075
rect 13275 4673 13287 7515
rect 13299 4433 13311 7515
rect 13347 6449 13359 7515
rect 13275 1793 13287 4395
rect 13323 1865 13335 6387
rect 13395 5561 13407 7515
rect 13419 4793 13431 7515
rect 13347 1793 13359 3315
rect 13371 1793 13383 3219
rect 13467 2681 13479 7515
rect 13395 1793 13407 1851
rect 13443 1793 13455 1971
rect 13491 1793 13503 7323
rect 13515 5705 13527 7515
rect 13539 6401 13551 7515
rect 13563 6065 13575 7515
rect 13587 4121 13599 7515
rect 13611 6449 13623 7515
rect 13659 7481 13671 7515
rect 13539 1793 13551 3819
rect 13563 1793 13575 2667
rect 13635 1793 13647 7155
rect 13659 1793 13671 4011
rect 13683 2057 13695 7515
rect 13707 6281 13719 7515
rect 13731 7505 13743 7515
rect 13731 1793 13743 7035
rect 13755 1841 13767 5091
rect 13779 5009 13791 7515
rect 13803 6281 13815 7515
rect 13779 1793 13791 2043
rect 13815 1817 13827 5907
rect 13851 2249 13863 7515
rect 13899 6305 13911 7515
rect 13923 6449 13935 7515
rect 13875 1793 13887 4491
rect 13899 1793 13911 3747
rect 13947 1793 13959 3915
rect 13971 1793 13983 3411
rect 13995 2921 14007 7515
rect 13995 1793 14007 2379
rect 14019 2225 14031 7515
rect 14043 4577 14055 7515
rect 14067 7097 14079 7515
rect 14043 1793 14055 3747
rect 14067 1793 14079 2379
rect 14091 1793 14103 3915
rect 14115 3209 14127 7515
rect 14139 2897 14151 7515
rect 14163 5009 14175 7515
rect 14163 1793 14175 4395
rect 14187 1793 14199 5691
rect 14211 3713 14223 4659
rect 14235 2825 14247 6387
rect 14283 6137 14295 7515
rect 14259 1793 14271 4659
rect 14283 1793 14295 4491
rect 14307 2681 14319 6075
rect 14343 3761 14355 5523
rect 14331 1793 14343 3387
rect 14379 1793 14391 2379
rect 14403 1793 14415 5523
rect 14427 1793 14439 5115
rect 14451 3089 14463 7467
rect 14643 7433 14655 7515
rect 14475 2057 14487 6819
rect 14499 1793 14511 5499
rect 14523 1793 14535 3747
rect 14547 2393 14559 7323
rect 14835 7097 14847 7515
rect 14571 1793 14583 6531
rect 14595 1793 14607 2451
rect 14619 1793 14631 6963
rect 14667 1793 14679 4587
rect 14691 1793 14703 3195
rect 14739 1793 14751 4587
rect 14787 1793 14799 5691
rect 14811 1793 14823 3219
rect 14835 1793 14847 7011
rect 14859 6833 14871 7515
rect 14883 5921 14895 7515
rect 14943 6185 14955 7083
rect 15003 5921 15015 7515
rect 14883 1793 14895 4491
rect 14907 1793 14919 3411
rect 14943 3305 14955 5907
rect 14931 1793 14943 2523
rect 15027 1793 15039 7131
rect 15099 1793 15111 3075
rect 15123 1793 15135 6003
rect 15363 5561 15375 7515
rect 15411 6017 15423 7515
rect 15147 1793 15159 2667
rect 15195 1793 15207 2523
rect 15243 1793 15255 2451
rect 15291 1793 15303 2283
rect 15315 1793 15327 3507
rect 15387 1793 15399 4179
rect 15411 1793 15423 3675
rect 15435 1793 15447 5403
rect 15483 1793 15495 2883
rect 15507 1793 15519 4779
rect 15555 4169 15567 7515
rect 15579 4193 15591 7515
rect 15627 6425 15639 7515
rect 15675 6065 15687 7515
rect 15531 1793 15543 3363
rect 15555 1793 15567 2379
rect 15603 1793 15615 3915
rect 15627 1793 15639 3243
rect 15651 1793 15663 4155
rect 15699 3161 15711 7515
rect 15699 1793 15711 2811
rect 15723 1793 15735 4491
rect 15747 4145 15759 7515
rect 15795 6665 15807 7515
rect 15819 3233 15831 7515
rect 15843 5417 15855 7515
rect 15891 3425 15903 7515
rect 15939 3257 15951 7515
rect 16011 6473 16023 7515
rect 16035 5681 16047 7515
rect 16083 5681 16095 7515
rect 16131 6137 16143 7515
rect 16155 6305 16167 7515
rect 16179 6401 16191 7515
rect 15771 1793 15783 2499
rect 16227 2465 16239 7515
rect 16275 6185 16287 7515
rect 16299 5825 16311 7515
rect 16323 6953 16335 7515
rect 16299 1793 16311 2091
rect 16371 1961 16383 7515
rect 16395 1889 16407 7515
rect 16419 6425 16431 7515
rect 16443 2393 16455 7515
rect 16467 6809 16479 7515
rect 16515 5633 16527 7515
rect 16539 7169 16551 7515
rect 16443 1793 16455 1995
rect 16467 1793 16479 5619
rect 16587 2921 16599 7515
rect 16515 1793 16527 2451
rect 16563 1793 16575 2379
rect 16611 1793 16623 7371
rect 16635 2753 16647 7515
rect 16659 6449 16671 7515
rect 16683 6473 16695 7515
rect 16707 4889 16719 7515
rect 16659 1793 16671 2787
rect 16683 1793 16695 4491
rect 16707 1793 16719 2883
rect 16731 2369 16743 6435
rect 16755 3737 16767 7515
rect 16779 3233 16791 7515
rect 16803 3881 16815 7515
rect 16851 7457 16863 7515
rect 16827 2849 16839 6339
rect 16875 2897 16887 7515
rect 16899 4889 16911 7515
rect 16755 1793 16767 2835
rect 16779 1793 16791 2739
rect 16803 1793 16815 2835
rect 16899 1793 16911 3867
rect 16923 1793 16935 4347
rect 16947 2465 16959 7515
rect 16995 6353 17007 7515
rect 16995 1793 17007 4227
rect 17019 1793 17031 3411
rect 17043 2033 17055 7515
rect 17067 2561 17079 6339
rect 17115 4145 17127 7515
rect 17139 5225 17151 7515
rect 17187 4625 17199 7515
rect 17307 7505 17319 7515
rect 17091 1793 17103 4011
rect 17211 1793 17223 5499
rect 17259 1793 17271 4227
rect 17331 1793 17343 3507
rect 17355 1793 17367 3411
rect 17379 1793 17391 6219
rect 17427 1793 17439 3387
rect 17475 1793 17487 5955
rect 17523 1793 17535 6003
rect 17571 1793 17583 2835
rect 17619 1793 17631 2547
rect 17691 1793 17703 5163
rect 17715 2081 17727 7515
rect 17739 1793 17751 5523
rect 17763 1793 17775 5547
rect 17859 4169 17871 7515
rect 17883 4433 17895 7515
rect 17907 5969 17919 7515
rect 17955 6065 17967 7515
rect 17787 1793 17799 2451
rect 17835 1793 17847 2931
rect 17859 1793 17871 3699
rect 17907 1793 17919 5043
rect 17931 1913 17943 5955
rect 17979 4361 17991 7515
rect 18003 2441 18015 7515
rect 18051 4217 18063 7515
rect 18075 4121 18087 7515
rect 18123 5321 18135 7515
rect 18171 6545 18183 7515
rect 18195 4049 18207 7515
rect 18219 6641 18231 7515
rect 18267 3401 18279 7515
rect 18291 5321 18303 7515
rect 18315 4313 18327 7515
rect 18363 2513 18375 7515
rect 18387 4985 18399 7515
rect 18411 3641 18423 7515
rect 18459 5609 18471 7515
rect 18483 2201 18495 7515
rect 18507 5801 18519 7515
rect 18579 5153 18591 7515
rect 18627 6353 18639 7515
rect 18699 6209 18711 7515
rect 18627 1793 18639 6171
rect 18723 5465 18735 7515
rect 18771 6617 18783 7515
rect 18699 1793 18711 4299
rect 18747 1793 18759 4155
rect 18819 3929 18831 7515
rect 18843 6089 18855 7515
rect 18819 1793 18831 3555
rect 18843 1793 18855 3387
rect 18867 3089 18879 7515
rect 18891 3401 18903 6507
rect 18915 5609 18927 7515
rect 18915 1793 18927 5475
rect 18939 3305 18951 7515
rect 18963 3761 18975 5595
rect 18987 2369 18999 7035
rect 19011 5153 19023 7515
rect 19035 5465 19047 7515
rect 19083 6137 19095 7515
rect 19131 5465 19143 7515
rect 19179 6785 19191 7515
rect 18939 1793 18951 2355
rect 19011 1793 19023 3747
rect 19035 1793 19047 3243
rect 19059 2321 19071 5451
rect 19083 1793 19095 3579
rect 19131 1793 19143 4683
rect 19155 1793 19167 5739
rect 19203 3857 19215 7515
rect 19227 5993 19239 7515
rect 19203 1793 19215 3579
rect 19251 1793 19263 4131
rect 19275 3881 19287 7515
rect 19275 1793 19287 3363
rect 19299 2441 19311 7515
rect 19323 4169 19335 5451
rect 19347 4673 19359 7515
rect 19347 1793 19359 3747
rect 19371 1793 19383 3651
rect 19395 2705 19407 7515
rect 19419 4385 19431 7515
rect 19443 2465 19455 7515
rect 19467 3977 19479 7515
rect 19467 1793 19479 3651
rect 19491 1793 19503 4395
rect 19515 3353 19527 7515
rect 19539 4505 19551 7515
rect 19563 4841 19575 7515
rect 19539 1793 19551 4371
rect 19587 1793 19599 5883
rect 19611 4457 19623 7515
rect 19635 4673 19647 7515
rect 19659 3833 19671 7515
rect 19683 3665 19695 5547
rect 19707 4985 19719 7515
rect 19707 1793 19719 4611
rect 19731 2825 19743 7515
rect 19755 4121 19767 7515
rect 19731 1793 19743 2691
rect 19755 1793 19767 3963
rect 19779 3881 19791 7515
rect 19827 4865 19839 7515
rect 19851 5465 19863 7515
rect 19803 1793 19815 4515
rect 19851 1793 19863 4923
rect 19875 4337 19887 7515
rect 19899 4385 19911 7443
rect 19923 5705 19935 7515
rect 19947 4433 19959 7515
rect 19971 7265 19983 7515
rect 19923 1793 19935 2715
rect 19983 2705 19995 4995
rect 20019 2681 20031 7515
rect 20043 4841 20055 7515
rect 20067 6449 20079 7515
rect 20043 1793 20055 3771
rect 20067 1793 20079 6315
rect 20091 6041 20103 7515
rect 20115 6641 20127 7515
rect 20163 7337 20175 7515
rect 20115 1793 20127 6555
rect 20139 1793 20151 5403
rect 20163 1793 20175 7227
rect 20187 3089 20199 7515
rect 20211 3977 20223 5931
rect 20235 4865 20247 7515
rect 20187 1793 20199 2691
rect 20235 1793 20247 2787
rect 20259 1793 20271 3219
rect 20283 2705 20295 7515
rect 20307 5921 20319 6627
rect 20307 2489 20319 5451
rect 20331 5009 20343 7515
rect 20355 6137 20367 7515
rect 20379 7289 20391 7515
rect 20331 1793 20343 4059
rect 20355 1793 20367 6051
rect 20379 1793 20391 2019
rect 20403 1793 20415 5259
rect 20427 2417 20439 7515
rect 20451 5897 20463 7515
rect 20475 5873 20487 7515
rect 20523 6329 20535 7515
rect 20451 1793 20463 5811
rect 20475 1793 20487 2715
rect 20499 1793 20511 4347
rect 20523 1793 20535 6147
rect 20547 4793 20559 7515
rect 20571 2345 20583 7515
rect 20595 1793 20607 4707
rect 20619 3641 20631 7515
rect 20643 6881 20655 7515
rect 20667 5777 20679 7515
rect 20691 1793 20703 6147
rect 20715 2609 20727 7515
rect 20739 6017 20751 7515
rect 20763 5273 20775 7515
rect 20787 5609 20799 7515
rect 20823 5561 20835 6123
rect 20715 1793 20727 2475
rect 20763 1793 20775 4419
rect 20787 1793 20799 5547
rect 20811 1793 20823 4467
rect 20835 3137 20847 4827
rect 20859 3593 20871 7323
rect 20907 5729 20919 7515
rect 20883 1793 20895 3699
rect 20907 1793 20919 2715
rect 20931 1793 20943 3435
rect 20955 1793 20967 5331
rect 20979 2129 20991 4851
rect 21003 1937 21015 5883
rect 21027 2945 21039 6315
rect 21051 1793 21063 4611
rect 21075 2489 21087 4299
rect 21099 3497 21111 5259
rect 21123 1793 21135 4083
rect 21171 1793 21183 7155
rect 21267 6329 21279 7515
rect 21195 1793 21207 3051
rect 21243 1793 21255 5571
rect 21267 1793 21279 6219
rect 21291 1793 21303 5091
rect 21315 3185 21327 7515
rect 21339 1793 21351 6507
rect 21459 5585 21471 7515
rect 21387 1793 21399 4035
rect 21459 1793 21471 5547
rect 21507 5393 21519 7515
rect 21531 4505 21543 7515
rect 21555 6425 21567 7515
rect 21603 5561 21615 7515
rect 21483 1793 21495 4083
rect 21507 1793 21519 4011
rect 21531 1793 21543 4443
rect 21579 1793 21591 2715
rect 21603 1793 21615 3915
rect 21627 2945 21639 7515
rect 21675 6137 21687 7515
rect 21723 6953 21735 7515
rect 21651 4313 21663 5571
rect 21675 1793 21687 6099
rect 21699 1793 21711 3171
rect 21723 1793 21735 6891
rect 21747 4457 21759 7059
rect 21771 4481 21783 7515
rect 21795 6209 21807 7515
rect 21819 4985 21831 7515
rect 21795 1793 21807 3411
rect 21843 2561 21855 7515
rect 21867 1793 21879 4131
rect 21891 4121 21903 7515
rect 21939 7169 21951 7515
rect 21891 1793 21903 4083
rect 21915 1793 21927 4251
rect 21963 1793 21975 6987
rect 22011 4505 22023 7515
rect 21987 1793 21999 3459
rect 22011 1793 22023 4443
rect 22035 2729 22047 6123
rect 22059 5705 22071 7515
rect 22131 7121 22143 7515
rect 22059 1793 22071 4515
rect 22083 1793 22095 4491
rect 22107 1793 22119 3747
rect 22155 1793 22167 4131
rect 22179 2537 22191 7515
rect 22215 4625 22227 6939
rect 22251 5273 22263 7515
rect 22275 6209 22287 7515
rect 22203 1793 22215 3267
rect 22251 1793 22263 5187
rect 22299 4937 22311 7515
rect 22323 5441 22335 7515
rect 22275 1793 22287 3411
rect 22347 1793 22359 3723
rect 22371 2513 22383 7515
rect 22395 7361 22407 7515
rect 22419 6281 22431 7515
rect 22467 3809 22479 7515
rect 22515 7193 22527 7515
rect 22491 4097 22503 5739
rect 22371 1793 22383 2475
rect 22443 1793 22455 3747
rect 22467 1793 22479 3507
rect 22515 1793 22527 4539
rect 22539 4529 22551 6531
rect 22587 4721 22599 7515
rect 22563 1793 22575 4611
rect 22587 1793 22599 4707
rect 22611 3713 22623 7515
rect 22635 6305 22647 7515
rect 22683 5345 22695 7515
rect 22731 6593 22743 7515
rect 22611 1793 22623 3651
rect 22659 1793 22671 4563
rect 22683 1793 22695 5211
rect 22707 1793 22719 4395
rect 22755 3473 22767 7515
rect 22755 1793 22767 3387
rect 22779 1793 22791 5691
rect 22803 2201 22815 7515
rect 22851 6833 22863 7515
rect 22827 2921 22839 5259
rect 22851 1793 22863 6051
rect 22875 4721 22887 7515
rect 22899 6689 22911 7515
rect 22875 1793 22887 4563
rect 22923 1793 22935 7251
rect 22947 3713 22959 7515
rect 22971 6089 22983 7515
rect 22995 7049 23007 7515
rect 22947 1793 22959 3627
rect 22995 1793 23007 5307
rect 23019 2489 23031 6339
rect 23043 4745 23055 7515
rect 23067 4937 23079 7515
rect 23091 5657 23103 7515
rect 23103 4457 23115 5331
rect 23043 1793 23055 2619
rect 23067 1793 23079 4275
rect 23139 4241 23151 7515
rect 23091 1793 23103 3891
rect 23163 2921 23175 7515
rect 23163 1793 23175 2787
rect 23187 1793 23199 3459
rect 23211 3209 23223 7515
rect 23235 3665 23247 5835
rect 23259 4793 23271 7515
rect 23283 4745 23295 7515
rect 23307 5369 23319 7515
rect 23355 6305 23367 7515
rect 23211 1793 23223 3171
rect 23259 1793 23271 3027
rect 23283 1793 23295 4467
rect 23319 3233 23331 4731
rect 23379 3161 23391 7515
rect 23403 5681 23415 7515
rect 23427 2345 23439 7515
rect 23451 5297 23463 7515
rect 23475 3401 23487 6195
rect 23499 5537 23511 7515
rect 23523 4721 23535 7515
rect 23571 7361 23583 7515
rect 23547 4577 23559 6915
rect 23583 3641 23595 6099
rect 23619 2777 23631 7515
rect 23643 2801 23655 6987
rect 23667 4745 23679 7515
rect 23739 6617 23751 7515
rect 23763 4937 23775 7515
rect 23787 3017 23799 7515
rect 23835 6857 23847 7515
rect 23859 6497 23871 7515
rect 23883 5033 23895 7515
rect 23787 1793 23799 2931
rect 23835 1793 23847 4707
rect 23931 2153 23943 7515
rect 23955 4889 23967 7515
rect 23979 2105 23991 7515
rect 24003 4625 24015 7515
rect 23979 1793 23991 2067
rect 24027 1793 24039 7299
rect 24051 7169 24063 7515
rect 24051 1793 24063 3603
rect 24075 3521 24087 7515
rect 24099 3497 24111 5139
rect 24075 1793 24087 3483
rect 24099 2081 24111 2667
rect 24123 2585 24135 7515
rect 24147 2561 24159 7035
rect 24171 5561 24183 7515
rect 24123 1793 24135 2547
rect 24171 1793 24183 4995
rect 24195 4961 24207 7515
rect 24219 5873 24231 7515
rect 24219 1793 24231 5835
rect 24267 5177 24279 7515
rect 24243 1793 24255 3843
rect 24267 1793 24279 4611
rect 24291 2201 24303 7515
rect 24315 7409 24327 7515
rect 24327 4673 24339 5859
rect 24351 4625 24363 6435
rect 24387 3761 24399 7515
rect 24411 1865 24423 7515
rect 24459 5513 24471 7515
rect 24507 6185 24519 7515
rect 24531 3449 24543 7515
rect 24555 2273 24567 7515
rect 24603 4193 24615 7515
rect 24627 3689 24639 7515
rect 24723 5633 24735 7515
rect 24795 6137 24807 7515
rect 24747 1793 24759 3435
rect 24795 1793 24807 6075
rect 24819 4601 24831 7515
rect 24843 5177 24855 7515
rect 24867 2201 24879 6123
rect 24915 2897 24927 7515
rect 24939 5201 24951 7515
rect 24963 6785 24975 7515
rect 24939 1793 24951 2235
rect 24963 1793 24975 6699
rect 24987 4673 24999 7515
rect 25011 4769 25023 7515
rect 24987 1793 24999 3459
rect 25011 1793 25023 4611
rect 25035 2849 25047 6771
rect 25059 4721 25071 7515
rect 25083 4769 25095 7515
rect 25107 6785 25119 7515
rect 25059 1793 25071 3555
rect 25083 1793 25095 4347
rect 25107 1793 25119 6747
rect 25131 3425 25143 4659
rect 25155 1793 25167 3147
rect 25179 2993 25191 7515
rect 25203 6377 25215 7515
rect 25179 1793 25191 2931
rect 25203 1793 25215 4659
rect 25227 2729 25239 4707
rect 25251 4145 25263 7515
rect 25275 4913 25287 7515
rect 25299 5513 25311 7515
rect 25347 6209 25359 7515
rect 25251 1793 25263 3435
rect 25275 1793 25287 4779
rect 25299 1793 25311 5475
rect 25323 2657 25335 4755
rect 25347 1793 25359 6171
rect 25371 5081 25383 7515
rect 25395 6785 25407 7515
rect 25371 1793 25383 4587
rect 25419 4001 25431 7515
rect 25443 4673 25455 6723
rect 25467 4625 25479 7515
rect 25515 5705 25527 7515
rect 25491 4649 25503 5499
rect 25539 2825 25551 7515
rect 25563 5057 25575 7515
rect 25587 7169 25599 7515
rect 25611 5273 25623 7515
rect 25611 1793 25623 5235
rect 25635 5129 25647 6195
rect 25659 3713 25671 7515
rect 25683 3449 25695 7515
rect 25707 6473 25719 7515
rect 25683 1793 25695 3411
rect 25707 1793 25719 3531
rect 25731 1793 25743 4731
rect 25755 4217 25767 7515
rect 25779 6329 25791 7515
rect 25755 1793 25767 3459
rect 25779 1793 25791 4659
rect 25803 4121 25815 7515
rect 25827 2753 25839 7515
rect 25875 7361 25887 7515
rect 25851 4601 25863 6075
rect 25899 4073 25911 7515
rect 25923 2873 25935 7515
rect 25971 6017 25983 7515
rect 25947 2393 25959 5259
rect 25995 5225 26007 7515
rect 26019 4697 26031 7515
rect 26043 3425 26055 5787
rect 26067 5609 26079 7515
rect 26091 3929 26103 7515
rect 26115 3113 26127 7515
rect 26163 6113 26175 7515
rect 26187 2969 26199 7515
rect 26211 6257 26223 7515
rect 26259 3329 26271 7515
rect 26283 7457 26295 7515
rect 26307 4505 26319 7515
rect 26331 7217 26343 7515
rect 26379 4673 26391 7515
rect 26427 3185 26439 7515
rect 26427 1865 26439 2163
rect 26451 1817 26463 3939
rect 26475 1841 26487 6387
rect 26570 1793 26770 7515
rect 26883 4804 26953 4816
rect 26883 1852 26953 1864
rect 26883 1828 26953 1840
rect 26883 1804 26953 1816
rect 0 131 70 143
rect 0 107 70 119
rect 123 0 323 994
rect 339 0 351 994
rect 363 0 375 994
rect 387 0 399 994
rect 411 0 423 994
rect 2331 168 2343 994
rect 2379 192 2391 994
rect 2427 120 2439 994
rect 2475 120 2487 994
rect 2571 216 2583 994
rect 2643 240 2655 994
rect 3723 264 3735 994
rect 3843 288 3855 994
rect 3987 192 3999 994
rect 4131 192 4143 994
rect 4347 168 4359 994
rect 4419 168 4431 994
rect 4635 168 4647 994
rect 5115 312 5127 994
rect 5283 336 5295 994
rect 6027 264 6039 994
rect 6075 360 6087 994
rect 6171 384 6183 994
rect 4432 154 4450 168
rect 4431 0 4443 154
rect 6267 96 6279 994
rect 6651 408 6663 994
rect 6699 432 6711 994
rect 6723 408 6735 994
rect 6771 336 6783 994
rect 6819 336 6831 994
rect 7035 408 7047 994
rect 7179 456 7191 994
rect 7491 72 7503 994
rect 7539 480 7551 994
rect 7563 504 7575 994
rect 7611 528 7623 994
rect 7827 552 7839 994
rect 8115 96 8127 994
rect 8163 576 8175 994
rect 8211 504 8223 994
rect 8427 384 8439 994
rect 8571 504 8583 994
rect 8643 600 8655 994
rect 8715 624 8727 994
rect 8739 648 8751 994
rect 8955 672 8967 994
rect 9003 696 9015 994
rect 9051 720 9063 994
rect 9483 744 9495 994
rect 9555 96 9567 994
rect 10347 96 10359 994
rect 10371 768 10383 994
rect 10395 792 10407 994
rect 10443 816 10455 994
rect 7815 0 7827 82
rect 10587 48 10599 994
rect 10779 840 10791 994
rect 10947 864 10959 994
rect 11043 888 11055 994
rect 11307 24 11319 994
rect 11403 384 11415 994
rect 11667 192 11679 994
rect 12387 480 12399 994
rect 12603 144 12615 994
rect 13035 480 13047 994
rect 13299 384 13311 994
rect 13467 336 13479 994
rect 13587 192 13599 994
rect 13683 144 13695 994
rect 13851 912 13863 994
rect 14115 840 14127 994
rect 14211 96 14223 994
rect 14475 840 14487 994
rect 14979 288 14991 994
rect 15003 96 15015 994
rect 15051 288 15063 994
rect 15219 816 15231 994
rect 15339 936 15351 994
rect 15891 960 15903 994
rect 16587 984 16599 994
rect 16827 312 16839 994
rect 16851 840 16863 994
rect 16947 840 16959 994
rect 17043 96 17055 994
rect 17139 600 17151 994
rect 17451 600 17463 994
rect 17547 936 17559 994
rect 17643 720 17655 994
rect 17464 586 17482 600
rect 17463 0 17475 586
rect 18027 120 18039 994
rect 18435 960 18447 994
rect 18579 456 18591 994
rect 18867 984 18879 994
rect 18963 600 18975 994
rect 19299 816 19311 994
rect 19419 432 19431 994
rect 19635 576 19647 994
rect 19947 600 19959 994
rect 19971 648 19983 994
rect 20019 552 20031 994
rect 20283 768 20295 994
rect 20571 240 20583 994
rect 20619 672 20631 994
rect 20667 744 20679 994
rect 20835 336 20847 994
rect 21003 504 21015 994
rect 21147 264 21159 994
rect 21627 456 21639 994
rect 21771 144 21783 994
rect 21819 408 21831 994
rect 22179 792 22191 994
rect 22299 480 22311 994
rect 22395 216 22407 994
rect 22803 720 22815 994
rect 22899 840 22911 994
rect 22995 504 23007 994
rect 23008 490 23026 504
rect 23007 0 23019 490
rect 23139 360 23151 994
rect 23307 912 23319 994
rect 23427 696 23439 994
rect 24003 192 24015 994
rect 24147 384 24159 994
rect 24387 528 24399 994
rect 25395 624 25407 994
rect 25443 288 25455 994
rect 25491 888 25503 994
rect 25563 864 25575 994
rect 25563 72 25575 82
rect 25587 48 25599 58
rect 25611 48 25623 154
rect 26570 0 26770 994
rect 26883 83 26953 95
rect 26883 59 26953 71
rect 26883 35 26953 47
rect 26883 11 26953 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7515
box 0 0 1464 799
use nand4 g8369
timestamp 1386234936
transform 1 0 1587 0 1 7515
box 0 0 144 799
use nor2 g8169
timestamp 1386235306
transform 1 0 1731 0 1 7515
box 0 0 120 799
use nand2 g8107
timestamp 1386234792
transform 1 0 1851 0 1 7515
box 0 0 96 799
use nand2 g8229
timestamp 1386234792
transform 1 0 1947 0 1 7515
box 0 0 96 799
use nand2 g8370
timestamp 1386234792
transform 1 0 2043 0 1 7515
box 0 0 96 799
use inv g8344
timestamp 1386238110
transform 1 0 2139 0 1 7515
box 0 0 120 799
use nand2 g8123
timestamp 1386234792
transform 1 0 2259 0 1 7515
box 0 0 96 799
use nand2 g8222
timestamp 1386234792
transform 1 0 2355 0 1 7515
box 0 0 96 799
use nand2 g8102
timestamp 1386234792
transform 1 0 2451 0 1 7515
box 0 0 96 799
use nand2 g8098
timestamp 1386234792
transform 1 0 2547 0 1 7515
box 0 0 96 799
use nand2 g8314
timestamp 1386234792
transform 1 0 2643 0 1 7515
box 0 0 96 799
use inv g8327
timestamp 1386238110
transform 1 0 2739 0 1 7515
box 0 0 120 799
use nand2 g8187
timestamp 1386234792
transform 1 0 2859 0 1 7515
box 0 0 96 799
use nand4 g8171
timestamp 1386234936
transform 1 0 2955 0 1 7515
box 0 0 144 799
use nand2 g8135
timestamp 1386234792
transform 1 0 3099 0 1 7515
box 0 0 96 799
use nand2 g8295
timestamp 1386234792
transform 1 0 3195 0 1 7515
box 0 0 96 799
use nor2 g8287
timestamp 1386235306
transform 1 0 3291 0 1 7515
box 0 0 120 799
use nor2 g8261
timestamp 1386235306
transform 1 0 3411 0 1 7515
box 0 0 120 799
use nand2 g8276
timestamp 1386234792
transform 1 0 3531 0 1 7515
box 0 0 96 799
use nand3 g8130
timestamp 1396952988
transform 1 0 3627 0 1 7515
box 0 0 120 799
use nor2 g8082
timestamp 1386235306
transform 1 0 3747 0 1 7515
box 0 0 120 799
use nand4 g8318
timestamp 1386234936
transform 1 0 3867 0 1 7515
box 0 0 144 799
use nor2 g8377
timestamp 1386235306
transform 1 0 4011 0 1 7515
box 0 0 120 799
use inv g8390
timestamp 1386238110
transform 1 0 4131 0 1 7515
box 0 0 120 799
use nand2 g8168
timestamp 1386234792
transform 1 0 4251 0 1 7515
box 0 0 96 799
use nand2 g8238
timestamp 1386234792
transform 1 0 4347 0 1 7515
box 0 0 96 799
use nand2 g8225
timestamp 1386234792
transform 1 0 4443 0 1 7515
box 0 0 96 799
use nand4 g8143
timestamp 1386234936
transform 1 0 4539 0 1 7515
box 0 0 144 799
use nand2 g8333
timestamp 1386234792
transform 1 0 4683 0 1 7515
box 0 0 96 799
use and2 g2
timestamp 1386234845
transform 1 0 4779 0 1 7515
box 0 0 120 799
use nor2 g8149
timestamp 1386235306
transform 1 0 4899 0 1 7515
box 0 0 120 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 5019 0 1 7515
box 0 0 48 799
use nand3 g8069
timestamp 1396952988
transform 1 0 5067 0 1 7515
box 0 0 120 799
use nand4 g8338
timestamp 1386234936
transform 1 0 5187 0 1 7515
box 0 0 144 799
use nand3 g8280
timestamp 1396952988
transform 1 0 5331 0 1 7515
box 0 0 120 799
use and2 g8249
timestamp 1386234845
transform 1 0 5451 0 1 7515
box 0 0 120 799
use nand2 g8064
timestamp 1386234792
transform 1 0 5571 0 1 7515
box 0 0 96 799
use nand2 g8310
timestamp 1386234792
transform 1 0 5667 0 1 7515
box 0 0 96 799
use inv g8235
timestamp 1386238110
transform 1 0 5763 0 1 7515
box 0 0 120 799
use nand2 g8362
timestamp 1386234792
transform 1 0 5883 0 1 7515
box 0 0 96 799
use mux2 g8055
timestamp 1386235218
transform 1 0 5979 0 1 7515
box 0 0 192 799
use nand3 g8088
timestamp 1396952988
transform 1 0 6171 0 1 7515
box 0 0 120 799
use nand3 g8214
timestamp 1396952988
transform 1 0 6291 0 1 7515
box 0 0 120 799
use nand2 g8056
timestamp 1386234792
transform 1 0 6411 0 1 7515
box 0 0 96 799
use nand3 g8281
timestamp 1396952988
transform 1 0 6507 0 1 7515
box 0 0 120 799
use nand3 g8366
timestamp 1396952988
transform 1 0 6627 0 1 7515
box 0 0 120 799
use nor2 g8269
timestamp 1386235306
transform 1 0 6747 0 1 7515
box 0 0 120 799
use nor2 g8183
timestamp 1386235306
transform 1 0 6867 0 1 7515
box 0 0 120 799
use nand3 g8170
timestamp 1396952988
transform 1 0 6987 0 1 7515
box 0 0 120 799
use nand2 g8124
timestamp 1386234792
transform 1 0 7107 0 1 7515
box 0 0 96 799
use nand2 g8106
timestamp 1386234792
transform 1 0 7203 0 1 7515
box 0 0 96 799
use nand2 g8414
timestamp 1386234792
transform 1 0 7299 0 1 7515
box 0 0 96 799
use inv g8119
timestamp 1386238110
transform 1 0 7395 0 1 7515
box 0 0 120 799
use inv g8275
timestamp 1386238110
transform 1 0 7515 0 1 7515
box 0 0 120 799
use nand2 g8146
timestamp 1386234792
transform 1 0 7635 0 1 7515
box 0 0 96 799
use nand2 g8127
timestamp 1386234792
transform 1 0 7731 0 1 7515
box 0 0 96 799
use nand2 g8155
timestamp 1386234792
transform 1 0 7827 0 1 7515
box 0 0 96 799
use inv g8290
timestamp 1386238110
transform 1 0 7923 0 1 7515
box 0 0 120 799
use nand3 g8252
timestamp 1396952988
transform 1 0 8043 0 1 7515
box 0 0 120 799
use nand2 g8334
timestamp 1386234792
transform 1 0 8163 0 1 7515
box 0 0 96 799
use nand2 g8244
timestamp 1386234792
transform 1 0 8259 0 1 7515
box 0 0 96 799
use nand2 g8240
timestamp 1386234792
transform 1 0 8355 0 1 7515
box 0 0 96 799
use inv g8054
timestamp 1386238110
transform 1 0 8451 0 1 7515
box 0 0 120 799
use nand3 g8407
timestamp 1396952988
transform 1 0 8571 0 1 7515
box 0 0 120 799
use and2 g8139
timestamp 1386234845
transform 1 0 8691 0 1 7515
box 0 0 120 799
use and2 g8118
timestamp 1386234845
transform 1 0 8811 0 1 7515
box 0 0 120 799
use nand4 g8363
timestamp 1386234936
transform 1 0 8931 0 1 7515
box 0 0 144 799
use nand2 g8111
timestamp 1386234792
transform 1 0 9075 0 1 7515
box 0 0 96 799
use nand2 g8381
timestamp 1386234792
transform 1 0 9171 0 1 7515
box 0 0 96 799
use nand2 g8403
timestamp 1386234792
transform 1 0 9267 0 1 7515
box 0 0 96 799
use inv g8357
timestamp 1386238110
transform 1 0 9363 0 1 7515
box 0 0 120 799
use rowcrosser PcWe
timestamp 1386086759
transform 1 0 9483 0 1 7515
box 0 0 48 799
use nand2 g8347
timestamp 1386234792
transform 1 0 9531 0 1 7515
box 0 0 96 799
use nand2 g8120
timestamp 1386234792
transform 1 0 9627 0 1 7515
box 0 0 96 799
use nand4 g8091
timestamp 1386234936
transform 1 0 9723 0 1 7515
box 0 0 144 799
use nand4 g8134
timestamp 1386234936
transform 1 0 9867 0 1 7515
box 0 0 144 799
use and2 g8386
timestamp 1386234845
transform 1 0 10011 0 1 7515
box 0 0 120 799
use nand2 g8425
timestamp 1386234792
transform 1 0 10131 0 1 7515
box 0 0 96 799
use inv g8320
timestamp 1386238110
transform 1 0 10227 0 1 7515
box 0 0 120 799
use rowcrosser AluOR_91_0_93_
timestamp 1386086759
transform 1 0 10347 0 1 7515
box 0 0 48 799
use rowcrosser ALE
timestamp 1386086759
transform 1 0 10395 0 1 7515
box 0 0 48 799
use and2 g8354
timestamp 1386234845
transform 1 0 10443 0 1 7515
box 0 0 120 799
use nand2 g8374
timestamp 1386234792
transform 1 0 10563 0 1 7515
box 0 0 96 799
use nand2 g8050
timestamp 1386234792
transform 1 0 10659 0 1 7515
box 0 0 96 799
use nand4 g8218
timestamp 1386234936
transform 1 0 10755 0 1 7515
box 0 0 144 799
use rowcrosser StatusRegEn
timestamp 1386086759
transform 1 0 10899 0 1 7515
box 0 0 48 799
use nand2 g8284
timestamp 1386234792
transform 1 0 10947 0 1 7515
box 0 0 96 799
use nand3 g8198
timestamp 1396952988
transform 1 0 11043 0 1 7515
box 0 0 120 799
use rowcrosser PcSel_91_2_93_
timestamp 1386086759
transform 1 0 11163 0 1 7515
box 0 0 48 799
use nand2 g8272
timestamp 1386234792
transform 1 0 11211 0 1 7515
box 0 0 96 799
use nor2 g8199
timestamp 1386235306
transform 1 0 11307 0 1 7515
box 0 0 120 799
use nand2 g8306
timestamp 1386234792
transform 1 0 11427 0 1 7515
box 0 0 96 799
use nand3 g8221
timestamp 1396952988
transform 1 0 11523 0 1 7515
box 0 0 120 799
use nand3 g8319
timestamp 1396952988
transform 1 0 11643 0 1 7515
box 0 0 120 799
use nand2 g8392
timestamp 1386234792
transform 1 0 11763 0 1 7515
box 0 0 96 799
use nand2 g8194
timestamp 1386234792
transform 1 0 11859 0 1 7515
box 0 0 96 799
use nand2 g8230
timestamp 1386234792
transform 1 0 11955 0 1 7515
box 0 0 96 799
use nor2 g8271
timestamp 1386235306
transform 1 0 12051 0 1 7515
box 0 0 120 799
use inv g8340
timestamp 1386238110
transform 1 0 12171 0 1 7515
box 0 0 120 799
use and2 rm_assigns_buf_StatusReg_1
timestamp 1386234845
transform 1 0 12291 0 1 7515
box 0 0 120 799
use buffer g8399
timestamp 1386236986
transform 1 0 12411 0 1 7515
box 0 0 120 799
use and2 g8074
timestamp 1386234845
transform 1 0 12531 0 1 7515
box 0 0 120 799
use nor2 g8209
timestamp 1386235306
transform 1 0 12651 0 1 7515
box 0 0 120 799
use nand2 g8103
timestamp 1386234792
transform 1 0 12771 0 1 7515
box 0 0 96 799
use nand2 g8268
timestamp 1386234792
transform 1 0 12867 0 1 7515
box 0 0 96 799
use nand2 g8283
timestamp 1386234792
transform 1 0 12963 0 1 7515
box 0 0 96 799
use nand2 g8411
timestamp 1386234792
transform 1 0 13059 0 1 7515
box 0 0 96 799
use nand2 g8321
timestamp 1386234792
transform 1 0 13155 0 1 7515
box 0 0 96 799
use nor2 g8379
timestamp 1386235306
transform 1 0 13251 0 1 7515
box 0 0 120 799
use and2 g8180
timestamp 1386234845
transform 1 0 13371 0 1 7515
box 0 0 120 799
use nand4 g8052
timestamp 1386234936
transform 1 0 13491 0 1 7515
box 0 0 144 799
use nand3 g8136
timestamp 1396952988
transform 1 0 13635 0 1 7515
box 0 0 120 799
use and2 g8110
timestamp 1386234845
transform 1 0 13755 0 1 7515
box 0 0 120 799
use nand2 g8153
timestamp 1386234792
transform 1 0 13875 0 1 7515
box 0 0 96 799
use nand3 g8361
timestamp 1396952988
transform 1 0 13971 0 1 7515
box 0 0 120 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 14091 0 1 7515
box 0 0 96 799
use scandtype g8308
timestamp 1386241841
transform 1 0 14187 0 1 7515
box 0 0 624 799
use nand2 stateSub_reg_91_2_93_
timestamp 1386234792
transform 1 0 14811 0 1 7515
box 0 0 96 799
use scandtype g8372
timestamp 1386241841
transform 1 0 14907 0 1 7515
box 0 0 624 799
use and2 g8294
timestamp 1386234845
transform 1 0 15531 0 1 7515
box 0 0 120 799
use and2 g8099
timestamp 1386234845
transform 1 0 15651 0 1 7515
box 0 0 120 799
use nand2 g8420
timestamp 1386234792
transform 1 0 15771 0 1 7515
box 0 0 96 799
use inv g8190
timestamp 1386238110
transform 1 0 15867 0 1 7515
box 0 0 120 799
use and2 g8045
timestamp 1386234845
transform 1 0 15987 0 1 7515
box 0 0 120 799
use nand2 g8304
timestamp 1386234792
transform 1 0 16107 0 1 7515
box 0 0 96 799
use rowcrosser RegWe
timestamp 1386086759
transform 1 0 16203 0 1 7515
box 0 0 48 799
use nand2 g8092
timestamp 1386234792
transform 1 0 16251 0 1 7515
box 0 0 96 799
use nand4 g8277
timestamp 1386234936
transform 1 0 16347 0 1 7515
box 0 0 144 799
use and2 g8081
timestamp 1386234845
transform 1 0 16491 0 1 7515
box 0 0 120 799
use nand3 g8243
timestamp 1396952988
transform 1 0 16611 0 1 7515
box 0 0 120 799
use nand2 g8296
timestamp 1386234792
transform 1 0 16731 0 1 7515
box 0 0 96 799
use nand2 g8348
timestamp 1386234792
transform 1 0 16827 0 1 7515
box 0 0 96 799
use rowcrosser MemEn
timestamp 1386086759
transform 1 0 16923 0 1 7515
box 0 0 48 799
use inv g8234
timestamp 1386238110
transform 1 0 16971 0 1 7515
box 0 0 120 799
use and2 StatusReg_reg_91_1_93_
timestamp 1386234845
transform 1 0 17091 0 1 7515
box 0 0 120 799
use scandtype g8324
timestamp 1386241841
transform 1 0 17211 0 1 7515
box 0 0 624 799
use nand2 g8293
timestamp 1386234792
transform 1 0 17835 0 1 7515
box 0 0 96 799
use nand2 g8312
timestamp 1386234792
transform 1 0 17931 0 1 7515
box 0 0 96 799
use nor2 g8213
timestamp 1386235306
transform 1 0 18027 0 1 7515
box 0 0 120 799
use nand2 g8096
timestamp 1386234792
transform 1 0 18147 0 1 7515
box 0 0 96 799
use nand2 g8212
timestamp 1386234792
transform 1 0 18243 0 1 7515
box 0 0 96 799
use nand2 g8084
timestamp 1386234792
transform 1 0 18339 0 1 7515
box 0 0 96 799
use nand3 g8265
timestamp 1396952988
transform 1 0 18435 0 1 7515
box 0 0 120 799
use inv g8200
timestamp 1386238110
transform 1 0 18555 0 1 7515
box 0 0 120 799
use and2 g8400
timestamp 1386234845
transform 1 0 18675 0 1 7515
box 0 0 120 799
use nand2 g8108
timestamp 1386234792
transform 1 0 18795 0 1 7515
box 0 0 96 799
use nand2 g8049
timestamp 1386234792
transform 1 0 18891 0 1 7515
box 0 0 96 799
use nor2 g8144
timestamp 1386235306
transform 1 0 18987 0 1 7515
box 0 0 120 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 19107 0 1 7515
box 0 0 48 799
use nand2 g8159
timestamp 1386234792
transform 1 0 19155 0 1 7515
box 0 0 96 799
use nor2 g8177
timestamp 1386235306
transform 1 0 19251 0 1 7515
box 0 0 120 799
use nand3 g8356
timestamp 1396952988
transform 1 0 19371 0 1 7515
box 0 0 120 799
use nand2 g8251
timestamp 1386234792
transform 1 0 19491 0 1 7515
box 0 0 96 799
use nand2 g8226
timestamp 1386234792
transform 1 0 19587 0 1 7515
box 0 0 96 799
use nand3 g8264
timestamp 1396952988
transform 1 0 19683 0 1 7515
box 0 0 120 799
use nand2 g8332
timestamp 1386234792
transform 1 0 19803 0 1 7515
box 0 0 96 799
use nand2 g8089
timestamp 1386234792
transform 1 0 19899 0 1 7515
box 0 0 96 799
use nand4 g8206
timestamp 1386234936
transform 1 0 19995 0 1 7515
box 0 0 144 799
use nor2 g8237
timestamp 1386235306
transform 1 0 20139 0 1 7515
box 0 0 120 799
use rowcrosser LrSel
timestamp 1386086759
transform 1 0 20259 0 1 7515
box 0 0 48 799
use nand2 g8278
timestamp 1386234792
transform 1 0 20307 0 1 7515
box 0 0 96 799
use nand2 g8376
timestamp 1386234792
transform 1 0 20403 0 1 7515
box 0 0 96 799
use nand2 g8181
timestamp 1386234792
transform 1 0 20499 0 1 7515
box 0 0 96 799
use nand2 g8216
timestamp 1386234792
transform 1 0 20595 0 1 7515
box 0 0 96 799
use nand3 StatusReg_reg_91_0_93_
timestamp 1396952988
transform 1 0 20691 0 1 7515
box 0 0 120 799
use scandtype g8253
timestamp 1386241841
transform 1 0 20811 0 1 7515
box 0 0 624 799
use rowcrosser AluOR_91_1_93_
timestamp 1386086759
transform 1 0 21435 0 1 7515
box 0 0 48 799
use nand2 g8373
timestamp 1386234792
transform 1 0 21483 0 1 7515
box 0 0 96 799
use and2 g8186
timestamp 1386234845
transform 1 0 21579 0 1 7515
box 0 0 120 799
use rowcrosser Op2Sel_91_1_93_
timestamp 1386086759
transform 1 0 21699 0 1 7515
box 0 0 48 799
use nand3 g8424
timestamp 1396952988
transform 1 0 21747 0 1 7515
box 0 0 120 799
use inv g8432
timestamp 1386238110
transform 1 0 21867 0 1 7515
box 0 0 120 799
use inv g8090
timestamp 1386238110
transform 1 0 21987 0 1 7515
box 0 0 120 799
use inv g8223
timestamp 1386238110
transform 1 0 22107 0 1 7515
box 0 0 120 799
use nand3 g8195
timestamp 1396952988
transform 1 0 22227 0 1 7515
box 0 0 120 799
use nand2 g8077
timestamp 1386234792
transform 1 0 22347 0 1 7515
box 0 0 96 799
use inv g8410
timestamp 1386238110
transform 1 0 22443 0 1 7515
box 0 0 120 799
use nand2 g8133
timestamp 1386234792
transform 1 0 22563 0 1 7515
box 0 0 96 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 22659 0 1 7515
box 0 0 48 799
use and2 g8341
timestamp 1386234845
transform 1 0 22707 0 1 7515
box 0 0 120 799
use nand2 g8406
timestamp 1386234792
transform 1 0 22827 0 1 7515
box 0 0 96 799
use nand2 g8289
timestamp 1386234792
transform 1 0 22923 0 1 7515
box 0 0 96 799
use nand2 g8128
timestamp 1386234792
transform 1 0 23019 0 1 7515
box 0 0 96 799
use nor2 g8397
timestamp 1386235306
transform 1 0 23115 0 1 7515
box 0 0 120 799
use nand2 g8100
timestamp 1386234792
transform 1 0 23235 0 1 7515
box 0 0 96 799
use nand4 g8350
timestamp 1386234936
transform 1 0 23331 0 1 7515
box 0 0 144 799
use and2 g8117
timestamp 1386234845
transform 1 0 23475 0 1 7515
box 0 0 120 799
use inv g8167
timestamp 1386238110
transform 1 0 23595 0 1 7515
box 0 0 120 799
use nand2 g8191
timestamp 1386234792
transform 1 0 23715 0 1 7515
box 0 0 96 799
use nand2 g8227
timestamp 1386234792
transform 1 0 23811 0 1 7515
box 0 0 96 799
use nand3 g8387
timestamp 1396952988
transform 1 0 23907 0 1 7515
box 0 0 120 799
use and2 g8270
timestamp 1386234845
transform 1 0 24027 0 1 7515
box 0 0 120 799
use nand2 g8073
timestamp 1386234792
transform 1 0 24147 0 1 7515
box 0 0 96 799
use nand3 g8163
timestamp 1396952988
transform 1 0 24243 0 1 7515
box 0 0 120 799
use nor2 g8273
timestamp 1386235306
transform 1 0 24363 0 1 7515
box 0 0 120 799
use nand2 g8337
timestamp 1386234792
transform 1 0 24483 0 1 7515
box 0 0 96 799
use xor2 g8051
timestamp 1396952988
transform 1 0 24579 0 1 7515
box 0 0 192 799
use nand3 g8147
timestamp 1396952988
transform 1 0 24771 0 1 7515
box 0 0 120 799
use nand4 g8353
timestamp 1386234936
transform 1 0 24891 0 1 7515
box 0 0 144 799
use nand2 g8367
timestamp 1386234792
transform 1 0 25035 0 1 7515
box 0 0 96 799
use nand2 g8248
timestamp 1386234792
transform 1 0 25131 0 1 7515
box 0 0 96 799
use nand2 g8114
timestamp 1386234792
transform 1 0 25227 0 1 7515
box 0 0 96 799
use nand3 g8174
timestamp 1396952988
transform 1 0 25323 0 1 7515
box 0 0 120 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 25443 0 1 7515
box 0 0 48 799
use nand4 g8393
timestamp 1386234936
transform 1 0 25491 0 1 7515
box 0 0 144 799
use nand2 g8305
timestamp 1386234792
transform 1 0 25635 0 1 7515
box 0 0 96 799
use nand3 g8241
timestamp 1396952988
transform 1 0 25731 0 1 7515
box 0 0 120 799
use nand2 g8382
timestamp 1386234792
transform 1 0 25851 0 1 7515
box 0 0 96 799
use nand2 g8158
timestamp 1386234792
transform 1 0 25947 0 1 7515
box 0 0 96 799
use nand2 g8063
timestamp 1386234792
transform 1 0 26043 0 1 7515
box 0 0 96 799
use nand2 g8257
timestamp 1386234792
transform 1 0 26139 0 1 7515
box 0 0 96 799
use nand3 ENB
timestamp 1396952988
transform 1 0 26235 0 1 7515
box 0 0 120 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 26355 0 1 7515
box 0 0 48 799
use rowcrosser Op2Sel_91_0_93_
timestamp 1386086759
transform 1 0 26403 0 1 7515
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 26451 0 1 7515
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 994
box 0 0 1464 799
use scandtype g8409
timestamp 1386241841
transform 1 0 1587 0 1 994
box 0 0 624 799
use nand2 g8352
timestamp 1386234792
transform 1 0 2211 0 1 994
box 0 0 96 799
use nand2 g8430
timestamp 1386234792
transform 1 0 2307 0 1 994
box 0 0 96 799
use inv g8150
timestamp 1386238110
transform 1 0 2403 0 1 994
box 0 0 120 799
use nand4 g8250
timestamp 1386234936
transform 1 0 2523 0 1 994
box 0 0 144 799
use inv state_reg_91_1_93_
timestamp 1386238110
transform 1 0 2667 0 1 994
box 0 0 120 799
use scandtype g8416
timestamp 1386241841
transform 1 0 2787 0 1 994
box 0 0 624 799
use inv g8148
timestamp 1386238110
transform 1 0 3411 0 1 994
box 0 0 120 799
use inv g8211
timestamp 1386238110
transform 1 0 3531 0 1 994
box 0 0 120 799
use inv g8196
timestamp 1386238110
transform 1 0 3651 0 1 994
box 0 0 120 799
use nand2 g8359
timestamp 1386234792
transform 1 0 3771 0 1 994
box 0 0 96 799
use nand2 g8300
timestamp 1386234792
transform 1 0 3867 0 1 994
box 0 0 96 799
use nand2 g8175
timestamp 1386234792
transform 1 0 3963 0 1 994
box 0 0 96 799
use nand2 g8078
timestamp 1386234792
transform 1 0 4059 0 1 994
box 0 0 96 799
use nand3 g8388
timestamp 1396952988
transform 1 0 4155 0 1 994
box 0 0 120 799
use nand2 g8093
timestamp 1386234792
transform 1 0 4275 0 1 994
box 0 0 96 799
use nand2 g8429
timestamp 1386234792
transform 1 0 4371 0 1 994
box 0 0 96 799
use inv g8104
timestamp 1386238110
transform 1 0 4467 0 1 994
box 0 0 120 799
use nand2 g8391
timestamp 1386234792
transform 1 0 4587 0 1 994
box 0 0 96 799
use inv g8307
timestamp 1386238110
transform 1 0 4683 0 1 994
box 0 0 120 799
use inv g8389
timestamp 1386238110
transform 1 0 4803 0 1 994
box 0 0 120 799
use nand2 g8335
timestamp 1386234792
transform 1 0 4923 0 1 994
box 0 0 96 799
use nand3 g8160
timestamp 1396952988
transform 1 0 5019 0 1 994
box 0 0 120 799
use nand2 g8076
timestamp 1386234792
transform 1 0 5139 0 1 994
box 0 0 96 799
use nand4 StatusReg_reg_91_2_93_
timestamp 1386234936
transform 1 0 5235 0 1 994
box 0 0 144 799
use scandtype g8161
timestamp 1386241841
transform 1 0 5379 0 1 994
box 0 0 624 799
use nand2 g8224
timestamp 1386234792
transform 1 0 6003 0 1 994
box 0 0 96 799
use nand3 g8094
timestamp 1396952988
transform 1 0 6099 0 1 994
box 0 0 120 799
use nand2 g8266
timestamp 1386234792
transform 1 0 6219 0 1 994
box 0 0 96 799
use nor2 g8401
timestamp 1386235306
transform 1 0 6315 0 1 994
box 0 0 120 799
use inv g8189
timestamp 1386238110
transform 1 0 6435 0 1 994
box 0 0 120 799
use nor2 g8125
timestamp 1386235306
transform 1 0 6555 0 1 994
box 0 0 120 799
use nor2 g8297
timestamp 1386235306
transform 1 0 6675 0 1 994
box 0 0 120 799
use inv g8232
timestamp 1386238110
transform 1 0 6795 0 1 994
box 0 0 120 799
use nand2 g8152
timestamp 1386234792
transform 1 0 6915 0 1 994
box 0 0 96 799
use nand4 g8303
timestamp 1386234936
transform 1 0 7011 0 1 994
box 0 0 144 799
use nand2 g8328
timestamp 1386234792
transform 1 0 7155 0 1 994
box 0 0 96 799
use nand2 g8394
timestamp 1386234792
transform 1 0 7251 0 1 994
box 0 0 96 799
use inv g8080
timestamp 1386238110
transform 1 0 7347 0 1 994
box 0 0 120 799
use rowcrosser g8182
timestamp 1386086759
transform 1 0 7467 0 1 994
box 0 0 48 799
use nand3 g8395
timestamp 1396952988
transform 1 0 7515 0 1 994
box 0 0 120 799
use nand2 g8282
timestamp 1386234792
transform 1 0 7635 0 1 994
box 0 0 96 799
use nand3 g8267
timestamp 1396952988
transform 1 0 7731 0 1 994
box 0 0 120 799
use nand2 g8274
timestamp 1386234792
transform 1 0 7851 0 1 994
box 0 0 96 799
use nand2 g8236
timestamp 1386234792
transform 1 0 7947 0 1 994
box 0 0 96 799
use nand2 g8101
timestamp 1386234792
transform 1 0 8043 0 1 994
box 0 0 96 799
use nand2 g8349
timestamp 1386234792
transform 1 0 8139 0 1 994
box 0 0 96 799
use nor2 g8412
timestamp 1386235306
transform 1 0 8235 0 1 994
box 0 0 120 799
use inv g8185
timestamp 1386238110
transform 1 0 8355 0 1 994
box 0 0 120 799
use nand3 g8365
timestamp 1396952988
transform 1 0 8475 0 1 994
box 0 0 120 799
use nand2 g8255
timestamp 1386234792
transform 1 0 8595 0 1 994
box 0 0 96 799
use and2 g8301
timestamp 1386234845
transform 1 0 8691 0 1 994
box 0 0 120 799
use and2 g8086
timestamp 1386234845
transform 1 0 8811 0 1 994
box 0 0 120 799
use nand2 g8192
timestamp 1386234792
transform 1 0 8931 0 1 994
box 0 0 96 799
use inv g8292
timestamp 1386238110
transform 1 0 9027 0 1 994
box 0 0 120 799
use inv g8254
timestamp 1386238110
transform 1 0 9147 0 1 994
box 0 0 120 799
use and2 g8116
timestamp 1386234845
transform 1 0 9267 0 1 994
box 0 0 120 799
use nand3 g8166
timestamp 1396952988
transform 1 0 9387 0 1 994
box 0 0 120 799
use nand2 g8145
timestamp 1386234792
transform 1 0 9507 0 1 994
box 0 0 96 799
use inv g8426
timestamp 1386238110
transform 1 0 9603 0 1 994
box 0 0 120 799
use inv g8315
timestamp 1386238110
transform 1 0 9723 0 1 994
box 0 0 120 799
use nor2 g8228
timestamp 1386235306
transform 1 0 9843 0 1 994
box 0 0 120 799
use and2 g8342
timestamp 1386234845
transform 1 0 9963 0 1 994
box 0 0 120 799
use and2 g8072
timestamp 1386234845
transform 1 0 10083 0 1 994
box 0 0 120 799
use nand3 g8279
timestamp 1396952988
transform 1 0 10203 0 1 994
box 0 0 120 799
use nand2 g8259
timestamp 1386234792
transform 1 0 10323 0 1 994
box 0 0 96 799
use inv g8105
timestamp 1386238110
transform 1 0 10419 0 1 994
box 0 0 120 799
use nand2 g8375
timestamp 1386234792
transform 1 0 10539 0 1 994
box 0 0 96 799
use inv g8122
timestamp 1386238110
transform 1 0 10635 0 1 994
box 0 0 120 799
use nand2 g8446
timestamp 1386234792
transform 1 0 10755 0 1 994
box 0 0 96 799
use nand3 g8059
timestamp 1396952988
transform 1 0 10851 0 1 994
box 0 0 120 799
use nand4 g8097
timestamp 1386234936
transform 1 0 10971 0 1 994
box 0 0 144 799
use nand4 g8062
timestamp 1386234936
transform 1 0 11115 0 1 994
box 0 0 144 799
use nand2 g8247
timestamp 1386234792
transform 1 0 11259 0 1 994
box 0 0 96 799
use and2 g8263
timestamp 1386234845
transform 1 0 11355 0 1 994
box 0 0 120 799
use nand3 IntStatus_reg
timestamp 1396952988
transform 1 0 11475 0 1 994
box 0 0 120 799
use scanreg g8256
timestamp 1386241447
transform 1 0 11595 0 1 994
box 0 0 720 799
use nand2 g8131
timestamp 1386234792
transform 1 0 12315 0 1 994
box 0 0 96 799
use nand2 g8087
timestamp 1386234792
transform 1 0 12411 0 1 994
box 0 0 96 799
use nand3 g8345
timestamp 1396952988
transform 1 0 12507 0 1 994
box 0 0 120 799
use nand2 g8322
timestamp 1386234792
transform 1 0 12627 0 1 994
box 0 0 96 799
use nand2 g8286
timestamp 1386234792
transform 1 0 12723 0 1 994
box 0 0 96 799
use nand2 g8368
timestamp 1386234792
transform 1 0 12819 0 1 994
box 0 0 96 799
use nand2 g8137
timestamp 1386234792
transform 1 0 12915 0 1 994
box 0 0 96 799
use nand3 g8201
timestamp 1396952988
transform 1 0 13011 0 1 994
box 0 0 120 799
use nand2 g8331
timestamp 1386234792
transform 1 0 13131 0 1 994
box 0 0 96 799
use nand2 g8336
timestamp 1386234792
transform 1 0 13227 0 1 994
box 0 0 96 799
use nand2 g8242
timestamp 1386234792
transform 1 0 13323 0 1 994
box 0 0 96 799
use nand2 g8207
timestamp 1386234792
transform 1 0 13419 0 1 994
box 0 0 96 799
use nand2 g8383
timestamp 1386234792
transform 1 0 13515 0 1 994
box 0 0 96 799
use nand2 g8405
timestamp 1386234792
transform 1 0 13611 0 1 994
box 0 0 96 799
use inv g8173
timestamp 1386238110
transform 1 0 13707 0 1 994
box 0 0 120 799
use nand2 g8398
timestamp 1386234792
transform 1 0 13827 0 1 994
box 0 0 96 799
use nand2 g8157
timestamp 1386234792
transform 1 0 13923 0 1 994
box 0 0 96 799
use nand3 g8325
timestamp 1396952988
transform 1 0 14019 0 1 994
box 0 0 120 799
use nand2 g8140
timestamp 1386234792
transform 1 0 14139 0 1 994
box 0 0 96 799
use and2 g8210
timestamp 1386234845
transform 1 0 14235 0 1 994
box 0 0 120 799
use nand2 g8141
timestamp 1386234792
transform 1 0 14355 0 1 994
box 0 0 96 799
use nand2 g8203
timestamp 1386234792
transform 1 0 14451 0 1 994
box 0 0 96 799
use nand2 g8065
timestamp 1386234792
transform 1 0 14547 0 1 994
box 0 0 96 799
use nor2 g8404
timestamp 1386235306
transform 1 0 14643 0 1 994
box 0 0 120 799
use nand2 g8413
timestamp 1386234792
transform 1 0 14763 0 1 994
box 0 0 96 799
use nand2 g8113
timestamp 1386234792
transform 1 0 14859 0 1 994
box 0 0 96 799
use nand3 g8358
timestamp 1396952988
transform 1 0 14955 0 1 994
box 0 0 120 799
use nand2 g8070
timestamp 1386234792
transform 1 0 15075 0 1 994
box 0 0 96 799
use nand2 g8323
timestamp 1386234792
transform 1 0 15171 0 1 994
box 0 0 96 799
use nand2 g8408
timestamp 1386234792
transform 1 0 15267 0 1 994
box 0 0 96 799
use nand2 g8309
timestamp 1386234792
transform 1 0 15363 0 1 994
box 0 0 96 799
use nand3 g8380
timestamp 1396952988
transform 1 0 15459 0 1 994
box 0 0 120 799
use nand2 g8233
timestamp 1386234792
transform 1 0 15579 0 1 994
box 0 0 96 799
use and2 IRQ2_reg
timestamp 1386234845
transform 1 0 15675 0 1 994
box 0 0 120 799
use scandtype g8151
timestamp 1386241841
transform 1 0 15795 0 1 994
box 0 0 624 799
use nor2 g8138
timestamp 1386235306
transform 1 0 16419 0 1 994
box 0 0 120 799
use nand2 g8402
timestamp 1386234792
transform 1 0 16539 0 1 994
box 0 0 96 799
use nand2 g8188
timestamp 1386234792
transform 1 0 16635 0 1 994
box 0 0 96 799
use nand4 g8176
timestamp 1386234936
transform 1 0 16731 0 1 994
box 0 0 144 799
use nand2 g8172
timestamp 1386234792
transform 1 0 16875 0 1 994
box 0 0 96 799
use nand2 g8422
timestamp 1386234792
transform 1 0 16971 0 1 994
box 0 0 96 799
use inv g8162
timestamp 1386238110
transform 1 0 17067 0 1 994
box 0 0 120 799
use inv g8415
timestamp 1386238110
transform 1 0 17187 0 1 994
box 0 0 120 799
use nand2 g8095
timestamp 1386234792
transform 1 0 17307 0 1 994
box 0 0 96 799
use nand2 g8299
timestamp 1386234792
transform 1 0 17403 0 1 994
box 0 0 96 799
use nand2 g8126
timestamp 1386234792
transform 1 0 17499 0 1 994
box 0 0 96 799
use and2 g8326
timestamp 1386234845
transform 1 0 17595 0 1 994
box 0 0 120 799
use nand2 g8396
timestamp 1386234792
transform 1 0 17715 0 1 994
box 0 0 96 799
use nor2 IRQ1_reg
timestamp 1386235306
transform 1 0 17811 0 1 994
box 0 0 120 799
use scandtype g8329
timestamp 1386241841
transform 1 0 17931 0 1 994
box 0 0 624 799
use inv rm_assigns_buf_MemEn
timestamp 1386238110
transform 1 0 18555 0 1 994
box 0 0 120 799
use buffer g8205
timestamp 1386236986
transform 1 0 18675 0 1 994
box 0 0 120 799
use nand2 g8339
timestamp 1386234792
transform 1 0 18795 0 1 994
box 0 0 96 799
use nand2 g8164
timestamp 1386234792
transform 1 0 18891 0 1 994
box 0 0 96 799
use nor2 g8245
timestamp 1386235306
transform 1 0 18987 0 1 994
box 0 0 120 799
use nor2 g8260
timestamp 1386235306
transform 1 0 19107 0 1 994
box 0 0 120 799
use nand2 g8165
timestamp 1386234792
transform 1 0 19227 0 1 994
box 0 0 96 799
use nor2 g8351
timestamp 1386235306
transform 1 0 19323 0 1 994
box 0 0 120 799
use nor2 g3
timestamp 1386235306
transform 1 0 19443 0 1 994
box 0 0 120 799
use inv g8215
timestamp 1386238110
transform 1 0 19563 0 1 994
box 0 0 120 799
use nand2 g8343
timestamp 1386234792
transform 1 0 19683 0 1 994
box 0 0 96 799
use inv g8288
timestamp 1386238110
transform 1 0 19779 0 1 994
box 0 0 120 799
use nand2 g8239
timestamp 1386234792
transform 1 0 19899 0 1 994
box 0 0 96 799
use nand2 g8079
timestamp 1386234792
transform 1 0 19995 0 1 994
box 0 0 96 799
use nand3 g8384
timestamp 1396952988
transform 1 0 20091 0 1 994
box 0 0 120 799
use nand2 g8262
timestamp 1386234792
transform 1 0 20211 0 1 994
box 0 0 96 799
use nand3 g8311
timestamp 1396952988
transform 1 0 20307 0 1 994
box 0 0 120 799
use nand3 g8109
timestamp 1396952988
transform 1 0 20427 0 1 994
box 0 0 120 799
use nand2 g8085
timestamp 1386234792
transform 1 0 20547 0 1 994
box 0 0 96 799
use nand2 g8298
timestamp 1386234792
transform 1 0 20643 0 1 994
box 0 0 96 799
use nand3 g8346
timestamp 1396952988
transform 1 0 20739 0 1 994
box 0 0 120 799
use nand3 g8184
timestamp 1396952988
transform 1 0 20859 0 1 994
box 0 0 120 799
use inv g8132
timestamp 1386238110
transform 1 0 20979 0 1 994
box 0 0 120 799
use nand3 g8355
timestamp 1396952988
transform 1 0 21099 0 1 994
box 0 0 120 799
use nand2 g8385
timestamp 1386234792
transform 1 0 21219 0 1 994
box 0 0 96 799
use inv g8219
timestamp 1386238110
transform 1 0 21315 0 1 994
box 0 0 120 799
use nand3 g8330
timestamp 1396952988
transform 1 0 21435 0 1 994
box 0 0 120 799
use nand2 g8061
timestamp 1386234792
transform 1 0 21555 0 1 994
box 0 0 96 799
use nand2 g8360
timestamp 1386234792
transform 1 0 21651 0 1 994
box 0 0 96 799
use nand2 g8258
timestamp 1386234792
transform 1 0 21747 0 1 994
box 0 0 96 799
use nand2 g8115
timestamp 1386234792
transform 1 0 21843 0 1 994
box 0 0 96 799
use nand2 g8202
timestamp 1386234792
transform 1 0 21939 0 1 994
box 0 0 96 799
use nand2 g8246
timestamp 1386234792
transform 1 0 22035 0 1 994
box 0 0 96 799
use nand2 g8208
timestamp 1386234792
transform 1 0 22131 0 1 994
box 0 0 96 799
use nand2 g8231
timestamp 1386234792
transform 1 0 22227 0 1 994
box 0 0 96 799
use nand2 g8156
timestamp 1386234792
transform 1 0 22323 0 1 994
box 0 0 96 799
use nor2 g8179
timestamp 1386235306
transform 1 0 22419 0 1 994
box 0 0 120 799
use nand2 g8371
timestamp 1386234792
transform 1 0 22539 0 1 994
box 0 0 96 799
use nand2 g8193
timestamp 1386234792
transform 1 0 22635 0 1 994
box 0 0 96 799
use nand2 g8071
timestamp 1386234792
transform 1 0 22731 0 1 994
box 0 0 96 799
use nand4 g8285
timestamp 1386234936
transform 1 0 22827 0 1 994
box 0 0 144 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 22971 0 1 994
box 0 0 48 799
use nand2 g8083
timestamp 1386234792
transform 1 0 23019 0 1 994
box 0 0 96 799
use nand3 g8204
timestamp 1396952988
transform 1 0 23115 0 1 994
box 0 0 120 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 23235 0 1 994
box 0 0 96 799
use scandtype g8053
timestamp 1386241841
transform 1 0 23331 0 1 994
box 0 0 624 799
use nand4 g8302
timestamp 1386234936
transform 1 0 23955 0 1 994
box 0 0 144 799
use nand2 g8142
timestamp 1386234792
transform 1 0 24099 0 1 994
box 0 0 96 799
use nand2 stateSub_reg_91_1_93_
timestamp 1386234792
transform 1 0 24195 0 1 994
box 0 0 96 799
use scandtype g8075
timestamp 1386241841
transform 1 0 24291 0 1 994
box 0 0 624 799
use nand3 g8197
timestamp 1396952988
transform 1 0 24915 0 1 994
box 0 0 120 799
use nand2 g8316
timestamp 1386234792
transform 1 0 25035 0 1 994
box 0 0 96 799
use nand2 g8378
timestamp 1386234792
transform 1 0 25131 0 1 994
box 0 0 96 799
use nand2 g8291
timestamp 1386234792
transform 1 0 25227 0 1 994
box 0 0 96 799
use nand2 g8112
timestamp 1386234792
transform 1 0 25323 0 1 994
box 0 0 96 799
use inv g8445
timestamp 1386238110
transform 1 0 25419 0 1 994
box 0 0 120 799
use inv g8060
timestamp 1386238110
transform 1 0 25539 0 1 994
box 0 0 120 799
use nand4 SysBus_91_3_93_
timestamp 1386234936
transform 1 0 25659 0 1 994
box 0 0 144 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 26450 0 1 994
box 0 0 320 799
<< labels >>
rlabel m2contact 26553 8451 26553 8451 6 RwSel[1]
rlabel m2contact 26553 8331 26553 8331 6 RwSel[1]
rlabel m2contact 26529 8379 26529 8379 6 AluOR[0]
rlabel m2contact 26529 8331 26529 8331 6 AluOR[0]
rlabel m2contact 26505 8403 26505 8403 6 AluOR[1]
rlabel m2contact 26505 8379 26505 8379 6 AluOR[1]
rlabel m2contact 26481 8427 26481 8427 6 ENB
rlabel m2contact 26481 8403 26481 8403 6 ENB
rlabel m2contact 26457 8427 26457 8427 6 RegWe
rlabel m2contact 26457 8355 26457 8355 6 RegWe
rlabel m2contact 26433 8379 26433 8379 6 AluOR[1]
rlabel m2contact 26385 8427 26385 8427 6 RegWe
rlabel m2contact 26193 8523 26193 8523 6 StatusReg[2]
rlabel m2contact 25473 8499 25473 8499 6 Op2Sel[1]
rlabel m2contact 25437 8379 25437 8379 6 StatusRegEn
rlabel m2contact 25161 8355 25161 8355 6 StatusReg[3]
rlabel m2contact 24873 8571 24873 8571 6 AluEn
rlabel m2contact 24621 8427 24621 8427 6 StatusReg[0]
rlabel m2contact 24345 8547 24345 8547 6 AluWe
rlabel m2contact 23805 8475 23805 8475 6 StatusReg[1]
rlabel m2contact 23781 8523 23781 8523 6 StatusReg[2]
rlabel m2contact 23217 8523 23217 8523 6 Op1Sel
rlabel m2contact 22689 8331 22689 8331 6 AluOR[0]
rlabel m2contact 22173 8355 22173 8355 6 StatusReg[3]
rlabel m2contact 22149 8571 22149 8571 6 AluEn
rlabel m2contact 21729 8379 21729 8379 6 StatusRegEn
rlabel m2contact 21465 8403 21465 8403 6 ENB
rlabel m2contact 21333 8547 21333 8547 6 AluWe
rlabel m2contact 21321 8427 21321 8427 6 StatusReg[0]
rlabel metal2 20307 8427 20307 8427 6 Op2Sel[0]
rlabel m2contact 20289 8427 20289 8427 6 Op2Sel[0]
rlabel m2contact 19701 8499 19701 8499 6 Op2Sel[1]
rlabel m2contact 19137 8571 19137 8571 6 MemEn
rlabel m2contact 18969 8499 18969 8499 6 PcSel[0]
rlabel m2contact 18885 8523 18885 8523 6 Op1Sel
rlabel m2contact 18537 8451 18537 8451 6 RwSel[1]
rlabel m2contact 17277 8451 17277 8451 6 WdSel
rlabel m2contact 16953 8451 16953 8451 6 WdSel
rlabel m2contact 16461 8547 16461 8547 6 PcEn
rlabel metal2 16251 8451 16251 8451 6 PcWe
rlabel m2contact 16233 8451 16233 8451 6 PcWe
rlabel m2contact 15621 8499 15621 8499 6 PcSel[0]
rlabel m2contact 14697 8355 14697 8355 6 StatusReg[3]
rlabel m2contact 14013 8403 14013 8403 6 PcSel[1]
rlabel m2contact 13953 8499 13953 8499 6 LrEn
rlabel m2contact 13197 8523 13197 8523 4 PcSel[2]
rlabel m2contact 13161 8499 13161 8499 4 LrEn
rlabel m2contact 12489 8475 12489 8475 4 StatusReg[1]
rlabel m2contact 11541 8427 11541 8427 4 LrWe
rlabel metal2 11211 8475 11211 8475 4 LrSel
rlabel m2contact 11193 8475 11193 8475 4 LrSel
rlabel m2contact 10929 8475 10929 8475 4 ALE
rlabel m2contact 10617 8499 10617 8499 4 OpcodeCondIn[4]
rlabel metal2 10443 8451 10443 8451 4 ImmSel
rlabel m2contact 10425 8451 10425 8451 4 ImmSel
rlabel m2contact 10377 8451 10377 8451 4 nME
rlabel metal2 9531 8379 9531 8379 4 IrWe
rlabel m2contact 9513 8379 9513 8379 4 IrWe
rlabel m2contact 9249 8427 9249 8427 4 LrWe
rlabel m2contact 9021 8571 9021 8571 4 MemEn
rlabel m2contact 8721 8379 8721 8379 4 OpcodeCondIn[3]
rlabel m2contact 7401 8427 7401 8427 4 OpcodeCondIn[0]
rlabel metal2 6819 8571 6819 8571 4 OpcodeCondIn[1]
rlabel m2contact 6801 8571 6801 8571 4 OpcodeCondIn[1]
rlabel m2contact 6777 8427 6777 8427 4 OpcodeCondIn[0]
rlabel m2contact 6465 8427 6465 8427 4 OpcodeCondIn[5]
rlabel m2contact 6393 8403 6393 8403 4 PcSel[1]
rlabel m2contact 5745 8403 5745 8403 4 OpcodeCondIn[2]
rlabel m2contact 5721 8355 5721 8355 4 StatusReg[3]
rlabel m2contact 5709 8379 5709 8379 4 OpcodeCondIn[3]
rlabel m2contact 5313 8547 5313 8547 4 PcEn
rlabel m2contact 5049 8523 5049 8523 4 PcSel[2]
rlabel m2contact 4881 8499 4881 8499 4 OpcodeCondIn[4]
rlabel m2contact 4305 8499 4305 8499 4 OpcodeCondIn[6]
rlabel m2contact 4065 8403 4065 8403 4 OpcodeCondIn[2]
rlabel m2contact 4053 8427 4053 8427 4 OpcodeCondIn[5]
rlabel m2contact 3225 8499 3225 8499 4 OpcodeCondIn[6]
rlabel metal2 2331 8499 2331 8499 4 OpcodeCondIn[7]
rlabel m2contact 2313 8499 2313 8499 4 OpcodeCondIn[7]
rlabel m2contact 25617 161 25617 161 8 Flags[0]
rlabel m2contact 25617 41 25617 41 8 Flags[0]
rlabel m2contact 25593 65 25593 65 8 Flags[1]
rlabel m2contact 25593 41 25593 41 8 Flags[1]
rlabel m2contact 25569 89 25569 89 8 Flags[2]
rlabel m2contact 25569 65 25569 65 8 Flags[2]
rlabel m2contact 25569 857 25569 857 6 n_397
rlabel m2contact 25497 881 25497 881 6 n_333
rlabel m2contact 25449 281 25449 281 8 n_320
rlabel m2contact 25401 617 25401 617 8 n_111
rlabel m2contact 24393 521 24393 521 8 n_349
rlabel m2contact 24153 377 24153 377 8 n_39
rlabel m2contact 24009 185 24009 185 8 n_144
rlabel m2contact 23433 689 23433 689 8 n_299
rlabel m2contact 23313 905 23313 905 6 n_169
rlabel m2contact 23145 353 23145 353 8 n_258
rlabel metal2 23019 497 23019 497 8 SysBus[3]
rlabel m2contact 23001 497 23001 497 8 SysBus[3]
rlabel m2contact 22905 833 22905 833 6 n_189
rlabel m2contact 22809 713 22809 713 8 n_246
rlabel m2contact 22401 209 22401 209 8 n_141
rlabel m2contact 22305 473 22305 473 8 n_167
rlabel m2contact 22185 785 22185 785 8 n_104
rlabel m2contact 21825 401 21825 401 8 n_60
rlabel m2contact 21777 137 21777 137 8 n_23
rlabel m2contact 21633 449 21633 449 8 n_68
rlabel m2contact 21153 257 21153 257 8 n_257
rlabel m2contact 21009 497 21009 497 8 n_186
rlabel m2contact 20841 329 20841 329 8 n_91
rlabel m2contact 20673 737 20673 737 8 n_287
rlabel m2contact 20625 665 20625 665 8 n_250
rlabel m2contact 20577 233 20577 233 8 n_198
rlabel m2contact 20289 761 20289 761 8 n_24
rlabel m2contact 20025 545 20025 545 8 n_103
rlabel m2contact 19977 641 19977 641 8 n_95
rlabel m2contact 19953 593 19953 593 8 n_54
rlabel m2contact 19641 569 19641 569 8 n_396
rlabel m2contact 19425 425 19425 425 8 n_271
rlabel m2contact 19305 809 19305 809 6 n_173
rlabel m2contact 18969 593 18969 593 8 n_54
rlabel m2contact 18873 977 18873 977 6 n_237
rlabel m2contact 18585 449 18585 449 8 n_68
rlabel m2contact 18441 953 18441 953 6 IRQ1
rlabel m2contact 18033 113 18033 113 8 n_1
rlabel m2contact 17649 713 17649 713 8 n_246
rlabel m2contact 17553 929 17553 929 6 n_41
rlabel metal2 17475 593 17475 593 8 SysBus[2]
rlabel m2contact 17457 593 17457 593 8 SysBus[2]
rlabel m2contact 17145 593 17145 593 8 n_0
rlabel m2contact 17049 89 17049 89 8 n_267
rlabel m2contact 16953 833 16953 833 6 n_189
rlabel m2contact 16857 833 16857 833 6 n_216
rlabel m2contact 16833 305 16833 305 8 n_16
rlabel m2contact 16593 977 16593 977 6 n_237
rlabel m2contact 15897 953 15897 953 6 IRQ1
rlabel m2contact 15345 929 15345 929 6 n_41
rlabel m2contact 15225 809 15225 809 6 n_173
rlabel m2contact 15057 281 15057 281 8 n_320
rlabel m2contact 15009 89 15009 89 8 n_267
rlabel m2contact 14985 281 14985 281 8 n_243
rlabel m2contact 14481 833 14481 833 6 n_216
rlabel m2contact 14217 89 14217 89 8 n_62
rlabel m2contact 14121 833 14121 833 6 n_259
rlabel m2contact 13857 905 13857 905 6 n_169
rlabel m2contact 13689 137 13689 137 8 n_23
rlabel m2contact 13593 185 13593 185 2 n_144
rlabel m2contact 13473 329 13473 329 2 n_91
rlabel m2contact 13305 377 13305 377 2 n_39
rlabel m2contact 13041 473 13041 473 2 n_167
rlabel m2contact 12609 137 12609 137 2 nWE
rlabel m2contact 12393 473 12393 473 2 n_133
rlabel m2contact 11673 185 11673 185 2 n_266
rlabel m2contact 11409 377 11409 377 2 n_156
rlabel m2contact 11313 17 11313 17 2 CFlag
rlabel m2contact 11049 881 11049 881 4 n_333
rlabel m2contact 10953 857 10953 857 4 n_397
rlabel m2contact 10785 833 10785 833 4 n_259
rlabel m2contact 10593 41 10593 41 2 Flags[1]
rlabel m2contact 10449 809 10449 809 4 n_173
rlabel m2contact 10401 785 10401 785 2 n_104
rlabel m2contact 10377 761 10377 761 2 n_24
rlabel m2contact 10353 89 10353 89 2 n_62
rlabel m2contact 9561 89 9561 89 2 n_161
rlabel m2contact 9489 737 9489 737 2 n_287
rlabel m2contact 9057 713 9057 713 2 n_246
rlabel m2contact 9009 689 9009 689 2 n_299
rlabel m2contact 8961 665 8961 665 2 n_250
rlabel m2contact 8745 641 8745 641 2 n_95
rlabel m2contact 8721 617 8721 617 2 n_111
rlabel m2contact 8649 593 8649 593 2 n_0
rlabel m2contact 8577 497 8577 497 2 n_186
rlabel m2contact 8433 377 8433 377 2 n_156
rlabel m2contact 8217 497 8217 497 2 n_306
rlabel m2contact 8169 569 8169 569 2 n_396
rlabel m2contact 8121 89 8121 89 2 n_161
rlabel m2contact 7833 545 7833 545 2 n_103
rlabel m2contact 7821 89 7821 89 2 SysBus[1]
rlabel m2contact 7617 521 7617 521 2 n_349
rlabel m2contact 7569 497 7569 497 2 n_306
rlabel m2contact 7545 473 7545 473 2 n_133
rlabel m2contact 7497 65 7497 65 2 Flags[2]
rlabel m2contact 7185 449 7185 449 2 n_68
rlabel m2contact 7041 401 7041 401 2 n_60
rlabel m2contact 6825 329 6825 329 2 n_91
rlabel m2contact 6777 329 6777 329 2 n_316
rlabel m2contact 6729 401 6729 401 2 n_215
rlabel m2contact 6705 425 6705 425 2 n_271
rlabel m2contact 6657 401 6657 401 2 n_215
rlabel m2contact 6273 89 6273 89 2 SysBus[1]
rlabel m2contact 6177 377 6177 377 2 n_156
rlabel m2contact 6081 353 6081 353 2 n_258
rlabel m2contact 6033 257 6033 257 2 n_257
rlabel m2contact 5289 329 5289 329 2 n_316
rlabel m2contact 5121 305 5121 305 2 n_16
rlabel m2contact 4641 161 4641 161 2 Flags[0]
rlabel metal2 4443 161 4443 161 2 SysBus[0]
rlabel m2contact 4425 161 4425 161 2 SysBus[0]
rlabel m2contact 4353 161 4353 161 2 n_21
rlabel m2contact 4137 185 4137 185 2 n_266
rlabel m2contact 3993 185 3993 185 2 n_65
rlabel m2contact 3849 281 3849 281 2 n_243
rlabel m2contact 3729 257 3729 257 2 n_257
rlabel m2contact 2649 233 2649 233 2 n_198
rlabel m2contact 2577 209 2577 209 2 n_141
rlabel m2contact 2481 113 2481 113 2 n_1
rlabel m2contact 2433 113 2433 113 2 nIRQ
rlabel m2contact 2385 185 2385 185 2 n_65
rlabel m2contact 2337 161 2337 161 2 n_21
rlabel m2contact 26481 6394 26481 6394 6 Rs1Sel[0]
rlabel m2contact 26481 1834 26481 1834 6 Rs1Sel[0]
rlabel m2contact 26457 3946 26457 3946 6 Flags[3]
rlabel m2contact 26457 1810 26457 1810 6 Flags[3]
rlabel m2contact 26433 2170 26433 2170 6 Rs1Sel[1]
rlabel m2contact 26433 1858 26433 1858 6 Rs1Sel[1]
rlabel m2contact 26433 3178 26433 3178 6 AluOR[1]
rlabel m2contact 26385 4666 26385 4666 6 RegWe
rlabel m2contact 26337 7210 26337 7210 6 n_124
rlabel m2contact 26313 4498 26313 4498 6 OpcodeCondIn[7]
rlabel m2contact 26289 7450 26289 7450 6 n_100
rlabel m2contact 26265 3322 26265 3322 6 n_102
rlabel m2contact 26217 6250 26217 6250 6 n_345
rlabel m2contact 26193 2962 26193 2962 6 StatusReg[2]
rlabel m2contact 26169 6106 26169 6106 6 n_346
rlabel m2contact 26121 3106 26121 3106 6 n_196
rlabel m2contact 26097 3922 26097 3922 6 n_195
rlabel m2contact 26073 5602 26073 5602 6 n_165
rlabel m2contact 26049 5794 26049 5794 6 n_334
rlabel m2contact 26049 3418 26049 3418 6 n_334
rlabel m2contact 26025 4690 26025 4690 6 n_94
rlabel m2contact 26001 5218 26001 5218 6 n_162
rlabel m2contact 25977 6010 25977 6010 6 stateSub[2]
rlabel m2contact 25953 5266 25953 5266 6 n_148
rlabel m2contact 25953 2386 25953 2386 6 n_148
rlabel m2contact 25929 2866 25929 2866 6 n_175
rlabel m2contact 25905 4066 25905 4066 6 n_192
rlabel m2contact 25881 7354 25881 7354 6 n_179
rlabel m2contact 25857 6082 25857 6082 6 stateSub[1]
rlabel m2contact 25857 4594 25857 4594 6 stateSub[1]
rlabel m2contact 25833 2746 25833 2746 6 n_49
rlabel m2contact 25809 4114 25809 4114 6 OpcodeCondIn[2]
rlabel m2contact 25785 4666 25785 4666 6 RegWe
rlabel m2contact 25785 6322 25785 6322 6 n_393
rlabel m2contact 25761 3466 25761 3466 6 n_353
rlabel m2contact 25761 4210 25761 4210 6 n_46
rlabel m2contact 25737 4738 25737 4738 6 n_302
rlabel m2contact 25713 6466 25713 6466 6 n_22
rlabel m2contact 25713 3538 25713 3538 6 n_313
rlabel m2contact 25689 3418 25689 3418 6 n_334
rlabel m2contact 25689 3442 25689 3442 6 n_119
rlabel m2contact 25665 3706 25665 3706 6 state[1]
rlabel m2contact 25641 6202 25641 6202 6 n_310
rlabel m2contact 25641 5122 25641 5122 6 n_310
rlabel m2contact 25617 5266 25617 5266 6 n_148
rlabel m2contact 25617 5242 25617 5242 6 n_398
rlabel m2contact 25593 7162 25593 7162 6 n_146
rlabel m2contact 25569 5050 25569 5050 6 n_171
rlabel m2contact 25545 2818 25545 2818 6 n_147
rlabel m2contact 25521 5698 25521 5698 6 n_170
rlabel m2contact 25497 5506 25497 5506 6 n_155
rlabel m2contact 25497 4642 25497 4642 6 n_155
rlabel m2contact 25473 4618 25473 4618 6 Op2Sel[1]
rlabel m2contact 25449 6730 25449 6730 6 n_45
rlabel m2contact 25449 4666 25449 4666 6 n_45
rlabel m2contact 25425 3994 25425 3994 6 nOE
rlabel m2contact 25401 6778 25401 6778 6 n_64
rlabel m2contact 25377 4594 25377 4594 6 stateSub[1]
rlabel m2contact 25377 5074 25377 5074 6 n_251
rlabel m2contact 25353 6202 25353 6202 6 n_310
rlabel m2contact 25353 6178 25353 6178 6 n_116
rlabel m2contact 25329 4762 25329 4762 6 n_29
rlabel m2contact 25329 2650 25329 2650 6 n_29
rlabel m2contact 25305 5506 25305 5506 6 n_155
rlabel m2contact 25305 5482 25305 5482 6 n_28
rlabel m2contact 25281 4906 25281 4906 6 n_154
rlabel m2contact 25281 4786 25281 4786 6 n_225
rlabel m2contact 25257 4138 25257 4138 6 n_157
rlabel m2contact 25257 3442 25257 3442 6 n_119
rlabel m2contact 25233 4714 25233 4714 6 n_79
rlabel m2contact 25233 2722 25233 2722 6 n_79
rlabel m2contact 25209 4666 25209 4666 6 n_45
rlabel m2contact 25209 6370 25209 6370 6 n_55
rlabel m2contact 25185 2938 25185 2938 6 n_44
rlabel m2contact 25185 2986 25185 2986 6 n_392
rlabel m2contact 25161 3154 25161 3154 6 n_110
rlabel m2contact 25137 4666 25137 4666 6 OpcodeCondIn[3]
rlabel m2contact 25137 3418 25137 3418 6 OpcodeCondIn[3]
rlabel m2contact 25113 6778 25113 6778 6 n_64
rlabel m2contact 25113 6754 25113 6754 6 n_242
rlabel m2contact 25089 4762 25089 4762 6 n_29
rlabel m2contact 25089 4354 25089 4354 6 stateSub[0]
rlabel m2contact 25065 4714 25065 4714 6 n_79
rlabel m2contact 25065 3562 25065 3562 6 n_241
rlabel m2contact 25041 6778 25041 6778 6 n_90
rlabel m2contact 25041 2842 25041 2842 6 n_90
rlabel m2contact 25017 4618 25017 4618 6 Op2Sel[1]
rlabel m2contact 25017 4762 25017 4762 6 n_174
rlabel m2contact 24993 4666 24993 4666 6 OpcodeCondIn[3]
rlabel m2contact 24993 3466 24993 3466 6 n_353
rlabel m2contact 24969 6778 24969 6778 6 n_90
rlabel m2contact 24969 6706 24969 6706 6 n_332
rlabel m2contact 24945 2242 24945 2242 6 n_364
rlabel m2contact 24945 5194 24945 5194 6 n_166
rlabel m2contact 24921 2890 24921 2890 6 n_92
rlabel m2contact 24873 6130 24873 6130 6 n_363
rlabel m2contact 24873 2194 24873 2194 6 n_363
rlabel m2contact 24849 5170 24849 5170 6 n_359
rlabel m2contact 24825 4594 24825 4594 6 n_369
rlabel m2contact 24801 6130 24801 6130 6 n_363
rlabel m2contact 24801 6082 24801 6082 6 stateSub[1]
rlabel m2contact 24753 3442 24753 3442 6 n_119
rlabel m2contact 24729 5626 24729 5626 6 n_13
rlabel m2contact 24633 3682 24633 3682 6 OpcodeCondIn[1]
rlabel m2contact 24609 4186 24609 4186 6 OpcodeCondIn[0]
rlabel m2contact 24561 2266 24561 2266 6 n_117
rlabel m2contact 24537 3442 24537 3442 6 n_119
rlabel m2contact 24513 6178 24513 6178 6 n_116
rlabel m2contact 24465 5506 24465 5506 6 n_308
rlabel m2contact 24417 1858 24417 1858 6 n_82
rlabel m2contact 24393 3754 24393 3754 6 n_273
rlabel m2contact 24357 6442 24357 6442 6 n_262
rlabel m2contact 24357 4618 24357 4618 6 n_262
rlabel m2contact 24333 5866 24333 5866 6 n_50
rlabel m2contact 24333 4666 24333 4666 6 n_50
rlabel m2contact 24321 7402 24321 7402 6 n_305
rlabel m2contact 24297 2194 24297 2194 6 n_363
rlabel m2contact 24273 4618 24273 4618 6 n_262
rlabel m2contact 24273 5170 24273 5170 6 n_359
rlabel m2contact 24249 3850 24249 3850 6 n_261
rlabel m2contact 24225 5866 24225 5866 6 n_50
rlabel m2contact 24225 5842 24225 5842 6 n_219
rlabel m2contact 24201 4954 24201 4954 6 n_14
rlabel m2contact 24177 5002 24177 5002 6 n_87
rlabel m2contact 24177 5554 24177 5554 6 n_137
rlabel m2contact 24153 7042 24153 7042 6 n_53
rlabel m2contact 24153 2554 24153 2554 6 n_53
rlabel m2contact 24129 2554 24129 2554 6 n_53
rlabel m2contact 24129 2578 24129 2578 6 n_36
rlabel m2contact 24105 5146 24105 5146 6 n_350
rlabel m2contact 24105 3490 24105 3490 6 n_350
rlabel m2contact 24105 2674 24105 2674 6 n_314
rlabel m2contact 24105 2074 24105 2074 6 n_314
rlabel m2contact 24081 3490 24081 3490 6 n_350
rlabel m2contact 24081 3514 24081 3514 6 OpcodeCondIn[6]
rlabel m2contact 24057 7162 24057 7162 6 n_146
rlabel m2contact 24057 3610 24057 3610 6 n_81
rlabel m2contact 24033 7306 24033 7306 6 n_304
rlabel m2contact 24009 4618 24009 4618 6 n_164
rlabel m2contact 23985 2074 23985 2074 6 n_314
rlabel m2contact 23985 2098 23985 2098 6 IRQ2
rlabel m2contact 23961 4882 23961 4882 6 n_93
rlabel m2contact 23937 2146 23937 2146 6 IntStatus
rlabel m2contact 23889 5026 23889 5026 6 n_212
rlabel m2contact 23865 6490 23865 6490 6 n_140
rlabel m2contact 23841 6850 23841 6850 6 n_153
rlabel m2contact 23841 4714 23841 4714 6 state[0]
rlabel m2contact 23793 3010 23793 3010 6 n_255
rlabel m2contact 23793 2938 23793 2938 6 n_44
rlabel m2contact 23769 4930 23769 4930 6 n_228
rlabel m2contact 23745 6610 23745 6610 6 n_253
rlabel m2contact 23673 4738 23673 4738 6 n_302
rlabel m2contact 23649 6994 23649 6994 6 n_329
rlabel m2contact 23649 2794 23649 2794 6 n_329
rlabel m2contact 23625 2770 23625 2770 6 n_284
rlabel m2contact 23589 6106 23589 6106 6 n_346
rlabel m2contact 23589 3634 23589 3634 6 n_346
rlabel m2contact 23577 7354 23577 7354 6 n_179
rlabel m2contact 23553 6922 23553 6922 6 n_263
rlabel m2contact 23553 4570 23553 4570 6 n_263
rlabel m2contact 23529 4714 23529 4714 6 state[0]
rlabel m2contact 23505 5530 23505 5530 6 n_232
rlabel m2contact 23481 6202 23481 6202 6 n_233
rlabel m2contact 23481 3394 23481 3394 6 n_233
rlabel m2contact 23457 5290 23457 5290 6 n_276
rlabel m2contact 23433 2338 23433 2338 6 n_274
rlabel m2contact 23409 5674 23409 5674 6 n_214
rlabel m2contact 23385 3154 23385 3154 6 n_110
rlabel m2contact 23361 6298 23361 6298 6 n_275
rlabel m2contact 23325 4738 23325 4738 6 OpcodeCondIn[4]
rlabel m2contact 23325 3226 23325 3226 6 OpcodeCondIn[4]
rlabel m2contact 23313 5362 23313 5362 6 n_11
rlabel m2contact 23289 4738 23289 4738 6 OpcodeCondIn[4]
rlabel m2contact 23289 4474 23289 4474 6 n_252
rlabel m2contact 23265 3034 23265 3034 6 n_127
rlabel m2contact 23265 4786 23265 4786 6 n_225
rlabel m2contact 23241 5842 23241 5842 6 n_219
rlabel m2contact 23241 3658 23241 3658 6 n_219
rlabel m2contact 23217 3178 23217 3178 6 AluOR[1]
rlabel m2contact 23217 3202 23217 3202 6 Op1Sel
rlabel m2contact 23193 3466 23193 3466 6 n_353
rlabel m2contact 23169 2794 23169 2794 6 n_329
rlabel m2contact 23169 2914 23169 2914 6 n_234
rlabel m2contact 23145 4234 23145 4234 6 n_288
rlabel m2contact 23109 5338 23109 5338 6 AluOR[0]
rlabel m2contact 23109 4450 23109 4450 6 AluOR[0]
rlabel m2contact 23097 5650 23097 5650 6 n_113
rlabel m2contact 23097 3898 23097 3898 6 n_99
rlabel m2contact 23073 4282 23073 4282 6 n_33
rlabel m2contact 23073 4930 23073 4930 6 n_228
rlabel m2contact 23049 4738 23049 4738 6 n_112
rlabel m2contact 23049 2626 23049 2626 6 n_98
rlabel m2contact 23025 6346 23025 6346 6 n_108
rlabel m2contact 23025 2482 23025 2482 6 n_108
rlabel m2contact 23001 5314 23001 5314 6 SysBus[3]
rlabel m2contact 23001 7042 23001 7042 6 n_53
rlabel m2contact 22977 6082 22977 6082 6 stateSub[1]
rlabel m2contact 22953 3634 22953 3634 6 n_346
rlabel m2contact 22953 3706 22953 3706 6 state[1]
rlabel m2contact 22929 7258 22929 7258 6 n_118
rlabel m2contact 22905 6682 22905 6682 6 n_35
rlabel m2contact 22881 4570 22881 4570 6 n_263
rlabel m2contact 22881 4714 22881 4714 6 state[0]
rlabel m2contact 22857 6826 22857 6826 6 n_78
rlabel m2contact 22857 6058 22857 6058 6 n_185
rlabel m2contact 22833 5266 22833 5266 6 n_234
rlabel m2contact 22833 2914 22833 2914 6 n_234
rlabel m2contact 22809 2194 22809 2194 6 n_363
rlabel m2contact 22785 5698 22785 5698 6 n_170
rlabel m2contact 22761 3394 22761 3394 6 n_233
rlabel m2contact 22761 3466 22761 3466 6 n_353
rlabel m2contact 22737 6586 22737 6586 6 n_254
rlabel m2contact 22713 4402 22713 4402 6 n_61
rlabel m2contact 22689 5338 22689 5338 6 AluOR[0]
rlabel m2contact 22689 5218 22689 5218 6 n_162
rlabel m2contact 22665 4570 22665 4570 6 n_223
rlabel m2contact 22641 6298 22641 6298 6 n_275
rlabel m2contact 22617 3658 22617 3658 6 n_219
rlabel m2contact 22617 3706 22617 3706 6 state[1]
rlabel m2contact 22593 4714 22593 4714 6 state[0]
rlabel m2contact 22569 4618 22569 4618 6 n_164
rlabel m2contact 22545 6538 22545 6538 6 n_239
rlabel m2contact 22545 4522 22545 4522 6 n_239
rlabel m2contact 22521 7186 22521 7186 6 n_303
rlabel m2contact 22521 4546 22521 4546 6 n_290
rlabel m2contact 22497 5746 22497 5746 6 n_128
rlabel m2contact 22497 4090 22497 4090 6 n_128
rlabel m2contact 22473 3802 22473 3802 6 n_285
rlabel m2contact 22473 3514 22473 3514 6 OpcodeCondIn[6]
rlabel m2contact 22449 3754 22449 3754 6 n_273
rlabel m2contact 22425 6274 22425 6274 6 n_181
rlabel m2contact 22401 7354 22401 7354 6 n_179
rlabel m2contact 22377 2482 22377 2482 6 n_108
rlabel m2contact 22377 2506 22377 2506 6 n_180
rlabel m2contact 22353 3730 22353 3730 6 n_135
rlabel m2contact 22329 5434 22329 5434 6 n_229
rlabel m2contact 22305 4930 22305 4930 6 n_228
rlabel m2contact 22281 6202 22281 6202 6 n_233
rlabel m2contact 22281 3418 22281 3418 6 OpcodeCondIn[3]
rlabel m2contact 22257 5266 22257 5266 6 n_234
rlabel m2contact 22257 5194 22257 5194 6 n_166
rlabel m2contact 22221 6946 22221 6946 6 StatusRegEn
rlabel m2contact 22221 4618 22221 4618 6 StatusRegEn
rlabel m2contact 22209 3274 22209 3274 6 n_158
rlabel m2contact 22185 2530 22185 2530 6 n_312
rlabel m2contact 22161 4138 22161 4138 6 n_157
rlabel m2contact 22137 7114 22137 7114 6 n_298
rlabel m2contact 22113 3754 22113 3754 6 n_273
rlabel m2contact 22089 4498 22089 4498 6 OpcodeCondIn[7]
rlabel m2contact 22065 4522 22065 4522 6 n_239
rlabel m2contact 22065 5698 22065 5698 6 n_170
rlabel m2contact 22041 6130 22041 6130 6 n_79
rlabel m2contact 22041 2722 22041 2722 6 n_79
rlabel m2contact 22017 4450 22017 4450 6 AluOR[0]
rlabel m2contact 22017 4498 22017 4498 6 OpcodeCondIn[7]
rlabel m2contact 21993 3466 21993 3466 6 n_353
rlabel m2contact 21969 6994 21969 6994 6 n_329
rlabel m2contact 21945 7162 21945 7162 6 n_146
rlabel m2contact 21921 4258 21921 4258 6 n_151
rlabel m2contact 21897 4090 21897 4090 6 n_128
rlabel m2contact 21897 4114 21897 4114 6 OpcodeCondIn[2]
rlabel m2contact 21873 4138 21873 4138 6 n_157
rlabel m2contact 21849 2554 21849 2554 6 n_247
rlabel m2contact 21825 4978 21825 4978 6 n_182
rlabel m2contact 21801 6202 21801 6202 6 n_233
rlabel m2contact 21801 3418 21801 3418 6 OpcodeCondIn[3]
rlabel m2contact 21777 4474 21777 4474 6 n_252
rlabel m2contact 21753 7066 21753 7066 6 n_203
rlabel m2contact 21753 4450 21753 4450 6 n_203
rlabel m2contact 21729 6946 21729 6946 6 StatusRegEn
rlabel m2contact 21729 6898 21729 6898 6 n_348
rlabel m2contact 21705 3178 21705 3178 6 StatusReg[0]
rlabel m2contact 21681 6130 21681 6130 6 n_79
rlabel m2contact 21681 6106 21681 6106 6 n_346
rlabel m2contact 21657 5578 21657 5578 6 ENB
rlabel m2contact 21657 4306 21657 4306 6 ENB
rlabel m2contact 21633 2938 21633 2938 6 n_44
rlabel m2contact 21609 5554 21609 5554 6 n_137
rlabel m2contact 21609 3922 21609 3922 6 n_195
rlabel m2contact 21585 2722 21585 2722 6 n_79
rlabel m2contact 21561 6418 21561 6418 6 n_134
rlabel m2contact 21537 4450 21537 4450 6 n_203
rlabel m2contact 21537 4498 21537 4498 6 OpcodeCondIn[7]
rlabel m2contact 21513 5386 21513 5386 6 n_89
rlabel m2contact 21513 4018 21513 4018 6 nWait
rlabel m2contact 21489 4090 21489 4090 6 n_202
rlabel m2contact 21465 5578 21465 5578 6 ENB
rlabel m2contact 21465 5554 21465 5554 6 n_137
rlabel m2contact 21393 4042 21393 4042 6 n_230
rlabel m2contact 21345 6514 21345 6514 6 n_236
rlabel m2contact 21321 3178 21321 3178 6 StatusReg[0]
rlabel m2contact 21297 5098 21297 5098 6 n_96
rlabel m2contact 21273 6322 21273 6322 6 n_393
rlabel m2contact 21273 6226 21273 6226 6 n_10
rlabel m2contact 21249 5578 21249 5578 6 n_19
rlabel m2contact 21201 3058 21201 3058 6 n_280
rlabel m2contact 21177 7162 21177 7162 6 n_146
rlabel m2contact 21129 4090 21129 4090 6 n_202
rlabel m2contact 21105 5266 21105 5266 6 n_83
rlabel m2contact 21105 3490 21105 3490 6 n_83
rlabel m2contact 21081 4306 21081 4306 6 ENB
rlabel m2contact 21081 2482 21081 2482 6 ENB
rlabel m2contact 21057 4618 21057 4618 6 StatusRegEn
rlabel m2contact 21033 6322 21033 6322 6 n_44
rlabel m2contact 21033 2938 21033 2938 6 n_44
rlabel m2contact 21009 5890 21009 5890 6 n_74
rlabel m2contact 21009 1930 21009 1930 6 n_74
rlabel m2contact 20985 4858 20985 4858 6 n_168
rlabel m2contact 20985 2122 20985 2122 6 n_168
rlabel m2contact 20961 5338 20961 5338 6 n_318
rlabel m2contact 20937 3442 20937 3442 6 n_119
rlabel m2contact 20913 5722 20913 5722 6 n_372
rlabel m2contact 20913 2722 20913 2722 6 n_79
rlabel m2contact 20889 3706 20889 3706 6 state[1]
rlabel m2contact 20865 7330 20865 7330 6 n_129
rlabel m2contact 20865 3586 20865 3586 6 n_129
rlabel m2contact 20841 4834 20841 4834 6 n_222
rlabel m2contact 20841 3130 20841 3130 6 n_222
rlabel m2contact 20829 6130 20829 6130 6 n_137
rlabel m2contact 20829 5554 20829 5554 6 n_137
rlabel m2contact 20817 4474 20817 4474 6 n_252
rlabel m2contact 20793 5602 20793 5602 6 n_165
rlabel m2contact 20793 5554 20793 5554 6 n_137
rlabel m2contact 20769 5266 20769 5266 6 n_83
rlabel m2contact 20769 4426 20769 4426 6 n_183
rlabel m2contact 20745 6010 20745 6010 6 stateSub[2]
rlabel m2contact 20721 2482 20721 2482 6 ENB
rlabel m2contact 20721 2602 20721 2602 6 n_120
rlabel m2contact 20697 6154 20697 6154 6 n_84
rlabel m2contact 20673 5770 20673 5770 6 n_218
rlabel m2contact 20649 6874 20649 6874 6 n_159
rlabel m2contact 20625 3634 20625 3634 6 n_217
rlabel m2contact 20601 4714 20601 4714 6 state[0]
rlabel m2contact 20577 2338 20577 2338 6 n_274
rlabel m2contact 20553 4786 20553 4786 6 n_225
rlabel m2contact 20529 6322 20529 6322 6 n_44
rlabel m2contact 20529 6154 20529 6154 6 n_84
rlabel m2contact 20505 4354 20505 4354 6 stateSub[0]
rlabel m2contact 20481 5866 20481 5866 6 n_115
rlabel m2contact 20481 2722 20481 2722 6 n_79
rlabel m2contact 20457 5890 20457 5890 6 n_74
rlabel m2contact 20457 5818 20457 5818 6 n_286
rlabel m2contact 20433 2410 20433 2410 6 n_66
rlabel m2contact 20409 5266 20409 5266 6 n_150
rlabel m2contact 20385 2026 20385 2026 6 n_149
rlabel m2contact 20385 7282 20385 7282 6 n_138
rlabel m2contact 20361 6130 20361 6130 6 n_137
rlabel m2contact 20361 6058 20361 6058 6 n_185
rlabel m2contact 20337 5002 20337 5002 6 n_87
rlabel m2contact 20337 4066 20337 4066 6 n_192
rlabel m2contact 20313 6634 20313 6634 6 n_315
rlabel m2contact 20313 5914 20313 5914 6 n_315
rlabel m2contact 20313 5458 20313 5458 6 n_27
rlabel m2contact 20313 2482 20313 2482 6 n_27
rlabel m2contact 20289 2698 20289 2698 6 Op2Sel[0]
rlabel m2contact 20265 3226 20265 3226 6 OpcodeCondIn[4]
rlabel m2contact 20241 4858 20241 4858 6 n_168
rlabel m2contact 20241 2794 20241 2794 6 n_191
rlabel m2contact 20217 5938 20217 5938 6 n_206
rlabel m2contact 20217 3970 20217 3970 6 n_206
rlabel m2contact 20193 2698 20193 2698 6 Op2Sel[0]
rlabel m2contact 20193 3082 20193 3082 6 n_51
rlabel m2contact 20169 7330 20169 7330 6 n_129
rlabel m2contact 20169 7234 20169 7234 6 n_211
rlabel m2contact 20145 5410 20145 5410 6 n_351
rlabel m2contact 20121 6634 20121 6634 6 n_315
rlabel m2contact 20121 6562 20121 6562 6 n_209
rlabel m2contact 20097 6034 20097 6034 6 n_20
rlabel m2contact 20073 6442 20073 6442 6 n_262
rlabel m2contact 20073 6322 20073 6322 6 n_136
rlabel m2contact 20049 4834 20049 4834 6 n_222
rlabel m2contact 20049 3778 20049 3778 6 n_69
rlabel m2contact 20025 2674 20025 2674 6 n_314
rlabel m2contact 19989 5002 19989 5002 6 n_59
rlabel m2contact 19989 2698 19989 2698 6 n_59
rlabel m2contact 19977 7258 19977 7258 6 n_118
rlabel m2contact 19953 4426 19953 4426 6 n_183
rlabel m2contact 19929 2722 19929 2722 6 n_79
rlabel m2contact 19929 5698 19929 5698 6 n_170
rlabel m2contact 19905 7450 19905 7450 6 n_100
rlabel m2contact 19905 4378 19905 4378 6 n_100
rlabel m2contact 19881 4330 19881 4330 6 n_122
rlabel m2contact 19857 5458 19857 5458 6 n_27
rlabel m2contact 19857 4930 19857 4930 6 n_228
rlabel m2contact 19833 4858 19833 4858 6 n_121
rlabel m2contact 19809 4522 19809 4522 6 n_67
rlabel m2contact 19785 3874 19785 3874 6 n_188
rlabel m2contact 19761 3970 19761 3970 6 n_206
rlabel m2contact 19761 4114 19761 4114 6 OpcodeCondIn[2]
rlabel m2contact 19737 2698 19737 2698 6 n_59
rlabel m2contact 19737 2818 19737 2818 6 n_147
rlabel m2contact 19713 4978 19713 4978 6 n_182
rlabel m2contact 19713 4618 19713 4618 6 n_207
rlabel m2contact 19689 5554 19689 5554 6 n_137
rlabel m2contact 19689 3658 19689 3658 6 n_137
rlabel m2contact 19665 3826 19665 3826 6 n_125
rlabel m2contact 19641 4666 19641 4666 6 n_50
rlabel m2contact 19617 4450 19617 4450 6 n_8
rlabel m2contact 19593 5890 19593 5890 6 n_395
rlabel m2contact 19569 4834 19569 4834 6 n_63
rlabel m2contact 19545 4378 19545 4378 6 n_100
rlabel m2contact 19545 4498 19545 4498 6 OpcodeCondIn[7]
rlabel m2contact 19521 3346 19521 3346 6 n_31
rlabel m2contact 19497 4402 19497 4402 6 n_61
rlabel m2contact 19473 3658 19473 3658 6 n_137
rlabel m2contact 19473 3970 19473 3970 6 n_221
rlabel m2contact 19449 2458 19449 2458 6 n_70
rlabel m2contact 19425 4378 19425 4378 6 n_163
rlabel m2contact 19401 2698 19401 2698 6 n_40
rlabel m2contact 19377 3658 19377 3658 6 n_97
rlabel m2contact 19353 3754 19353 3754 6 n_273
rlabel m2contact 19353 4666 19353 4666 6 n_194
rlabel m2contact 19329 5458 19329 5458 6 MemEn
rlabel m2contact 19329 4162 19329 4162 6 MemEn
rlabel m2contact 19305 2434 19305 2434 6 n_131
rlabel m2contact 19281 3874 19281 3874 6 n_188
rlabel m2contact 19281 3370 19281 3370 6 OpcodeCondIn[5]
rlabel m2contact 19257 4138 19257 4138 6 n_157
rlabel m2contact 19233 5986 19233 5986 6 n_277
rlabel m2contact 19209 3586 19209 3586 6 n_129
rlabel m2contact 19209 3850 19209 3850 6 n_261
rlabel m2contact 19185 6778 19185 6778 6 n_282
rlabel m2contact 19161 5746 19161 5746 6 n_128
rlabel m2contact 19137 5458 19137 5458 6 MemEn
rlabel m2contact 19137 4690 19137 4690 6 n_94
rlabel m2contact 19089 6130 19089 6130 6 n_367
rlabel m2contact 19089 3586 19089 3586 6 n_272
rlabel m2contact 19065 5458 19065 5458 6 n_32
rlabel m2contact 19065 2314 19065 2314 6 n_32
rlabel m2contact 19041 5458 19041 5458 6 n_32
rlabel m2contact 19041 3250 19041 3250 6 n_72
rlabel m2contact 19017 3754 19017 3754 6 n_273
rlabel m2contact 19017 5146 19017 5146 6 n_350
rlabel m2contact 18993 7042 18993 7042 6 n_53
rlabel m2contact 18993 2362 18993 2362 6 n_53
rlabel m2contact 18969 5602 18969 5602 6 n_309
rlabel m2contact 18969 3754 18969 3754 6 n_309
rlabel m2contact 18945 2362 18945 2362 6 n_53
rlabel m2contact 18945 3298 18945 3298 6 n_338
rlabel m2contact 18921 5602 18921 5602 6 n_309
rlabel m2contact 18921 5482 18921 5482 6 n_28
rlabel m2contact 18897 6514 18897 6514 6 n_236
rlabel m2contact 18897 3394 18897 3394 6 n_236
rlabel m2contact 18873 3082 18873 3082 6 n_51
rlabel m2contact 18849 3394 18849 3394 6 n_236
rlabel m2contact 18849 6082 18849 6082 6 stateSub[1]
rlabel m2contact 18825 3562 18825 3562 6 n_241
rlabel m2contact 18825 3922 18825 3922 6 n_195
rlabel m2contact 18777 6610 18777 6610 6 n_253
rlabel m2contact 18753 4162 18753 4162 6 MemEn
rlabel m2contact 18729 5458 18729 5458 6 n_210
rlabel m2contact 18705 4306 18705 4306 6 ENB
rlabel m2contact 18705 6202 18705 6202 6 n_233
rlabel m2contact 18633 6346 18633 6346 6 n_108
rlabel m2contact 18633 6178 18633 6178 6 n_116
rlabel m2contact 18585 5146 18585 5146 6 n_123
rlabel m2contact 18513 5794 18513 5794 6 n_334
rlabel m2contact 18489 2194 18489 2194 6 n_363
rlabel m2contact 18465 5602 18465 5602 6 n_270
rlabel m2contact 18417 3634 18417 3634 6 n_217
rlabel m2contact 18393 4978 18393 4978 6 n_182
rlabel m2contact 18369 2506 18369 2506 6 n_180
rlabel m2contact 18321 4306 18321 4306 6 n_292
rlabel m2contact 18297 5314 18297 5314 6 SysBus[3]
rlabel m2contact 18273 3394 18273 3394 6 n_294
rlabel m2contact 18225 6634 18225 6634 6 n_231
rlabel m2contact 18201 4042 18201 4042 6 n_230
rlabel m2contact 18177 6538 18177 6538 6 n_239
rlabel m2contact 18129 5314 18129 5314 6 n_47
rlabel m2contact 18081 4114 18081 4114 6 OpcodeCondIn[2]
rlabel m2contact 18057 4210 18057 4210 6 n_46
rlabel m2contact 18009 2434 18009 2434 6 n_131
rlabel m2contact 17985 4354 17985 4354 6 stateSub[0]
rlabel m2contact 17961 6058 17961 6058 6 n_185
rlabel m2contact 17937 5962 17937 5962 6 n_71
rlabel m2contact 17937 1906 17937 1906 6 n_71
rlabel m2contact 17913 5962 17913 5962 6 n_71
rlabel m2contact 17913 5050 17913 5050 6 n_171
rlabel m2contact 17889 4426 17889 4426 6 n_183
rlabel m2contact 17865 4162 17865 4162 6 n_9
rlabel m2contact 17865 3706 17865 3706 6 state[1]
rlabel m2contact 17841 2938 17841 2938 6 n_44
rlabel m2contact 17793 2458 17793 2458 6 n_70
rlabel m2contact 17769 5554 17769 5554 6 n_137
rlabel m2contact 17745 5530 17745 5530 6 n_232
rlabel m2contact 17721 2074 17721 2074 6 CFlag
rlabel m2contact 17697 5170 17697 5170 6 n_359
rlabel m2contact 17625 2554 17625 2554 6 n_247
rlabel m2contact 17577 2842 17577 2842 6 n_90
rlabel m2contact 17529 6010 17529 6010 6 stateSub[2]
rlabel m2contact 17481 5962 17481 5962 6 n_293
rlabel m2contact 17433 3394 17433 3394 6 n_294
rlabel m2contact 17385 6226 17385 6226 6 n_10
rlabel m2contact 17361 3418 17361 3418 6 OpcodeCondIn[3]
rlabel m2contact 17337 3514 17337 3514 6 OpcodeCondIn[6]
rlabel m2contact 17313 7498 17313 7498 6 n_370
rlabel m2contact 17265 4234 17265 4234 6 n_288
rlabel m2contact 17217 5506 17217 5506 6 n_308
rlabel m2contact 17193 4618 17193 4618 6 n_207
rlabel m2contact 17145 5218 17145 5218 6 n_162
rlabel m2contact 17121 4138 17121 4138 6 n_157
rlabel m2contact 17097 4018 17097 4018 6 nWait
rlabel m2contact 17073 6346 17073 6346 6 n_77
rlabel m2contact 17073 2554 17073 2554 6 n_77
rlabel m2contact 17049 2026 17049 2026 6 n_149
rlabel m2contact 17025 3418 17025 3418 6 OpcodeCondIn[3]
rlabel m2contact 17001 6346 17001 6346 6 n_77
rlabel m2contact 17001 4234 17001 4234 6 n_268
rlabel m2contact 16953 2458 16953 2458 6 WdSel
rlabel m2contact 16929 4354 16929 4354 6 stateSub[0]
rlabel m2contact 16905 3874 16905 3874 6 n_188
rlabel m2contact 16905 4882 16905 4882 6 n_93
rlabel m2contact 16881 2890 16881 2890 6 n_92
rlabel m2contact 16857 7450 16857 7450 6 n_100
rlabel m2contact 16833 6346 16833 6346 6 n_142
rlabel m2contact 16833 2842 16833 2842 6 n_142
rlabel m2contact 16809 2842 16809 2842 6 n_142
rlabel m2contact 16809 3874 16809 3874 6 n_176
rlabel m2contact 16785 2746 16785 2746 6 n_49
rlabel m2contact 16785 3226 16785 3226 6 OpcodeCondIn[4]
rlabel m2contact 16761 2842 16761 2842 6 n_80
rlabel m2contact 16761 3730 16761 3730 6 n_135
rlabel m2contact 16737 6442 16737 6442 6 n_227
rlabel m2contact 16737 2362 16737 2362 6 n_227
rlabel m2contact 16713 2890 16713 2890 6 n_92
rlabel m2contact 16713 4882 16713 4882 6 n_301
rlabel m2contact 16689 6466 16689 6466 6 n_22
rlabel m2contact 16689 4498 16689 4498 6 OpcodeCondIn[7]
rlabel m2contact 16665 6442 16665 6442 6 n_227
rlabel m2contact 16665 2794 16665 2794 6 n_191
rlabel m2contact 16641 2746 16641 2746 6 n_86
rlabel m2contact 16617 7378 16617 7378 6 n_278
rlabel m2contact 16593 2914 16593 2914 6 n_234
rlabel m2contact 16569 2386 16569 2386 6 n_148
rlabel m2contact 16545 7162 16545 7162 6 n_146
rlabel m2contact 16521 2458 16521 2458 6 WdSel
rlabel m2contact 16521 5626 16521 5626 6 n_13
rlabel m2contact 16473 6802 16473 6802 6 n_279
rlabel m2contact 16473 5626 16473 5626 6 n_7
rlabel m2contact 16449 2386 16449 2386 6 n_48
rlabel m2contact 16449 2002 16449 2002 6 n_193
rlabel m2contact 16425 6418 16425 6418 6 n_134
rlabel m2contact 16401 1882 16401 1882 6 n_114
rlabel m2contact 16377 1954 16377 1954 6 n_199
rlabel m2contact 16329 6946 16329 6946 6 n_109
rlabel m2contact 16305 2098 16305 2098 6 IRQ2
rlabel m2contact 16305 5818 16305 5818 6 n_286
rlabel m2contact 16281 6178 16281 6178 6 n_116
rlabel m2contact 16233 2458 16233 2458 6 PcWe
rlabel m2contact 16185 6394 16185 6394 6 Rs1Sel[0]
rlabel m2contact 16161 6298 16161 6298 6 n_275
rlabel m2contact 16137 6130 16137 6130 6 n_367
rlabel m2contact 16089 5674 16089 5674 6 n_214
rlabel m2contact 16041 5674 16041 5674 6 n_160
rlabel m2contact 16017 6466 16017 6466 6 n_213
rlabel m2contact 15945 3250 15945 3250 6 n_72
rlabel m2contact 15897 3418 15897 3418 6 OpcodeCondIn[3]
rlabel m2contact 15849 5410 15849 5410 6 n_351
rlabel m2contact 15825 3226 15825 3226 6 OpcodeCondIn[4]
rlabel m2contact 15801 6658 15801 6658 6 n_331
rlabel m2contact 15777 2506 15777 2506 6 n_180
rlabel m2contact 15753 4138 15753 4138 6 n_157
rlabel m2contact 15729 4498 15729 4498 6 OpcodeCondIn[7]
rlabel m2contact 15705 3154 15705 3154 6 n_110
rlabel m2contact 15705 2818 15705 2818 6 n_147
rlabel m2contact 15681 6058 15681 6058 6 n_185
rlabel m2contact 15657 4162 15657 4162 6 n_9
rlabel m2contact 15633 6418 15633 6418 6 n_37
rlabel m2contact 15633 3250 15633 3250 6 n_72
rlabel m2contact 15609 3922 15609 3922 6 n_195
rlabel m2contact 15585 4186 15585 4186 6 OpcodeCondIn[0]
rlabel m2contact 15561 2386 15561 2386 6 n_48
rlabel m2contact 15561 4162 15561 4162 6 n_17
rlabel m2contact 15537 3370 15537 3370 6 OpcodeCondIn[5]
rlabel m2contact 15513 4786 15513 4786 6 n_225
rlabel m2contact 15489 2890 15489 2890 6 n_92
rlabel m2contact 15441 5410 15441 5410 6 n_6
rlabel m2contact 15417 6010 15417 6010 6 stateSub[2]
rlabel m2contact 15417 3682 15417 3682 6 OpcodeCondIn[1]
rlabel m2contact 15393 4186 15393 4186 6 OpcodeCondIn[0]
rlabel m2contact 15369 5554 15369 5554 6 n_137
rlabel m2contact 15321 3514 15321 3514 6 OpcodeCondIn[6]
rlabel m2contact 15297 2290 15297 2290 6 n_18
rlabel m2contact 15249 2458 15249 2458 6 PcWe
rlabel m2contact 15201 2530 15201 2530 6 n_312
rlabel m2contact 15153 2674 15153 2674 6 n_314
rlabel m2contact 15129 6010 15129 6010 6 stateSub[2]
rlabel m2contact 15105 3082 15105 3082 6 n_51
rlabel m2contact 15033 7138 15033 7138 6 n_300
rlabel m2contact 15009 5914 15009 5914 6 n_315
rlabel m2contact 14949 5914 14949 5914 6 n_338
rlabel m2contact 14949 3298 14949 3298 6 n_338
rlabel m2contact 14949 7090 14949 7090 6 n_116
rlabel m2contact 14949 6178 14949 6178 6 n_116
rlabel m2contact 14937 2530 14937 2530 6 n_12
rlabel m2contact 14913 3418 14913 3418 6 OpcodeCondIn[3]
rlabel m2contact 14889 5914 14889 5914 6 n_338
rlabel m2contact 14889 4498 14889 4498 6 OpcodeCondIn[7]
rlabel m2contact 14865 6826 14865 6826 6 n_78
rlabel m2contact 14841 7090 14841 7090 6 n_116
rlabel m2contact 14841 7018 14841 7018 6 n_30
rlabel m2contact 14817 3226 14817 3226 6 OpcodeCondIn[4]
rlabel m2contact 14793 5698 14793 5698 6 n_170
rlabel m2contact 14745 4594 14745 4594 6 n_369
rlabel m2contact 14697 3202 14697 3202 6 Op1Sel
rlabel m2contact 14673 4594 14673 4594 6 n_361
rlabel m2contact 14649 7426 14649 7426 6 n_394
rlabel m2contact 14625 6970 14625 6970 6 n_238
rlabel m2contact 14601 2458 14601 2458 6 n_42
rlabel m2contact 14577 6538 14577 6538 6 n_239
rlabel m2contact 14553 7330 14553 7330 6 n_244
rlabel m2contact 14553 2386 14553 2386 6 n_244
rlabel m2contact 14529 3754 14529 3754 6 n_309
rlabel m2contact 14505 5506 14505 5506 6 n_308
rlabel m2contact 14481 6826 14481 6826 6 n_78
rlabel m2contact 14481 2050 14481 2050 6 n_78
rlabel m2contact 14457 7474 14457 7474 6 n_324
rlabel m2contact 14457 3082 14457 3082 6 n_324
rlabel m2contact 14433 5122 14433 5122 6 n_310
rlabel m2contact 14409 5530 14409 5530 6 n_232
rlabel m2contact 14385 2386 14385 2386 6 n_244
rlabel m2contact 14349 5530 14349 5530 6 n_232
rlabel m2contact 14349 3754 14349 3754 6 n_232
rlabel m2contact 14337 3394 14337 3394 6 n_294
rlabel m2contact 14313 6082 14313 6082 6 stateSub[1]
rlabel m2contact 14313 2674 14313 2674 6 stateSub[1]
rlabel m2contact 14289 6130 14289 6130 6 n_362
rlabel m2contact 14289 4498 14289 4498 6 OpcodeCondIn[7]
rlabel m2contact 14265 4666 14265 4666 6 n_194
rlabel m2contact 14241 6394 14241 6394 6 n_147
rlabel m2contact 14241 2818 14241 2818 6 n_147
rlabel m2contact 14217 4666 14217 4666 6 state[1]
rlabel m2contact 14217 3706 14217 3706 6 state[1]
rlabel m2contact 14193 5698 14193 5698 6 n_170
rlabel m2contact 14169 5002 14169 5002 6 n_59
rlabel m2contact 14169 4402 14169 4402 6 n_61
rlabel m2contact 14145 2890 14145 2890 6 n_92
rlabel m2contact 14121 3202 14121 3202 6 n_58
rlabel m2contact 14097 3922 14097 3922 6 n_195
rlabel m2contact 14073 2386 14073 2386 6 n_244
rlabel m2contact 14073 7090 14073 7090 6 n_224
rlabel m2contact 14049 3754 14049 3754 6 n_232
rlabel m2contact 14049 4570 14049 4570 6 n_223
rlabel m2contact 14025 2218 14025 2218 6 n_200
rlabel m2contact 14001 2386 14001 2386 6 n_15
rlabel m2contact 14001 2914 14001 2914 6 n_234
rlabel m2contact 13977 3418 13977 3418 6 OpcodeCondIn[3]
rlabel m2contact 13953 3922 13953 3922 6 n_195
rlabel m2contact 13929 6442 13929 6442 6 n_145
rlabel m2contact 13905 6298 13905 6298 6 n_341
rlabel m2contact 13905 3754 13905 3754 6 n_190
rlabel m2contact 13881 4498 13881 4498 6 OpcodeCondIn[7]
rlabel m2contact 13857 2242 13857 2242 6 n_364
rlabel m2contact 13821 5914 13821 5914 6 n_240
rlabel m2contact 13821 1810 13821 1810 6 n_240
rlabel m2contact 13809 6274 13809 6274 6 n_181
rlabel m2contact 13785 2050 13785 2050 6 n_78
rlabel m2contact 13785 5002 13785 5002 6 n_184
rlabel m2contact 13761 5098 13761 5098 6 n_96
rlabel m2contact 13761 1834 13761 1834 6 n_96
rlabel m2contact 13737 7498 13737 7498 6 n_370
rlabel m2contact 13737 7042 13737 7042 6 n_53
rlabel m2contact 13713 6274 13713 6274 6 n_295
rlabel m2contact 13689 2050 13689 2050 6 n_347
rlabel m2contact 13665 7474 13665 7474 6 n_324
rlabel m2contact 13665 4018 13665 4018 6 nWait
rlabel m2contact 13641 7162 13641 7162 6 n_146
rlabel m2contact 13617 6442 13617 6442 4 n_145
rlabel m2contact 13593 4114 13593 4114 4 OpcodeCondIn[2]
rlabel m2contact 13569 2674 13569 2674 4 stateSub[1]
rlabel m2contact 13569 6058 13569 6058 4 n_185
rlabel m2contact 13545 6394 13545 6394 4 n_147
rlabel m2contact 13545 3826 13545 3826 4 n_125
rlabel m2contact 13521 5698 13521 5698 4 n_170
rlabel m2contact 13497 7330 13497 7330 4 n_244
rlabel m2contact 13473 2674 13473 2674 4 n_26
rlabel m2contact 13449 1978 13449 1978 4 n_132
rlabel m2contact 13425 4786 13425 4786 4 n_225
rlabel m2contact 13401 1858 13401 1858 4 n_82
rlabel m2contact 13401 5554 13401 5554 4 n_137
rlabel m2contact 13377 3226 13377 3226 4 OpcodeCondIn[4]
rlabel m2contact 13353 6442 13353 6442 4 n_75
rlabel m2contact 13353 3322 13353 3322 4 n_102
rlabel m2contact 13329 6394 13329 6394 4 n_56
rlabel m2contact 13329 1858 13329 1858 4 n_56
rlabel m2contact 13305 4426 13305 4426 4 n_183
rlabel m2contact 13281 4666 13281 4666 4 state[1]
rlabel m2contact 13281 4402 13281 4402 4 n_61
rlabel m2contact 13257 6082 13257 6082 4 stateSub[1]
rlabel m2contact 13233 5554 13233 5554 4 n_5
rlabel m2contact 13209 1810 13209 1810 4 n_240
rlabel m2contact 13209 3514 13209 3514 4 OpcodeCondIn[6]
rlabel m2contact 13185 1834 13185 1834 4 n_96
rlabel m2contact 13185 4354 13185 4354 4 stateSub[0]
rlabel m2contact 13161 6538 13161 6538 4 n_239
rlabel m2contact 13137 4666 13137 4666 4 n_101
rlabel m2contact 13113 1954 13113 1954 4 n_199
rlabel m2contact 13113 4834 13113 4834 4 n_63
rlabel m2contact 13089 7450 13089 7450 4 n_100
rlabel m2contact 13089 5218 13089 5218 4 n_162
rlabel m2contact 13065 5818 13065 5818 4 n_286
rlabel m2contact 13041 1954 13041 1954 4 n_107
rlabel m2contact 13017 3442 13017 3442 4 n_119
rlabel m2contact 12993 1858 12993 1858 4 n_56
rlabel m2contact 12993 4834 12993 4834 4 n_76
rlabel m2contact 12969 7426 12969 7426 4 n_394
rlabel m2contact 12945 7402 12945 7402 4 n_305
rlabel m2contact 12945 2962 12945 2962 4 StatusReg[2]
rlabel m2contact 12921 4354 12921 4354 4 stateSub[0]
rlabel m2contact 12897 1882 12897 1882 4 n_114
rlabel m2contact 12897 7378 12897 7378 4 n_278
rlabel m2contact 12873 5530 12873 5530 4 n_232
rlabel m2contact 12849 1906 12849 1906 4 n_71
rlabel m2contact 12849 6562 12849 6562 4 n_209
rlabel m2contact 12825 4906 12825 4906 4 n_154
rlabel m2contact 12801 1930 12801 1930 4 n_74
rlabel m2contact 12801 6202 12801 6202 4 n_233
rlabel m2contact 12777 3250 12777 3250 4 n_72
rlabel m2contact 12753 7306 12753 7306 4 n_304
rlabel m2contact 12753 6562 12753 6562 4 n_73
rlabel m2contact 12705 2410 12705 2410 4 n_66
rlabel m2contact 12705 7306 12705 7306 4 n_178
rlabel m2contact 12681 6802 12681 6802 4 n_279
rlabel m2contact 12681 4498 12681 4498 4 OpcodeCondIn[7]
rlabel m2contact 12657 4042 12657 4042 4 n_230
rlabel m2contact 12633 3154 12633 3154 4 n_110
rlabel m2contact 12609 6802 12609 6802 4 n_283
rlabel m2contact 12609 1930 12609 1930 4 n_283
rlabel m2contact 12585 2410 12585 2410 4 n_52
rlabel m2contact 12585 3922 12585 3922 4 n_195
rlabel m2contact 12561 1930 12561 1930 4 n_283
rlabel m2contact 12561 6010 12561 6010 4 stateSub[2]
rlabel m2contact 12537 5122 12537 5122 4 n_310
rlabel m2contact 12513 7378 12513 7378 4 CFlag
rlabel m2contact 12513 2074 12513 2074 4 CFlag
rlabel m2contact 12489 6298 12489 6298 4 n_341
rlabel m2contact 12465 4738 12465 4738 4 n_112
rlabel m2contact 12441 7378 12441 7378 4 CFlag
rlabel m2contact 12441 5506 12441 5506 4 n_308
rlabel m2contact 12393 5122 12393 5122 4 n_38
rlabel m2contact 12369 4354 12369 4354 4 stateSub[0]
rlabel m2contact 12345 1954 12345 1954 4 n_107
rlabel m2contact 12345 2578 12345 2578 4 n_36
rlabel m2contact 12321 6418 12321 6418 4 n_37
rlabel m2contact 12249 1978 12249 1978 4 n_132
rlabel m2contact 12201 2146 12201 2146 4 IntStatus
rlabel m2contact 12201 4066 12201 4066 4 n_192
rlabel m2contact 12153 6346 12153 6346 4 n_142
rlabel m2contact 12105 5314 12105 5314 4 n_47
rlabel m2contact 12081 6346 12081 6346 4 n_88
rlabel m2contact 12033 5314 12033 5314 4 n_245
rlabel m2contact 12009 7354 12009 7354 4 n_179
rlabel m2contact 11985 7330 11985 7330 4 n_244
rlabel m2contact 11937 3346 11937 3346 4 n_31
rlabel m2contact 11913 3514 11913 3514 4 OpcodeCondIn[6]
rlabel m2contact 11889 3250 11889 3250 4 n_72
rlabel m2contact 11841 2458 11841 2458 4 n_42
rlabel m2contact 11817 3226 11817 3226 4 OpcodeCondIn[4]
rlabel m2contact 11793 2458 11793 2458 4 n_25
rlabel m2contact 11745 2002 11745 2002 4 n_193
rlabel m2contact 11721 2794 11721 2794 4 n_191
rlabel m2contact 11697 4090 11697 4090 4 n_202
rlabel m2contact 11673 4066 11673 4066 4 n_192
rlabel m2contact 11625 5290 11625 5290 4 n_276
rlabel m2contact 11625 7138 11625 7138 4 n_300
rlabel m2contact 11601 3442 11601 3442 4 n_119
rlabel m2contact 11577 6178 11577 6178 4 n_116
rlabel m2contact 11577 5290 11577 5290 4 n_172
rlabel m2contact 11553 2026 11553 2026 4 n_149
rlabel m2contact 11553 3706 11553 3706 4 state[1]
rlabel m2contact 11529 4066 11529 4066 4 n_192
rlabel m2contact 11505 7306 11505 7306 4 n_178
rlabel m2contact 11505 5050 11505 5050 4 n_171
rlabel m2contact 11481 6178 11481 6178 4 n_139
rlabel m2contact 11457 7282 11457 7282 4 n_138
rlabel m2contact 11457 2218 11457 2218 4 n_200
rlabel m2contact 11409 4066 11409 4066 4 n_192
rlabel m2contact 11385 4138 11385 4138 4 n_157
rlabel m2contact 11361 7258 11361 7258 4 n_118
rlabel m2contact 11337 2050 11337 2050 4 n_347
rlabel m2contact 11337 6010 11337 6010 4 stateSub[2]
rlabel m2contact 11313 2074 11313 2074 4 CFlag
rlabel m2contact 11289 7234 11289 7234 4 n_211
rlabel m2contact 11289 6106 11289 6106 4 n_346
rlabel m2contact 11265 5866 11265 5866 4 n_115
rlabel m2contact 11241 2362 11241 2362 4 n_227
rlabel m2contact 11241 4618 11241 4618 4 n_207
rlabel m2contact 11217 2098 11217 2098 4 IRQ2
rlabel m2contact 11217 5866 11217 5866 4 n_58
rlabel m2contact 11217 3202 11217 3202 4 n_58
rlabel m2contact 11193 2122 11193 2122 4 n_168
rlabel m2contact 11193 2362 11193 2362 4 LrSel
rlabel m2contact 11169 4714 11169 4714 4 state[0]
rlabel m2contact 11145 2146 11145 2146 4 IntStatus
rlabel m2contact 11145 5746 11145 5746 4 n_128
rlabel m2contact 11121 2890 11121 2890 4 n_92
rlabel m2contact 11097 2170 11097 2170 4 Rs1Sel[1]
rlabel m2contact 11097 7018 11097 7018 4 n_30
rlabel m2contact 11073 5866 11073 5866 4 n_58
rlabel m2contact 11073 5746 11073 5746 4 n_357
rlabel m2contact 11025 2194 11025 2194 4 n_363
rlabel m2contact 11025 5866 11025 5866 4 n_204
rlabel m2contact 11001 2242 11001 2242 4 n_364
rlabel m2contact 11001 7210 11001 7210 4 n_124
rlabel m2contact 10977 3874 10977 3874 4 n_176
rlabel m2contact 10953 7210 10953 7210 4 ALE
rlabel m2contact 10953 2242 10953 2242 4 ALE
rlabel m2contact 10929 7210 10929 7210 4 ALE
rlabel m2contact 10929 5458 10929 5458 4 n_210
rlabel m2contact 10905 4570 10905 4570 4 n_223
rlabel m2contact 10881 2218 10881 2218 4 n_200
rlabel m2contact 10881 4810 10881 4810 4 RwSel[0]
rlabel m2contact 10857 2338 10857 2338 4 n_274
rlabel m2contact 10833 2242 10833 2242 4 ALE
rlabel m2contact 10833 7186 10833 7186 4 n_303
rlabel m2contact 10809 2266 10809 2266 4 n_117
rlabel m2contact 10809 4810 10809 4810 4 n_126
rlabel m2contact 10785 6466 10785 6466 4 n_213
rlabel m2contact 10737 2290 10737 2290 4 n_18
rlabel m2contact 10713 2314 10713 2314 4 n_32
rlabel m2contact 10713 4498 10713 4498 4 OpcodeCondIn[7]
rlabel m2contact 10689 4162 10689 4162 4 n_17
rlabel m2contact 10665 2338 10665 2338 4 n_274
rlabel m2contact 10641 4282 10641 4282 4 n_33
rlabel m2contact 10617 3082 10617 3082 4 n_324
rlabel m2contact 10617 3226 10617 3226 4 OpcodeCondIn[4]
rlabel m2contact 10593 2530 10593 2530 4 n_12
rlabel m2contact 10569 4282 10569 4282 4 n_323
rlabel m2contact 10545 4738 10545 4738 4 n_112
rlabel m2contact 10497 7162 10497 7162 4 n_146
rlabel m2contact 10497 6538 10497 6538 4 n_239
rlabel m2contact 10473 4210 10473 4210 4 n_46
rlabel m2contact 10425 3082 10425 3082 4 ImmSel
rlabel m2contact 10377 2314 10377 2314 4 nME
rlabel m2contact 10353 7162 10353 7162 4 OpcodeCondIn[6]
rlabel m2contact 10353 3514 10353 3514 4 OpcodeCondIn[6]
rlabel m2contact 10329 6058 10329 6058 4 n_185
rlabel m2contact 10329 2338 10329 2338 4 n_185
rlabel m2contact 10305 2314 10305 2314 4 nME
rlabel m2contact 10305 2794 10305 2794 4 n_191
rlabel m2contact 10281 4354 10281 4354 4 stateSub[0]
rlabel m2contact 10257 7162 10257 7162 4 OpcodeCondIn[6]
rlabel m2contact 10257 4738 10257 4738 4 n_289
rlabel m2contact 10233 4858 10233 4858 4 n_121
rlabel m2contact 10209 6514 10209 6514 4 n_236
rlabel m2contact 10185 2338 10185 2338 4 n_185
rlabel m2contact 10185 3418 10185 3418 4 OpcodeCondIn[3]
rlabel m2contact 10161 2794 10161 2794 4 n_191
rlabel m2contact 10137 4714 10137 4714 4 state[0]
rlabel m2contact 10113 6994 10113 6994 4 n_329
rlabel m2contact 10113 5818 10113 5818 4 n_286
rlabel m2contact 10065 7138 10065 7138 4 n_300
rlabel m2contact 10065 6994 10065 6994 4 IrWe
rlabel m2contact 10041 3010 10041 3010 4 n_255
rlabel m2contact 10017 4018 10017 4018 4 nWait
rlabel m2contact 9993 7114 9993 7114 4 n_298
rlabel m2contact 9993 3010 9993 3010 4 n_85
rlabel m2contact 9969 3298 9969 3298 4 n_338
rlabel m2contact 9945 7090 9945 7090 4 n_224
rlabel m2contact 9945 4834 9945 4834 4 n_76
rlabel m2contact 9921 7066 9921 7066 4 n_203
rlabel m2contact 9921 4570 9921 4570 4 n_223
rlabel m2contact 9921 2338 9921 2338 4 n_223
rlabel m2contact 9897 2674 9897 2674 4 n_26
rlabel m2contact 9897 4258 9897 4258 4 n_151
rlabel m2contact 9873 2722 9873 2722 4 n_79
rlabel m2contact 9849 2674 9849 2674 4 n_319
rlabel m2contact 9825 5338 9825 5338 4 n_318
rlabel m2contact 9801 2338 9801 2338 4 n_223
rlabel m2contact 9801 4258 9801 4258 4 n_269
rlabel m2contact 9777 6754 9777 6754 4 n_242
rlabel m2contact 9753 5266 9753 5266 4 n_150
rlabel m2contact 9753 3226 9753 3226 4 OpcodeCondIn[4]
rlabel m2contact 9705 5266 9705 5266 4 n_34
rlabel m2contact 9681 2362 9681 2362 4 LrSel
rlabel m2contact 9681 6514 9681 6514 4 n_236
rlabel m2contact 9657 2386 9657 2386 4 n_15
rlabel m2contact 9633 6754 9633 6754 4 n_326
rlabel m2contact 9609 2410 9609 2410 4 n_52
rlabel m2contact 9585 7042 9585 7042 4 n_53
rlabel m2contact 9585 6778 9585 6778 4 n_282
rlabel m2contact 9561 2722 9561 2722 4 n_79
rlabel m2contact 9537 3634 9537 3634 4 n_217
rlabel m2contact 9513 6994 9513 6994 4 IrWe
rlabel m2contact 9489 6778 9489 6778 4 n_282
rlabel m2contact 9489 2410 9489 2410 4 n_282
rlabel m2contact 9465 4354 9465 4354 4 stateSub[0]
rlabel m2contact 9441 2410 9441 2410 4 n_282
rlabel m2contact 9441 6562 9441 6562 4 n_73
rlabel m2contact 9417 5818 9417 5818 4 n_286
rlabel m2contact 9393 7018 9393 7018 4 n_30
rlabel m2contact 9393 6994 9393 6994 4 n_72
rlabel m2contact 9393 3250 9393 3250 4 n_72
rlabel m2contact 9369 6202 9369 6202 4 n_233
rlabel m2contact 9345 2458 9345 2458 4 n_25
rlabel m2contact 9321 6994 9321 6994 4 n_72
rlabel m2contact 9321 4426 9321 4426 4 n_183
rlabel m2contact 9297 4138 9297 4138 4 n_157
rlabel m2contact 9297 5698 9297 5698 4 n_170
rlabel m2contact 9225 4138 9225 4138 4 n_187
rlabel m2contact 9225 4090 9225 4090 4 n_202
rlabel m2contact 9201 6754 9201 6754 4 n_326
rlabel m2contact 9177 2434 9177 2434 4 n_131
rlabel m2contact 9153 2458 9153 2458 4 n_57
rlabel m2contact 9129 6370 9129 6370 4 n_55
rlabel m2contact 9105 6394 9105 6394 4 n_56
rlabel m2contact 9105 4234 9105 4234 4 n_268
rlabel m2contact 9057 2770 9057 2770 4 n_284
rlabel m2contact 9033 4642 9033 4642 4 n_155
rlabel m2contact 9009 2770 9009 2770 4 n_197
rlabel m2contact 8985 6970 8985 6970 4 n_238
rlabel m2contact 8985 6946 8985 6946 4 n_109
rlabel m2contact 8961 4642 8961 4642 4 n_208
rlabel m2contact 8913 6922 8913 6922 4 n_263
rlabel m2contact 8913 6346 8913 6346 4 n_88
rlabel m2contact 8865 6346 8865 6346 4 n_177
rlabel m2contact 8865 4978 8865 4978 4 n_182
rlabel m2contact 8841 2458 8841 2458 4 n_57
rlabel m2contact 8841 3106 8841 3106 4 n_196
rlabel m2contact 8793 5626 8793 5626 4 n_7
rlabel m2contact 8793 3106 8793 3106 4 n_152
rlabel m2contact 8745 4114 8745 4114 4 OpcodeCondIn[2]
rlabel m2contact 8721 3418 8721 3418 4 OpcodeCondIn[3]
rlabel m2contact 8673 2482 8673 2482 4 n_27
rlabel m2contact 8673 5722 8673 5722 4 n_372
rlabel m2contact 8649 5626 8649 5626 4 n_296
rlabel m2contact 8625 6898 8625 6898 4 n_348
rlabel m2contact 8625 4786 8625 4786 4 n_225
rlabel m2contact 8601 5722 8601 5722 4 n_325
rlabel m2contact 8553 5458 8553 5458 4 n_210
rlabel m2contact 8529 2506 8529 2506 4 n_180
rlabel m2contact 8529 3562 8529 3562 4 n_241
rlabel m2contact 8505 6058 8505 6058 4 n_185
rlabel m2contact 8481 2866 8481 2866 4 n_175
rlabel m2contact 8433 6874 8433 6874 4 n_159
rlabel m2contact 8409 4042 8409 4042 4 n_230
rlabel m2contact 8385 2530 8385 2530 4 n_12
rlabel m2contact 8385 4066 8385 4066 4 n_192
rlabel m2contact 8337 2554 8337 2554 4 n_77
rlabel m2contact 8337 2626 8337 2626 4 n_98
rlabel m2contact 8313 4474 8313 4474 4 n_252
rlabel m2contact 8289 2578 8289 2578 4 n_36
rlabel m2contact 8289 5698 8289 5698 4 n_170
rlabel m2contact 8265 3322 8265 3322 4 n_102
rlabel m2contact 8241 6850 8241 6850 4 n_153
rlabel m2contact 8241 5818 8241 5818 4 n_286
rlabel m2contact 8241 2578 8241 2578 4 n_286
rlabel m2contact 8217 3514 8217 3514 4 OpcodeCondIn[6]
rlabel m2contact 8193 2578 8193 2578 4 n_286
rlabel m2contact 8193 4066 8193 4066 4 n_192
rlabel m2contact 8145 3466 8145 3466 4 n_353
rlabel m2contact 8121 2938 8121 2938 4 n_44
rlabel m2contact 8097 3154 8097 3154 4 n_110
rlabel m2contact 8097 2794 8097 2794 4 n_191
rlabel m2contact 8073 6826 8073 6826 4 n_78
rlabel m2contact 8073 4066 8073 4066 4 n_192
rlabel m2contact 8025 2938 8025 2938 4 n_106
rlabel m2contact 8001 2626 8001 2626 4 n_98
rlabel m2contact 8001 3154 8001 3154 4 n_291
rlabel m2contact 7977 4786 7977 4786 4 n_225
rlabel m2contact 7953 4546 7953 4546 4 n_290
rlabel m2contact 7929 2602 7929 2602 4 n_120
rlabel m2contact 7929 4930 7929 4930 4 n_228
rlabel m2contact 7929 2626 7929 2626 4 n_228
rlabel m2contact 7905 6802 7905 6802 4 n_283
rlabel m2contact 7905 5218 7905 5218 4 n_162
rlabel m2contact 7881 2626 7881 2626 4 n_228
rlabel m2contact 7881 4786 7881 4786 4 n_225
rlabel m2contact 7857 6778 7857 6778 4 n_282
rlabel m2contact 7809 6754 7809 6754 4 n_326
rlabel m2contact 7809 3226 7809 3226 4 OpcodeCondIn[4]
rlabel m2contact 7785 3322 7785 3322 4 n_102
rlabel m2contact 7785 5458 7785 5458 4 n_210
rlabel m2contact 7761 5506 7761 5506 4 n_308
rlabel m2contact 7761 4498 7761 4498 4 OpcodeCondIn[7]
rlabel m2contact 7737 6754 7737 6754 4 state[1]
rlabel m2contact 7737 3706 7737 3706 4 state[1]
rlabel m2contact 7713 2650 7713 2650 4 n_29
rlabel m2contact 7713 5506 7713 5506 4 n_105
rlabel m2contact 7689 6754 7689 6754 4 state[1]
rlabel m2contact 7689 4786 7689 4786 4 n_225
rlabel m2contact 7665 6730 7665 6730 4 n_45
rlabel m2contact 7665 6082 7665 6082 4 stateSub[1]
rlabel m2contact 7593 6706 7593 6706 4 n_332
rlabel m2contact 7593 6682 7593 6682 4 n_35
rlabel m2contact 7545 2674 7545 2674 4 n_319
rlabel m2contact 7497 2674 7497 2674 4 Flags[2]
rlabel m2contact 7473 4474 7473 4474 4 n_252
rlabel m2contact 7425 6226 7425 6226 4 n_10
rlabel m2contact 7425 5818 7425 5818 4 n_286
rlabel m2contact 7377 2650 7377 2650 4 n_29
rlabel m2contact 7377 6226 7377 6226 4 n_322
rlabel m2contact 7353 2674 7353 2674 4 Flags[2]
rlabel m2contact 7329 2698 7329 2698 4 n_40
rlabel m2contact 7329 4282 7329 4282 4 n_323
rlabel m2contact 7305 3442 7305 3442 4 n_119
rlabel m2contact 7281 2722 7281 2722 4 n_79
rlabel m2contact 7281 6658 7281 6658 4 n_331
rlabel m2contact 7257 6634 7257 6634 4 n_231
rlabel m2contact 7233 2746 7233 2746 4 n_86
rlabel m2contact 7233 3154 7233 3154 4 n_291
rlabel m2contact 7209 3706 7209 3706 4 state[1]
rlabel m2contact 7185 6586 7185 6586 4 n_254
rlabel m2contact 7161 4474 7161 4474 4 n_252
rlabel m2contact 7137 2770 7137 2770 4 n_197
rlabel m2contact 7137 6610 7137 6610 4 n_253
rlabel m2contact 7113 2794 7113 2794 4 n_191
rlabel m2contact 7113 6586 7113 6586 4 n_249
rlabel m2contact 7113 3154 7113 3154 4 n_249
rlabel m2contact 7089 6586 7089 6586 4 n_249
rlabel m2contact 7089 4090 7089 4090 4 n_202
rlabel m2contact 7065 6562 7065 6562 4 n_73
rlabel m2contact 7065 4066 7065 4066 4 n_192
rlabel m2contact 7041 6538 7041 6538 4 n_239
rlabel m2contact 7017 6514 7017 6514 4 n_236
rlabel m2contact 6993 6490 6993 6490 4 n_140
rlabel m2contact 6969 6466 6969 6466 4 n_213
rlabel m2contact 6969 5458 6969 5458 4 n_210
rlabel m2contact 6945 2818 6945 2818 4 n_147
rlabel m2contact 6921 3442 6921 3442 4 n_119
rlabel m2contact 6897 6442 6897 6442 4 n_75
rlabel m2contact 6873 2818 6873 2818 4 n_147
rlabel m2contact 6849 4978 6849 4978 4 n_182
rlabel m2contact 6801 3682 6801 3682 4 OpcodeCondIn[1]
rlabel m2contact 6777 4186 6777 4186 4 OpcodeCondIn[0]
rlabel m2contact 6729 2842 6729 2842 4 n_80
rlabel m2contact 6705 6418 6705 6418 4 n_37
rlabel m2contact 6681 6394 6681 6394 4 n_56
rlabel m2contact 6657 6370 6657 6370 4 n_55
rlabel m2contact 6609 6130 6609 6130 4 n_362
rlabel m2contact 6609 4354 6609 4354 4 stateSub[0]
rlabel m2contact 6585 2866 6585 2866 4 n_175
rlabel m2contact 6585 4306 6585 4306 4 n_292
rlabel m2contact 6561 6130 6561 6130 4 n_344
rlabel m2contact 6537 4306 6537 4306 4 n_321
rlabel m2contact 6513 4906 6513 4906 4 n_154
rlabel m2contact 6489 6346 6489 6346 4 n_177
rlabel m2contact 6465 2890 6465 2890 4 n_92
rlabel m2contact 6465 3370 6465 3370 4 OpcodeCondIn[5]
rlabel m2contact 6441 6322 6441 6322 4 n_136
rlabel m2contact 6417 5146 6417 5146 4 n_123
rlabel m2contact 6393 6322 6393 6322 4 n_338
rlabel m2contact 6393 3298 6393 3298 4 n_338
rlabel m2contact 6369 6322 6369 6322 4 n_338
rlabel m2contact 6369 4978 6369 4978 4 n_182
rlabel m2contact 6345 6298 6345 6298 4 n_341
rlabel m2contact 6345 5458 6345 5458 4 n_210
rlabel m2contact 6321 3058 6321 3058 4 n_280
rlabel m2contact 6297 6274 6297 6274 4 n_295
rlabel m2contact 6273 3058 6273 3058 4 n_371
rlabel m2contact 6249 5962 6249 5962 4 n_293
rlabel m2contact 6249 3394 6249 3394 4 n_294
rlabel m2contact 6225 6250 6225 6250 4 n_345
rlabel m2contact 6201 6226 6201 6226 4 n_322
rlabel m2contact 6201 5962 6201 5962 4 n_235
rlabel m2contact 6153 6202 6153 6202 4 n_233
rlabel m2contact 6129 2914 6129 2914 4 n_234
rlabel m2contact 6129 4954 6129 4954 4 n_14
rlabel m2contact 6105 3682 6105 3682 4 OpcodeCondIn[1]
rlabel m2contact 6081 6202 6081 6202 4 OpcodeCondIn[6]
rlabel m2contact 6081 3514 6081 3514 4 OpcodeCondIn[6]
rlabel m2contact 6057 6202 6057 6202 4 OpcodeCondIn[6]
rlabel m2contact 6057 4954 6057 4954 4 n_256
rlabel m2contact 6033 4498 6033 4498 4 OpcodeCondIn[7]
rlabel m2contact 5961 6178 5961 6178 4 n_139
rlabel m2contact 5937 4354 5937 4354 4 stateSub[0]
rlabel m2contact 5913 2938 5913 2938 4 n_106
rlabel m2contact 5889 2962 5889 2962 4 StatusReg[2]
rlabel m2contact 5841 2986 5841 2986 4 n_392
rlabel m2contact 5841 3010 5841 3010 4 n_85
rlabel m2contact 5793 6154 5793 6154 4 n_84
rlabel m2contact 5745 6130 5745 6130 4 n_344
rlabel m2contact 5697 6106 5697 6106 4 n_346
rlabel m2contact 5649 3034 5649 3034 4 n_127
rlabel m2contact 5625 5146 5625 5146 4 n_123
rlabel m2contact 5601 6082 5601 6082 4 stateSub[1]
rlabel m2contact 5553 4954 5553 4954 4 n_256
rlabel m2contact 5505 3922 5505 3922 4 n_195
rlabel m2contact 5481 3058 5481 3058 4 n_371
rlabel m2contact 5481 6058 5481 6058 4 n_185
rlabel m2contact 5433 6034 5433 6034 4 n_20
rlabel m2contact 5409 3706 5409 3706 4 state[1]
rlabel m2contact 5385 6010 5385 6010 4 stateSub[2]
rlabel m2contact 5361 3082 5361 3082 4 ImmSel
rlabel m2contact 5361 4714 5361 4714 4 state[0]
rlabel m2contact 5337 5746 5337 5746 4 n_357
rlabel m2contact 5313 5170 5313 5170 4 n_359
rlabel m2contact 5289 3106 5289 3106 4 n_152
rlabel m2contact 5265 3154 5265 3154 4 n_249
rlabel m2contact 5265 5170 5265 5170 4 n_307
rlabel m2contact 5241 5986 5241 5986 4 n_277
rlabel m2contact 5217 3130 5217 3130 4 n_222
rlabel m2contact 5217 5962 5217 5962 4 n_235
rlabel m2contact 5217 5866 5217 5866 4 n_204
rlabel m2contact 5217 3154 5217 3154 4 n_204
rlabel m2contact 5193 4786 5193 4786 4 n_225
rlabel m2contact 5169 3154 5169 3154 4 n_204
rlabel m2contact 5169 4282 5169 4282 4 n_323
rlabel m2contact 5145 3274 5145 3274 4 n_158
rlabel m2contact 5121 5914 5121 5914 4 n_240
rlabel m2contact 5097 5938 5097 5938 4 n_206
rlabel m2contact 5097 3682 5097 3682 4 OpcodeCondIn[1]
rlabel m2contact 5073 3178 5073 3178 4 StatusReg[0]
rlabel m2contact 5073 5914 5073 5914 4 PcSel[2]
rlabel m2contact 5073 3274 5073 3274 4 PcSel[2]
rlabel m2contact 5049 5914 5049 5914 4 PcSel[2]
rlabel m2contact 5049 4186 5049 4186 4 OpcodeCondIn[0]
rlabel m2contact 5001 5890 5001 5890 4 n_395
rlabel m2contact 5001 3202 5001 3202 4 n_58
rlabel m2contact 4977 3226 4977 3226 4 OpcodeCondIn[4]
rlabel m2contact 4953 5866 4953 5866 4 n_204
rlabel m2contact 4953 3250 4953 3250 4 n_72
rlabel m2contact 4929 5842 4929 5842 4 n_219
rlabel m2contact 4881 3274 4881 3274 4 PcSel[2]
rlabel m2contact 4881 3850 4881 3850 4 n_261
rlabel m2contact 4833 3298 4833 3298 4 n_338
rlabel m2contact 4833 3922 4833 3922 4 n_195
rlabel m2contact 4809 5818 4809 5818 4 n_286
rlabel m2contact 4761 5794 4761 5794 4 n_334
rlabel m2contact 4761 3322 4761 3322 4 n_102
rlabel m2contact 4737 4954 4737 4954 4 n_256
rlabel m2contact 4713 3346 4713 3346 4 n_31
rlabel m2contact 4713 5770 4713 5770 4 n_218
rlabel m2contact 4665 5746 4665 5746 4 n_357
rlabel m2contact 4665 5722 4665 5722 4 n_325
rlabel m2contact 4641 4426 4641 4426 4 n_183
rlabel m2contact 4617 4954 4617 4954 4 n_256
rlabel m2contact 4617 4282 4617 4282 4 n_323
rlabel m2contact 4593 4042 4593 4042 4 n_230
rlabel m2contact 4569 5698 4569 5698 4 n_170
rlabel m2contact 4545 5218 4545 5218 4 n_162
rlabel m2contact 4521 5674 4521 5674 4 n_160
rlabel m2contact 4497 3370 4497 3370 4 OpcodeCondIn[5]
rlabel m2contact 4497 5650 4497 5650 4 n_113
rlabel m2contact 4473 4786 4473 4786 4 n_225
rlabel m2contact 4449 5626 4449 5626 4 n_296
rlabel m2contact 4425 5602 4425 5602 4 n_270
rlabel m2contact 4401 3394 4401 3394 4 n_294
rlabel m2contact 4401 4474 4401 4474 4 n_252
rlabel m2contact 4377 4234 4377 4234 4 n_268
rlabel m2contact 4329 5578 4329 5578 4 n_19
rlabel m2contact 4329 3418 4329 3418 4 OpcodeCondIn[3]
rlabel m2contact 4305 3442 4305 3442 4 n_119
rlabel m2contact 4305 3514 4305 3514 4 OpcodeCondIn[6]
rlabel m2contact 4281 4570 4281 4570 4 n_223
rlabel m2contact 4257 3802 4257 3802 4 n_285
rlabel m2contact 4233 5554 4233 5554 4 n_5
rlabel m2contact 4209 5530 4209 5530 4 n_232
rlabel m2contact 4209 3802 4209 3802 4 n_226
rlabel m2contact 4185 5506 4185 5506 4 n_105
rlabel m2contact 4161 5482 4161 5482 4 n_28
rlabel m2contact 4113 5458 4113 5458 4 n_210
rlabel m2contact 4113 3466 4113 3466 4 n_353
rlabel m2contact 4089 5434 4089 5434 4 n_229
rlabel m2contact 4065 4114 4065 4114 4 OpcodeCondIn[2]
rlabel m2contact 4041 5410 4041 5410 4 n_6
rlabel m2contact 4041 5386 4041 5386 4 n_89
rlabel m2contact 4017 5362 4017 5362 4 n_11
rlabel m2contact 3993 4594 3993 4594 4 n_361
rlabel m2contact 3969 5338 3969 5338 4 n_318
rlabel m2contact 3945 3490 3945 3490 4 n_83
rlabel m2contact 3945 4594 3945 4594 4 n_317
rlabel m2contact 3921 3514 3921 3514 4 OpcodeCondIn[6]
rlabel m2contact 3921 5314 3921 5314 4 n_245
rlabel m2contact 3897 5290 3897 5290 4 n_172
rlabel m2contact 3897 4426 3897 4426 4 n_183
rlabel m2contact 3849 3538 3849 3538 4 n_313
rlabel m2contact 3825 5266 3825 5266 4 n_34
rlabel m2contact 3801 5242 3801 5242 4 n_398
rlabel m2contact 3801 3562 3801 3562 4 n_241
rlabel m2contact 3777 3586 3777 3586 4 n_272
rlabel m2contact 3729 3610 3729 3610 4 n_81
rlabel m2contact 3705 5218 3705 5218 4 n_162
rlabel m2contact 3681 3634 3681 3634 4 n_217
rlabel m2contact 3681 4786 3681 4786 4 n_225
rlabel m2contact 3657 4906 3657 4906 4 n_154
rlabel m2contact 3609 5194 3609 5194 4 n_166
rlabel m2contact 3609 5170 3609 5170 4 n_307
rlabel m2contact 3585 4498 3585 4498 4 OpcodeCondIn[7]
rlabel m2contact 3561 5146 3561 5146 4 n_123
rlabel m2contact 3561 4282 3561 4282 4 n_323
rlabel m2contact 3513 3658 3513 3658 4 n_97
rlabel m2contact 3489 4162 3489 4162 4 n_17
rlabel m2contact 3465 5122 3465 5122 4 n_38
rlabel m2contact 3441 5098 3441 5098 4 n_96
rlabel m2contact 3441 3682 3441 3682 4 OpcodeCondIn[1]
rlabel m2contact 3393 3730 3393 3730 4 n_135
rlabel m2contact 3345 4522 3345 4522 4 n_67
rlabel m2contact 3321 4690 3321 4690 4 n_94
rlabel m2contact 3297 3706 3297 3706 4 state[1]
rlabel m2contact 3297 4786 3297 4786 4 n_225
rlabel m2contact 3297 3730 3297 3730 4 n_225
rlabel m2contact 3273 4690 3273 4690 4 n_265
rlabel m2contact 3249 3730 3249 3730 4 n_225
rlabel m2contact 3249 4426 3249 4426 4 n_183
rlabel m2contact 3225 3754 3225 3754 4 n_190
rlabel m2contact 3177 5074 3177 5074 4 n_251
rlabel m2contact 3153 5050 3153 5050 4 n_171
rlabel m2contact 3129 5026 3129 5026 4 n_212
rlabel m2contact 3081 5002 3081 5002 4 n_184
rlabel m2contact 3057 4978 3057 4978 4 n_182
rlabel m2contact 3033 4954 3033 4954 4 n_256
rlabel m2contact 3009 4930 3009 4930 4 n_228
rlabel m2contact 2985 4426 2985 4426 4 n_183
rlabel m2contact 2937 3778 2937 3778 4 n_69
rlabel m2contact 2913 4570 2913 4570 4 n_223
rlabel m2contact 2889 4906 2889 4906 4 n_154
rlabel m2contact 2889 4882 2889 4882 4 n_301
rlabel m2contact 2817 4858 2817 4858 4 n_121
rlabel m2contact 2769 4834 2769 4834 4 n_76
rlabel m2contact 2745 4810 2745 4810 4 n_126
rlabel m2contact 2721 3802 2721 3802 4 n_226
rlabel m2contact 2697 4786 2697 4786 4 n_225
rlabel m2contact 2697 3826 2697 3826 4 n_125
rlabel m2contact 2673 4762 2673 4762 4 n_174
rlabel m2contact 2625 4738 2625 4738 4 n_289
rlabel m2contact 2625 3850 2625 3850 4 n_261
rlabel m2contact 2601 4714 2601 4714 4 state[0]
rlabel m2contact 2601 3874 2601 3874 4 n_176
rlabel m2contact 2577 4690 2577 4690 4 n_265
rlabel m2contact 2553 4666 2553 4666 4 n_101
rlabel m2contact 2529 4642 2529 4642 4 n_208
rlabel m2contact 2505 3898 2505 3898 4 n_99
rlabel m2contact 2481 4618 2481 4618 4 n_207
rlabel m2contact 2433 4594 2433 4594 4 n_317
rlabel m2contact 2409 4570 2409 4570 4 n_223
rlabel m2contact 2385 4546 2385 4546 4 n_290
rlabel m2contact 2361 4354 2361 4354 4 stateSub[0]
rlabel m2contact 2337 4522 2337 4522 4 n_67
rlabel m2contact 2313 4498 2313 4498 4 OpcodeCondIn[7]
rlabel m2contact 2289 4474 2289 4474 4 n_252
rlabel m2contact 2289 4450 2289 4450 4 n_8
rlabel m2contact 2265 4114 2265 4114 4 OpcodeCondIn[2]
rlabel m2contact 2241 4354 2241 4354 4 stateSub[0]
rlabel m2contact 2217 4426 2217 4426 4 n_183
rlabel m2contact 2169 4402 2169 4402 4 n_61
rlabel m2contact 2121 4378 2121 4378 4 n_163
rlabel m2contact 2097 4354 2097 4354 4 stateSub[0]
rlabel m2contact 2073 4330 2073 4330 4 n_122
rlabel m2contact 2049 3922 2049 3922 4 n_195
rlabel m2contact 2025 4306 2025 4306 4 n_321
rlabel m2contact 2001 3946 2001 3946 4 Flags[3]
rlabel m2contact 1977 4282 1977 4282 4 n_323
rlabel m2contact 1929 4258 1929 4258 4 n_269
rlabel m2contact 1905 4042 1905 4042 4 n_230
rlabel m2contact 1881 4234 1881 4234 4 n_268
rlabel m2contact 1833 4210 1833 4210 4 n_46
rlabel m2contact 1785 4186 1785 4186 4 OpcodeCondIn[0]
rlabel m2contact 1761 4162 1761 4162 4 n_17
rlabel m2contact 1713 4138 1713 4138 4 n_187
rlabel m2contact 1689 3970 1689 3970 4 n_221
rlabel m2contact 1689 4114 1689 4114 4 OpcodeCondIn[2]
rlabel m2contact 1665 4090 1665 4090 4 n_202
rlabel m2contact 1641 4066 1641 4066 4 n_192
rlabel m2contact 1617 4042 1617 4042 4 n_230
rlabel metal2 25431 8588 25443 8588 6 StatusRegEn
rlabel metal2 24615 8588 24627 8588 6 StatusReg[0]
rlabel metal2 23799 8588 23811 8588 6 StatusReg[1]
rlabel metal2 23775 8588 23787 8588 6 StatusReg[2]
rlabel metal2 22167 8588 22179 8588 6 StatusReg[3]
rlabel metal2 22143 8588 22155 8588 6 AluEn
rlabel metal2 21327 8588 21339 8588 6 AluWe
rlabel metal2 20295 8588 20307 8588 6 Op2Sel[0]
rlabel metal2 19695 8588 19707 8588 6 Op2Sel[1]
rlabel metal2 18879 8588 18891 8588 6 Op1Sel
rlabel metal2 17271 8588 17283 8588 6 WdSel
rlabel metal2 16455 8588 16467 8588 6 PcEn
rlabel metal2 16239 8588 16251 8588 6 PcWe
rlabel metal2 15615 8588 15627 8588 6 PcSel[0]
rlabel metal2 14007 8588 14019 8588 6 PcSel[1]
rlabel metal2 13191 8588 13203 8588 4 PcSel[2]
rlabel metal2 13155 8588 13167 8588 4 LrEn
rlabel metal2 11535 8588 11547 8588 4 LrWe
rlabel metal2 11199 8588 11211 8588 4 LrSel
rlabel metal2 10431 8588 10443 8588 4 ImmSel
rlabel metal2 9519 8588 9531 8588 4 IrWe
rlabel metal2 9015 8588 9027 8588 4 MemEn
rlabel metal2 7395 8588 7407 8588 4 OpcodeCondIn[0]
rlabel metal2 6807 8588 6819 8588 4 OpcodeCondIn[1]
rlabel metal2 5739 8588 5751 8588 4 OpcodeCondIn[2]
rlabel metal2 5703 8588 5715 8588 4 OpcodeCondIn[3]
rlabel metal2 4875 8588 4887 8588 4 OpcodeCondIn[4]
rlabel metal2 4047 8588 4059 8588 4 OpcodeCondIn[5]
rlabel metal2 3219 8588 3231 8588 4 OpcodeCondIn[6]
rlabel metal2 2319 8588 2331 8588 4 OpcodeCondIn[7]
rlabel metal2 23007 0 23019 0 8 SysBus[3]
rlabel metal2 17463 0 17475 0 8 SysBus[2]
rlabel metal2 7815 0 7827 0 2 SysBus[1]
rlabel metal2 4431 0 4443 0 2 SysBus[0]
rlabel metal2 26953 83 26953 95 8 Flags[2]
rlabel metal2 26953 59 26953 71 8 Flags[1]
rlabel metal2 26953 35 26953 47 8 Flags[0]
rlabel metal2 26953 11 26953 23 8 CFlag
rlabel metal2 26953 4804 26953 4816 6 RwSel[0]
rlabel metal2 26953 1852 26953 1864 6 Rs1Sel[1]
rlabel metal2 26953 1828 26953 1840 6 Rs1Sel[0]
rlabel metal2 26953 1804 26953 1816 6 Flags[3]
rlabel metal2 26953 8421 26953 8433 6 ENB
rlabel metal2 26953 8397 26953 8409 6 AluOR[1]
rlabel metal2 26953 8373 26953 8385 6 AluOR[0]
rlabel metal2 26953 8349 26953 8361 6 RegWe
rlabel metal2 26953 8325 26953 8337 6 RwSel[1]
rlabel metal2 0 131 0 143 2 nWE
rlabel metal2 0 107 0 119 2 nIRQ
rlabel metal2 0 4012 0 4024 4 nWait
rlabel metal2 0 3988 0 4000 4 nOE
rlabel metal2 0 8469 0 8481 4 ALE
rlabel metal2 0 8445 0 8457 4 nME
rlabel metal2 26570 0 26770 0 1 GND!
rlabel metal2 26571 8588 26771 8588 5 GND!
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 123 8588 323 8588 5 Vdd!
rlabel metal2 411 8588 423 8588 5 nReset
rlabel metal2 363 8588 375 8588 5 Test
rlabel metal2 387 8588 399 8588 5 Clock
rlabel metal2 339 8588 351 8588 5 SDO
<< end >>
