magic
tech c035u
timestamp 1394117868
<< metal1 >>
rect 0 920 71 930
rect 85 920 191 930
rect 205 920 431 930
rect 445 920 767 930
rect 781 920 1007 930
rect 1021 920 1127 930
rect 1141 920 1343 930
rect 1357 920 1679 930
rect 0 898 47 908
rect 61 898 167 908
rect 181 898 551 908
rect 565 898 671 908
rect 685 898 887 908
rect 901 898 1223 908
rect 1237 898 1319 908
rect 1333 898 1559 908
rect 1573 898 1693 908
rect 0 875 23 885
rect 37 875 311 885
rect 325 875 407 885
rect 421 875 647 885
rect 661 875 863 885
rect 877 875 1103 885
rect 1117 875 1439 885
rect 1453 875 1535 885
rect 1549 875 1693 885
<< m2contact >>
rect 71 918 85 932
rect 191 918 205 932
rect 431 918 445 932
rect 767 918 781 932
rect 1007 918 1021 932
rect 1127 918 1141 932
rect 1343 918 1357 932
rect 1679 918 1693 932
rect 47 896 61 910
rect 167 896 181 910
rect 551 896 565 910
rect 671 896 685 910
rect 887 896 901 910
rect 1223 896 1237 910
rect 1319 896 1333 910
rect 1559 896 1573 910
rect 23 873 37 887
rect 311 873 325 887
rect 407 873 421 887
rect 647 873 661 887
rect 863 873 877 887
rect 1103 873 1117 887
rect 1439 873 1453 887
rect 1535 873 1549 887
<< metal2 >>
rect 24 844 36 873
rect 48 844 60 896
rect 72 844 84 918
rect 168 844 180 896
rect 192 844 204 918
rect 312 844 324 873
rect 408 844 420 873
rect 432 844 444 918
rect 552 844 564 896
rect 648 844 660 873
rect 672 844 684 896
rect 768 844 780 918
rect 864 844 876 873
rect 888 844 900 896
rect 1008 844 1020 918
rect 1104 844 1116 873
rect 1128 844 1140 918
rect 1224 844 1236 896
rect 1320 844 1332 896
rect 1344 844 1356 918
rect 1440 844 1452 873
rect 1536 844 1548 873
rect 1560 844 1572 896
rect 1680 844 1692 918
rect 120 0 132 45
rect 240 33 300 45
rect 360 0 372 45
rect 480 33 540 45
rect 600 0 612 45
rect 696 33 756 45
rect 816 0 828 45
rect 936 33 996 45
rect 1056 0 1068 45
rect 1152 33 1212 45
rect 1272 0 1284 45
rect 1368 33 1428 45
rect 1488 0 1500 45
rect 1608 33 1668 45
rect 1728 0 1740 45
use nor3 nor3_0
timestamp 1386235396
transform 1 0 0 0 1 45
box 0 0 144 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 144 0 1 45
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 264 0 1 45
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 384 0 1 45
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 504 0 1 45
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 624 0 1 45
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 720 0 1 45
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 840 0 1 45
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 960 0 1 45
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1080 0 1 45
box 0 0 96 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 1176 0 1 45
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 1296 0 1 45
box 0 0 96 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 1392 0 1 45
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 1512 0 1 45
box 0 0 120 799
use and2 and2_4
timestamp 1386234845
transform 1 0 1632 0 1 45
box 0 0 120 799
<< labels >>
rlabel metal1 0 920 0 930 4 In[2]
rlabel metal1 0 898 0 908 3 In[1]
rlabel metal1 0 875 0 885 3 In[0]
rlabel metal2 1728 0 1740 0 1 Out[7]
rlabel metal2 1488 0 1500 0 1 Out[6]
rlabel metal2 1272 0 1284 0 1 Out[5]
rlabel metal2 1056 0 1068 0 1 Out[4]
rlabel metal2 816 0 828 0 1 Out[3]
rlabel metal2 600 0 612 0 1 Out[2]
rlabel metal2 360 0 372 0 1 Out[1]
rlabel metal2 120 0 132 0 1 Out[0]
<< end >>
