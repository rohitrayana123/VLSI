magic
tech c035u
timestamp 1394299567
<< metal1 >>
rect 4045 1081 5495 1091
rect 5509 1081 14832 1091
rect -5 174 1464 184
rect -5 114 1487 124
rect 1501 114 5375 124
rect 5389 114 5543 124
rect 5557 114 14836 124
rect 2437 92 14836 102
rect 5101 70 14836 80
rect 14581 48 14836 58
rect 14797 26 14836 36
<< m2contact >>
rect 4031 1079 4045 1093
rect 5495 1079 5509 1093
rect 1487 112 1501 126
rect 5375 112 5389 126
rect 5543 112 5557 126
rect 2423 90 2437 104
rect 5087 68 5101 82
rect 14567 46 14581 60
rect 14783 24 14797 38
<< metal2 >>
rect 0 911 200 1098
rect 216 989 228 1098
rect 240 989 252 1098
rect 264 989 276 1098
rect 288 989 300 1098
rect 1536 1069 1548 1098
rect 2208 1069 2220 1098
rect 2256 1069 2268 1098
rect 2328 1069 2340 1098
rect 2688 1069 2700 1098
rect 2832 1069 2844 1098
rect 3048 1069 3060 1098
rect 3792 1069 3804 1098
rect 3960 1069 3972 1098
rect 4032 1069 4044 1079
rect 4344 1069 4356 1098
rect 4560 1069 4572 1098
rect 5304 1069 5316 1098
rect 5472 989 5484 1098
rect 5496 989 5508 1079
rect 5568 1069 5652 1081
rect 5688 1069 5700 1098
rect 6432 1069 6444 1098
rect 6648 1069 6660 1098
rect 6840 1069 6852 1098
rect 7584 1069 7596 1098
rect 7800 1069 7812 1098
rect 5568 989 5580 1069
rect 7992 1068 8004 1098
rect 8736 1069 8748 1098
rect 8952 1069 8964 1098
rect 9144 1069 9156 1098
rect 9888 1069 9900 1098
rect 10104 1069 10116 1098
rect 10296 1069 10308 1098
rect 11040 1069 11052 1098
rect 11256 1069 11268 1098
rect 11448 1069 11460 1098
rect 12192 1069 12204 1098
rect 12408 1069 12420 1098
rect 12600 1069 12612 1098
rect 13344 1069 13356 1098
rect 13560 1069 13572 1098
rect 13752 1068 13764 1098
rect 14496 1069 14508 1098
rect 14712 1068 14724 1098
rect 0 19 200 190
rect 216 19 228 190
rect 240 19 252 190
rect 264 19 276 190
rect 288 19 300 190
rect 1488 126 1500 130
rect 1536 19 1548 132
rect 2208 19 2220 131
rect 2256 19 2268 130
rect 2328 19 2340 130
rect 2424 104 2436 130
rect 2688 19 2700 130
rect 2832 19 2844 130
rect 3048 19 3060 130
rect 3792 19 3804 130
rect 3960 19 3972 133
rect 4344 19 4356 132
rect 4560 19 4572 132
rect 5088 82 5100 130
rect 5304 19 5316 130
rect 5376 126 5388 130
rect 5472 19 5484 190
rect 5544 126 5556 190
rect 5688 19 5700 141
rect 6432 19 6444 130
rect 6648 19 6660 130
rect 6840 19 6852 130
rect 7584 19 7596 130
rect 7800 19 7812 130
rect 7992 19 8004 130
rect 8736 19 8748 130
rect 8952 19 8964 130
rect 9144 19 9156 130
rect 9888 19 9900 130
rect 10104 19 10116 130
rect 10296 19 10308 130
rect 11040 19 11052 130
rect 11256 19 11268 130
rect 11448 19 11460 130
rect 12192 19 12204 131
rect 12408 19 12420 130
rect 12600 19 12612 131
rect 13344 19 13356 130
rect 13560 19 13572 130
rect 13752 19 13764 130
rect 14496 19 14508 130
rect 14568 60 14580 130
rect 14712 19 14724 130
rect 14784 38 14796 131
use leftbuf  leftbuf_0
timestamp 1386242881
transform 1 0 0 0 1 190
box 0 0 1464 799
use IrAA  IrAA_0
timestamp 1394294731
transform 1 0 1464 0 1 130
box 0 0 1008 939
use Pc_slice  Pc_slice_0
timestamp 1394294966
transform 1 0 2472 0 1 130
box 0 0 2952 939
use mux2  mux2_0
timestamp 1386235218
transform 1 0 5424 0 1 190
box 0 0 192 799
use regBlock_slice  regBlock_slice_0
timestamp 1394295027
transform 1 0 5616 0 1 130
box 0 0 9216 939
<< labels >>
rlabel metal1 5568 119 5568 119 1 SysBus
rlabel metal1 14830 1086 14830 1086 6 AluOut
rlabel metal1 14825 53 14825 53 1 Rd1
rlabel metal1 14827 30 14827 30 1 Rd2
rlabel metal2 0 19 200 19 1 Vdd!
rlabel metal2 216 19 228 19 1 SDI
rlabel metal2 240 19 252 19 1 Test
rlabel metal2 264 19 276 19 1 Clock
rlabel metal2 288 19 300 19 1 nReset
rlabel metal2 2328 19 2340 19 1 ImmSel
rlabel metal2 2256 19 2268 19 1 Ext1
rlabel metal2 2208 19 2220 19 1 Ext0
rlabel metal2 2688 19 2700 19 1 PcIncCin
rlabel metal2 2832 19 2844 19 1 LrSel
rlabel metal2 3048 19 3060 19 1 LrWe
rlabel metal2 3792 19 3804 19 1 LrEn
rlabel metal2 3960 19 3972 19 1 PcSel[0]
rlabel metal2 4344 19 4356 19 1 PcSel[1]
rlabel metal2 4560 19 4572 19 1 PcWe
rlabel metal2 5304 19 5316 19 1 PcEn
rlabel metal2 5472 19 5484 19 1 WdSel
rlabel metal2 5688 19 5700 19 1 Rq[0]
rlabel metal2 6432 19 6444 19 1 Rs1[0]
rlabel metal2 6648 19 6660 19 1 Ps2[0]
rlabel metal2 6840 19 6852 19 1 Rw[1]
rlabel metal2 7584 19 7596 19 1 Rs1[1]
rlabel metal2 7800 19 7812 19 1 Rs2[1]
rlabel metal2 7992 19 8004 19 1 Rw[2]
rlabel metal2 8736 19 8748 19 1 Rs1[2]
rlabel metal2 8952 19 8964 19 1 Rs2[2]
rlabel metal2 9144 19 9156 19 1 Rw[3]
rlabel metal2 9888 19 9900 19 1 Rs1[3]
rlabel metal2 10104 19 10116 19 1 Rs2[3]
rlabel metal2 10296 19 10308 19 1 Rw[4]
rlabel metal2 11040 19 11052 19 1 Rs1[4]
rlabel metal2 11256 19 11268 19 1 Rs2[4]
rlabel metal2 11448 19 11460 19 1 Rw[5]
rlabel metal2 12192 19 12204 19 1 Rs1[5]
rlabel metal2 12408 19 12420 19 1 Rs2[5]
rlabel metal2 12600 19 12612 19 1 Rw[6]
rlabel metal2 13344 19 13356 19 1 Rs1[6]
rlabel metal2 13560 19 13572 19 1 Rs2[6]
rlabel metal2 13752 19 13764 19 1 Rw[7]
rlabel metal2 14496 19 14508 19 1 Rs1[7]
rlabel metal2 14712 19 14724 19 1 Rs2[7]
rlabel metal2 1536 19 1548 19 1 IrWe
rlabel metal1 14824 119 14824 119 1 SysBus
rlabel metal1 14825 97 14825 97 1 Imm
rlabel metal1 14826 75 14826 75 1 Pc
rlabel metal2 14712 1098 14724 1098 5 Rs2[7]
rlabel metal2 14496 1098 14508 1098 5 Rs1[7]
rlabel metal2 13752 1098 13764 1098 5 Rw[7]
rlabel metal2 13560 1098 13572 1098 5 Rs2[6]
rlabel metal2 13344 1098 13356 1098 5 Rs1[6]
rlabel metal2 12600 1098 12612 1098 5 Rw[6]
rlabel metal2 12192 1098 12204 1098 5 Rs1[5]
rlabel metal2 12408 1098 12420 1098 5 Rs2[5]
rlabel metal2 11448 1098 11460 1098 5 Rw[5]
rlabel metal2 11256 1098 11268 1098 5 Rs2[4]
rlabel metal2 11040 1098 11052 1098 5 Rs1[4]
rlabel metal2 10296 1098 10308 1098 5 Rw[4]
rlabel metal2 10104 1098 10116 1098 5 Rs2[3]
rlabel metal2 9888 1098 9900 1098 5 Rs1[3]
rlabel metal2 9144 1098 9156 1098 5 Rw[3]
rlabel metal2 8952 1098 8964 1098 5 Rs2[2]
rlabel metal2 8736 1098 8748 1098 5 Rs1[2]
rlabel metal2 7992 1098 8004 1098 5 Rw[2]
rlabel metal2 7800 1098 7812 1098 5 Rs2[1]
rlabel metal2 7584 1098 7596 1098 5 Rs1[1]
rlabel metal2 6840 1098 6852 1098 5 Rw[1]
rlabel metal2 6648 1098 6660 1098 5 Rs2[0]
rlabel metal2 6432 1098 6444 1098 5 Rs1[0]
rlabel metal2 5688 1098 5700 1098 5 Rw[0]
rlabel metal2 5472 1098 5484 1098 5 WdSel
rlabel metal2 5304 1098 5316 1098 5 PcEn
rlabel metal2 4560 1098 4572 1098 5 PcWe
rlabel metal2 4344 1098 4356 1098 5 PcSel[1]
rlabel metal2 3960 1098 3972 1098 5 PcSel[0]
rlabel metal2 3792 1098 3804 1098 5 LrEn
rlabel metal2 3048 1098 3060 1098 5 LrWe
rlabel metal2 2832 1098 2844 1098 5 LrSel
rlabel metal2 2688 1098 2700 1098 5 PcIncCout
rlabel metal2 2328 1098 2340 1098 5 ImmSel
rlabel metal2 2256 1098 2268 1098 5 Ext1
rlabel metal2 2208 1098 2220 1098 5 Ext0
rlabel metal2 1536 1098 1548 1098 5 IrWe
rlabel metal2 0 1098 200 1098 5 Vdd!
rlabel metal2 216 1098 228 1098 5 SDO
rlabel metal2 240 1098 252 1098 5 Test
rlabel metal2 264 1098 276 1098 5 Clock
rlabel metal2 288 1098 300 1098 5 nReset
rlabel metal1 -5 114 -5 124 3 SysBus
rlabel metal1 -5 174 -5 184 3 Ir
<< end >>
