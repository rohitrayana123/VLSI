magic
tech c035u
timestamp 1395324901
<< nwell >>
rect 27769 7676 27842 8074
<< pwell >>
rect 27769 7275 27842 7676
<< metal1 >>
rect 18038 8228 18056 8242
rect 20390 8230 23520 8240
rect 2990 8206 3816 8216
rect 4814 8206 16464 8216
rect 16478 8206 17496 8216
rect 17510 8206 28196 8216
rect 84 8182 7872 8192
rect 8606 8182 14784 8192
rect 17630 8182 26808 8192
rect 84 8158 9960 8168
rect 10382 8158 11208 8168
rect 12578 8158 23688 8168
rect 24494 8158 26160 8168
rect 26174 8158 26784 8168
rect 84 8134 1752 8144
rect 2750 8134 12600 8144
rect 16622 8134 19152 8144
rect 19790 8134 28196 8144
rect 84 8110 5736 8120
rect 6662 8108 6680 8122
rect 6998 8110 21336 8120
rect 26750 8108 26768 8122
rect 26822 8110 28196 8120
rect 3794 8086 25008 8096
rect 26798 8086 28196 8096
rect 27769 8057 27842 8067
rect 27769 8034 27842 8044
rect 27769 7996 27842 8021
rect 27769 7351 27842 7376
rect 14270 7253 14472 7263
rect 18326 7253 25968 7263
rect 13622 7229 21000 7239
rect 21014 7229 21336 7239
rect 21350 7229 24120 7239
rect 24134 7229 26448 7239
rect 13142 7205 19536 7215
rect 12950 7181 15840 7191
rect 17870 7181 21744 7191
rect 12614 7157 14496 7167
rect 14510 7157 16104 7167
rect 16430 7157 23760 7167
rect 12518 7133 22296 7143
rect 12374 7109 19656 7119
rect 12278 7085 22704 7095
rect 22718 7085 24024 7095
rect 24038 7085 25560 7095
rect 12086 7061 18432 7071
rect 11582 7037 17664 7047
rect 17678 7037 19632 7047
rect 19646 7037 22992 7047
rect 11558 7013 11568 7023
rect 12014 7013 16416 7023
rect 17294 7013 17616 7023
rect 17702 7013 18312 7023
rect 11438 6989 27744 6999
rect 11390 6965 17016 6975
rect 17222 6965 21648 6975
rect 21662 6965 26112 6975
rect 11078 6941 13608 6951
rect 13910 6941 24144 6951
rect 11030 6917 14424 6927
rect 17150 6917 27288 6927
rect 10910 6893 19848 6903
rect 10526 6869 15480 6879
rect 15494 6869 21984 6879
rect 21998 6869 23832 6879
rect 10310 6845 13176 6855
rect 13382 6845 18144 6855
rect 18158 6845 24192 6855
rect 10190 6821 23448 6831
rect 23462 6821 23856 6831
rect 9830 6797 10032 6807
rect 10142 6797 11424 6807
rect 11438 6797 15984 6807
rect 15998 6797 18936 6807
rect 9662 6773 9672 6783
rect 9806 6773 18024 6783
rect 21326 6773 21456 6783
rect 21470 6773 21840 6783
rect 9182 6749 10680 6759
rect 10766 6749 24960 6759
rect 9158 6725 13896 6735
rect 13910 6725 14256 6735
rect 14270 6725 19056 6735
rect 19070 6725 21312 6735
rect 21326 6725 23760 6735
rect 23774 6725 26232 6735
rect 8966 6701 13008 6711
rect 13118 6701 13128 6711
rect 13214 6701 13344 6711
rect 13478 6701 19680 6711
rect 8798 6677 20328 6687
rect 8750 6653 23736 6663
rect 8414 6629 22128 6639
rect 7886 6605 7944 6615
rect 7958 6605 10488 6615
rect 10502 6605 11208 6615
rect 11222 6605 19512 6615
rect 19526 6605 25800 6615
rect 7838 6581 10296 6591
rect 10358 6581 25296 6591
rect 7742 6557 10944 6567
rect 11006 6557 24528 6567
rect 7646 6533 8208 6543
rect 8318 6533 13920 6543
rect 14078 6533 14400 6543
rect 15182 6533 16752 6543
rect 16766 6533 25872 6543
rect 7622 6509 9504 6519
rect 9590 6509 11136 6519
rect 11366 6509 23520 6519
rect 23534 6509 24456 6519
rect 7622 6485 24240 6495
rect 7598 6461 24864 6471
rect 7406 6437 13416 6447
rect 13430 6437 16824 6447
rect 16838 6437 19872 6447
rect 7286 6413 7776 6423
rect 7790 6413 8688 6423
rect 8702 6413 12360 6423
rect 12374 6413 16368 6423
rect 16382 6413 18960 6423
rect 18974 6413 19320 6423
rect 19334 6413 22032 6423
rect 22064 6413 22368 6423
rect 24830 6413 24876 6423
rect 7214 6389 24816 6399
rect 24830 6389 25776 6399
rect 7094 6365 10440 6375
rect 10454 6365 17784 6375
rect 17798 6365 19560 6375
rect 19574 6365 21696 6375
rect 21710 6365 23928 6375
rect 23942 6365 25392 6375
rect 6974 6341 16056 6351
rect 16694 6341 20616 6351
rect 6806 6317 6816 6327
rect 6926 6317 7320 6327
rect 7382 6317 15192 6327
rect 16262 6317 22536 6327
rect 6758 6293 10008 6303
rect 10022 6293 25296 6303
rect 6734 6269 11376 6279
rect 11390 6269 21408 6279
rect 21422 6269 21792 6279
rect 21806 6269 23856 6279
rect 6710 6245 7920 6255
rect 7934 6245 12504 6255
rect 12518 6245 14328 6255
rect 14342 6245 25104 6255
rect 6614 6221 14064 6231
rect 14078 6221 23592 6231
rect 6590 6197 13248 6207
rect 13262 6197 27336 6207
rect 6446 6173 7296 6183
rect 7310 6173 12480 6183
rect 12494 6173 13272 6183
rect 13286 6173 16392 6183
rect 16406 6173 19344 6183
rect 19358 6173 25680 6183
rect 25694 6173 26784 6183
rect 6326 6149 10632 6159
rect 10646 6149 24552 6159
rect 26294 6149 26328 6159
rect 6206 6125 26280 6135
rect 6206 6101 21264 6111
rect 6158 6077 12600 6087
rect 12614 6077 13056 6087
rect 13070 6077 14016 6087
rect 15158 6077 15216 6087
rect 16214 6077 16224 6087
rect 16646 6077 23616 6087
rect 6038 6053 21624 6063
rect 5990 6029 13728 6039
rect 14006 6029 14184 6039
rect 14990 6029 22944 6039
rect 5942 6005 21528 6015
rect 25622 6005 25980 6015
rect 5894 5981 11160 5991
rect 11270 5981 19968 5991
rect 25478 5981 25752 5991
rect 5846 5957 27456 5967
rect 5822 5933 13488 5943
rect 13502 5933 13512 5943
rect 13526 5933 13968 5943
rect 13982 5933 19248 5943
rect 19262 5933 21912 5943
rect 21926 5933 25464 5943
rect 25478 5933 25608 5943
rect 25622 5933 27024 5943
rect 5270 5909 25896 5919
rect 5174 5885 16776 5895
rect 16790 5885 17880 5895
rect 5126 5861 7056 5871
rect 7070 5861 7176 5871
rect 7190 5861 7368 5871
rect 7382 5861 13800 5871
rect 13814 5861 13992 5871
rect 14006 5861 15696 5871
rect 15710 5861 23160 5871
rect 23174 5861 24312 5871
rect 5030 5837 8784 5847
rect 8798 5837 9912 5847
rect 10118 5837 25008 5847
rect 4982 5813 8184 5823
rect 8246 5813 18192 5823
rect 24782 5813 24792 5823
rect 4934 5789 5400 5799
rect 5750 5789 5880 5799
rect 5942 5789 15000 5799
rect 15014 5789 25128 5799
rect 25142 5789 27264 5799
rect 27278 5789 27672 5799
rect 4886 5765 9432 5775
rect 9446 5765 13176 5775
rect 13190 5765 17424 5775
rect 17438 5765 26040 5775
rect 4862 5741 4968 5751
rect 4982 5741 8160 5751
rect 8174 5741 9240 5751
rect 9254 5741 11880 5751
rect 11894 5741 12096 5751
rect 12110 5741 13632 5751
rect 13646 5741 24768 5751
rect 4742 5717 9444 5727
rect 9458 5717 24336 5727
rect 4742 5693 11808 5703
rect 11966 5693 21384 5703
rect 21398 5693 23532 5703
rect 4694 5669 7872 5679
rect 8078 5669 25824 5679
rect 4694 5645 11112 5655
rect 11198 5645 27480 5655
rect 4670 5621 6216 5631
rect 6230 5621 16128 5631
rect 16142 5621 19728 5631
rect 19742 5621 23088 5631
rect 4646 5597 7416 5607
rect 7478 5597 9624 5607
rect 9638 5597 18912 5607
rect 4598 5573 10872 5583
rect 10886 5573 15168 5583
rect 15902 5573 27528 5583
rect 4598 5549 10728 5559
rect 10790 5549 19416 5559
rect 4550 5525 5664 5535
rect 5678 5525 5952 5535
rect 5966 5525 8808 5535
rect 8822 5525 11304 5535
rect 11318 5525 21192 5535
rect 4550 5501 15048 5511
rect 15110 5501 18744 5511
rect 18758 5501 24096 5511
rect 24110 5501 26472 5511
rect 4526 5477 17976 5487
rect 18182 5477 28196 5487
rect 4502 5453 12768 5463
rect 12830 5453 23352 5463
rect 4454 5429 19128 5439
rect 4358 5405 7248 5415
rect 7262 5405 24696 5415
rect 4310 5381 12240 5391
rect 12254 5381 21768 5391
rect 4262 5357 5352 5367
rect 5366 5357 15552 5367
rect 15566 5357 26136 5367
rect 4142 5333 9120 5343
rect 9134 5333 17904 5343
rect 18086 5333 19584 5343
rect 23270 5333 23496 5343
rect 4046 5309 5640 5319
rect 5654 5309 9576 5319
rect 9590 5309 9648 5319
rect 9710 5309 18048 5319
rect 18062 5309 22296 5319
rect 22310 5309 24504 5319
rect 24518 5309 25032 5319
rect 4022 5285 14832 5295
rect 14846 5285 23256 5295
rect 23270 5285 26016 5295
rect 3974 5261 12912 5271
rect 12926 5261 22416 5271
rect 3926 5237 3960 5247
rect 4022 5237 14040 5247
rect 14222 5237 18264 5247
rect 19094 5237 22608 5247
rect 22622 5237 25704 5247
rect 3854 5213 4440 5223
rect 4454 5213 7488 5223
rect 7502 5213 8712 5223
rect 8726 5213 13368 5223
rect 13382 5213 14208 5223
rect 14222 5213 18072 5223
rect 18086 5213 18576 5223
rect 18590 5213 19080 5223
rect 19094 5213 22848 5223
rect 22862 5213 24936 5223
rect 24950 5213 25080 5223
rect 3830 5189 12960 5199
rect 12974 5189 14232 5199
rect 14246 5189 18984 5199
rect 18998 5189 27072 5199
rect 27086 5189 27240 5199
rect 3806 5165 19224 5175
rect 3758 5141 5496 5151
rect 5558 5141 11544 5151
rect 11654 5141 22824 5151
rect 22838 5141 22992 5151
rect 3662 5117 11616 5127
rect 11774 5117 15312 5127
rect 15326 5117 19224 5127
rect 21566 5117 22068 5127
rect 23486 5117 23556 5127
rect 3590 5093 3624 5103
rect 3638 5093 4752 5103
rect 4766 5093 6432 5103
rect 6446 5093 10824 5103
rect 10838 5093 11232 5103
rect 11246 5093 12216 5103
rect 12230 5093 17376 5103
rect 17390 5093 20664 5103
rect 20678 5093 21888 5103
rect 21902 5093 23136 5103
rect 23150 5093 23616 5103
rect 23630 5093 25368 5103
rect 3542 5069 23472 5079
rect 23486 5069 23664 5079
rect 3446 5045 4416 5055
rect 4478 5045 9936 5055
rect 9950 5045 20112 5055
rect 21062 5045 21168 5055
rect 21374 5045 21960 5055
rect 3422 5021 3504 5031
rect 3518 5021 3720 5031
rect 3734 5021 5328 5031
rect 5342 5021 8376 5031
rect 8390 5021 12576 5031
rect 12590 5021 15384 5031
rect 15398 5021 20520 5031
rect 20534 5021 20712 5031
rect 20726 5021 25584 5031
rect 25598 5021 26160 5031
rect 26174 5021 26568 5031
rect 26582 5021 27552 5031
rect 3326 4997 19008 5007
rect 21038 4997 21840 5007
rect 21854 4997 25536 5007
rect 3278 4973 10560 4983
rect 10574 4973 24000 4983
rect 3254 4949 14088 4959
rect 14318 4949 19344 4959
rect 19478 4949 19488 4959
rect 20414 4949 23784 4959
rect 3182 4925 24432 4935
rect 3158 4901 7968 4911
rect 8030 4901 16320 4911
rect 16622 4901 16836 4911
rect 16982 4901 26196 4911
rect 3110 4877 4992 4887
rect 5054 4877 6576 4887
rect 6590 4877 19464 4887
rect 19478 4877 26592 4887
rect 2918 4853 5520 4863
rect 5534 4853 6384 4863
rect 6494 4853 6984 4863
rect 6998 4853 11280 4863
rect 11294 4853 13320 4863
rect 13334 4853 13464 4863
rect 13478 4853 13872 4863
rect 13886 4853 26256 4863
rect 2870 4829 11328 4839
rect 11342 4829 21552 4839
rect 22406 4829 22560 4839
rect 25238 4829 25440 4839
rect 2798 4805 13824 4815
rect 13838 4805 16200 4815
rect 16214 4805 21360 4815
rect 22358 4805 25752 4815
rect 2726 4781 5856 4791
rect 5870 4781 16512 4791
rect 16526 4781 16776 4791
rect 16934 4781 19008 4791
rect 19790 4781 22272 4791
rect 22334 4781 22464 4791
rect 25070 4781 25944 4791
rect 2702 4757 19800 4767
rect 19814 4757 27816 4767
rect 2678 4733 2976 4743
rect 2990 4733 7512 4743
rect 7574 4733 16800 4743
rect 16910 4733 20448 4743
rect 20846 4733 20868 4743
rect 20942 4733 21120 4743
rect 22118 4733 26952 4743
rect 2630 4709 13440 4719
rect 13598 4709 27384 4719
rect 2606 4685 12144 4695
rect 12158 4685 15912 4695
rect 16046 4685 16080 4695
rect 16166 4685 19392 4695
rect 19454 4685 20904 4695
rect 20918 4685 22200 4695
rect 22214 4685 23904 4695
rect 23918 4685 27768 4695
rect 2606 4661 6000 4671
rect 6062 4661 7848 4671
rect 7910 4661 10608 4671
rect 10622 4661 15264 4671
rect 15278 4661 21048 4671
rect 21062 4661 21288 4671
rect 21302 4661 22224 4671
rect 22238 4661 27696 4671
rect 2582 4637 25632 4647
rect 2534 4613 3048 4623
rect 3110 4613 7920 4623
rect 7934 4613 8016 4623
rect 8030 4613 9744 4623
rect 9758 4613 17688 4623
rect 17702 4613 18384 4623
rect 18398 4613 22392 4623
rect 22406 4613 25272 4623
rect 25934 4613 26400 4623
rect 27614 4613 27648 4623
rect 2510 4589 7056 4599
rect 7070 4589 15120 4599
rect 15134 4589 15240 4599
rect 15254 4589 15360 4599
rect 15374 4589 21432 4599
rect 21590 4589 23208 4599
rect 24326 4589 26736 4599
rect 26846 4589 26856 4599
rect 27086 4589 27840 4599
rect 2486 4565 13032 4575
rect 13238 4565 22068 4575
rect 22118 4565 27120 4575
rect 2414 4541 13824 4551
rect 13838 4541 18120 4551
rect 19166 4541 20280 4551
rect 20534 4541 25980 4551
rect 26078 4541 27168 4551
rect 2366 4517 19368 4527
rect 20990 4517 27624 4527
rect 2294 4493 2328 4503
rect 2390 4493 15960 4503
rect 16118 4493 24720 4503
rect 24950 4493 25512 4503
rect 25814 4493 26112 4503
rect 2270 4469 3936 4479
rect 3950 4469 9552 4479
rect 9566 4469 19944 4479
rect 19958 4469 20424 4479
rect 20438 4469 21456 4479
rect 21470 4469 24600 4479
rect 24614 4469 25488 4479
rect 2222 4445 26688 4455
rect 2174 4421 18480 4431
rect 18494 4421 21096 4431
rect 21446 4421 22044 4431
rect 23174 4421 23448 4431
rect 2150 4397 14448 4407
rect 14462 4397 23184 4407
rect 23198 4397 25656 4407
rect 25670 4397 26784 4407
rect 2126 4373 6408 4383
rect 6422 4373 6528 4383
rect 6542 4373 11856 4383
rect 11870 4373 12888 4383
rect 12902 4373 14136 4383
rect 14150 4373 15648 4383
rect 15662 4373 16176 4383
rect 16190 4373 17352 4383
rect 17366 4373 17904 4383
rect 17918 4373 20544 4383
rect 20558 4373 24072 4383
rect 2078 4349 5208 4359
rect 5222 4349 7680 4359
rect 7694 4349 12768 4359
rect 12782 4349 13080 4359
rect 13094 4349 17592 4359
rect 17870 4349 26904 4359
rect 2054 4325 9360 4335
rect 9494 4325 20784 4335
rect 21110 4325 21192 4335
rect 21614 4325 23640 4335
rect 1958 4301 9864 4311
rect 9974 4301 18720 4311
rect 18734 4301 26376 4311
rect 1934 4277 13776 4287
rect 14102 4277 16728 4287
rect 17438 4277 24840 4287
rect 1910 4253 2232 4263
rect 2246 4253 8136 4263
rect 8150 4253 16368 4263
rect 16382 4253 21072 4263
rect 21086 4253 21672 4263
rect 21686 4253 25248 4263
rect 25262 4253 27000 4263
rect 1910 4229 22152 4239
rect 1862 4205 8448 4215
rect 8510 4205 23424 4215
rect 1838 4181 6792 4191
rect 6806 4181 7992 4191
rect 8006 4181 19104 4191
rect 19118 4181 22008 4191
rect 22022 4181 25152 4191
rect 1814 4157 3984 4167
rect 3998 4157 4080 4167
rect 4094 4157 5136 4167
rect 5150 4157 12336 4167
rect 12350 4157 12456 4167
rect 12470 4157 17040 4167
rect 17054 4157 20592 4167
rect 20606 4157 21864 4167
rect 21878 4157 23064 4167
rect 23078 4157 26832 4167
rect 1790 4133 5568 4143
rect 5798 4133 26304 4143
rect 1766 4109 2832 4119
rect 2846 4109 3288 4119
rect 3302 4109 9768 4119
rect 9782 4109 10248 4119
rect 10262 4109 12480 4119
rect 12494 4109 12648 4119
rect 12662 4109 13536 4119
rect 13550 4109 13656 4119
rect 13670 4109 14280 4119
rect 14294 4109 16056 4119
rect 16070 4109 19296 4119
rect 19310 4109 21240 4119
rect 21254 4109 24576 4119
rect 1742 4085 5064 4095
rect 5126 4085 16296 4095
rect 16526 4085 16752 4095
rect 17606 4085 17664 4095
rect 21878 4085 22416 4095
rect 1718 4061 22584 4071
rect 1670 4037 11592 4047
rect 11966 4037 17304 4047
rect 17318 4037 24912 4047
rect 24926 4037 25056 4047
rect 1646 4013 17640 4023
rect 84 3989 16608 3999
rect 16694 3989 23304 3999
rect 84 3965 6240 3975
rect 6302 3965 25224 3975
rect 84 3941 6360 3951
rect 6542 3941 10896 3951
rect 10910 3941 12096 3951
rect 12110 3941 16536 3951
rect 16550 3941 18864 3951
rect 84 3917 7704 3927
rect 7766 3917 10848 3927
rect 10862 3917 15144 3927
rect 15422 3917 20304 3927
rect 1670 3893 11904 3903
rect 12014 3893 13392 3903
rect 13406 3893 19176 3903
rect 19190 3893 25440 3903
rect 1694 3869 22320 3879
rect 1694 3845 3384 3855
rect 3398 3845 25344 3855
rect 2006 3821 25320 3831
rect 2030 3797 21480 3807
rect 2270 3773 3600 3783
rect 3614 3773 9168 3783
rect 9182 3773 10536 3783
rect 10550 3773 11664 3783
rect 11678 3773 20688 3783
rect 2318 3749 2664 3759
rect 2678 3749 3480 3759
rect 3494 3749 4392 3759
rect 4406 3749 9528 3759
rect 9542 3749 11520 3759
rect 11534 3749 12432 3759
rect 12446 3749 13200 3759
rect 13214 3749 26928 3759
rect 2438 3725 25680 3735
rect 2462 3701 5064 3711
rect 5078 3701 13680 3711
rect 13694 3701 20832 3711
rect 2486 3677 4560 3687
rect 4574 3677 4896 3687
rect 4910 3677 12384 3687
rect 12398 3677 23400 3687
rect 23414 3677 23808 3687
rect 23822 3677 26856 3687
rect 2558 3653 4200 3663
rect 4214 3653 4296 3663
rect 4310 3653 9408 3663
rect 9422 3653 11496 3663
rect 11510 3653 12192 3663
rect 12206 3653 18240 3663
rect 18254 3653 21144 3663
rect 21158 3653 27576 3663
rect 2582 3629 7464 3639
rect 7478 3629 17832 3639
rect 17846 3629 20736 3639
rect 23414 3629 23532 3639
rect 2654 3605 2808 3615
rect 2822 3605 4656 3615
rect 4670 3605 6552 3615
rect 6566 3605 6864 3615
rect 6878 3605 7824 3615
rect 7838 3605 10512 3615
rect 10526 3605 11784 3615
rect 11798 3605 16440 3615
rect 16454 3605 19200 3615
rect 19214 3605 20760 3615
rect 20774 3605 22800 3615
rect 22814 3605 23376 3615
rect 23390 3605 25944 3615
rect 25958 3605 27600 3615
rect 2702 3581 2928 3591
rect 2942 3581 6072 3591
rect 6086 3581 18696 3591
rect 18710 3581 22464 3591
rect 2750 3557 10416 3567
rect 10430 3557 21216 3567
rect 2774 3533 7320 3543
rect 7334 3533 10152 3543
rect 10166 3533 22200 3543
rect 22214 3533 22512 3543
rect 22526 3533 23904 3543
rect 23918 3533 24408 3543
rect 24422 3533 24648 3543
rect 2846 3509 3360 3519
rect 3374 3509 7008 3519
rect 7022 3509 21936 3519
rect 21950 3509 22944 3519
rect 22958 3509 24048 3519
rect 24062 3509 24408 3519
rect 2870 3485 3912 3495
rect 3926 3485 4320 3495
rect 4334 3485 6840 3495
rect 6854 3485 9000 3495
rect 9086 3485 16584 3495
rect 16598 3485 17988 3495
rect 21230 3485 21744 3495
rect 24062 3485 24096 3495
rect 2918 3461 7152 3471
rect 7166 3461 12072 3471
rect 12086 3461 13296 3471
rect 13310 3461 15864 3471
rect 15878 3461 19104 3471
rect 3038 3437 12936 3447
rect 12998 3437 14184 3447
rect 14294 3437 16272 3447
rect 16574 3437 19032 3447
rect 3062 3413 7800 3423
rect 7814 3413 12168 3423
rect 12182 3413 13680 3423
rect 13694 3413 13848 3423
rect 13862 3413 20376 3423
rect 20390 3413 23832 3423
rect 3206 3389 13704 3399
rect 13790 3389 13920 3399
rect 14126 3389 22440 3399
rect 3230 3365 25968 3375
rect 3614 3341 3624 3351
rect 3710 3341 24504 3351
rect 24518 3341 25416 3351
rect 3662 3317 4224 3327
rect 4238 3317 9384 3327
rect 9398 3317 12552 3327
rect 12566 3317 17712 3327
rect 17726 3317 18504 3327
rect 18518 3317 23040 3327
rect 23054 3317 24624 3327
rect 25430 3317 26664 3327
rect 3806 3293 16704 3303
rect 16718 3293 17736 3303
rect 17846 3293 17880 3303
rect 22454 3293 22488 3303
rect 22502 3293 22608 3303
rect 3854 3269 3960 3279
rect 3974 3269 7248 3279
rect 7262 3269 14352 3279
rect 14366 3269 16032 3279
rect 16046 3269 24720 3279
rect 3878 3245 21672 3255
rect 3950 3221 7104 3231
rect 7166 3221 8664 3231
rect 8726 3221 8856 3231
rect 8942 3221 14160 3231
rect 14174 3221 15216 3231
rect 15230 3221 15720 3231
rect 15734 3221 18168 3231
rect 18182 3221 24168 3231
rect 4070 3197 6816 3207
rect 6830 3197 8904 3207
rect 8918 3197 10560 3207
rect 10574 3197 12312 3207
rect 12326 3197 13968 3207
rect 13982 3197 20088 3207
rect 4142 3173 20160 3183
rect 20174 3173 20640 3183
rect 20654 3173 24288 3183
rect 24302 3173 24600 3183
rect 4430 3149 6888 3159
rect 6902 3149 21504 3159
rect 4766 3125 5616 3135
rect 5630 3125 12672 3135
rect 12686 3125 13560 3135
rect 14438 3125 14496 3135
rect 14966 3125 24876 3135
rect 4814 3101 9720 3111
rect 9734 3101 10032 3111
rect 10046 3101 19704 3111
rect 19718 3101 26088 3111
rect 4886 3077 14376 3087
rect 14390 3077 23556 3087
rect 5006 3053 9024 3063
rect 9038 3053 12144 3063
rect 12158 3053 12456 3063
rect 12470 3053 13344 3063
rect 13358 3053 19992 3063
rect 5030 3029 13752 3039
rect 13766 3029 15672 3039
rect 15686 3029 18840 3039
rect 5102 3005 7512 3015
rect 7526 3005 11736 3015
rect 11750 3005 13944 3015
rect 13958 3005 22728 3015
rect 22742 3005 24528 3015
rect 5246 2981 5784 2991
rect 5846 2981 19488 2991
rect 5438 2957 20928 2967
rect 6038 2933 20952 2943
rect 20966 2933 23328 2943
rect 6086 2909 27864 2919
rect 6110 2885 27192 2895
rect 6182 2861 25008 2871
rect 6230 2837 18816 2847
rect 18830 2837 26496 2847
rect 6254 2813 17472 2823
rect 17726 2813 17784 2823
rect 6326 2789 17760 2799
rect 17774 2789 17808 2799
rect 6350 2765 22752 2775
rect 6374 2741 6384 2751
rect 6614 2741 6648 2751
rect 6710 2741 17256 2751
rect 17270 2741 27792 2751
rect 6662 2717 8592 2727
rect 8606 2717 8856 2727
rect 8870 2717 17568 2727
rect 17582 2717 23688 2727
rect 23702 2717 23976 2727
rect 6830 2693 6936 2703
rect 7046 2693 10080 2703
rect 10094 2693 23496 2703
rect 6926 2669 7392 2679
rect 7406 2669 8256 2679
rect 8270 2669 9672 2679
rect 9686 2669 10368 2679
rect 10382 2669 13296 2679
rect 13310 2669 16836 2679
rect 16850 2669 17952 2679
rect 17966 2669 18024 2679
rect 18038 2669 24216 2679
rect 24230 2669 26328 2679
rect 7118 2645 8616 2655
rect 8630 2645 11976 2655
rect 11990 2645 17928 2655
rect 7238 2621 9216 2631
rect 9230 2621 9312 2631
rect 9326 2621 10464 2631
rect 10478 2621 16296 2631
rect 16310 2621 16656 2631
rect 16670 2621 21984 2631
rect 21998 2621 24864 2631
rect 7358 2597 8568 2607
rect 8582 2597 10224 2607
rect 10334 2597 21720 2607
rect 7598 2573 22248 2583
rect 22262 2573 24264 2583
rect 7646 2549 28196 2559
rect 7814 2525 7872 2535
rect 7958 2525 26640 2535
rect 8174 2501 8208 2511
rect 8366 2501 20868 2511
rect 8486 2477 9192 2487
rect 9278 2477 17160 2487
rect 17942 2477 17988 2487
rect 8534 2453 10416 2463
rect 10694 2453 16872 2463
rect 16886 2453 21168 2463
rect 8750 2429 11712 2439
rect 12206 2429 12240 2439
rect 12350 2429 12408 2439
rect 12422 2429 12696 2439
rect 12710 2429 16080 2439
rect 16094 2429 18984 2439
rect 18998 2429 24696 2439
rect 24710 2429 25368 2439
rect 25382 2429 25488 2439
rect 8846 2405 18648 2415
rect 18662 2405 23952 2415
rect 23966 2405 27744 2415
rect 8966 2381 24384 2391
rect 9158 2357 14472 2367
rect 14486 2357 22176 2367
rect 22190 2357 25728 2367
rect 9350 2333 11064 2343
rect 11174 2333 11208 2343
rect 11270 2333 20856 2343
rect 20870 2333 21792 2343
rect 21806 2333 23520 2343
rect 23534 2333 25200 2343
rect 25214 2333 27648 2343
rect 9374 2309 9444 2319
rect 9566 2309 11568 2319
rect 11582 2309 15936 2319
rect 15950 2309 23232 2319
rect 23246 2309 26352 2319
rect 9422 2285 14400 2295
rect 15470 2285 17544 2295
rect 24398 2285 24456 2295
rect 9878 2261 16008 2271
rect 16022 2261 25272 2271
rect 25286 2261 25848 2271
rect 9902 2237 22656 2247
rect 25862 2237 26196 2247
rect 9902 2213 21816 2223
rect 10718 2189 17640 2199
rect 10862 2165 22560 2175
rect 10982 2141 23280 2151
rect 11030 2117 24792 2127
rect 11102 2093 26184 2103
rect 11486 2069 12912 2079
rect 13046 2069 19896 2079
rect 11606 2045 17088 2055
rect 11726 2021 15600 2031
rect 15614 2021 20064 2031
rect 20078 2021 25176 2031
rect 25190 2021 26544 2031
rect 12566 1997 20208 2007
rect 12590 1973 12600 1983
rect 12902 1973 12960 1983
rect 13094 1973 15288 1983
rect 16166 1973 16224 1983
rect 13334 1949 21960 1959
rect 13430 1925 21120 1935
rect 27878 1925 28196 1935
rect 13574 1901 13800 1911
rect 27854 1901 28196 1911
rect 12662 1068 13920 1078
rect 14150 1068 22224 1078
rect 11918 1044 15912 1054
rect 16478 1044 22584 1054
rect 11870 1020 12408 1030
rect 12614 1020 23592 1030
rect 11822 996 22128 1006
rect 11678 972 19320 982
rect 19766 972 26424 982
rect 11342 948 21168 958
rect 11150 924 23184 934
rect 9926 900 11832 910
rect 11894 900 22032 910
rect 22118 900 28196 910
rect 9614 876 19560 886
rect 19718 876 23640 886
rect 9494 852 17376 862
rect 17798 852 26088 862
rect 9470 828 17016 838
rect 17030 828 20376 838
rect 21830 828 27000 838
rect 9302 804 10608 814
rect 10622 804 20592 814
rect 20894 804 22608 814
rect 9038 780 18888 790
rect 18902 780 22080 790
rect 8150 756 25896 766
rect 7718 732 24216 742
rect 7430 708 10752 718
rect 10838 708 14472 718
rect 15518 708 19056 718
rect 19286 708 20952 718
rect 21734 708 23376 718
rect 23390 708 27024 718
rect 7286 684 10344 694
rect 10670 684 15840 694
rect 16262 684 25584 694
rect 6950 660 19824 670
rect 20558 660 24648 670
rect 24974 660 25992 670
rect 6782 636 10368 646
rect 10478 636 10800 646
rect 10934 636 25752 646
rect 6566 612 19440 622
rect 19454 612 21120 622
rect 21470 612 28196 622
rect 6422 588 12048 598
rect 12062 588 12720 598
rect 12734 588 22920 598
rect 24110 588 25572 598
rect 6302 564 6480 574
rect 6494 564 20736 574
rect 20798 564 21192 574
rect 21254 564 28196 574
rect 6182 540 22872 550
rect 23438 540 28196 550
rect 6158 516 16704 526
rect 16910 516 21768 526
rect 5966 492 19488 502
rect 5246 468 19608 478
rect 4934 444 7680 454
rect 8054 444 23136 454
rect 4646 420 24456 430
rect 4478 396 26976 406
rect 4358 372 12984 382
rect 14174 372 26232 382
rect 4262 348 13752 358
rect 14702 348 16152 358
rect 17822 348 18528 358
rect 4214 324 13272 334
rect 13286 324 16224 334
rect 16238 324 16320 334
rect 16334 324 19128 334
rect 19142 324 23400 334
rect 23414 324 23952 334
rect 23966 324 24432 334
rect 4190 300 9072 310
rect 9254 300 12816 310
rect 13022 300 20688 310
rect 3974 276 4848 286
rect 4862 276 8568 286
rect 8582 276 16752 286
rect 18374 276 23976 286
rect 23990 276 24168 286
rect 3782 252 10704 262
rect 10790 252 17976 262
rect 3014 228 12240 238
rect 12302 228 14592 238
rect 15806 228 21000 238
rect 2966 204 15000 214
rect 1646 180 13512 190
rect 84 156 19848 166
rect 84 132 1728 142
rect 2510 132 16848 142
rect 84 108 13128 118
rect 84 84 1776 94
rect 2798 84 9264 94
rect 9326 84 10356 94
rect 10958 84 11760 94
rect 11774 84 12264 94
rect 12278 84 16584 94
rect 16598 84 27048 94
rect 5798 60 16884 70
rect 9974 34 9992 48
rect 10190 36 17616 46
rect 17630 36 18600 46
rect 18614 36 21228 46
rect 21242 36 23712 46
rect 10982 12 14712 22
<< m2contact >>
rect 18024 8228 18038 8242
rect 20376 8228 20390 8242
rect 23520 8228 23534 8242
rect 2976 8204 2990 8218
rect 3816 8204 3830 8218
rect 4800 8204 4814 8218
rect 16464 8204 16478 8218
rect 17496 8204 17510 8218
rect 28196 8204 28210 8218
rect 70 8180 84 8194
rect 7872 8180 7886 8194
rect 8592 8180 8606 8194
rect 14784 8180 14798 8194
rect 17616 8180 17630 8194
rect 26808 8180 26822 8194
rect 70 8156 84 8170
rect 9960 8156 9974 8170
rect 10368 8156 10382 8170
rect 11208 8156 11222 8170
rect 12564 8156 12578 8170
rect 23688 8156 23702 8170
rect 24480 8156 24494 8170
rect 26160 8156 26174 8170
rect 26784 8156 26798 8170
rect 70 8132 84 8146
rect 1752 8132 1766 8146
rect 2736 8132 2750 8146
rect 12600 8132 12614 8146
rect 16608 8132 16622 8146
rect 19152 8132 19166 8146
rect 19776 8132 19790 8146
rect 28196 8132 28210 8146
rect 70 8108 84 8122
rect 5736 8108 5750 8122
rect 6648 8108 6662 8122
rect 6984 8108 6998 8122
rect 21336 8108 21350 8122
rect 26736 8108 26750 8122
rect 26808 8108 26822 8122
rect 28196 8108 28210 8122
rect 3780 8084 3794 8098
rect 25008 8084 25022 8098
rect 26784 8084 26798 8098
rect 28196 8084 28210 8098
rect 14256 7251 14270 7265
rect 14472 7251 14486 7265
rect 18312 7251 18326 7265
rect 25968 7251 25982 7265
rect 13608 7227 13622 7241
rect 21000 7227 21014 7241
rect 21336 7227 21350 7241
rect 24120 7227 24134 7241
rect 26448 7227 26462 7241
rect 13128 7203 13142 7217
rect 19536 7203 19550 7217
rect 12936 7179 12950 7193
rect 15840 7179 15854 7193
rect 17856 7179 17870 7193
rect 21744 7179 21758 7193
rect 12600 7155 12614 7169
rect 14496 7155 14510 7169
rect 16104 7155 16118 7169
rect 16416 7155 16430 7169
rect 23760 7155 23774 7169
rect 12504 7131 12518 7145
rect 22296 7131 22310 7145
rect 12360 7107 12374 7121
rect 19656 7107 19670 7121
rect 12264 7083 12278 7097
rect 22704 7083 22718 7097
rect 24024 7083 24038 7097
rect 25560 7083 25574 7097
rect 12072 7059 12086 7073
rect 18432 7059 18446 7073
rect 11568 7035 11582 7049
rect 17664 7035 17678 7049
rect 19632 7035 19646 7049
rect 22992 7035 23006 7049
rect 11544 7011 11558 7025
rect 11568 7011 11582 7025
rect 12000 7011 12014 7025
rect 16416 7011 16430 7025
rect 17280 7011 17294 7025
rect 17616 7011 17630 7025
rect 17688 7011 17702 7025
rect 18312 7011 18326 7025
rect 11424 6987 11438 7001
rect 27744 6987 27758 7001
rect 11376 6963 11390 6977
rect 17016 6963 17030 6977
rect 17208 6963 17222 6977
rect 21648 6963 21662 6977
rect 26112 6963 26126 6977
rect 11064 6939 11078 6953
rect 13608 6939 13622 6953
rect 13896 6939 13910 6953
rect 24144 6939 24158 6953
rect 11016 6915 11030 6929
rect 14424 6915 14438 6929
rect 17136 6915 17150 6929
rect 27288 6915 27302 6929
rect 10896 6891 10910 6905
rect 19848 6891 19862 6905
rect 10512 6867 10526 6881
rect 15480 6867 15494 6881
rect 21984 6867 21998 6881
rect 23832 6867 23846 6881
rect 10296 6843 10310 6857
rect 13176 6843 13190 6857
rect 13368 6843 13382 6857
rect 18144 6843 18158 6857
rect 24192 6843 24206 6857
rect 10176 6819 10190 6833
rect 23448 6819 23462 6833
rect 23856 6819 23870 6833
rect 9816 6795 9830 6809
rect 10032 6795 10046 6809
rect 10128 6795 10142 6809
rect 11424 6795 11438 6809
rect 15984 6795 15998 6809
rect 18936 6795 18950 6809
rect 9648 6771 9662 6785
rect 9672 6771 9686 6785
rect 9792 6771 9806 6785
rect 18024 6771 18038 6785
rect 21312 6771 21326 6785
rect 21456 6771 21470 6785
rect 21840 6771 21854 6785
rect 9168 6747 9182 6761
rect 10680 6747 10694 6761
rect 10752 6747 10766 6761
rect 24960 6747 24974 6761
rect 9144 6723 9158 6737
rect 13896 6723 13910 6737
rect 14256 6723 14270 6737
rect 19056 6723 19070 6737
rect 21312 6723 21326 6737
rect 23760 6723 23774 6737
rect 26232 6723 26246 6737
rect 8952 6699 8966 6713
rect 13008 6699 13022 6713
rect 13104 6699 13118 6713
rect 13128 6699 13142 6713
rect 13200 6699 13214 6713
rect 13344 6699 13358 6713
rect 13464 6699 13478 6713
rect 19680 6699 19694 6713
rect 8784 6675 8798 6689
rect 20328 6675 20342 6689
rect 8736 6651 8750 6665
rect 23736 6651 23750 6665
rect 8400 6627 8414 6641
rect 22128 6627 22142 6641
rect 7872 6603 7886 6617
rect 7944 6603 7958 6617
rect 10488 6603 10502 6617
rect 11208 6603 11222 6617
rect 19512 6603 19526 6617
rect 25800 6603 25814 6617
rect 7824 6579 7838 6593
rect 10296 6579 10310 6593
rect 10344 6579 10358 6593
rect 25296 6579 25310 6593
rect 7728 6555 7742 6569
rect 10944 6555 10958 6569
rect 10992 6555 11006 6569
rect 24528 6555 24542 6569
rect 7632 6531 7646 6545
rect 8208 6531 8222 6545
rect 8304 6531 8318 6545
rect 13920 6531 13934 6545
rect 14064 6531 14078 6545
rect 14400 6531 14414 6545
rect 15168 6531 15182 6545
rect 16752 6531 16766 6545
rect 25872 6531 25886 6545
rect 7608 6507 7622 6521
rect 9504 6507 9518 6521
rect 9576 6507 9590 6521
rect 11136 6507 11150 6521
rect 11352 6507 11366 6521
rect 23520 6507 23534 6521
rect 24456 6507 24470 6521
rect 7608 6483 7622 6497
rect 24240 6483 24254 6497
rect 7584 6459 7598 6473
rect 24864 6459 24878 6473
rect 7392 6435 7406 6449
rect 13416 6435 13430 6449
rect 16824 6435 16838 6449
rect 19872 6435 19886 6449
rect 7272 6411 7286 6425
rect 7776 6411 7790 6425
rect 8688 6411 8702 6425
rect 12360 6411 12374 6425
rect 16368 6411 16382 6425
rect 18960 6411 18974 6425
rect 19320 6411 19334 6425
rect 22032 6411 22064 6425
rect 22368 6411 22382 6425
rect 24816 6411 24830 6425
rect 24876 6411 24890 6425
rect 7200 6387 7214 6401
rect 24816 6387 24830 6401
rect 25776 6387 25790 6401
rect 7080 6363 7094 6377
rect 10440 6363 10454 6377
rect 17784 6363 17798 6377
rect 19560 6363 19574 6377
rect 21696 6363 21710 6377
rect 23928 6363 23942 6377
rect 25392 6363 25406 6377
rect 6960 6339 6974 6353
rect 16056 6339 16070 6353
rect 16680 6339 16694 6353
rect 20616 6339 20630 6353
rect 6792 6315 6806 6329
rect 6816 6315 6830 6329
rect 6912 6315 6926 6329
rect 7320 6315 7334 6329
rect 7368 6315 7382 6329
rect 15192 6315 15206 6329
rect 16248 6315 16262 6329
rect 22536 6315 22550 6329
rect 6744 6291 6758 6305
rect 10008 6291 10022 6305
rect 25296 6291 25310 6305
rect 6720 6267 6734 6281
rect 11376 6267 11390 6281
rect 21408 6267 21422 6281
rect 21792 6267 21806 6281
rect 23856 6267 23870 6281
rect 6696 6243 6710 6257
rect 7920 6243 7934 6257
rect 12504 6243 12518 6257
rect 14328 6243 14342 6257
rect 25104 6243 25118 6257
rect 6600 6219 6614 6233
rect 14064 6219 14078 6233
rect 23592 6219 23606 6233
rect 6576 6195 6590 6209
rect 13248 6195 13262 6209
rect 27336 6195 27350 6209
rect 6432 6171 6446 6185
rect 7296 6171 7310 6185
rect 12480 6171 12494 6185
rect 13272 6171 13286 6185
rect 16392 6171 16406 6185
rect 19344 6171 19358 6185
rect 25680 6171 25694 6185
rect 26784 6171 26798 6185
rect 6312 6147 6326 6161
rect 10632 6147 10646 6161
rect 24552 6147 24566 6161
rect 26280 6147 26294 6161
rect 26328 6147 26342 6161
rect 6192 6123 6206 6137
rect 26280 6123 26294 6137
rect 6192 6099 6206 6113
rect 21264 6099 21278 6113
rect 6144 6075 6158 6089
rect 12600 6075 12614 6089
rect 13056 6075 13070 6089
rect 14016 6075 14030 6089
rect 15144 6075 15158 6089
rect 15216 6075 15230 6089
rect 16200 6075 16214 6089
rect 16224 6075 16238 6089
rect 16632 6075 16646 6089
rect 23616 6075 23630 6089
rect 6024 6051 6038 6065
rect 21624 6051 21638 6065
rect 5976 6027 5990 6041
rect 13728 6027 13742 6041
rect 13992 6027 14006 6041
rect 14184 6027 14198 6041
rect 14976 6027 14990 6041
rect 22944 6027 22958 6041
rect 5928 6003 5942 6017
rect 21528 6003 21542 6017
rect 25608 6003 25622 6017
rect 25980 6003 25994 6017
rect 5880 5979 5894 5993
rect 11160 5979 11174 5993
rect 11256 5979 11270 5993
rect 19968 5979 19982 5993
rect 25464 5979 25478 5993
rect 25752 5979 25766 5993
rect 5832 5955 5846 5969
rect 27456 5955 27470 5969
rect 5808 5931 5822 5945
rect 13488 5931 13502 5945
rect 13512 5931 13526 5945
rect 13968 5931 13982 5945
rect 19248 5931 19262 5945
rect 21912 5931 21926 5945
rect 25464 5931 25478 5945
rect 25608 5931 25622 5945
rect 27024 5931 27038 5945
rect 5256 5907 5270 5921
rect 25896 5907 25910 5921
rect 5160 5883 5174 5897
rect 16776 5883 16790 5897
rect 17880 5883 17894 5897
rect 5112 5859 5126 5873
rect 7056 5859 7070 5873
rect 7176 5859 7190 5873
rect 7368 5859 7382 5873
rect 13800 5859 13814 5873
rect 13992 5859 14006 5873
rect 15696 5859 15710 5873
rect 23160 5859 23174 5873
rect 24312 5859 24326 5873
rect 5016 5835 5030 5849
rect 8784 5835 8798 5849
rect 9912 5835 9926 5849
rect 10104 5835 10118 5849
rect 25008 5835 25022 5849
rect 4968 5811 4982 5825
rect 8184 5811 8198 5825
rect 8232 5811 8246 5825
rect 18192 5811 18206 5825
rect 24768 5811 24782 5825
rect 24792 5811 24806 5825
rect 4920 5787 4934 5801
rect 5400 5787 5414 5801
rect 5736 5787 5750 5801
rect 5880 5787 5894 5801
rect 5928 5787 5942 5801
rect 15000 5787 15014 5801
rect 25128 5787 25142 5801
rect 27264 5787 27278 5801
rect 27672 5787 27686 5801
rect 4872 5763 4886 5777
rect 9432 5763 9446 5777
rect 13176 5763 13190 5777
rect 17424 5763 17438 5777
rect 26040 5763 26054 5777
rect 4848 5739 4862 5753
rect 4968 5739 4982 5753
rect 8160 5739 8174 5753
rect 9240 5739 9254 5753
rect 11880 5739 11894 5753
rect 12096 5739 12110 5753
rect 13632 5739 13646 5753
rect 24768 5739 24782 5753
rect 4728 5715 4742 5729
rect 9444 5715 9458 5729
rect 24336 5715 24350 5729
rect 4728 5691 4742 5705
rect 11808 5691 11822 5705
rect 11952 5691 11966 5705
rect 21384 5691 21398 5705
rect 23532 5691 23546 5705
rect 4680 5667 4694 5681
rect 7872 5667 7886 5681
rect 8064 5667 8078 5681
rect 25824 5667 25838 5681
rect 4680 5643 4694 5657
rect 11112 5643 11126 5657
rect 11184 5643 11198 5657
rect 27480 5643 27494 5657
rect 4656 5619 4670 5633
rect 6216 5619 6230 5633
rect 16128 5619 16142 5633
rect 19728 5619 19742 5633
rect 23088 5619 23102 5633
rect 4632 5595 4646 5609
rect 7416 5595 7430 5609
rect 7464 5595 7478 5609
rect 9624 5595 9638 5609
rect 18912 5595 18926 5609
rect 4584 5571 4598 5585
rect 10872 5571 10886 5585
rect 15168 5571 15182 5585
rect 15888 5571 15902 5585
rect 27528 5571 27542 5585
rect 4584 5547 4598 5561
rect 10728 5547 10742 5561
rect 10776 5547 10790 5561
rect 19416 5547 19430 5561
rect 4536 5523 4550 5537
rect 5664 5523 5678 5537
rect 5952 5523 5966 5537
rect 8808 5523 8822 5537
rect 11304 5523 11318 5537
rect 21192 5523 21206 5537
rect 4536 5499 4550 5513
rect 15048 5499 15062 5513
rect 15096 5499 15110 5513
rect 18744 5499 18758 5513
rect 24096 5499 24110 5513
rect 26472 5499 26486 5513
rect 4512 5475 4526 5489
rect 17976 5475 17990 5489
rect 18168 5475 18182 5489
rect 28196 5475 28210 5489
rect 4488 5451 4502 5465
rect 12768 5451 12782 5465
rect 12816 5451 12830 5465
rect 23352 5451 23366 5465
rect 4440 5427 4454 5441
rect 19128 5427 19142 5441
rect 4344 5403 4358 5417
rect 7248 5403 7262 5417
rect 24696 5403 24710 5417
rect 4296 5379 4310 5393
rect 12240 5379 12254 5393
rect 21768 5379 21782 5393
rect 4248 5355 4262 5369
rect 5352 5355 5366 5369
rect 15552 5355 15566 5369
rect 26136 5355 26150 5369
rect 4128 5331 4142 5345
rect 9120 5331 9134 5345
rect 17904 5331 17918 5345
rect 18072 5331 18086 5345
rect 19584 5331 19598 5345
rect 23256 5331 23270 5345
rect 23496 5331 23510 5345
rect 4032 5307 4046 5321
rect 5640 5307 5654 5321
rect 9576 5307 9590 5321
rect 9648 5307 9662 5321
rect 9696 5307 9710 5321
rect 18048 5307 18062 5321
rect 22296 5307 22310 5321
rect 24504 5307 24518 5321
rect 25032 5307 25046 5321
rect 4008 5283 4022 5297
rect 14832 5283 14846 5297
rect 23256 5283 23270 5297
rect 26016 5283 26030 5297
rect 3960 5259 3974 5273
rect 12912 5259 12926 5273
rect 22416 5259 22430 5273
rect 3912 5235 3926 5249
rect 3960 5235 3974 5249
rect 4008 5235 4022 5249
rect 14040 5235 14054 5249
rect 14208 5235 14222 5249
rect 18264 5235 18278 5249
rect 19080 5235 19094 5249
rect 22608 5235 22622 5249
rect 25704 5235 25718 5249
rect 3840 5211 3854 5225
rect 4440 5211 4454 5225
rect 7488 5211 7502 5225
rect 8712 5211 8726 5225
rect 13368 5211 13382 5225
rect 14208 5211 14222 5225
rect 18072 5211 18086 5225
rect 18576 5211 18590 5225
rect 19080 5211 19094 5225
rect 22848 5211 22862 5225
rect 24936 5211 24950 5225
rect 25080 5211 25094 5225
rect 3816 5187 3830 5201
rect 12960 5187 12974 5201
rect 14232 5187 14246 5201
rect 18984 5187 18998 5201
rect 27072 5187 27086 5201
rect 27240 5187 27254 5201
rect 3792 5163 3806 5177
rect 19224 5163 19238 5177
rect 3744 5139 3758 5153
rect 5496 5139 5510 5153
rect 5544 5139 5558 5153
rect 11544 5139 11558 5153
rect 11640 5139 11654 5153
rect 22824 5139 22838 5153
rect 22992 5139 23006 5153
rect 3648 5115 3662 5129
rect 11616 5115 11630 5129
rect 11760 5115 11774 5129
rect 15312 5115 15326 5129
rect 19224 5115 19238 5129
rect 21552 5115 21566 5129
rect 22068 5115 22082 5129
rect 23472 5115 23486 5129
rect 23556 5115 23570 5129
rect 3576 5091 3590 5105
rect 3624 5091 3638 5105
rect 4752 5091 4766 5105
rect 6432 5091 6446 5105
rect 10824 5091 10838 5105
rect 11232 5091 11246 5105
rect 12216 5091 12230 5105
rect 17376 5091 17390 5105
rect 20664 5091 20678 5105
rect 21888 5091 21902 5105
rect 23136 5091 23150 5105
rect 23616 5091 23630 5105
rect 25368 5091 25382 5105
rect 3528 5067 3542 5081
rect 23472 5067 23486 5081
rect 23664 5067 23678 5081
rect 3432 5043 3446 5057
rect 4416 5043 4430 5057
rect 4464 5043 4478 5057
rect 9936 5043 9950 5057
rect 20112 5043 20126 5057
rect 21048 5043 21062 5057
rect 21168 5043 21182 5057
rect 21360 5043 21374 5057
rect 21960 5043 21974 5057
rect 3408 5019 3422 5033
rect 3504 5019 3518 5033
rect 3720 5019 3734 5033
rect 5328 5019 5342 5033
rect 8376 5019 8390 5033
rect 12576 5019 12590 5033
rect 15384 5019 15398 5033
rect 20520 5019 20534 5033
rect 20712 5019 20726 5033
rect 25584 5019 25598 5033
rect 26160 5019 26174 5033
rect 26568 5019 26582 5033
rect 27552 5019 27566 5033
rect 3312 4995 3326 5009
rect 19008 4995 19022 5009
rect 21024 4995 21038 5009
rect 21840 4995 21854 5009
rect 25536 4995 25550 5009
rect 3264 4971 3278 4985
rect 10560 4971 10574 4985
rect 24000 4971 24014 4985
rect 3240 4947 3254 4961
rect 14088 4947 14102 4961
rect 14304 4947 14318 4961
rect 19344 4947 19358 4961
rect 19464 4947 19478 4961
rect 19488 4947 19502 4961
rect 20400 4947 20414 4961
rect 23784 4947 23798 4961
rect 3168 4923 3182 4937
rect 24432 4923 24446 4937
rect 3144 4899 3158 4913
rect 7968 4899 7982 4913
rect 8016 4899 8030 4913
rect 16320 4899 16334 4913
rect 16608 4899 16622 4913
rect 16836 4899 16850 4913
rect 16968 4899 16982 4913
rect 26196 4899 26210 4913
rect 3096 4875 3110 4889
rect 4992 4875 5006 4889
rect 5040 4875 5054 4889
rect 6576 4875 6590 4889
rect 19464 4875 19478 4889
rect 26592 4875 26606 4889
rect 2904 4851 2918 4865
rect 5520 4851 5534 4865
rect 6384 4851 6398 4865
rect 6480 4851 6494 4865
rect 6984 4851 6998 4865
rect 11280 4851 11294 4865
rect 13320 4851 13334 4865
rect 13464 4851 13478 4865
rect 13872 4851 13886 4865
rect 26256 4851 26270 4865
rect 2856 4827 2870 4841
rect 11328 4827 11342 4841
rect 21552 4827 21566 4841
rect 22392 4827 22406 4841
rect 22560 4827 22574 4841
rect 25224 4827 25238 4841
rect 25440 4827 25454 4841
rect 2784 4803 2798 4817
rect 13824 4803 13838 4817
rect 16200 4803 16214 4817
rect 21360 4803 21374 4817
rect 22344 4803 22358 4817
rect 25752 4803 25766 4817
rect 2712 4779 2726 4793
rect 5856 4779 5870 4793
rect 16512 4779 16526 4793
rect 16776 4779 16790 4793
rect 16920 4779 16934 4793
rect 19008 4779 19022 4793
rect 19776 4779 19790 4793
rect 22272 4779 22286 4793
rect 22320 4779 22334 4793
rect 22464 4779 22478 4793
rect 25056 4779 25070 4793
rect 25944 4779 25958 4793
rect 2688 4755 2702 4769
rect 19800 4755 19814 4769
rect 27816 4755 27830 4769
rect 2664 4731 2678 4745
rect 2976 4731 2990 4745
rect 7512 4731 7526 4745
rect 7560 4731 7574 4745
rect 16800 4731 16814 4745
rect 16896 4731 16910 4745
rect 20448 4731 20462 4745
rect 20832 4731 20846 4745
rect 20868 4731 20882 4745
rect 20928 4731 20942 4745
rect 21120 4731 21134 4745
rect 22104 4731 22118 4745
rect 26952 4731 26966 4745
rect 2616 4707 2630 4721
rect 13440 4707 13454 4721
rect 13584 4707 13598 4721
rect 27384 4707 27398 4721
rect 2592 4683 2606 4697
rect 12144 4683 12158 4697
rect 15912 4683 15926 4697
rect 16032 4683 16046 4697
rect 16080 4683 16094 4697
rect 16152 4683 16166 4697
rect 19392 4683 19406 4697
rect 19440 4683 19454 4697
rect 20904 4683 20918 4697
rect 22200 4683 22214 4697
rect 23904 4683 23918 4697
rect 27768 4683 27782 4697
rect 2592 4659 2606 4673
rect 6000 4659 6014 4673
rect 6048 4659 6062 4673
rect 7848 4659 7862 4673
rect 7896 4659 7910 4673
rect 10608 4659 10622 4673
rect 15264 4659 15278 4673
rect 21048 4659 21062 4673
rect 21288 4659 21302 4673
rect 22224 4659 22238 4673
rect 27696 4659 27710 4673
rect 2568 4635 2582 4649
rect 25632 4635 25646 4649
rect 2520 4611 2534 4625
rect 3048 4611 3062 4625
rect 3096 4611 3110 4625
rect 7920 4611 7934 4625
rect 8016 4611 8030 4625
rect 9744 4611 9758 4625
rect 17688 4611 17702 4625
rect 18384 4611 18398 4625
rect 22392 4611 22406 4625
rect 25272 4611 25286 4625
rect 25920 4611 25934 4625
rect 26400 4611 26414 4625
rect 27600 4611 27614 4625
rect 27648 4611 27662 4625
rect 2496 4587 2510 4601
rect 7056 4587 7070 4601
rect 15120 4587 15134 4601
rect 15240 4587 15254 4601
rect 15360 4587 15374 4601
rect 21432 4587 21446 4601
rect 21576 4587 21590 4601
rect 23208 4587 23222 4601
rect 24312 4587 24326 4601
rect 26736 4587 26750 4601
rect 26832 4587 26846 4601
rect 26856 4587 26870 4601
rect 27072 4587 27086 4601
rect 27840 4587 27854 4601
rect 2472 4563 2486 4577
rect 13032 4563 13046 4577
rect 13224 4563 13238 4577
rect 22068 4563 22082 4577
rect 22104 4563 22118 4577
rect 27120 4563 27134 4577
rect 2400 4539 2414 4553
rect 13824 4539 13838 4553
rect 18120 4539 18134 4553
rect 19152 4539 19166 4553
rect 20280 4539 20294 4553
rect 20520 4539 20534 4553
rect 25980 4539 25994 4553
rect 26064 4539 26078 4553
rect 27168 4539 27182 4553
rect 2352 4515 2366 4529
rect 19368 4515 19382 4529
rect 20976 4515 20990 4529
rect 27624 4515 27638 4529
rect 2280 4491 2294 4505
rect 2328 4491 2342 4505
rect 2376 4491 2390 4505
rect 15960 4491 15974 4505
rect 16104 4491 16118 4505
rect 24720 4491 24734 4505
rect 24936 4491 24950 4505
rect 25512 4491 25526 4505
rect 25800 4491 25814 4505
rect 26112 4491 26126 4505
rect 2256 4467 2270 4481
rect 3936 4467 3950 4481
rect 9552 4467 9566 4481
rect 19944 4467 19958 4481
rect 20424 4467 20438 4481
rect 21456 4467 21470 4481
rect 24600 4467 24614 4481
rect 25488 4467 25502 4481
rect 2208 4443 2222 4457
rect 26688 4443 26702 4457
rect 2160 4419 2174 4433
rect 18480 4419 18494 4433
rect 21096 4419 21110 4433
rect 21432 4419 21446 4433
rect 22044 4419 22058 4433
rect 23160 4419 23174 4433
rect 23448 4419 23462 4433
rect 2136 4395 2150 4409
rect 14448 4395 14462 4409
rect 23184 4395 23198 4409
rect 25656 4395 25670 4409
rect 26784 4395 26798 4409
rect 2112 4371 2126 4385
rect 6408 4371 6422 4385
rect 6528 4371 6542 4385
rect 11856 4371 11870 4385
rect 12888 4371 12902 4385
rect 14136 4371 14150 4385
rect 15648 4371 15662 4385
rect 16176 4371 16190 4385
rect 17352 4371 17366 4385
rect 17904 4371 17918 4385
rect 20544 4371 20558 4385
rect 24072 4371 24086 4385
rect 2064 4347 2078 4361
rect 5208 4347 5222 4361
rect 7680 4347 7694 4361
rect 12768 4347 12782 4361
rect 13080 4347 13094 4361
rect 17592 4347 17606 4361
rect 17856 4347 17870 4361
rect 26904 4347 26918 4361
rect 2040 4323 2054 4337
rect 9360 4323 9374 4337
rect 9480 4323 9494 4337
rect 20784 4323 20798 4337
rect 21096 4323 21110 4337
rect 21192 4323 21206 4337
rect 21600 4323 21614 4337
rect 23640 4323 23654 4337
rect 1944 4299 1958 4313
rect 9864 4299 9878 4313
rect 9960 4299 9974 4313
rect 18720 4299 18734 4313
rect 26376 4299 26390 4313
rect 1920 4275 1934 4289
rect 13776 4275 13790 4289
rect 14088 4275 14102 4289
rect 16728 4275 16742 4289
rect 17424 4275 17438 4289
rect 24840 4275 24854 4289
rect 1896 4251 1910 4265
rect 2232 4251 2246 4265
rect 8136 4251 8150 4265
rect 16368 4251 16382 4265
rect 21072 4251 21086 4265
rect 21672 4251 21686 4265
rect 25248 4251 25262 4265
rect 27000 4251 27014 4265
rect 1896 4227 1910 4241
rect 22152 4227 22166 4241
rect 1848 4203 1862 4217
rect 8448 4203 8462 4217
rect 8496 4203 8510 4217
rect 23424 4203 23438 4217
rect 1824 4179 1838 4193
rect 6792 4179 6806 4193
rect 7992 4179 8006 4193
rect 19104 4179 19118 4193
rect 22008 4179 22022 4193
rect 25152 4179 25166 4193
rect 1800 4155 1814 4169
rect 3984 4155 3998 4169
rect 4080 4155 4094 4169
rect 5136 4155 5150 4169
rect 12336 4155 12350 4169
rect 12456 4155 12470 4169
rect 17040 4155 17054 4169
rect 20592 4155 20606 4169
rect 21864 4155 21878 4169
rect 23064 4155 23078 4169
rect 26832 4155 26846 4169
rect 1776 4131 1790 4145
rect 5568 4131 5582 4145
rect 5784 4131 5798 4145
rect 26304 4131 26318 4145
rect 1752 4107 1766 4121
rect 2832 4107 2846 4121
rect 3288 4107 3302 4121
rect 9768 4107 9782 4121
rect 10248 4107 10262 4121
rect 12480 4107 12494 4121
rect 12648 4107 12662 4121
rect 13536 4107 13550 4121
rect 13656 4107 13670 4121
rect 14280 4107 14294 4121
rect 16056 4107 16070 4121
rect 19296 4107 19310 4121
rect 21240 4107 21254 4121
rect 24576 4107 24590 4121
rect 1728 4083 1742 4097
rect 5064 4083 5078 4097
rect 5112 4083 5126 4097
rect 16296 4083 16310 4097
rect 16512 4083 16526 4097
rect 16752 4083 16766 4097
rect 17592 4083 17606 4097
rect 17664 4083 17678 4097
rect 21864 4083 21878 4097
rect 22416 4083 22430 4097
rect 1704 4059 1718 4073
rect 22584 4059 22598 4073
rect 1656 4035 1670 4049
rect 11592 4035 11606 4049
rect 11952 4035 11966 4049
rect 17304 4035 17318 4049
rect 24912 4035 24926 4049
rect 25056 4035 25070 4049
rect 1632 4011 1646 4025
rect 17640 4011 17654 4025
rect 70 3987 84 4001
rect 16608 3987 16622 4001
rect 16680 3987 16694 4001
rect 23304 3987 23318 4001
rect 70 3963 84 3977
rect 6240 3963 6254 3977
rect 6288 3963 6302 3977
rect 25224 3963 25238 3977
rect 70 3939 84 3953
rect 6360 3939 6374 3953
rect 6528 3939 6542 3953
rect 10896 3939 10910 3953
rect 12096 3939 12110 3953
rect 16536 3939 16550 3953
rect 18864 3939 18878 3953
rect 70 3915 84 3929
rect 7704 3915 7718 3929
rect 7752 3915 7766 3929
rect 10848 3915 10862 3929
rect 15144 3915 15158 3929
rect 15408 3915 15422 3929
rect 20304 3915 20318 3929
rect 1656 3891 1670 3905
rect 11904 3891 11918 3905
rect 12000 3891 12014 3905
rect 13392 3891 13406 3905
rect 19176 3891 19190 3905
rect 25440 3891 25454 3905
rect 1680 3867 1694 3881
rect 22320 3867 22334 3881
rect 1680 3843 1694 3857
rect 3384 3843 3398 3857
rect 25344 3843 25358 3857
rect 1992 3819 2006 3833
rect 25320 3819 25334 3833
rect 2016 3795 2030 3809
rect 21480 3795 21494 3809
rect 2256 3771 2270 3785
rect 3600 3771 3614 3785
rect 9168 3771 9182 3785
rect 10536 3771 10550 3785
rect 11664 3771 11678 3785
rect 20688 3771 20702 3785
rect 2304 3747 2318 3761
rect 2664 3747 2678 3761
rect 3480 3747 3494 3761
rect 4392 3747 4406 3761
rect 9528 3747 9542 3761
rect 11520 3747 11534 3761
rect 12432 3747 12446 3761
rect 13200 3747 13214 3761
rect 26928 3747 26942 3761
rect 2424 3723 2438 3737
rect 25680 3723 25694 3737
rect 2448 3699 2462 3713
rect 5064 3699 5078 3713
rect 13680 3699 13694 3713
rect 20832 3699 20846 3713
rect 2472 3675 2486 3689
rect 4560 3675 4574 3689
rect 4896 3675 4910 3689
rect 12384 3675 12398 3689
rect 23400 3675 23414 3689
rect 23808 3675 23822 3689
rect 26856 3675 26870 3689
rect 2544 3651 2558 3665
rect 4200 3651 4214 3665
rect 4296 3651 4310 3665
rect 9408 3651 9422 3665
rect 11496 3651 11510 3665
rect 12192 3651 12206 3665
rect 18240 3651 18254 3665
rect 21144 3651 21158 3665
rect 27576 3651 27590 3665
rect 2568 3627 2582 3641
rect 7464 3627 7478 3641
rect 17832 3627 17846 3641
rect 20736 3627 20750 3641
rect 23400 3627 23414 3641
rect 23532 3627 23546 3641
rect 2640 3603 2654 3617
rect 2808 3603 2822 3617
rect 4656 3603 4670 3617
rect 6552 3603 6566 3617
rect 6864 3603 6878 3617
rect 7824 3603 7838 3617
rect 10512 3603 10526 3617
rect 11784 3603 11798 3617
rect 16440 3603 16454 3617
rect 19200 3603 19214 3617
rect 20760 3603 20774 3617
rect 22800 3603 22814 3617
rect 23376 3603 23390 3617
rect 25944 3603 25958 3617
rect 27600 3603 27614 3617
rect 2688 3579 2702 3593
rect 2928 3579 2942 3593
rect 6072 3579 6086 3593
rect 18696 3579 18710 3593
rect 22464 3579 22478 3593
rect 2736 3555 2750 3569
rect 10416 3555 10430 3569
rect 21216 3555 21230 3569
rect 2760 3531 2774 3545
rect 7320 3531 7334 3545
rect 10152 3531 10166 3545
rect 22200 3531 22214 3545
rect 22512 3531 22526 3545
rect 23904 3531 23918 3545
rect 24408 3531 24422 3545
rect 24648 3531 24662 3545
rect 2832 3507 2846 3521
rect 3360 3507 3374 3521
rect 7008 3507 7022 3521
rect 21936 3507 21950 3521
rect 22944 3507 22958 3521
rect 24048 3507 24062 3521
rect 24408 3507 24422 3521
rect 2856 3483 2870 3497
rect 3912 3483 3926 3497
rect 4320 3483 4334 3497
rect 6840 3483 6854 3497
rect 9000 3483 9014 3497
rect 9072 3483 9086 3497
rect 16584 3483 16598 3497
rect 17988 3483 18002 3497
rect 21216 3483 21230 3497
rect 21744 3483 21758 3497
rect 24048 3483 24062 3497
rect 24096 3483 24110 3497
rect 2904 3459 2918 3473
rect 7152 3459 7166 3473
rect 12072 3459 12086 3473
rect 13296 3459 13310 3473
rect 15864 3459 15878 3473
rect 19104 3459 19118 3473
rect 3024 3435 3038 3449
rect 12936 3435 12950 3449
rect 12984 3435 12998 3449
rect 14184 3435 14198 3449
rect 14280 3435 14294 3449
rect 16272 3435 16286 3449
rect 16560 3435 16574 3449
rect 19032 3435 19046 3449
rect 3048 3411 3062 3425
rect 7800 3411 7814 3425
rect 12168 3411 12182 3425
rect 13680 3411 13694 3425
rect 13848 3411 13862 3425
rect 20376 3411 20390 3425
rect 23832 3411 23846 3425
rect 3192 3387 3206 3401
rect 13704 3387 13718 3401
rect 13776 3387 13790 3401
rect 13920 3387 13934 3401
rect 14112 3387 14126 3401
rect 22440 3387 22454 3401
rect 3216 3363 3230 3377
rect 25968 3363 25982 3377
rect 3600 3339 3614 3353
rect 3624 3339 3638 3353
rect 3696 3339 3710 3353
rect 24504 3339 24518 3353
rect 25416 3339 25430 3353
rect 3648 3315 3662 3329
rect 4224 3315 4238 3329
rect 9384 3315 9398 3329
rect 12552 3315 12566 3329
rect 17712 3315 17726 3329
rect 18504 3315 18518 3329
rect 23040 3315 23054 3329
rect 24624 3315 24638 3329
rect 25416 3315 25430 3329
rect 26664 3315 26678 3329
rect 3792 3291 3806 3305
rect 16704 3291 16718 3305
rect 17736 3291 17750 3305
rect 17832 3291 17846 3305
rect 17880 3291 17894 3305
rect 22440 3291 22454 3305
rect 22488 3291 22502 3305
rect 22608 3291 22622 3305
rect 3840 3267 3854 3281
rect 3960 3267 3974 3281
rect 7248 3267 7262 3281
rect 14352 3267 14366 3281
rect 16032 3267 16046 3281
rect 24720 3267 24734 3281
rect 3864 3243 3878 3257
rect 21672 3243 21686 3257
rect 3936 3219 3950 3233
rect 7104 3219 7118 3233
rect 7152 3219 7166 3233
rect 8664 3219 8678 3233
rect 8712 3219 8726 3233
rect 8856 3219 8870 3233
rect 8928 3219 8942 3233
rect 14160 3219 14174 3233
rect 15216 3219 15230 3233
rect 15720 3219 15734 3233
rect 18168 3219 18182 3233
rect 24168 3219 24182 3233
rect 4056 3195 4070 3209
rect 6816 3195 6830 3209
rect 8904 3195 8918 3209
rect 10560 3195 10574 3209
rect 12312 3195 12326 3209
rect 13968 3195 13982 3209
rect 20088 3195 20102 3209
rect 4128 3171 4142 3185
rect 20160 3171 20174 3185
rect 20640 3171 20654 3185
rect 24288 3171 24302 3185
rect 24600 3171 24614 3185
rect 4416 3147 4430 3161
rect 6888 3147 6902 3161
rect 21504 3147 21518 3161
rect 4752 3123 4766 3137
rect 5616 3123 5630 3137
rect 12672 3123 12686 3137
rect 13560 3123 13574 3137
rect 14424 3123 14438 3137
rect 14496 3123 14510 3137
rect 14952 3123 14966 3137
rect 24876 3123 24890 3137
rect 4800 3099 4814 3113
rect 9720 3099 9734 3113
rect 10032 3099 10046 3113
rect 19704 3099 19718 3113
rect 26088 3099 26102 3113
rect 4872 3075 4886 3089
rect 14376 3075 14390 3089
rect 23556 3075 23570 3089
rect 4992 3051 5006 3065
rect 9024 3051 9038 3065
rect 12144 3051 12158 3065
rect 12456 3051 12470 3065
rect 13344 3051 13358 3065
rect 19992 3051 20006 3065
rect 5016 3027 5030 3041
rect 13752 3027 13766 3041
rect 15672 3027 15686 3041
rect 18840 3027 18854 3041
rect 5088 3003 5102 3017
rect 7512 3003 7526 3017
rect 11736 3003 11750 3017
rect 13944 3003 13958 3017
rect 22728 3003 22742 3017
rect 24528 3003 24542 3017
rect 5232 2979 5246 2993
rect 5784 2979 5798 2993
rect 5832 2979 5846 2993
rect 19488 2979 19502 2993
rect 5424 2955 5438 2969
rect 20928 2955 20942 2969
rect 6024 2931 6038 2945
rect 20952 2931 20966 2945
rect 23328 2931 23342 2945
rect 6072 2907 6086 2921
rect 27864 2907 27878 2921
rect 6096 2883 6110 2897
rect 27192 2883 27206 2897
rect 6168 2859 6182 2873
rect 25008 2859 25022 2873
rect 6216 2835 6230 2849
rect 18816 2835 18830 2849
rect 26496 2835 26510 2849
rect 6240 2811 6254 2825
rect 17472 2811 17486 2825
rect 17712 2811 17726 2825
rect 17784 2811 17798 2825
rect 6312 2787 6326 2801
rect 17760 2787 17774 2801
rect 17808 2787 17822 2801
rect 6336 2763 6350 2777
rect 22752 2763 22766 2777
rect 6360 2739 6374 2753
rect 6384 2739 6398 2753
rect 6600 2739 6614 2753
rect 6648 2739 6662 2753
rect 6696 2739 6710 2753
rect 17256 2739 17270 2753
rect 27792 2739 27806 2753
rect 6648 2715 6662 2729
rect 8592 2715 8606 2729
rect 8856 2715 8870 2729
rect 17568 2715 17582 2729
rect 23688 2715 23702 2729
rect 23976 2715 23990 2729
rect 6816 2691 6830 2705
rect 6936 2691 6950 2705
rect 7032 2691 7046 2705
rect 10080 2691 10094 2705
rect 23496 2691 23510 2705
rect 6912 2667 6926 2681
rect 7392 2667 7406 2681
rect 8256 2667 8270 2681
rect 9672 2667 9686 2681
rect 10368 2667 10382 2681
rect 13296 2667 13310 2681
rect 16836 2667 16850 2681
rect 17952 2667 17966 2681
rect 18024 2667 18038 2681
rect 24216 2667 24230 2681
rect 26328 2667 26342 2681
rect 7104 2643 7118 2657
rect 8616 2643 8630 2657
rect 11976 2643 11990 2657
rect 17928 2643 17942 2657
rect 7224 2619 7238 2633
rect 9216 2619 9230 2633
rect 9312 2619 9326 2633
rect 10464 2619 10478 2633
rect 16296 2619 16310 2633
rect 16656 2619 16670 2633
rect 21984 2619 21998 2633
rect 24864 2619 24878 2633
rect 7344 2595 7358 2609
rect 8568 2595 8582 2609
rect 10224 2595 10238 2609
rect 10320 2595 10334 2609
rect 21720 2595 21734 2609
rect 7584 2571 7598 2585
rect 22248 2571 22262 2585
rect 24264 2571 24278 2585
rect 7632 2547 7646 2561
rect 28196 2547 28210 2561
rect 7800 2523 7814 2537
rect 7872 2523 7886 2537
rect 7944 2523 7958 2537
rect 26640 2523 26654 2537
rect 8160 2499 8174 2513
rect 8208 2499 8222 2513
rect 8352 2499 8366 2513
rect 20868 2499 20882 2513
rect 8472 2475 8486 2489
rect 9192 2475 9206 2489
rect 9264 2475 9278 2489
rect 17160 2475 17174 2489
rect 17928 2475 17942 2489
rect 17988 2475 18002 2489
rect 8520 2451 8534 2465
rect 10416 2451 10430 2465
rect 10680 2451 10694 2465
rect 16872 2451 16886 2465
rect 21168 2451 21182 2465
rect 8736 2427 8750 2441
rect 11712 2427 11726 2441
rect 12192 2427 12206 2441
rect 12240 2427 12254 2441
rect 12336 2427 12350 2441
rect 12408 2427 12422 2441
rect 12696 2427 12710 2441
rect 16080 2427 16094 2441
rect 18984 2427 18998 2441
rect 24696 2427 24710 2441
rect 25368 2427 25382 2441
rect 25488 2427 25502 2441
rect 8832 2403 8846 2417
rect 18648 2403 18662 2417
rect 23952 2403 23966 2417
rect 27744 2403 27758 2417
rect 8952 2379 8966 2393
rect 24384 2379 24398 2393
rect 9144 2355 9158 2369
rect 14472 2355 14486 2369
rect 22176 2355 22190 2369
rect 25728 2355 25742 2369
rect 9336 2331 9350 2345
rect 11064 2331 11078 2345
rect 11160 2331 11174 2345
rect 11208 2331 11222 2345
rect 11256 2331 11270 2345
rect 20856 2331 20870 2345
rect 21792 2331 21806 2345
rect 23520 2331 23534 2345
rect 25200 2331 25214 2345
rect 27648 2331 27662 2345
rect 9360 2307 9374 2321
rect 9444 2307 9458 2321
rect 9552 2307 9566 2321
rect 11568 2307 11582 2321
rect 15936 2307 15950 2321
rect 23232 2307 23246 2321
rect 26352 2307 26366 2321
rect 9408 2283 9422 2297
rect 14400 2283 14414 2297
rect 15456 2283 15470 2297
rect 17544 2283 17558 2297
rect 24384 2283 24398 2297
rect 24456 2283 24470 2297
rect 9864 2259 9878 2273
rect 16008 2259 16022 2273
rect 25272 2259 25286 2273
rect 25848 2259 25862 2273
rect 9888 2235 9902 2249
rect 22656 2235 22670 2249
rect 25848 2235 25862 2249
rect 26196 2235 26210 2249
rect 9888 2211 9902 2225
rect 21816 2211 21830 2225
rect 10704 2187 10718 2201
rect 17640 2187 17654 2201
rect 10848 2163 10862 2177
rect 22560 2163 22574 2177
rect 10968 2139 10982 2153
rect 23280 2139 23294 2153
rect 11016 2115 11030 2129
rect 24792 2115 24806 2129
rect 11088 2091 11102 2105
rect 26184 2091 26198 2105
rect 11472 2067 11486 2081
rect 12912 2067 12926 2081
rect 13032 2067 13046 2081
rect 19896 2067 19910 2081
rect 11592 2043 11606 2057
rect 17088 2043 17102 2057
rect 11712 2019 11726 2033
rect 15600 2019 15614 2033
rect 20064 2019 20078 2033
rect 25176 2019 25190 2033
rect 26544 2019 26558 2033
rect 12552 1995 12566 2009
rect 20208 1995 20222 2009
rect 12576 1971 12590 1985
rect 12600 1971 12614 1985
rect 12888 1971 12902 1985
rect 12960 1971 12974 1985
rect 13080 1971 13094 1985
rect 15288 1971 15302 1985
rect 16152 1971 16166 1985
rect 16224 1971 16238 1985
rect 13320 1947 13334 1961
rect 21960 1947 21974 1961
rect 13416 1923 13430 1937
rect 21120 1923 21134 1937
rect 27864 1923 27878 1937
rect 28196 1923 28210 1937
rect 13560 1899 13574 1913
rect 13800 1899 13814 1913
rect 27840 1899 27854 1913
rect 28196 1899 28210 1913
rect 12648 1066 12662 1080
rect 13920 1066 13934 1080
rect 14136 1066 14150 1080
rect 22224 1066 22238 1080
rect 11904 1042 11918 1056
rect 15912 1042 15926 1056
rect 16464 1042 16478 1056
rect 22584 1042 22598 1056
rect 11856 1018 11870 1032
rect 12408 1018 12422 1032
rect 12600 1018 12614 1032
rect 23592 1018 23606 1032
rect 11808 994 11822 1008
rect 22128 994 22142 1008
rect 11664 970 11678 984
rect 19320 970 19334 984
rect 19752 970 19766 984
rect 26424 970 26438 984
rect 11328 946 11342 960
rect 21168 946 21182 960
rect 11136 922 11150 936
rect 23184 922 23198 936
rect 9912 898 9926 912
rect 11832 898 11846 912
rect 11880 898 11894 912
rect 22032 898 22046 912
rect 22104 898 22118 912
rect 28196 898 28210 912
rect 9600 874 9614 888
rect 19560 874 19574 888
rect 19704 874 19718 888
rect 23640 874 23654 888
rect 9480 850 9494 864
rect 17376 850 17390 864
rect 17784 850 17798 864
rect 26088 850 26102 864
rect 9456 826 9470 840
rect 17016 826 17030 840
rect 20376 826 20390 840
rect 21816 826 21830 840
rect 27000 826 27014 840
rect 9288 802 9302 816
rect 10608 802 10622 816
rect 20592 802 20606 816
rect 20880 802 20894 816
rect 22608 802 22622 816
rect 9024 778 9038 792
rect 18888 778 18902 792
rect 22080 778 22094 792
rect 8136 754 8150 768
rect 25896 754 25910 768
rect 7704 730 7718 744
rect 24216 730 24230 744
rect 7416 706 7430 720
rect 10752 706 10766 720
rect 10824 706 10838 720
rect 14472 706 14486 720
rect 15504 706 15518 720
rect 19056 706 19070 720
rect 19272 706 19286 720
rect 20952 706 20966 720
rect 21720 706 21734 720
rect 23376 706 23390 720
rect 27024 706 27038 720
rect 7272 682 7286 696
rect 10344 682 10358 696
rect 10656 682 10670 696
rect 15840 682 15854 696
rect 16248 682 16262 696
rect 25584 682 25598 696
rect 6936 658 6950 672
rect 19824 658 19838 672
rect 20544 658 20558 672
rect 24648 658 24662 672
rect 24960 658 24974 672
rect 25992 658 26006 672
rect 6768 634 6782 648
rect 10368 634 10382 648
rect 10464 634 10478 648
rect 10800 634 10814 648
rect 10920 634 10934 648
rect 25752 634 25766 648
rect 6552 610 6566 624
rect 19440 610 19454 624
rect 21120 610 21134 624
rect 21456 610 21470 624
rect 28196 610 28210 624
rect 6408 586 6422 600
rect 12048 586 12062 600
rect 12720 586 12734 600
rect 22920 586 22934 600
rect 24096 586 24110 600
rect 25572 586 25586 600
rect 6288 562 6302 576
rect 6480 562 6494 576
rect 20736 562 20750 576
rect 20784 562 20798 576
rect 21192 562 21206 576
rect 21240 562 21254 576
rect 28196 562 28210 576
rect 6168 538 6182 552
rect 22872 538 22886 552
rect 23424 538 23438 552
rect 28196 538 28210 552
rect 6144 514 6158 528
rect 16704 514 16718 528
rect 16896 514 16910 528
rect 21768 514 21782 528
rect 5952 490 5966 504
rect 19488 490 19502 504
rect 5232 466 5246 480
rect 19608 466 19622 480
rect 4920 442 4934 456
rect 7680 442 7694 456
rect 8040 442 8054 456
rect 23136 442 23150 456
rect 4632 418 4646 432
rect 24456 418 24470 432
rect 4464 394 4478 408
rect 26976 394 26990 408
rect 4344 370 4358 384
rect 12984 370 12998 384
rect 14160 370 14174 384
rect 26232 370 26246 384
rect 4248 346 4262 360
rect 13752 346 13766 360
rect 14688 346 14702 360
rect 16152 346 16166 360
rect 17808 346 17822 360
rect 18528 346 18542 360
rect 4200 322 4214 336
rect 13272 322 13286 336
rect 16224 322 16238 336
rect 16320 322 16334 336
rect 19128 322 19142 336
rect 23400 322 23414 336
rect 23952 322 23966 336
rect 24432 322 24446 336
rect 4176 298 4190 312
rect 9072 298 9086 312
rect 9240 298 9254 312
rect 12816 298 12830 312
rect 13008 298 13022 312
rect 20688 298 20702 312
rect 3960 274 3974 288
rect 4848 274 4862 288
rect 8568 274 8582 288
rect 16752 274 16766 288
rect 18360 274 18374 288
rect 23976 274 23990 288
rect 24168 274 24182 288
rect 3768 250 3782 264
rect 10704 250 10718 264
rect 10776 250 10790 264
rect 17976 250 17990 264
rect 3000 226 3014 240
rect 12240 226 12254 240
rect 12288 226 12302 240
rect 14592 226 14606 240
rect 15792 226 15806 240
rect 21000 226 21014 240
rect 2952 202 2966 216
rect 15000 202 15014 216
rect 1632 178 1646 192
rect 13512 178 13526 192
rect 70 154 84 168
rect 19848 154 19862 168
rect 70 130 84 144
rect 1728 130 1742 144
rect 2496 130 2510 144
rect 16848 130 16862 144
rect 70 106 84 120
rect 13128 106 13142 120
rect 70 82 84 96
rect 1776 82 1790 96
rect 2784 82 2798 96
rect 9264 82 9278 96
rect 9312 82 9326 96
rect 10356 82 10370 96
rect 10944 82 10958 96
rect 11760 82 11774 96
rect 12264 82 12278 96
rect 16584 82 16598 96
rect 27048 82 27062 96
rect 5784 58 5798 72
rect 16884 58 16898 72
rect 9960 34 9974 48
rect 10176 34 10190 48
rect 17616 34 17630 48
rect 18600 34 18614 48
rect 21228 34 21242 48
rect 23712 34 23726 48
rect 10968 10 10982 24
rect 14712 10 14726 24
<< metal2 >>
rect 0 8181 70 8193
rect 0 8157 70 8169
rect 0 8133 70 8145
rect 0 8109 70 8121
rect 145 8074 345 8252
rect 361 8074 373 8252
rect 385 8074 397 8252
rect 409 8074 421 8252
rect 433 8074 445 8252
rect 1753 8074 1765 8132
rect 2737 8074 2749 8132
rect 2977 8074 2989 8204
rect 3781 8098 3793 8252
rect 3817 8218 3829 8252
rect 4801 8074 4813 8204
rect 6661 8122 6673 8252
rect 6662 8108 6680 8122
rect 5737 8074 5749 8108
rect 6649 8074 6661 8108
rect 6985 8074 6997 8108
rect 7873 8074 7885 8180
rect 8593 8074 8605 8180
rect 10369 8170 10381 8252
rect 12565 8170 12577 8252
rect 9961 8074 9973 8156
rect 11209 8074 11221 8156
rect 12601 8146 12613 8252
rect 14785 8194 14797 8252
rect 18037 8242 18049 8252
rect 18038 8228 18056 8242
rect 16465 8074 16477 8204
rect 16609 8074 16621 8132
rect 17497 8074 17509 8204
rect 17617 8074 17629 8180
rect 18025 8074 18037 8228
rect 19153 8146 19165 8252
rect 19777 8074 19789 8132
rect 20377 8074 20389 8228
rect 21337 8122 21349 8252
rect 23521 8242 23533 8252
rect 23689 8074 23701 8156
rect 24481 8074 24493 8156
rect 25009 8074 25021 8084
rect 26161 8074 26173 8156
rect 26749 8122 26761 8252
rect 26750 8108 26768 8122
rect 26737 8074 26749 8108
rect 26785 8098 26797 8156
rect 26809 8122 26821 8180
rect 27961 8074 28161 8252
rect 28210 8205 28280 8217
rect 28210 8133 28280 8145
rect 28210 8109 28280 8121
rect 28210 8085 28280 8097
rect 0 3988 70 4000
rect 0 3964 70 3976
rect 0 3940 70 3952
rect 0 3916 70 3928
rect 145 1889 345 7275
rect 361 1889 373 7275
rect 385 1889 397 7275
rect 409 1889 421 7275
rect 433 1889 445 7275
rect 1633 4025 1645 7275
rect 1657 4049 1669 7275
rect 1657 1889 1669 3891
rect 1681 3881 1693 7275
rect 1705 4073 1717 7275
rect 1753 4121 1765 7275
rect 1801 4169 1813 7275
rect 1825 4193 1837 7275
rect 1849 4217 1861 7275
rect 1897 4265 1909 7275
rect 1921 4289 1933 7275
rect 1945 4313 1957 7275
rect 1681 1889 1693 3843
rect 1729 1889 1741 4083
rect 1777 1889 1789 4131
rect 1897 1889 1909 4227
rect 1993 3833 2005 7275
rect 2017 3809 2029 7275
rect 2041 4337 2053 7275
rect 2065 4361 2077 7275
rect 2113 4385 2125 7275
rect 2137 4409 2149 7275
rect 2161 4433 2173 7275
rect 2209 4457 2221 7275
rect 2233 4265 2245 7275
rect 2257 4481 2269 7275
rect 2281 4505 2293 7275
rect 2329 4505 2341 7275
rect 2353 4529 2365 7275
rect 2377 4505 2389 7275
rect 2401 4553 2413 7275
rect 2257 1889 2269 3771
rect 2305 1889 2317 3747
rect 2425 3737 2437 7275
rect 2473 4577 2485 7275
rect 2497 4601 2509 7275
rect 2521 4625 2533 7275
rect 2569 4649 2581 7275
rect 2593 4697 2605 7275
rect 2617 4721 2629 7275
rect 2665 4745 2677 7275
rect 2689 4769 2701 7275
rect 2713 4793 2725 7275
rect 2785 4817 2797 7275
rect 2449 1889 2461 3699
rect 2473 1889 2485 3675
rect 2545 1889 2557 3651
rect 2569 1889 2581 3627
rect 2593 1889 2605 4659
rect 2641 1889 2653 3603
rect 2665 1889 2677 3747
rect 2809 3617 2821 7275
rect 2833 4121 2845 7275
rect 2857 4841 2869 7275
rect 2905 4865 2917 7275
rect 2929 3593 2941 7275
rect 2689 1889 2701 3579
rect 2737 1889 2749 3555
rect 2761 1889 2773 3531
rect 2833 1889 2845 3507
rect 2857 1889 2869 3483
rect 2905 1889 2917 3459
rect 2977 1889 2989 4731
rect 3025 3449 3037 7275
rect 3049 4625 3061 7275
rect 3097 4889 3109 7275
rect 3145 4913 3157 7275
rect 3169 4937 3181 7275
rect 3049 1889 3061 3411
rect 3097 1889 3109 4611
rect 3193 3401 3205 7275
rect 3217 3377 3229 7275
rect 3265 4985 3277 7275
rect 3241 1889 3253 4947
rect 3289 4121 3301 7275
rect 3313 5009 3325 7275
rect 3361 3521 3373 7275
rect 3385 3857 3397 7275
rect 3409 5033 3421 7275
rect 3433 5057 3445 7275
rect 3481 3761 3493 7275
rect 3505 5033 3517 7275
rect 3529 5081 3541 7275
rect 3577 5105 3589 7275
rect 3601 3785 3613 7275
rect 3649 5129 3661 7275
rect 3625 3353 3637 5091
rect 3697 3353 3709 7275
rect 3721 5033 3733 7275
rect 3745 5153 3757 7275
rect 3793 5177 3805 7275
rect 3817 5201 3829 7275
rect 3841 5225 3853 7275
rect 3601 1889 3613 3339
rect 3649 1889 3661 3315
rect 3793 1889 3805 3291
rect 3841 1889 3853 3267
rect 3865 3257 3877 7275
rect 3913 5249 3925 7275
rect 3937 4481 3949 7275
rect 3961 5273 3973 7275
rect 4009 5297 4021 7275
rect 4033 5321 4045 7275
rect 4129 5345 4141 7275
rect 3913 1889 3925 3483
rect 3961 3281 3973 5235
rect 3937 1889 3949 3219
rect 3985 1889 3997 4155
rect 4009 1889 4021 5235
rect 4057 1889 4069 3195
rect 4081 1889 4093 4155
rect 4201 3665 4213 7275
rect 4225 3329 4237 7275
rect 4249 5369 4261 7275
rect 4297 5393 4309 7275
rect 4345 5417 4357 7275
rect 4417 5057 4429 7275
rect 4441 5441 4453 7275
rect 4129 1889 4141 3171
rect 4297 1889 4309 3651
rect 4321 1889 4333 3483
rect 4393 1889 4405 3747
rect 4417 1889 4429 3147
rect 4441 1889 4453 5211
rect 4465 5057 4477 7275
rect 4489 5465 4501 7275
rect 4537 5537 4549 7275
rect 4513 1889 4525 5475
rect 4537 1889 4549 5499
rect 4561 3689 4573 7275
rect 4585 5585 4597 7275
rect 4633 5609 4645 7275
rect 4657 5633 4669 7275
rect 4681 5681 4693 7275
rect 4729 5729 4741 7275
rect 4585 1889 4597 5547
rect 4657 1889 4669 3603
rect 4681 1889 4693 5643
rect 4729 1889 4741 5691
rect 4753 5105 4765 7275
rect 4849 5753 4861 7275
rect 4873 5777 4885 7275
rect 4897 3689 4909 7275
rect 4921 5801 4933 7275
rect 4969 5825 4981 7275
rect 4753 1889 4765 3123
rect 4801 1889 4813 3099
rect 4873 1889 4885 3075
rect 4969 1889 4981 5739
rect 4993 4889 5005 7275
rect 5017 5849 5029 7275
rect 5041 4889 5053 7275
rect 5065 4097 5077 7275
rect 5113 5873 5125 7275
rect 5137 4169 5149 7275
rect 5161 5897 5173 7275
rect 5209 4361 5221 7275
rect 4993 1889 5005 3051
rect 5017 1889 5029 3027
rect 5065 1889 5077 3699
rect 5089 1889 5101 3003
rect 5113 1889 5125 4083
rect 5233 2993 5245 7275
rect 5257 5921 5269 7275
rect 5329 5033 5341 7275
rect 5353 5369 5365 7275
rect 5401 5801 5413 7275
rect 5425 2969 5437 7275
rect 5497 5153 5509 7275
rect 5521 4865 5533 7275
rect 5545 5153 5557 7275
rect 5569 4145 5581 7275
rect 5617 3137 5629 7275
rect 5665 5537 5677 7275
rect 5737 5801 5749 7275
rect 5641 1889 5653 5307
rect 5785 4145 5797 7275
rect 5809 5945 5821 7275
rect 5833 5969 5845 7275
rect 5881 5993 5893 7275
rect 5929 6017 5941 7275
rect 5785 1889 5797 2979
rect 5833 1889 5845 2979
rect 5857 1889 5869 4779
rect 5881 1889 5893 5787
rect 5929 1889 5941 5787
rect 5953 1889 5965 5523
rect 5977 1889 5989 6027
rect 6001 4673 6013 7275
rect 6025 6065 6037 7275
rect 6049 4673 6061 7275
rect 6073 3593 6085 7275
rect 6025 1889 6037 2931
rect 6073 1889 6085 2907
rect 6097 2897 6109 7275
rect 6145 6089 6157 7275
rect 6169 2873 6181 7275
rect 6193 6137 6205 7275
rect 6193 1889 6205 6099
rect 6217 5633 6229 7275
rect 6241 3977 6253 7275
rect 6289 3977 6301 7275
rect 6313 6161 6325 7275
rect 6217 1889 6229 2835
rect 6241 1889 6253 2811
rect 6313 1889 6325 2787
rect 6337 2777 6349 7275
rect 6361 3953 6373 7275
rect 6385 2753 6397 4851
rect 6409 4385 6421 7275
rect 6433 6185 6445 7275
rect 6361 1889 6373 2739
rect 6433 1889 6445 5091
rect 6481 4865 6493 7275
rect 6529 4385 6541 7275
rect 6529 1889 6541 3939
rect 6553 3617 6565 7275
rect 6577 6209 6589 7275
rect 6601 6233 6613 7275
rect 6577 1889 6589 4875
rect 6649 2753 6661 7275
rect 6697 6257 6709 7275
rect 6721 6281 6733 7275
rect 6745 6305 6757 7275
rect 6793 6329 6805 7275
rect 6601 1889 6613 2739
rect 6649 1889 6661 2715
rect 6697 1889 6709 2739
rect 6793 1889 6805 4179
rect 6817 3209 6829 6315
rect 6841 3497 6853 7275
rect 6913 6329 6925 7275
rect 6817 1889 6829 2691
rect 6865 1889 6877 3603
rect 6889 1889 6901 3147
rect 6937 2705 6949 7275
rect 6961 6353 6973 7275
rect 6913 1889 6925 2667
rect 6985 1889 6997 4851
rect 7009 1889 7021 3507
rect 7033 2705 7045 7275
rect 7057 5873 7069 7275
rect 7081 6377 7093 7275
rect 7057 1889 7069 4587
rect 7105 3233 7117 7275
rect 7153 3473 7165 7275
rect 7177 5873 7189 7275
rect 7201 6401 7213 7275
rect 7249 5417 7261 7275
rect 7273 6425 7285 7275
rect 7297 6185 7309 7275
rect 7321 6329 7333 7275
rect 7369 6329 7381 7275
rect 7393 6449 7405 7275
rect 7105 1889 7117 2643
rect 7153 1889 7165 3219
rect 7225 1889 7237 2619
rect 7249 1889 7261 3267
rect 7321 1889 7333 3531
rect 7345 1889 7357 2595
rect 7369 1889 7381 5859
rect 7417 5609 7429 7275
rect 7465 5609 7477 7275
rect 7489 5225 7501 7275
rect 7513 4745 7525 7275
rect 7561 4745 7573 7275
rect 7585 6473 7597 7275
rect 7609 6521 7621 7275
rect 7633 6545 7645 7275
rect 7393 1889 7405 2667
rect 7465 1889 7477 3627
rect 7513 1889 7525 3003
rect 7585 1889 7597 2571
rect 7609 1889 7621 6483
rect 7681 4361 7693 7275
rect 7705 3929 7717 7275
rect 7729 6569 7741 7275
rect 7777 6425 7789 7275
rect 7633 1889 7645 2547
rect 7753 1889 7765 3915
rect 7801 3425 7813 7275
rect 7825 6593 7837 7275
rect 7873 6617 7885 7275
rect 7921 6257 7933 7275
rect 7945 6617 7957 7275
rect 7801 1889 7813 2523
rect 7825 1889 7837 3603
rect 7849 1889 7861 4659
rect 7873 2537 7885 5667
rect 7969 4913 7981 7275
rect 8017 4913 8029 7275
rect 8065 5681 8077 7275
rect 7897 1889 7909 4659
rect 7921 1889 7933 4611
rect 7945 1889 7957 2523
rect 7993 1889 8005 4179
rect 8017 1889 8029 4611
rect 8137 4265 8149 7275
rect 8161 5753 8173 7275
rect 8185 5825 8197 7275
rect 8209 2513 8221 6531
rect 8233 5825 8245 7275
rect 8257 2681 8269 7275
rect 8305 6545 8317 7275
rect 8353 2513 8365 7275
rect 8377 5033 8389 7275
rect 8401 6641 8413 7275
rect 8449 4217 8461 7275
rect 8161 1889 8173 2499
rect 8473 2489 8485 7275
rect 8497 4217 8509 7275
rect 8521 2465 8533 7275
rect 8569 2609 8581 7275
rect 8593 2729 8605 7275
rect 8617 2657 8629 7275
rect 8665 3233 8677 7275
rect 8689 6425 8701 7275
rect 8713 5225 8725 7275
rect 8737 6665 8749 7275
rect 8785 6689 8797 7275
rect 8713 1889 8725 3219
rect 8737 1889 8749 2427
rect 8785 1889 8797 5835
rect 8809 5537 8821 7275
rect 8857 3233 8869 7275
rect 8905 3209 8917 7275
rect 8929 3233 8941 7275
rect 8953 6713 8965 7275
rect 9001 3497 9013 7275
rect 9025 3065 9037 7275
rect 9073 3497 9085 7275
rect 9121 5345 9133 7275
rect 9145 6737 9157 7275
rect 9169 6761 9181 7275
rect 8833 1889 8845 2403
rect 8857 1889 8869 2715
rect 8953 1889 8965 2379
rect 9145 1889 9157 2355
rect 9169 1889 9181 3771
rect 9217 2633 9229 7275
rect 9241 5753 9253 7275
rect 9265 2489 9277 7275
rect 9313 2633 9325 7275
rect 9193 1889 9205 2475
rect 9337 2345 9349 7275
rect 9361 4337 9373 7275
rect 9409 3665 9421 7275
rect 9433 5777 9445 7275
rect 9361 1889 9373 2307
rect 9385 1889 9397 3315
rect 9445 2321 9457 5715
rect 9481 4337 9493 7275
rect 9409 1889 9421 2283
rect 9505 1889 9517 6507
rect 9529 3761 9541 7275
rect 9553 4481 9565 7275
rect 9577 6521 9589 7275
rect 9625 5609 9637 7275
rect 9649 6785 9661 7275
rect 9553 1889 9565 2307
rect 9577 1889 9589 5307
rect 9649 1889 9661 5307
rect 9673 2681 9685 6771
rect 9697 5321 9709 7275
rect 9745 4625 9757 7275
rect 9769 4121 9781 7275
rect 9817 6809 9829 7275
rect 9721 1889 9733 3099
rect 9793 1889 9805 6771
rect 9865 4313 9877 7275
rect 9865 1889 9877 2259
rect 9889 2249 9901 7275
rect 9913 5849 9925 7275
rect 9937 5057 9949 7275
rect 10009 6305 10021 7275
rect 10033 6809 10045 7275
rect 9889 1889 9901 2211
rect 9961 1889 9973 4299
rect 10033 1889 10045 3099
rect 10081 2705 10093 7275
rect 10129 6809 10141 7275
rect 10105 1889 10117 5835
rect 10153 3545 10165 7275
rect 10177 6833 10189 7275
rect 10225 2609 10237 7275
rect 10249 4121 10261 7275
rect 10297 6857 10309 7275
rect 10345 6593 10357 7275
rect 10225 1889 10237 2595
rect 10297 1889 10309 6579
rect 10369 2681 10381 7275
rect 10417 3569 10429 7275
rect 10321 1889 10333 2595
rect 10417 1889 10429 2451
rect 10441 1889 10453 6363
rect 10465 2633 10477 7275
rect 10489 6617 10501 7275
rect 10513 6881 10525 7275
rect 10561 4985 10573 7275
rect 10609 4673 10621 7275
rect 10681 6761 10693 7275
rect 10513 1889 10525 3603
rect 10537 1889 10549 3771
rect 10561 1889 10573 3195
rect 10633 1889 10645 6147
rect 10681 1889 10693 2451
rect 10705 2201 10717 7275
rect 10729 5561 10741 7275
rect 10753 6761 10765 7275
rect 10777 5561 10789 7275
rect 10825 5105 10837 7275
rect 10849 3929 10861 7275
rect 10873 5585 10885 7275
rect 10897 6905 10909 7275
rect 10945 6569 10957 7275
rect 10849 1889 10861 2163
rect 10897 1889 10909 3939
rect 10969 2153 10981 7275
rect 10993 6569 11005 7275
rect 11017 6929 11029 7275
rect 11065 6953 11077 7275
rect 11017 1889 11029 2115
rect 11065 1889 11077 2331
rect 11089 2105 11101 7275
rect 11113 5657 11125 7275
rect 11137 6521 11149 7275
rect 11161 5993 11173 7275
rect 11161 1889 11173 2331
rect 11185 1889 11197 5643
rect 11209 2345 11221 6603
rect 11257 5993 11269 7275
rect 11233 1889 11245 5091
rect 11257 1889 11269 2331
rect 11281 1889 11293 4851
rect 11305 1889 11317 5523
rect 11329 4841 11341 7275
rect 11353 6521 11365 7275
rect 11377 6977 11389 7275
rect 11425 7001 11437 7275
rect 11377 1889 11389 6267
rect 11425 1889 11437 6795
rect 11473 2081 11485 7275
rect 11545 7025 11557 7275
rect 11569 7049 11581 7275
rect 11497 1889 11509 3651
rect 11521 1889 11533 3747
rect 11545 1889 11557 5139
rect 11569 2321 11581 7011
rect 11593 4049 11605 7275
rect 11641 5153 11653 7275
rect 11593 1889 11605 2043
rect 11617 1889 11629 5115
rect 11665 3785 11677 7275
rect 11713 2441 11725 7275
rect 11761 5129 11773 7275
rect 11785 3617 11797 7275
rect 11809 5705 11821 7275
rect 11857 4385 11869 7275
rect 11881 5753 11893 7275
rect 11905 3905 11917 7275
rect 11953 5705 11965 7275
rect 12001 7025 12013 7275
rect 12073 7073 12085 7275
rect 12097 5753 12109 7275
rect 12145 4697 12157 7275
rect 11713 1889 11725 2019
rect 11737 1889 11749 3003
rect 11953 1889 11965 4035
rect 11977 1889 11989 2643
rect 12001 1889 12013 3891
rect 12073 1889 12085 3459
rect 12097 1889 12109 3939
rect 12193 3665 12205 7275
rect 12217 5105 12229 7275
rect 12265 7097 12277 7275
rect 12145 1889 12157 3051
rect 12169 1889 12181 3411
rect 12241 2441 12253 5379
rect 12313 3209 12325 7275
rect 12337 4169 12349 7275
rect 12361 7121 12373 7275
rect 12193 1889 12205 2427
rect 12337 1889 12349 2427
rect 12361 1889 12373 6411
rect 12385 1889 12397 3675
rect 12409 2441 12421 7275
rect 12433 3761 12445 7275
rect 12457 4169 12469 7275
rect 12481 6185 12493 7275
rect 12505 7145 12517 7275
rect 12457 1889 12469 3051
rect 12481 1889 12493 4107
rect 12505 1889 12517 6243
rect 12553 3329 12565 7275
rect 12577 5033 12589 7275
rect 12601 7169 12613 7275
rect 12553 1889 12565 1995
rect 12601 1985 12613 6075
rect 12649 4121 12661 7275
rect 12577 1889 12589 1971
rect 12673 1889 12685 3123
rect 12697 2441 12709 7275
rect 12769 5465 12781 7275
rect 12817 5465 12829 7275
rect 12889 4385 12901 7275
rect 12913 5273 12925 7275
rect 12937 7193 12949 7275
rect 12769 1889 12781 4347
rect 12889 1889 12901 1971
rect 12913 1889 12925 2067
rect 12937 1889 12949 3435
rect 12961 1985 12973 5187
rect 12985 3449 12997 7275
rect 13009 6713 13021 7275
rect 13033 4577 13045 7275
rect 13033 1889 13045 2067
rect 13057 1889 13069 6075
rect 13081 4361 13093 7275
rect 13105 6713 13117 7275
rect 13129 7217 13141 7275
rect 13177 6857 13189 7275
rect 13201 6713 13213 7275
rect 13081 1889 13093 1971
rect 13129 1889 13141 6699
rect 13249 6209 13261 7275
rect 13177 1889 13189 5763
rect 13201 1889 13213 3747
rect 13225 1889 13237 4563
rect 13273 1889 13285 6171
rect 13297 3473 13309 7275
rect 13321 4865 13333 7275
rect 13369 6857 13381 7275
rect 13345 3065 13357 6699
rect 13417 6449 13429 7275
rect 13297 1889 13309 2667
rect 13321 1889 13333 1947
rect 13369 1889 13381 5211
rect 13441 4721 13453 7275
rect 13465 6713 13477 7275
rect 13513 5945 13525 7275
rect 13393 1889 13405 3891
rect 13417 1889 13429 1923
rect 13465 1889 13477 4851
rect 13489 1889 13501 5931
rect 13537 4121 13549 7275
rect 13561 3137 13573 7275
rect 13609 7241 13621 7275
rect 13561 1889 13573 1899
rect 13585 1889 13597 4707
rect 13609 1889 13621 6939
rect 13633 5753 13645 7275
rect 13657 1889 13669 4107
rect 13681 3713 13693 7275
rect 13729 6041 13741 7275
rect 13681 1889 13693 3411
rect 13705 1889 13717 3387
rect 13753 3041 13765 7275
rect 13777 4289 13789 7275
rect 13777 1889 13789 3387
rect 13801 1913 13813 5859
rect 13825 4817 13837 7275
rect 13825 1889 13837 4539
rect 13849 3425 13861 7275
rect 13897 6953 13909 7275
rect 13873 1889 13885 4851
rect 13897 1889 13909 6723
rect 13921 3401 13933 6531
rect 13945 3017 13957 7275
rect 13969 5945 13981 7275
rect 13993 6041 14005 7275
rect 13969 1889 13981 3195
rect 13993 1889 14005 5859
rect 14017 1889 14029 6075
rect 14041 5249 14053 7275
rect 14065 6545 14077 7275
rect 14065 1889 14077 6219
rect 14089 4961 14101 7275
rect 14137 4385 14149 7275
rect 14089 1889 14101 4275
rect 14113 1889 14125 3387
rect 14161 3233 14173 7275
rect 14185 3449 14197 6027
rect 14209 5249 14221 7275
rect 14257 7265 14269 7275
rect 14209 1889 14221 5211
rect 14233 1889 14245 5187
rect 14257 1889 14269 6723
rect 14281 4121 14293 7275
rect 14305 4961 14317 7275
rect 14425 6929 14437 7275
rect 14281 1889 14293 3435
rect 14329 1889 14341 6243
rect 14353 1889 14365 3267
rect 14377 1889 14389 3075
rect 14401 2297 14413 6531
rect 14425 1889 14437 3123
rect 14449 1889 14461 4395
rect 14473 2369 14485 7251
rect 14497 3137 14509 7155
rect 14833 5297 14845 7275
rect 14977 6041 14989 7275
rect 15001 5801 15013 7275
rect 15049 5513 15061 7275
rect 15097 5513 15109 7275
rect 15121 4601 15133 7275
rect 15145 6089 15157 7275
rect 15169 6545 15181 7275
rect 14953 1889 14965 3123
rect 15145 1889 15157 3915
rect 15169 1889 15181 5571
rect 15193 1889 15205 6315
rect 15217 3233 15229 6075
rect 15241 1889 15253 4587
rect 15265 1889 15277 4659
rect 15289 1985 15301 7275
rect 15313 1889 15325 5115
rect 15361 1889 15373 4587
rect 15385 1889 15397 5019
rect 15409 1889 15421 3915
rect 15457 1889 15469 2283
rect 15481 1889 15493 6867
rect 15553 1889 15565 5355
rect 15649 4385 15661 7275
rect 15697 5873 15709 7275
rect 15841 7193 15853 7275
rect 15865 3473 15877 7275
rect 15889 5585 15901 7275
rect 15913 4697 15925 7275
rect 15601 1889 15613 2019
rect 15673 1889 15685 3027
rect 15721 1889 15733 3219
rect 15937 2321 15949 7275
rect 15985 6809 15997 7275
rect 15961 1889 15973 4491
rect 16009 2273 16021 7275
rect 16033 4697 16045 7275
rect 16057 6353 16069 7275
rect 16105 7169 16117 7275
rect 16129 5633 16141 7275
rect 16153 4697 16165 7275
rect 16033 1889 16045 3267
rect 16057 1889 16069 4107
rect 16081 2441 16093 4683
rect 16105 1889 16117 4491
rect 16177 4385 16189 7275
rect 16201 6089 16213 7275
rect 16249 6329 16261 7275
rect 16153 1889 16165 1971
rect 16201 1889 16213 4803
rect 16225 1985 16237 6075
rect 16273 3449 16285 7275
rect 16297 4097 16309 7275
rect 16321 4913 16333 7275
rect 16369 6425 16381 7275
rect 16393 6185 16405 7275
rect 16417 7169 16429 7275
rect 16297 1889 16309 2619
rect 16369 1889 16381 4251
rect 16417 1889 16429 7011
rect 16513 4793 16525 7275
rect 16441 1889 16453 3603
rect 16513 1889 16525 4083
rect 16537 1889 16549 3939
rect 16585 3497 16597 7275
rect 16609 4913 16621 7275
rect 16633 6089 16645 7275
rect 16681 6353 16693 7275
rect 16561 1889 16573 3435
rect 16609 1889 16621 3987
rect 16657 1889 16669 2619
rect 16681 1889 16693 3987
rect 16705 3305 16717 7275
rect 16729 4289 16741 7275
rect 16753 4097 16765 6531
rect 16777 5897 16789 7275
rect 16825 6449 16837 7275
rect 16777 1889 16789 4779
rect 16801 1889 16813 4731
rect 16837 2681 16849 4899
rect 16897 4745 16909 7275
rect 16921 4793 16933 7275
rect 16969 4913 16981 7275
rect 17017 6977 17029 7275
rect 17041 4169 17053 7275
rect 16873 1889 16885 2451
rect 17089 2057 17101 7275
rect 17137 6929 17149 7275
rect 17161 2489 17173 7275
rect 17209 6977 17221 7275
rect 17257 2753 17269 7275
rect 17281 7025 17293 7275
rect 17305 4049 17317 7275
rect 17353 4385 17365 7275
rect 17377 5105 17389 7275
rect 17425 5777 17437 7275
rect 17425 1889 17437 4275
rect 17473 2825 17485 7275
rect 17545 2297 17557 7275
rect 17593 4361 17605 7275
rect 17569 1889 17581 2715
rect 17593 1889 17605 4083
rect 17617 1889 17629 7011
rect 17641 4025 17653 7275
rect 17665 4097 17677 7035
rect 17689 7025 17701 7275
rect 17641 1889 17653 2187
rect 17689 1889 17701 4611
rect 17713 3329 17725 7275
rect 17713 1889 17725 2811
rect 17737 1889 17749 3291
rect 17761 2801 17773 7275
rect 17785 2825 17797 6363
rect 17809 2801 17821 7275
rect 17833 3641 17845 7275
rect 17857 7193 17869 7275
rect 17833 1889 17845 3291
rect 17857 1889 17869 4347
rect 17881 3305 17893 5883
rect 17905 5345 17917 7275
rect 17905 1889 17917 4371
rect 17929 2657 17941 7275
rect 17977 5489 17989 7275
rect 18025 6785 18037 7275
rect 18049 5321 18061 7275
rect 18073 5345 18085 7275
rect 17929 1889 17941 2475
rect 17953 1889 17965 2667
rect 17989 2489 18001 3483
rect 18025 1889 18037 2667
rect 18073 1889 18085 5211
rect 18121 4553 18133 7275
rect 18145 1889 18157 6843
rect 18169 5489 18181 7275
rect 18313 7265 18325 7275
rect 18169 1889 18181 3219
rect 18193 1889 18205 5811
rect 18241 1889 18253 3651
rect 18265 1889 18277 5235
rect 18313 1889 18325 7011
rect 18385 1889 18397 4611
rect 18433 1889 18445 7059
rect 18481 1889 18493 4419
rect 18505 1889 18517 3315
rect 18577 1889 18589 5211
rect 18721 4313 18733 7275
rect 18649 1889 18661 2403
rect 18697 1889 18709 3579
rect 18745 1889 18757 5499
rect 18865 3953 18877 7275
rect 18913 5609 18925 7275
rect 18817 1889 18829 2835
rect 18841 1889 18853 3027
rect 18937 1889 18949 6795
rect 18961 1889 18973 6411
rect 18985 5201 18997 7275
rect 19009 5009 19021 7275
rect 18985 1889 18997 2427
rect 19009 1889 19021 4779
rect 19033 3449 19045 7275
rect 19057 1889 19069 6723
rect 19081 5249 19093 7275
rect 19081 1889 19093 5211
rect 19105 4193 19117 7275
rect 19129 5441 19141 7275
rect 19105 1889 19117 3459
rect 19153 1889 19165 4539
rect 19177 3905 19189 7275
rect 19225 5177 19237 7275
rect 19201 1889 19213 3603
rect 19225 1889 19237 5115
rect 19249 1889 19261 5931
rect 19297 4121 19309 7275
rect 19321 6425 19333 7275
rect 19345 6185 19357 7275
rect 19345 1889 19357 4947
rect 19369 4529 19381 7275
rect 19417 5561 19429 7275
rect 19441 4697 19453 7275
rect 19465 4961 19477 7275
rect 19513 6617 19525 7275
rect 19393 1889 19405 4683
rect 19465 1889 19477 4875
rect 19489 2993 19501 4947
rect 19537 1889 19549 7203
rect 19561 6377 19573 7275
rect 19633 7049 19645 7275
rect 19585 1889 19597 5331
rect 19657 1889 19669 7107
rect 19681 1889 19693 6699
rect 19705 3113 19717 7275
rect 19729 1889 19741 5619
rect 19777 4793 19789 7275
rect 19849 6905 19861 7275
rect 19873 6449 19885 7275
rect 19801 1889 19813 4755
rect 19897 2081 19909 7275
rect 19945 4481 19957 7275
rect 19969 1889 19981 5979
rect 19993 3065 20005 7275
rect 20065 2033 20077 7275
rect 20089 3209 20101 7275
rect 20113 5057 20125 7275
rect 20161 3185 20173 7275
rect 20209 2009 20221 7275
rect 20281 4553 20293 7275
rect 20305 3929 20317 7275
rect 20329 6689 20341 7275
rect 20377 3425 20389 7275
rect 20401 4961 20413 7275
rect 20425 4481 20437 7275
rect 20449 4745 20461 7275
rect 20521 5033 20533 7275
rect 20521 1889 20533 4539
rect 20545 4385 20557 7275
rect 20593 4169 20605 7275
rect 20617 6353 20629 7275
rect 20641 1889 20653 3171
rect 20665 1889 20677 5091
rect 20689 3785 20701 7275
rect 20713 5033 20725 7275
rect 20737 3641 20749 7275
rect 20785 4337 20797 7275
rect 20833 4745 20845 7275
rect 20761 1889 20773 3603
rect 20833 1889 20845 3699
rect 20869 2513 20881 4731
rect 20905 4697 20917 7275
rect 20929 4745 20941 7275
rect 20857 1889 20869 2331
rect 20929 1889 20941 2955
rect 20953 2945 20965 7275
rect 21001 7241 21013 7275
rect 21025 5009 21037 7275
rect 21049 5057 21061 7275
rect 20977 1889 20989 4515
rect 21049 1889 21061 4659
rect 21097 4433 21109 7275
rect 21073 1889 21085 4251
rect 21097 1889 21109 4323
rect 21121 1937 21133 4731
rect 21145 3665 21157 7275
rect 21169 2465 21181 5043
rect 21193 4337 21205 5523
rect 21217 3569 21229 7275
rect 21241 4121 21253 7275
rect 21265 6113 21277 7275
rect 21313 6785 21325 7275
rect 21337 7241 21349 7275
rect 21217 1889 21229 3483
rect 21289 1889 21301 4659
rect 21313 1889 21325 6723
rect 21361 5057 21373 7275
rect 21385 5705 21397 7275
rect 21361 1889 21373 4803
rect 21409 1889 21421 6267
rect 21433 4601 21445 7275
rect 21457 6785 21469 7275
rect 21433 1889 21445 4419
rect 21457 1889 21469 4467
rect 21481 1889 21493 3795
rect 21505 3161 21517 7275
rect 21529 1889 21541 6003
rect 21553 5129 21565 7275
rect 21553 1889 21565 4827
rect 21577 4601 21589 7275
rect 21625 6065 21637 7275
rect 21601 1889 21613 4323
rect 21649 1889 21661 6963
rect 21673 4265 21685 7275
rect 21697 6377 21709 7275
rect 21673 1889 21685 3243
rect 21721 2609 21733 7275
rect 21745 3497 21757 7179
rect 21769 5393 21781 7275
rect 21793 6281 21805 7275
rect 21793 1889 21805 2331
rect 21817 2225 21829 7275
rect 21841 5009 21853 6771
rect 21865 4169 21877 7275
rect 21889 5105 21901 7275
rect 21865 1889 21877 4083
rect 21913 1889 21925 5931
rect 21937 3521 21949 7275
rect 21985 6881 21997 7275
rect 22033 6425 22045 7275
rect 21961 1961 21973 5043
rect 22045 4433 22057 6411
rect 22069 4577 22081 5115
rect 22105 4745 22117 7275
rect 22129 6641 22141 7275
rect 21985 1889 21997 2619
rect 22009 1889 22021 4179
rect 22105 1889 22117 4563
rect 22153 4241 22165 7275
rect 22201 4697 22213 7275
rect 22225 4673 22237 7275
rect 22177 1889 22189 2355
rect 22201 1889 22213 3531
rect 22249 2585 22261 7275
rect 22297 7145 22309 7275
rect 22273 1889 22285 4779
rect 22297 1889 22309 5307
rect 22321 4793 22333 7275
rect 22345 4817 22357 7275
rect 22321 1889 22333 3867
rect 22369 1889 22381 6411
rect 22393 4841 22405 7275
rect 22393 1889 22405 4611
rect 22417 4097 22429 5259
rect 22441 3401 22453 7275
rect 22465 3593 22477 4779
rect 22441 1889 22453 3291
rect 22489 1889 22501 3291
rect 22513 1889 22525 3531
rect 22537 1889 22549 6315
rect 22561 2177 22573 4827
rect 22585 4073 22597 7275
rect 22609 3305 22621 5235
rect 22657 1889 22669 2235
rect 22705 1889 22717 7083
rect 22945 6041 22957 7275
rect 22993 7049 23005 7275
rect 22729 1889 22741 3003
rect 22753 1889 22765 2763
rect 22801 1889 22813 3603
rect 22825 1889 22837 5139
rect 22849 1889 22861 5211
rect 22945 1889 22957 3507
rect 22993 1889 23005 5139
rect 23041 1889 23053 3315
rect 23065 1889 23077 4155
rect 23089 1889 23101 5619
rect 23137 5105 23149 7275
rect 23161 5873 23173 7275
rect 23161 1889 23173 4419
rect 23185 4409 23197 7275
rect 23209 4601 23221 7275
rect 23257 5345 23269 7275
rect 23233 1889 23245 2307
rect 23257 1889 23269 5283
rect 23305 4001 23317 7275
rect 23281 1889 23293 2139
rect 23329 1889 23341 2931
rect 23353 1889 23365 5451
rect 23377 3617 23389 7275
rect 23401 3689 23413 7275
rect 23425 4217 23437 7275
rect 23449 4433 23461 6819
rect 23473 5129 23485 7275
rect 23521 6521 23533 7275
rect 23593 6233 23605 7275
rect 23617 6089 23629 7275
rect 23401 1889 23413 3627
rect 23473 1889 23485 5067
rect 23497 2705 23509 5331
rect 23533 3641 23545 5691
rect 23557 3089 23569 5115
rect 23521 1889 23533 2331
rect 23617 1889 23629 5091
rect 23641 4337 23653 7275
rect 23665 5081 23677 7275
rect 23737 6665 23749 7275
rect 23761 7169 23773 7275
rect 23689 1889 23701 2715
rect 23761 1889 23773 6723
rect 23785 4961 23797 7275
rect 23833 6881 23845 7275
rect 23857 6833 23869 7275
rect 23809 1889 23821 3675
rect 23833 1889 23845 3411
rect 23857 1889 23869 6267
rect 23905 4697 23917 7275
rect 23905 1889 23917 3531
rect 23929 1889 23941 6363
rect 23953 2417 23965 7275
rect 23977 2729 23989 7275
rect 24001 4985 24013 7275
rect 24025 1889 24037 7083
rect 24049 3521 24061 7275
rect 24073 4385 24085 7275
rect 24121 7241 24133 7275
rect 24097 3497 24109 5499
rect 24049 1889 24061 3483
rect 24145 1889 24157 6939
rect 24169 3233 24181 7275
rect 24193 6857 24205 7275
rect 24217 2681 24229 7275
rect 24241 6497 24253 7275
rect 24289 3185 24301 7275
rect 24313 5873 24325 7275
rect 24337 5729 24349 7275
rect 24265 1889 24277 2571
rect 24313 1889 24325 4587
rect 24385 2393 24397 7275
rect 24409 3545 24421 7275
rect 24433 4937 24445 7275
rect 24385 1889 24397 2283
rect 24409 1889 24421 3507
rect 24457 2297 24469 6507
rect 24505 5321 24517 7275
rect 24529 6569 24541 7275
rect 24505 1889 24517 3339
rect 24529 1889 24541 3003
rect 24553 1889 24565 6147
rect 24577 4121 24589 7275
rect 24601 4481 24613 7275
rect 24649 3545 24661 7275
rect 24697 5417 24709 7275
rect 24721 4505 24733 7275
rect 24769 5825 24781 7275
rect 24817 6425 24829 7275
rect 24601 1889 24613 3171
rect 24625 1889 24637 3315
rect 24697 1889 24709 2427
rect 24721 1889 24733 3267
rect 24769 1889 24781 5739
rect 24793 2129 24805 5811
rect 24817 1889 24829 6387
rect 24841 4289 24853 7275
rect 24865 6473 24877 7275
rect 24877 3137 24889 6411
rect 24913 4049 24925 7275
rect 24937 5225 24949 7275
rect 24961 6761 24973 7275
rect 25009 5849 25021 7275
rect 25033 5321 25045 7275
rect 25057 4793 25069 7275
rect 25105 6257 25117 7275
rect 24865 1889 24877 2619
rect 24937 1889 24949 4491
rect 25009 1889 25021 2859
rect 25057 1889 25069 4035
rect 25081 1889 25093 5211
rect 25129 1889 25141 5787
rect 25153 4193 25165 7275
rect 25225 4841 25237 7275
rect 25249 4265 25261 7275
rect 25273 4625 25285 7275
rect 25297 6593 25309 7275
rect 25177 1889 25189 2019
rect 25201 1889 25213 2331
rect 25225 1889 25237 3963
rect 25273 1889 25285 2259
rect 25297 1889 25309 6291
rect 25345 3857 25357 7275
rect 25369 5105 25381 7275
rect 25321 1889 25333 3819
rect 25369 1889 25381 2427
rect 25393 1889 25405 6363
rect 25417 3353 25429 7275
rect 25465 5993 25477 7275
rect 25441 3905 25453 4827
rect 25417 1889 25429 3315
rect 25465 1889 25477 5931
rect 25489 4481 25501 7275
rect 25513 4505 25525 7275
rect 25561 7097 25573 7275
rect 25585 5033 25597 7275
rect 25609 6017 25621 7275
rect 25489 1889 25501 2427
rect 25537 1889 25549 4995
rect 25609 1889 25621 5931
rect 25633 1889 25645 4635
rect 25657 4409 25669 7275
rect 25681 6185 25693 7275
rect 25681 1889 25693 3723
rect 25705 1889 25717 5235
rect 25729 2369 25741 7275
rect 25777 6401 25789 7275
rect 25801 6617 25813 7275
rect 25753 4817 25765 5979
rect 25801 1889 25813 4491
rect 25825 1889 25837 5667
rect 25849 2273 25861 7275
rect 25849 1889 25861 2235
rect 25873 1889 25885 6531
rect 25897 5921 25909 7275
rect 25921 4625 25933 7275
rect 25945 4793 25957 7275
rect 25969 7265 25981 7275
rect 25981 4553 25993 6003
rect 26017 5297 26029 7275
rect 25945 1889 25957 3603
rect 25969 1889 25981 3363
rect 26041 1889 26053 5763
rect 26065 1889 26077 4539
rect 26089 3113 26101 7275
rect 26113 4505 26125 6963
rect 26233 6737 26245 7275
rect 26137 1889 26149 5355
rect 26161 1889 26173 5019
rect 26197 2249 26209 4899
rect 26257 4865 26269 7275
rect 26281 6161 26293 7275
rect 26185 1889 26197 2091
rect 26281 1889 26293 6123
rect 26305 4145 26317 7275
rect 26329 2681 26341 6147
rect 26353 2321 26365 7275
rect 26377 4313 26389 7275
rect 26401 4625 26413 7275
rect 26449 7241 26461 7275
rect 26473 5513 26485 7275
rect 26497 2849 26509 7275
rect 26545 2033 26557 7275
rect 26569 5033 26581 7275
rect 26593 4889 26605 7275
rect 26641 2537 26653 7275
rect 26665 3329 26677 7275
rect 26689 4457 26701 7275
rect 26737 4601 26749 7275
rect 26785 6185 26797 7275
rect 26833 4601 26845 7275
rect 26785 1889 26797 4395
rect 26833 1889 26845 4155
rect 26857 3689 26869 4587
rect 26905 4361 26917 7275
rect 26929 3761 26941 7275
rect 26953 4745 26965 7275
rect 27001 4265 27013 7275
rect 27025 5945 27037 7275
rect 27073 5201 27085 7275
rect 27073 1889 27085 4587
rect 27121 4577 27133 7275
rect 27169 4553 27181 7275
rect 27241 5201 27253 7275
rect 27265 5801 27277 7275
rect 27289 6929 27301 7275
rect 27337 6209 27349 7275
rect 27385 4721 27397 7275
rect 27457 5969 27469 7275
rect 27481 5657 27493 7275
rect 27529 5585 27541 7275
rect 27193 1889 27205 2883
rect 27553 1889 27565 5019
rect 27577 3665 27589 7275
rect 27601 4625 27613 7275
rect 27625 4529 27637 7275
rect 27673 5801 27685 7275
rect 27697 4673 27709 7275
rect 27745 7001 27757 7275
rect 27601 1889 27613 3603
rect 27649 2345 27661 4611
rect 27745 1889 27757 2403
rect 27769 1889 27781 4683
rect 27793 1889 27805 2739
rect 27817 1889 27829 4755
rect 27841 1913 27853 4587
rect 27865 1937 27877 2907
rect 27961 1889 28161 7275
rect 28210 5476 28280 5488
rect 28210 2548 28280 2560
rect 28210 1924 28280 1936
rect 28210 1900 28280 1912
rect 0 155 70 167
rect 0 131 70 143
rect 0 107 70 119
rect 0 83 70 95
rect 145 0 345 1090
rect 361 0 373 1090
rect 385 0 397 1090
rect 409 0 421 1090
rect 433 0 445 1090
rect 1633 192 1645 1090
rect 1729 144 1741 1090
rect 1777 96 1789 1090
rect 2497 144 2509 1090
rect 2785 96 2797 1090
rect 2953 216 2965 1090
rect 3001 240 3013 1090
rect 3961 288 3973 1090
rect 4177 312 4189 1090
rect 4201 336 4213 1090
rect 4249 360 4261 1090
rect 4345 384 4357 1090
rect 4465 408 4477 1090
rect 4633 432 4645 1090
rect 4849 288 4861 1090
rect 4921 456 4933 1090
rect 5233 480 5245 1090
rect 3769 0 3781 250
rect 5785 72 5797 1090
rect 6145 528 6157 1090
rect 6169 552 6181 1090
rect 6289 576 6301 1090
rect 6409 600 6421 1090
rect 6481 576 6493 1090
rect 6553 624 6565 1090
rect 6769 648 6781 1090
rect 6937 672 6949 1090
rect 7273 696 7285 1090
rect 7417 720 7429 1090
rect 5953 0 5965 490
rect 7681 456 7693 1090
rect 7705 744 7717 1090
rect 8041 456 8053 1090
rect 8137 0 8149 754
rect 8569 288 8581 1090
rect 9025 792 9037 1090
rect 9073 312 9085 1090
rect 9241 312 9253 1090
rect 9265 96 9277 1090
rect 9289 816 9301 1090
rect 9313 96 9325 1090
rect 9457 840 9469 1090
rect 9481 864 9493 1090
rect 9601 888 9613 1090
rect 9913 912 9925 1090
rect 9961 48 9973 1090
rect 10177 48 10189 1090
rect 10345 696 10357 1090
rect 10369 648 10381 1090
rect 10465 648 10477 1090
rect 10609 816 10621 1090
rect 10657 696 10669 1090
rect 10705 264 10717 1090
rect 10753 720 10765 1090
rect 10777 264 10789 1090
rect 10801 648 10813 1090
rect 10825 720 10837 1090
rect 10921 648 10933 1090
rect 10945 96 10957 1090
rect 9974 34 9992 48
rect 9973 0 9985 34
rect 10357 0 10369 82
rect 10969 24 10981 1090
rect 11137 936 11149 1090
rect 11329 960 11341 1090
rect 11665 984 11677 1090
rect 11761 96 11773 1090
rect 11809 1008 11821 1090
rect 11833 912 11845 1090
rect 11857 1032 11869 1090
rect 11881 912 11893 1090
rect 11905 1056 11917 1090
rect 12049 600 12061 1090
rect 12241 240 12253 1090
rect 12265 96 12277 1090
rect 12289 240 12301 1090
rect 12409 1032 12421 1090
rect 12601 1032 12613 1090
rect 12649 1080 12661 1090
rect 12721 600 12733 1090
rect 12817 312 12829 1090
rect 12985 384 12997 1090
rect 13009 312 13021 1090
rect 13129 120 13141 1090
rect 13273 336 13285 1090
rect 13513 192 13525 1090
rect 13753 360 13765 1090
rect 13921 1080 13933 1090
rect 14137 1080 14149 1090
rect 14161 384 14173 1090
rect 14473 720 14485 1090
rect 14593 240 14605 1090
rect 14689 0 14701 346
rect 15001 216 15013 1090
rect 15505 720 15517 1090
rect 15793 240 15805 1090
rect 15841 696 15853 1090
rect 15913 1056 15925 1090
rect 16153 360 16165 1090
rect 16225 336 16237 1090
rect 16249 696 16261 1090
rect 16321 336 16333 1090
rect 16465 1056 16477 1090
rect 16585 96 16597 1090
rect 16705 528 16717 1090
rect 16753 288 16765 1090
rect 16849 144 16861 1090
rect 16897 528 16909 1090
rect 17017 840 17029 1090
rect 17377 864 17389 1090
rect 14713 0 14725 10
rect 16885 0 16897 58
rect 17617 48 17629 1090
rect 17785 864 17797 1090
rect 17809 360 17821 1090
rect 17977 264 17989 1090
rect 18361 288 18373 1090
rect 18529 360 18541 1090
rect 18601 48 18613 1090
rect 18889 792 18901 1090
rect 19057 0 19069 706
rect 19129 336 19141 1090
rect 19273 720 19285 1090
rect 19321 984 19333 1090
rect 19441 624 19453 1090
rect 19489 504 19501 1090
rect 19561 888 19573 1090
rect 19609 480 19621 1090
rect 19705 888 19717 1090
rect 19753 984 19765 1090
rect 19825 672 19837 1090
rect 19849 168 19861 1090
rect 20377 840 20389 1090
rect 20545 672 20557 1090
rect 20593 816 20605 1090
rect 20689 312 20701 1090
rect 20737 576 20749 1090
rect 20785 576 20797 1090
rect 20881 816 20893 1090
rect 20953 720 20965 1090
rect 21001 240 21013 1090
rect 21121 624 21133 1090
rect 21169 960 21181 1090
rect 21193 576 21205 1090
rect 21241 576 21253 1090
rect 21457 624 21469 1090
rect 21721 720 21733 1090
rect 21769 528 21781 1090
rect 21817 840 21829 1090
rect 22033 912 22045 1090
rect 22081 792 22093 1090
rect 22105 912 22117 1090
rect 22129 1008 22141 1090
rect 22225 1080 22237 1090
rect 22585 1056 22597 1090
rect 22609 816 22621 1090
rect 22873 552 22885 1090
rect 22921 600 22933 1090
rect 23137 456 23149 1090
rect 23185 936 23197 1090
rect 23377 720 23389 1090
rect 23425 552 23437 1090
rect 23593 1032 23605 1090
rect 23641 888 23653 1090
rect 21229 0 21241 34
rect 23401 0 23413 322
rect 23713 48 23725 1090
rect 23953 336 23965 1090
rect 23977 288 23989 1090
rect 24097 600 24109 1090
rect 24169 288 24181 1090
rect 24217 744 24229 1090
rect 24433 336 24445 1090
rect 24457 432 24469 1090
rect 24649 672 24661 1090
rect 24961 672 24973 1090
rect 25585 696 25597 1090
rect 25753 648 25765 1090
rect 25897 768 25909 1090
rect 25993 672 26005 1090
rect 26089 864 26101 1090
rect 25573 0 25585 586
rect 26233 384 26245 1090
rect 26425 984 26437 1090
rect 26977 408 26989 1090
rect 27001 840 27013 1090
rect 27025 720 27037 1090
rect 27049 96 27061 1090
rect 27961 0 28161 1090
rect 28210 899 28280 911
rect 28210 611 28280 623
rect 28210 563 28280 575
rect 28210 539 28280 551
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 145 0 1 7275
box 0 0 1464 799
use nand3 g9738
timestamp 1386234893
transform 1 0 1609 0 1 7275
box 0 0 120 799
use rowcrosser OpcodeCondIn_91_5_93_
timestamp 1386086759
transform 1 0 1729 0 1 7275
box 0 0 48 799
use nand2 g9544
timestamp 1386234792
transform 1 0 1777 0 1 7275
box 0 0 96 799
use nand2 g9509
timestamp 1386234792
transform 1 0 1873 0 1 7275
box 0 0 96 799
use nand3 g9758
timestamp 1386234893
transform 1 0 1969 0 1 7275
box 0 0 120 799
use nand2 g9539
timestamp 1386234792
transform 1 0 2089 0 1 7275
box 0 0 96 799
use nand3 g9429
timestamp 1386234893
transform 1 0 2185 0 1 7275
box 0 0 120 799
use nand4 g9535
timestamp 1386234936
transform 1 0 2305 0 1 7275
box 0 0 144 799
use nand2 g9527
timestamp 1386234792
transform 1 0 2449 0 1 7275
box 0 0 96 799
use nand2 g9452
timestamp 1386234792
transform 1 0 2545 0 1 7275
box 0 0 96 799
use nand3 g9597
timestamp 1386234893
transform 1 0 2641 0 1 7275
box 0 0 120 799
use nand3 g9463
timestamp 1386234893
transform 1 0 2761 0 1 7275
box 0 0 120 799
use nor2 g9497
timestamp 1386235306
transform 1 0 2881 0 1 7275
box 0 0 120 799
use and2 g9552
timestamp 1386234845
transform 1 0 3001 0 1 7275
box 0 0 120 799
use nand3 g9687
timestamp 1386234893
transform 1 0 3121 0 1 7275
box 0 0 120 799
use nand2 g9540
timestamp 1386234792
transform 1 0 3241 0 1 7275
box 0 0 96 799
use nand3 g9777
timestamp 1386234893
transform 1 0 3337 0 1 7275
box 0 0 120 799
use nand2 g9756
timestamp 1386234792
transform 1 0 3457 0 1 7275
box 0 0 96 799
use and2 g9521
timestamp 1386234845
transform 1 0 3553 0 1 7275
box 0 0 120 799
use nand2 g9493
timestamp 1386234792
transform 1 0 3673 0 1 7275
box 0 0 96 799
use nand3 g9736
timestamp 1386234893
transform 1 0 3769 0 1 7275
box 0 0 120 799
use nand2 g9747
timestamp 1386234792
transform 1 0 3889 0 1 7275
box 0 0 96 799
use xor2 g9741
timestamp 1386237344
transform 1 0 3985 0 1 7275
box 0 0 192 799
use nand2 g9763
timestamp 1386234792
transform 1 0 4177 0 1 7275
box 0 0 96 799
use inv g9479
timestamp 1386238110
transform 1 0 4273 0 1 7275
box 0 0 120 799
use nand3 g9605
timestamp 1386234893
transform 1 0 4393 0 1 7275
box 0 0 120 799
use nand2 g9446
timestamp 1386234792
transform 1 0 4513 0 1 7275
box 0 0 96 799
use nand2 g9613
timestamp 1386234792
transform 1 0 4609 0 1 7275
box 0 0 96 799
use nor2 g9633
timestamp 1386235306
transform 1 0 4705 0 1 7275
box 0 0 120 799
use nand3 g9425
timestamp 1386234893
transform 1 0 4825 0 1 7275
box 0 0 120 799
use nand4 g9786
timestamp 1386234936
transform 1 0 4945 0 1 7275
box 0 0 144 799
use nand2 g9469
timestamp 1386234792
transform 1 0 5089 0 1 7275
box 0 0 96 799
use nand2 g9555
timestamp 1386234792
transform 1 0 5185 0 1 7275
box 0 0 96 799
use mux2 g9474
timestamp 1386235218
transform 1 0 5281 0 1 7275
box 0 0 192 799
use nand3 g9674
timestamp 1386234893
transform 1 0 5473 0 1 7275
box 0 0 120 799
use inv g9626
timestamp 1386238110
transform 1 0 5593 0 1 7275
box 0 0 120 799
use rowcrosser OpcodeCondIn_91_7_93_
timestamp 1386086759
transform 1 0 5713 0 1 7275
box 0 0 48 799
use nand2 g9512
timestamp 1386234792
transform 1 0 5761 0 1 7275
box 0 0 96 799
use inv g9405
timestamp 1386238110
transform 1 0 5857 0 1 7275
box 0 0 120 799
use nand4 g9411
timestamp 1386234936
transform 1 0 5977 0 1 7275
box 0 0 144 799
use nand4 g9507
timestamp 1386234936
transform 1 0 6121 0 1 7275
box 0 0 144 799
use nand3 g9768
timestamp 1386234893
transform 1 0 6265 0 1 7275
box 0 0 120 799
use and2 g2
timestamp 1386234845
transform 1 0 6385 0 1 7275
box 0 0 120 799
use nand3 g9730
timestamp 1386234893
transform 1 0 6505 0 1 7275
box 0 0 120 799
use rowcrosser LrSel
timestamp 1386086759
transform 1 0 6625 0 1 7275
box 0 0 48 799
use nand2 g9774
timestamp 1386234792
transform 1 0 6673 0 1 7275
box 0 0 96 799
use inv g9431
timestamp 1386238110
transform 1 0 6769 0 1 7275
box 0 0 120 799
use nand3 g9594
timestamp 1386234893
transform 1 0 6889 0 1 7275
box 0 0 120 799
use nand3 g9672
timestamp 1386234893
transform 1 0 7009 0 1 7275
box 0 0 120 799
use nand2 g9528
timestamp 1386234792
transform 1 0 7129 0 1 7275
box 0 0 96 799
use nand3 g9462
timestamp 1386234893
transform 1 0 7225 0 1 7275
box 0 0 120 799
use nand2 g9522
timestamp 1386234792
transform 1 0 7345 0 1 7275
box 0 0 96 799
use nand2 g9500
timestamp 1386234792
transform 1 0 7441 0 1 7275
box 0 0 96 799
use nand3 g9471
timestamp 1386234893
transform 1 0 7537 0 1 7275
box 0 0 120 799
use nand2 g9578
timestamp 1386234792
transform 1 0 7657 0 1 7275
box 0 0 96 799
use nand2 g9727
timestamp 1386234792
transform 1 0 7753 0 1 7275
box 0 0 96 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 7849 0 1 7275
box 0 0 48 799
use nand2 g9475
timestamp 1386234792
transform 1 0 7897 0 1 7275
box 0 0 96 799
use inv g9583
timestamp 1386238110
transform 1 0 7993 0 1 7275
box 0 0 120 799
use nand2 g9562
timestamp 1386234792
transform 1 0 8113 0 1 7275
box 0 0 96 799
use nor2 g9644
timestamp 1386235306
transform 1 0 8209 0 1 7275
box 0 0 120 799
use nand2 g9632
timestamp 1386234792
transform 1 0 8329 0 1 7275
box 0 0 96 799
use nand3 g9755
timestamp 1386234893
transform 1 0 8425 0 1 7275
box 0 0 120 799
use nand2 g9549
timestamp 1386234792
transform 1 0 8545 0 1 7275
box 0 0 96 799
use nand3 g9492
timestamp 1386234893
transform 1 0 8641 0 1 7275
box 0 0 120 799
use and2 g9627
timestamp 1386234845
transform 1 0 8761 0 1 7275
box 0 0 120 799
use nand2 g9704
timestamp 1386234792
transform 1 0 8881 0 1 7275
box 0 0 96 799
use and2 g9694
timestamp 1386234845
transform 1 0 8977 0 1 7275
box 0 0 120 799
use nand2 g9635
timestamp 1386234792
transform 1 0 9097 0 1 7275
box 0 0 96 799
use nand2 g9607
timestamp 1386234792
transform 1 0 9193 0 1 7275
box 0 0 96 799
use nand2 g9701
timestamp 1386234792
transform 1 0 9289 0 1 7275
box 0 0 96 799
use nor2 g9784
timestamp 1386235306
transform 1 0 9385 0 1 7275
box 0 0 120 799
use nand2 g9530
timestamp 1386234792
transform 1 0 9505 0 1 7275
box 0 0 96 799
use and2 g9772
timestamp 1386234845
transform 1 0 9601 0 1 7275
box 0 0 120 799
use nor2 g9440
timestamp 1386235306
transform 1 0 9721 0 1 7275
box 0 0 120 799
use nand4 g9659
timestamp 1386234936
transform 1 0 9841 0 1 7275
box 0 0 144 799
use nor2 g9737
timestamp 1386235306
transform 1 0 9985 0 1 7275
box 0 0 120 799
use nand2 g9759
timestamp 1386234792
transform 1 0 10105 0 1 7275
box 0 0 96 799
use and2 g9502
timestamp 1386234845
transform 1 0 10201 0 1 7275
box 0 0 120 799
use nor2 g9622
timestamp 1386235306
transform 1 0 10321 0 1 7275
box 0 0 120 799
use nand2 g9717
timestamp 1386234792
transform 1 0 10441 0 1 7275
box 0 0 96 799
use inv g9556
timestamp 1386238110
transform 1 0 10537 0 1 7275
box 0 0 120 799
use nand4 g9458
timestamp 1386234936
transform 1 0 10657 0 1 7275
box 0 0 144 799
use nand3 g9422
timestamp 1386234893
transform 1 0 10801 0 1 7275
box 0 0 120 799
use nand3 g9513
timestamp 1386234893
transform 1 0 10921 0 1 7275
box 0 0 120 799
use nand4 g9805
timestamp 1386234936
transform 1 0 11041 0 1 7275
box 0 0 144 799
use inv g9525
timestamp 1386238110
transform 1 0 11185 0 1 7275
box 0 0 120 799
use nand2 g9682
timestamp 1386234792
transform 1 0 11305 0 1 7275
box 0 0 96 799
use inv g9441
timestamp 1386238110
transform 1 0 11401 0 1 7275
box 0 0 120 799
use nand2 g9518
timestamp 1386234792
transform 1 0 11521 0 1 7275
box 0 0 96 799
use and2 g9641
timestamp 1386234845
transform 1 0 11617 0 1 7275
box 0 0 120 799
use nand2 g9652
timestamp 1386234792
transform 1 0 11737 0 1 7275
box 0 0 96 799
use nand2 g9568
timestamp 1386234792
transform 1 0 11833 0 1 7275
box 0 0 96 799
use inv g9588
timestamp 1386238110
transform 1 0 11929 0 1 7275
box 0 0 120 799
use nor2 g9715
timestamp 1386235306
transform 1 0 12049 0 1 7275
box 0 0 120 799
use and2 g9724
timestamp 1386234845
transform 1 0 12169 0 1 7275
box 0 0 120 799
use nand2 g9686
timestamp 1386234792
transform 1 0 12289 0 1 7275
box 0 0 96 799
use nand4 g9778
timestamp 1386234936
transform 1 0 12385 0 1 7275
box 0 0 144 799
use nand2 g9795
timestamp 1386234792
transform 1 0 12529 0 1 7275
box 0 0 96 799
use inv g9478
timestamp 1386238110
transform 1 0 12625 0 1 7275
box 0 0 120 799
use inv g9655
timestamp 1386238110
transform 1 0 12745 0 1 7275
box 0 0 120 799
use nand2 g9584
timestamp 1386234792
transform 1 0 12865 0 1 7275
box 0 0 96 799
use nand2 g9470
timestamp 1386234792
transform 1 0 12961 0 1 7275
box 0 0 96 799
use nand2 g9712
timestamp 1386234792
transform 1 0 13057 0 1 7275
box 0 0 96 799
use nor2 g9679
timestamp 1386235306
transform 1 0 13153 0 1 7275
box 0 0 120 799
use and2 g9487
timestamp 1386234845
transform 1 0 13273 0 1 7275
box 0 0 120 799
use nand2 g9675
timestamp 1386234792
transform 1 0 13393 0 1 7275
box 0 0 96 799
use nand2 g9669
timestamp 1386234792
transform 1 0 13489 0 1 7275
box 0 0 96 799
use and2 g9572
timestamp 1386234845
transform 1 0 13585 0 1 7275
box 0 0 120 799
use nand2 g9600
timestamp 1386234792
transform 1 0 13705 0 1 7275
box 0 0 96 799
use nor2 g9673
timestamp 1386235306
transform 1 0 13801 0 1 7275
box 0 0 120 799
use nand2 g9447
timestamp 1386234792
transform 1 0 13921 0 1 7275
box 0 0 96 799
use nand2 g9606
timestamp 1386234792
transform 1 0 14017 0 1 7275
box 0 0 96 799
use and2 g9719
timestamp 1386234845
transform 1 0 14113 0 1 7275
box 0 0 120 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 14233 0 1 7275
box 0 0 96 799
use scandtype g9643
timestamp 1386241841
transform 1 0 14329 0 1 7275
box 0 0 624 799
use and2 g9595
timestamp 1386234845
transform 1 0 14953 0 1 7275
box 0 0 120 799
use nand3 stateSub_reg_91_2_93_
timestamp 1386234893
transform 1 0 15073 0 1 7275
box 0 0 120 799
use scandtype g9464
timestamp 1386241841
transform 1 0 15193 0 1 7275
box 0 0 624 799
use nand4 g9545
timestamp 1386234936
transform 1 0 15817 0 1 7275
box 0 0 144 799
use nand3 g9410
timestamp 1386234893
transform 1 0 15961 0 1 7275
box 0 0 120 799
use nand4 g9476
timestamp 1386234936
transform 1 0 16081 0 1 7275
box 0 0 144 799
use nand3 g9579
timestamp 1386234893
transform 1 0 16225 0 1 7275
box 0 0 120 799
use nand2 g9612
timestamp 1386234792
transform 1 0 16345 0 1 7275
box 0 0 96 799
use inv g9690
timestamp 1386238110
transform 1 0 16441 0 1 7275
box 0 0 120 799
use nand2 g9653
timestamp 1386234792
transform 1 0 16561 0 1 7275
box 0 0 96 799
use nand2 g9785
timestamp 1386234792
transform 1 0 16657 0 1 7275
box 0 0 96 799
use inv g9427
timestamp 1386238110
transform 1 0 16753 0 1 7275
box 0 0 120 799
use and2 g9499
timestamp 1386234845
transform 1 0 16873 0 1 7275
box 0 0 120 799
use and2 g9494
timestamp 1386234845
transform 1 0 16993 0 1 7275
box 0 0 120 799
use and2 g9753
timestamp 1386234845
transform 1 0 17113 0 1 7275
box 0 0 120 799
use nand2 g9762
timestamp 1386234792
transform 1 0 17233 0 1 7275
box 0 0 96 799
use and2 g9416
timestamp 1386234845
transform 1 0 17329 0 1 7275
box 0 0 120 799
use nor2 g9468
timestamp 1386235306
transform 1 0 17449 0 1 7275
box 0 0 120 799
use nand2 g9520
timestamp 1386234792
transform 1 0 17569 0 1 7275
box 0 0 96 799
use nor2 g9486
timestamp 1386235306
transform 1 0 17665 0 1 7275
box 0 0 120 799
use nand2 g9666
timestamp 1386234792
transform 1 0 17785 0 1 7275
box 0 0 96 799
use nor2 g9438
timestamp 1386235306
transform 1 0 17881 0 1 7275
box 0 0 120 799
use nand2 g9515
timestamp 1386234792
transform 1 0 18001 0 1 7275
box 0 0 96 799
use inv StatusReg_reg_91_1_93_
timestamp 1386238110
transform 1 0 18097 0 1 7275
box 0 0 120 799
use scandtype g9575
timestamp 1386241841
transform 1 0 18217 0 1 7275
box 0 0 624 799
use inv g9534
timestamp 1386238110
transform 1 0 18841 0 1 7275
box 0 0 120 799
use nand2 g9538
timestamp 1386234792
transform 1 0 18961 0 1 7275
box 0 0 96 799
use nand2 g9731
timestamp 1386234792
transform 1 0 19057 0 1 7275
box 0 0 96 799
use inv g9524
timestamp 1386238110
transform 1 0 19153 0 1 7275
box 0 0 120 799
use nand3 g9489
timestamp 1386234893
transform 1 0 19273 0 1 7275
box 0 0 120 799
use nand2 g9803
timestamp 1386234792
transform 1 0 19393 0 1 7275
box 0 0 96 799
use inv g459
timestamp 1386238110
transform 1 0 19489 0 1 7275
box 0 0 120 799
use trisbuf g9435
timestamp 1386237216
transform 1 0 19609 0 1 7275
box 0 0 216 799
use nand2 g9799
timestamp 1386234792
transform 1 0 19825 0 1 7275
box 0 0 96 799
use inv g9677
timestamp 1386238110
transform 1 0 19921 0 1 7275
box 0 0 120 799
use nand2 g9707
timestamp 1386234792
transform 1 0 20041 0 1 7275
box 0 0 96 799
use inv g9529
timestamp 1386238110
transform 1 0 20137 0 1 7275
box 0 0 120 799
use nand2 g9453
timestamp 1386234792
transform 1 0 20257 0 1 7275
box 0 0 96 799
use nand3 g9746
timestamp 1386234893
transform 1 0 20353 0 1 7275
box 0 0 120 799
use mux2 g9761
timestamp 1386235218
transform 1 0 20473 0 1 7275
box 0 0 192 799
use nand2 g9700
timestamp 1386234792
transform 1 0 20665 0 1 7275
box 0 0 96 799
use inv g9551
timestamp 1386238110
transform 1 0 20761 0 1 7275
box 0 0 120 799
use nand2 g9636
timestamp 1386234792
transform 1 0 20881 0 1 7275
box 0 0 96 799
use nand2 g9757
timestamp 1386234792
transform 1 0 20977 0 1 7275
box 0 0 96 799
use inv g9457
timestamp 1386238110
transform 1 0 21073 0 1 7275
box 0 0 120 799
use nand2 g9569
timestamp 1386234792
transform 1 0 21193 0 1 7275
box 0 0 96 799
use nand3 g9628
timestamp 1386234893
transform 1 0 21289 0 1 7275
box 0 0 120 799
use and2 g9693
timestamp 1386234845
transform 1 0 21409 0 1 7275
box 0 0 120 799
use and2 g9559
timestamp 1386234845
transform 1 0 21529 0 1 7275
box 0 0 120 799
use nand2 g9733
timestamp 1386234792
transform 1 0 21649 0 1 7275
box 0 0 96 799
use nand2 g9771
timestamp 1386234792
transform 1 0 21745 0 1 7275
box 0 0 96 799
use and2 g9621
timestamp 1386234845
transform 1 0 21841 0 1 7275
box 0 0 120 799
use inv g9517
timestamp 1386238110
transform 1 0 21961 0 1 7275
box 0 0 120 799
use nand2 g9537
timestamp 1386234792
transform 1 0 22081 0 1 7275
box 0 0 96 799
use nand2 g9631
timestamp 1386234792
transform 1 0 22177 0 1 7275
box 0 0 96 799
use nand2 g9510
timestamp 1386234792
transform 1 0 22273 0 1 7275
box 0 0 96 799
use inv StatusReg_reg_91_0_93_
timestamp 1386238110
transform 1 0 22369 0 1 7275
box 0 0 120 799
use scandtype g9742
timestamp 1386241841
transform 1 0 22489 0 1 7275
box 0 0 624 799
use nand3 g9658
timestamp 1386234893
transform 1 0 23113 0 1 7275
box 0 0 120 799
use inv g9779
timestamp 1386238110
transform 1 0 23233 0 1 7275
box 0 0 120 799
use nand2 g9728
timestamp 1386234792
transform 1 0 23353 0 1 7275
box 0 0 96 799
use inv g9417
timestamp 1386238110
transform 1 0 23449 0 1 7275
box 0 0 120 799
use nand4 g9503
timestamp 1386234936
transform 1 0 23569 0 1 7275
box 0 0 144 799
use nand2 g9580
timestamp 1386234792
transform 1 0 23713 0 1 7275
box 0 0 96 799
use nor2 g9718
timestamp 1386235306
transform 1 0 23809 0 1 7275
box 0 0 120 799
use nand2 g9710
timestamp 1386234792
transform 1 0 23929 0 1 7275
box 0 0 96 799
use and2 g9563
timestamp 1386234845
transform 1 0 24025 0 1 7275
box 0 0 120 799
use nand3 g9678
timestamp 1386234893
transform 1 0 24145 0 1 7275
box 0 0 120 799
use nand2 g9618
timestamp 1386234792
transform 1 0 24265 0 1 7275
box 0 0 96 799
use nand2 g9439
timestamp 1386234792
transform 1 0 24361 0 1 7275
box 0 0 96 799
use nand2 g9781
timestamp 1386234792
transform 1 0 24457 0 1 7275
box 0 0 96 799
use and2 g9647
timestamp 1386234845
transform 1 0 24553 0 1 7275
box 0 0 120 799
use nor2 g9642
timestamp 1386235306
transform 1 0 24673 0 1 7275
box 0 0 120 799
use nand2 g9716
timestamp 1386234792
transform 1 0 24793 0 1 7275
box 0 0 96 799
use nand2 g9437
timestamp 1386234792
transform 1 0 24889 0 1 7275
box 0 0 96 799
use nand2 g9769
timestamp 1386234792
transform 1 0 24985 0 1 7275
box 0 0 96 799
use inv g9546
timestamp 1386238110
transform 1 0 25081 0 1 7275
box 0 0 120 799
use nand3 g9564
timestamp 1386234893
transform 1 0 25201 0 1 7275
box 0 0 120 799
use and2 g9585
timestamp 1386234845
transform 1 0 25321 0 1 7275
box 0 0 120 799
use nand2 g9663
timestamp 1386234792
transform 1 0 25441 0 1 7275
box 0 0 96 799
use nand2 g9765
timestamp 1386234792
transform 1 0 25537 0 1 7275
box 0 0 96 799
use nor2 g9601
timestamp 1386235306
transform 1 0 25633 0 1 7275
box 0 0 120 799
use nor2 g9420
timestamp 1386235306
transform 1 0 25753 0 1 7275
box 0 0 120 799
use nand3 g1
timestamp 1386234893
transform 1 0 25873 0 1 7275
box 0 0 120 799
use trisbuf g9660
timestamp 1386237216
transform 1 0 25993 0 1 7275
box 0 0 216 799
use nand3 g9442
timestamp 1386234893
transform 1 0 26209 0 1 7275
box 0 0 120 799
use nand2 g9668
timestamp 1386234792
transform 1 0 26329 0 1 7275
box 0 0 96 799
use nand2 g9656
timestamp 1386234792
transform 1 0 26425 0 1 7275
box 0 0 96 799
use nand2 g9598
timestamp 1386234792
transform 1 0 26521 0 1 7275
box 0 0 96 799
use nand2 g9796
timestamp 1386234792
transform 1 0 26617 0 1 7275
box 0 0 96 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 26713 0 1 7275
box 0 0 48 799
use inv g9591
timestamp 1386238110
transform 1 0 26761 0 1 7275
box 0 0 120 799
use nand2 g9589
timestamp 1386234792
transform 1 0 26881 0 1 7275
box 0 0 96 799
use and2 g9800
timestamp 1386234845
transform 1 0 26977 0 1 7275
box 0 0 120 799
use inv g9533
timestamp 1386238110
transform 1 0 27097 0 1 7275
box 0 0 120 799
use nand2 g9711
timestamp 1386234792
transform 1 0 27217 0 1 7275
box 0 0 96 799
use inv g9592
timestamp 1386238110
transform 1 0 27313 0 1 7275
box 0 0 120 799
use and2 g9722
timestamp 1386234845
transform 1 0 27433 0 1 7275
box 0 0 120 799
use nand2 g9683
timestamp 1386234792
transform 1 0 27553 0 1 7275
box 0 0 96 799
use nor2 AluOR_91_1_93_
timestamp 1386235306
transform 1 0 27649 0 1 7275
box 0 0 120 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27842 0 1 7275
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 145 0 1 1090
box 0 0 1464 799
use nand2 stateSub_reg_91_0_93_
timestamp 1386234792
transform 1 0 1609 0 1 1090
box 0 0 96 799
use rowcrosser g9419
timestamp 1386086759
transform 1 0 1705 0 1 1090
box 0 0 48 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 1753 0 1 1090
box 0 0 48 799
use scandtype g9603
timestamp 1386241841
transform 1 0 1801 0 1 1090
box 0 0 624 799
use nand2 g9713
timestamp 1386234792
transform 1 0 2425 0 1 1090
box 0 0 96 799
use nand2 g9788
timestamp 1386234792
transform 1 0 2521 0 1 1090
box 0 0 96 799
use nand2 g9455
timestamp 1386234792
transform 1 0 2617 0 1 1090
box 0 0 96 799
use nand2 g9725
timestamp 1386234792
transform 1 0 2713 0 1 1090
box 0 0 96 799
use and2 g9484
timestamp 1386234845
transform 1 0 2809 0 1 1090
box 0 0 120 799
use nand2 g9791
timestamp 1386234792
transform 1 0 2929 0 1 1090
box 0 0 96 799
use inv state_reg_91_1_93_
timestamp 1386238110
transform 1 0 3025 0 1 1090
box 0 0 120 799
use scandtype g9750
timestamp 1386241841
transform 1 0 3145 0 1 1090
box 0 0 624 799
use inv g9477
timestamp 1386238110
transform 1 0 3769 0 1 1090
box 0 0 120 799
use nand4 g9708
timestamp 1386234936
transform 1 0 3889 0 1 1090
box 0 0 144 799
use nor2 g9560
timestamp 1386235306
transform 1 0 4033 0 1 1090
box 0 0 120 799
use nor2 g9744
timestamp 1386235306
transform 1 0 4153 0 1 1090
box 0 0 120 799
use nand2 g9542
timestamp 1386234792
transform 1 0 4273 0 1 1090
box 0 0 96 799
use nand3 g9599
timestamp 1386234893
transform 1 0 4369 0 1 1090
box 0 0 120 799
use nor2 g9586
timestamp 1386235306
transform 1 0 4489 0 1 1090
box 0 0 120 799
use nand2 g9570
timestamp 1386234792
transform 1 0 4609 0 1 1090
box 0 0 96 799
use nor2 g9689
timestamp 1386235306
transform 1 0 4705 0 1 1090
box 0 0 120 799
use and2 g9649
timestamp 1386234845
transform 1 0 4825 0 1 1090
box 0 0 120 799
use nand2 g9611
timestamp 1386234792
transform 1 0 4945 0 1 1090
box 0 0 96 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 5041 0 1 1090
box 0 0 96 799
use scandtype g9472
timestamp 1386241841
transform 1 0 5137 0 1 1090
box 0 0 624 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 5761 0 1 1090
box 0 0 48 799
use nand2 g9620
timestamp 1386234792
transform 1 0 5809 0 1 1090
box 0 0 96 799
use nand2 g9550
timestamp 1386234792
transform 1 0 5905 0 1 1090
box 0 0 96 799
use inv g9433
timestamp 1386238110
transform 1 0 6001 0 1 1090
box 0 0 120 799
use nand4 g9485
timestamp 1386234936
transform 1 0 6121 0 1 1090
box 0 0 144 799
use nor2 g9566
timestamp 1386235306
transform 1 0 6265 0 1 1090
box 0 0 120 799
use and2 g9490
timestamp 1386234845
transform 1 0 6385 0 1 1090
box 0 0 120 799
use nand3 g9793
timestamp 1386234893
transform 1 0 6505 0 1 1090
box 0 0 120 799
use inv g9467
timestamp 1386238110
transform 1 0 6625 0 1 1090
box 0 0 120 799
use nand2 g9554
timestamp 1386234792
transform 1 0 6745 0 1 1090
box 0 0 96 799
use nand3 g9734
timestamp 1386234893
transform 1 0 6841 0 1 1090
box 0 0 120 799
use and2 g9754
timestamp 1386234845
transform 1 0 6961 0 1 1090
box 0 0 120 799
use inv g9624
timestamp 1386238110
transform 1 0 7081 0 1 1090
box 0 0 120 799
use nand2 g9640
timestamp 1386234792
transform 1 0 7201 0 1 1090
box 0 0 96 799
use nand4 g9760
timestamp 1386234936
transform 1 0 7297 0 1 1090
box 0 0 144 799
use inv g9495
timestamp 1386238110
transform 1 0 7441 0 1 1090
box 0 0 120 799
use nand2 g9514
timestamp 1386234792
transform 1 0 7561 0 1 1090
box 0 0 96 799
use nor2 g9428
timestamp 1386235306
transform 1 0 7657 0 1 1090
box 0 0 120 799
use nand2 g9650
timestamp 1386234792
transform 1 0 7777 0 1 1090
box 0 0 96 799
use nand2 g9706
timestamp 1386234792
transform 1 0 7873 0 1 1090
box 0 0 96 799
use nand2 IntReq_reg
timestamp 1386234792
transform 1 0 7969 0 1 1090
box 0 0 96 799
use scandtype g9460
timestamp 1386241841
transform 1 0 8065 0 1 1090
box 0 0 624 799
use nor2 g9696
timestamp 1386235306
transform 1 0 8689 0 1 1090
box 0 0 120 799
use xor2 g9609
timestamp 1386237344
transform 1 0 8809 0 1 1090
box 0 0 192 799
use inv g9703
timestamp 1386238110
transform 1 0 9001 0 1 1090
box 0 0 120 799
use nand2 g9424
timestamp 1386234792
transform 1 0 9121 0 1 1090
box 0 0 96 799
use nand3 g9637
timestamp 1386234893
transform 1 0 9217 0 1 1090
box 0 0 120 799
use nand2 g9680
timestamp 1386234792
transform 1 0 9337 0 1 1090
box 0 0 96 799
use nand2 g9443
timestamp 1386234792
transform 1 0 9433 0 1 1090
box 0 0 96 799
use nand2 g457
timestamp 1386234792
transform 1 0 9529 0 1 1090
box 0 0 96 799
use trisbuf g9582
timestamp 1386237216
transform 1 0 9625 0 1 1090
box 0 0 216 799
use nand2 g458
timestamp 1386234792
transform 1 0 9841 0 1 1090
box 0 0 96 799
use trisbuf g9801
timestamp 1386237216
transform 1 0 9937 0 1 1090
box 0 0 216 799
use inv g9501
timestamp 1386238110
transform 1 0 10153 0 1 1090
box 0 0 120 799
use nand3 g9558
timestamp 1386234893
transform 1 0 10273 0 1 1090
box 0 0 120 799
use nand2 g9775
timestamp 1386234792
transform 1 0 10393 0 1 1090
box 0 0 96 799
use nand2 g9426
timestamp 1386234792
transform 1 0 10489 0 1 1090
box 0 0 96 799
use nand4 g9511
timestamp 1386234936
transform 1 0 10585 0 1 1090
box 0 0 144 799
use nand4 g9404
timestamp 1386234936
transform 1 0 10729 0 1 1090
box 0 0 144 799
use nand3 g9646
timestamp 1386234893
transform 1 0 10873 0 1 1090
box 0 0 120 799
use inv g9615
timestamp 1386238110
transform 1 0 10993 0 1 1090
box 0 0 120 799
use nand2 g9581
timestamp 1386234792
transform 1 0 11113 0 1 1090
box 0 0 96 799
use nand4 g9766
timestamp 1386234936
transform 1 0 11209 0 1 1090
box 0 0 144 799
use inv g9743
timestamp 1386238110
transform 1 0 11353 0 1 1090
box 0 0 120 799
use nand2 g9459
timestamp 1386234792
transform 1 0 11473 0 1 1090
box 0 0 96 799
use nor2 g9667
timestamp 1386235306
transform 1 0 11569 0 1 1090
box 0 0 120 799
use nand2 g9481
timestamp 1386234792
transform 1 0 11689 0 1 1090
box 0 0 96 799
use nand4 g9732
timestamp 1386234936
transform 1 0 11785 0 1 1090
box 0 0 144 799
use nand2 g9576
timestamp 1386234792
transform 1 0 11929 0 1 1090
box 0 0 96 799
use nand2 g9764
timestamp 1386234792
transform 1 0 12025 0 1 1090
box 0 0 96 799
use nand2 g9466
timestamp 1386234792
transform 1 0 12121 0 1 1090
box 0 0 96 799
use nand2 g9519
timestamp 1386234792
transform 1 0 12217 0 1 1090
box 0 0 96 799
use nand3 g9770
timestamp 1386234893
transform 1 0 12313 0 1 1090
box 0 0 120 799
use nand2 g9661
timestamp 1386234792
transform 1 0 12433 0 1 1090
box 0 0 96 799
use nand2 g9619
timestamp 1386234792
transform 1 0 12529 0 1 1090
box 0 0 96 799
use nor2 g9508
timestamp 1386235306
transform 1 0 12625 0 1 1090
box 0 0 120 799
use inv g9532
timestamp 1386238110
transform 1 0 12745 0 1 1090
box 0 0 120 799
use nand2 g9413
timestamp 1386234792
transform 1 0 12865 0 1 1090
box 0 0 96 799
use nand4 g9739
timestamp 1386234936
transform 1 0 12961 0 1 1090
box 0 0 144 799
use rowcrosser Rs1Sel_91_1_93_
timestamp 1386086759
transform 1 0 13105 0 1 1090
box 0 0 48 799
use nand2 g9782
timestamp 1386234792
transform 1 0 13153 0 1 1090
box 0 0 96 799
use nand2 g9657
timestamp 1386234792
transform 1 0 13249 0 1 1090
box 0 0 96 799
use nand2 g9692
timestamp 1386234792
transform 1 0 13345 0 1 1090
box 0 0 96 799
use nand2 g9684
timestamp 1386234792
transform 1 0 13441 0 1 1090
box 0 0 96 799
use nand2 g9789
timestamp 1386234792
transform 1 0 13537 0 1 1090
box 0 0 96 799
use nand2 g9516
timestamp 1386234792
transform 1 0 13633 0 1 1090
box 0 0 96 799
use nor2 g9721
timestamp 1386235306
transform 1 0 13729 0 1 1090
box 0 0 120 799
use nand2 g9726
timestamp 1386234792
transform 1 0 13849 0 1 1090
box 0 0 96 799
use nand2 g9449
timestamp 1386234792
transform 1 0 13945 0 1 1090
box 0 0 96 799
use nand4 g9504
timestamp 1386234936
transform 1 0 14041 0 1 1090
box 0 0 144 799
use nand3 g9729
timestamp 1386234893
transform 1 0 14185 0 1 1090
box 0 0 120 799
use nand2 g9709
timestamp 1386234792
transform 1 0 14305 0 1 1090
box 0 0 96 799
use nand2 InISR_reg
timestamp 1386234792
transform 1 0 14401 0 1 1090
box 0 0 96 799
use scandtype g9483
timestamp 1386241841
transform 1 0 14497 0 1 1090
box 0 0 624 799
use nand2 g9688
timestamp 1386234792
transform 1 0 15121 0 1 1090
box 0 0 96 799
use and2 g9664
timestamp 1386234845
transform 1 0 15217 0 1 1090
box 0 0 120 799
use nand2 g9412
timestamp 1386234792
transform 1 0 15337 0 1 1090
box 0 0 96 799
use nand2 g9740
timestamp 1386234792
transform 1 0 15433 0 1 1090
box 0 0 96 799
use inv g9648
timestamp 1386238110
transform 1 0 15529 0 1 1090
box 0 0 120 799
use inv g9505
timestamp 1386238110
transform 1 0 15649 0 1 1090
box 0 0 120 799
use inv g9480
timestamp 1386238110
transform 1 0 15769 0 1 1090
box 0 0 120 799
use inv g9702
timestamp 1386238110
transform 1 0 15889 0 1 1090
box 0 0 120 799
use nor2 g9630
timestamp 1386235306
transform 1 0 16009 0 1 1090
box 0 0 120 799
use rowcrosser nWE
timestamp 1386086759
transform 1 0 16129 0 1 1090
box 0 0 48 799
use nand2 g9623
timestamp 1386234792
transform 1 0 16177 0 1 1090
box 0 0 96 799
use and2 g9526
timestamp 1386234845
transform 1 0 16273 0 1 1090
box 0 0 120 799
use nand2 g9451
timestamp 1386234792
transform 1 0 16393 0 1 1090
box 0 0 96 799
use nand4 g9625
timestamp 1386234936
transform 1 0 16489 0 1 1090
box 0 0 144 799
use nand2 g9593
timestamp 1386234792
transform 1 0 16633 0 1 1090
box 0 0 96 799
use nand2 g9565
timestamp 1386234792
transform 1 0 16729 0 1 1090
box 0 0 96 799
use nand2 IRQ2_reg
timestamp 1386234792
transform 1 0 16825 0 1 1090
box 0 0 96 799
use scandtype g9745
timestamp 1386241841
transform 1 0 16921 0 1 1090
box 0 0 624 799
use nand3 g9751
timestamp 1386234893
transform 1 0 17545 0 1 1090
box 0 0 120 799
use nand2 g9634
timestamp 1386234792
transform 1 0 17665 0 1 1090
box 0 0 96 799
use nand3 g9604
timestamp 1386234893
transform 1 0 17761 0 1 1090
box 0 0 120 799
use nand3 g9792
timestamp 1386234893
transform 1 0 17881 0 1 1090
box 0 0 120 799
use inv g9639
timestamp 1386238110
transform 1 0 18001 0 1 1090
box 0 0 120 799
use nand2 g9573
timestamp 1386234792
transform 1 0 18121 0 1 1090
box 0 0 96 799
use nor2 g9602
timestamp 1386235306
transform 1 0 18217 0 1 1090
box 0 0 120 799
use nor2 g9714
timestamp 1386235306
transform 1 0 18337 0 1 1090
box 0 0 120 799
use nand2 g9773
timestamp 1386234792
transform 1 0 18457 0 1 1090
box 0 0 96 799
use and2 g9787
timestamp 1386234845
transform 1 0 18553 0 1 1090
box 0 0 120 799
use inv g9610
timestamp 1386238110
transform 1 0 18673 0 1 1090
box 0 0 120 799
use nor2 g9547
timestamp 1386235306
transform 1 0 18793 0 1 1090
box 0 0 120 799
use nand3 g9587
timestamp 1386234893
transform 1 0 18913 0 1 1090
box 0 0 120 799
use nand4 g9571
timestamp 1386234936
transform 1 0 19033 0 1 1090
box 0 0 144 799
use nand3 g9445
timestamp 1386234893
transform 1 0 19177 0 1 1090
box 0 0 120 799
use and2 g9523
timestamp 1386234845
transform 1 0 19297 0 1 1090
box 0 0 120 799
use nand2 g9421
timestamp 1386234792
transform 1 0 19417 0 1 1090
box 0 0 96 799
use nand3 g9432
timestamp 1386234893
transform 1 0 19513 0 1 1090
box 0 0 120 799
use nand4 g9473
timestamp 1386234936
transform 1 0 19633 0 1 1090
box 0 0 144 799
use nand2 IRQ1_reg
timestamp 1386234792
transform 1 0 19777 0 1 1090
box 0 0 96 799
use scandtype g9614
timestamp 1386241841
transform 1 0 19873 0 1 1090
box 0 0 624 799
use and2 g9651
timestamp 1386234845
transform 1 0 20497 0 1 1090
box 0 0 120 799
use nand2 g9541
timestamp 1386234792
transform 1 0 20617 0 1 1090
box 0 0 96 799
use nand2 g9617
timestamp 1386234792
transform 1 0 20713 0 1 1090
box 0 0 96 799
use nand2 g9506
timestamp 1386234792
transform 1 0 20809 0 1 1090
box 0 0 96 799
use nand3 g9596
timestamp 1386234893
transform 1 0 20905 0 1 1090
box 0 0 120 799
use nand3 g9450
timestamp 1386234893
transform 1 0 21025 0 1 1090
box 0 0 120 799
use nand3 g9645
timestamp 1386234893
transform 1 0 21145 0 1 1090
box 0 0 120 799
use nor2 g9553
timestamp 1386235306
transform 1 0 21265 0 1 1090
box 0 0 120 799
use nand3 g9454
timestamp 1386234893
transform 1 0 21385 0 1 1090
box 0 0 120 799
use and2 g9461
timestamp 1386234845
transform 1 0 21505 0 1 1090
box 0 0 120 799
use and2 g9543
timestamp 1386234845
transform 1 0 21625 0 1 1090
box 0 0 120 799
use nand2 g9735
timestamp 1386234792
transform 1 0 21745 0 1 1090
box 0 0 96 799
use inv g9629
timestamp 1386238110
transform 1 0 21841 0 1 1090
box 0 0 120 799
use nand2 g9567
timestamp 1386234792
transform 1 0 21961 0 1 1090
box 0 0 96 799
use nand2 g9723
timestamp 1386234792
transform 1 0 22057 0 1 1090
box 0 0 96 799
use nand2 g9436
timestamp 1386234792
transform 1 0 22153 0 1 1090
box 0 0 96 799
use nand2 g9561
timestamp 1386234792
transform 1 0 22249 0 1 1090
box 0 0 96 799
use and2 g9531
timestamp 1386234845
transform 1 0 22345 0 1 1090
box 0 0 120 799
use nand2 g9491
timestamp 1386234792
transform 1 0 22465 0 1 1090
box 0 0 96 799
use and2 g9676
timestamp 1386234845
transform 1 0 22561 0 1 1090
box 0 0 120 799
use nand2 g9496
timestamp 1386234792
transform 1 0 22681 0 1 1090
box 0 0 96 799
use nand3 g9574
timestamp 1386234893
transform 1 0 22777 0 1 1090
box 0 0 120 799
use and2 g9783
timestamp 1386234845
transform 1 0 22897 0 1 1090
box 0 0 120 799
use nand2 g9662
timestamp 1386234792
transform 1 0 23017 0 1 1090
box 0 0 96 799
use nand2 g9444
timestamp 1386234792
transform 1 0 23113 0 1 1090
box 0 0 96 799
use nand2 g9418
timestamp 1386234792
transform 1 0 23209 0 1 1090
box 0 0 96 799
use nand4 g9776
timestamp 1386234936
transform 1 0 23305 0 1 1090
box 0 0 144 799
use inv g9608
timestamp 1386238110
transform 1 0 23449 0 1 1090
box 0 0 120 799
use nand2 g9749
timestamp 1386234792
transform 1 0 23569 0 1 1090
box 0 0 96 799
use nor2 g9767
timestamp 1386235306
transform 1 0 23665 0 1 1090
box 0 0 120 799
use nand2 g9681
timestamp 1386234792
transform 1 0 23785 0 1 1090
box 0 0 96 799
use nand3 g9695
timestamp 1386234893
transform 1 0 23881 0 1 1090
box 0 0 120 799
use and2 g9557
timestamp 1386234845
transform 1 0 24001 0 1 1090
box 0 0 120 799
use nor2 g9536
timestamp 1386235306
transform 1 0 24121 0 1 1090
box 0 0 120 799
use inv g9638
timestamp 1386238110
transform 1 0 24241 0 1 1090
box 0 0 120 799
use nand3 g9548
timestamp 1386234893
transform 1 0 24361 0 1 1090
box 0 0 120 799
use nand2 g9685
timestamp 1386234792
transform 1 0 24481 0 1 1090
box 0 0 96 799
use nand2 g9705
timestamp 1386234792
transform 1 0 24577 0 1 1090
box 0 0 96 799
use and2 g9671
timestamp 1386234845
transform 1 0 24673 0 1 1090
box 0 0 120 799
use inv g9465
timestamp 1386238110
transform 1 0 24793 0 1 1090
box 0 0 120 799
use and2 g9720
timestamp 1386234845
transform 1 0 24913 0 1 1090
box 0 0 120 799
use nor2 g9691
timestamp 1386235306
transform 1 0 25033 0 1 1090
box 0 0 120 799
use nand2 g9590
timestamp 1386234792
transform 1 0 25153 0 1 1090
box 0 0 96 799
use nand2 g9752
timestamp 1386234792
transform 1 0 25249 0 1 1090
box 0 0 96 799
use nand2 g9654
timestamp 1386234792
transform 1 0 25345 0 1 1090
box 0 0 96 799
use and2 g9577
timestamp 1386234845
transform 1 0 25441 0 1 1090
box 0 0 120 799
use nand2 g9415
timestamp 1386234792
transform 1 0 25561 0 1 1090
box 0 0 96 799
use nor2 g9403
timestamp 1386235306
transform 1 0 25657 0 1 1090
box 0 0 120 799
use nand4 g9498
timestamp 1386234936
transform 1 0 25777 0 1 1090
box 0 0 144 799
use nand2 g9697
timestamp 1386234792
transform 1 0 25921 0 1 1090
box 0 0 96 799
use nand2 g9665
timestamp 1386234792
transform 1 0 26017 0 1 1090
box 0 0 96 799
use nand2 g9448
timestamp 1386234792
transform 1 0 26113 0 1 1090
box 0 0 96 799
use inv state_reg_91_0_93_
timestamp 1386238110
transform 1 0 26209 0 1 1090
box 0 0 120 799
use scandtype g9430
timestamp 1386241841
transform 1 0 26329 0 1 1090
box 0 0 624 799
use nand4 stateSub_reg_91_1_93_
timestamp 1386234936
transform 1 0 26953 0 1 1090
box 0 0 144 799
use scandtype g9488
timestamp 1386241841
transform 1 0 27097 0 1 1090
box 0 0 624 799
use nand3 Flags_91_1_93_
timestamp 1386234893
transform 1 0 27721 0 1 1090
box 0 0 120 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27841 0 1 1090
box 0 0 320 799
<< labels >>
rlabel m2contact 26815 8187 26815 8187 6 Flags[0]
rlabel m2contact 26815 8115 26815 8115 6 Flags[0]
rlabel m2contact 26791 8163 26791 8163 6 SysBus[3]
rlabel m2contact 26791 8091 26791 8091 6 SysBus[3]
rlabel metal2 26761 8115 26761 8115 6 LrSel
rlabel m2contact 26743 8115 26743 8115 6 LrSel
rlabel m2contact 26167 8163 26167 8163 6 SysBus[3]
rlabel m2contact 25015 8091 25015 8091 6 SysBus[1]
rlabel m2contact 24487 8163 24487 8163 6 SysBus[3]
rlabel m2contact 23695 8163 23695 8163 6 RwSel[0]
rlabel m2contact 23527 8235 23527 8235 6 OpcodeCondIn[4]
rlabel m2contact 21343 8115 21343 8115 6 Op2Sel[0]
rlabel m2contact 20383 8235 20383 8235 6 OpcodeCondIn[4]
rlabel m2contact 19783 8139 19783 8139 6 SysBus[0]
rlabel m2contact 19159 8139 19159 8139 6 OpcodeCondIn[2]
rlabel metal2 18049 8235 18049 8235 6 SysBus[2]
rlabel m2contact 18031 8235 18031 8235 6 SysBus[2]
rlabel m2contact 17623 8187 17623 8187 6 Flags[0]
rlabel m2contact 17503 8211 17503 8211 6 PcSel[2]
rlabel m2contact 16615 8139 16615 8139 6 OpcodeCondIn[2]
rlabel m2contact 16471 8211 16471 8211 6 PcSel[2]
rlabel m2contact 14791 8187 14791 8187 6 OpcodeCondIn[0]
rlabel m2contact 12607 8139 12607 8139 4 PcSel[1]
rlabel m2contact 12571 8163 12571 8163 4 RwSel[0]
rlabel m2contact 11215 8163 11215 8163 4 nIRQ
rlabel m2contact 10375 8163 10375 8163 4 nIRQ
rlabel m2contact 9967 8163 9967 8163 4 Op2Sel[1]
rlabel m2contact 8599 8187 8599 8187 4 OpcodeCondIn[0]
rlabel m2contact 7879 8187 7879 8187 4 OpcodeCondIn[5]
rlabel m2contact 6991 8115 6991 8115 4 Op2Sel[0]
rlabel metal2 6673 8115 6673 8115 4 AluOR[1]
rlabel m2contact 6655 8115 6655 8115 4 AluOR[1]
rlabel m2contact 5743 8115 5743 8115 4 PcSel[0]
rlabel m2contact 4807 8211 4807 8211 4 PcSel[2]
rlabel m2contact 3823 8211 3823 8211 4 ENB
rlabel m2contact 3787 8091 3787 8091 4 SysBus[1]
rlabel m2contact 2983 8211 2983 8211 4 ENB
rlabel m2contact 2743 8139 2743 8139 4 PcSel[1]
rlabel m2contact 1759 8139 1759 8139 4 OpcodeCondIn[7]
rlabel m2contact 27055 89 27055 89 8 n_382
rlabel m2contact 27031 713 27031 713 8 n_383
rlabel m2contact 27007 833 27007 833 6 n_245
rlabel m2contact 26983 401 26983 401 8 n_223
rlabel m2contact 26431 977 26431 977 6 n_350
rlabel m2contact 26239 377 26239 377 8 n_300
rlabel m2contact 26095 857 26095 857 6 n_28
rlabel m2contact 25999 665 25999 665 8 n_203
rlabel m2contact 25903 761 25903 761 8 ImmSel
rlabel m2contact 25759 641 25759 641 8 n_388
rlabel m2contact 25591 689 25591 689 8 n_140
rlabel m2contact 25579 593 25579 593 8 IrWe
rlabel m2contact 24967 665 24967 665 8 n_203
rlabel m2contact 24655 665 24655 665 8 n_78
rlabel m2contact 24463 425 24463 425 8 n_129
rlabel m2contact 24439 329 24439 329 8 OpcodeCondIn[3]
rlabel m2contact 24223 737 24223 737 8 n_197
rlabel m2contact 24175 281 24175 281 8 n_53
rlabel m2contact 24103 593 24103 593 8 IrWe
rlabel m2contact 23983 281 23983 281 8 n_53
rlabel m2contact 23959 329 23959 329 8 OpcodeCondIn[3]
rlabel m2contact 23719 41 23719 41 8 OpcodeCondIn[1]
rlabel m2contact 23647 881 23647 881 6 n_148
rlabel m2contact 23599 1025 23599 1025 6 n_103
rlabel m2contact 23431 545 23431 545 8 AluEn
rlabel m2contact 23407 329 23407 329 8 OpcodeCondIn[3]
rlabel m2contact 23383 713 23383 713 8 n_383
rlabel m2contact 23191 929 23191 929 6 n_102
rlabel m2contact 23143 449 23143 449 8 n_67
rlabel m2contact 22927 593 22927 593 8 n_213
rlabel m2contact 22879 545 22879 545 8 n_286
rlabel m2contact 22615 809 22615 809 6 n_141
rlabel m2contact 22591 1049 22591 1049 6 n_229
rlabel m2contact 22231 1073 22231 1073 6 n_43
rlabel m2contact 22135 1001 22135 1001 6 n_196
rlabel m2contact 22111 905 22111 905 6 nWait
rlabel m2contact 22087 785 22087 785 8 n_170
rlabel m2contact 22039 905 22039 905 6 n_162
rlabel m2contact 21823 833 21823 833 6 n_245
rlabel m2contact 21775 521 21775 521 8 n_216
rlabel m2contact 21727 713 21727 713 8 n_383
rlabel m2contact 21463 617 21463 617 8 OpcodeCondIn[6]
rlabel m2contact 21247 569 21247 569 8 MemEn
rlabel m2contact 21235 41 21235 41 8 OpcodeCondIn[1]
rlabel m2contact 21199 569 21199 569 8 n_247
rlabel m2contact 21175 953 21175 953 6 n_209
rlabel m2contact 21127 617 21127 617 8 n_287
rlabel m2contact 21007 233 21007 233 8 n_232
rlabel m2contact 20959 713 20959 713 8 n_175
rlabel m2contact 20887 809 20887 809 6 n_141
rlabel m2contact 20791 569 20791 569 8 n_247
rlabel m2contact 20743 569 20743 569 8 n_246
rlabel m2contact 20695 305 20695 305 8 n_84
rlabel m2contact 20599 809 20599 809 6 n_326
rlabel m2contact 20551 665 20551 665 8 n_78
rlabel m2contact 20383 833 20383 833 6 IRQ1
rlabel m2contact 19855 161 19855 161 8 LrEn
rlabel m2contact 19831 665 19831 665 8 n_242
rlabel m2contact 19759 977 19759 977 6 n_350
rlabel m2contact 19711 881 19711 881 6 n_148
rlabel m2contact 19615 473 19615 473 8 n_379
rlabel m2contact 19567 881 19567 881 6 n_308
rlabel m2contact 19495 497 19495 497 8 AluOR[0]
rlabel m2contact 19447 617 19447 617 8 n_287
rlabel m2contact 19327 977 19327 977 6 n_280
rlabel m2contact 19279 713 19279 713 8 n_175
rlabel m2contact 19135 329 19135 329 8 OpcodeCondIn[3]
rlabel m2contact 19063 713 19063 713 8 PcWe
rlabel m2contact 18895 785 18895 785 8 n_170
rlabel m2contact 18607 41 18607 41 8 OpcodeCondIn[1]
rlabel m2contact 18535 353 18535 353 8 n_36
rlabel m2contact 18367 281 18367 281 8 n_53
rlabel m2contact 17983 257 17983 257 8 n_133
rlabel m2contact 17815 353 17815 353 8 n_36
rlabel m2contact 17791 857 17791 857 6 n_28
rlabel m2contact 17623 41 17623 41 8 OpcodeCondIn[1]
rlabel m2contact 17383 857 17383 857 6 n_498
rlabel m2contact 17023 833 17023 833 6 IRQ1
rlabel m2contact 16903 521 16903 521 8 n_216
rlabel m2contact 16891 65 16891 65 8 Flags[1]
rlabel m2contact 16855 137 16855 137 8 n_149
rlabel m2contact 16759 281 16759 281 8 IntReq
rlabel m2contact 16711 521 16711 521 8 n_165
rlabel m2contact 16591 89 16591 89 8 n_382
rlabel m2contact 16471 1049 16471 1049 6 n_229
rlabel m2contact 16327 329 16327 329 8 OpcodeCondIn[3]
rlabel m2contact 16255 689 16255 689 8 n_140
rlabel m2contact 16231 329 16231 329 8 OpcodeCondIn[3]
rlabel m2contact 16159 353 16159 353 8 nME
rlabel m2contact 15919 1049 15919 1049 6 n_338
rlabel m2contact 15847 689 15847 689 8 n_262
rlabel m2contact 15799 233 15799 233 8 n_232
rlabel m2contact 15511 713 15511 713 8 PcWe
rlabel m2contact 15007 209 15007 209 8 n_401
rlabel m2contact 14719 17 14719 17 8 RegWe
rlabel m2contact 14695 353 14695 353 8 nME
rlabel m2contact 14599 233 14599 233 8 n_353
rlabel m2contact 14479 713 14479 713 2 n_48
rlabel m2contact 14167 377 14167 377 2 n_300
rlabel m2contact 14143 1073 14143 1073 4 n_43
rlabel m2contact 13927 1073 13927 1073 4 n_29
rlabel m2contact 13759 353 13759 353 2 n_221
rlabel m2contact 13519 185 13519 185 2 n_119
rlabel m2contact 13279 329 13279 329 2 OpcodeCondIn[3]
rlabel m2contact 13135 113 13135 113 2 Flags[2]
rlabel m2contact 13015 305 13015 305 2 n_84
rlabel m2contact 12991 377 12991 377 2 n_55
rlabel m2contact 12823 305 12823 305 2 n_340
rlabel m2contact 12727 593 12727 593 2 n_213
rlabel m2contact 12655 1073 12655 1073 4 n_29
rlabel m2contact 12607 1025 12607 1025 4 n_103
rlabel m2contact 12415 1025 12415 1025 4 n_258
rlabel m2contact 12295 233 12295 233 2 n_353
rlabel m2contact 12271 89 12271 89 2 n_382
rlabel m2contact 12247 233 12247 233 2 n_337
rlabel m2contact 12055 593 12055 593 2 n_213
rlabel m2contact 11911 1049 11911 1049 4 n_338
rlabel m2contact 11887 905 11887 905 4 n_162
rlabel m2contact 11863 1025 11863 1025 4 n_258
rlabel m2contact 11839 905 11839 905 4 n_185
rlabel m2contact 11815 1001 11815 1001 4 n_196
rlabel m2contact 11767 89 11767 89 2 n_382
rlabel m2contact 11671 977 11671 977 4 n_280
rlabel m2contact 11335 953 11335 953 4 n_209
rlabel m2contact 11143 929 11143 929 4 n_102
rlabel m2contact 10975 17 10975 17 2 RegWe
rlabel m2contact 10951 89 10951 89 2 n_382
rlabel m2contact 10927 641 10927 641 2 n_388
rlabel m2contact 10831 713 10831 713 2 n_48
rlabel m2contact 10807 641 10807 641 2 n_155
rlabel m2contact 10783 257 10783 257 2 n_133
rlabel m2contact 10759 713 10759 713 2 n_33
rlabel m2contact 10711 257 10711 257 2 nOE
rlabel m2contact 10663 689 10663 689 2 n_262
rlabel m2contact 10615 809 10615 809 4 n_326
rlabel m2contact 10471 641 10471 641 2 n_155
rlabel m2contact 10375 641 10375 641 2 n_285
rlabel m2contact 10363 89 10363 89 2 PcEn
rlabel m2contact 10351 689 10351 689 2 n_166
rlabel m2contact 10183 41 10183 41 2 OpcodeCondIn[1]
rlabel metal2 9985 41 9985 41 2 CFlag
rlabel m2contact 9967 41 9967 41 2 CFlag
rlabel m2contact 9919 905 9919 905 4 n_185
rlabel m2contact 9607 881 9607 881 4 n_308
rlabel m2contact 9487 857 9487 857 4 n_498
rlabel m2contact 9463 833 9463 833 4 IRQ1
rlabel m2contact 9319 89 9319 89 2 PcEn
rlabel m2contact 9295 809 9295 809 4 n_326
rlabel m2contact 9271 89 9271 89 2 n_319
rlabel m2contact 9247 305 9247 305 2 n_340
rlabel m2contact 9079 305 9079 305 2 n_171
rlabel m2contact 9031 785 9031 785 2 n_170
rlabel m2contact 8575 281 8575 281 2 IntReq
rlabel m2contact 8143 761 8143 761 2 ImmSel
rlabel m2contact 8047 449 8047 449 2 n_67
rlabel m2contact 7711 737 7711 737 2 n_197
rlabel m2contact 7687 449 7687 449 2 n_92
rlabel m2contact 7423 713 7423 713 2 n_33
rlabel m2contact 7279 689 7279 689 2 n_166
rlabel m2contact 6943 665 6943 665 2 n_242
rlabel m2contact 6775 641 6775 641 2 n_285
rlabel m2contact 6559 617 6559 617 2 n_287
rlabel m2contact 6487 569 6487 569 2 n_246
rlabel m2contact 6415 593 6415 593 2 n_213
rlabel m2contact 6295 569 6295 569 2 n_246
rlabel m2contact 6175 545 6175 545 2 n_286
rlabel m2contact 6151 521 6151 521 2 n_165
rlabel m2contact 5959 497 5959 497 2 AluOR[0]
rlabel m2contact 5791 65 5791 65 2 Flags[1]
rlabel m2contact 5239 473 5239 473 2 n_379
rlabel m2contact 4927 449 4927 449 2 n_92
rlabel m2contact 4855 281 4855 281 2 IntReq
rlabel m2contact 4639 425 4639 425 2 n_129
rlabel m2contact 4471 401 4471 401 2 n_223
rlabel m2contact 4351 377 4351 377 2 n_55
rlabel m2contact 4255 353 4255 353 2 n_221
rlabel m2contact 4207 329 4207 329 2 OpcodeCondIn[3]
rlabel m2contact 4183 305 4183 305 2 n_171
rlabel m2contact 3967 281 3967 281 2 IntReq
rlabel m2contact 3775 257 3775 257 2 nOE
rlabel m2contact 3007 233 3007 233 2 n_337
rlabel m2contact 2959 209 2959 209 2 n_401
rlabel m2contact 2791 89 2791 89 2 n_319
rlabel m2contact 2503 137 2503 137 2 n_149
rlabel m2contact 1783 89 1783 89 2 nWE
rlabel m2contact 1735 137 1735 137 2 Rs1Sel[1]
rlabel m2contact 1639 185 1639 185 2 n_119
rlabel m2contact 27871 2914 27871 2914 6 Op1Sel
rlabel m2contact 27871 1930 27871 1930 6 Op1Sel
rlabel m2contact 27847 4594 27847 4594 6 AluWe
rlabel m2contact 27847 1906 27847 1906 6 AluWe
rlabel m2contact 27823 4762 27823 4762 6 n_328
rlabel m2contact 27799 2746 27799 2746 6 n_16
rlabel m2contact 27775 4690 27775 4690 6 n_265
rlabel m2contact 27751 6994 27751 6994 6 n_94
rlabel m2contact 27751 2410 27751 2410 6 n_49
rlabel m2contact 27703 4666 27703 4666 6 n_234
rlabel m2contact 27679 5794 27679 5794 6 n_183
rlabel m2contact 27655 4618 27655 4618 6 n_208
rlabel m2contact 27655 2338 27655 2338 6 n_208
rlabel m2contact 27631 4522 27631 4522 6 n_59
rlabel m2contact 27607 4618 27607 4618 6 n_208
rlabel m2contact 27607 3610 27607 3610 6 stateSub[1]
rlabel m2contact 27583 3658 27583 3658 6 n_73
rlabel m2contact 27559 5026 27559 5026 6 n_224
rlabel m2contact 27535 5578 27535 5578 6 n_189
rlabel m2contact 27487 5650 27487 5650 6 n_142
rlabel m2contact 27463 5962 27463 5962 6 n_132
rlabel m2contact 27391 4714 27391 4714 6 n_65
rlabel m2contact 27343 6202 27343 6202 6 n_64
rlabel m2contact 27295 6922 27295 6922 6 n_251
rlabel m2contact 27271 5794 27271 5794 6 n_183
rlabel m2contact 27247 5194 27247 5194 6 n_278
rlabel m2contact 27199 2890 27199 2890 6 n_390
rlabel m2contact 27175 4546 27175 4546 6 n_1
rlabel m2contact 27127 4570 27127 4570 6 nWait
rlabel m2contact 27079 4594 27079 4594 6 AluWe
rlabel m2contact 27079 5194 27079 5194 6 n_278
rlabel m2contact 27031 5938 27031 5938 6 n_192
rlabel m2contact 27007 4258 27007 4258 6 n_243
rlabel m2contact 26959 4738 26959 4738 6 n_153
rlabel m2contact 26935 3754 26935 3754 6 stateSub[0]
rlabel m2contact 26911 4354 26911 4354 6 n_111
rlabel m2contact 26863 4594 26863 4594 6 n_186
rlabel m2contact 26863 3682 26863 3682 6 n_186
rlabel m2contact 26839 4594 26839 4594 6 n_186
rlabel m2contact 26839 4162 26839 4162 6 state[0]
rlabel m2contact 26791 6178 26791 6178 6 OpcodeCondIn[3]
rlabel m2contact 26791 4402 26791 4402 6 n_18
rlabel m2contact 26743 4594 26743 4594 6 LrSel
rlabel m2contact 26695 4450 26695 4450 6 n_152
rlabel m2contact 26671 3322 26671 3322 6 n_15
rlabel m2contact 26647 2530 26647 2530 6 n_108
rlabel m2contact 26599 4882 26599 4882 6 n_306
rlabel m2contact 26575 5026 26575 5026 6 n_224
rlabel m2contact 26551 2026 26551 2026 6 n_125
rlabel m2contact 26503 2842 26503 2842 6 n_147
rlabel m2contact 26479 5506 26479 5506 6 n_116
rlabel m2contact 26455 7234 26455 7234 6 n_159
rlabel m2contact 26407 4618 26407 4618 6 n_310
rlabel m2contact 26383 4306 26383 4306 6 CFlag
rlabel m2contact 26359 2314 26359 2314 6 n_309
rlabel m2contact 26335 6154 26335 6154 6 OpcodeCondIn[2]
rlabel m2contact 26335 2674 26335 2674 6 OpcodeCondIn[2]
rlabel m2contact 26311 4138 26311 4138 6 n_51
rlabel m2contact 26287 6154 26287 6154 6 OpcodeCondIn[2]
rlabel m2contact 26287 6130 26287 6130 6 n_320
rlabel m2contact 26263 4858 26263 4858 6 n_118
rlabel m2contact 26239 6730 26239 6730 6 n_136
rlabel m2contact 26203 4906 26203 4906 6 n_376
rlabel m2contact 26203 2242 26203 2242 6 n_376
rlabel m2contact 26191 2098 26191 2098 6 n_98
rlabel m2contact 26167 5026 26167 5026 6 n_224
rlabel m2contact 26143 5362 26143 5362 6 n_97
rlabel m2contact 26119 6970 26119 6970 6 n_339
rlabel m2contact 26119 4498 26119 4498 6 n_339
rlabel m2contact 26095 3106 26095 3106 6 n_237
rlabel m2contact 26071 4546 26071 4546 6 n_1
rlabel m2contact 26047 5770 26047 5770 6 n_72
rlabel m2contact 26023 5290 26023 5290 6 StatusReg[3]
rlabel m2contact 25987 6010 25987 6010 6 n_100
rlabel m2contact 25987 4546 25987 4546 6 n_100
rlabel m2contact 25975 7258 25975 7258 6 n_380
rlabel m2contact 25975 3370 25975 3370 6 n_179
rlabel m2contact 25951 4786 25951 4786 6 n_334
rlabel m2contact 25951 3610 25951 3610 6 stateSub[1]
rlabel m2contact 25927 4618 25927 4618 6 n_310
rlabel m2contact 25903 5914 25903 5914 6 n_351
rlabel m2contact 25879 6538 25879 6538 6 n_322
rlabel m2contact 25855 2242 25855 2242 6 n_376
rlabel m2contact 25855 2266 25855 2266 6 n_190
rlabel m2contact 25831 5674 25831 5674 6 n_363
rlabel m2contact 25807 4498 25807 4498 6 n_339
rlabel m2contact 25807 6610 25807 6610 6 OpcodeCondIn[5]
rlabel m2contact 25783 6394 25783 6394 6 n_124
rlabel m2contact 25759 5986 25759 5986 6 n_52
rlabel m2contact 25759 4810 25759 4810 6 n_52
rlabel m2contact 25735 2362 25735 2362 6 n_42
rlabel m2contact 25711 5242 25711 5242 6 n_275
rlabel m2contact 25687 6178 25687 6178 6 OpcodeCondIn[3]
rlabel m2contact 25687 3730 25687 3730 6 n_374
rlabel m2contact 25663 4402 25663 4402 6 n_18
rlabel m2contact 25639 4642 25639 4642 6 n_193
rlabel m2contact 25615 6010 25615 6010 6 n_100
rlabel m2contact 25615 5938 25615 5938 6 n_192
rlabel m2contact 25591 5026 25591 5026 6 n_224
rlabel m2contact 25567 7090 25567 7090 6 n_99
rlabel m2contact 25543 5002 25543 5002 6 n_163
rlabel m2contact 25519 4498 25519 4498 6 n_115
rlabel m2contact 25495 2434 25495 2434 6 n_257
rlabel m2contact 25495 4474 25495 4474 6 OpcodeCondIn[6]
rlabel m2contact 25471 5986 25471 5986 6 n_52
rlabel m2contact 25471 5938 25471 5938 6 n_192
rlabel m2contact 25447 4834 25447 4834 6 n_81
rlabel m2contact 25447 3898 25447 3898 6 n_81
rlabel m2contact 25423 3322 25423 3322 6 n_15
rlabel m2contact 25423 3346 25423 3346 6 n_255
rlabel m2contact 25399 6370 25399 6370 6 n_154
rlabel m2contact 25375 2434 25375 2434 6 n_257
rlabel m2contact 25375 5098 25375 5098 6 n_217
rlabel m2contact 25351 3850 25351 3850 6 n_218
rlabel m2contact 25327 3826 25327 3826 6 n_191
rlabel m2contact 25303 6586 25303 6586 6 n_244
rlabel m2contact 25303 6298 25303 6298 6 n_80
rlabel m2contact 25279 2266 25279 2266 6 n_190
rlabel m2contact 25279 4618 25279 4618 6 n_241
rlabel m2contact 25255 4258 25255 4258 6 n_243
rlabel m2contact 25231 4834 25231 4834 6 n_81
rlabel m2contact 25231 3970 25231 3970 6 n_120
rlabel m2contact 25207 2338 25207 2338 6 n_208
rlabel m2contact 25183 2026 25183 2026 6 n_125
rlabel m2contact 25159 4186 25159 4186 6 n_270
rlabel m2contact 25135 5794 25135 5794 6 n_183
rlabel m2contact 25111 6250 25111 6250 6 n_40
rlabel m2contact 25087 5218 25087 5218 6 n_283
rlabel m2contact 25063 4786 25063 4786 6 n_334
rlabel m2contact 25063 4042 25063 4042 6 n_44
rlabel m2contact 25039 5314 25039 5314 6 n_333
rlabel m2contact 25015 5842 25015 5842 6 SysBus[1]
rlabel m2contact 25015 2866 25015 2866 6 n_249
rlabel m2contact 24967 6754 24967 6754 6 n_46
rlabel m2contact 24943 4498 24943 4498 6 n_115
rlabel m2contact 24943 5218 24943 5218 6 n_283
rlabel m2contact 24919 4042 24919 4042 6 n_44
rlabel m2contact 24883 6418 24883 6418 6 n_500
rlabel m2contact 24883 3130 24883 3130 6 n_500
rlabel m2contact 24871 6466 24871 6466 6 n_86
rlabel m2contact 24871 2626 24871 2626 6 n_167
rlabel m2contact 24847 4282 24847 4282 6 n_400
rlabel m2contact 24823 6418 24823 6418 6 n_500
rlabel m2contact 24823 6394 24823 6394 6 n_124
rlabel m2contact 24799 5818 24799 5818 6 n_110
rlabel m2contact 24799 2122 24799 2122 6 n_110
rlabel m2contact 24775 5818 24775 5818 6 n_110
rlabel m2contact 24775 5746 24775 5746 6 n_160
rlabel m2contact 24727 4498 24727 4498 6 n_71
rlabel m2contact 24727 3274 24727 3274 6 n_70
rlabel m2contact 24703 2434 24703 2434 6 n_257
rlabel m2contact 24703 5410 24703 5410 6 n_109
rlabel m2contact 24655 3538 24655 3538 6 n_274
rlabel m2contact 24631 3322 24631 3322 6 state[1]
rlabel m2contact 24607 3178 24607 3178 6 n_83
rlabel m2contact 24607 4474 24607 4474 6 OpcodeCondIn[6]
rlabel m2contact 24583 4114 24583 4114 6 OpcodeCondIn[7]
rlabel m2contact 24559 6154 24559 6154 6 n_325
rlabel m2contact 24535 6562 24535 6562 6 n_331
rlabel m2contact 24535 3010 24535 3010 6 n_143
rlabel m2contact 24511 5314 24511 5314 6 n_333
rlabel m2contact 24511 3346 24511 3346 6 n_255
rlabel m2contact 24463 6514 24463 6514 6 n_128
rlabel m2contact 24463 2290 24463 2290 6 n_128
rlabel m2contact 24439 4930 24439 4930 6 n_114
rlabel m2contact 24415 3514 24415 3514 6 n_212
rlabel m2contact 24415 3538 24415 3538 6 n_274
rlabel m2contact 24391 2290 24391 2290 6 n_128
rlabel m2contact 24391 2386 24391 2386 6 n_50
rlabel m2contact 24343 5722 24343 5722 6 n_130
rlabel m2contact 24319 4594 24319 4594 6 LrSel
rlabel m2contact 24319 5866 24319 5866 6 stateSub[2]
rlabel m2contact 24295 3178 24295 3178 6 n_83
rlabel m2contact 24271 2578 24271 2578 6 n_272
rlabel m2contact 24247 6490 24247 6490 6 n_177
rlabel m2contact 24223 2674 24223 2674 6 OpcodeCondIn[2]
rlabel m2contact 24199 6850 24199 6850 6 n_157
rlabel m2contact 24175 3226 24175 3226 6 n_176
rlabel m2contact 24151 6946 24151 6946 6 n_151
rlabel m2contact 24127 7234 24127 7234 6 n_159
rlabel m2contact 24103 5506 24103 5506 6 n_116
rlabel m2contact 24103 3490 24103 3490 6 n_116
rlabel m2contact 24079 4378 24079 4378 6 n_173
rlabel m2contact 24055 3490 24055 3490 6 n_116
rlabel m2contact 24055 3514 24055 3514 6 n_212
rlabel m2contact 24031 7090 24031 7090 6 n_99
rlabel m2contact 24007 4978 24007 4978 6 n_60
rlabel m2contact 23983 2722 23983 2722 6 OpcodeCondIn[0]
rlabel m2contact 23959 2410 23959 2410 6 n_49
rlabel m2contact 23935 6370 23935 6370 6 n_154
rlabel m2contact 23911 4690 23911 4690 6 n_265
rlabel m2contact 23911 3538 23911 3538 6 n_274
rlabel m2contact 23863 6826 23863 6826 6 n_101
rlabel m2contact 23863 6274 23863 6274 6 n_39
rlabel m2contact 23839 6874 23839 6874 6 n_210
rlabel m2contact 23839 3418 23839 3418 6 OpcodeCondIn[4]
rlabel m2contact 23815 3682 23815 3682 6 n_186
rlabel m2contact 23791 4954 23791 4954 6 n_298
rlabel m2contact 23767 7162 23767 7162 6 n_238
rlabel m2contact 23767 6730 23767 6730 6 n_136
rlabel m2contact 23743 6658 23743 6658 6 n_267
rlabel m2contact 23695 2722 23695 2722 6 OpcodeCondIn[0]
rlabel m2contact 23671 5074 23671 5074 6 n_20
rlabel m2contact 23647 4330 23647 4330 6 n_297
rlabel m2contact 23623 6082 23623 6082 6 n_91
rlabel m2contact 23623 5098 23623 5098 6 n_217
rlabel m2contact 23599 6226 23599 6226 6 n_501
rlabel m2contact 23563 5122 23563 5122 6 n_88
rlabel m2contact 23563 3082 23563 3082 6 n_88
rlabel m2contact 23539 5698 23539 5698 6 n_194
rlabel m2contact 23539 3634 23539 3634 6 n_194
rlabel m2contact 23527 6514 23527 6514 6 n_128
rlabel m2contact 23527 2338 23527 2338 6 n_208
rlabel m2contact 23503 5338 23503 5338 6 n_104
rlabel m2contact 23503 2698 23503 2698 6 n_104
rlabel m2contact 23479 5122 23479 5122 6 n_88
rlabel m2contact 23479 5074 23479 5074 6 n_20
rlabel m2contact 23455 6826 23455 6826 6 n_101
rlabel m2contact 23455 4426 23455 4426 6 n_101
rlabel m2contact 23431 4210 23431 4210 6 n_11
rlabel m2contact 23407 3634 23407 3634 6 n_194
rlabel m2contact 23407 3682 23407 3682 6 n_186
rlabel m2contact 23383 3610 23383 3610 6 stateSub[1]
rlabel m2contact 23359 5458 23359 5458 6 n_362
rlabel m2contact 23335 2938 23335 2938 6 n_294
rlabel m2contact 23311 3994 23311 3994 6 n_105
rlabel m2contact 23287 2146 23287 2146 6 n_302
rlabel m2contact 23263 5338 23263 5338 6 n_104
rlabel m2contact 23263 5290 23263 5290 6 StatusReg[3]
rlabel m2contact 23239 2314 23239 2314 6 n_309
rlabel m2contact 23215 4594 23215 4594 6 n_19
rlabel m2contact 23191 4402 23191 4402 6 n_18
rlabel m2contact 23167 4426 23167 4426 6 n_101
rlabel m2contact 23167 5866 23167 5866 6 stateSub[2]
rlabel m2contact 23143 5098 23143 5098 6 n_217
rlabel m2contact 23095 5626 23095 5626 6 n_367
rlabel m2contact 23071 4162 23071 4162 6 state[0]
rlabel m2contact 23047 3322 23047 3322 6 state[1]
rlabel m2contact 22999 5146 22999 5146 6 n_259
rlabel m2contact 22999 7042 22999 7042 6 StatusReg[0]
rlabel m2contact 22951 6034 22951 6034 6 n_499
rlabel m2contact 22951 3514 22951 3514 6 n_212
rlabel m2contact 22855 5218 22855 5218 6 n_283
rlabel m2contact 22831 5146 22831 5146 6 n_259
rlabel m2contact 22807 3610 22807 3610 6 stateSub[1]
rlabel m2contact 22759 2770 22759 2770 6 n_96
rlabel m2contact 22735 3010 22735 3010 6 n_143
rlabel m2contact 22711 7090 22711 7090 6 n_99
rlabel m2contact 22663 2242 22663 2242 6 n_289
rlabel m2contact 22615 5242 22615 5242 6 n_275
rlabel m2contact 22615 3298 22615 3298 6 n_275
rlabel m2contact 22591 4066 22591 4066 6 n_381
rlabel m2contact 22567 4834 22567 4834 6 n_202
rlabel m2contact 22567 2170 22567 2170 6 n_202
rlabel m2contact 22543 6322 22543 6322 6 n_276
rlabel m2contact 22519 3538 22519 3538 6 n_274
rlabel m2contact 22495 3298 22495 3298 6 n_275
rlabel m2contact 22471 4786 22471 4786 6 n_342
rlabel m2contact 22471 3586 22471 3586 6 n_342
rlabel m2contact 22447 3298 22447 3298 6 n_275
rlabel m2contact 22447 3394 22447 3394 6 n_231
rlabel m2contact 22423 5266 22423 5266 6 n_87
rlabel m2contact 22423 4090 22423 4090 6 n_87
rlabel m2contact 22399 4834 22399 4834 6 n_202
rlabel m2contact 22399 4618 22399 4618 6 n_241
rlabel m2contact 22375 6418 22375 6418 6 n_266
rlabel m2contact 22351 4810 22351 4810 6 n_52
rlabel m2contact 22327 4786 22327 4786 6 n_342
rlabel m2contact 22327 3874 22327 3874 6 n_335
rlabel m2contact 22303 7138 22303 7138 6 n_17
rlabel m2contact 22303 5314 22303 5314 6 n_333
rlabel m2contact 22279 4786 22279 4786 6 SysBus[0]
rlabel m2contact 22255 2578 22255 2578 6 n_272
rlabel m2contact 22231 4666 22231 4666 6 n_234
rlabel m2contact 22207 4690 22207 4690 6 n_265
rlabel m2contact 22207 3538 22207 3538 6 n_274
rlabel m2contact 22183 2362 22183 2362 6 n_42
rlabel m2contact 22159 4234 22159 4234 6 n_182
rlabel m2contact 22135 6634 22135 6634 6 n_127
rlabel m2contact 22111 4738 22111 4738 6 n_153
rlabel m2contact 22111 4570 22111 4570 6 nWait
rlabel m2contact 22075 5122 22075 5122 6 n_37
rlabel m2contact 22075 4570 22075 4570 6 n_37
rlabel m2contact 22057 6418 22057 6418 6 n_266
rlabel m2contact 22051 4426 22051 4426 6 n_266
rlabel m2contact 22039 6418 22039 6418 6 n_266
rlabel m2contact 22015 4186 22015 4186 6 n_270
rlabel m2contact 21991 6874 21991 6874 6 n_210
rlabel m2contact 21991 2626 21991 2626 6 n_167
rlabel m2contact 21967 5050 21967 5050 6 n_5
rlabel m2contact 21967 1954 21967 1954 6 n_5
rlabel m2contact 21943 3514 21943 3514 6 n_212
rlabel m2contact 21919 5938 21919 5938 6 n_192
rlabel m2contact 21895 5098 21895 5098 6 n_217
rlabel m2contact 21871 4090 21871 4090 6 n_87
rlabel m2contact 21871 4162 21871 4162 6 state[0]
rlabel m2contact 21847 6778 21847 6778 6 n_163
rlabel m2contact 21847 5002 21847 5002 6 n_163
rlabel m2contact 21823 2218 21823 2218 6 n_38
rlabel m2contact 21799 2338 21799 2338 6 n_208
rlabel m2contact 21799 6274 21799 6274 6 n_39
rlabel m2contact 21775 5386 21775 5386 6 n_21
rlabel m2contact 21751 7186 21751 7186 6 n_313
rlabel m2contact 21751 3490 21751 3490 6 n_313
rlabel m2contact 21727 2602 21727 2602 6 n_220
rlabel m2contact 21703 6370 21703 6370 6 n_154
rlabel m2contact 21679 3250 21679 3250 6 n_279
rlabel m2contact 21679 4258 21679 4258 6 n_243
rlabel m2contact 21655 6970 21655 6970 6 n_339
rlabel m2contact 21631 6058 21631 6058 6 n_76
rlabel m2contact 21607 4330 21607 4330 6 n_297
rlabel m2contact 21583 4594 21583 4594 6 n_19
rlabel m2contact 21559 5122 21559 5122 6 n_37
rlabel m2contact 21559 4834 21559 4834 6 n_180
rlabel m2contact 21535 6010 21535 6010 6 n_261
rlabel m2contact 21511 3154 21511 3154 6 n_222
rlabel m2contact 21487 3802 21487 3802 6 n_264
rlabel m2contact 21463 6778 21463 6778 6 n_163
rlabel m2contact 21463 4474 21463 4474 6 OpcodeCondIn[6]
rlabel m2contact 21439 4426 21439 4426 6 n_266
rlabel m2contact 21439 4594 21439 4594 6 n_187
rlabel m2contact 21415 6274 21415 6274 6 n_39
rlabel m2contact 21391 5698 21391 5698 6 n_194
rlabel m2contact 21367 5050 21367 5050 6 n_5
rlabel m2contact 21367 4810 21367 4810 6 n_150
rlabel m2contact 21343 7234 21343 7234 6 n_159
rlabel m2contact 21319 6778 21319 6778 6 n_163
rlabel m2contact 21319 6730 21319 6730 6 n_136
rlabel m2contact 21295 4666 21295 4666 6 n_234
rlabel m2contact 21271 6106 21271 6106 6 n_318
rlabel m2contact 21247 4114 21247 4114 6 OpcodeCondIn[7]
rlabel m2contact 21223 3490 21223 3490 6 n_313
rlabel m2contact 21223 3562 21223 3562 6 n_317
rlabel m2contact 21199 5530 21199 5530 6 n_207
rlabel m2contact 21199 4330 21199 4330 6 n_207
rlabel m2contact 21175 5050 21175 5050 6 n_215
rlabel m2contact 21175 2458 21175 2458 6 n_215
rlabel m2contact 21151 3658 21151 3658 6 n_73
rlabel m2contact 21127 4738 21127 4738 6 n_82
rlabel m2contact 21127 1930 21127 1930 6 n_82
rlabel m2contact 21103 4330 21103 4330 6 n_207
rlabel m2contact 21103 4426 21103 4426 6 n_22
rlabel m2contact 21079 4258 21079 4258 6 n_243
rlabel m2contact 21055 5050 21055 5050 6 n_215
rlabel m2contact 21055 4666 21055 4666 6 n_234
rlabel m2contact 21031 5002 21031 5002 6 n_163
rlabel m2contact 21007 7234 21007 7234 6 n_159
rlabel m2contact 20983 4522 20983 4522 6 n_59
rlabel m2contact 20959 2938 20959 2938 6 n_294
rlabel m2contact 20935 4738 20935 4738 6 n_82
rlabel m2contact 20935 2962 20935 2962 6 n_178
rlabel m2contact 20911 4690 20911 4690 6 n_265
rlabel m2contact 20875 4738 20875 4738 6 n_89
rlabel m2contact 20875 2506 20875 2506 6 n_89
rlabel m2contact 20863 2338 20863 2338 6 n_208
rlabel m2contact 20839 4738 20839 4738 6 n_89
rlabel m2contact 20839 3706 20839 3706 6 n_144
rlabel m2contact 20791 4330 20791 4330 6 n_74
rlabel m2contact 20767 3610 20767 3610 6 stateSub[1]
rlabel m2contact 20743 3634 20743 3634 6 n_62
rlabel m2contact 20719 5026 20719 5026 6 n_224
rlabel m2contact 20695 3778 20695 3778 6 n_31
rlabel m2contact 20671 5098 20671 5098 6 n_217
rlabel m2contact 20647 3178 20647 3178 6 n_83
rlabel m2contact 20623 6346 20623 6346 6 n_25
rlabel m2contact 20599 4162 20599 4162 6 state[0]
rlabel m2contact 20551 4378 20551 4378 6 n_173
rlabel m2contact 20527 4546 20527 4546 6 n_100
rlabel m2contact 20527 5026 20527 5026 6 n_224
rlabel m2contact 20455 4738 20455 4738 6 n_354
rlabel m2contact 20431 4474 20431 4474 6 OpcodeCondIn[6]
rlabel m2contact 20407 4954 20407 4954 6 n_298
rlabel m2contact 20383 3418 20383 3418 6 OpcodeCondIn[4]
rlabel m2contact 20335 6682 20335 6682 6 n_156
rlabel m2contact 20311 3922 20311 3922 6 n_79
rlabel m2contact 20287 4546 20287 4546 6 n_137
rlabel m2contact 20215 2002 20215 2002 6 n_66
rlabel m2contact 20167 3178 20167 3178 6 n_83
rlabel m2contact 20119 5050 20119 5050 6 n_347
rlabel m2contact 20095 3202 20095 3202 6 n_122
rlabel m2contact 20071 2026 20071 2026 6 n_125
rlabel m2contact 19999 3058 19999 3058 6 n_68
rlabel m2contact 19975 5986 19975 5986 6 n_0
rlabel m2contact 19951 4474 19951 4474 6 OpcodeCondIn[6]
rlabel m2contact 19903 2074 19903 2074 6 n_345
rlabel m2contact 19879 6442 19879 6442 6 n_315
rlabel m2contact 19855 6898 19855 6898 6 n_296
rlabel m2contact 19807 4762 19807 4762 6 n_328
rlabel m2contact 19783 4786 19783 4786 6 SysBus[0]
rlabel m2contact 19735 5626 19735 5626 6 n_367
rlabel m2contact 19711 3106 19711 3106 6 n_237
rlabel m2contact 19687 6706 19687 6706 6 n_290
rlabel m2contact 19663 7114 19663 7114 6 n_41
rlabel m2contact 19639 7042 19639 7042 6 StatusReg[0]
rlabel m2contact 19591 5338 19591 5338 6 n_332
rlabel m2contact 19567 6370 19567 6370 6 n_154
rlabel m2contact 19543 7210 19543 7210 6 n_366
rlabel m2contact 19519 6610 19519 6610 6 OpcodeCondIn[5]
rlabel m2contact 19495 4954 19495 4954 6 n_263
rlabel m2contact 19495 2986 19495 2986 6 n_263
rlabel m2contact 19471 4954 19471 4954 6 n_263
rlabel m2contact 19471 4882 19471 4882 6 n_306
rlabel m2contact 19447 4690 19447 4690 6 n_265
rlabel m2contact 19423 5554 19423 5554 6 n_198
rlabel m2contact 19399 4690 19399 4690 6 n_324
rlabel m2contact 19375 4522 19375 4522 6 n_254
rlabel m2contact 19351 4954 19351 4954 6 n_45
rlabel m2contact 19351 6178 19351 6178 6 OpcodeCondIn[3]
rlabel m2contact 19327 6418 19327 6418 6 n_266
rlabel m2contact 19303 4114 19303 4114 6 OpcodeCondIn[7]
rlabel m2contact 19255 5938 19255 5938 6 n_192
rlabel m2contact 19231 5122 19231 5122 6 n_138
rlabel m2contact 19231 5170 19231 5170 6 n_58
rlabel m2contact 19207 3610 19207 3610 6 stateSub[1]
rlabel m2contact 19183 3898 19183 3898 6 n_81
rlabel m2contact 19159 4546 19159 4546 6 n_137
rlabel m2contact 19135 5434 19135 5434 6 n_271
rlabel m2contact 19111 3466 19111 3466 6 n_211
rlabel m2contact 19111 4186 19111 4186 6 n_270
rlabel m2contact 19087 5242 19087 5242 6 n_275
rlabel m2contact 19087 5218 19087 5218 6 n_283
rlabel m2contact 19063 6730 19063 6730 6 n_136
rlabel m2contact 19039 3442 19039 3442 6 n_250
rlabel m2contact 19015 4786 19015 4786 6 n_268
rlabel m2contact 19015 5002 19015 5002 6 n_77
rlabel m2contact 18991 2434 18991 2434 6 n_257
rlabel m2contact 18991 5194 18991 5194 6 n_278
rlabel m2contact 18967 6418 18967 6418 6 n_266
rlabel m2contact 18943 6802 18943 6802 6 n_200
rlabel m2contact 18919 5602 18919 5602 6 n_277
rlabel m2contact 18871 3946 18871 3946 6 n_321
rlabel m2contact 18847 3034 18847 3034 6 n_146
rlabel m2contact 18823 2842 18823 2842 6 n_147
rlabel m2contact 18751 5506 18751 5506 6 n_116
rlabel m2contact 18727 4306 18727 4306 6 CFlag
rlabel m2contact 18703 3586 18703 3586 6 n_342
rlabel m2contact 18655 2410 18655 2410 6 n_49
rlabel m2contact 18583 5218 18583 5218 6 n_283
rlabel m2contact 18511 3322 18511 3322 6 state[1]
rlabel m2contact 18487 4426 18487 4426 6 n_22
rlabel m2contact 18439 7066 18439 7066 6 n_54
rlabel m2contact 18391 4618 18391 4618 6 n_241
rlabel m2contact 18319 7258 18319 7258 6 n_380
rlabel m2contact 18319 7018 18319 7018 6 n_214
rlabel m2contact 18271 5242 18271 5242 6 n_174
rlabel m2contact 18247 3658 18247 3658 6 n_73
rlabel m2contact 18199 5818 18199 5818 6 n_158
rlabel m2contact 18175 5482 18175 5482 6 WdSel
rlabel m2contact 18175 3226 18175 3226 6 n_176
rlabel m2contact 18151 6850 18151 6850 6 n_157
rlabel m2contact 18127 4546 18127 4546 6 n_281
rlabel m2contact 18079 5338 18079 5338 6 n_332
rlabel m2contact 18079 5218 18079 5218 6 n_283
rlabel m2contact 18055 5314 18055 5314 6 n_333
rlabel m2contact 18031 6778 18031 6778 6 SysBus[2]
rlabel m2contact 18031 2674 18031 2674 6 OpcodeCondIn[2]
rlabel m2contact 17995 3490 17995 3490 6 n_90
rlabel m2contact 17995 2482 17995 2482 6 n_90
rlabel m2contact 17983 5482 17983 5482 6 n_35
rlabel m2contact 17959 2674 17959 2674 6 OpcodeCondIn[2]
rlabel m2contact 17935 2482 17935 2482 6 n_90
rlabel m2contact 17935 2650 17935 2650 6 n_34
rlabel m2contact 17911 5338 17911 5338 6 n_26
rlabel m2contact 17911 4378 17911 4378 6 n_173
rlabel m2contact 17887 5890 17887 5890 6 n_10
rlabel m2contact 17887 3298 17887 3298 6 n_10
rlabel m2contact 17863 7186 17863 7186 6 n_313
rlabel m2contact 17863 4354 17863 4354 6 n_111
rlabel m2contact 17839 3298 17839 3298 6 n_10
rlabel m2contact 17839 3634 17839 3634 6 n_62
rlabel m2contact 17815 2794 17815 2794 6 n_312
rlabel m2contact 17791 6370 17791 6370 6 n_154
rlabel m2contact 17791 2818 17791 2818 6 n_154
rlabel m2contact 17767 2794 17767 2794 6 n_312
rlabel m2contact 17743 3298 17743 3298 6 n_24
rlabel m2contact 17719 2818 17719 2818 6 n_154
rlabel m2contact 17719 3322 17719 3322 6 state[1]
rlabel m2contact 17695 7018 17695 7018 6 n_214
rlabel m2contact 17695 4618 17695 4618 6 n_241
rlabel m2contact 17671 7042 17671 7042 6 StatusReg[0]
rlabel m2contact 17671 4090 17671 4090 6 StatusReg[0]
rlabel m2contact 17647 2194 17647 2194 6 n_9
rlabel m2contact 17647 4018 17647 4018 6 n_352
rlabel m2contact 17623 7018 17623 7018 6 OpcodeCondIn[1]
rlabel m2contact 17599 4090 17599 4090 6 StatusReg[0]
rlabel m2contact 17599 4354 17599 4354 6 n_364
rlabel m2contact 17575 2722 17575 2722 6 OpcodeCondIn[0]
rlabel m2contact 17551 2290 17551 2290 6 n_386
rlabel m2contact 17479 2818 17479 2818 6 n_373
rlabel m2contact 17431 4282 17431 4282 6 n_400
rlabel m2contact 17431 5770 17431 5770 6 n_72
rlabel m2contact 17383 5098 17383 5098 6 n_217
rlabel m2contact 17359 4378 17359 4378 6 n_173
rlabel m2contact 17311 4042 17311 4042 6 n_44
rlabel m2contact 17287 7018 17287 7018 6 OpcodeCondIn[1]
rlabel m2contact 17263 2746 17263 2746 6 n_16
rlabel m2contact 17215 6970 17215 6970 6 n_339
rlabel m2contact 17167 2482 17167 2482 6 n_161
rlabel m2contact 17143 6922 17143 6922 6 n_251
rlabel m2contact 17095 2050 17095 2050 6 n_236
rlabel m2contact 17047 4162 17047 4162 6 state[0]
rlabel m2contact 17023 6970 17023 6970 6 n_181
rlabel m2contact 16975 4906 16975 4906 6 n_376
rlabel m2contact 16927 4786 16927 4786 6 n_268
rlabel m2contact 16903 4738 16903 4738 6 n_354
rlabel m2contact 16879 2458 16879 2458 6 n_215
rlabel m2contact 16843 4906 16843 4906 6 OpcodeCondIn[2]
rlabel m2contact 16843 2674 16843 2674 6 OpcodeCondIn[2]
rlabel m2contact 16831 6442 16831 6442 6 n_315
rlabel m2contact 16807 4738 16807 4738 6 n_188
rlabel m2contact 16783 5890 16783 5890 6 n_10
rlabel m2contact 16783 4786 16783 4786 6 n_303
rlabel m2contact 16759 6538 16759 6538 6 n_322
rlabel m2contact 16759 4090 16759 4090 6 n_322
rlabel m2contact 16735 4282 16735 4282 6 n_57
rlabel m2contact 16711 3298 16711 3298 6 n_24
rlabel m2contact 16687 6346 16687 6346 6 n_25
rlabel m2contact 16687 3994 16687 3994 6 n_105
rlabel m2contact 16663 2626 16663 2626 6 n_167
rlabel m2contact 16639 6082 16639 6082 6 n_91
rlabel m2contact 16615 4906 16615 4906 6 OpcodeCondIn[2]
rlabel m2contact 16615 3994 16615 3994 6 RwSel[1]
rlabel m2contact 16591 3490 16591 3490 6 n_90
rlabel m2contact 16567 3442 16567 3442 6 n_250
rlabel m2contact 16543 3946 16543 3946 6 n_321
rlabel m2contact 16519 4090 16519 4090 6 n_322
rlabel m2contact 16519 4786 16519 4786 6 n_303
rlabel m2contact 16447 3610 16447 3610 6 stateSub[1]
rlabel m2contact 16423 7162 16423 7162 6 n_238
rlabel m2contact 16423 7018 16423 7018 6 n_195
rlabel m2contact 16399 6178 16399 6178 6 OpcodeCondIn[3]
rlabel m2contact 16375 6418 16375 6418 6 n_266
rlabel m2contact 16375 4258 16375 4258 6 n_243
rlabel m2contact 16327 4906 16327 4906 6 n_349
rlabel m2contact 16303 2626 16303 2626 6 n_167
rlabel m2contact 16303 4090 16303 4090 6 n_145
rlabel m2contact 16279 3442 16279 3442 6 n_284
rlabel m2contact 16255 6322 16255 6322 6 n_276
rlabel m2contact 16231 6082 16231 6082 6 nME
rlabel m2contact 16231 1978 16231 1978 6 nME
rlabel m2contact 16207 6082 16207 6082 6 nME
rlabel m2contact 16207 4810 16207 4810 6 n_150
rlabel m2contact 16183 4378 16183 4378 6 n_173
rlabel m2contact 16159 4690 16159 4690 6 n_324
rlabel m2contact 16159 1978 16159 1978 6 nME
rlabel m2contact 16135 5626 16135 5626 6 n_367
rlabel m2contact 16111 4498 16111 4498 6 n_71
rlabel m2contact 16111 7162 16111 7162 6 n_47
rlabel m2contact 16087 4690 16087 4690 6 n_257
rlabel m2contact 16087 2434 16087 2434 6 n_257
rlabel m2contact 16063 6346 16063 6346 6 n_201
rlabel m2contact 16063 4114 16063 4114 6 OpcodeCondIn[7]
rlabel m2contact 16039 4690 16039 4690 6 n_257
rlabel m2contact 16039 3274 16039 3274 6 n_70
rlabel m2contact 16015 2266 16015 2266 6 n_190
rlabel m2contact 15991 6802 15991 6802 6 n_200
rlabel m2contact 15967 4498 15967 4498 6 n_346
rlabel m2contact 15943 2314 15943 2314 6 n_309
rlabel m2contact 15919 4690 15919 4690 6 n_227
rlabel m2contact 15895 5578 15895 5578 6 n_189
rlabel m2contact 15871 3466 15871 3466 6 n_211
rlabel m2contact 15847 7186 15847 7186 6 n_106
rlabel m2contact 15727 3226 15727 3226 6 n_176
rlabel m2contact 15703 5866 15703 5866 6 stateSub[2]
rlabel m2contact 15679 3034 15679 3034 6 n_146
rlabel m2contact 15655 4378 15655 4378 6 n_173
rlabel m2contact 15607 2026 15607 2026 6 n_125
rlabel m2contact 15559 5362 15559 5362 6 n_97
rlabel m2contact 15487 6874 15487 6874 6 n_210
rlabel m2contact 15463 2290 15463 2290 6 n_386
rlabel m2contact 15415 3922 15415 3922 6 n_79
rlabel m2contact 15391 5026 15391 5026 6 n_224
rlabel m2contact 15367 4594 15367 4594 6 n_187
rlabel m2contact 15319 5122 15319 5122 6 n_138
rlabel m2contact 15295 1978 15295 1978 6 n_377
rlabel m2contact 15271 4666 15271 4666 6 n_234
rlabel m2contact 15247 4594 15247 4594 6 n_187
rlabel m2contact 15223 6082 15223 6082 6 n_176
rlabel m2contact 15223 3226 15223 3226 6 n_176
rlabel m2contact 15199 6322 15199 6322 6 n_293
rlabel m2contact 15175 6538 15175 6538 6 n_322
rlabel m2contact 15175 5578 15175 5578 6 n_291
rlabel m2contact 15151 6082 15151 6082 6 n_176
rlabel m2contact 15151 3922 15151 3922 6 n_292
rlabel m2contact 15127 4594 15127 4594 6 n_187
rlabel m2contact 15103 5506 15103 5506 6 n_116
rlabel m2contact 15055 5506 15055 5506 6 n_85
rlabel m2contact 15007 5794 15007 5794 6 n_183
rlabel m2contact 14983 6034 14983 6034 6 n_499
rlabel m2contact 14959 3130 14959 3130 6 n_500
rlabel m2contact 14839 5290 14839 5290 6 StatusReg[3]
rlabel m2contact 14503 7162 14503 7162 4 n_47
rlabel m2contact 14503 3130 14503 3130 4 n_47
rlabel m2contact 14479 7258 14479 7258 4 n_42
rlabel m2contact 14479 2362 14479 2362 4 n_42
rlabel m2contact 14455 4402 14455 4402 4 n_18
rlabel m2contact 14431 3130 14431 3130 4 n_47
rlabel m2contact 14431 6922 14431 6922 4 n_378
rlabel m2contact 14407 6538 14407 6538 4 n_131
rlabel m2contact 14407 2290 14407 2290 4 n_131
rlabel m2contact 14383 3082 14383 3082 4 n_88
rlabel m2contact 14359 3274 14359 3274 4 n_70
rlabel m2contact 14335 6250 14335 6250 4 n_40
rlabel m2contact 14311 4954 14311 4954 4 n_45
rlabel m2contact 14287 3442 14287 3442 4 n_284
rlabel m2contact 14287 4114 14287 4114 4 OpcodeCondIn[7]
rlabel m2contact 14263 7258 14263 7258 4 n_42
rlabel m2contact 14263 6730 14263 6730 4 n_136
rlabel m2contact 14239 5194 14239 5194 4 n_278
rlabel m2contact 14215 5242 14215 5242 4 n_174
rlabel m2contact 14215 5218 14215 5218 4 n_283
rlabel m2contact 14191 6034 14191 6034 4 n_123
rlabel m2contact 14191 3442 14191 3442 4 n_123
rlabel m2contact 14167 3226 14167 3226 4 n_176
rlabel m2contact 14143 4378 14143 4378 4 n_173
rlabel m2contact 14119 3394 14119 3394 4 n_231
rlabel m2contact 14095 4282 14095 4282 4 n_57
rlabel m2contact 14095 4954 14095 4954 4 n_233
rlabel m2contact 14071 6538 14071 6538 4 n_131
rlabel m2contact 14071 6226 14071 6226 4 n_501
rlabel m2contact 14047 5242 14047 5242 4 n_199
rlabel m2contact 14023 6082 14023 6082 4 n_368
rlabel m2contact 13999 6034 13999 6034 4 n_123
rlabel m2contact 13999 5866 13999 5866 4 stateSub[2]
rlabel m2contact 13975 5938 13975 5938 4 n_192
rlabel m2contact 13975 3202 13975 3202 4 n_122
rlabel m2contact 13951 3010 13951 3010 4 n_143
rlabel m2contact 13927 6538 13927 6538 4 n_219
rlabel m2contact 13927 3394 13927 3394 4 n_219
rlabel m2contact 13903 6946 13903 6946 4 n_151
rlabel m2contact 13903 6730 13903 6730 4 n_136
rlabel m2contact 13879 4858 13879 4858 4 n_118
rlabel m2contact 13855 3418 13855 3418 4 OpcodeCondIn[4]
rlabel m2contact 13831 4810 13831 4810 4 n_150
rlabel m2contact 13831 4546 13831 4546 4 n_281
rlabel m2contact 13807 5866 13807 5866 4 stateSub[2]
rlabel m2contact 13807 1906 13807 1906 4 stateSub[2]
rlabel m2contact 13783 3394 13783 3394 4 n_219
rlabel m2contact 13783 4282 13783 4282 4 n_240
rlabel m2contact 13759 3034 13759 3034 4 n_146
rlabel m2contact 13735 6034 13735 6034 4 n_184
rlabel m2contact 13711 3394 13711 3394 4 n_6
rlabel m2contact 13687 3418 13687 3418 4 OpcodeCondIn[4]
rlabel m2contact 13687 3706 13687 3706 4 n_144
rlabel m2contact 13663 4114 13663 4114 4 OpcodeCondIn[7]
rlabel m2contact 13639 5746 13639 5746 4 n_160
rlabel m2contact 13615 7234 13615 7234 4 n_159
rlabel m2contact 13615 6946 13615 6946 4 n_93
rlabel m2contact 13591 4714 13591 4714 4 n_65
rlabel m2contact 13567 1906 13567 1906 4 stateSub[2]
rlabel m2contact 13567 3130 13567 3130 4 n_168
rlabel m2contact 13543 4114 13543 4114 4 OpcodeCondIn[7]
rlabel m2contact 13519 5938 13519 5938 4 n_192
rlabel m2contact 13495 5938 13495 5938 4 n_192
rlabel m2contact 13471 6706 13471 6706 4 n_290
rlabel m2contact 13471 4858 13471 4858 4 n_118
rlabel m2contact 13447 4714 13447 4714 4 n_228
rlabel m2contact 13423 1930 13423 1930 4 n_82
rlabel m2contact 13423 6442 13423 6442 4 n_315
rlabel m2contact 13399 3898 13399 3898 4 n_81
rlabel m2contact 13375 6850 13375 6850 4 n_157
rlabel m2contact 13375 5218 13375 5218 4 n_283
rlabel m2contact 13351 6706 13351 6706 4 n_68
rlabel m2contact 13351 3058 13351 3058 4 n_68
rlabel m2contact 13327 1954 13327 1954 4 n_5
rlabel m2contact 13327 4858 13327 4858 4 n_118
rlabel m2contact 13303 2674 13303 2674 4 OpcodeCondIn[2]
rlabel m2contact 13303 3466 13303 3466 4 n_211
rlabel m2contact 13279 6178 13279 6178 4 OpcodeCondIn[3]
rlabel m2contact 13255 6202 13255 6202 4 n_64
rlabel m2contact 13231 4570 13231 4570 4 n_37
rlabel m2contact 13207 6706 13207 6706 4 n_68
rlabel m2contact 13207 3754 13207 3754 4 stateSub[0]
rlabel m2contact 13183 6850 13183 6850 4 n_13
rlabel m2contact 13183 5770 13183 5770 4 n_72
rlabel m2contact 13135 7210 13135 7210 4 n_366
rlabel m2contact 13135 6706 13135 6706 4 Flags[2]
rlabel m2contact 13111 6706 13111 6706 4 Flags[2]
rlabel m2contact 13087 1978 13087 1978 4 n_377
rlabel m2contact 13087 4354 13087 4354 4 n_364
rlabel m2contact 13063 6082 13063 6082 4 n_368
rlabel m2contact 13039 2074 13039 2074 4 n_345
rlabel m2contact 13039 4570 13039 4570 4 n_204
rlabel m2contact 13015 6706 13015 6706 4 n_164
rlabel m2contact 12991 3442 12991 3442 4 n_123
rlabel m2contact 12967 5194 12967 5194 4 n_278
rlabel m2contact 12967 1978 12967 1978 4 n_278
rlabel m2contact 12943 7186 12943 7186 4 n_106
rlabel m2contact 12943 3442 12943 3442 4 n_252
rlabel m2contact 12919 2074 12919 2074 4 n_121
rlabel m2contact 12919 5266 12919 5266 4 n_87
rlabel m2contact 12895 1978 12895 1978 4 n_278
rlabel m2contact 12895 4378 12895 4378 4 n_173
rlabel m2contact 12823 5458 12823 5458 4 n_362
rlabel m2contact 12775 5458 12775 5458 4 n_348
rlabel m2contact 12775 4354 12775 4354 4 n_364
rlabel m2contact 12703 2434 12703 2434 4 n_257
rlabel m2contact 12679 3130 12679 3130 4 n_168
rlabel m2contact 12655 4114 12655 4114 4 OpcodeCondIn[7]
rlabel m2contact 12607 7162 12607 7162 4 n_47
rlabel m2contact 12607 6082 12607 6082 4 n_368
rlabel m2contact 12607 1978 12607 1978 4 n_368
rlabel m2contact 12583 1978 12583 1978 4 n_368
rlabel m2contact 12583 5026 12583 5026 4 n_224
rlabel m2contact 12559 2002 12559 2002 4 n_66
rlabel m2contact 12559 3322 12559 3322 4 state[1]
rlabel m2contact 12511 7138 12511 7138 4 n_17
rlabel m2contact 12511 6250 12511 6250 4 n_40
rlabel m2contact 12487 6178 12487 6178 4 OpcodeCondIn[3]
rlabel m2contact 12487 4114 12487 4114 4 OpcodeCondIn[7]
rlabel m2contact 12463 3058 12463 3058 4 n_68
rlabel m2contact 12463 4162 12463 4162 4 state[0]
rlabel m2contact 12439 3754 12439 3754 4 stateSub[0]
rlabel m2contact 12415 2434 12415 2434 4 n_257
rlabel m2contact 12391 3682 12391 3682 4 n_186
rlabel m2contact 12367 7114 12367 7114 4 n_41
rlabel m2contact 12367 6418 12367 6418 4 n_266
rlabel m2contact 12343 2434 12343 2434 4 n_257
rlabel m2contact 12343 4162 12343 4162 4 state[0]
rlabel m2contact 12319 3202 12319 3202 4 n_122
rlabel m2contact 12271 7090 12271 7090 4 n_99
rlabel m2contact 12247 5386 12247 5386 4 n_21
rlabel m2contact 12247 2434 12247 2434 4 n_21
rlabel m2contact 12223 5098 12223 5098 4 n_217
rlabel m2contact 12199 2434 12199 2434 4 n_21
rlabel m2contact 12199 3658 12199 3658 4 n_73
rlabel m2contact 12175 3418 12175 3418 4 OpcodeCondIn[4]
rlabel m2contact 12151 3058 12151 3058 4 n_68
rlabel m2contact 12151 4690 12151 4690 4 n_227
rlabel m2contact 12103 3946 12103 3946 4 n_321
rlabel m2contact 12103 5746 12103 5746 4 n_160
rlabel m2contact 12079 7066 12079 7066 4 n_54
rlabel m2contact 12079 3466 12079 3466 4 n_211
rlabel m2contact 12007 3898 12007 3898 4 n_81
rlabel m2contact 12007 7018 12007 7018 4 n_195
rlabel m2contact 11983 2650 11983 2650 4 n_34
rlabel m2contact 11959 4042 11959 4042 4 n_44
rlabel m2contact 11959 5698 11959 5698 4 n_194
rlabel m2contact 11911 3898 11911 3898 4 n_107
rlabel m2contact 11887 5746 11887 5746 4 n_160
rlabel m2contact 11863 4378 11863 4378 4 n_173
rlabel m2contact 11815 5698 11815 5698 4 n_139
rlabel m2contact 11791 3610 11791 3610 4 stateSub[1]
rlabel m2contact 11767 5122 11767 5122 4 n_138
rlabel m2contact 11743 3010 11743 3010 4 n_143
rlabel m2contact 11719 2026 11719 2026 4 n_125
rlabel m2contact 11719 2434 11719 2434 4 n_260
rlabel m2contact 11671 3778 11671 3778 4 n_31
rlabel m2contact 11647 5146 11647 5146 4 n_259
rlabel m2contact 11623 5122 11623 5122 4 n_8
rlabel m2contact 11599 2050 11599 2050 4 n_236
rlabel m2contact 11599 4042 11599 4042 4 n_311
rlabel m2contact 11575 7042 11575 7042 4 StatusReg[0]
rlabel m2contact 11575 7018 11575 7018 4 n_309
rlabel m2contact 11575 2314 11575 2314 4 n_309
rlabel m2contact 11551 7018 11551 7018 4 n_309
rlabel m2contact 11551 5146 11551 5146 4 n_56
rlabel m2contact 11527 3754 11527 3754 4 stateSub[0]
rlabel m2contact 11503 3658 11503 3658 4 n_73
rlabel m2contact 11479 2074 11479 2074 4 n_121
rlabel m2contact 11431 6994 11431 6994 4 n_94
rlabel m2contact 11431 6802 11431 6802 4 n_200
rlabel m2contact 11383 6970 11383 6970 4 n_181
rlabel m2contact 11383 6274 11383 6274 4 n_39
rlabel m2contact 11359 6514 11359 6514 4 n_128
rlabel m2contact 11335 4834 11335 4834 4 n_180
rlabel m2contact 11311 5530 11311 5530 4 n_207
rlabel m2contact 11287 4858 11287 4858 4 n_118
rlabel m2contact 11263 2338 11263 2338 4 n_208
rlabel m2contact 11263 5986 11263 5986 4 n_0
rlabel m2contact 11239 5098 11239 5098 4 n_217
rlabel m2contact 11215 6610 11215 6610 4 OpcodeCondIn[5]
rlabel m2contact 11215 2338 11215 2338 4 OpcodeCondIn[5]
rlabel m2contact 11191 5650 11191 5650 4 n_142
rlabel m2contact 11167 2338 11167 2338 4 OpcodeCondIn[5]
rlabel m2contact 11167 5986 11167 5986 4 n_230
rlabel m2contact 11143 6514 11143 6514 4 n_4
rlabel m2contact 11119 5650 11119 5650 4 n_169
rlabel m2contact 11095 2098 11095 2098 4 n_98
rlabel m2contact 11071 6946 11071 6946 4 n_93
rlabel m2contact 11071 2338 11071 2338 4 n_126
rlabel m2contact 11023 2122 11023 2122 4 n_110
rlabel m2contact 11023 6922 11023 6922 4 n_378
rlabel m2contact 10999 6562 10999 6562 4 n_331
rlabel m2contact 10975 2146 10975 2146 4 n_302
rlabel m2contact 10951 6562 10951 6562 4 n_365
rlabel m2contact 10903 6898 10903 6898 4 n_296
rlabel m2contact 10903 3946 10903 3946 4 n_321
rlabel m2contact 10879 5578 10879 5578 4 n_291
rlabel m2contact 10855 2170 10855 2170 4 n_202
rlabel m2contact 10855 3922 10855 3922 4 n_292
rlabel m2contact 10831 5098 10831 5098 4 n_217
rlabel m2contact 10783 5554 10783 5554 4 n_198
rlabel m2contact 10759 6754 10759 6754 4 n_46
rlabel m2contact 10735 5554 10735 5554 4 n_134
rlabel m2contact 10711 2194 10711 2194 4 n_9
rlabel m2contact 10687 2458 10687 2458 4 n_215
rlabel m2contact 10687 6754 10687 6754 4 n_27
rlabel m2contact 10639 6154 10639 6154 4 n_325
rlabel m2contact 10615 4666 10615 4666 4 n_234
rlabel m2contact 10567 3202 10567 3202 4 n_122
rlabel m2contact 10567 4978 10567 4978 4 n_60
rlabel m2contact 10543 3778 10543 3778 4 n_31
rlabel m2contact 10519 6874 10519 6874 4 n_210
rlabel m2contact 10519 3610 10519 3610 4 stateSub[1]
rlabel m2contact 10495 6610 10495 6610 4 OpcodeCondIn[5]
rlabel m2contact 10471 2626 10471 2626 4 n_167
rlabel m2contact 10447 6370 10447 6370 4 n_154
rlabel m2contact 10423 2458 10423 2458 4 n_113
rlabel m2contact 10423 3562 10423 3562 4 n_317
rlabel m2contact 10375 2674 10375 2674 4 OpcodeCondIn[2]
rlabel m2contact 10351 6586 10351 6586 4 n_244
rlabel m2contact 10327 2602 10327 2602 4 n_220
rlabel m2contact 10303 6850 10303 6850 4 n_13
rlabel m2contact 10303 6586 10303 6586 4 n_239
rlabel m2contact 10255 4114 10255 4114 4 OpcodeCondIn[7]
rlabel m2contact 10231 2602 10231 2602 4 n_14
rlabel m2contact 10183 6826 10183 6826 4 n_101
rlabel m2contact 10159 3538 10159 3538 4 n_274
rlabel m2contact 10135 6802 10135 6802 4 n_200
rlabel m2contact 10111 5842 10111 5842 4 SysBus[1]
rlabel m2contact 10087 2698 10087 2698 4 n_104
rlabel m2contact 10039 6802 10039 6802 4 n_7
rlabel m2contact 10039 3106 10039 3106 4 n_237
rlabel m2contact 10015 6298 10015 6298 4 n_80
rlabel m2contact 9967 4306 9967 4306 4 CFlag
rlabel m2contact 9943 5050 9943 5050 4 n_347
rlabel m2contact 9919 5842 9919 5842 4 n_357
rlabel m2contact 9895 2218 9895 2218 4 n_38
rlabel m2contact 9895 2242 9895 2242 4 n_289
rlabel m2contact 9871 2266 9871 2266 4 n_190
rlabel m2contact 9871 4306 9871 4306 4 n_269
rlabel m2contact 9823 6802 9823 6802 4 n_7
rlabel m2contact 9799 6778 9799 6778 4 SysBus[2]
rlabel m2contact 9775 4114 9775 4114 4 OpcodeCondIn[7]
rlabel m2contact 9751 4618 9751 4618 4 n_241
rlabel m2contact 9727 3106 9727 3106 4 n_237
rlabel m2contact 9703 5314 9703 5314 4 n_333
rlabel m2contact 9679 6778 9679 6778 4 OpcodeCondIn[2]
rlabel m2contact 9679 2674 9679 2674 4 OpcodeCondIn[2]
rlabel m2contact 9655 6778 9655 6778 4 OpcodeCondIn[2]
rlabel m2contact 9655 5314 9655 5314 4 StatusReg[2]
rlabel m2contact 9631 5602 9631 5602 4 n_277
rlabel m2contact 9583 6514 9583 6514 4 n_4
rlabel m2contact 9583 5314 9583 5314 4 StatusReg[2]
rlabel m2contact 9559 2314 9559 2314 4 n_309
rlabel m2contact 9559 4474 9559 4474 4 OpcodeCondIn[6]
rlabel m2contact 9535 3754 9535 3754 4 stateSub[0]
rlabel m2contact 9511 6514 9511 6514 4 n_95
rlabel m2contact 9487 4330 9487 4330 4 n_74
rlabel m2contact 9451 5722 9451 5722 4 n_130
rlabel m2contact 9451 2314 9451 2314 4 n_130
rlabel m2contact 9439 5770 9439 5770 4 n_72
rlabel m2contact 9415 2290 9415 2290 4 n_131
rlabel m2contact 9415 3658 9415 3658 4 n_73
rlabel m2contact 9391 3322 9391 3322 4 state[1]
rlabel m2contact 9367 2314 9367 2314 4 n_130
rlabel m2contact 9367 4330 9367 4330 4 n_172
rlabel m2contact 9343 2338 9343 2338 4 n_126
rlabel m2contact 9319 2626 9319 2626 4 n_167
rlabel m2contact 9271 2482 9271 2482 4 n_161
rlabel m2contact 9247 5746 9247 5746 4 n_160
rlabel m2contact 9223 2626 9223 2626 4 n_167
rlabel m2contact 9199 2482 9199 2482 4 n_32
rlabel m2contact 9175 6754 9175 6754 4 n_27
rlabel m2contact 9175 3778 9175 3778 4 n_31
rlabel m2contact 9151 2362 9151 2362 4 n_42
rlabel m2contact 9151 6730 9151 6730 4 n_136
rlabel m2contact 9127 5338 9127 5338 4 n_26
rlabel m2contact 9079 3490 9079 3490 4 n_90
rlabel m2contact 9031 3058 9031 3058 4 n_68
rlabel m2contact 9007 3490 9007 3490 4 n_69
rlabel m2contact 8959 2386 8959 2386 4 n_50
rlabel m2contact 8959 6706 8959 6706 4 n_164
rlabel m2contact 8935 3226 8935 3226 4 n_176
rlabel m2contact 8911 3202 8911 3202 4 n_122
rlabel m2contact 8863 3226 8863 3226 4 n_206
rlabel m2contact 8863 2722 8863 2722 4 OpcodeCondIn[0]
rlabel m2contact 8839 2410 8839 2410 4 n_49
rlabel m2contact 8815 5530 8815 5530 4 n_207
rlabel m2contact 8791 6682 8791 6682 4 n_156
rlabel m2contact 8791 5842 8791 5842 4 n_357
rlabel m2contact 8743 2434 8743 2434 4 n_260
rlabel m2contact 8743 6658 8743 6658 4 n_267
rlabel m2contact 8719 3226 8719 3226 4 n_206
rlabel m2contact 8719 5218 8719 5218 4 n_283
rlabel m2contact 8695 6418 8695 6418 4 n_266
rlabel m2contact 8671 3226 8671 3226 4 n_23
rlabel m2contact 8623 2650 8623 2650 4 n_34
rlabel m2contact 8599 2722 8599 2722 4 OpcodeCondIn[0]
rlabel m2contact 8575 2602 8575 2602 4 n_14
rlabel m2contact 8527 2458 8527 2458 4 n_113
rlabel m2contact 8503 4210 8503 4210 4 n_11
rlabel m2contact 8479 2482 8479 2482 4 n_32
rlabel m2contact 8455 4210 8455 4210 4 n_61
rlabel m2contact 8407 6634 8407 6634 4 n_127
rlabel m2contact 8383 5026 8383 5026 4 n_224
rlabel m2contact 8359 2506 8359 2506 4 n_89
rlabel m2contact 8311 6538 8311 6538 4 n_219
rlabel m2contact 8263 2674 8263 2674 4 OpcodeCondIn[2]
rlabel m2contact 8239 5818 8239 5818 4 n_158
rlabel m2contact 8215 6538 8215 6538 4 n_235
rlabel m2contact 8215 2506 8215 2506 4 n_235
rlabel m2contact 8191 5818 8191 5818 4 n_205
rlabel m2contact 8167 2506 8167 2506 4 n_235
rlabel m2contact 8167 5746 8167 5746 4 n_160
rlabel m2contact 8143 4258 8143 4258 4 n_243
rlabel m2contact 8071 5674 8071 5674 4 n_363
rlabel m2contact 8023 4906 8023 4906 4 n_349
rlabel m2contact 8023 4618 8023 4618 4 n_241
rlabel m2contact 7999 4186 7999 4186 4 n_270
rlabel m2contact 7975 4906 7975 4906 4 n_30
rlabel m2contact 7951 2530 7951 2530 4 n_108
rlabel m2contact 7951 6610 7951 6610 4 OpcodeCondIn[5]
rlabel m2contact 7927 6250 7927 6250 4 n_40
rlabel m2contact 7927 4618 7927 4618 4 n_241
rlabel m2contact 7903 4666 7903 4666 4 n_234
rlabel m2contact 7879 6610 7879 6610 4 OpcodeCondIn[5]
rlabel m2contact 7879 5674 7879 5674 4 n_355
rlabel m2contact 7879 2530 7879 2530 4 n_355
rlabel m2contact 7855 4666 7855 4666 4 n_375
rlabel m2contact 7831 6586 7831 6586 4 n_239
rlabel m2contact 7831 3610 7831 3610 4 stateSub[1]
rlabel m2contact 7807 2530 7807 2530 4 n_355
rlabel m2contact 7807 3418 7807 3418 4 OpcodeCondIn[4]
rlabel m2contact 7783 6418 7783 6418 4 n_266
rlabel m2contact 7759 3922 7759 3922 4 n_292
rlabel m2contact 7735 6562 7735 6562 4 n_365
rlabel m2contact 7711 3922 7711 3922 4 Flags[3]
rlabel m2contact 7687 4354 7687 4354 4 n_364
rlabel m2contact 7639 6538 7639 6538 4 n_235
rlabel m2contact 7639 2554 7639 2554 4 LrWe
rlabel m2contact 7615 6514 7615 6514 4 n_95
rlabel m2contact 7615 6490 7615 6490 4 n_177
rlabel m2contact 7591 2578 7591 2578 4 n_272
rlabel m2contact 7591 6466 7591 6466 4 n_86
rlabel m2contact 7567 4738 7567 4738 4 n_188
rlabel m2contact 7519 3010 7519 3010 4 n_143
rlabel m2contact 7519 4738 7519 4738 4 n_336
rlabel m2contact 7495 5218 7495 5218 4 n_283
rlabel m2contact 7471 5602 7471 5602 4 n_277
rlabel m2contact 7471 3634 7471 3634 4 n_62
rlabel m2contact 7423 5602 7423 5602 4 n_316
rlabel m2contact 7399 6442 7399 6442 4 n_315
rlabel m2contact 7399 2674 7399 2674 4 OpcodeCondIn[2]
rlabel m2contact 7375 6322 7375 6322 4 n_293
rlabel m2contact 7375 5866 7375 5866 4 stateSub[2]
rlabel m2contact 7351 2602 7351 2602 4 n_14
rlabel m2contact 7327 6322 7327 6322 4 n_253
rlabel m2contact 7327 3538 7327 3538 4 n_274
rlabel m2contact 7303 6178 7303 6178 4 OpcodeCondIn[3]
rlabel m2contact 7279 6418 7279 6418 4 n_266
rlabel m2contact 7255 5410 7255 5410 4 n_109
rlabel m2contact 7255 3274 7255 3274 4 n_70
rlabel m2contact 7231 2626 7231 2626 4 n_167
rlabel m2contact 7207 6394 7207 6394 4 n_124
rlabel m2contact 7183 5866 7183 5866 4 stateSub[2]
rlabel m2contact 7159 3226 7159 3226 4 n_23
rlabel m2contact 7159 3466 7159 3466 4 n_211
rlabel m2contact 7111 2650 7111 2650 4 n_34
rlabel m2contact 7111 3226 7111 3226 4 n_135
rlabel m2contact 7087 6370 7087 6370 4 n_154
rlabel m2contact 7063 5866 7063 5866 4 stateSub[2]
rlabel m2contact 7063 4594 7063 4594 4 n_187
rlabel m2contact 7039 2698 7039 2698 4 n_104
rlabel m2contact 7015 3514 7015 3514 4 n_212
rlabel m2contact 6991 4858 6991 4858 4 n_118
rlabel m2contact 6967 6346 6967 6346 4 n_201
rlabel m2contact 6943 2698 6943 2698 4 n_314
rlabel m2contact 6919 2674 6919 2674 4 OpcodeCondIn[2]
rlabel m2contact 6919 6322 6919 6322 4 n_253
rlabel m2contact 6895 3154 6895 3154 4 n_222
rlabel m2contact 6871 3610 6871 3610 4 stateSub[1]
rlabel m2contact 6847 3490 6847 3490 4 n_69
rlabel m2contact 6823 2698 6823 2698 4 n_314
rlabel m2contact 6823 6322 6823 6322 4 n_122
rlabel m2contact 6823 3202 6823 3202 4 n_122
rlabel m2contact 6799 6322 6799 6322 4 n_122
rlabel m2contact 6799 4186 6799 4186 4 n_270
rlabel m2contact 6751 6298 6751 6298 4 n_80
rlabel m2contact 6727 6274 6727 6274 4 n_39
rlabel m2contact 6703 6250 6703 6250 4 n_40
rlabel m2contact 6703 2746 6703 2746 4 n_16
rlabel m2contact 6655 2722 6655 2722 4 OpcodeCondIn[0]
rlabel m2contact 6655 2746 6655 2746 4 AluOR[1]
rlabel m2contact 6607 6226 6607 6226 4 n_501
rlabel m2contact 6607 2746 6607 2746 4 AluOR[1]
rlabel m2contact 6583 6202 6583 6202 4 n_64
rlabel m2contact 6583 4882 6583 4882 4 n_306
rlabel m2contact 6559 3610 6559 3610 4 stateSub[1]
rlabel m2contact 6535 3946 6535 3946 4 n_321
rlabel m2contact 6535 4378 6535 4378 4 n_173
rlabel m2contact 6487 4858 6487 4858 4 n_118
rlabel m2contact 6439 6178 6439 6178 4 OpcodeCondIn[3]
rlabel m2contact 6439 5098 6439 5098 4 n_217
rlabel m2contact 6415 4378 6415 4378 4 n_173
rlabel m2contact 6391 4858 6391 4858 4 n_343
rlabel m2contact 6391 2746 6391 2746 4 n_343
rlabel m2contact 6367 2746 6367 2746 4 n_343
rlabel m2contact 6367 3946 6367 3946 4 ALE
rlabel m2contact 6343 2770 6343 2770 4 n_96
rlabel m2contact 6319 6154 6319 6154 4 n_325
rlabel m2contact 6319 2794 6319 2794 4 n_312
rlabel m2contact 6295 3970 6295 3970 4 n_120
rlabel m2contact 6247 2818 6247 2818 4 n_373
rlabel m2contact 6247 3970 6247 3970 4 Rs1Sel[0]
rlabel m2contact 6223 2842 6223 2842 4 n_147
rlabel m2contact 6223 5626 6223 5626 4 n_367
rlabel m2contact 6199 6130 6199 6130 4 n_320
rlabel m2contact 6199 6106 6199 6106 4 n_318
rlabel m2contact 6175 2866 6175 2866 4 n_249
rlabel m2contact 6151 6082 6151 6082 4 n_368
rlabel m2contact 6103 2890 6103 2890 4 n_390
rlabel m2contact 6079 2914 6079 2914 4 Op1Sel
rlabel m2contact 6079 3586 6079 3586 4 n_342
rlabel m2contact 6055 4666 6055 4666 4 n_375
rlabel m2contact 6031 6058 6031 6058 4 n_76
rlabel m2contact 6031 2938 6031 2938 4 n_294
rlabel m2contact 6007 4666 6007 4666 4 n_63
rlabel m2contact 5983 6034 5983 6034 4 n_184
rlabel m2contact 5959 5530 5959 5530 4 n_207
rlabel m2contact 5935 6010 5935 6010 4 n_261
rlabel m2contact 5935 5794 5935 5794 4 n_183
rlabel m2contact 5887 5986 5887 5986 4 n_230
rlabel m2contact 5887 5794 5887 5794 4 PcSel[0]
rlabel m2contact 5863 4786 5863 4786 4 n_303
rlabel m2contact 5839 5962 5839 5962 4 n_132
rlabel m2contact 5839 2986 5839 2986 4 n_263
rlabel m2contact 5815 5938 5815 5938 4 n_192
rlabel m2contact 5791 4138 5791 4138 4 n_51
rlabel m2contact 5791 2986 5791 2986 4 Flags[1]
rlabel m2contact 5743 5794 5743 5794 4 PcSel[0]
rlabel m2contact 5671 5530 5671 5530 4 n_207
rlabel m2contact 5647 5314 5647 5314 4 StatusReg[2]
rlabel m2contact 5623 3130 5623 3130 4 n_168
rlabel m2contact 5575 4138 5575 4138 4 nWE
rlabel m2contact 5551 5146 5551 5146 4 n_56
rlabel m2contact 5527 4858 5527 4858 4 n_343
rlabel m2contact 5503 5146 5503 5146 4 n_256
rlabel m2contact 5431 2962 5431 2962 4 n_178
rlabel m2contact 5407 5794 5407 5794 4 n_112
rlabel m2contact 5359 5362 5359 5362 4 n_97
rlabel m2contact 5335 5026 5335 5026 4 n_224
rlabel m2contact 5263 5914 5263 5914 4 n_351
rlabel m2contact 5239 2986 5239 2986 4 Flags[1]
rlabel m2contact 5215 4354 5215 4354 4 n_364
rlabel m2contact 5167 5890 5167 5890 4 n_10
rlabel m2contact 5143 4162 5143 4162 4 state[0]
rlabel m2contact 5119 5866 5119 5866 4 stateSub[2]
rlabel m2contact 5119 4090 5119 4090 4 n_145
rlabel m2contact 5095 3010 5095 3010 4 n_143
rlabel m2contact 5071 3706 5071 3706 4 n_144
rlabel m2contact 5071 4090 5071 4090 4 Rs1Sel[1]
rlabel m2contact 5047 4882 5047 4882 4 n_306
rlabel m2contact 5023 5842 5023 5842 4 n_357
rlabel m2contact 5023 3034 5023 3034 4 n_146
rlabel m2contact 4999 3058 4999 3058 4 n_68
rlabel m2contact 4999 4882 4999 4882 4 n_301
rlabel m2contact 4975 5818 4975 5818 4 n_205
rlabel m2contact 4975 5746 4975 5746 4 n_160
rlabel m2contact 4927 5794 4927 5794 4 n_112
rlabel m2contact 4903 3682 4903 3682 4 n_186
rlabel m2contact 4879 5770 4879 5770 4 n_72
rlabel m2contact 4879 3082 4879 3082 4 n_88
rlabel m2contact 4855 5746 4855 5746 4 n_160
rlabel m2contact 4807 3106 4807 3106 4 n_237
rlabel m2contact 4759 3130 4759 3130 4 n_168
rlabel m2contact 4759 5098 4759 5098 4 n_217
rlabel m2contact 4735 5722 4735 5722 4 n_130
rlabel m2contact 4735 5698 4735 5698 4 n_139
rlabel m2contact 4687 5674 4687 5674 4 n_355
rlabel m2contact 4687 5650 4687 5650 4 n_169
rlabel m2contact 4663 5626 4663 5626 4 n_367
rlabel m2contact 4663 3610 4663 3610 4 stateSub[1]
rlabel m2contact 4639 5602 4639 5602 4 n_316
rlabel m2contact 4591 5578 4591 5578 4 n_291
rlabel m2contact 4591 5554 4591 5554 4 n_134
rlabel m2contact 4567 3682 4567 3682 4 n_186
rlabel m2contact 4543 5530 4543 5530 4 n_207
rlabel m2contact 4543 5506 4543 5506 4 n_85
rlabel m2contact 4519 5482 4519 5482 4 n_35
rlabel m2contact 4495 5458 4495 5458 4 n_348
rlabel m2contact 4471 5050 4471 5050 4 n_347
rlabel m2contact 4447 5434 4447 5434 4 n_271
rlabel m2contact 4447 5218 4447 5218 4 n_283
rlabel m2contact 4423 3154 4423 3154 4 n_222
rlabel m2contact 4423 5050 4423 5050 4 n_225
rlabel m2contact 4399 3754 4399 3754 4 stateSub[0]
rlabel m2contact 4351 5410 4351 5410 4 n_109
rlabel m2contact 4327 3490 4327 3490 4 n_69
rlabel m2contact 4303 5386 4303 5386 4 n_21
rlabel m2contact 4303 3658 4303 3658 4 n_73
rlabel m2contact 4255 5362 4255 5362 4 n_97
rlabel m2contact 4231 3322 4231 3322 4 state[1]
rlabel m2contact 4207 3658 4207 3658 4 n_73
rlabel m2contact 4135 5338 4135 5338 4 n_26
rlabel m2contact 4135 3178 4135 3178 4 n_83
rlabel m2contact 4087 4162 4087 4162 4 state[0]
rlabel m2contact 4063 3202 4063 3202 4 n_122
rlabel m2contact 4039 5314 4039 5314 4 StatusReg[2]
rlabel m2contact 4015 5290 4015 5290 4 StatusReg[3]
rlabel m2contact 4015 5242 4015 5242 4 n_199
rlabel m2contact 3991 4162 3991 4162 4 state[0]
rlabel m2contact 3967 5266 3967 5266 4 n_87
rlabel m2contact 3967 5242 3967 5242 4 n_70
rlabel m2contact 3967 3274 3967 3274 4 n_70
rlabel m2contact 3943 3226 3943 3226 4 n_135
rlabel m2contact 3943 4474 3943 4474 4 OpcodeCondIn[6]
rlabel m2contact 3919 5242 3919 5242 4 n_70
rlabel m2contact 3919 3490 3919 3490 4 n_69
rlabel m2contact 3871 3250 3871 3250 4 n_279
rlabel m2contact 3847 5218 3847 5218 4 n_283
rlabel m2contact 3847 3274 3847 3274 4 n_70
rlabel m2contact 3823 5194 3823 5194 4 n_278
rlabel m2contact 3799 5170 3799 5170 4 n_58
rlabel m2contact 3799 3298 3799 3298 4 n_24
rlabel m2contact 3751 5146 3751 5146 4 n_256
rlabel m2contact 3727 5026 3727 5026 4 n_224
rlabel m2contact 3703 3346 3703 3346 4 n_255
rlabel m2contact 3655 5122 3655 5122 4 n_8
rlabel m2contact 3655 3322 3655 3322 4 state[1]
rlabel m2contact 3631 5098 3631 5098 4 n_217
rlabel m2contact 3631 3346 3631 3346 4 n_217
rlabel m2contact 3607 3346 3607 3346 4 n_217
rlabel m2contact 3607 3778 3607 3778 4 n_31
rlabel m2contact 3583 5098 3583 5098 4 n_217
rlabel m2contact 3535 5074 3535 5074 4 n_20
rlabel m2contact 3511 5026 3511 5026 4 n_224
rlabel m2contact 3487 3754 3487 3754 4 stateSub[0]
rlabel m2contact 3439 5050 3439 5050 4 n_225
rlabel m2contact 3415 5026 3415 5026 4 n_224
rlabel m2contact 3391 3850 3391 3850 4 n_218
rlabel m2contact 3367 3514 3367 3514 4 n_212
rlabel m2contact 3319 5002 3319 5002 4 n_77
rlabel m2contact 3295 4114 3295 4114 4 OpcodeCondIn[7]
rlabel m2contact 3271 4978 3271 4978 4 n_60
rlabel m2contact 3247 4954 3247 4954 4 n_233
rlabel m2contact 3223 3370 3223 3370 4 n_179
rlabel m2contact 3199 3394 3199 3394 4 n_6
rlabel m2contact 3175 4930 3175 4930 4 n_114
rlabel m2contact 3151 4906 3151 4906 4 n_30
rlabel m2contact 3103 4882 3103 4882 4 n_301
rlabel m2contact 3103 4618 3103 4618 4 n_241
rlabel m2contact 3055 3418 3055 3418 4 OpcodeCondIn[4]
rlabel m2contact 3055 4618 3055 4618 4 n_248
rlabel m2contact 3031 3442 3031 3442 4 n_252
rlabel m2contact 2983 4738 2983 4738 4 n_336
rlabel m2contact 2935 3586 2935 3586 4 n_342
rlabel m2contact 2911 4858 2911 4858 4 n_343
rlabel m2contact 2911 3466 2911 3466 4 n_211
rlabel m2contact 2863 4834 2863 4834 4 n_180
rlabel m2contact 2863 3490 2863 3490 4 n_69
rlabel m2contact 2839 3514 2839 3514 4 n_212
rlabel m2contact 2839 4114 2839 4114 4 OpcodeCondIn[7]
rlabel m2contact 2815 3610 2815 3610 4 stateSub[1]
rlabel m2contact 2791 4810 2791 4810 4 n_150
rlabel m2contact 2767 3538 2767 3538 4 n_274
rlabel m2contact 2743 3562 2743 3562 4 n_317
rlabel m2contact 2719 4786 2719 4786 4 n_303
rlabel m2contact 2695 4762 2695 4762 4 n_328
rlabel m2contact 2695 3586 2695 3586 4 n_342
rlabel m2contact 2671 4738 2671 4738 4 n_336
rlabel m2contact 2671 3754 2671 3754 4 stateSub[0]
rlabel m2contact 2647 3610 2647 3610 4 stateSub[1]
rlabel m2contact 2623 4714 2623 4714 4 n_228
rlabel m2contact 2599 4690 2599 4690 4 n_227
rlabel m2contact 2599 4666 2599 4666 4 n_63
rlabel m2contact 2575 4642 2575 4642 4 n_193
rlabel m2contact 2575 3634 2575 3634 4 n_62
rlabel m2contact 2551 3658 2551 3658 4 n_73
rlabel m2contact 2527 4618 2527 4618 4 n_248
rlabel m2contact 2503 4594 2503 4594 4 n_187
rlabel m2contact 2479 4570 2479 4570 4 n_204
rlabel m2contact 2479 3682 2479 3682 4 n_186
rlabel m2contact 2455 3706 2455 3706 4 n_144
rlabel m2contact 2431 3730 2431 3730 4 n_374
rlabel m2contact 2407 4546 2407 4546 4 n_281
rlabel m2contact 2383 4498 2383 4498 4 n_346
rlabel m2contact 2359 4522 2359 4522 4 n_254
rlabel m2contact 2335 4498 2335 4498 4 n_226
rlabel m2contact 2311 3754 2311 3754 4 stateSub[0]
rlabel m2contact 2287 4498 2287 4498 4 n_226
rlabel m2contact 2263 4474 2263 4474 4 OpcodeCondIn[6]
rlabel m2contact 2263 3778 2263 3778 4 n_31
rlabel m2contact 2239 4258 2239 4258 4 n_243
rlabel m2contact 2215 4450 2215 4450 4 n_152
rlabel m2contact 2167 4426 2167 4426 4 n_22
rlabel m2contact 2143 4402 2143 4402 4 n_18
rlabel m2contact 2119 4378 2119 4378 4 n_173
rlabel m2contact 2071 4354 2071 4354 4 n_364
rlabel m2contact 2047 4330 2047 4330 4 n_172
rlabel m2contact 2023 3802 2023 3802 4 n_264
rlabel m2contact 1999 3826 1999 3826 4 n_191
rlabel m2contact 1951 4306 1951 4306 4 n_269
rlabel m2contact 1927 4282 1927 4282 4 n_240
rlabel m2contact 1903 4258 1903 4258 4 n_243
rlabel m2contact 1903 4234 1903 4234 4 n_182
rlabel m2contact 1855 4210 1855 4210 4 n_61
rlabel m2contact 1831 4186 1831 4186 4 n_270
rlabel m2contact 1807 4162 1807 4162 4 state[0]
rlabel m2contact 1783 4138 1783 4138 4 nWE
rlabel m2contact 1759 4114 1759 4114 4 OpcodeCondIn[7]
rlabel m2contact 1735 4090 1735 4090 4 Rs1Sel[1]
rlabel m2contact 1711 4066 1711 4066 4 n_381
rlabel m2contact 1687 3850 1687 3850 4 n_218
rlabel m2contact 1687 3874 1687 3874 4 n_335
rlabel m2contact 1663 3898 1663 3898 4 n_107
rlabel m2contact 1663 4042 1663 4042 4 n_311
rlabel m2contact 1639 4018 1639 4018 4 n_352
rlabel metal2 26749 8252 26761 8252 6 LrSel
rlabel metal2 23521 8252 23533 8252 6 OpcodeCondIn[4]
rlabel metal2 21337 8252 21349 8252 6 Op2Sel[0]
rlabel metal2 19153 8252 19165 8252 6 OpcodeCondIn[2]
rlabel metal2 18037 8252 18049 8252 6 SysBus[2]
rlabel metal2 14785 8252 14797 8252 6 OpcodeCondIn[0]
rlabel metal2 12601 8252 12613 8252 4 PcSel[1]
rlabel metal2 12565 8252 12577 8252 4 RwSel[0]
rlabel metal2 10369 8252 10381 8252 4 nIRQ
rlabel metal2 6661 8252 6673 8252 4 AluOR[1]
rlabel metal2 3817 8252 3829 8252 4 ENB
rlabel metal2 3781 8252 3793 8252 4 SysBus[1]
rlabel metal2 25573 0 25585 0 8 IrWe
rlabel metal2 23401 0 23413 0 8 OpcodeCondIn[3]
rlabel metal2 21229 0 21241 0 8 OpcodeCondIn[1]
rlabel metal2 19057 0 19069 0 8 PcWe
rlabel metal2 16885 0 16897 0 8 Flags[1]
rlabel metal2 14713 0 14725 0 8 RegWe
rlabel metal2 14689 0 14701 0 8 nME
rlabel metal2 10357 0 10369 0 2 PcEn
rlabel metal2 9973 0 9985 0 2 CFlag
rlabel metal2 8137 0 8149 0 2 ImmSel
rlabel metal2 5953 0 5965 0 2 AluOR[0]
rlabel metal2 3769 0 3781 0 2 nOE
rlabel metal2 28280 8085 28280 8097 6 SysBus[3]
rlabel metal2 28280 8109 28280 8121 6 Flags[0]
rlabel metal2 28280 8133 28280 8145 6 SysBus[0]
rlabel metal2 28280 8205 28280 8217 6 PcSel[2]
rlabel metal2 28280 1900 28280 1912 6 AluWe
rlabel metal2 28280 1924 28280 1936 6 Op1Sel
rlabel metal2 28280 2548 28280 2560 6 LrWe
rlabel metal2 28280 5476 28280 5488 6 WdSel
rlabel metal2 28280 539 28280 551 8 AluEn
rlabel metal2 28280 563 28280 575 8 MemEn
rlabel metal2 28280 611 28280 623 8 OpcodeCondIn[6]
rlabel metal2 28280 899 28280 911 6 nWait
rlabel metal2 27961 0 28161 0 1 GND!
rlabel metal2 0 8181 0 8193 4 OpcodeCondIn[5]
rlabel metal2 0 8157 0 8169 4 Op2Sel[1]
rlabel metal2 0 8133 0 8145 4 OpcodeCondIn[7]
rlabel metal2 0 8109 0 8121 4 PcSel[0]
rlabel metal2 0 3988 0 4000 4 RwSel[1]
rlabel metal2 0 3964 0 3976 4 Rs1Sel[0]
rlabel metal2 0 3940 0 3952 4 ALE
rlabel metal2 0 3916 0 3928 4 Flags[3]
rlabel metal2 0 155 0 167 2 LrEn
rlabel metal2 0 131 0 143 2 Rs1Sel[1]
rlabel metal2 0 107 0 119 2 Flags[2]
rlabel metal2 0 83 0 95 2 nWE
rlabel metal2 145 0 345 0 1 Vdd!
rlabel metal2 27961 8252 28161 8252 5 GND!
rlabel metal2 145 8252 345 8252 5 Vdd!
rlabel metal2 361 0 373 0 1 SDI
rlabel metal2 385 0 397 0 1 Test
rlabel metal2 409 0 421 0 1 Clock
rlabel metal2 433 0 445 0 1 nReset
rlabel metal2 433 8252 445 8252 5 nReset
rlabel metal2 385 8252 397 8252 5 Test
rlabel metal2 409 8252 421 8252 5 Clock
rlabel metal2 361 8252 373 8252 5 SDO
<< end >>
