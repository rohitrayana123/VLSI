magic
tech c035u
timestamp 1394990067
<< metal1 >>
rect 32232 31758 32266 31762
rect 32221 31752 32266 31758
rect 32221 31748 32242 31752
rect 32256 31597 32266 31752
rect 32232 31566 32290 31570
rect 32221 31560 32290 31566
rect 32221 31556 32242 31560
rect 32256 30805 32266 31535
rect 32280 30802 32290 31560
rect 32280 30792 32314 30802
rect 32232 30774 32290 30778
rect 32221 30768 32290 30774
rect 32221 30764 32242 30768
rect 32256 30037 32266 30743
rect 32280 30037 32290 30768
rect 32304 30034 32314 30792
rect 32304 30024 32338 30034
rect 32232 30006 32314 30010
rect 32221 30000 32314 30006
rect 32221 29996 32242 30000
rect 32256 29293 32266 29975
rect 32280 29293 32290 29975
rect 32304 29293 32314 30000
rect 32328 29290 32338 30024
rect 32328 29280 32362 29290
rect 32232 29262 32338 29266
rect 32221 29256 32338 29262
rect 32221 29252 32242 29256
rect 32256 28333 32266 29231
rect 32280 28333 32290 29231
rect 32304 28333 32314 29231
rect 32328 28333 32338 29256
rect 32352 28330 32362 29280
rect 32352 28320 32386 28330
rect 32232 28302 32362 28306
rect 32221 28296 32362 28302
rect 32221 28292 32242 28296
rect 32256 27589 32266 28271
rect 32280 27589 32290 28271
rect 32304 27589 32314 28271
rect 32328 27589 32338 28271
rect 32352 27589 32362 28296
rect 32376 27586 32386 28320
rect 32376 27576 32410 27586
rect 32232 27558 32386 27562
rect 32221 27552 32386 27558
rect 32221 27548 32242 27552
rect 32256 27421 32266 27527
rect 32280 27421 32290 27527
rect 32304 27421 32314 27527
rect 32328 27421 32338 27527
rect 32352 27421 32362 27527
rect 32376 27421 32386 27552
rect 32400 27418 32410 27576
rect 32400 27408 32434 27418
rect 32232 27390 32410 27394
rect 32221 27384 32410 27390
rect 32221 27380 32242 27384
rect 32256 18013 32266 27359
rect 32280 18013 32290 27359
rect 32304 18013 32314 27359
rect 32328 18013 32338 27359
rect 32352 18013 32362 27359
rect 32376 18013 32386 27359
rect 32400 18013 32410 27384
rect 32424 18010 32434 27408
rect 66696 23386 66735 23390
rect 32688 23380 66735 23386
rect 32688 23376 66706 23380
rect 32424 18000 32458 18010
rect 32232 17982 32434 17986
rect 32221 17976 32434 17982
rect 32221 17972 32242 17976
rect 32256 17821 32266 17951
rect 32280 17821 32290 17951
rect 32304 17821 32314 17951
rect 32328 17821 32338 17951
rect 32352 17821 32362 17951
rect 32376 17821 32386 17951
rect 32400 17821 32410 17951
rect 32424 17821 32434 17976
rect 32448 17818 32458 18000
rect 32448 17808 32482 17818
rect 32232 17790 32458 17794
rect 32221 17784 32458 17790
rect 32221 17780 32242 17784
rect 32256 17581 32266 17759
rect 32280 17581 32290 17759
rect 32304 17581 32314 17759
rect 32328 17581 32338 17759
rect 32352 17581 32362 17759
rect 32376 17581 32386 17759
rect 32400 17581 32410 17759
rect 32424 17581 32434 17759
rect 32448 17578 32458 17784
rect 32472 17602 32482 17808
rect 32472 17592 32506 17602
rect 32448 17568 32482 17578
rect 32232 17550 32458 17554
rect 32221 17544 32458 17550
rect 32221 17540 32242 17544
rect 32256 17341 32266 17519
rect 32280 17341 32290 17519
rect 32304 17341 32314 17519
rect 32328 17341 32338 17519
rect 32352 17341 32362 17519
rect 32376 17341 32386 17519
rect 32400 17341 32410 17519
rect 32424 17341 32434 17519
rect 32448 17341 32458 17544
rect 32472 17338 32482 17568
rect 32496 17362 32506 17592
rect 32496 17352 32530 17362
rect 32472 17328 32506 17338
rect 32221 17304 32482 17314
rect 32256 16861 32266 17279
rect 32280 16861 32290 17279
rect 32304 16861 32314 17279
rect 32328 16861 32338 17279
rect 32352 16861 32362 17279
rect 32376 16861 32386 17279
rect 32400 16861 32410 17279
rect 32424 16861 32434 17279
rect 32448 16861 32458 17279
rect 32472 16861 32482 17304
rect 32496 16861 32506 17328
rect 32520 16858 32530 17352
rect 32520 16848 32554 16858
rect 32221 16824 32530 16834
rect 32256 16621 32266 16799
rect 32280 16621 32290 16799
rect 32304 16621 32314 16799
rect 32328 16621 32338 16799
rect 32352 16621 32362 16799
rect 32376 16621 32386 16799
rect 32400 16621 32410 16799
rect 32424 16621 32434 16799
rect 32448 16621 32458 16799
rect 32472 16621 32482 16799
rect 32496 16621 32506 16799
rect 32520 16621 32530 16824
rect 32544 16618 32554 16848
rect 32544 16608 32578 16618
rect 32221 16584 32554 16594
rect 32256 16381 32266 16559
rect 32280 16381 32290 16559
rect 32304 16381 32314 16559
rect 32328 16381 32338 16559
rect 32352 16381 32362 16559
rect 32376 16381 32386 16559
rect 32400 16381 32410 16559
rect 32424 16381 32434 16559
rect 32448 16381 32458 16559
rect 32472 16381 32482 16559
rect 32496 16378 32506 16559
rect 32520 16405 32530 16559
rect 32544 16405 32554 16584
rect 32568 16402 32578 16608
rect 32568 16392 32602 16402
rect 32496 16368 32578 16378
rect 32221 16344 32506 16354
rect 32256 16141 32266 16319
rect 32280 16141 32290 16319
rect 32304 16141 32314 16319
rect 32328 16141 32338 16319
rect 32352 16141 32362 16319
rect 32376 16138 32386 16319
rect 32400 16165 32410 16319
rect 32424 16165 32434 16319
rect 32448 16165 32458 16319
rect 32472 16165 32482 16319
rect 32496 16165 32506 16344
rect 32520 16165 32530 16343
rect 32544 16165 32554 16343
rect 32568 16165 32578 16368
rect 32592 16162 32602 16392
rect 32592 16152 32626 16162
rect 32376 16128 32602 16138
rect 32221 16104 32386 16114
rect 32256 9877 32266 16079
rect 32280 9877 32290 16079
rect 32304 9877 32314 16079
rect 32328 9877 32338 16079
rect 32352 9877 32362 16079
rect 32376 9877 32386 16104
rect 32400 9877 32410 16103
rect 32424 9877 32434 16103
rect 32448 9877 32458 16103
rect 32472 9877 32482 16103
rect 32496 9877 32506 16103
rect 32520 9874 32530 16103
rect 32544 9901 32554 16103
rect 32568 9901 32578 16103
rect 32592 9901 32602 16128
rect 32616 9898 32626 16152
rect 32616 9888 32650 9898
rect 32520 9864 32626 9874
rect 32232 9846 32530 9850
rect 32221 9840 32530 9846
rect 32221 9836 32242 9840
rect 32256 9133 32266 9815
rect 32280 9133 32290 9815
rect 32304 9133 32314 9815
rect 32328 9133 32338 9815
rect 32352 9133 32362 9815
rect 32376 9133 32386 9815
rect 32400 9133 32410 9815
rect 32424 9130 32434 9815
rect 32448 9157 32458 9815
rect 32472 9157 32482 9815
rect 32496 9157 32506 9815
rect 32520 9157 32530 9840
rect 32544 9157 32554 9839
rect 32568 9154 32578 9839
rect 32592 9178 32602 9839
rect 32616 9205 32626 9864
rect 32640 9202 32650 9888
rect 32640 9192 32674 9202
rect 32592 9168 32650 9178
rect 32568 9144 32602 9154
rect 32424 9120 32578 9130
rect 32232 9102 32434 9106
rect 32221 9096 32434 9102
rect 32221 9092 32242 9096
rect 32256 8701 32266 9071
rect 32280 8701 32290 9071
rect 32304 8701 32314 9071
rect 32328 8701 32338 9071
rect 32352 8701 32362 9071
rect 32376 8701 32386 9071
rect 32400 8701 32410 9071
rect 32424 8701 32434 9096
rect 32448 8701 32458 9095
rect 32472 8701 32482 9095
rect 32496 8701 32506 9095
rect 32520 8701 32530 9095
rect 32544 8701 32554 9095
rect 32568 8701 32578 9120
rect 32592 8701 32602 9144
rect 32616 8701 32626 9143
rect 32640 8698 32650 9168
rect 32664 8722 32674 9192
rect 32688 8749 32698 23376
rect 66696 17434 66735 17442
rect 32856 17432 66735 17434
rect 32856 17424 66706 17432
rect 32856 17221 32866 17424
rect 66696 17194 66735 17202
rect 32712 17192 66735 17194
rect 32712 17184 66706 17192
rect 32712 8749 32722 17184
rect 32856 15541 32866 17159
rect 66696 16954 66735 16962
rect 32904 16952 66735 16954
rect 32904 16944 66706 16952
rect 32904 15541 32914 16944
rect 66696 16714 66735 16722
rect 32928 16712 66735 16714
rect 32928 16704 66706 16712
rect 32928 15541 32938 16704
rect 66696 16474 66735 16482
rect 32952 16472 66735 16474
rect 32952 16464 66706 16472
rect 32952 15541 32962 16464
rect 66696 16234 66735 16242
rect 32976 16232 66735 16234
rect 32976 16224 66706 16232
rect 32976 15541 32986 16224
rect 66696 15994 66735 16002
rect 33000 15992 66735 15994
rect 33000 15984 66706 15992
rect 33000 15541 33010 15984
rect 66696 15754 66735 15762
rect 33024 15752 66735 15754
rect 33024 15744 66706 15752
rect 33024 15541 33034 15744
rect 66696 15514 66735 15522
rect 32760 15512 66735 15514
rect 32760 15504 66706 15512
rect 32760 14341 32770 15504
rect 32856 14341 32866 15479
rect 32904 14341 32914 15479
rect 32928 14341 32938 15479
rect 32952 14341 32962 15479
rect 32976 14341 32986 15479
rect 33000 14341 33010 15479
rect 33024 14341 33034 15479
rect 66696 15274 66735 15282
rect 33048 15272 66735 15274
rect 33048 15264 66706 15272
rect 33048 14341 33058 15264
rect 66696 15034 66735 15042
rect 33072 15032 66735 15034
rect 33072 15024 66706 15032
rect 33072 14341 33082 15024
rect 66696 14794 66735 14802
rect 33096 14792 66735 14794
rect 33096 14784 66706 14792
rect 33096 14341 33106 14784
rect 66696 14554 66735 14562
rect 33120 14552 66735 14554
rect 33120 14544 66706 14552
rect 33120 14341 33130 14544
rect 66696 14314 66735 14322
rect 32736 14312 66735 14314
rect 32736 14304 66706 14312
rect 32736 8749 32746 14304
rect 32760 8749 32770 14279
rect 32856 14101 32866 14279
rect 32904 14101 32914 14279
rect 32928 14101 32938 14279
rect 32952 14101 32962 14279
rect 32976 14101 32986 14279
rect 33000 14101 33010 14279
rect 33024 14101 33034 14279
rect 33048 14101 33058 14279
rect 33072 14101 33082 14279
rect 33096 14101 33106 14279
rect 33120 14101 33130 14279
rect 66696 14074 66735 14082
rect 32808 14072 66735 14074
rect 32808 14064 66706 14072
rect 32808 12181 32818 14064
rect 32856 13621 32866 14039
rect 32904 13621 32914 14039
rect 32928 13621 32938 14039
rect 32952 13621 32962 14039
rect 32976 13621 32986 14039
rect 33000 13621 33010 14039
rect 33024 13621 33034 14039
rect 33048 13621 33058 14039
rect 33072 13621 33082 14039
rect 33096 13621 33106 14039
rect 33120 13621 33130 14039
rect 66696 13834 66735 13842
rect 33144 13832 66735 13834
rect 33144 13824 66706 13832
rect 33144 13621 33154 13824
rect 66696 13594 66735 13602
rect 32832 13592 66735 13594
rect 32832 13584 66706 13592
rect 32832 12181 32842 13584
rect 32856 12181 32866 13559
rect 32904 12181 32914 13559
rect 32928 12181 32938 13559
rect 32952 12181 32962 13559
rect 32976 12181 32986 13559
rect 33000 12181 33010 13559
rect 33024 12181 33034 13559
rect 33048 12181 33058 13559
rect 33072 12181 33082 13559
rect 33096 12181 33106 13559
rect 33120 12181 33130 13559
rect 33144 12181 33154 13559
rect 66696 13354 66735 13362
rect 33168 13352 66735 13354
rect 33168 13344 66706 13352
rect 33168 12181 33178 13344
rect 66696 13114 66735 13122
rect 41160 13112 66735 13114
rect 41160 13104 66706 13112
rect 41160 12901 41170 13104
rect 66696 12874 66735 12882
rect 33192 12872 66735 12874
rect 33192 12864 66706 12872
rect 33192 12181 33202 12864
rect 41160 12661 41170 12839
rect 66696 12634 66735 12642
rect 33240 12632 66735 12634
rect 33240 12624 66706 12632
rect 33240 12181 33250 12624
rect 41160 12421 41170 12599
rect 66696 12394 66735 12402
rect 33264 12392 66735 12394
rect 33264 12384 66706 12392
rect 33264 12181 33274 12384
rect 41160 12181 41170 12359
rect 66696 12154 66735 12162
rect 32784 12152 66735 12154
rect 32784 12144 66706 12152
rect 32784 8749 32794 12144
rect 32808 8749 32818 12119
rect 32832 8749 32842 12119
rect 32856 8749 32866 12119
rect 32664 8712 32890 8722
rect 32640 8688 32674 8698
rect 32221 8664 32650 8674
rect 32640 8626 32650 8664
rect 32664 8629 32674 8688
rect 32688 8629 32698 8687
rect 32712 8629 32722 8687
rect 32736 8629 32746 8687
rect 32760 8629 32770 8687
rect 32784 8629 32794 8687
rect 32808 8629 32818 8687
rect 32832 8629 32842 8687
rect 32856 8629 32866 8687
rect 32880 8629 32890 8712
rect 32904 8629 32914 12119
rect 32928 8629 32938 12119
rect 32952 8629 32962 12119
rect 32976 8629 32986 12119
rect 33000 8629 33010 12119
rect 33024 8629 33034 12119
rect 33048 8629 33058 12119
rect 33072 8629 33082 12119
rect 33096 8629 33106 12119
rect 33120 8629 33130 12119
rect 33144 8629 33154 12119
rect 32173 8616 32650 8626
rect 33168 8602 33178 12119
rect 32149 8592 33178 8602
rect 32125 8568 32351 8578
rect 32640 8568 32663 8578
rect 32616 8554 32626 8567
rect 32101 8544 32626 8554
rect 32077 8520 32591 8530
rect 32640 8530 32650 8568
rect 33192 8578 33202 12119
rect 33240 8821 33250 12119
rect 33264 8821 33274 12119
rect 41160 11941 41170 12119
rect 66696 11914 66735 11922
rect 33288 11912 66735 11914
rect 33288 11904 66706 11912
rect 33288 8821 33298 11904
rect 41160 11701 41170 11879
rect 66696 11674 66735 11682
rect 33312 11672 66735 11674
rect 33312 11664 66706 11672
rect 33312 8821 33322 11664
rect 41160 8821 41170 11639
rect 66696 8794 66735 8802
rect 33216 8792 66735 8794
rect 33216 8784 66706 8792
rect 33216 8581 33226 8784
rect 33168 8568 33202 8578
rect 32688 8554 32698 8567
rect 32664 8544 32698 8554
rect 32664 8533 32674 8544
rect 32629 8520 32650 8530
rect 33072 8530 33082 8567
rect 32701 8520 33082 8530
rect 32053 8496 32927 8506
rect 33096 8506 33106 8567
rect 33120 8509 33130 8567
rect 33144 8509 33154 8567
rect 33168 8509 33178 8568
rect 33240 8554 33250 8759
rect 33192 8544 33250 8554
rect 33192 8509 33202 8544
rect 33264 8530 33274 8759
rect 33240 8520 33274 8530
rect 33240 8509 33250 8520
rect 33085 8496 33106 8506
rect 33288 8506 33298 8759
rect 33264 8496 33298 8506
rect 33264 8482 33274 8496
rect 33312 8482 33322 8759
rect 32029 8472 33274 8482
rect 33288 8472 33322 8482
rect 32005 8448 33239 8458
rect 33288 8458 33298 8472
rect 33264 8448 33298 8458
rect 31981 8424 33023 8434
rect 33096 8424 33119 8434
rect 33096 8410 33106 8424
rect 33264 8434 33274 8448
rect 33240 8424 33274 8434
rect 33144 8410 33154 8423
rect 31957 8400 33106 8410
rect 33120 8400 33154 8410
rect 31933 8376 32567 8386
rect 32605 8376 32615 8386
rect 32653 8376 32663 8386
rect 32941 8376 32951 8386
rect 33037 8376 33047 8386
rect 33120 8386 33130 8400
rect 33168 8386 33178 8423
rect 33096 8376 33130 8386
rect 33144 8376 33178 8386
rect 33072 8362 33082 8375
rect 31909 8352 33082 8362
rect 33096 8338 33106 8376
rect 33144 8362 33154 8376
rect 33192 8362 33202 8423
rect 33216 8365 33226 8423
rect 31885 8328 33106 8338
rect 33120 8352 33154 8362
rect 33168 8352 33202 8362
rect 31861 8304 32543 8314
rect 32581 8304 32591 8314
rect 32629 8304 32903 8314
rect 32952 8304 32975 8314
rect 32928 8290 32938 8303
rect 32952 8293 32962 8304
rect 33120 8314 33130 8352
rect 33168 8338 33178 8352
rect 33240 8338 33250 8424
rect 33048 8304 33130 8314
rect 33144 8328 33178 8338
rect 33192 8328 33250 8338
rect 31824 8280 32938 8290
rect 31824 8269 31834 8280
rect 33000 8290 33010 8303
rect 32976 8280 33010 8290
rect 32352 8256 32519 8266
rect 32328 8242 32338 8255
rect 32352 8245 32362 8256
rect 32544 8256 32567 8266
rect 31800 8232 32338 8242
rect 31800 8221 31810 8232
rect 32544 8242 32554 8256
rect 32592 8256 32639 8266
rect 32520 8232 32554 8242
rect 32496 8218 32506 8231
rect 32520 8221 32530 8232
rect 32592 8242 32602 8256
rect 32976 8266 32986 8280
rect 33024 8266 33034 8303
rect 32677 8256 32986 8266
rect 33000 8256 33034 8266
rect 32581 8232 32602 8242
rect 33000 8242 33010 8256
rect 33048 8242 33058 8304
rect 33144 8290 33154 8328
rect 33192 8314 33202 8328
rect 32653 8232 33010 8242
rect 33024 8232 33058 8242
rect 33072 8280 33154 8290
rect 33168 8304 33202 8314
rect 32341 8208 32506 8218
rect 32557 8208 32855 8218
rect 32917 8208 32951 8218
rect 33024 8218 33034 8232
rect 33072 8218 33082 8280
rect 33168 8266 33178 8304
rect 32976 8208 33034 8218
rect 33048 8208 33082 8218
rect 33096 8256 33178 8266
rect 32976 8194 32986 8208
rect 33048 8194 33058 8208
rect 33096 8194 33106 8256
rect 31776 8184 32986 8194
rect 33000 8184 33058 8194
rect 33072 8184 33106 8194
rect 31776 6421 31786 8184
rect 32592 8160 32903 8170
rect 31800 6421 31810 8159
rect 31824 6421 31834 8159
rect 31848 6421 31858 8159
rect 31872 6421 31882 8159
rect 31896 6421 31906 8159
rect 31920 6421 31930 8159
rect 31944 6421 31954 8159
rect 31968 6421 31978 8159
rect 31992 6421 32002 8159
rect 32016 6421 32026 8159
rect 32040 6421 32050 8159
rect 32064 6421 32074 8159
rect 32088 6421 32098 8159
rect 32112 6421 32122 8159
rect 32136 6421 32146 8159
rect 32160 6421 32170 8159
rect 32256 6421 32266 8159
rect 32280 6421 32290 8159
rect 32304 6421 32314 8159
rect 32328 6421 32338 8159
rect 32352 6421 32362 8159
rect 32376 6421 32386 8159
rect 32400 6421 32410 8159
rect 32424 6421 32434 8159
rect 32448 6421 32458 8159
rect 32472 6421 32482 8159
rect 32520 6421 32530 8159
rect 32544 6421 32554 8159
rect 32568 6421 32578 8159
rect 32592 6421 32602 8160
rect 33000 8170 33010 8184
rect 33072 8170 33082 8184
rect 32928 8160 33010 8170
rect 33024 8160 33082 8170
rect 32928 8146 32938 8160
rect 33024 8146 33034 8160
rect 32856 8136 32938 8146
rect 32952 8136 33034 8146
rect 32616 6421 32626 8135
rect 32640 6421 32650 8135
rect 32664 6421 32674 8135
rect 32688 6421 32698 8135
rect 32712 6421 32722 8135
rect 32736 6421 32746 8135
rect 32760 6421 32770 8135
rect 32784 6421 32794 8135
rect 32808 6421 32818 8135
rect 32832 6421 32842 8135
rect 32856 6421 32866 8136
rect 32952 8122 32962 8136
rect 32904 8112 32962 8122
rect 32880 6421 32890 8111
rect 32904 6421 32914 8112
rect 33216 6421 33226 8303
rect 41160 6421 41170 8759
rect 66696 6394 66735 6402
rect 31752 6392 66735 6394
rect 31752 6384 66706 6392
rect 31752 6181 31762 6384
rect 31776 6181 31786 6359
rect 31800 6181 31810 6359
rect 31824 6181 31834 6359
rect 31848 6181 31858 6359
rect 31872 6181 31882 6359
rect 31896 6181 31906 6359
rect 31920 6181 31930 6359
rect 31944 6181 31954 6359
rect 31968 6181 31978 6359
rect 31992 6181 32002 6359
rect 32016 6181 32026 6359
rect 32040 6181 32050 6359
rect 32064 6181 32074 6359
rect 32088 6181 32098 6359
rect 32112 6181 32122 6359
rect 32136 6181 32146 6359
rect 32160 6181 32170 6359
rect 32256 6181 32266 6359
rect 32280 6181 32290 6359
rect 32304 6181 32314 6359
rect 32328 6181 32338 6359
rect 32352 6181 32362 6359
rect 32376 6181 32386 6359
rect 32400 6181 32410 6359
rect 32424 6181 32434 6359
rect 32448 6181 32458 6359
rect 32472 6181 32482 6359
rect 32520 6181 32530 6359
rect 32544 6181 32554 6359
rect 32568 6181 32578 6359
rect 32592 6181 32602 6359
rect 32616 6181 32626 6359
rect 32640 6181 32650 6359
rect 32664 6181 32674 6359
rect 32688 6181 32698 6359
rect 32712 6181 32722 6359
rect 32736 6181 32746 6359
rect 32760 6181 32770 6359
rect 32784 6181 32794 6359
rect 32808 6181 32818 6359
rect 32832 6181 32842 6359
rect 32856 6181 32866 6359
rect 32880 6181 32890 6359
rect 32904 6181 32914 6359
rect 33216 6181 33226 6359
rect 41160 6181 41170 6359
rect 66696 6154 66735 6162
rect 31728 6152 66735 6154
rect 31728 6144 66706 6152
rect 31728 5461 31738 6144
rect 31752 5461 31762 6119
rect 31776 5461 31786 6119
rect 31800 5461 31810 6119
rect 31824 5461 31834 6119
rect 31848 5461 31858 6119
rect 31872 5461 31882 6119
rect 31896 5461 31906 6119
rect 31920 5461 31930 6119
rect 31944 5461 31954 6119
rect 31968 5461 31978 6119
rect 31992 5461 32002 6119
rect 32016 5461 32026 6119
rect 32040 5461 32050 6119
rect 32064 5461 32074 6119
rect 32088 5461 32098 6119
rect 32112 5461 32122 6119
rect 32136 5461 32146 6119
rect 32160 5461 32170 6119
rect 32256 5461 32266 6119
rect 32280 5461 32290 6119
rect 32304 5461 32314 6119
rect 32328 5461 32338 6119
rect 32352 5461 32362 6119
rect 32376 5461 32386 6119
rect 32400 5461 32410 6119
rect 32424 5461 32434 6119
rect 32448 5461 32458 6119
rect 32472 5461 32482 6119
rect 32520 5461 32530 6119
rect 32544 5461 32554 6119
rect 32568 5461 32578 6119
rect 32592 5461 32602 6119
rect 32616 5461 32626 6119
rect 32640 5461 32650 6119
rect 32664 5461 32674 6119
rect 32688 5461 32698 6119
rect 32712 5461 32722 6119
rect 32736 5461 32746 6119
rect 32760 5461 32770 6119
rect 32784 5461 32794 6119
rect 32808 5461 32818 6119
rect 32832 5461 32842 6119
rect 32856 5461 32866 6119
rect 32880 5461 32890 6119
rect 32904 5461 32914 6119
rect 33216 5461 33226 6119
rect 41160 5941 41170 6119
rect 66696 5914 66735 5922
rect 33336 5912 66735 5914
rect 33336 5904 66706 5912
rect 33336 5461 33346 5904
rect 41160 5701 41170 5879
rect 66696 5674 66735 5682
rect 33384 5672 66735 5674
rect 33384 5664 66706 5672
rect 33384 5461 33394 5664
rect 41160 5461 41170 5639
rect 66696 5434 66735 5442
rect 31704 5432 66735 5434
rect 31704 5424 66706 5432
rect 27613 5400 27647 5410
rect 27877 5400 27935 5410
rect 27973 5400 28031 5410
rect 28093 5400 28127 5410
rect 27565 5376 27743 5386
rect 27805 5376 28247 5386
rect 27541 5352 28343 5362
rect 28405 5352 28439 5362
rect 26989 5328 27071 5338
rect 27253 5328 27287 5338
rect 27325 5328 27407 5338
rect 27469 5328 28535 5338
rect 28597 5328 28631 5338
rect 28693 5328 28727 5338
rect 28765 5328 28823 5338
rect 30469 5328 30527 5338
rect 26869 5304 27191 5314
rect 27229 5304 28919 5314
rect 30253 5304 30287 5314
rect 30325 5304 30383 5314
rect 30445 5304 30647 5314
rect 30685 5304 30767 5314
rect 24565 5280 24599 5290
rect 26461 5280 26495 5290
rect 26797 5280 29015 5290
rect 30013 5280 30071 5290
rect 30109 5280 30167 5290
rect 30229 5280 30887 5290
rect 30949 5280 31007 5290
rect 31453 5280 31487 5290
rect 31525 5280 31583 5290
rect 24541 5256 24695 5266
rect 26413 5256 26591 5266
rect 26653 5256 26711 5266
rect 26749 5256 29111 5266
rect 29989 5256 31127 5266
rect 31165 5256 31247 5266
rect 31704 5266 31714 5424
rect 31405 5256 31714 5266
rect 31728 5245 31738 5399
rect 31752 5245 31762 5399
rect 24517 5232 24815 5242
rect 24853 5232 24935 5242
rect 24973 5232 25031 5242
rect 26389 5232 29231 5242
rect 29269 5232 29327 5242
rect 29437 5232 31703 5242
rect 24397 5208 24455 5218
rect 24493 5208 25127 5218
rect 25189 5208 25223 5218
rect 25261 5208 25343 5218
rect 25381 5208 25439 5218
rect 25477 5208 25535 5218
rect 25645 5208 26255 5218
rect 31776 5218 31786 5399
rect 26317 5208 31786 5218
rect 24277 5184 24335 5194
rect 31800 5194 31810 5399
rect 31824 5197 31834 5399
rect 24373 5184 31810 5194
rect 31848 5170 31858 5399
rect 24253 5160 31858 5170
rect 24037 5136 24095 5146
rect 31872 5146 31882 5399
rect 24133 5136 31882 5146
rect 23917 5112 23975 5122
rect 31896 5122 31906 5399
rect 24013 5112 31906 5122
rect 31920 5101 31930 5399
rect 31944 5101 31954 5399
rect 31968 5101 31978 5399
rect 23701 5088 23735 5098
rect 23821 5088 23855 5098
rect 23893 5088 31895 5098
rect 23557 5064 23615 5074
rect 31992 5074 32002 5399
rect 23653 5064 32002 5074
rect 32016 5050 32026 5399
rect 23533 5040 32026 5050
rect 23413 5016 29423 5026
rect 29461 5016 32015 5026
rect 32040 5002 32050 5399
rect 32064 5005 32074 5399
rect 23317 4992 32050 5002
rect 32088 4978 32098 5399
rect 32112 4981 32122 5399
rect 32136 4981 32146 5399
rect 32160 4981 32170 5399
rect 32256 4981 32266 5399
rect 32280 4981 32290 5399
rect 32304 4981 32314 5399
rect 32328 4981 32338 5399
rect 32352 4981 32362 5399
rect 32376 4981 32386 5399
rect 32400 4981 32410 5399
rect 32424 4981 32434 5399
rect 32448 4981 32458 5399
rect 32472 4981 32482 5399
rect 23293 4968 32098 4978
rect 23269 4944 28391 4954
rect 28429 4944 32506 4954
rect 23173 4920 32111 4930
rect 23149 4896 27791 4906
rect 27829 4896 32194 4906
rect 23029 4872 23087 4882
rect 23125 4872 32111 4882
rect 32184 4882 32194 4896
rect 32256 4885 32266 4919
rect 32280 4885 32290 4919
rect 32304 4885 32314 4919
rect 32328 4885 32338 4919
rect 32352 4885 32362 4919
rect 32376 4885 32386 4919
rect 32400 4885 32410 4919
rect 32424 4885 32434 4919
rect 32448 4885 32458 4919
rect 32472 4885 32482 4919
rect 32496 4885 32506 4944
rect 32520 4885 32530 5399
rect 32544 4885 32554 5399
rect 32568 4885 32578 5399
rect 32592 4885 32602 5399
rect 32616 4885 32626 5399
rect 32640 4885 32650 5399
rect 32664 4885 32674 5399
rect 32688 4885 32698 5399
rect 32712 4885 32722 5399
rect 32736 4885 32746 5399
rect 32760 4885 32770 5399
rect 32784 4885 32794 5399
rect 32808 4885 32818 5399
rect 32832 4885 32842 5399
rect 32856 4885 32866 5399
rect 32184 4872 32218 4882
rect 22813 4848 22895 4858
rect 22957 4848 24959 4858
rect 24997 4848 25295 4858
rect 25309 4848 26567 4858
rect 26581 4848 27119 4858
rect 27133 4848 30935 4858
rect 30973 4848 31223 4858
rect 31237 4848 31679 4858
rect 32208 4858 32218 4872
rect 32880 4882 32890 5399
rect 32904 4909 32914 5399
rect 32880 4872 32927 4882
rect 31693 4848 32194 4858
rect 32208 4848 32951 4858
rect 22789 4824 32159 4834
rect 32197 4824 32231 4834
rect 32509 4824 32975 4834
rect 22429 4800 22535 4810
rect 22573 4800 22631 4810
rect 22693 4800 29255 4810
rect 29293 4800 33010 4810
rect 33000 4789 33010 4800
rect 22357 4776 32879 4786
rect 22261 4752 22295 4762
rect 22333 4752 22991 4762
rect 23053 4752 26735 4762
rect 26773 4752 33023 4762
rect 33216 4741 33226 5399
rect 33336 4741 33346 5399
rect 33384 4741 33394 5399
rect 41160 4741 41170 5399
rect 66696 5194 66735 5202
rect 59760 5192 66735 5194
rect 59760 5184 66706 5192
rect 59760 4981 59770 5184
rect 66696 4954 66735 4962
rect 59040 4952 66735 4954
rect 59040 4944 66706 4952
rect 59040 4741 59050 4944
rect 59760 4741 59770 4919
rect 22213 4728 23783 4738
rect 23797 4728 32207 4738
rect 32244 4728 33047 4738
rect 21637 4704 21671 4714
rect 21733 4704 21791 4714
rect 21853 4704 21911 4714
rect 21949 4704 22031 4714
rect 22069 4704 22127 4714
rect 22189 4704 32495 4714
rect 66696 4714 66735 4722
rect 32893 4712 66735 4714
rect 32893 4704 66706 4712
rect 21589 4680 32063 4690
rect 32101 4680 32172 4690
rect 32221 4680 32879 4690
rect 21085 4656 21143 4666
rect 21565 4656 32207 4666
rect 32244 4656 33071 4666
rect 20461 4632 20543 4642
rect 20581 4632 20639 4642
rect 20725 4632 20759 4642
rect 20821 4632 20855 4642
rect 20989 4632 21239 4642
rect 21277 4632 21335 4642
rect 21493 4632 32375 4642
rect 32509 4632 33095 4642
rect 20437 4608 21431 4618
rect 21469 4608 23159 4618
rect 23197 4608 31151 4618
rect 31189 4608 32172 4618
rect 32221 4608 33119 4618
rect 20365 4584 33143 4594
rect 20341 4560 27503 4570
rect 27589 4560 32207 4570
rect 32244 4560 33178 4570
rect 20221 4536 32351 4546
rect 32389 4536 32543 4546
rect 33168 4525 33178 4560
rect 19405 4512 19463 4522
rect 19501 4512 19559 4522
rect 19621 4512 19703 4522
rect 19813 4512 26951 4522
rect 27013 4512 27719 4522
rect 27733 4512 32172 4522
rect 32221 4512 32543 4522
rect 19285 4488 19343 4498
rect 19381 4488 33202 4498
rect 33192 4477 33202 4488
rect 19165 4464 19223 4474
rect 19261 4464 32759 4474
rect 33216 4450 33226 4679
rect 19093 4440 33226 4450
rect 19069 4416 32375 4426
rect 32509 4416 32807 4426
rect 32965 4416 33215 4426
rect 18949 4392 20423 4402
rect 20485 4392 31175 4402
rect 31213 4392 31655 4402
rect 31669 4392 32207 4402
rect 32244 4392 32951 4402
rect 33037 4392 33239 4402
rect 18781 4368 18815 4378
rect 18877 4368 24023 4378
rect 24061 4368 33263 4378
rect 18637 4344 18719 4354
rect 18757 4344 32183 4354
rect 32221 4344 33287 4354
rect 18565 4320 33322 4330
rect 33312 4309 33322 4320
rect 33336 4309 33346 4679
rect 18469 4296 18503 4306
rect 18541 4296 33023 4306
rect 33384 4285 33394 4679
rect 41160 4501 41170 4679
rect 59040 4501 59050 4679
rect 59760 4501 59770 4679
rect 66696 4474 66735 4482
rect 33480 4472 66735 4474
rect 33480 4464 66706 4472
rect 18445 4272 32495 4282
rect 32557 4272 33359 4282
rect 33480 4261 33490 4464
rect 41160 4261 41170 4439
rect 59040 4261 59050 4439
rect 59760 4261 59770 4439
rect 18349 4248 18383 4258
rect 18421 4248 32207 4258
rect 32245 4248 33407 4258
rect 66696 4234 66735 4242
rect 18301 4232 66735 4234
rect 18301 4224 66706 4232
rect 18277 4200 27599 4210
rect 27637 4200 32194 4210
rect 32221 4200 33431 4210
rect 33469 4200 33503 4210
rect 17365 4176 17447 4186
rect 17581 4176 33527 4186
rect 33565 4176 33599 4186
rect 35413 4176 35447 4186
rect 17149 4152 33695 4162
rect 35389 4152 35567 4162
rect 16933 4128 17087 4138
rect 17101 4128 17303 4138
rect 17317 4128 17519 4138
rect 17533 4128 17735 4138
rect 17749 4128 17951 4138
rect 17965 4128 18167 4138
rect 18181 4128 22055 4138
rect 22093 4128 23903 4138
rect 23941 4128 24047 4138
rect 24085 4128 27383 4138
rect 27397 4128 32207 4138
rect 32232 4128 33815 4138
rect 35269 4128 35327 4138
rect 35365 4128 35663 4138
rect 16717 4104 32172 4114
rect 32184 4104 32231 4114
rect 32184 4093 32194 4104
rect 32245 4104 33935 4114
rect 33973 4104 34031 4114
rect 34069 4104 34127 4114
rect 34165 4104 34223 4114
rect 35149 4104 35207 4114
rect 35245 4104 35759 4114
rect 16501 4080 22751 4090
rect 22837 4080 32172 4090
rect 32221 4080 34343 4090
rect 34861 4080 34895 4090
rect 34933 4080 34991 4090
rect 35029 4080 35087 4090
rect 35125 4080 35855 4090
rect 16285 4056 33479 4066
rect 33541 4056 34439 4066
rect 34477 4056 34535 4066
rect 34741 4056 34799 4066
rect 34837 4056 35951 4066
rect 35989 4056 36047 4066
rect 16069 4032 21575 4042
rect 21613 4032 32543 4042
rect 32773 4032 32831 4042
rect 33277 4032 34199 4042
rect 34237 4032 34631 4042
rect 34693 4032 34943 4042
rect 34957 4032 36143 4042
rect 41160 4021 41170 4199
rect 59040 4021 59050 4199
rect 59760 4021 59770 4199
rect 15853 4008 32135 4018
rect 32173 4008 34775 4018
rect 34813 4008 36263 4018
rect 36301 4008 36359 4018
rect 15397 3984 15455 3994
rect 15637 3984 23231 3994
rect 23341 3984 32495 3994
rect 66696 3994 66735 4002
rect 33277 3992 66735 3994
rect 33277 3984 66706 3992
rect 15373 3960 32327 3970
rect 32365 3960 36455 3970
rect 15085 3936 15119 3946
rect 15325 3936 32663 3946
rect 32821 3936 32855 3946
rect 33253 3936 36551 3946
rect 15037 3912 32303 3922
rect 32341 3912 32855 3922
rect 33216 3922 33226 3935
rect 33216 3912 36671 3922
rect 14677 3888 14711 3898
rect 14749 3888 14807 3898
rect 14845 3888 14903 3898
rect 14941 3888 32207 3898
rect 32244 3888 36791 3898
rect 14581 3864 14615 3874
rect 14653 3864 19607 3874
rect 19645 3864 36887 3874
rect 36925 3864 37031 3874
rect 37069 3864 37127 3874
rect 37165 3864 37223 3874
rect 14485 3840 14519 3850
rect 14557 3840 17807 3850
rect 17821 3840 23303 3850
rect 23365 3840 37343 3850
rect 37405 3840 37463 3850
rect 37501 3840 37583 3850
rect 14269 3816 14327 3826
rect 14389 3816 14423 3826
rect 14461 3816 14831 3826
rect 14869 3816 21839 3826
rect 21877 3816 37679 3826
rect 37741 3816 37775 3826
rect 14245 3792 32759 3802
rect 32845 3792 32903 3802
rect 33205 3792 37871 3802
rect 14173 3768 19031 3778
rect 19117 3768 23255 3778
rect 23317 3768 32172 3778
rect 32221 3768 32903 3778
rect 33168 3778 33178 3791
rect 33168 3768 35807 3778
rect 35821 3768 37511 3778
rect 37525 3768 37967 3778
rect 14029 3744 18455 3754
rect 18493 3744 28679 3754
rect 28717 3744 38087 3754
rect 38125 3744 38183 3754
rect 13597 3720 13655 3730
rect 13693 3720 13751 3730
rect 13885 3720 14159 3730
rect 14197 3720 32687 3730
rect 32773 3720 32807 3730
rect 33133 3720 38303 3730
rect 13501 3696 13535 3706
rect 13573 3696 30455 3706
rect 30493 3696 32207 3706
rect 32244 3696 35183 3706
rect 35221 3696 38423 3706
rect 13477 3672 38519 3682
rect 13453 3648 19391 3658
rect 19429 3648 26639 3658
rect 26677 3648 32172 3658
rect 32221 3648 38663 3658
rect 13405 3624 25175 3634
rect 25213 3624 25511 3634
rect 25525 3624 26231 3634
rect 26245 3624 31367 3634
rect 31429 3624 38759 3634
rect 38917 3624 38951 3634
rect 39709 3624 39767 3634
rect 39805 3624 39863 3634
rect 39901 3624 39959 3634
rect 40501 3624 40559 3634
rect 40597 3624 40655 3634
rect 41160 3613 41170 3959
rect 13381 3600 20327 3610
rect 20389 3600 25631 3610
rect 25669 3600 31439 3610
rect 31477 3600 38855 3610
rect 38893 3600 39047 3610
rect 39229 3600 39263 3610
rect 39301 3600 39359 3610
rect 39517 3600 39551 3610
rect 39613 3600 39647 3610
rect 39685 3600 40055 3610
rect 40405 3600 40439 3610
rect 40477 3600 40775 3610
rect 40813 3600 40871 3610
rect 41053 3600 41087 3610
rect 41245 3600 41303 3610
rect 41341 3600 41399 3610
rect 13021 3576 13103 3586
rect 13141 3576 13199 3586
rect 13285 3576 15839 3586
rect 15877 3576 18431 3586
rect 18469 3576 26831 3586
rect 26893 3576 30671 3586
rect 30709 3576 34967 3586
rect 35005 3576 39167 3586
rect 39205 3576 39455 3586
rect 39493 3576 40151 3586
rect 40189 3576 40247 3586
rect 40285 3576 40343 3586
rect 40381 3576 40991 3586
rect 41029 3576 41495 3586
rect 41869 3576 41903 3586
rect 12997 3552 30431 3562
rect 30469 3552 32207 3562
rect 32244 3552 32687 3562
rect 32821 3552 32831 3562
rect 33109 3552 41615 3562
rect 41677 3552 41711 3562
rect 41749 3552 41807 3562
rect 41845 3552 41999 3562
rect 42037 3552 42119 3562
rect 12829 3528 12863 3538
rect 12949 3528 13583 3538
rect 13621 3528 32831 3538
rect 33072 3538 33082 3551
rect 59040 3541 59050 3959
rect 59760 3781 59770 3959
rect 66696 3754 66735 3762
rect 59640 3752 66735 3754
rect 59640 3744 66706 3752
rect 59640 3541 59650 3744
rect 59760 3541 59770 3719
rect 33072 3528 40415 3538
rect 40453 3528 42215 3538
rect 12709 3504 12767 3514
rect 12805 3504 26975 3514
rect 27037 3504 27695 3514
rect 27709 3504 34511 3514
rect 34549 3504 35471 3514
rect 35485 3504 39431 3514
rect 39469 3504 42335 3514
rect 66696 3514 66735 3522
rect 58920 3512 66735 3514
rect 58920 3504 66706 3512
rect 12637 3480 19079 3490
rect 19141 3480 33383 3490
rect 33445 3480 42455 3490
rect 12589 3456 13487 3466
rect 13525 3456 25415 3466
rect 25429 3456 30743 3466
rect 30757 3456 34079 3466
rect 34093 3456 39095 3466
rect 39109 3456 40895 3466
rect 40909 3456 42599 3466
rect 12373 3432 12431 3442
rect 12565 3432 20567 3442
rect 20605 3432 22799 3442
rect 22861 3432 31799 3442
rect 31861 3432 32172 3442
rect 32221 3432 35543 3442
rect 35581 3432 42695 3442
rect 12277 3408 12311 3418
rect 12349 3408 32759 3418
rect 33085 3408 35423 3418
rect 35461 3408 42815 3418
rect 12181 3384 12215 3394
rect 12253 3384 13127 3394
rect 13165 3384 32218 3394
rect 32244 3384 37103 3394
rect 12109 3360 24647 3370
rect 24661 3360 27839 3370
rect 32208 3370 32218 3384
rect 37141 3384 42935 3394
rect 27901 3360 32172 3370
rect 32208 3360 33575 3370
rect 33613 3360 43055 3370
rect 43429 3360 43463 3370
rect 12061 3336 27551 3346
rect 27613 3336 34871 3346
rect 34909 3336 43151 3346
rect 43213 3336 43271 3346
rect 43333 3336 43367 3346
rect 43405 3336 43559 3346
rect 43621 3336 43655 3346
rect 12013 3312 23687 3322
rect 23725 3312 31631 3322
rect 31645 3312 32207 3322
rect 32244 3312 35735 3322
rect 35773 3312 40223 3322
rect 40261 3312 43751 3322
rect 58920 3301 58930 3504
rect 59040 3301 59050 3479
rect 59640 3301 59650 3479
rect 59760 3301 59770 3479
rect 11965 3288 18095 3298
rect 18109 3288 43871 3298
rect 44029 3288 44063 3298
rect 11941 3264 43967 3274
rect 44005 3264 44183 3274
rect 66696 3274 66735 3282
rect 58800 3272 66735 3274
rect 58800 3264 66706 3272
rect 11917 3240 15071 3250
rect 15109 3240 44351 3250
rect 44413 3240 44471 3250
rect 11893 3216 22343 3226
rect 22381 3216 44567 3226
rect 11869 3192 12359 3202
rect 12397 3192 28079 3202
rect 28117 3192 28319 3202
rect 28333 3192 44711 3202
rect 11821 3168 13391 3178
rect 13429 3168 22775 3178
rect 22813 3168 44807 3178
rect 11797 3144 21479 3154
rect 21517 3144 32172 3154
rect 32221 3144 35039 3154
rect 35053 3144 38039 3154
rect 38053 3144 44903 3154
rect 11725 3120 12671 3130
rect 12733 3120 33431 3130
rect 33445 3120 36527 3130
rect 36565 3120 40631 3130
rect 40669 3120 44447 3130
rect 44485 3120 44999 3130
rect 11701 3096 20711 3106
rect 20749 3096 45119 3106
rect 11677 3072 11711 3082
rect 11749 3072 21935 3082
rect 21973 3072 30095 3082
rect 30133 3072 33671 3082
rect 33709 3072 45215 3082
rect 11629 3048 17135 3058
rect 17173 3048 31967 3058
rect 32005 3048 32207 3058
rect 32244 3048 33791 3058
rect 33829 3048 39335 3058
rect 39373 3048 45335 3058
rect 11605 3024 22679 3034
rect 22717 3024 27863 3034
rect 27925 3024 34415 3034
rect 34453 3024 45455 3034
rect 11581 3000 30575 3010
rect 30589 3000 32172 3010
rect 32221 3000 39239 3010
rect 39277 3000 45551 3010
rect 11533 2976 22175 2986
rect 22237 2976 30311 2986
rect 30349 2976 32375 2986
rect 32664 2976 32735 2986
rect 11461 2952 16703 2962
rect 32640 2962 32650 2975
rect 16741 2952 32650 2962
rect 11437 2928 16055 2938
rect 32664 2938 32674 2976
rect 32760 2976 32807 2986
rect 32760 2962 32770 2976
rect 33061 2976 33191 2986
rect 33205 2976 33863 2986
rect 33877 2976 34751 2986
rect 34765 2976 42551 2986
rect 42565 2976 44639 2986
rect 44653 2976 45647 2986
rect 16093 2928 32674 2938
rect 32736 2952 32770 2962
rect 11413 2904 32279 2914
rect 32317 2904 32639 2914
rect 32736 2914 32746 2952
rect 32821 2952 33263 2962
rect 33325 2952 45767 2962
rect 45829 2952 45863 2962
rect 45901 2952 45959 2962
rect 32760 2928 33335 2938
rect 32760 2917 32770 2928
rect 33373 2928 46055 2938
rect 46093 2928 46151 2938
rect 32677 2904 32746 2914
rect 33013 2904 33383 2914
rect 33421 2904 43487 2914
rect 43525 2904 46247 2914
rect 11365 2880 32255 2890
rect 32293 2880 46367 2890
rect 46909 2880 46943 2890
rect 11293 2856 16271 2866
rect 16309 2856 31943 2866
rect 31981 2856 32218 2866
rect 32244 2856 33623 2866
rect 11269 2832 12935 2842
rect 12973 2832 31919 2842
rect 32208 2842 32218 2856
rect 33637 2856 35927 2866
rect 35965 2856 40319 2866
rect 40357 2856 46463 2866
rect 46501 2856 46559 2866
rect 46885 2856 47063 2866
rect 47101 2856 47159 2866
rect 31957 2832 32172 2842
rect 32208 2832 43535 2842
rect 43573 2832 46679 2842
rect 46717 2832 46823 2842
rect 46861 2832 47255 2842
rect 47557 2832 47591 2842
rect 11245 2808 32447 2818
rect 32653 2808 39935 2818
rect 39973 2808 44327 2818
rect 44365 2808 44615 2818
rect 44629 2808 44951 2818
rect 44965 2808 45047 2818
rect 45061 2808 47375 2818
rect 47533 2808 47711 2818
rect 47749 2808 47831 2818
rect 47965 2808 47999 2818
rect 11197 2784 19367 2794
rect 19405 2784 29999 2794
rect 30037 2784 36407 2794
rect 36421 2784 47471 2794
rect 47509 2784 48119 2794
rect 11149 2760 27527 2770
rect 27565 2760 41783 2770
rect 41821 2760 48263 2770
rect 11053 2736 11231 2746
rect 11317 2736 24215 2746
rect 24301 2736 32207 2746
rect 32244 2736 37847 2746
rect 37909 2736 43679 2746
rect 43693 2736 43847 2746
rect 43885 2736 48383 2746
rect 48421 2736 48479 2746
rect 11029 2712 11879 2722
rect 11989 2712 18767 2722
rect 18805 2712 20927 2722
rect 20941 2712 25367 2722
rect 25405 2712 31511 2722
rect 31549 2712 36119 2722
rect 36157 2712 37919 2722
rect 37933 2712 38327 2722
rect 38341 2712 38783 2722
rect 38797 2712 42791 2722
rect 42829 2712 48575 2722
rect 10957 2688 31751 2698
rect 31789 2688 32172 2698
rect 32221 2688 33479 2698
rect 33517 2688 35495 2698
rect 35509 2688 44135 2698
rect 44149 2688 48671 2698
rect 48733 2688 48767 2698
rect 10861 2664 10895 2674
rect 10933 2664 31391 2674
rect 31453 2664 37199 2674
rect 37237 2664 43439 2674
rect 43477 2664 48863 2674
rect 10837 2640 12815 2650
rect 12853 2640 13367 2650
rect 13405 2640 32207 2650
rect 32244 2640 36959 2650
rect 36973 2640 39911 2650
rect 39925 2640 46751 2650
rect 46765 2640 48599 2650
rect 48613 2640 48959 2650
rect 10789 2616 41375 2626
rect 41413 2616 41543 2626
rect 41557 2616 42863 2626
rect 42877 2616 42959 2626
rect 42973 2616 44495 2626
rect 44509 2616 48359 2626
rect 48397 2616 49055 2626
rect 49093 2616 49151 2626
rect 10693 2592 12623 2602
rect 12661 2592 32172 2602
rect 32221 2592 36863 2602
rect 36901 2592 41591 2602
rect 41629 2592 42911 2602
rect 42949 2592 43343 2602
rect 43381 2592 47975 2602
rect 48013 2592 49247 2602
rect 10645 2568 15383 2578
rect 15421 2568 21383 2578
rect 21397 2568 24839 2578
rect 24877 2568 43799 2578
rect 43813 2568 46967 2578
rect 46981 2568 49343 2578
rect 10309 2544 10391 2554
rect 10621 2544 12527 2554
rect 12613 2544 21719 2554
rect 21757 2544 22487 2554
rect 22501 2544 24767 2554
rect 24781 2544 25079 2554
rect 25093 2544 26639 2554
rect 26653 2544 29975 2554
rect 30013 2544 34007 2554
rect 34045 2544 36647 2554
rect 36685 2544 39815 2554
rect 39829 2544 42503 2554
rect 42517 2544 48623 2554
rect 48637 2544 49439 2554
rect 10189 2520 10247 2530
rect 10285 2520 10487 2530
rect 10525 2520 11903 2530
rect 12037 2520 16487 2530
rect 16525 2520 23999 2530
rect 24037 2520 26999 2530
rect 27061 2520 29207 2530
rect 29221 2520 32999 2530
rect 33013 2520 49535 2530
rect 10141 2496 32207 2506
rect 32244 2496 38735 2506
rect 38773 2496 40847 2506
rect 40885 2496 46535 2506
rect 46573 2496 49631 2506
rect 10093 2472 11783 2482
rect 11845 2472 32639 2482
rect 32749 2472 32759 2482
rect 32989 2472 37367 2482
rect 37381 2472 41879 2482
rect 41917 2472 49727 2482
rect 10069 2448 32759 2458
rect 32989 2448 38927 2458
rect 38965 2448 41423 2458
rect 41437 2448 46031 2458
rect 46069 2448 49847 2458
rect 50029 2448 50063 2458
rect 9973 2424 11855 2434
rect 11893 2424 19487 2434
rect 19525 2424 22247 2434
rect 22285 2424 22871 2434
rect 22885 2424 42311 2434
rect 42349 2424 49967 2434
rect 50005 2424 50159 2434
rect 9949 2400 32172 2410
rect 32221 2400 45311 2410
rect 45349 2400 45623 2410
rect 45661 2400 50255 2410
rect 9925 2376 10847 2386
rect 10885 2376 17567 2386
rect 17605 2376 31823 2386
rect 31885 2376 48839 2386
rect 48877 2376 50351 2386
rect 9877 2352 14735 2362
rect 14773 2352 18263 2362
rect 18325 2352 32207 2362
rect 32244 2352 44543 2362
rect 44581 2352 50831 2362
rect 9853 2328 10583 2338
rect 10669 2328 20351 2338
rect 20413 2328 38279 2338
rect 38317 2328 46799 2338
rect 46837 2328 49271 2338
rect 49285 2328 50879 2338
rect 51037 2328 51071 2338
rect 9829 2304 13823 2314
rect 13837 2304 51167 2314
rect 51229 2304 51263 2314
rect 9781 2280 10127 2290
rect 10165 2280 23279 2290
rect 23389 2280 31727 2290
rect 31765 2280 35063 2290
rect 35101 2280 40031 2290
rect 40069 2280 47039 2290
rect 47077 2280 50087 2290
rect 50101 2280 51383 2290
rect 9709 2256 13679 2266
rect 13717 2256 14015 2266
rect 14053 2256 15167 2266
rect 15181 2256 15503 2266
rect 15517 2256 15719 2266
rect 15733 2256 15935 2266
rect 15949 2256 16151 2266
rect 16165 2256 16367 2266
rect 16381 2256 16583 2266
rect 16597 2256 16799 2266
rect 16813 2256 17015 2266
rect 17029 2256 17231 2266
rect 17245 2256 17351 2266
rect 17389 2256 32591 2266
rect 32917 2256 47687 2266
rect 47725 2256 49367 2266
rect 49381 2256 51503 2266
rect 8701 2232 8735 2242
rect 8773 2232 8831 2242
rect 9685 2232 11015 2242
rect 11077 2232 23807 2242
rect 23845 2232 24191 2242
rect 24205 2232 32183 2242
rect 32221 2232 35831 2242
rect 35869 2232 43943 2242
rect 43981 2232 48167 2242
rect 48181 2232 49751 2242
rect 49765 2232 51599 2242
rect 51685 2232 51719 2242
rect 8581 2208 8639 2218
rect 8677 2208 8927 2218
rect 8965 2208 9023 2218
rect 9661 2208 37703 2218
rect 37717 2208 41639 2218
rect 41653 2208 43295 2218
rect 43309 2208 51791 2218
rect 51805 2208 51863 2218
rect 8557 2184 9119 2194
rect 9181 2184 9215 2194
rect 9445 2184 9527 2194
rect 9565 2184 9839 2194
rect 9901 2184 14999 2194
rect 15061 2184 22199 2194
rect 22261 2184 35303 2194
rect 35341 2184 49223 2194
rect 49261 2184 51983 2194
rect 8317 2160 8399 2170
rect 8533 2160 9311 2170
rect 9349 2160 11159 2170
rect 11221 2160 18599 2170
rect 18661 2160 24551 2170
rect 24589 2160 41687 2170
rect 41725 2160 50039 2170
rect 50077 2160 52103 2170
rect 8221 2136 32207 2146
rect 32245 2136 45407 2146
rect 45421 2136 52199 2146
rect 8197 2112 14663 2122
rect 14701 2112 48095 2122
rect 48133 2112 49391 2122
rect 49405 2112 52319 2122
rect 8125 2088 8759 2098
rect 8797 2088 8879 2098
rect 8893 2088 9071 2098
rect 9085 2088 9263 2098
rect 9277 2088 12575 2098
rect 12637 2088 32903 2098
rect 32965 2088 34391 2098
rect 34405 2088 38399 2098
rect 38437 2088 39839 2098
rect 39877 2088 44039 2098
rect 44077 2088 49463 2098
rect 49477 2088 49895 2098
rect 49909 2088 52439 2098
rect 8101 2064 9335 2074
rect 9373 2064 10823 2074
rect 10861 2064 18623 2074
rect 18685 2064 23879 2074
rect 23917 2064 24887 2074
rect 24901 2064 24983 2074
rect 25021 2064 27167 2074
rect 27181 2064 30863 2074
rect 30877 2064 41759 2074
rect 41773 2064 51911 2074
rect 51925 2064 52559 2074
rect 8077 2040 22727 2050
rect 22741 2040 52679 2050
rect 8053 2016 8567 2026
rect 8605 2016 13559 2026
rect 13597 2016 20951 2026
rect 21013 2016 22943 2026
rect 22981 2016 37991 2026
rect 38005 2016 46991 2026
rect 47005 2016 47279 2026
rect 47293 2016 52799 2026
rect 8029 1992 8903 2002
rect 8917 1992 17879 2002
rect 17893 1992 32471 2002
rect 32605 1992 32663 2002
rect 32941 1992 43031 2002
rect 43069 1992 51143 2002
rect 51181 1992 52895 2002
rect 32880 1981 32890 1991
rect 7981 1968 9287 1978
rect 9301 1968 17663 1978
rect 17677 1968 32663 1978
rect 32893 1968 35711 1978
rect 35725 1968 40607 1978
rect 40621 1968 47303 1978
rect 47317 1968 51743 1978
rect 51757 1968 53015 1978
rect 7957 1944 10679 1954
rect 10717 1944 19271 1954
rect 19309 1944 48239 1954
rect 48277 1944 50135 1954
rect 50173 1944 53135 1954
rect 7909 1920 11039 1930
rect 11101 1920 13871 1930
rect 13909 1920 14111 1930
rect 14125 1920 15239 1930
rect 15253 1920 15575 1930
rect 15589 1920 15791 1930
rect 15805 1920 16007 1930
rect 16021 1920 16223 1930
rect 16237 1920 16439 1930
rect 16453 1920 16655 1930
rect 16669 1920 16871 1930
rect 16885 1920 16919 1930
rect 16957 1920 19247 1930
rect 19285 1920 19799 1930
rect 19837 1920 24263 1930
rect 24325 1920 49127 1930
rect 49165 1920 53231 1930
rect 7885 1896 12263 1906
rect 12301 1896 26015 1906
rect 26029 1896 35615 1906
rect 35629 1896 37607 1906
rect 37621 1896 38255 1906
rect 38269 1896 47111 1906
rect 47125 1896 50303 1906
rect 50317 1896 51767 1906
rect 51781 1896 53375 1906
rect 7837 1872 10751 1882
rect 10813 1872 18551 1882
rect 18589 1872 22391 1882
rect 22453 1872 33335 1882
rect 33349 1872 38351 1882
rect 38365 1872 44927 1882
rect 44941 1872 47207 1882
rect 47221 1872 47879 1882
rect 47893 1872 48431 1882
rect 48445 1872 51647 1882
rect 51661 1872 53471 1882
rect 7741 1848 8543 1858
rect 8581 1848 11255 1858
rect 11341 1848 11687 1858
rect 11725 1848 28583 1858
rect 28621 1848 30815 1858
rect 30829 1848 30935 1858
rect 30949 1848 31079 1858
rect 31093 1848 31319 1858
rect 31333 1848 31535 1858
rect 31573 1848 37631 1858
rect 37645 1848 43127 1858
rect 43165 1848 44231 1858
rect 44245 1848 44423 1858
rect 44437 1848 53591 1858
rect 7597 1824 9959 1834
rect 9997 1824 36767 1834
rect 36805 1824 50327 1834
rect 50365 1824 51239 1834
rect 51277 1824 53639 1834
rect 7189 1800 11615 1810
rect 11653 1800 24239 1810
rect 24277 1800 36023 1810
rect 36061 1800 41063 1810
rect 41101 1800 44783 1810
rect 44821 1800 45935 1810
rect 45973 1800 53663 1810
rect 6973 1776 32591 1786
rect 32773 1776 44159 1786
rect 44197 1776 51695 1786
rect 51733 1776 53687 1786
rect 6925 1752 8063 1762
rect 8149 1752 12239 1762
rect 12277 1752 18335 1762
rect 18373 1752 33983 1762
rect 33997 1752 40679 1762
rect 40693 1752 42623 1762
rect 42637 1752 46223 1762
rect 46261 1752 50855 1762
rect 50893 1752 53711 1762
rect 6277 1728 6359 1738
rect 6397 1728 6455 1738
rect 6565 1728 22199 1738
rect 22213 1728 38159 1738
rect 38197 1728 40535 1738
rect 40573 1728 48455 1738
rect 48493 1728 49175 1738
rect 49189 1728 50183 1738
rect 50197 1728 53783 1738
rect 6085 1704 6143 1714
rect 6181 1704 10511 1714
rect 10549 1704 11663 1714
rect 11701 1704 11807 1714
rect 11869 1704 11927 1714
rect 12085 1704 20207 1714
rect 20245 1704 36215 1714
rect 36229 1704 39575 1714
rect 39589 1704 43895 1714
rect 43909 1704 48791 1714
rect 48805 1704 49007 1714
rect 49021 1704 49103 1714
rect 49117 1704 51311 1714
rect 51325 1704 51887 1714
rect 51901 1704 52031 1714
rect 52045 1704 53903 1714
rect 5845 1680 5927 1690
rect 5965 1680 9623 1690
rect 9733 1680 21263 1690
rect 21301 1680 24527 1690
rect 24565 1680 33119 1690
rect 33157 1680 45743 1690
rect 45781 1680 49703 1690
rect 49741 1680 53999 1690
rect 5797 1656 36431 1666
rect 36469 1656 54095 1666
rect 5773 1632 11855 1642
rect 11917 1632 13463 1642
rect 13501 1632 22559 1642
rect 22597 1632 26447 1642
rect 26485 1632 42575 1642
rect 42613 1632 44975 1642
rect 45013 1632 46583 1642
rect 46597 1632 52415 1642
rect 52453 1632 52943 1642
rect 52957 1632 54119 1642
rect 5725 1608 26855 1618
rect 26917 1608 51191 1618
rect 51205 1608 51407 1618
rect 51421 1608 54215 1618
rect 5701 1584 11111 1594
rect 11125 1584 11999 1594
rect 12133 1584 27455 1594
rect 27493 1584 32591 1594
rect 32677 1584 53615 1594
rect 53677 1584 54263 1594
rect 5677 1560 9863 1570
rect 9973 1560 14567 1570
rect 14605 1560 21623 1570
rect 21661 1560 53111 1570
rect 53149 1560 54287 1570
rect 5653 1536 8039 1546
rect 8077 1536 11351 1546
rect 11389 1536 11591 1546
rect 11629 1536 20183 1546
rect 20197 1536 38591 1546
rect 38605 1536 44303 1546
rect 44317 1536 46727 1546
rect 46741 1536 48911 1546
rect 48925 1536 52631 1546
rect 52645 1536 54311 1546
rect 5605 1512 9167 1522
rect 9205 1512 18287 1522
rect 18349 1512 24503 1522
rect 24541 1512 37007 1522
rect 37045 1512 40007 1522
rect 40021 1512 40079 1522
rect 40093 1512 43079 1522
rect 43093 1512 47567 1522
rect 47605 1512 54407 1522
rect 5557 1488 9407 1498
rect 9469 1488 15431 1498
rect 15445 1488 22511 1498
rect 22525 1488 43583 1498
rect 43597 1488 54551 1498
rect 5533 1464 6959 1474
rect 6997 1464 9647 1474
rect 9757 1464 12911 1474
rect 12925 1464 14375 1474
rect 14413 1464 37247 1474
rect 37261 1464 43631 1474
rect 43669 1464 49415 1474
rect 49453 1464 51287 1474
rect 51301 1464 51431 1474
rect 51445 1464 52007 1474
rect 52021 1464 54671 1474
rect 5509 1440 13271 1450
rect 13309 1440 32567 1450
rect 32677 1440 37655 1450
rect 37693 1440 44831 1450
rect 44845 1440 45383 1450
rect 45397 1440 52991 1450
rect 53029 1440 54791 1450
rect 5485 1416 7943 1426
rect 8005 1416 10775 1426
rect 10837 1416 18407 1426
rect 18445 1416 28751 1426
rect 28789 1416 30119 1426
rect 30157 1416 36743 1426
rect 36757 1416 38999 1426
rect 39013 1416 42983 1426
rect 42997 1416 44735 1426
rect 44749 1416 45719 1426
rect 45733 1416 45791 1426
rect 45805 1416 45911 1426
rect 45925 1416 52871 1426
rect 52909 1416 54239 1426
rect 54277 1416 54335 1426
rect 54349 1416 54887 1426
rect 5461 1392 10943 1402
rect 10981 1392 20375 1402
rect 20437 1392 26303 1402
rect 26341 1392 30239 1402
rect 30277 1392 53159 1402
rect 53173 1392 54983 1402
rect 5413 1368 5471 1378
rect 5581 1368 32735 1378
rect 32773 1368 37751 1378
rect 37789 1368 41975 1378
rect 42013 1368 49511 1378
rect 49549 1368 55079 1378
rect 5389 1344 5663 1354
rect 5749 1344 12047 1354
rect 12157 1344 18911 1354
rect 18973 1344 27959 1354
rect 27997 1344 28079 1354
rect 28093 1344 34319 1354
rect 34357 1344 43823 1354
rect 43837 1344 55151 1354
rect 5269 1320 5327 1330
rect 5365 1320 5759 1330
rect 5821 1320 15359 1330
rect 15397 1320 45983 1330
rect 45997 1320 48887 1330
rect 48901 1320 54647 1330
rect 54685 1320 54815 1330
rect 54829 1320 54911 1330
rect 54925 1320 55295 1330
rect 5245 1296 11567 1306
rect 11605 1296 12551 1306
rect 12589 1296 25463 1306
rect 25501 1296 27359 1306
rect 27373 1296 29183 1306
rect 29197 1296 34607 1306
rect 34645 1296 36479 1306
rect 36493 1296 39023 1306
rect 39061 1296 39071 1306
rect 39085 1296 45143 1306
rect 45157 1296 48935 1306
rect 48973 1296 49559 1306
rect 49573 1296 49655 1306
rect 49669 1296 55391 1306
rect 5149 1272 7799 1282
rect 7861 1272 35639 1282
rect 35677 1272 41279 1282
rect 41317 1272 42263 1282
rect 42277 1272 45095 1282
rect 45133 1272 51047 1282
rect 51085 1272 55535 1282
rect 5125 1248 8279 1258
rect 8341 1248 9911 1258
rect 10021 1248 37823 1258
rect 37885 1248 40295 1258
rect 40309 1248 52055 1258
rect 52069 1248 55631 1258
rect 5053 1224 7895 1234
rect 7933 1224 30215 1234
rect 30253 1224 38063 1234
rect 38101 1224 42431 1234
rect 42469 1224 49607 1234
rect 49645 1224 53447 1234
rect 53485 1224 55007 1234
rect 55021 1224 55343 1234
rect 55357 1224 55751 1234
rect 5005 1200 6239 1210
rect 6301 1200 7871 1210
rect 7909 1200 9695 1210
rect 9792 1200 32423 1210
rect 4933 1176 8303 1186
rect 9768 1186 9778 1199
rect 9792 1189 9802 1200
rect 32461 1200 37559 1210
rect 37597 1200 42095 1210
rect 42133 1200 47807 1210
rect 47845 1200 49871 1210
rect 49885 1200 55055 1210
rect 55093 1200 55103 1210
rect 55117 1200 55847 1210
rect 8365 1176 9778 1186
rect 9853 1176 33527 1186
rect 33541 1176 34175 1186
rect 34189 1176 34487 1186
rect 34501 1176 34559 1186
rect 34573 1176 36239 1186
rect 36277 1176 43727 1186
rect 43765 1176 47231 1186
rect 47269 1176 50111 1186
rect 50125 1176 53663 1186
rect 53725 1176 54767 1186
rect 54805 1176 55775 1186
rect 55789 1176 55943 1186
rect 56053 1176 56471 1186
rect 4909 1152 5543 1162
rect 5629 1152 9431 1162
rect 9493 1152 12479 1162
rect 12493 1152 14255 1162
rect 14293 1152 54143 1162
rect 54157 1152 56663 1162
rect 4861 1128 6551 1138
rect 6589 1128 7823 1138
rect 7885 1128 22319 1138
rect 22357 1128 27239 1138
rect 27277 1128 30719 1138
rect 30733 1128 36311 1138
rect 36325 1128 36935 1138
rect 36949 1128 41567 1138
rect 41581 1128 46007 1138
rect 46021 1128 46103 1138
rect 46117 1128 46295 1138
rect 46309 1128 51575 1138
rect 51613 1128 55271 1138
rect 55309 1128 55463 1138
rect 55477 1128 55871 1138
rect 55885 1128 56687 1138
rect 4789 1104 6263 1114
rect 6325 1104 24479 1114
rect 24517 1104 51839 1114
rect 51877 1104 56783 1114
rect 4765 1080 11735 1090
rect 11773 1080 18935 1090
rect 18997 1080 26351 1090
rect 26437 1080 39623 1090
rect 39661 1080 42743 1090
rect 42757 1080 47447 1090
rect 47485 1080 52823 1090
rect 52837 1080 53578 1090
rect 53568 1069 53578 1080
rect 53653 1080 56879 1090
rect 4741 1056 21719 1066
rect 21733 1056 28799 1066
rect 28813 1056 30599 1066
rect 30613 1056 39983 1066
rect 39997 1056 40703 1066
rect 40717 1056 41255 1066
rect 41269 1056 47663 1066
rect 47677 1056 53543 1066
rect 53592 1066 53602 1079
rect 53592 1056 56711 1066
rect 56725 1056 56975 1066
rect 4717 1032 4895 1042
rect 4957 1032 5711 1042
rect 5773 1032 9551 1042
rect 9589 1032 11015 1042
rect 11029 1032 12335 1042
rect 12373 1032 14471 1042
rect 14509 1032 33239 1042
rect 33253 1032 36983 1042
rect 36997 1032 40919 1042
rect 40933 1032 47423 1042
rect 47437 1032 47759 1042
rect 47773 1032 53327 1042
rect 53341 1032 57095 1042
rect 4693 1008 11903 1018
rect 11941 1008 23639 1018
rect 23677 1008 41951 1018
rect 41965 1008 44855 1018
rect 44869 1008 51815 1018
rect 51829 1008 53303 1018
rect 53317 1008 53855 1018
rect 53869 1008 54695 1018
rect 54709 1008 57191 1018
rect 4597 984 4919 994
rect 4981 984 5039 994
rect 5077 984 8951 994
rect 8989 984 9167 994
rect 9181 984 9359 994
rect 9397 984 32807 994
rect 32869 984 47135 994
rect 47173 984 47183 994
rect 47197 984 51479 994
rect 51517 984 54191 994
rect 54229 984 57250 994
rect 4549 960 5087 970
rect 5173 960 8111 970
rect 8173 960 9935 970
rect 10045 960 19631 970
rect 19669 960 24383 970
rect 24421 960 31055 970
rect 31069 960 32807 970
rect 32832 970 32842 983
rect 32832 960 46127 970
rect 46165 960 46175 970
rect 46189 960 52295 970
rect 52333 960 56759 970
rect 56797 960 57215 970
rect 57240 970 57250 984
rect 57240 960 57287 970
rect 4189 936 5399 946
rect 5437 936 10919 946
rect 10957 936 20399 946
rect 20509 936 21839 946
rect 21853 936 22943 946
rect 22957 936 23135 946
rect 23173 936 41927 946
rect 41941 936 49943 946
rect 49981 936 50447 946
rect 50461 936 56447 946
rect 56485 936 57383 946
rect 3973 912 53639 922
rect 53701 912 55559 922
rect 55573 912 57407 922
rect 3925 888 6047 898
rect 6109 888 18023 898
rect 18037 888 32711 898
rect 32749 888 48647 898
rect 48685 888 57479 898
rect 3397 864 3455 874
rect 3565 864 8495 874
rect 8557 864 10055 874
rect 10117 864 12695 874
rect 12757 864 13175 874
rect 13189 864 21047 874
rect 21109 864 21215 874
rect 21229 864 25247 874
rect 25285 864 28871 874
rect 28885 864 32831 874
rect 32869 864 35591 874
rect 35605 864 35687 874
rect 35701 864 35783 874
rect 35797 864 35879 874
rect 35893 864 36599 874
rect 36613 864 39143 874
rect 39181 864 40127 874
rect 40165 864 49319 874
rect 49357 864 51959 874
rect 51997 864 53711 874
rect 53725 864 57599 874
rect 3373 840 5999 850
rect 6013 840 8807 850
rect 8821 840 11951 850
rect 12013 840 22415 850
rect 22477 840 26063 850
rect 26077 840 37079 850
rect 37093 840 37175 850
rect 37189 840 39407 850
rect 39421 840 40199 850
rect 40213 840 48695 850
rect 48709 840 51119 850
rect 51133 840 53519 850
rect 53557 840 57503 850
rect 57517 840 57695 850
rect 3325 816 11183 826
rect 11245 816 11447 826
rect 11485 816 27311 826
rect 27349 816 29159 826
rect 29173 816 38447 826
rect 38461 816 40967 826
rect 41005 816 46439 826
rect 46477 816 46919 826
rect 46957 816 49199 826
rect 49213 816 56639 826
rect 56677 816 57815 826
rect 3205 792 3239 802
rect 3277 792 4679 802
rect 4813 792 8471 802
rect 8485 792 10991 802
rect 11005 792 11759 802
rect 11797 792 32783 802
rect 32845 792 42887 802
rect 42901 792 44087 802
rect 44101 792 52607 802
rect 52621 792 52727 802
rect 52741 792 57575 802
rect 57613 792 57863 802
rect 3181 768 5375 778
rect 5413 768 9719 778
rect 9781 768 18527 778
rect 18565 768 29855 778
rect 29869 768 37799 778
rect 37837 768 41111 778
rect 41125 768 43247 778
rect 43285 768 45575 778
rect 45589 768 49823 778
rect 49861 768 56663 778
rect 56701 768 57887 778
rect 3085 744 5255 754
rect 5293 744 7727 754
rect 7765 744 18239 754
rect 18253 744 19055 754
rect 19093 744 23543 754
rect 23581 744 26207 754
rect 26221 744 27791 754
rect 27805 744 28175 754
rect 28189 744 28295 754
rect 28309 744 28391 754
rect 28405 744 33911 754
rect 33949 744 44255 754
rect 44269 744 52367 754
rect 52381 744 56855 754
rect 56893 744 57935 754
rect 3037 720 3335 730
rect 3408 720 8519 730
rect 3384 706 3394 719
rect 3408 709 3418 720
rect 8629 720 14927 730
rect 14965 720 21407 730
rect 21421 720 23279 730
rect 23293 720 27143 730
rect 27157 720 34703 730
rect 34717 720 36191 730
rect 36205 720 38567 730
rect 38581 720 41471 730
rect 41509 720 45263 730
rect 45277 720 49031 730
rect 49069 720 56615 730
rect 56653 720 56735 730
rect 56749 720 56831 730
rect 56845 720 57719 730
rect 57733 720 58042 730
rect 3013 696 3394 706
rect 3445 696 4703 706
rect 4837 696 5447 706
rect 5485 696 7871 706
rect 7957 696 11399 706
rect 11461 696 13247 706
rect 13261 696 14447 706
rect 14485 696 21527 706
rect 21589 696 30215 706
rect 30229 696 32567 706
rect 32581 696 42143 706
rect 42157 696 44879 706
rect 44917 696 46775 706
rect 46789 696 53759 706
rect 53797 696 55511 706
rect 55549 696 58007 706
rect 58032 706 58042 720
rect 58032 696 58127 706
rect 2989 672 3191 682
rect 3229 672 9455 682
rect 9517 672 12503 682
rect 12517 672 46607 682
rect 46621 672 50207 682
rect 50221 672 54167 682
rect 54181 672 56591 682
rect 56605 672 57743 682
rect 57757 672 58223 682
rect 2941 648 7175 658
rect 7213 648 11255 658
rect 11365 648 19079 658
rect 19189 648 26399 658
rect 26461 648 37943 658
rect 37981 648 38807 658
rect 38821 648 40103 658
rect 40117 648 45503 658
rect 45517 648 47903 658
rect 47917 648 49295 658
rect 49309 648 54839 658
rect 54853 648 57431 658
rect 57445 648 58055 658
rect 58069 648 58319 658
rect 2917 624 3167 634
rect 3205 624 3551 634
rect 3589 624 5639 634
rect 5677 624 24359 634
rect 24397 624 25103 634
rect 25117 624 26543 634
rect 26557 624 36839 634
rect 36853 624 40823 634
rect 40837 624 52703 634
rect 52717 624 57911 634
rect 57949 624 58391 634
rect 2893 600 2975 610
rect 3061 600 5351 610
rect 5389 600 5951 610
rect 5989 600 8447 610
rect 8461 600 10607 610
rect 10693 600 21551 610
rect 21637 600 23399 610
rect 23437 600 26375 610
rect 26413 600 33263 610
rect 33301 600 37319 610
rect 37357 600 45527 610
rect 45565 600 50807 610
rect 50845 600 57359 610
rect 57421 600 57455 610
rect 57493 600 58439 610
rect 2869 576 2927 586
rect 2965 576 4775 586
rect 4885 576 5783 586
rect 5869 576 8087 586
rect 8125 576 8183 586
rect 8245 576 10271 586
rect 10333 576 12983 586
rect 13045 576 19151 586
rect 19213 576 27215 586
rect 27253 576 32783 586
rect 32821 576 34367 586
rect 34381 576 38975 586
rect 38989 576 39383 586
rect 39397 576 45191 586
rect 45229 576 54263 586
rect 54301 576 57071 586
rect 57109 576 58175 586
rect 58189 576 58463 586
rect 58477 576 58559 586
rect 2808 552 5207 562
rect 2808 538 2818 552
rect 5269 552 6383 562
rect 6421 552 13967 562
rect 13981 552 32615 562
rect 32653 552 48047 562
rect 48061 552 52775 562
rect 52813 552 53831 562
rect 53845 552 55679 562
rect 55693 552 58655 562
rect 2760 528 2818 538
rect 2760 493 2770 528
rect 2845 528 4799 538
rect 4909 528 12791 538
rect 12829 528 20807 538
rect 20845 528 23207 538
rect 23221 528 23591 538
rect 23605 528 23663 538
rect 23701 528 23807 538
rect 23821 528 28487 538
rect 28501 528 28583 538
rect 28597 528 28679 538
rect 28693 528 28967 538
rect 28981 528 29279 538
rect 29317 528 33767 538
rect 33781 528 42191 538
rect 42229 528 47351 538
rect 47389 528 47399 538
rect 47413 528 52175 538
rect 52213 528 55703 538
rect 55717 528 57047 538
rect 57061 528 57407 538
rect 57421 528 57959 538
rect 57973 528 58151 538
rect 58165 528 58487 538
rect 58501 528 58727 538
rect 2784 504 4751 514
rect 2784 493 2794 504
rect 4789 504 10175 514
rect 10213 504 12167 514
rect 12205 504 23111 514
rect 23149 504 54959 514
rect 54997 504 55727 514
rect 55765 504 57023 514
rect 57037 504 58786 514
rect 58776 493 58786 504
rect 58800 493 58810 3264
rect 2821 480 5831 490
rect 5893 480 23471 490
rect 23485 480 32399 490
rect 32437 480 39743 490
rect 39781 480 43919 490
rect 43933 480 53351 490
rect 53389 480 54071 490
rect 54109 480 57263 490
rect 57301 480 58751 490
rect 2749 456 8015 466
rect 8053 456 21071 466
rect 21133 456 29063 466
rect 29077 456 44111 466
rect 44125 456 45695 466
rect 45709 456 46271 466
rect 46285 456 51095 466
rect 51109 456 53399 466
rect 53413 456 54527 466
rect 54565 456 56807 466
rect 56821 456 58823 466
rect 58920 445 58930 3239
rect 2725 432 2855 442
rect 2928 432 5231 442
rect 2904 418 2914 431
rect 2928 421 2938 432
rect 5317 432 5591 442
rect 5653 432 18863 442
rect 18901 432 33215 442
rect 33229 432 39527 442
rect 39565 432 42383 442
rect 42397 432 45431 442
rect 45469 432 45839 442
rect 45877 432 52487 442
rect 52501 432 54863 442
rect 54901 432 58415 442
rect 58453 432 58871 442
rect 2677 408 2914 418
rect 2989 408 4943 418
rect 5029 408 6071 418
rect 6133 408 6215 418
rect 6229 408 6431 418
rect 6445 408 7775 418
rect 7789 408 8207 418
rect 8269 408 12047 418
rect 12061 408 21983 418
rect 21997 408 36335 418
rect 36373 408 36383 418
rect 36397 408 36719 418
rect 36733 408 36815 418
rect 36829 408 38231 418
rect 38245 408 38687 418
rect 38701 408 42671 418
rect 42709 408 50231 418
rect 50269 408 51335 418
rect 51349 408 53087 418
rect 53101 408 53279 418
rect 53293 408 54935 418
rect 54949 408 58943 418
rect 59040 397 59050 3239
rect 59640 3061 59650 3239
rect 59760 3061 59770 3239
rect 66696 3034 66735 3042
rect 59160 3032 66735 3034
rect 59160 3024 66706 3032
rect 2653 384 9095 394
rect 9109 384 9815 394
rect 9877 384 10007 394
rect 10069 384 32519 394
rect 32557 384 37439 394
rect 37477 384 44687 394
rect 44725 384 55607 394
rect 55645 384 58079 394
rect 58093 384 58247 394
rect 58261 384 58799 394
rect 58837 384 58847 394
rect 58885 384 58991 394
rect 2616 360 7967 370
rect 2616 349 2626 360
rect 8029 360 8135 370
rect 8197 360 10079 370
rect 10141 360 11519 370
rect 11557 360 40511 370
rect 40525 360 53927 370
rect 53941 360 57671 370
rect 57709 360 57839 370
rect 57877 360 58631 370
rect 58669 360 59074 370
rect 2688 336 5783 346
rect 2640 322 2650 335
rect 2688 325 2698 336
rect 5797 336 9863 346
rect 9925 336 21455 346
rect 21493 336 26783 346
rect 26821 336 28199 346
rect 28213 336 47327 346
rect 47341 336 49487 346
rect 49501 336 56951 346
rect 56989 336 58967 346
rect 59005 336 59039 346
rect 59064 346 59074 360
rect 59160 349 59170 3024
rect 59640 2821 59650 2999
rect 59760 2821 59770 2999
rect 66696 2794 66735 2802
rect 59520 2792 66735 2794
rect 59520 2784 66706 2792
rect 59520 2341 59530 2784
rect 59640 2341 59650 2759
rect 59760 2341 59770 2759
rect 66696 2554 66735 2562
rect 59880 2552 66735 2554
rect 59880 2544 66706 2552
rect 59880 2341 59890 2544
rect 66696 2314 66735 2322
rect 59400 2312 66735 2314
rect 59400 2304 66706 2312
rect 59400 2101 59410 2304
rect 59520 2101 59530 2279
rect 59640 2101 59650 2279
rect 59760 2101 59770 2279
rect 59880 2101 59890 2279
rect 66696 2074 66735 2082
rect 59280 2072 66735 2074
rect 59280 2064 66706 2072
rect 59064 336 59111 346
rect 2581 312 2650 322
rect 2856 312 4175 322
rect 2712 298 2722 311
rect 2856 301 2866 312
rect 4213 312 5111 322
rect 5197 312 8687 322
rect 8725 312 9671 322
rect 9709 312 13439 322
rect 13477 312 14951 322
rect 14989 312 15623 322
rect 15661 312 24119 322
rect 24157 312 35903 322
rect 35917 312 46391 322
rect 46405 312 52535 322
rect 52573 312 57791 322
rect 57829 312 59194 322
rect 2557 288 2722 298
rect 2917 288 20975 298
rect 21037 288 38495 298
rect 38533 288 50279 298
rect 50293 288 54383 298
rect 54421 288 58295 298
rect 58333 288 58607 298
rect 58621 288 59159 298
rect 59184 298 59194 312
rect 59280 301 59290 2064
rect 59184 288 59231 298
rect 2533 264 2999 274
rect 3109 264 4583 274
rect 4621 264 10439 274
rect 10477 264 10631 274
rect 10741 264 11543 274
rect 11581 264 38711 274
rect 38725 264 41351 274
rect 41365 264 48983 274
rect 48997 264 49775 274
rect 49789 264 51527 274
rect 51541 264 54095 274
rect 54133 264 55823 274
rect 55861 264 58103 274
rect 58141 264 59303 274
rect 59400 253 59410 2039
rect 2389 240 2759 250
rect 3013 240 5519 250
rect 5557 240 5687 250
rect 5725 240 13367 250
rect 13381 240 14639 250
rect 14677 240 23015 250
rect 23077 240 46511 250
rect 46525 240 47639 250
rect 47653 240 48287 250
rect 48301 240 48503 250
rect 48517 240 52247 250
rect 52261 240 57167 250
rect 57229 240 57335 250
rect 57397 240 59351 250
rect 2328 216 2567 226
rect 2328 202 2338 216
rect 2605 216 5495 226
rect 5533 216 7583 226
rect 7621 216 35999 226
rect 36013 216 39311 226
rect 39325 216 43223 226
rect 43237 216 46199 226
rect 46213 216 47615 226
rect 47629 216 48191 226
rect 48205 216 48311 226
rect 48325 216 48527 226
rect 48541 216 54479 226
rect 54493 216 54575 226
rect 54589 216 57647 226
rect 57661 216 58367 226
rect 58405 216 59087 226
rect 59125 216 59423 226
rect 59520 205 59530 2039
rect 1981 192 2338 202
rect 2365 192 2543 202
rect 2581 192 2687 202
rect 2725 192 14231 202
rect 14269 192 14375 202
rect 14389 192 14783 202
rect 14797 192 14855 202
rect 14893 192 21767 202
rect 21781 192 23951 202
rect 23965 192 24791 202
rect 24805 192 31295 202
rect 31309 192 38015 202
rect 38029 192 46655 202
rect 46693 192 48551 202
rect 48589 192 48743 202
rect 48781 192 48815 202
rect 48829 192 50999 202
rect 51013 192 52127 202
rect 52141 192 53879 202
rect 53917 192 54455 202
rect 54469 192 55223 202
rect 55237 192 57311 202
rect 57349 192 57623 202
rect 57637 192 58343 202
rect 58357 192 58703 202
rect 58789 192 59327 202
rect 59365 192 59471 202
rect 1765 168 3359 178
rect 3397 168 4991 178
rect 5053 168 8663 178
rect 8701 168 8975 178
rect 9013 168 11279 178
rect 11413 168 11423 178
rect 11509 168 15023 178
rect 15085 168 18863 178
rect 18877 168 20711 178
rect 20725 168 20807 178
rect 20821 168 21287 178
rect 21325 168 28511 178
rect 28525 168 42527 178
rect 42541 168 45479 178
rect 45493 168 46415 178
rect 46429 168 53207 178
rect 53245 168 53975 178
rect 54013 168 55919 178
rect 55957 168 57239 178
rect 57253 168 59207 178
rect 59245 168 59543 178
rect 59640 157 59650 2039
rect 1717 144 3071 154
rect 3133 144 3263 154
rect 3301 144 3911 154
rect 3949 144 6911 154
rect 6949 144 44759 154
rect 44773 144 45023 154
rect 45037 144 54599 154
rect 54613 144 55247 154
rect 55261 144 55319 154
rect 55333 144 57143 154
rect 57205 144 59591 154
rect 1344 120 1751 130
rect 1344 106 1354 120
rect 1789 120 1967 130
rect 2005 120 2519 130
rect 2557 120 2879 130
rect 3085 120 4847 130
rect 4933 120 10295 130
rect 10357 120 13007 130
rect 13069 120 21191 130
rect 21205 120 24407 130
rect 24445 120 28895 130
rect 28909 120 29087 130
rect 29101 120 34103 130
rect 34141 120 36071 130
rect 36085 120 38831 130
rect 38869 120 52655 130
rect 52693 120 54047 130
rect 54085 120 57527 130
rect 57541 120 57863 130
rect 57901 120 59447 130
rect 59485 120 59663 130
rect 59760 109 59770 2039
rect 1141 96 1354 106
rect 1381 96 1703 106
rect 1741 96 3959 106
rect 3997 96 4727 106
rect 4765 96 5495 106
rect 5509 96 6167 106
rect 6205 96 14543 106
rect 14581 96 20903 106
rect 20917 96 46343 106
rect 46381 96 51359 106
rect 51397 96 54287 106
rect 54325 96 55439 106
rect 55453 96 57119 106
rect 57133 96 58679 106
rect 58741 96 59711 106
rect 59880 85 59890 2039
rect 757 72 4535 82
rect 4573 72 18743 82
rect 18781 72 25175 82
rect 25189 72 26303 82
rect 26317 72 27455 82
rect 27469 72 30839 82
rect 30853 72 32063 82
rect 32077 72 33311 82
rect 33325 72 33743 82
rect 33757 72 33839 82
rect 33853 72 34247 82
rect 34261 72 38639 82
rect 38677 72 40751 82
rect 40789 72 52079 82
rect 52117 72 56903 82
rect 56917 72 58199 82
rect 58237 72 58271 82
rect 58285 72 58919 82
rect 58957 72 59279 82
rect 59317 72 59639 82
rect 59677 72 59807 82
rect 504 48 2375 58
rect 504 34 514 48
rect 2413 48 2615 58
rect 2653 48 3023 58
rect 3157 48 23519 58
rect 23557 48 24143 58
rect 24181 48 26783 58
rect 26797 48 27983 58
rect 28021 48 42047 58
rect 42061 48 49679 58
rect 49693 48 53063 58
rect 53077 48 58535 58
rect 58573 48 58583 58
rect 58597 48 59399 58
rect 59437 48 59567 58
rect 59605 48 59914 58
rect 120 24 514 34
rect 528 24 1127 34
rect 120 13 130 24
rect 528 13 538 24
rect 1152 24 2735 34
rect 1152 13 1162 24
rect 2760 24 12095 34
rect 2760 13 2770 24
rect 12168 24 20447 34
rect 12120 13 12130 23
rect 12144 13 12154 23
rect 12168 13 12178 24
rect 20520 24 59519 34
rect 20472 13 20482 23
rect 20496 13 20506 23
rect 20520 13 20530 24
rect 28992 13 29002 24
rect 34272 13 34282 24
rect 37272 13 37282 24
rect 49584 13 49594 24
rect 54720 13 54730 24
rect 55032 13 55042 24
rect 55800 13 55810 24
rect 55896 13 55906 24
rect 57984 13 57994 24
rect 59557 24 59698 34
rect 59520 13 59530 23
rect 59688 13 59698 24
rect 59725 24 59879 34
rect 59904 34 59914 48
rect 59904 24 59938 34
rect 59880 13 59890 23
rect 59928 13 59938 24
<< m2contact >>
rect 32255 31583 32269 31597
rect 32255 31535 32269 31549
rect 32255 30791 32269 30805
rect 32255 30743 32269 30757
rect 32255 30023 32269 30037
rect 32279 30023 32293 30037
rect 32255 29975 32269 29989
rect 32279 29975 32293 29989
rect 32255 29279 32269 29293
rect 32279 29279 32293 29293
rect 32303 29279 32317 29293
rect 32255 29231 32269 29245
rect 32279 29231 32293 29245
rect 32303 29231 32317 29245
rect 32255 28319 32269 28333
rect 32279 28319 32293 28333
rect 32303 28319 32317 28333
rect 32327 28319 32341 28333
rect 32255 28271 32269 28285
rect 32279 28271 32293 28285
rect 32303 28271 32317 28285
rect 32327 28271 32341 28285
rect 32255 27575 32269 27589
rect 32279 27575 32293 27589
rect 32303 27575 32317 27589
rect 32327 27575 32341 27589
rect 32351 27575 32365 27589
rect 32255 27527 32269 27541
rect 32279 27527 32293 27541
rect 32303 27527 32317 27541
rect 32327 27527 32341 27541
rect 32351 27527 32365 27541
rect 32255 27407 32269 27421
rect 32279 27407 32293 27421
rect 32303 27407 32317 27421
rect 32327 27407 32341 27421
rect 32351 27407 32365 27421
rect 32375 27407 32389 27421
rect 32255 27359 32269 27373
rect 32279 27359 32293 27373
rect 32303 27359 32317 27373
rect 32327 27359 32341 27373
rect 32351 27359 32365 27373
rect 32375 27359 32389 27373
rect 32255 17999 32269 18013
rect 32279 17999 32293 18013
rect 32303 17999 32317 18013
rect 32327 17999 32341 18013
rect 32351 17999 32365 18013
rect 32375 17999 32389 18013
rect 32399 17999 32413 18013
rect 32255 17951 32269 17965
rect 32279 17951 32293 17965
rect 32303 17951 32317 17965
rect 32327 17951 32341 17965
rect 32351 17951 32365 17965
rect 32375 17951 32389 17965
rect 32399 17951 32413 17965
rect 32255 17807 32269 17821
rect 32279 17807 32293 17821
rect 32303 17807 32317 17821
rect 32327 17807 32341 17821
rect 32351 17807 32365 17821
rect 32375 17807 32389 17821
rect 32399 17807 32413 17821
rect 32423 17807 32437 17821
rect 32255 17759 32269 17773
rect 32279 17759 32293 17773
rect 32303 17759 32317 17773
rect 32327 17759 32341 17773
rect 32351 17759 32365 17773
rect 32375 17759 32389 17773
rect 32399 17759 32413 17773
rect 32423 17759 32437 17773
rect 32255 17567 32269 17581
rect 32279 17567 32293 17581
rect 32303 17567 32317 17581
rect 32327 17567 32341 17581
rect 32351 17567 32365 17581
rect 32375 17567 32389 17581
rect 32399 17567 32413 17581
rect 32423 17567 32437 17581
rect 32255 17519 32269 17533
rect 32279 17519 32293 17533
rect 32303 17519 32317 17533
rect 32327 17519 32341 17533
rect 32351 17519 32365 17533
rect 32375 17519 32389 17533
rect 32399 17519 32413 17533
rect 32423 17519 32437 17533
rect 32255 17327 32269 17341
rect 32279 17327 32293 17341
rect 32303 17327 32317 17341
rect 32327 17327 32341 17341
rect 32351 17327 32365 17341
rect 32375 17327 32389 17341
rect 32399 17327 32413 17341
rect 32423 17327 32437 17341
rect 32447 17327 32461 17341
rect 32255 17279 32269 17293
rect 32279 17279 32293 17293
rect 32303 17279 32317 17293
rect 32327 17279 32341 17293
rect 32351 17279 32365 17293
rect 32375 17279 32389 17293
rect 32399 17279 32413 17293
rect 32423 17279 32437 17293
rect 32447 17279 32461 17293
rect 32255 16847 32269 16861
rect 32279 16847 32293 16861
rect 32303 16847 32317 16861
rect 32327 16847 32341 16861
rect 32351 16847 32365 16861
rect 32375 16847 32389 16861
rect 32399 16847 32413 16861
rect 32423 16847 32437 16861
rect 32447 16847 32461 16861
rect 32471 16847 32485 16861
rect 32495 16847 32509 16861
rect 32255 16799 32269 16813
rect 32279 16799 32293 16813
rect 32303 16799 32317 16813
rect 32327 16799 32341 16813
rect 32351 16799 32365 16813
rect 32375 16799 32389 16813
rect 32399 16799 32413 16813
rect 32423 16799 32437 16813
rect 32447 16799 32461 16813
rect 32471 16799 32485 16813
rect 32495 16799 32509 16813
rect 32255 16607 32269 16621
rect 32279 16607 32293 16621
rect 32303 16607 32317 16621
rect 32327 16607 32341 16621
rect 32351 16607 32365 16621
rect 32375 16607 32389 16621
rect 32399 16607 32413 16621
rect 32423 16607 32437 16621
rect 32447 16607 32461 16621
rect 32471 16607 32485 16621
rect 32495 16607 32509 16621
rect 32519 16607 32533 16621
rect 32255 16559 32269 16573
rect 32279 16559 32293 16573
rect 32303 16559 32317 16573
rect 32327 16559 32341 16573
rect 32351 16559 32365 16573
rect 32375 16559 32389 16573
rect 32399 16559 32413 16573
rect 32423 16559 32437 16573
rect 32447 16559 32461 16573
rect 32471 16559 32485 16573
rect 32495 16559 32509 16573
rect 32519 16559 32533 16573
rect 32255 16367 32269 16381
rect 32279 16367 32293 16381
rect 32303 16367 32317 16381
rect 32327 16367 32341 16381
rect 32351 16367 32365 16381
rect 32375 16367 32389 16381
rect 32399 16367 32413 16381
rect 32423 16367 32437 16381
rect 32447 16367 32461 16381
rect 32471 16367 32485 16381
rect 32519 16391 32533 16405
rect 32543 16391 32557 16405
rect 32255 16319 32269 16333
rect 32279 16319 32293 16333
rect 32303 16319 32317 16333
rect 32327 16319 32341 16333
rect 32351 16319 32365 16333
rect 32375 16319 32389 16333
rect 32399 16319 32413 16333
rect 32423 16319 32437 16333
rect 32447 16319 32461 16333
rect 32471 16319 32485 16333
rect 32255 16127 32269 16141
rect 32279 16127 32293 16141
rect 32303 16127 32317 16141
rect 32327 16127 32341 16141
rect 32351 16127 32365 16141
rect 32519 16343 32533 16357
rect 32543 16343 32557 16357
rect 32399 16151 32413 16165
rect 32423 16151 32437 16165
rect 32447 16151 32461 16165
rect 32471 16151 32485 16165
rect 32495 16151 32509 16165
rect 32519 16151 32533 16165
rect 32543 16151 32557 16165
rect 32567 16151 32581 16165
rect 32255 16079 32269 16093
rect 32279 16079 32293 16093
rect 32303 16079 32317 16093
rect 32327 16079 32341 16093
rect 32351 16079 32365 16093
rect 32399 16103 32413 16117
rect 32423 16103 32437 16117
rect 32447 16103 32461 16117
rect 32471 16103 32485 16117
rect 32495 16103 32509 16117
rect 32519 16103 32533 16117
rect 32543 16103 32557 16117
rect 32567 16103 32581 16117
rect 32255 9863 32269 9877
rect 32279 9863 32293 9877
rect 32303 9863 32317 9877
rect 32327 9863 32341 9877
rect 32351 9863 32365 9877
rect 32375 9863 32389 9877
rect 32399 9863 32413 9877
rect 32423 9863 32437 9877
rect 32447 9863 32461 9877
rect 32471 9863 32485 9877
rect 32495 9863 32509 9877
rect 32543 9887 32557 9901
rect 32567 9887 32581 9901
rect 32591 9887 32605 9901
rect 32255 9815 32269 9829
rect 32279 9815 32293 9829
rect 32303 9815 32317 9829
rect 32327 9815 32341 9829
rect 32351 9815 32365 9829
rect 32375 9815 32389 9829
rect 32399 9815 32413 9829
rect 32423 9815 32437 9829
rect 32447 9815 32461 9829
rect 32471 9815 32485 9829
rect 32495 9815 32509 9829
rect 32255 9119 32269 9133
rect 32279 9119 32293 9133
rect 32303 9119 32317 9133
rect 32327 9119 32341 9133
rect 32351 9119 32365 9133
rect 32375 9119 32389 9133
rect 32399 9119 32413 9133
rect 32543 9839 32557 9853
rect 32567 9839 32581 9853
rect 32591 9839 32605 9853
rect 32447 9143 32461 9157
rect 32471 9143 32485 9157
rect 32495 9143 32509 9157
rect 32519 9143 32533 9157
rect 32543 9143 32557 9157
rect 32615 9191 32629 9205
rect 32255 9071 32269 9085
rect 32279 9071 32293 9085
rect 32303 9071 32317 9085
rect 32327 9071 32341 9085
rect 32351 9071 32365 9085
rect 32375 9071 32389 9085
rect 32399 9071 32413 9085
rect 32447 9095 32461 9109
rect 32471 9095 32485 9109
rect 32495 9095 32509 9109
rect 32519 9095 32533 9109
rect 32543 9095 32557 9109
rect 32615 9143 32629 9157
rect 32255 8687 32269 8701
rect 32279 8687 32293 8701
rect 32303 8687 32317 8701
rect 32327 8687 32341 8701
rect 32351 8687 32365 8701
rect 32375 8687 32389 8701
rect 32399 8687 32413 8701
rect 32423 8687 32437 8701
rect 32447 8687 32461 8701
rect 32471 8687 32485 8701
rect 32495 8687 32509 8701
rect 32519 8687 32533 8701
rect 32543 8687 32557 8701
rect 32567 8687 32581 8701
rect 32591 8687 32605 8701
rect 32615 8687 32629 8701
rect 32855 17207 32869 17221
rect 32855 17159 32869 17173
rect 32855 15527 32869 15541
rect 32903 15527 32917 15541
rect 32927 15527 32941 15541
rect 32951 15527 32965 15541
rect 32975 15527 32989 15541
rect 32999 15527 33013 15541
rect 33023 15527 33037 15541
rect 32855 15479 32869 15493
rect 32903 15479 32917 15493
rect 32927 15479 32941 15493
rect 32951 15479 32965 15493
rect 32975 15479 32989 15493
rect 32999 15479 33013 15493
rect 33023 15479 33037 15493
rect 32759 14327 32773 14341
rect 32855 14327 32869 14341
rect 32903 14327 32917 14341
rect 32927 14327 32941 14341
rect 32951 14327 32965 14341
rect 32975 14327 32989 14341
rect 32999 14327 33013 14341
rect 33023 14327 33037 14341
rect 33047 14327 33061 14341
rect 33071 14327 33085 14341
rect 33095 14327 33109 14341
rect 33119 14327 33133 14341
rect 32759 14279 32773 14293
rect 32855 14279 32869 14293
rect 32903 14279 32917 14293
rect 32927 14279 32941 14293
rect 32951 14279 32965 14293
rect 32975 14279 32989 14293
rect 32999 14279 33013 14293
rect 33023 14279 33037 14293
rect 33047 14279 33061 14293
rect 33071 14279 33085 14293
rect 33095 14279 33109 14293
rect 33119 14279 33133 14293
rect 32855 14087 32869 14101
rect 32903 14087 32917 14101
rect 32927 14087 32941 14101
rect 32951 14087 32965 14101
rect 32975 14087 32989 14101
rect 32999 14087 33013 14101
rect 33023 14087 33037 14101
rect 33047 14087 33061 14101
rect 33071 14087 33085 14101
rect 33095 14087 33109 14101
rect 33119 14087 33133 14101
rect 32855 14039 32869 14053
rect 32903 14039 32917 14053
rect 32927 14039 32941 14053
rect 32951 14039 32965 14053
rect 32975 14039 32989 14053
rect 32999 14039 33013 14053
rect 33023 14039 33037 14053
rect 33047 14039 33061 14053
rect 33071 14039 33085 14053
rect 33095 14039 33109 14053
rect 33119 14039 33133 14053
rect 32855 13607 32869 13621
rect 32903 13607 32917 13621
rect 32927 13607 32941 13621
rect 32951 13607 32965 13621
rect 32975 13607 32989 13621
rect 32999 13607 33013 13621
rect 33023 13607 33037 13621
rect 33047 13607 33061 13621
rect 33071 13607 33085 13621
rect 33095 13607 33109 13621
rect 33119 13607 33133 13621
rect 33143 13607 33157 13621
rect 32855 13559 32869 13573
rect 32903 13559 32917 13573
rect 32927 13559 32941 13573
rect 32951 13559 32965 13573
rect 32975 13559 32989 13573
rect 32999 13559 33013 13573
rect 33023 13559 33037 13573
rect 33047 13559 33061 13573
rect 33071 13559 33085 13573
rect 33095 13559 33109 13573
rect 33119 13559 33133 13573
rect 33143 13559 33157 13573
rect 41159 12887 41173 12901
rect 41159 12839 41173 12853
rect 41159 12647 41173 12661
rect 41159 12599 41173 12613
rect 41159 12407 41173 12421
rect 41159 12359 41173 12373
rect 32807 12167 32821 12181
rect 32831 12167 32845 12181
rect 32855 12167 32869 12181
rect 32903 12167 32917 12181
rect 32927 12167 32941 12181
rect 32951 12167 32965 12181
rect 32975 12167 32989 12181
rect 32999 12167 33013 12181
rect 33023 12167 33037 12181
rect 33047 12167 33061 12181
rect 33071 12167 33085 12181
rect 33095 12167 33109 12181
rect 33119 12167 33133 12181
rect 33143 12167 33157 12181
rect 33167 12167 33181 12181
rect 33191 12167 33205 12181
rect 33239 12167 33253 12181
rect 33263 12167 33277 12181
rect 41159 12167 41173 12181
rect 32807 12119 32821 12133
rect 32831 12119 32845 12133
rect 32855 12119 32869 12133
rect 32903 12119 32917 12133
rect 32927 12119 32941 12133
rect 32951 12119 32965 12133
rect 32975 12119 32989 12133
rect 32999 12119 33013 12133
rect 33023 12119 33037 12133
rect 33047 12119 33061 12133
rect 33071 12119 33085 12133
rect 33095 12119 33109 12133
rect 33119 12119 33133 12133
rect 33143 12119 33157 12133
rect 33167 12119 33181 12133
rect 33191 12119 33205 12133
rect 33239 12119 33253 12133
rect 33263 12119 33277 12133
rect 41159 12119 41173 12133
rect 32687 8735 32701 8749
rect 32711 8735 32725 8749
rect 32735 8735 32749 8749
rect 32759 8735 32773 8749
rect 32783 8735 32797 8749
rect 32807 8735 32821 8749
rect 32831 8735 32845 8749
rect 32855 8735 32869 8749
rect 32159 8615 32173 8629
rect 32687 8687 32701 8701
rect 32711 8687 32725 8701
rect 32735 8687 32749 8701
rect 32759 8687 32773 8701
rect 32783 8687 32797 8701
rect 32807 8687 32821 8701
rect 32831 8687 32845 8701
rect 32855 8687 32869 8701
rect 32663 8615 32677 8629
rect 32687 8615 32701 8629
rect 32711 8615 32725 8629
rect 32735 8615 32749 8629
rect 32759 8615 32773 8629
rect 32783 8615 32797 8629
rect 32807 8615 32821 8629
rect 32831 8615 32845 8629
rect 32855 8615 32869 8629
rect 32879 8615 32893 8629
rect 32903 8615 32917 8629
rect 32927 8615 32941 8629
rect 32951 8615 32965 8629
rect 32975 8615 32989 8629
rect 32999 8615 33013 8629
rect 33023 8615 33037 8629
rect 33047 8615 33061 8629
rect 33071 8615 33085 8629
rect 33095 8615 33109 8629
rect 33119 8615 33133 8629
rect 33143 8615 33157 8629
rect 32135 8591 32149 8605
rect 32111 8567 32125 8581
rect 32351 8567 32365 8581
rect 32615 8567 32629 8581
rect 32087 8543 32101 8557
rect 32063 8519 32077 8533
rect 32591 8519 32605 8533
rect 32615 8519 32629 8533
rect 32663 8567 32677 8581
rect 32687 8567 32701 8581
rect 33071 8567 33085 8581
rect 33095 8567 33109 8581
rect 33119 8567 33133 8581
rect 33143 8567 33157 8581
rect 41159 11927 41173 11941
rect 41159 11879 41173 11893
rect 41159 11687 41173 11701
rect 41159 11639 41173 11653
rect 33239 8807 33253 8821
rect 33263 8807 33277 8821
rect 33287 8807 33301 8821
rect 33311 8807 33325 8821
rect 41159 8807 41173 8821
rect 33239 8759 33253 8773
rect 33263 8759 33277 8773
rect 33287 8759 33301 8773
rect 33311 8759 33325 8773
rect 41159 8759 41173 8773
rect 32663 8519 32677 8533
rect 32687 8519 32701 8533
rect 32039 8495 32053 8509
rect 32927 8495 32941 8509
rect 33071 8495 33085 8509
rect 33215 8567 33229 8581
rect 33119 8495 33133 8509
rect 33143 8495 33157 8509
rect 33167 8495 33181 8509
rect 33191 8495 33205 8509
rect 33239 8495 33253 8509
rect 32015 8471 32029 8485
rect 31991 8447 32005 8461
rect 33239 8447 33253 8461
rect 31967 8423 31981 8437
rect 33023 8423 33037 8437
rect 31943 8399 31957 8413
rect 33119 8423 33133 8437
rect 33143 8423 33157 8437
rect 33167 8423 33181 8437
rect 33191 8423 33205 8437
rect 33215 8423 33229 8437
rect 31919 8375 31933 8389
rect 32567 8375 32581 8389
rect 32591 8375 32605 8389
rect 32615 8375 32629 8389
rect 32639 8375 32653 8389
rect 32663 8375 32677 8389
rect 32927 8375 32941 8389
rect 32951 8375 32965 8389
rect 33023 8375 33037 8389
rect 33047 8375 33061 8389
rect 33071 8375 33085 8389
rect 31895 8351 31909 8365
rect 31871 8327 31885 8341
rect 31847 8303 31861 8317
rect 32543 8303 32557 8317
rect 32567 8303 32581 8317
rect 32591 8303 32605 8317
rect 32615 8303 32629 8317
rect 32903 8303 32917 8317
rect 32927 8303 32941 8317
rect 32975 8303 32989 8317
rect 32999 8303 33013 8317
rect 33023 8303 33037 8317
rect 33215 8351 33229 8365
rect 32951 8279 32965 8293
rect 31823 8255 31837 8269
rect 32327 8255 32341 8269
rect 32519 8255 32533 8269
rect 32351 8231 32365 8245
rect 32495 8231 32509 8245
rect 32567 8255 32581 8269
rect 31799 8207 31813 8221
rect 32327 8207 32341 8221
rect 32567 8231 32581 8245
rect 32639 8255 32653 8269
rect 32663 8255 32677 8269
rect 32639 8231 32653 8245
rect 32519 8207 32533 8221
rect 32543 8207 32557 8221
rect 32855 8207 32869 8221
rect 32903 8207 32917 8221
rect 32951 8207 32965 8221
rect 33215 8303 33229 8317
rect 31799 8159 31813 8173
rect 31823 8159 31837 8173
rect 31847 8159 31861 8173
rect 31871 8159 31885 8173
rect 31895 8159 31909 8173
rect 31919 8159 31933 8173
rect 31943 8159 31957 8173
rect 31967 8159 31981 8173
rect 31991 8159 32005 8173
rect 32015 8159 32029 8173
rect 32039 8159 32053 8173
rect 32063 8159 32077 8173
rect 32087 8159 32101 8173
rect 32111 8159 32125 8173
rect 32135 8159 32149 8173
rect 32159 8159 32173 8173
rect 32255 8159 32269 8173
rect 32279 8159 32293 8173
rect 32303 8159 32317 8173
rect 32327 8159 32341 8173
rect 32351 8159 32365 8173
rect 32375 8159 32389 8173
rect 32399 8159 32413 8173
rect 32423 8159 32437 8173
rect 32447 8159 32461 8173
rect 32471 8159 32485 8173
rect 32519 8159 32533 8173
rect 32543 8159 32557 8173
rect 32567 8159 32581 8173
rect 32903 8159 32917 8173
rect 32615 8135 32629 8149
rect 32639 8135 32653 8149
rect 32663 8135 32677 8149
rect 32687 8135 32701 8149
rect 32711 8135 32725 8149
rect 32735 8135 32749 8149
rect 32759 8135 32773 8149
rect 32783 8135 32797 8149
rect 32807 8135 32821 8149
rect 32831 8135 32845 8149
rect 32879 8111 32893 8125
rect 31775 6407 31789 6421
rect 31799 6407 31813 6421
rect 31823 6407 31837 6421
rect 31847 6407 31861 6421
rect 31871 6407 31885 6421
rect 31895 6407 31909 6421
rect 31919 6407 31933 6421
rect 31943 6407 31957 6421
rect 31967 6407 31981 6421
rect 31991 6407 32005 6421
rect 32015 6407 32029 6421
rect 32039 6407 32053 6421
rect 32063 6407 32077 6421
rect 32087 6407 32101 6421
rect 32111 6407 32125 6421
rect 32135 6407 32149 6421
rect 32159 6407 32173 6421
rect 32255 6407 32269 6421
rect 32279 6407 32293 6421
rect 32303 6407 32317 6421
rect 32327 6407 32341 6421
rect 32351 6407 32365 6421
rect 32375 6407 32389 6421
rect 32399 6407 32413 6421
rect 32423 6407 32437 6421
rect 32447 6407 32461 6421
rect 32471 6407 32485 6421
rect 32519 6407 32533 6421
rect 32543 6407 32557 6421
rect 32567 6407 32581 6421
rect 32591 6407 32605 6421
rect 32615 6407 32629 6421
rect 32639 6407 32653 6421
rect 32663 6407 32677 6421
rect 32687 6407 32701 6421
rect 32711 6407 32725 6421
rect 32735 6407 32749 6421
rect 32759 6407 32773 6421
rect 32783 6407 32797 6421
rect 32807 6407 32821 6421
rect 32831 6407 32845 6421
rect 32855 6407 32869 6421
rect 32879 6407 32893 6421
rect 32903 6407 32917 6421
rect 33215 6407 33229 6421
rect 41159 6407 41173 6421
rect 31775 6359 31789 6373
rect 31799 6359 31813 6373
rect 31823 6359 31837 6373
rect 31847 6359 31861 6373
rect 31871 6359 31885 6373
rect 31895 6359 31909 6373
rect 31919 6359 31933 6373
rect 31943 6359 31957 6373
rect 31967 6359 31981 6373
rect 31991 6359 32005 6373
rect 32015 6359 32029 6373
rect 32039 6359 32053 6373
rect 32063 6359 32077 6373
rect 32087 6359 32101 6373
rect 32111 6359 32125 6373
rect 32135 6359 32149 6373
rect 32159 6359 32173 6373
rect 32255 6359 32269 6373
rect 32279 6359 32293 6373
rect 32303 6359 32317 6373
rect 32327 6359 32341 6373
rect 32351 6359 32365 6373
rect 32375 6359 32389 6373
rect 32399 6359 32413 6373
rect 32423 6359 32437 6373
rect 32447 6359 32461 6373
rect 32471 6359 32485 6373
rect 32519 6359 32533 6373
rect 32543 6359 32557 6373
rect 32567 6359 32581 6373
rect 32591 6359 32605 6373
rect 32615 6359 32629 6373
rect 32639 6359 32653 6373
rect 32663 6359 32677 6373
rect 32687 6359 32701 6373
rect 32711 6359 32725 6373
rect 32735 6359 32749 6373
rect 32759 6359 32773 6373
rect 32783 6359 32797 6373
rect 32807 6359 32821 6373
rect 32831 6359 32845 6373
rect 32855 6359 32869 6373
rect 32879 6359 32893 6373
rect 32903 6359 32917 6373
rect 33215 6359 33229 6373
rect 41159 6359 41173 6373
rect 31751 6167 31765 6181
rect 31775 6167 31789 6181
rect 31799 6167 31813 6181
rect 31823 6167 31837 6181
rect 31847 6167 31861 6181
rect 31871 6167 31885 6181
rect 31895 6167 31909 6181
rect 31919 6167 31933 6181
rect 31943 6167 31957 6181
rect 31967 6167 31981 6181
rect 31991 6167 32005 6181
rect 32015 6167 32029 6181
rect 32039 6167 32053 6181
rect 32063 6167 32077 6181
rect 32087 6167 32101 6181
rect 32111 6167 32125 6181
rect 32135 6167 32149 6181
rect 32159 6167 32173 6181
rect 32255 6167 32269 6181
rect 32279 6167 32293 6181
rect 32303 6167 32317 6181
rect 32327 6167 32341 6181
rect 32351 6167 32365 6181
rect 32375 6167 32389 6181
rect 32399 6167 32413 6181
rect 32423 6167 32437 6181
rect 32447 6167 32461 6181
rect 32471 6167 32485 6181
rect 32519 6167 32533 6181
rect 32543 6167 32557 6181
rect 32567 6167 32581 6181
rect 32591 6167 32605 6181
rect 32615 6167 32629 6181
rect 32639 6167 32653 6181
rect 32663 6167 32677 6181
rect 32687 6167 32701 6181
rect 32711 6167 32725 6181
rect 32735 6167 32749 6181
rect 32759 6167 32773 6181
rect 32783 6167 32797 6181
rect 32807 6167 32821 6181
rect 32831 6167 32845 6181
rect 32855 6167 32869 6181
rect 32879 6167 32893 6181
rect 32903 6167 32917 6181
rect 33215 6167 33229 6181
rect 41159 6167 41173 6181
rect 31751 6119 31765 6133
rect 31775 6119 31789 6133
rect 31799 6119 31813 6133
rect 31823 6119 31837 6133
rect 31847 6119 31861 6133
rect 31871 6119 31885 6133
rect 31895 6119 31909 6133
rect 31919 6119 31933 6133
rect 31943 6119 31957 6133
rect 31967 6119 31981 6133
rect 31991 6119 32005 6133
rect 32015 6119 32029 6133
rect 32039 6119 32053 6133
rect 32063 6119 32077 6133
rect 32087 6119 32101 6133
rect 32111 6119 32125 6133
rect 32135 6119 32149 6133
rect 32159 6119 32173 6133
rect 32255 6119 32269 6133
rect 32279 6119 32293 6133
rect 32303 6119 32317 6133
rect 32327 6119 32341 6133
rect 32351 6119 32365 6133
rect 32375 6119 32389 6133
rect 32399 6119 32413 6133
rect 32423 6119 32437 6133
rect 32447 6119 32461 6133
rect 32471 6119 32485 6133
rect 32519 6119 32533 6133
rect 32543 6119 32557 6133
rect 32567 6119 32581 6133
rect 32591 6119 32605 6133
rect 32615 6119 32629 6133
rect 32639 6119 32653 6133
rect 32663 6119 32677 6133
rect 32687 6119 32701 6133
rect 32711 6119 32725 6133
rect 32735 6119 32749 6133
rect 32759 6119 32773 6133
rect 32783 6119 32797 6133
rect 32807 6119 32821 6133
rect 32831 6119 32845 6133
rect 32855 6119 32869 6133
rect 32879 6119 32893 6133
rect 32903 6119 32917 6133
rect 33215 6119 33229 6133
rect 41159 6119 41173 6133
rect 41159 5927 41173 5941
rect 41159 5879 41173 5893
rect 41159 5687 41173 5701
rect 41159 5639 41173 5653
rect 31727 5447 31741 5461
rect 31751 5447 31765 5461
rect 31775 5447 31789 5461
rect 31799 5447 31813 5461
rect 31823 5447 31837 5461
rect 31847 5447 31861 5461
rect 31871 5447 31885 5461
rect 31895 5447 31909 5461
rect 31919 5447 31933 5461
rect 31943 5447 31957 5461
rect 31967 5447 31981 5461
rect 31991 5447 32005 5461
rect 32015 5447 32029 5461
rect 32039 5447 32053 5461
rect 32063 5447 32077 5461
rect 32087 5447 32101 5461
rect 32111 5447 32125 5461
rect 32135 5447 32149 5461
rect 32159 5447 32173 5461
rect 32255 5447 32269 5461
rect 32279 5447 32293 5461
rect 32303 5447 32317 5461
rect 32327 5447 32341 5461
rect 32351 5447 32365 5461
rect 32375 5447 32389 5461
rect 32399 5447 32413 5461
rect 32423 5447 32437 5461
rect 32447 5447 32461 5461
rect 32471 5447 32485 5461
rect 32519 5447 32533 5461
rect 32543 5447 32557 5461
rect 32567 5447 32581 5461
rect 32591 5447 32605 5461
rect 32615 5447 32629 5461
rect 32639 5447 32653 5461
rect 32663 5447 32677 5461
rect 32687 5447 32701 5461
rect 32711 5447 32725 5461
rect 32735 5447 32749 5461
rect 32759 5447 32773 5461
rect 32783 5447 32797 5461
rect 32807 5447 32821 5461
rect 32831 5447 32845 5461
rect 32855 5447 32869 5461
rect 32879 5447 32893 5461
rect 32903 5447 32917 5461
rect 33215 5447 33229 5461
rect 33335 5447 33349 5461
rect 33383 5447 33397 5461
rect 41159 5447 41173 5461
rect 27599 5399 27613 5413
rect 27647 5399 27661 5413
rect 27863 5399 27877 5413
rect 27935 5399 27949 5413
rect 27959 5399 27973 5413
rect 28031 5399 28045 5413
rect 28079 5399 28093 5413
rect 28127 5399 28141 5413
rect 27551 5375 27565 5389
rect 27743 5375 27757 5389
rect 27791 5375 27805 5389
rect 28247 5375 28261 5389
rect 27527 5351 27541 5365
rect 28343 5351 28357 5365
rect 28391 5351 28405 5365
rect 28439 5351 28453 5365
rect 26975 5327 26989 5341
rect 27071 5327 27085 5341
rect 27239 5327 27253 5341
rect 27287 5327 27301 5341
rect 27311 5327 27325 5341
rect 27407 5327 27421 5341
rect 27455 5327 27469 5341
rect 28535 5327 28549 5341
rect 28583 5327 28597 5341
rect 28631 5327 28645 5341
rect 28679 5327 28693 5341
rect 28727 5327 28741 5341
rect 28751 5327 28765 5341
rect 28823 5327 28837 5341
rect 30455 5327 30469 5341
rect 30527 5327 30541 5341
rect 26855 5303 26869 5317
rect 27191 5303 27205 5317
rect 27215 5303 27229 5317
rect 28919 5303 28933 5317
rect 30239 5303 30253 5317
rect 30287 5303 30301 5317
rect 30311 5303 30325 5317
rect 30383 5303 30397 5317
rect 30431 5303 30445 5317
rect 30647 5303 30661 5317
rect 30671 5303 30685 5317
rect 30767 5303 30781 5317
rect 24551 5279 24565 5293
rect 24599 5279 24613 5293
rect 26447 5279 26461 5293
rect 26495 5279 26509 5293
rect 26783 5279 26797 5293
rect 29015 5279 29029 5293
rect 29999 5279 30013 5293
rect 30071 5279 30085 5293
rect 30095 5279 30109 5293
rect 30167 5279 30181 5293
rect 30215 5279 30229 5293
rect 30887 5279 30901 5293
rect 30935 5279 30949 5293
rect 31007 5279 31021 5293
rect 31439 5279 31453 5293
rect 31487 5279 31501 5293
rect 31511 5279 31525 5293
rect 31583 5279 31597 5293
rect 24527 5255 24541 5269
rect 24695 5255 24709 5269
rect 26399 5255 26413 5269
rect 26591 5255 26605 5269
rect 26639 5255 26653 5269
rect 26711 5255 26725 5269
rect 26735 5255 26749 5269
rect 29111 5255 29125 5269
rect 29975 5255 29989 5269
rect 31127 5255 31141 5269
rect 31151 5255 31165 5269
rect 31247 5255 31261 5269
rect 31391 5255 31405 5269
rect 31727 5399 31741 5413
rect 31751 5399 31765 5413
rect 31775 5399 31789 5413
rect 31799 5399 31813 5413
rect 31823 5399 31837 5413
rect 31847 5399 31861 5413
rect 31871 5399 31885 5413
rect 31895 5399 31909 5413
rect 31919 5399 31933 5413
rect 31943 5399 31957 5413
rect 31967 5399 31981 5413
rect 31991 5399 32005 5413
rect 32015 5399 32029 5413
rect 32039 5399 32053 5413
rect 32063 5399 32077 5413
rect 32087 5399 32101 5413
rect 32111 5399 32125 5413
rect 32135 5399 32149 5413
rect 32159 5399 32173 5413
rect 32255 5399 32269 5413
rect 32279 5399 32293 5413
rect 32303 5399 32317 5413
rect 32327 5399 32341 5413
rect 32351 5399 32365 5413
rect 32375 5399 32389 5413
rect 32399 5399 32413 5413
rect 32423 5399 32437 5413
rect 32447 5399 32461 5413
rect 32471 5399 32485 5413
rect 32519 5399 32533 5413
rect 32543 5399 32557 5413
rect 32567 5399 32581 5413
rect 32591 5399 32605 5413
rect 32615 5399 32629 5413
rect 32639 5399 32653 5413
rect 32663 5399 32677 5413
rect 32687 5399 32701 5413
rect 32711 5399 32725 5413
rect 32735 5399 32749 5413
rect 32759 5399 32773 5413
rect 32783 5399 32797 5413
rect 32807 5399 32821 5413
rect 32831 5399 32845 5413
rect 32855 5399 32869 5413
rect 32879 5399 32893 5413
rect 32903 5399 32917 5413
rect 33215 5399 33229 5413
rect 33335 5399 33349 5413
rect 33383 5399 33397 5413
rect 41159 5399 41173 5413
rect 24503 5231 24517 5245
rect 24815 5231 24829 5245
rect 24839 5231 24853 5245
rect 24935 5231 24949 5245
rect 24959 5231 24973 5245
rect 25031 5231 25045 5245
rect 26375 5231 26389 5245
rect 29231 5231 29245 5245
rect 29255 5231 29269 5245
rect 29327 5231 29341 5245
rect 29423 5231 29437 5245
rect 31703 5231 31717 5245
rect 31727 5231 31741 5245
rect 31751 5231 31765 5245
rect 24383 5207 24397 5221
rect 24455 5207 24469 5221
rect 24479 5207 24493 5221
rect 25127 5207 25141 5221
rect 25175 5207 25189 5221
rect 25223 5207 25237 5221
rect 25247 5207 25261 5221
rect 25343 5207 25357 5221
rect 25367 5207 25381 5221
rect 25439 5207 25453 5221
rect 25463 5207 25477 5221
rect 25535 5207 25549 5221
rect 25631 5207 25645 5221
rect 26255 5207 26269 5221
rect 26303 5207 26317 5221
rect 24263 5183 24277 5197
rect 24335 5183 24349 5197
rect 24359 5183 24373 5197
rect 31823 5183 31837 5197
rect 24239 5159 24253 5173
rect 24023 5135 24037 5149
rect 24095 5135 24109 5149
rect 24119 5135 24133 5149
rect 23903 5111 23917 5125
rect 23975 5111 23989 5125
rect 23999 5111 24013 5125
rect 23687 5087 23701 5101
rect 23735 5087 23749 5101
rect 23807 5087 23821 5101
rect 23855 5087 23869 5101
rect 23879 5087 23893 5101
rect 31895 5087 31909 5101
rect 31919 5087 31933 5101
rect 31943 5087 31957 5101
rect 31967 5087 31981 5101
rect 23543 5063 23557 5077
rect 23615 5063 23629 5077
rect 23639 5063 23653 5077
rect 23519 5039 23533 5053
rect 23399 5015 23413 5029
rect 29423 5015 29437 5029
rect 29447 5015 29461 5029
rect 32015 5015 32029 5029
rect 23303 4991 23317 5005
rect 32063 4991 32077 5005
rect 23279 4967 23293 4981
rect 32111 4967 32125 4981
rect 32135 4967 32149 4981
rect 32159 4967 32173 4981
rect 32255 4967 32269 4981
rect 32279 4967 32293 4981
rect 32303 4967 32317 4981
rect 32327 4967 32341 4981
rect 32351 4967 32365 4981
rect 32375 4967 32389 4981
rect 32399 4967 32413 4981
rect 32423 4967 32437 4981
rect 32447 4967 32461 4981
rect 32471 4967 32485 4981
rect 23255 4943 23269 4957
rect 28391 4943 28405 4957
rect 28415 4943 28429 4957
rect 23159 4919 23173 4933
rect 32111 4919 32125 4933
rect 32255 4919 32269 4933
rect 32279 4919 32293 4933
rect 32303 4919 32317 4933
rect 32327 4919 32341 4933
rect 32351 4919 32365 4933
rect 32375 4919 32389 4933
rect 32399 4919 32413 4933
rect 32423 4919 32437 4933
rect 32447 4919 32461 4933
rect 32471 4919 32485 4933
rect 23135 4895 23149 4909
rect 27791 4895 27805 4909
rect 27815 4895 27829 4909
rect 23015 4871 23029 4885
rect 23087 4871 23101 4885
rect 23111 4871 23125 4885
rect 32111 4871 32125 4885
rect 22799 4847 22813 4861
rect 22895 4847 22909 4861
rect 22943 4847 22957 4861
rect 24959 4847 24973 4861
rect 24983 4847 24997 4861
rect 25295 4847 25309 4861
rect 26567 4847 26581 4861
rect 27119 4847 27133 4861
rect 30935 4847 30949 4861
rect 30959 4847 30973 4861
rect 31223 4847 31237 4861
rect 31679 4847 31693 4861
rect 32255 4871 32269 4885
rect 32279 4871 32293 4885
rect 32303 4871 32317 4885
rect 32327 4871 32341 4885
rect 32351 4871 32365 4885
rect 32375 4871 32389 4885
rect 32399 4871 32413 4885
rect 32423 4871 32437 4885
rect 32447 4871 32461 4885
rect 32471 4871 32485 4885
rect 32495 4871 32509 4885
rect 32519 4871 32533 4885
rect 32543 4871 32557 4885
rect 32567 4871 32581 4885
rect 32591 4871 32605 4885
rect 32615 4871 32629 4885
rect 32639 4871 32653 4885
rect 32663 4871 32677 4885
rect 32687 4871 32701 4885
rect 32711 4871 32725 4885
rect 32735 4871 32749 4885
rect 32759 4871 32773 4885
rect 32783 4871 32797 4885
rect 32807 4871 32821 4885
rect 32831 4871 32845 4885
rect 32855 4871 32869 4885
rect 32903 4895 32917 4909
rect 32927 4871 32941 4885
rect 32951 4847 32965 4861
rect 22775 4823 22789 4837
rect 32159 4823 32173 4837
rect 32183 4823 32197 4837
rect 32231 4823 32245 4837
rect 32495 4823 32509 4837
rect 32975 4823 32989 4837
rect 22415 4799 22429 4813
rect 22535 4799 22549 4813
rect 22559 4799 22573 4813
rect 22631 4799 22645 4813
rect 22679 4799 22693 4813
rect 29255 4799 29269 4813
rect 29279 4799 29293 4813
rect 22343 4775 22357 4789
rect 32879 4775 32893 4789
rect 32999 4775 33013 4789
rect 22247 4751 22261 4765
rect 22295 4751 22309 4765
rect 22319 4751 22333 4765
rect 22991 4751 23005 4765
rect 23039 4751 23053 4765
rect 26735 4751 26749 4765
rect 26759 4751 26773 4765
rect 33023 4751 33037 4765
rect 59759 4967 59773 4981
rect 59759 4919 59773 4933
rect 22199 4727 22213 4741
rect 23783 4727 23797 4741
rect 32207 4727 32221 4741
rect 33047 4727 33061 4741
rect 33215 4727 33229 4741
rect 33335 4727 33349 4741
rect 33383 4727 33397 4741
rect 41159 4727 41173 4741
rect 59039 4727 59053 4741
rect 59759 4727 59773 4741
rect 21623 4703 21637 4717
rect 21671 4703 21685 4717
rect 21719 4703 21733 4717
rect 21791 4703 21805 4717
rect 21839 4703 21853 4717
rect 21911 4703 21925 4717
rect 21935 4703 21949 4717
rect 22031 4703 22045 4717
rect 22055 4703 22069 4717
rect 22127 4703 22141 4717
rect 22175 4703 22189 4717
rect 32495 4703 32509 4717
rect 32879 4703 32893 4717
rect 21575 4679 21589 4693
rect 32063 4679 32077 4693
rect 32087 4679 32101 4693
rect 32207 4679 32221 4693
rect 32879 4679 32893 4693
rect 33215 4679 33229 4693
rect 33335 4679 33349 4693
rect 33383 4679 33397 4693
rect 41159 4679 41173 4693
rect 59039 4679 59053 4693
rect 59759 4679 59773 4693
rect 21071 4655 21085 4669
rect 21143 4655 21157 4669
rect 21551 4655 21565 4669
rect 32207 4655 32221 4669
rect 33071 4655 33085 4669
rect 20447 4631 20461 4645
rect 20543 4631 20557 4645
rect 20567 4631 20581 4645
rect 20639 4631 20653 4645
rect 20711 4631 20725 4645
rect 20759 4631 20773 4645
rect 20807 4631 20821 4645
rect 20855 4631 20869 4645
rect 20975 4631 20989 4645
rect 21239 4631 21253 4645
rect 21263 4631 21277 4645
rect 21335 4631 21349 4645
rect 21479 4631 21493 4645
rect 32375 4631 32389 4645
rect 32495 4631 32509 4645
rect 33095 4631 33109 4645
rect 20423 4607 20437 4621
rect 21431 4607 21445 4621
rect 21455 4607 21469 4621
rect 23159 4607 23173 4621
rect 23183 4607 23197 4621
rect 31151 4607 31165 4621
rect 31175 4607 31189 4621
rect 32207 4607 32221 4621
rect 33119 4607 33133 4621
rect 20351 4583 20365 4597
rect 33143 4583 33157 4597
rect 20327 4559 20341 4573
rect 27503 4559 27517 4573
rect 27575 4559 27589 4573
rect 32207 4559 32221 4573
rect 20207 4535 20221 4549
rect 32351 4535 32365 4549
rect 32375 4535 32389 4549
rect 32543 4535 32557 4549
rect 19391 4511 19405 4525
rect 19463 4511 19477 4525
rect 19487 4511 19501 4525
rect 19559 4511 19573 4525
rect 19607 4511 19621 4525
rect 19703 4511 19717 4525
rect 19799 4511 19813 4525
rect 26951 4511 26965 4525
rect 26999 4511 27013 4525
rect 27719 4511 27733 4525
rect 32207 4511 32221 4525
rect 32543 4511 32557 4525
rect 33167 4511 33181 4525
rect 19271 4487 19285 4501
rect 19343 4487 19357 4501
rect 19367 4487 19381 4501
rect 19151 4463 19165 4477
rect 19223 4463 19237 4477
rect 19247 4463 19261 4477
rect 32759 4463 32773 4477
rect 33191 4463 33205 4477
rect 19079 4439 19093 4453
rect 19055 4415 19069 4429
rect 32375 4415 32389 4429
rect 32495 4415 32509 4429
rect 32807 4415 32821 4429
rect 32951 4415 32965 4429
rect 33215 4415 33229 4429
rect 18935 4391 18949 4405
rect 20423 4391 20437 4405
rect 20471 4391 20485 4405
rect 31175 4391 31189 4405
rect 31199 4391 31213 4405
rect 31655 4391 31669 4405
rect 32207 4391 32221 4405
rect 32951 4391 32965 4405
rect 33023 4391 33037 4405
rect 33239 4391 33253 4405
rect 18767 4367 18781 4381
rect 18815 4367 18829 4381
rect 18863 4367 18877 4381
rect 24023 4367 24037 4381
rect 24047 4367 24061 4381
rect 33263 4367 33277 4381
rect 18623 4343 18637 4357
rect 18719 4343 18733 4357
rect 18743 4343 18757 4357
rect 32183 4343 32197 4357
rect 32207 4343 32221 4357
rect 33287 4343 33301 4357
rect 18551 4319 18565 4333
rect 18455 4295 18469 4309
rect 18503 4295 18517 4309
rect 18527 4295 18541 4309
rect 33023 4295 33037 4309
rect 33311 4295 33325 4309
rect 33335 4295 33349 4309
rect 41159 4487 41173 4501
rect 59039 4487 59053 4501
rect 59759 4487 59773 4501
rect 18431 4271 18445 4285
rect 32495 4271 32509 4285
rect 32543 4271 32557 4285
rect 33359 4271 33373 4285
rect 33383 4271 33397 4285
rect 41159 4439 41173 4453
rect 59039 4439 59053 4453
rect 59759 4439 59773 4453
rect 18335 4247 18349 4261
rect 18383 4247 18397 4261
rect 18407 4247 18421 4261
rect 32207 4247 32221 4261
rect 32231 4247 32245 4261
rect 33407 4247 33421 4261
rect 33479 4247 33493 4261
rect 41159 4247 41173 4261
rect 59039 4247 59053 4261
rect 59759 4247 59773 4261
rect 18287 4223 18301 4237
rect 18263 4199 18277 4213
rect 27599 4199 27613 4213
rect 27623 4199 27637 4213
rect 32207 4199 32221 4213
rect 33431 4199 33445 4213
rect 33455 4199 33469 4213
rect 33503 4199 33517 4213
rect 41159 4199 41173 4213
rect 59039 4199 59053 4213
rect 59759 4199 59773 4213
rect 17351 4175 17365 4189
rect 17447 4175 17461 4189
rect 17567 4175 17581 4189
rect 33527 4175 33541 4189
rect 33551 4175 33565 4189
rect 33599 4175 33613 4189
rect 35399 4175 35413 4189
rect 35447 4175 35461 4189
rect 17135 4151 17149 4165
rect 33695 4151 33709 4165
rect 35375 4151 35389 4165
rect 35567 4151 35581 4165
rect 16919 4127 16933 4141
rect 17087 4127 17101 4141
rect 17303 4127 17317 4141
rect 17519 4127 17533 4141
rect 17735 4127 17749 4141
rect 17951 4127 17965 4141
rect 18167 4127 18181 4141
rect 22055 4127 22069 4141
rect 22079 4127 22093 4141
rect 23903 4127 23917 4141
rect 23927 4127 23941 4141
rect 24047 4127 24061 4141
rect 24071 4127 24085 4141
rect 27383 4127 27397 4141
rect 32207 4127 32221 4141
rect 33815 4127 33829 4141
rect 35255 4127 35269 4141
rect 35327 4127 35341 4141
rect 35351 4127 35365 4141
rect 35663 4127 35677 4141
rect 16703 4103 16717 4117
rect 32231 4103 32245 4117
rect 33935 4103 33949 4117
rect 33959 4103 33973 4117
rect 34031 4103 34045 4117
rect 34055 4103 34069 4117
rect 34127 4103 34141 4117
rect 34151 4103 34165 4117
rect 34223 4103 34237 4117
rect 35135 4103 35149 4117
rect 35207 4103 35221 4117
rect 35231 4103 35245 4117
rect 35759 4103 35773 4117
rect 16487 4079 16501 4093
rect 22751 4079 22765 4093
rect 22823 4079 22837 4093
rect 32183 4079 32197 4093
rect 32207 4079 32221 4093
rect 34343 4079 34357 4093
rect 34847 4079 34861 4093
rect 34895 4079 34909 4093
rect 34919 4079 34933 4093
rect 34991 4079 35005 4093
rect 35015 4079 35029 4093
rect 35087 4079 35101 4093
rect 35111 4079 35125 4093
rect 35855 4079 35869 4093
rect 16271 4055 16285 4069
rect 33479 4055 33493 4069
rect 33527 4055 33541 4069
rect 34439 4055 34453 4069
rect 34463 4055 34477 4069
rect 34535 4055 34549 4069
rect 34727 4055 34741 4069
rect 34799 4055 34813 4069
rect 34823 4055 34837 4069
rect 35951 4055 35965 4069
rect 35975 4055 35989 4069
rect 36047 4055 36061 4069
rect 16055 4031 16069 4045
rect 21575 4031 21589 4045
rect 21599 4031 21613 4045
rect 32543 4031 32557 4045
rect 32759 4031 32773 4045
rect 32831 4031 32845 4045
rect 33263 4031 33277 4045
rect 34199 4031 34213 4045
rect 34223 4031 34237 4045
rect 34631 4031 34645 4045
rect 34679 4031 34693 4045
rect 34943 4031 34957 4045
rect 36143 4031 36157 4045
rect 15839 4007 15853 4021
rect 32135 4007 32149 4021
rect 32159 4007 32173 4021
rect 34775 4007 34789 4021
rect 34799 4007 34813 4021
rect 36263 4007 36277 4021
rect 36287 4007 36301 4021
rect 36359 4007 36373 4021
rect 41159 4007 41173 4021
rect 59039 4007 59053 4021
rect 59759 4007 59773 4021
rect 15383 3983 15397 3997
rect 15455 3983 15469 3997
rect 15623 3983 15637 3997
rect 23231 3983 23245 3997
rect 23327 3983 23341 3997
rect 32495 3983 32509 3997
rect 33263 3983 33277 3997
rect 15359 3959 15373 3973
rect 32327 3959 32341 3973
rect 32351 3959 32365 3973
rect 36455 3959 36469 3973
rect 41159 3959 41173 3973
rect 59039 3959 59053 3973
rect 59759 3959 59773 3973
rect 15071 3935 15085 3949
rect 15119 3935 15133 3949
rect 15311 3935 15325 3949
rect 32663 3935 32677 3949
rect 32807 3935 32821 3949
rect 32855 3935 32869 3949
rect 33215 3935 33229 3949
rect 33239 3935 33253 3949
rect 36551 3935 36565 3949
rect 15023 3911 15037 3925
rect 32303 3911 32317 3925
rect 32327 3911 32341 3925
rect 32855 3911 32869 3925
rect 36671 3911 36685 3925
rect 14663 3887 14677 3901
rect 14711 3887 14725 3901
rect 14735 3887 14749 3901
rect 14807 3887 14821 3901
rect 14831 3887 14845 3901
rect 14903 3887 14917 3901
rect 14927 3887 14941 3901
rect 32207 3887 32221 3901
rect 36791 3887 36805 3901
rect 14567 3863 14581 3877
rect 14615 3863 14629 3877
rect 14639 3863 14653 3877
rect 19607 3863 19621 3877
rect 19631 3863 19645 3877
rect 36887 3863 36901 3877
rect 36911 3863 36925 3877
rect 37031 3863 37045 3877
rect 37055 3863 37069 3877
rect 37127 3863 37141 3877
rect 37151 3863 37165 3877
rect 37223 3863 37237 3877
rect 14471 3839 14485 3853
rect 14519 3839 14533 3853
rect 14543 3839 14557 3853
rect 17807 3839 17821 3853
rect 23303 3839 23317 3853
rect 23351 3839 23365 3853
rect 37343 3839 37357 3853
rect 37391 3839 37405 3853
rect 37463 3839 37477 3853
rect 37487 3839 37501 3853
rect 37583 3839 37597 3853
rect 14255 3815 14269 3829
rect 14327 3815 14341 3829
rect 14375 3815 14389 3829
rect 14423 3815 14437 3829
rect 14447 3815 14461 3829
rect 14831 3815 14845 3829
rect 14855 3815 14869 3829
rect 21839 3815 21853 3829
rect 21863 3815 21877 3829
rect 37679 3815 37693 3829
rect 37727 3815 37741 3829
rect 37775 3815 37789 3829
rect 14231 3791 14245 3805
rect 32759 3791 32773 3805
rect 32831 3791 32845 3805
rect 32903 3791 32917 3805
rect 33167 3791 33181 3805
rect 33191 3791 33205 3805
rect 37871 3791 37885 3805
rect 14159 3767 14173 3781
rect 19031 3767 19045 3781
rect 19103 3767 19117 3781
rect 23255 3767 23269 3781
rect 23303 3767 23317 3781
rect 32207 3767 32221 3781
rect 32903 3767 32917 3781
rect 35807 3767 35821 3781
rect 37511 3767 37525 3781
rect 37967 3767 37981 3781
rect 14015 3743 14029 3757
rect 18455 3743 18469 3757
rect 18479 3743 18493 3757
rect 28679 3743 28693 3757
rect 28703 3743 28717 3757
rect 38087 3743 38101 3757
rect 38111 3743 38125 3757
rect 38183 3743 38197 3757
rect 13583 3719 13597 3733
rect 13655 3719 13669 3733
rect 13679 3719 13693 3733
rect 13751 3719 13765 3733
rect 13871 3719 13885 3733
rect 14159 3719 14173 3733
rect 14183 3719 14197 3733
rect 32687 3719 32701 3733
rect 32759 3719 32773 3733
rect 32807 3719 32821 3733
rect 33119 3719 33133 3733
rect 38303 3719 38317 3733
rect 13487 3695 13501 3709
rect 13535 3695 13549 3709
rect 13559 3695 13573 3709
rect 30455 3695 30469 3709
rect 30479 3695 30493 3709
rect 32207 3695 32221 3709
rect 35183 3695 35197 3709
rect 35207 3695 35221 3709
rect 38423 3695 38437 3709
rect 13463 3671 13477 3685
rect 38519 3671 38533 3685
rect 13439 3647 13453 3661
rect 19391 3647 19405 3661
rect 19415 3647 19429 3661
rect 26639 3647 26653 3661
rect 26663 3647 26677 3661
rect 32207 3647 32221 3661
rect 38663 3647 38677 3661
rect 13391 3623 13405 3637
rect 25175 3623 25189 3637
rect 25199 3623 25213 3637
rect 25511 3623 25525 3637
rect 26231 3623 26245 3637
rect 31367 3623 31381 3637
rect 31415 3623 31429 3637
rect 38759 3623 38773 3637
rect 38903 3623 38917 3637
rect 38951 3623 38965 3637
rect 39695 3623 39709 3637
rect 39767 3623 39781 3637
rect 39791 3623 39805 3637
rect 39863 3623 39877 3637
rect 39887 3623 39901 3637
rect 39959 3623 39973 3637
rect 40487 3623 40501 3637
rect 40559 3623 40573 3637
rect 40583 3623 40597 3637
rect 40655 3623 40669 3637
rect 13367 3599 13381 3613
rect 20327 3599 20341 3613
rect 20375 3599 20389 3613
rect 25631 3599 25645 3613
rect 25655 3599 25669 3613
rect 31439 3599 31453 3613
rect 31463 3599 31477 3613
rect 38855 3599 38869 3613
rect 38879 3599 38893 3613
rect 39047 3599 39061 3613
rect 39215 3599 39229 3613
rect 39263 3599 39277 3613
rect 39287 3599 39301 3613
rect 39359 3599 39373 3613
rect 39503 3599 39517 3613
rect 39551 3599 39565 3613
rect 39599 3599 39613 3613
rect 39647 3599 39661 3613
rect 39671 3599 39685 3613
rect 40055 3599 40069 3613
rect 40391 3599 40405 3613
rect 40439 3599 40453 3613
rect 40463 3599 40477 3613
rect 40775 3599 40789 3613
rect 40799 3599 40813 3613
rect 40871 3599 40885 3613
rect 41039 3599 41053 3613
rect 41087 3599 41101 3613
rect 41159 3599 41173 3613
rect 41231 3599 41245 3613
rect 41303 3599 41317 3613
rect 41327 3599 41341 3613
rect 41399 3599 41413 3613
rect 13007 3575 13021 3589
rect 13103 3575 13117 3589
rect 13127 3575 13141 3589
rect 13199 3575 13213 3589
rect 13271 3575 13285 3589
rect 15839 3575 15853 3589
rect 15863 3575 15877 3589
rect 18431 3575 18445 3589
rect 18455 3575 18469 3589
rect 26831 3575 26845 3589
rect 26879 3575 26893 3589
rect 30671 3575 30685 3589
rect 30695 3575 30709 3589
rect 34967 3575 34981 3589
rect 34991 3575 35005 3589
rect 39167 3575 39181 3589
rect 39191 3575 39205 3589
rect 39455 3575 39469 3589
rect 39479 3575 39493 3589
rect 40151 3575 40165 3589
rect 40175 3575 40189 3589
rect 40247 3575 40261 3589
rect 40271 3575 40285 3589
rect 40343 3575 40357 3589
rect 40367 3575 40381 3589
rect 40991 3575 41005 3589
rect 41015 3575 41029 3589
rect 41495 3575 41509 3589
rect 41855 3575 41869 3589
rect 41903 3575 41917 3589
rect 12983 3551 12997 3565
rect 30431 3551 30445 3565
rect 30455 3551 30469 3565
rect 32207 3551 32221 3565
rect 32687 3551 32701 3565
rect 32807 3551 32821 3565
rect 32831 3551 32845 3565
rect 33071 3551 33085 3565
rect 33095 3551 33109 3565
rect 41615 3551 41629 3565
rect 41663 3551 41677 3565
rect 41711 3551 41725 3565
rect 41735 3551 41749 3565
rect 41807 3551 41821 3565
rect 41831 3551 41845 3565
rect 41999 3551 42013 3565
rect 42023 3551 42037 3565
rect 42119 3551 42133 3565
rect 12815 3527 12829 3541
rect 12863 3527 12877 3541
rect 12935 3527 12949 3541
rect 13583 3527 13597 3541
rect 13607 3527 13621 3541
rect 32831 3527 32845 3541
rect 59759 3767 59773 3781
rect 59759 3719 59773 3733
rect 40415 3527 40429 3541
rect 40439 3527 40453 3541
rect 42215 3527 42229 3541
rect 59039 3527 59053 3541
rect 59639 3527 59653 3541
rect 59759 3527 59773 3541
rect 12695 3503 12709 3517
rect 12767 3503 12781 3517
rect 12791 3503 12805 3517
rect 26975 3503 26989 3517
rect 27023 3503 27037 3517
rect 27695 3503 27709 3517
rect 34511 3503 34525 3517
rect 34535 3503 34549 3517
rect 35471 3503 35485 3517
rect 39431 3503 39445 3517
rect 39455 3503 39469 3517
rect 42335 3503 42349 3517
rect 12623 3479 12637 3493
rect 19079 3479 19093 3493
rect 19127 3479 19141 3493
rect 33383 3479 33397 3493
rect 33431 3479 33445 3493
rect 42455 3479 42469 3493
rect 12575 3455 12589 3469
rect 13487 3455 13501 3469
rect 13511 3455 13525 3469
rect 25415 3455 25429 3469
rect 30743 3455 30757 3469
rect 34079 3455 34093 3469
rect 39095 3455 39109 3469
rect 40895 3455 40909 3469
rect 42599 3455 42613 3469
rect 12359 3431 12373 3445
rect 12431 3431 12445 3445
rect 12551 3431 12565 3445
rect 20567 3431 20581 3445
rect 20591 3431 20605 3445
rect 22799 3431 22813 3445
rect 22847 3431 22861 3445
rect 31799 3431 31813 3445
rect 31847 3431 31861 3445
rect 32207 3431 32221 3445
rect 35543 3431 35557 3445
rect 35567 3431 35581 3445
rect 42695 3431 42709 3445
rect 12263 3407 12277 3421
rect 12311 3407 12325 3421
rect 12335 3407 12349 3421
rect 32759 3407 32773 3421
rect 33071 3407 33085 3421
rect 35423 3407 35437 3421
rect 35447 3407 35461 3421
rect 42815 3407 42829 3421
rect 12167 3383 12181 3397
rect 12215 3383 12229 3397
rect 12239 3383 12253 3397
rect 13127 3383 13141 3397
rect 13151 3383 13165 3397
rect 12095 3359 12109 3373
rect 24647 3359 24661 3373
rect 27839 3359 27853 3373
rect 27887 3359 27901 3373
rect 37103 3383 37117 3397
rect 37127 3383 37141 3397
rect 42935 3383 42949 3397
rect 33575 3359 33589 3373
rect 33599 3359 33613 3373
rect 43055 3359 43069 3373
rect 43415 3359 43429 3373
rect 43463 3359 43477 3373
rect 12047 3335 12061 3349
rect 27551 3335 27565 3349
rect 27599 3335 27613 3349
rect 34871 3335 34885 3349
rect 34895 3335 34909 3349
rect 43151 3335 43165 3349
rect 43199 3335 43213 3349
rect 43271 3335 43285 3349
rect 43319 3335 43333 3349
rect 43367 3335 43381 3349
rect 43391 3335 43405 3349
rect 43559 3335 43573 3349
rect 43607 3335 43621 3349
rect 43655 3335 43669 3349
rect 11999 3311 12013 3325
rect 23687 3311 23701 3325
rect 23711 3311 23725 3325
rect 31631 3311 31645 3325
rect 32207 3311 32221 3325
rect 35735 3311 35749 3325
rect 35759 3311 35773 3325
rect 40223 3311 40237 3325
rect 40247 3311 40261 3325
rect 43751 3311 43765 3325
rect 59039 3479 59053 3493
rect 59639 3479 59653 3493
rect 59759 3479 59773 3493
rect 11951 3287 11965 3301
rect 18095 3287 18109 3301
rect 43871 3287 43885 3301
rect 44015 3287 44029 3301
rect 44063 3287 44077 3301
rect 58919 3287 58933 3301
rect 59039 3287 59053 3301
rect 59639 3287 59653 3301
rect 59759 3287 59773 3301
rect 11927 3263 11941 3277
rect 43967 3263 43981 3277
rect 43991 3263 44005 3277
rect 44183 3263 44197 3277
rect 11903 3239 11917 3253
rect 15071 3239 15085 3253
rect 15095 3239 15109 3253
rect 44351 3239 44365 3253
rect 44399 3239 44413 3253
rect 44471 3239 44485 3253
rect 11879 3215 11893 3229
rect 22343 3215 22357 3229
rect 22367 3215 22381 3229
rect 44567 3215 44581 3229
rect 11855 3191 11869 3205
rect 12359 3191 12373 3205
rect 12383 3191 12397 3205
rect 28079 3191 28093 3205
rect 28103 3191 28117 3205
rect 28319 3191 28333 3205
rect 44711 3191 44725 3205
rect 11807 3167 11821 3181
rect 13391 3167 13405 3181
rect 13415 3167 13429 3181
rect 22775 3167 22789 3181
rect 22799 3167 22813 3181
rect 44807 3167 44821 3181
rect 11783 3143 11797 3157
rect 21479 3143 21493 3157
rect 21503 3143 21517 3157
rect 32207 3143 32221 3157
rect 35039 3143 35053 3157
rect 38039 3143 38053 3157
rect 44903 3143 44917 3157
rect 11711 3119 11725 3133
rect 12671 3119 12685 3133
rect 12719 3119 12733 3133
rect 33431 3119 33445 3133
rect 36527 3119 36541 3133
rect 36551 3119 36565 3133
rect 40631 3119 40645 3133
rect 40655 3119 40669 3133
rect 44447 3119 44461 3133
rect 44471 3119 44485 3133
rect 44999 3119 45013 3133
rect 11687 3095 11701 3109
rect 20711 3095 20725 3109
rect 20735 3095 20749 3109
rect 45119 3095 45133 3109
rect 11663 3071 11677 3085
rect 11711 3071 11725 3085
rect 11735 3071 11749 3085
rect 21935 3071 21949 3085
rect 21959 3071 21973 3085
rect 30095 3071 30109 3085
rect 30119 3071 30133 3085
rect 33671 3071 33685 3085
rect 33695 3071 33709 3085
rect 45215 3071 45229 3085
rect 11615 3047 11629 3061
rect 17135 3047 17149 3061
rect 17159 3047 17173 3061
rect 31967 3047 31981 3061
rect 31991 3047 32005 3061
rect 32207 3047 32221 3061
rect 33791 3047 33805 3061
rect 33815 3047 33829 3061
rect 39335 3047 39349 3061
rect 39359 3047 39373 3061
rect 45335 3047 45349 3061
rect 11591 3023 11605 3037
rect 22679 3023 22693 3037
rect 22703 3023 22717 3037
rect 27863 3023 27877 3037
rect 27911 3023 27925 3037
rect 34415 3023 34429 3037
rect 34439 3023 34453 3037
rect 45455 3023 45469 3037
rect 11567 2999 11581 3013
rect 30575 2999 30589 3013
rect 32207 2999 32221 3013
rect 39239 2999 39253 3013
rect 39263 2999 39277 3013
rect 45551 2999 45565 3013
rect 11519 2975 11533 2989
rect 22175 2975 22189 2989
rect 22223 2975 22237 2989
rect 30311 2975 30325 2989
rect 30335 2975 30349 2989
rect 32375 2975 32389 2989
rect 32639 2975 32653 2989
rect 11447 2951 11461 2965
rect 16703 2951 16717 2965
rect 16727 2951 16741 2965
rect 11423 2927 11437 2941
rect 16055 2927 16069 2941
rect 16079 2927 16093 2941
rect 32735 2975 32749 2989
rect 32807 2975 32821 2989
rect 33047 2975 33061 2989
rect 33191 2975 33205 2989
rect 33863 2975 33877 2989
rect 34751 2975 34765 2989
rect 42551 2975 42565 2989
rect 44639 2975 44653 2989
rect 45647 2975 45661 2989
rect 11399 2903 11413 2917
rect 32279 2903 32293 2917
rect 32303 2903 32317 2917
rect 32639 2903 32653 2917
rect 32663 2903 32677 2917
rect 32807 2951 32821 2965
rect 33263 2951 33277 2965
rect 33311 2951 33325 2965
rect 45767 2951 45781 2965
rect 45815 2951 45829 2965
rect 45863 2951 45877 2965
rect 45887 2951 45901 2965
rect 45959 2951 45973 2965
rect 33335 2927 33349 2941
rect 33359 2927 33373 2941
rect 46055 2927 46069 2941
rect 46079 2927 46093 2941
rect 46151 2927 46165 2941
rect 32759 2903 32773 2917
rect 32999 2903 33013 2917
rect 33383 2903 33397 2917
rect 33407 2903 33421 2917
rect 43487 2903 43501 2917
rect 43511 2903 43525 2917
rect 46247 2903 46261 2917
rect 11351 2879 11365 2893
rect 32255 2879 32269 2893
rect 32279 2879 32293 2893
rect 46367 2879 46381 2893
rect 46895 2879 46909 2893
rect 46943 2879 46957 2893
rect 11279 2855 11293 2869
rect 16271 2855 16285 2869
rect 16295 2855 16309 2869
rect 31943 2855 31957 2869
rect 31967 2855 31981 2869
rect 11255 2831 11269 2845
rect 12935 2831 12949 2845
rect 12959 2831 12973 2845
rect 31919 2831 31933 2845
rect 31943 2831 31957 2845
rect 33623 2855 33637 2869
rect 35927 2855 35941 2869
rect 35951 2855 35965 2869
rect 40319 2855 40333 2869
rect 40343 2855 40357 2869
rect 46463 2855 46477 2869
rect 46487 2855 46501 2869
rect 46559 2855 46573 2869
rect 46871 2855 46885 2869
rect 47063 2855 47077 2869
rect 47087 2855 47101 2869
rect 47159 2855 47173 2869
rect 43535 2831 43549 2845
rect 43559 2831 43573 2845
rect 46679 2831 46693 2845
rect 46703 2831 46717 2845
rect 46823 2831 46837 2845
rect 46847 2831 46861 2845
rect 47255 2831 47269 2845
rect 47543 2831 47557 2845
rect 47591 2831 47605 2845
rect 11231 2807 11245 2821
rect 32447 2807 32461 2821
rect 32639 2807 32653 2821
rect 39935 2807 39949 2821
rect 39959 2807 39973 2821
rect 44327 2807 44341 2821
rect 44351 2807 44365 2821
rect 44615 2807 44629 2821
rect 44951 2807 44965 2821
rect 45047 2807 45061 2821
rect 47375 2807 47389 2821
rect 47519 2807 47533 2821
rect 47711 2807 47725 2821
rect 47735 2807 47749 2821
rect 47831 2807 47845 2821
rect 47951 2807 47965 2821
rect 47999 2807 48013 2821
rect 11183 2783 11197 2797
rect 19367 2783 19381 2797
rect 19391 2783 19405 2797
rect 29999 2783 30013 2797
rect 30023 2783 30037 2797
rect 36407 2783 36421 2797
rect 47471 2783 47485 2797
rect 47495 2783 47509 2797
rect 48119 2783 48133 2797
rect 11135 2759 11149 2773
rect 27527 2759 27541 2773
rect 27551 2759 27565 2773
rect 41783 2759 41797 2773
rect 41807 2759 41821 2773
rect 48263 2759 48277 2773
rect 11039 2735 11053 2749
rect 11231 2735 11245 2749
rect 11303 2735 11317 2749
rect 24215 2735 24229 2749
rect 24287 2735 24301 2749
rect 32207 2735 32221 2749
rect 37847 2735 37861 2749
rect 37895 2735 37909 2749
rect 43679 2735 43693 2749
rect 43847 2735 43861 2749
rect 43871 2735 43885 2749
rect 48383 2735 48397 2749
rect 48407 2735 48421 2749
rect 48479 2735 48493 2749
rect 11015 2711 11029 2725
rect 11879 2711 11893 2725
rect 11975 2711 11989 2725
rect 18767 2711 18781 2725
rect 18791 2711 18805 2725
rect 20927 2711 20941 2725
rect 25367 2711 25381 2725
rect 25391 2711 25405 2725
rect 31511 2711 31525 2725
rect 31535 2711 31549 2725
rect 36119 2711 36133 2725
rect 36143 2711 36157 2725
rect 37919 2711 37933 2725
rect 38327 2711 38341 2725
rect 38783 2711 38797 2725
rect 42791 2711 42805 2725
rect 42815 2711 42829 2725
rect 48575 2711 48589 2725
rect 10943 2687 10957 2701
rect 31751 2687 31765 2701
rect 31775 2687 31789 2701
rect 32207 2687 32221 2701
rect 33479 2687 33493 2701
rect 33503 2687 33517 2701
rect 35495 2687 35509 2701
rect 44135 2687 44149 2701
rect 48671 2687 48685 2701
rect 48719 2687 48733 2701
rect 48767 2687 48781 2701
rect 10847 2663 10861 2677
rect 10895 2663 10909 2677
rect 10919 2663 10933 2677
rect 31391 2663 31405 2677
rect 31439 2663 31453 2677
rect 37199 2663 37213 2677
rect 37223 2663 37237 2677
rect 43439 2663 43453 2677
rect 43463 2663 43477 2677
rect 48863 2663 48877 2677
rect 10823 2639 10837 2653
rect 12815 2639 12829 2653
rect 12839 2639 12853 2653
rect 13367 2639 13381 2653
rect 13391 2639 13405 2653
rect 32207 2639 32221 2653
rect 36959 2639 36973 2653
rect 39911 2639 39925 2653
rect 46751 2639 46765 2653
rect 48599 2639 48613 2653
rect 48959 2639 48973 2653
rect 10775 2615 10789 2629
rect 41375 2615 41389 2629
rect 41399 2615 41413 2629
rect 41543 2615 41557 2629
rect 42863 2615 42877 2629
rect 42959 2615 42973 2629
rect 44495 2615 44509 2629
rect 48359 2615 48373 2629
rect 48383 2615 48397 2629
rect 49055 2615 49069 2629
rect 49079 2615 49093 2629
rect 49151 2615 49165 2629
rect 10679 2591 10693 2605
rect 12623 2591 12637 2605
rect 12647 2591 12661 2605
rect 32207 2591 32221 2605
rect 36863 2591 36877 2605
rect 36887 2591 36901 2605
rect 41591 2591 41605 2605
rect 41615 2591 41629 2605
rect 42911 2591 42925 2605
rect 42935 2591 42949 2605
rect 43343 2591 43357 2605
rect 43367 2591 43381 2605
rect 47975 2591 47989 2605
rect 47999 2591 48013 2605
rect 49247 2591 49261 2605
rect 10631 2567 10645 2581
rect 15383 2567 15397 2581
rect 15407 2567 15421 2581
rect 21383 2567 21397 2581
rect 24839 2567 24853 2581
rect 24863 2567 24877 2581
rect 43799 2567 43813 2581
rect 46967 2567 46981 2581
rect 49343 2567 49357 2581
rect 10295 2543 10309 2557
rect 10391 2543 10405 2557
rect 10607 2543 10621 2557
rect 12527 2543 12541 2557
rect 12599 2543 12613 2557
rect 21719 2543 21733 2557
rect 21743 2543 21757 2557
rect 22487 2543 22501 2557
rect 24767 2543 24781 2557
rect 25079 2543 25093 2557
rect 26639 2543 26653 2557
rect 29975 2543 29989 2557
rect 29999 2543 30013 2557
rect 34007 2543 34021 2557
rect 34031 2543 34045 2557
rect 36647 2543 36661 2557
rect 36671 2543 36685 2557
rect 39815 2543 39829 2557
rect 42503 2543 42517 2557
rect 48623 2543 48637 2557
rect 49439 2543 49453 2557
rect 10175 2519 10189 2533
rect 10247 2519 10261 2533
rect 10271 2519 10285 2533
rect 10487 2519 10501 2533
rect 10511 2519 10525 2533
rect 11903 2519 11917 2533
rect 12023 2519 12037 2533
rect 16487 2519 16501 2533
rect 16511 2519 16525 2533
rect 23999 2519 24013 2533
rect 24023 2519 24037 2533
rect 26999 2519 27013 2533
rect 27047 2519 27061 2533
rect 29207 2519 29221 2533
rect 32999 2519 33013 2533
rect 49535 2519 49549 2533
rect 10127 2495 10141 2509
rect 32207 2495 32221 2509
rect 38735 2495 38749 2509
rect 38759 2495 38773 2509
rect 40847 2495 40861 2509
rect 40871 2495 40885 2509
rect 46535 2495 46549 2509
rect 46559 2495 46573 2509
rect 49631 2495 49645 2509
rect 10079 2471 10093 2485
rect 11783 2471 11797 2485
rect 11831 2471 11845 2485
rect 32639 2471 32653 2485
rect 32735 2471 32749 2485
rect 32759 2471 32773 2485
rect 32975 2471 32989 2485
rect 37367 2471 37381 2485
rect 41879 2471 41893 2485
rect 41903 2471 41917 2485
rect 49727 2471 49741 2485
rect 10055 2447 10069 2461
rect 32759 2447 32773 2461
rect 32975 2447 32989 2461
rect 38927 2447 38941 2461
rect 38951 2447 38965 2461
rect 41423 2447 41437 2461
rect 46031 2447 46045 2461
rect 46055 2447 46069 2461
rect 49847 2447 49861 2461
rect 50015 2447 50029 2461
rect 50063 2447 50077 2461
rect 9959 2423 9973 2437
rect 11855 2423 11869 2437
rect 11879 2423 11893 2437
rect 19487 2423 19501 2437
rect 19511 2423 19525 2437
rect 22247 2423 22261 2437
rect 22271 2423 22285 2437
rect 22871 2423 22885 2437
rect 42311 2423 42325 2437
rect 42335 2423 42349 2437
rect 49967 2423 49981 2437
rect 49991 2423 50005 2437
rect 50159 2423 50173 2437
rect 9935 2399 9949 2413
rect 32207 2399 32221 2413
rect 45311 2399 45325 2413
rect 45335 2399 45349 2413
rect 45623 2399 45637 2413
rect 45647 2399 45661 2413
rect 50255 2399 50269 2413
rect 9911 2375 9925 2389
rect 10847 2375 10861 2389
rect 10871 2375 10885 2389
rect 17567 2375 17581 2389
rect 17591 2375 17605 2389
rect 31823 2375 31837 2389
rect 31871 2375 31885 2389
rect 48839 2375 48853 2389
rect 48863 2375 48877 2389
rect 50351 2375 50365 2389
rect 9863 2351 9877 2365
rect 14735 2351 14749 2365
rect 14759 2351 14773 2365
rect 18263 2351 18277 2365
rect 18311 2351 18325 2365
rect 32207 2351 32221 2365
rect 44543 2351 44557 2365
rect 44567 2351 44581 2365
rect 50831 2351 50845 2365
rect 9839 2327 9853 2341
rect 10583 2327 10597 2341
rect 10655 2327 10669 2341
rect 20351 2327 20365 2341
rect 20399 2327 20413 2341
rect 38279 2327 38293 2341
rect 38303 2327 38317 2341
rect 46799 2327 46813 2341
rect 46823 2327 46837 2341
rect 49271 2327 49285 2341
rect 50879 2327 50893 2341
rect 51023 2327 51037 2341
rect 51071 2327 51085 2341
rect 9815 2303 9829 2317
rect 13823 2303 13837 2317
rect 51167 2303 51181 2317
rect 51215 2303 51229 2317
rect 51263 2303 51277 2317
rect 9767 2279 9781 2293
rect 10127 2279 10141 2293
rect 10151 2279 10165 2293
rect 23279 2279 23293 2293
rect 23375 2279 23389 2293
rect 31727 2279 31741 2293
rect 31751 2279 31765 2293
rect 35063 2279 35077 2293
rect 35087 2279 35101 2293
rect 40031 2279 40045 2293
rect 40055 2279 40069 2293
rect 47039 2279 47053 2293
rect 47063 2279 47077 2293
rect 50087 2279 50101 2293
rect 51383 2279 51397 2293
rect 9695 2255 9709 2269
rect 13679 2255 13693 2269
rect 13703 2255 13717 2269
rect 14015 2255 14029 2269
rect 14039 2255 14053 2269
rect 15167 2255 15181 2269
rect 15503 2255 15517 2269
rect 15719 2255 15733 2269
rect 15935 2255 15949 2269
rect 16151 2255 16165 2269
rect 16367 2255 16381 2269
rect 16583 2255 16597 2269
rect 16799 2255 16813 2269
rect 17015 2255 17029 2269
rect 17231 2255 17245 2269
rect 17351 2255 17365 2269
rect 17375 2255 17389 2269
rect 32591 2255 32605 2269
rect 32903 2255 32917 2269
rect 47687 2255 47701 2269
rect 47711 2255 47725 2269
rect 49367 2255 49381 2269
rect 51503 2255 51517 2269
rect 8687 2231 8701 2245
rect 8735 2231 8749 2245
rect 8759 2231 8773 2245
rect 8831 2231 8845 2245
rect 9671 2231 9685 2245
rect 11015 2231 11029 2245
rect 11063 2231 11077 2245
rect 23807 2231 23821 2245
rect 23831 2231 23845 2245
rect 24191 2231 24205 2245
rect 32183 2231 32197 2245
rect 32207 2231 32221 2245
rect 35831 2231 35845 2245
rect 35855 2231 35869 2245
rect 43943 2231 43957 2245
rect 43967 2231 43981 2245
rect 48167 2231 48181 2245
rect 49751 2231 49765 2245
rect 51599 2231 51613 2245
rect 51671 2231 51685 2245
rect 51719 2231 51733 2245
rect 8567 2207 8581 2221
rect 8639 2207 8653 2221
rect 8663 2207 8677 2221
rect 8927 2207 8941 2221
rect 8951 2207 8965 2221
rect 9023 2207 9037 2221
rect 9647 2207 9661 2221
rect 37703 2207 37717 2221
rect 41639 2207 41653 2221
rect 43295 2207 43309 2221
rect 51791 2207 51805 2221
rect 51863 2207 51877 2221
rect 8543 2183 8557 2197
rect 9119 2183 9133 2197
rect 9167 2183 9181 2197
rect 9215 2183 9229 2197
rect 9431 2183 9445 2197
rect 9527 2183 9541 2197
rect 9551 2183 9565 2197
rect 9839 2183 9853 2197
rect 9887 2183 9901 2197
rect 14999 2183 15013 2197
rect 15047 2183 15061 2197
rect 22199 2183 22213 2197
rect 22247 2183 22261 2197
rect 35303 2183 35317 2197
rect 35327 2183 35341 2197
rect 49223 2183 49237 2197
rect 49247 2183 49261 2197
rect 51983 2183 51997 2197
rect 8303 2159 8317 2173
rect 8399 2159 8413 2173
rect 8519 2159 8533 2173
rect 9311 2159 9325 2173
rect 9335 2159 9349 2173
rect 11159 2159 11173 2173
rect 11207 2159 11221 2173
rect 18599 2159 18613 2173
rect 18647 2159 18661 2173
rect 24551 2159 24565 2173
rect 24575 2159 24589 2173
rect 41687 2159 41701 2173
rect 41711 2159 41725 2173
rect 50039 2159 50053 2173
rect 50063 2159 50077 2173
rect 52103 2159 52117 2173
rect 8207 2135 8221 2149
rect 32207 2135 32221 2149
rect 32231 2135 32245 2149
rect 45407 2135 45421 2149
rect 52199 2135 52213 2149
rect 8183 2111 8197 2125
rect 14663 2111 14677 2125
rect 14687 2111 14701 2125
rect 48095 2111 48109 2125
rect 48119 2111 48133 2125
rect 49391 2111 49405 2125
rect 52319 2111 52333 2125
rect 8111 2087 8125 2101
rect 8759 2087 8773 2101
rect 8783 2087 8797 2101
rect 8879 2087 8893 2101
rect 9071 2087 9085 2101
rect 9263 2087 9277 2101
rect 12575 2087 12589 2101
rect 12623 2087 12637 2101
rect 32903 2087 32917 2101
rect 32951 2087 32965 2101
rect 34391 2087 34405 2101
rect 38399 2087 38413 2101
rect 38423 2087 38437 2101
rect 39839 2087 39853 2101
rect 39863 2087 39877 2101
rect 44039 2087 44053 2101
rect 44063 2087 44077 2101
rect 49463 2087 49477 2101
rect 49895 2087 49909 2101
rect 52439 2087 52453 2101
rect 8087 2063 8101 2077
rect 9335 2063 9349 2077
rect 9359 2063 9373 2077
rect 10823 2063 10837 2077
rect 10847 2063 10861 2077
rect 18623 2063 18637 2077
rect 18671 2063 18685 2077
rect 23879 2063 23893 2077
rect 23903 2063 23917 2077
rect 24887 2063 24901 2077
rect 24983 2063 24997 2077
rect 25007 2063 25021 2077
rect 27167 2063 27181 2077
rect 30863 2063 30877 2077
rect 41759 2063 41773 2077
rect 51911 2063 51925 2077
rect 52559 2063 52573 2077
rect 8063 2039 8077 2053
rect 22727 2039 22741 2053
rect 52679 2039 52693 2053
rect 8039 2015 8053 2029
rect 8567 2015 8581 2029
rect 8591 2015 8605 2029
rect 13559 2015 13573 2029
rect 13583 2015 13597 2029
rect 20951 2015 20965 2029
rect 20999 2015 21013 2029
rect 22943 2015 22957 2029
rect 22967 2015 22981 2029
rect 37991 2015 38005 2029
rect 46991 2015 47005 2029
rect 47279 2015 47293 2029
rect 52799 2015 52813 2029
rect 8015 1991 8029 2005
rect 8903 1991 8917 2005
rect 17879 1991 17893 2005
rect 32471 1991 32485 2005
rect 32591 1991 32605 2005
rect 32663 1991 32677 2005
rect 32879 1991 32893 2005
rect 32927 1991 32941 2005
rect 43031 1991 43045 2005
rect 43055 1991 43069 2005
rect 51143 1991 51157 2005
rect 51167 1991 51181 2005
rect 52895 1991 52909 2005
rect 7967 1967 7981 1981
rect 9287 1967 9301 1981
rect 17663 1967 17677 1981
rect 32663 1967 32677 1981
rect 32879 1967 32893 1981
rect 35711 1967 35725 1981
rect 40607 1967 40621 1981
rect 47303 1967 47317 1981
rect 51743 1967 51757 1981
rect 53015 1967 53029 1981
rect 7943 1943 7957 1957
rect 10679 1943 10693 1957
rect 10703 1943 10717 1957
rect 19271 1943 19285 1957
rect 19295 1943 19309 1957
rect 48239 1943 48253 1957
rect 48263 1943 48277 1957
rect 50135 1943 50149 1957
rect 50159 1943 50173 1957
rect 53135 1943 53149 1957
rect 7895 1919 7909 1933
rect 11039 1919 11053 1933
rect 11087 1919 11101 1933
rect 13871 1919 13885 1933
rect 13895 1919 13909 1933
rect 14111 1919 14125 1933
rect 15239 1919 15253 1933
rect 15575 1919 15589 1933
rect 15791 1919 15805 1933
rect 16007 1919 16021 1933
rect 16223 1919 16237 1933
rect 16439 1919 16453 1933
rect 16655 1919 16669 1933
rect 16871 1919 16885 1933
rect 16919 1919 16933 1933
rect 16943 1919 16957 1933
rect 19247 1919 19261 1933
rect 19271 1919 19285 1933
rect 19799 1919 19813 1933
rect 19823 1919 19837 1933
rect 24263 1919 24277 1933
rect 24311 1919 24325 1933
rect 49127 1919 49141 1933
rect 49151 1919 49165 1933
rect 53231 1919 53245 1933
rect 7871 1895 7885 1909
rect 12263 1895 12277 1909
rect 12287 1895 12301 1909
rect 26015 1895 26029 1909
rect 35615 1895 35629 1909
rect 37607 1895 37621 1909
rect 38255 1895 38269 1909
rect 47111 1895 47125 1909
rect 50303 1895 50317 1909
rect 51767 1895 51781 1909
rect 53375 1895 53389 1909
rect 7823 1871 7837 1885
rect 10751 1871 10765 1885
rect 10799 1871 10813 1885
rect 18551 1871 18565 1885
rect 18575 1871 18589 1885
rect 22391 1871 22405 1885
rect 22439 1871 22453 1885
rect 33335 1871 33349 1885
rect 38351 1871 38365 1885
rect 44927 1871 44941 1885
rect 47207 1871 47221 1885
rect 47879 1871 47893 1885
rect 48431 1871 48445 1885
rect 51647 1871 51661 1885
rect 53471 1871 53485 1885
rect 7727 1847 7741 1861
rect 8543 1847 8557 1861
rect 8567 1847 8581 1861
rect 11255 1847 11269 1861
rect 11327 1847 11341 1861
rect 11687 1847 11701 1861
rect 11711 1847 11725 1861
rect 28583 1847 28597 1861
rect 28607 1847 28621 1861
rect 30815 1847 30829 1861
rect 30935 1847 30949 1861
rect 31079 1847 31093 1861
rect 31319 1847 31333 1861
rect 31535 1847 31549 1861
rect 31559 1847 31573 1861
rect 37631 1847 37645 1861
rect 43127 1847 43141 1861
rect 43151 1847 43165 1861
rect 44231 1847 44245 1861
rect 44423 1847 44437 1861
rect 53591 1847 53605 1861
rect 7583 1823 7597 1837
rect 9959 1823 9973 1837
rect 9983 1823 9997 1837
rect 36767 1823 36781 1837
rect 36791 1823 36805 1837
rect 50327 1823 50341 1837
rect 50351 1823 50365 1837
rect 51239 1823 51253 1837
rect 51263 1823 51277 1837
rect 53639 1823 53653 1837
rect 7175 1799 7189 1813
rect 11615 1799 11629 1813
rect 11639 1799 11653 1813
rect 24239 1799 24253 1813
rect 24263 1799 24277 1813
rect 36023 1799 36037 1813
rect 36047 1799 36061 1813
rect 41063 1799 41077 1813
rect 41087 1799 41101 1813
rect 44783 1799 44797 1813
rect 44807 1799 44821 1813
rect 45935 1799 45949 1813
rect 45959 1799 45973 1813
rect 53663 1799 53677 1813
rect 6959 1775 6973 1789
rect 32591 1775 32605 1789
rect 32759 1775 32773 1789
rect 44159 1775 44173 1789
rect 44183 1775 44197 1789
rect 51695 1775 51709 1789
rect 51719 1775 51733 1789
rect 53687 1775 53701 1789
rect 6911 1751 6925 1765
rect 8063 1751 8077 1765
rect 8135 1751 8149 1765
rect 12239 1751 12253 1765
rect 12263 1751 12277 1765
rect 18335 1751 18349 1765
rect 18359 1751 18373 1765
rect 33983 1751 33997 1765
rect 40679 1751 40693 1765
rect 42623 1751 42637 1765
rect 46223 1751 46237 1765
rect 46247 1751 46261 1765
rect 50855 1751 50869 1765
rect 50879 1751 50893 1765
rect 53711 1751 53725 1765
rect 6263 1727 6277 1741
rect 6359 1727 6373 1741
rect 6383 1727 6397 1741
rect 6455 1727 6469 1741
rect 6551 1727 6565 1741
rect 22199 1727 22213 1741
rect 38159 1727 38173 1741
rect 38183 1727 38197 1741
rect 40535 1727 40549 1741
rect 40559 1727 40573 1741
rect 48455 1727 48469 1741
rect 48479 1727 48493 1741
rect 49175 1727 49189 1741
rect 50183 1727 50197 1741
rect 53783 1727 53797 1741
rect 6071 1703 6085 1717
rect 6143 1703 6157 1717
rect 6167 1703 6181 1717
rect 10511 1703 10525 1717
rect 10535 1703 10549 1717
rect 11663 1703 11677 1717
rect 11687 1703 11701 1717
rect 11807 1703 11821 1717
rect 11855 1703 11869 1717
rect 11927 1703 11941 1717
rect 12071 1703 12085 1717
rect 20207 1703 20221 1717
rect 20231 1703 20245 1717
rect 36215 1703 36229 1717
rect 39575 1703 39589 1717
rect 43895 1703 43909 1717
rect 48791 1703 48805 1717
rect 49007 1703 49021 1717
rect 49103 1703 49117 1717
rect 51311 1703 51325 1717
rect 51887 1703 51901 1717
rect 52031 1703 52045 1717
rect 53903 1703 53917 1717
rect 5831 1679 5845 1693
rect 5927 1679 5941 1693
rect 5951 1679 5965 1693
rect 9623 1679 9637 1693
rect 9719 1679 9733 1693
rect 21263 1679 21277 1693
rect 21287 1679 21301 1693
rect 24527 1679 24541 1693
rect 24551 1679 24565 1693
rect 33119 1679 33133 1693
rect 33143 1679 33157 1693
rect 45743 1679 45757 1693
rect 45767 1679 45781 1693
rect 49703 1679 49717 1693
rect 49727 1679 49741 1693
rect 53999 1679 54013 1693
rect 5783 1655 5797 1669
rect 36431 1655 36445 1669
rect 36455 1655 36469 1669
rect 54095 1655 54109 1669
rect 5759 1631 5773 1645
rect 11855 1631 11869 1645
rect 11903 1631 11917 1645
rect 13463 1631 13477 1645
rect 13487 1631 13501 1645
rect 22559 1631 22573 1645
rect 22583 1631 22597 1645
rect 26447 1631 26461 1645
rect 26471 1631 26485 1645
rect 42575 1631 42589 1645
rect 42599 1631 42613 1645
rect 44975 1631 44989 1645
rect 44999 1631 45013 1645
rect 46583 1631 46597 1645
rect 52415 1631 52429 1645
rect 52439 1631 52453 1645
rect 52943 1631 52957 1645
rect 54119 1631 54133 1645
rect 5711 1607 5725 1621
rect 26855 1607 26869 1621
rect 26903 1607 26917 1621
rect 51191 1607 51205 1621
rect 51407 1607 51421 1621
rect 54215 1607 54229 1621
rect 5687 1583 5701 1597
rect 11111 1583 11125 1597
rect 11999 1583 12013 1597
rect 12119 1583 12133 1597
rect 27455 1583 27469 1597
rect 27479 1583 27493 1597
rect 32591 1583 32605 1597
rect 32663 1583 32677 1597
rect 53615 1583 53629 1597
rect 53663 1583 53677 1597
rect 54263 1583 54277 1597
rect 5663 1559 5677 1573
rect 9863 1559 9877 1573
rect 9959 1559 9973 1573
rect 14567 1559 14581 1573
rect 14591 1559 14605 1573
rect 21623 1559 21637 1573
rect 21647 1559 21661 1573
rect 53111 1559 53125 1573
rect 53135 1559 53149 1573
rect 54287 1559 54301 1573
rect 5639 1535 5653 1549
rect 8039 1535 8053 1549
rect 8063 1535 8077 1549
rect 11351 1535 11365 1549
rect 11375 1535 11389 1549
rect 11591 1535 11605 1549
rect 11615 1535 11629 1549
rect 20183 1535 20197 1549
rect 38591 1535 38605 1549
rect 44303 1535 44317 1549
rect 46727 1535 46741 1549
rect 48911 1535 48925 1549
rect 52631 1535 52645 1549
rect 54311 1535 54325 1549
rect 5591 1511 5605 1525
rect 9167 1511 9181 1525
rect 9191 1511 9205 1525
rect 18287 1511 18301 1525
rect 18335 1511 18349 1525
rect 24503 1511 24517 1525
rect 24527 1511 24541 1525
rect 37007 1511 37021 1525
rect 37031 1511 37045 1525
rect 40007 1511 40021 1525
rect 40079 1511 40093 1525
rect 43079 1511 43093 1525
rect 47567 1511 47581 1525
rect 47591 1511 47605 1525
rect 54407 1511 54421 1525
rect 5543 1487 5557 1501
rect 9407 1487 9421 1501
rect 9455 1487 9469 1501
rect 15431 1487 15445 1501
rect 22511 1487 22525 1501
rect 43583 1487 43597 1501
rect 54551 1487 54565 1501
rect 5519 1463 5533 1477
rect 6959 1463 6973 1477
rect 6983 1463 6997 1477
rect 9647 1463 9661 1477
rect 9743 1463 9757 1477
rect 12911 1463 12925 1477
rect 14375 1463 14389 1477
rect 14399 1463 14413 1477
rect 37247 1463 37261 1477
rect 43631 1463 43645 1477
rect 43655 1463 43669 1477
rect 49415 1463 49429 1477
rect 49439 1463 49453 1477
rect 51287 1463 51301 1477
rect 51431 1463 51445 1477
rect 52007 1463 52021 1477
rect 54671 1463 54685 1477
rect 5495 1439 5509 1453
rect 13271 1439 13285 1453
rect 13295 1439 13309 1453
rect 32567 1439 32581 1453
rect 32663 1439 32677 1453
rect 37655 1439 37669 1453
rect 37679 1439 37693 1453
rect 44831 1439 44845 1453
rect 45383 1439 45397 1453
rect 52991 1439 53005 1453
rect 53015 1439 53029 1453
rect 54791 1439 54805 1453
rect 5471 1415 5485 1429
rect 7943 1415 7957 1429
rect 7991 1415 8005 1429
rect 10775 1415 10789 1429
rect 10823 1415 10837 1429
rect 18407 1415 18421 1429
rect 18431 1415 18445 1429
rect 28751 1415 28765 1429
rect 28775 1415 28789 1429
rect 30119 1415 30133 1429
rect 30143 1415 30157 1429
rect 36743 1415 36757 1429
rect 38999 1415 39013 1429
rect 42983 1415 42997 1429
rect 44735 1415 44749 1429
rect 45719 1415 45733 1429
rect 45791 1415 45805 1429
rect 45911 1415 45925 1429
rect 52871 1415 52885 1429
rect 52895 1415 52909 1429
rect 54239 1415 54253 1429
rect 54263 1415 54277 1429
rect 54335 1415 54349 1429
rect 54887 1415 54901 1429
rect 5447 1391 5461 1405
rect 10943 1391 10957 1405
rect 10967 1391 10981 1405
rect 20375 1391 20389 1405
rect 20423 1391 20437 1405
rect 26303 1391 26317 1405
rect 26327 1391 26341 1405
rect 30239 1391 30253 1405
rect 30263 1391 30277 1405
rect 53159 1391 53173 1405
rect 54983 1391 54997 1405
rect 5399 1367 5413 1381
rect 5471 1367 5485 1381
rect 5567 1367 5581 1381
rect 32735 1367 32749 1381
rect 32759 1367 32773 1381
rect 37751 1367 37765 1381
rect 37775 1367 37789 1381
rect 41975 1367 41989 1381
rect 41999 1367 42013 1381
rect 49511 1367 49525 1381
rect 49535 1367 49549 1381
rect 55079 1367 55093 1381
rect 5375 1343 5389 1357
rect 5663 1343 5677 1357
rect 5735 1343 5749 1357
rect 12047 1343 12061 1357
rect 12143 1343 12157 1357
rect 18911 1343 18925 1357
rect 18959 1343 18973 1357
rect 27959 1343 27973 1357
rect 27983 1343 27997 1357
rect 28079 1343 28093 1357
rect 34319 1343 34333 1357
rect 34343 1343 34357 1357
rect 43823 1343 43837 1357
rect 55151 1343 55165 1357
rect 5255 1319 5269 1333
rect 5327 1319 5341 1333
rect 5351 1319 5365 1333
rect 5759 1319 5773 1333
rect 5807 1319 5821 1333
rect 15359 1319 15373 1333
rect 15383 1319 15397 1333
rect 45983 1319 45997 1333
rect 48887 1319 48901 1333
rect 54647 1319 54661 1333
rect 54671 1319 54685 1333
rect 54815 1319 54829 1333
rect 54911 1319 54925 1333
rect 55295 1319 55309 1333
rect 5231 1295 5245 1309
rect 11567 1295 11581 1309
rect 11591 1295 11605 1309
rect 12551 1295 12565 1309
rect 12575 1295 12589 1309
rect 25463 1295 25477 1309
rect 25487 1295 25501 1309
rect 27359 1295 27373 1309
rect 29183 1295 29197 1309
rect 34607 1295 34621 1309
rect 34631 1295 34645 1309
rect 36479 1295 36493 1309
rect 39023 1295 39037 1309
rect 39047 1295 39061 1309
rect 39071 1295 39085 1309
rect 45143 1295 45157 1309
rect 48935 1295 48949 1309
rect 48959 1295 48973 1309
rect 49559 1295 49573 1309
rect 49655 1295 49669 1309
rect 55391 1295 55405 1309
rect 5135 1271 5149 1285
rect 7799 1271 7813 1285
rect 7847 1271 7861 1285
rect 35639 1271 35653 1285
rect 35663 1271 35677 1285
rect 41279 1271 41293 1285
rect 41303 1271 41317 1285
rect 42263 1271 42277 1285
rect 45095 1271 45109 1285
rect 45119 1271 45133 1285
rect 51047 1271 51061 1285
rect 51071 1271 51085 1285
rect 55535 1271 55549 1285
rect 5111 1247 5125 1261
rect 8279 1247 8293 1261
rect 8327 1247 8341 1261
rect 9911 1247 9925 1261
rect 10007 1247 10021 1261
rect 37823 1247 37837 1261
rect 37871 1247 37885 1261
rect 40295 1247 40309 1261
rect 52055 1247 52069 1261
rect 55631 1247 55645 1261
rect 5039 1223 5053 1237
rect 7895 1223 7909 1237
rect 7919 1223 7933 1237
rect 30215 1223 30229 1237
rect 30239 1223 30253 1237
rect 38063 1223 38077 1237
rect 38087 1223 38101 1237
rect 42431 1223 42445 1237
rect 42455 1223 42469 1237
rect 49607 1223 49621 1237
rect 49631 1223 49645 1237
rect 53447 1223 53461 1237
rect 53471 1223 53485 1237
rect 55007 1223 55021 1237
rect 55343 1223 55357 1237
rect 55751 1223 55765 1237
rect 4991 1199 5005 1213
rect 6239 1199 6253 1213
rect 6287 1199 6301 1213
rect 7871 1199 7885 1213
rect 7895 1199 7909 1213
rect 9695 1199 9709 1213
rect 9767 1199 9781 1213
rect 4919 1175 4933 1189
rect 8303 1175 8317 1189
rect 8351 1175 8365 1189
rect 32423 1199 32437 1213
rect 32447 1199 32461 1213
rect 37559 1199 37573 1213
rect 37583 1199 37597 1213
rect 42095 1199 42109 1213
rect 42119 1199 42133 1213
rect 47807 1199 47821 1213
rect 47831 1199 47845 1213
rect 49871 1199 49885 1213
rect 55055 1199 55069 1213
rect 55079 1199 55093 1213
rect 55103 1199 55117 1213
rect 55847 1199 55861 1213
rect 9791 1175 9805 1189
rect 9839 1175 9853 1189
rect 33527 1175 33541 1189
rect 34175 1175 34189 1189
rect 34487 1175 34501 1189
rect 34559 1175 34573 1189
rect 36239 1175 36253 1189
rect 36263 1175 36277 1189
rect 43727 1175 43741 1189
rect 43751 1175 43765 1189
rect 47231 1175 47245 1189
rect 47255 1175 47269 1189
rect 50111 1175 50125 1189
rect 53663 1175 53677 1189
rect 53711 1175 53725 1189
rect 54767 1175 54781 1189
rect 54791 1175 54805 1189
rect 55775 1175 55789 1189
rect 55943 1175 55957 1189
rect 56039 1175 56053 1189
rect 56471 1175 56485 1189
rect 4895 1151 4909 1165
rect 5543 1151 5557 1165
rect 5615 1151 5629 1165
rect 9431 1151 9445 1165
rect 9479 1151 9493 1165
rect 12479 1151 12493 1165
rect 14255 1151 14269 1165
rect 14279 1151 14293 1165
rect 54143 1151 54157 1165
rect 56663 1151 56677 1165
rect 4847 1127 4861 1141
rect 6551 1127 6565 1141
rect 6575 1127 6589 1141
rect 7823 1127 7837 1141
rect 7871 1127 7885 1141
rect 22319 1127 22333 1141
rect 22343 1127 22357 1141
rect 27239 1127 27253 1141
rect 27263 1127 27277 1141
rect 30719 1127 30733 1141
rect 36311 1127 36325 1141
rect 36935 1127 36949 1141
rect 41567 1127 41581 1141
rect 46007 1127 46021 1141
rect 46103 1127 46117 1141
rect 46295 1127 46309 1141
rect 51575 1127 51589 1141
rect 51599 1127 51613 1141
rect 55271 1127 55285 1141
rect 55295 1127 55309 1141
rect 55463 1127 55477 1141
rect 55871 1127 55885 1141
rect 56687 1127 56701 1141
rect 4775 1103 4789 1117
rect 6263 1103 6277 1117
rect 6311 1103 6325 1117
rect 24479 1103 24493 1117
rect 24503 1103 24517 1117
rect 51839 1103 51853 1117
rect 51863 1103 51877 1117
rect 56783 1103 56797 1117
rect 4751 1079 4765 1093
rect 11735 1079 11749 1093
rect 11759 1079 11773 1093
rect 18935 1079 18949 1093
rect 18983 1079 18997 1093
rect 26351 1079 26365 1093
rect 26423 1079 26437 1093
rect 39623 1079 39637 1093
rect 39647 1079 39661 1093
rect 42743 1079 42757 1093
rect 47447 1079 47461 1093
rect 47471 1079 47485 1093
rect 52823 1079 52837 1093
rect 53591 1079 53605 1093
rect 53639 1079 53653 1093
rect 56879 1079 56893 1093
rect 4727 1055 4741 1069
rect 21719 1055 21733 1069
rect 28799 1055 28813 1069
rect 30599 1055 30613 1069
rect 39983 1055 39997 1069
rect 40703 1055 40717 1069
rect 41255 1055 41269 1069
rect 47663 1055 47677 1069
rect 53543 1055 53557 1069
rect 53567 1055 53581 1069
rect 56711 1055 56725 1069
rect 56975 1055 56989 1069
rect 4703 1031 4717 1045
rect 4895 1031 4909 1045
rect 4943 1031 4957 1045
rect 5711 1031 5725 1045
rect 5759 1031 5773 1045
rect 9551 1031 9565 1045
rect 9575 1031 9589 1045
rect 11015 1031 11029 1045
rect 12335 1031 12349 1045
rect 12359 1031 12373 1045
rect 14471 1031 14485 1045
rect 14495 1031 14509 1045
rect 33239 1031 33253 1045
rect 36983 1031 36997 1045
rect 40919 1031 40933 1045
rect 47423 1031 47437 1045
rect 47759 1031 47773 1045
rect 53327 1031 53341 1045
rect 57095 1031 57109 1045
rect 4679 1007 4693 1021
rect 11903 1007 11917 1021
rect 11927 1007 11941 1021
rect 23639 1007 23653 1021
rect 23663 1007 23677 1021
rect 41951 1007 41965 1021
rect 44855 1007 44869 1021
rect 51815 1007 51829 1021
rect 53303 1007 53317 1021
rect 53855 1007 53869 1021
rect 54695 1007 54709 1021
rect 57191 1007 57205 1021
rect 4583 983 4597 997
rect 4919 983 4933 997
rect 4967 983 4981 997
rect 5039 983 5053 997
rect 5063 983 5077 997
rect 8951 983 8965 997
rect 8975 983 8989 997
rect 9167 983 9181 997
rect 9359 983 9373 997
rect 9383 983 9397 997
rect 32807 983 32821 997
rect 32831 983 32845 997
rect 32855 983 32869 997
rect 47135 983 47149 997
rect 47159 983 47173 997
rect 47183 983 47197 997
rect 51479 983 51493 997
rect 51503 983 51517 997
rect 54191 983 54205 997
rect 54215 983 54229 997
rect 4535 959 4549 973
rect 5087 959 5101 973
rect 5159 959 5173 973
rect 8111 959 8125 973
rect 8159 959 8173 973
rect 9935 959 9949 973
rect 10031 959 10045 973
rect 19631 959 19645 973
rect 19655 959 19669 973
rect 24383 959 24397 973
rect 24407 959 24421 973
rect 31055 959 31069 973
rect 32807 959 32821 973
rect 46127 959 46141 973
rect 46151 959 46165 973
rect 46175 959 46189 973
rect 52295 959 52309 973
rect 52319 959 52333 973
rect 56759 959 56773 973
rect 56783 959 56797 973
rect 57215 959 57229 973
rect 57287 959 57301 973
rect 4175 935 4189 949
rect 5399 935 5413 949
rect 5423 935 5437 949
rect 10919 935 10933 949
rect 10943 935 10957 949
rect 20399 935 20413 949
rect 20495 935 20509 949
rect 21839 935 21853 949
rect 22943 935 22957 949
rect 23135 935 23149 949
rect 23159 935 23173 949
rect 41927 935 41941 949
rect 49943 935 49957 949
rect 49967 935 49981 949
rect 50447 935 50461 949
rect 56447 935 56461 949
rect 56471 935 56485 949
rect 57383 935 57397 949
rect 3959 911 3973 925
rect 53639 911 53653 925
rect 53687 911 53701 925
rect 55559 911 55573 925
rect 57407 911 57421 925
rect 3911 887 3925 901
rect 6047 887 6061 901
rect 6095 887 6109 901
rect 18023 887 18037 901
rect 32711 887 32725 901
rect 32735 887 32749 901
rect 48647 887 48661 901
rect 48671 887 48685 901
rect 57479 887 57493 901
rect 3383 863 3397 877
rect 3455 863 3469 877
rect 3551 863 3565 877
rect 8495 863 8509 877
rect 8543 863 8557 877
rect 10055 863 10069 877
rect 10103 863 10117 877
rect 12695 863 12709 877
rect 12743 863 12757 877
rect 13175 863 13189 877
rect 21047 863 21061 877
rect 21095 863 21109 877
rect 21215 863 21229 877
rect 25247 863 25261 877
rect 25271 863 25285 877
rect 28871 863 28885 877
rect 32831 863 32845 877
rect 32855 863 32869 877
rect 35591 863 35605 877
rect 35687 863 35701 877
rect 35783 863 35797 877
rect 35879 863 35893 877
rect 36599 863 36613 877
rect 39143 863 39157 877
rect 39167 863 39181 877
rect 40127 863 40141 877
rect 40151 863 40165 877
rect 49319 863 49333 877
rect 49343 863 49357 877
rect 51959 863 51973 877
rect 51983 863 51997 877
rect 53711 863 53725 877
rect 57599 863 57613 877
rect 3359 839 3373 853
rect 5999 839 6013 853
rect 8807 839 8821 853
rect 11951 839 11965 853
rect 11999 839 12013 853
rect 22415 839 22429 853
rect 22463 839 22477 853
rect 26063 839 26077 853
rect 37079 839 37093 853
rect 37175 839 37189 853
rect 39407 839 39421 853
rect 40199 839 40213 853
rect 48695 839 48709 853
rect 51119 839 51133 853
rect 53519 839 53533 853
rect 53543 839 53557 853
rect 57503 839 57517 853
rect 57695 839 57709 853
rect 3311 815 3325 829
rect 11183 815 11197 829
rect 11231 815 11245 829
rect 11447 815 11461 829
rect 11471 815 11485 829
rect 27311 815 27325 829
rect 27335 815 27349 829
rect 29159 815 29173 829
rect 38447 815 38461 829
rect 40967 815 40981 829
rect 40991 815 41005 829
rect 46439 815 46453 829
rect 46463 815 46477 829
rect 46919 815 46933 829
rect 46943 815 46957 829
rect 49199 815 49213 829
rect 56639 815 56653 829
rect 56663 815 56677 829
rect 57815 815 57829 829
rect 3191 791 3205 805
rect 3239 791 3253 805
rect 3263 791 3277 805
rect 4679 791 4693 805
rect 4799 791 4813 805
rect 8471 791 8485 805
rect 10991 791 11005 805
rect 11759 791 11773 805
rect 11783 791 11797 805
rect 32783 791 32797 805
rect 32831 791 32845 805
rect 42887 791 42901 805
rect 44087 791 44101 805
rect 52607 791 52621 805
rect 52727 791 52741 805
rect 57575 791 57589 805
rect 57599 791 57613 805
rect 57863 791 57877 805
rect 3167 767 3181 781
rect 5375 767 5389 781
rect 5399 767 5413 781
rect 9719 767 9733 781
rect 9767 767 9781 781
rect 18527 767 18541 781
rect 18551 767 18565 781
rect 29855 767 29869 781
rect 37799 767 37813 781
rect 37823 767 37837 781
rect 41111 767 41125 781
rect 43247 767 43261 781
rect 43271 767 43285 781
rect 45575 767 45589 781
rect 49823 767 49837 781
rect 49847 767 49861 781
rect 56663 767 56677 781
rect 56687 767 56701 781
rect 57887 767 57901 781
rect 3071 743 3085 757
rect 5255 743 5269 757
rect 5279 743 5293 757
rect 7727 743 7741 757
rect 7751 743 7765 757
rect 18239 743 18253 757
rect 19055 743 19069 757
rect 19079 743 19093 757
rect 23543 743 23557 757
rect 23567 743 23581 757
rect 26207 743 26221 757
rect 27791 743 27805 757
rect 28175 743 28189 757
rect 28295 743 28309 757
rect 28391 743 28405 757
rect 33911 743 33925 757
rect 33935 743 33949 757
rect 44255 743 44269 757
rect 52367 743 52381 757
rect 56855 743 56869 757
rect 56879 743 56893 757
rect 57935 743 57949 757
rect 3023 719 3037 733
rect 3335 719 3349 733
rect 3383 719 3397 733
rect 2999 695 3013 709
rect 8519 719 8533 733
rect 8615 719 8629 733
rect 14927 719 14941 733
rect 14951 719 14965 733
rect 21407 719 21421 733
rect 23279 719 23293 733
rect 27143 719 27157 733
rect 34703 719 34717 733
rect 36191 719 36205 733
rect 38567 719 38581 733
rect 41471 719 41485 733
rect 41495 719 41509 733
rect 45263 719 45277 733
rect 49031 719 49045 733
rect 49055 719 49069 733
rect 56615 719 56629 733
rect 56639 719 56653 733
rect 56735 719 56749 733
rect 56831 719 56845 733
rect 57719 719 57733 733
rect 3407 695 3421 709
rect 3431 695 3445 709
rect 4703 695 4717 709
rect 4823 695 4837 709
rect 5447 695 5461 709
rect 5471 695 5485 709
rect 7871 695 7885 709
rect 7943 695 7957 709
rect 11399 695 11413 709
rect 11447 695 11461 709
rect 13247 695 13261 709
rect 14447 695 14461 709
rect 14471 695 14485 709
rect 21527 695 21541 709
rect 21575 695 21589 709
rect 30215 695 30229 709
rect 32567 695 32581 709
rect 42143 695 42157 709
rect 44879 695 44893 709
rect 44903 695 44917 709
rect 46775 695 46789 709
rect 53759 695 53773 709
rect 53783 695 53797 709
rect 55511 695 55525 709
rect 55535 695 55549 709
rect 58007 695 58021 709
rect 58127 695 58141 709
rect 2975 671 2989 685
rect 3191 671 3205 685
rect 3215 671 3229 685
rect 9455 671 9469 685
rect 9503 671 9517 685
rect 12503 671 12517 685
rect 46607 671 46621 685
rect 50207 671 50221 685
rect 54167 671 54181 685
rect 56591 671 56605 685
rect 57743 671 57757 685
rect 58223 671 58237 685
rect 2927 647 2941 661
rect 7175 647 7189 661
rect 7199 647 7213 661
rect 11255 647 11269 661
rect 11351 647 11365 661
rect 19079 647 19093 661
rect 19175 647 19189 661
rect 26399 647 26413 661
rect 26447 647 26461 661
rect 37943 647 37957 661
rect 37967 647 37981 661
rect 38807 647 38821 661
rect 40103 647 40117 661
rect 45503 647 45517 661
rect 47903 647 47917 661
rect 49295 647 49309 661
rect 54839 647 54853 661
rect 57431 647 57445 661
rect 58055 647 58069 661
rect 58319 647 58333 661
rect 2903 623 2917 637
rect 3167 623 3181 637
rect 3191 623 3205 637
rect 3551 623 3565 637
rect 3575 623 3589 637
rect 5639 623 5653 637
rect 5663 623 5677 637
rect 24359 623 24373 637
rect 24383 623 24397 637
rect 25103 623 25117 637
rect 26543 623 26557 637
rect 36839 623 36853 637
rect 40823 623 40837 637
rect 52703 623 52717 637
rect 57911 623 57925 637
rect 57935 623 57949 637
rect 58391 623 58405 637
rect 2879 599 2893 613
rect 2975 599 2989 613
rect 3047 599 3061 613
rect 5351 599 5365 613
rect 5375 599 5389 613
rect 5951 599 5965 613
rect 5975 599 5989 613
rect 8447 599 8461 613
rect 10607 599 10621 613
rect 10679 599 10693 613
rect 21551 599 21565 613
rect 21623 599 21637 613
rect 23399 599 23413 613
rect 23423 599 23437 613
rect 26375 599 26389 613
rect 26399 599 26413 613
rect 33263 599 33277 613
rect 33287 599 33301 613
rect 37319 599 37333 613
rect 37343 599 37357 613
rect 45527 599 45541 613
rect 45551 599 45565 613
rect 50807 599 50821 613
rect 50831 599 50845 613
rect 57359 599 57373 613
rect 57407 599 57421 613
rect 57455 599 57469 613
rect 57479 599 57493 613
rect 58439 599 58453 613
rect 2855 575 2869 589
rect 2927 575 2941 589
rect 2951 575 2965 589
rect 4775 575 4789 589
rect 4871 575 4885 589
rect 5783 575 5797 589
rect 5855 575 5869 589
rect 8087 575 8101 589
rect 8111 575 8125 589
rect 8183 575 8197 589
rect 8231 575 8245 589
rect 10271 575 10285 589
rect 10319 575 10333 589
rect 12983 575 12997 589
rect 13031 575 13045 589
rect 19151 575 19165 589
rect 19199 575 19213 589
rect 27215 575 27229 589
rect 27239 575 27253 589
rect 32783 575 32797 589
rect 32807 575 32821 589
rect 34367 575 34381 589
rect 38975 575 38989 589
rect 39383 575 39397 589
rect 45191 575 45205 589
rect 45215 575 45229 589
rect 54263 575 54277 589
rect 54287 575 54301 589
rect 57071 575 57085 589
rect 57095 575 57109 589
rect 58175 575 58189 589
rect 58463 575 58477 589
rect 58559 575 58573 589
rect 5207 551 5221 565
rect 5255 551 5269 565
rect 6383 551 6397 565
rect 6407 551 6421 565
rect 13967 551 13981 565
rect 32615 551 32629 565
rect 32639 551 32653 565
rect 48047 551 48061 565
rect 52775 551 52789 565
rect 52799 551 52813 565
rect 53831 551 53845 565
rect 55679 551 55693 565
rect 58655 551 58669 565
rect 2831 527 2845 541
rect 4799 527 4813 541
rect 4895 527 4909 541
rect 12791 527 12805 541
rect 12815 527 12829 541
rect 20807 527 20821 541
rect 20831 527 20845 541
rect 23207 527 23221 541
rect 23591 527 23605 541
rect 23663 527 23677 541
rect 23687 527 23701 541
rect 23807 527 23821 541
rect 28487 527 28501 541
rect 28583 527 28597 541
rect 28679 527 28693 541
rect 28967 527 28981 541
rect 29279 527 29293 541
rect 29303 527 29317 541
rect 33767 527 33781 541
rect 42191 527 42205 541
rect 42215 527 42229 541
rect 47351 527 47365 541
rect 47375 527 47389 541
rect 47399 527 47413 541
rect 52175 527 52189 541
rect 52199 527 52213 541
rect 55703 527 55717 541
rect 57047 527 57061 541
rect 57407 527 57421 541
rect 57959 527 57973 541
rect 58151 527 58165 541
rect 58487 527 58501 541
rect 58727 527 58741 541
rect 4751 503 4765 517
rect 4775 503 4789 517
rect 10175 503 10189 517
rect 10199 503 10213 517
rect 12167 503 12181 517
rect 12191 503 12205 517
rect 23111 503 23125 517
rect 23135 503 23149 517
rect 54959 503 54973 517
rect 54983 503 54997 517
rect 55727 503 55741 517
rect 55751 503 55765 517
rect 57023 503 57037 517
rect 58919 3239 58933 3253
rect 59039 3239 59053 3253
rect 59639 3239 59653 3253
rect 59759 3239 59773 3253
rect 2759 479 2773 493
rect 2783 479 2797 493
rect 2807 479 2821 493
rect 5831 479 5845 493
rect 5879 479 5893 493
rect 23471 479 23485 493
rect 32399 479 32413 493
rect 32423 479 32437 493
rect 39743 479 39757 493
rect 39767 479 39781 493
rect 43919 479 43933 493
rect 53351 479 53365 493
rect 53375 479 53389 493
rect 54071 479 54085 493
rect 54095 479 54109 493
rect 57263 479 57277 493
rect 57287 479 57301 493
rect 58751 479 58765 493
rect 58775 479 58789 493
rect 58799 479 58813 493
rect 2735 455 2749 469
rect 8015 455 8029 469
rect 8039 455 8053 469
rect 21071 455 21085 469
rect 21119 455 21133 469
rect 29063 455 29077 469
rect 44111 455 44125 469
rect 45695 455 45709 469
rect 46271 455 46285 469
rect 51095 455 51109 469
rect 53399 455 53413 469
rect 54527 455 54541 469
rect 54551 455 54565 469
rect 56807 455 56821 469
rect 58823 455 58837 469
rect 2711 431 2725 445
rect 2855 431 2869 445
rect 2903 431 2917 445
rect 2663 407 2677 421
rect 5231 431 5245 445
rect 5303 431 5317 445
rect 5591 431 5605 445
rect 5639 431 5653 445
rect 18863 431 18877 445
rect 18887 431 18901 445
rect 33215 431 33229 445
rect 39527 431 39541 445
rect 39551 431 39565 445
rect 42383 431 42397 445
rect 45431 431 45445 445
rect 45455 431 45469 445
rect 45839 431 45853 445
rect 45863 431 45877 445
rect 52487 431 52501 445
rect 54863 431 54877 445
rect 54887 431 54901 445
rect 58415 431 58429 445
rect 58439 431 58453 445
rect 58871 431 58885 445
rect 58919 431 58933 445
rect 2927 407 2941 421
rect 2975 407 2989 421
rect 4943 407 4957 421
rect 5015 407 5029 421
rect 6071 407 6085 421
rect 6119 407 6133 421
rect 6215 407 6229 421
rect 6431 407 6445 421
rect 7775 407 7789 421
rect 8207 407 8221 421
rect 8255 407 8269 421
rect 12047 407 12061 421
rect 21983 407 21997 421
rect 36335 407 36349 421
rect 36359 407 36373 421
rect 36383 407 36397 421
rect 36719 407 36733 421
rect 36815 407 36829 421
rect 38231 407 38245 421
rect 38687 407 38701 421
rect 42671 407 42685 421
rect 42695 407 42709 421
rect 50231 407 50245 421
rect 50255 407 50269 421
rect 51335 407 51349 421
rect 53087 407 53101 421
rect 53279 407 53293 421
rect 54935 407 54949 421
rect 58943 407 58957 421
rect 59639 3047 59653 3061
rect 59759 3047 59773 3061
rect 2639 383 2653 397
rect 9095 383 9109 397
rect 9815 383 9829 397
rect 9863 383 9877 397
rect 10007 383 10021 397
rect 10055 383 10069 397
rect 32519 383 32533 397
rect 32543 383 32557 397
rect 37439 383 37453 397
rect 37463 383 37477 397
rect 44687 383 44701 397
rect 44711 383 44725 397
rect 55607 383 55621 397
rect 55631 383 55645 397
rect 58079 383 58093 397
rect 58247 383 58261 397
rect 58799 383 58813 397
rect 58823 383 58837 397
rect 58847 383 58861 397
rect 58871 383 58885 397
rect 58991 383 59005 397
rect 59039 383 59053 397
rect 7967 359 7981 373
rect 8015 359 8029 373
rect 8135 359 8149 373
rect 8183 359 8197 373
rect 10079 359 10093 373
rect 10127 359 10141 373
rect 11519 359 11533 373
rect 11543 359 11557 373
rect 40511 359 40525 373
rect 53927 359 53941 373
rect 57671 359 57685 373
rect 57695 359 57709 373
rect 57839 359 57853 373
rect 57863 359 57877 373
rect 58631 359 58645 373
rect 58655 359 58669 373
rect 2615 335 2629 349
rect 2639 335 2653 349
rect 2567 311 2581 325
rect 5783 335 5797 349
rect 9863 335 9877 349
rect 9911 335 9925 349
rect 21455 335 21469 349
rect 21479 335 21493 349
rect 26783 335 26797 349
rect 26807 335 26821 349
rect 28199 335 28213 349
rect 47327 335 47341 349
rect 49487 335 49501 349
rect 56951 335 56965 349
rect 56975 335 56989 349
rect 58967 335 58981 349
rect 58991 335 59005 349
rect 59039 335 59053 349
rect 59639 2999 59653 3013
rect 59759 2999 59773 3013
rect 59639 2807 59653 2821
rect 59759 2807 59773 2821
rect 59639 2759 59653 2773
rect 59759 2759 59773 2773
rect 59519 2327 59533 2341
rect 59639 2327 59653 2341
rect 59759 2327 59773 2341
rect 59879 2327 59893 2341
rect 59519 2279 59533 2293
rect 59639 2279 59653 2293
rect 59759 2279 59773 2293
rect 59879 2279 59893 2293
rect 59399 2087 59413 2101
rect 59519 2087 59533 2101
rect 59639 2087 59653 2101
rect 59759 2087 59773 2101
rect 59879 2087 59893 2101
rect 59111 335 59125 349
rect 59159 335 59173 349
rect 2687 311 2701 325
rect 2711 311 2725 325
rect 2543 287 2557 301
rect 4175 311 4189 325
rect 4199 311 4213 325
rect 5111 311 5125 325
rect 5183 311 5197 325
rect 8687 311 8701 325
rect 8711 311 8725 325
rect 9671 311 9685 325
rect 9695 311 9709 325
rect 13439 311 13453 325
rect 13463 311 13477 325
rect 14951 311 14965 325
rect 14975 311 14989 325
rect 15623 311 15637 325
rect 15647 311 15661 325
rect 24119 311 24133 325
rect 24143 311 24157 325
rect 35903 311 35917 325
rect 46391 311 46405 325
rect 52535 311 52549 325
rect 52559 311 52573 325
rect 57791 311 57805 325
rect 57815 311 57829 325
rect 2855 287 2869 301
rect 2903 287 2917 301
rect 20975 287 20989 301
rect 21023 287 21037 301
rect 38495 287 38509 301
rect 38519 287 38533 301
rect 50279 287 50293 301
rect 54383 287 54397 301
rect 54407 287 54421 301
rect 58295 287 58309 301
rect 58319 287 58333 301
rect 58607 287 58621 301
rect 59159 287 59173 301
rect 59399 2039 59413 2053
rect 59519 2039 59533 2053
rect 59639 2039 59653 2053
rect 59759 2039 59773 2053
rect 59879 2039 59893 2053
rect 59231 287 59245 301
rect 59279 287 59293 301
rect 2519 263 2533 277
rect 2999 263 3013 277
rect 3095 263 3109 277
rect 4583 263 4597 277
rect 4607 263 4621 277
rect 10439 263 10453 277
rect 10463 263 10477 277
rect 10631 263 10645 277
rect 10727 263 10741 277
rect 11543 263 11557 277
rect 11567 263 11581 277
rect 38711 263 38725 277
rect 41351 263 41365 277
rect 48983 263 48997 277
rect 49775 263 49789 277
rect 51527 263 51541 277
rect 54095 263 54109 277
rect 54119 263 54133 277
rect 55823 263 55837 277
rect 55847 263 55861 277
rect 58103 263 58117 277
rect 58127 263 58141 277
rect 59303 263 59317 277
rect 2375 239 2389 253
rect 2759 239 2773 253
rect 2999 239 3013 253
rect 5519 239 5533 253
rect 5543 239 5557 253
rect 5687 239 5701 253
rect 5711 239 5725 253
rect 13367 239 13381 253
rect 14639 239 14653 253
rect 14663 239 14677 253
rect 23015 239 23029 253
rect 23063 239 23077 253
rect 46511 239 46525 253
rect 47639 239 47653 253
rect 48287 239 48301 253
rect 48503 239 48517 253
rect 52247 239 52261 253
rect 57167 239 57181 253
rect 57215 239 57229 253
rect 57335 239 57349 253
rect 57383 239 57397 253
rect 59351 239 59365 253
rect 59399 239 59413 253
rect 1967 191 1981 205
rect 2567 215 2581 229
rect 2591 215 2605 229
rect 5495 215 5509 229
rect 5519 215 5533 229
rect 7583 215 7597 229
rect 7607 215 7621 229
rect 35999 215 36013 229
rect 39311 215 39325 229
rect 43223 215 43237 229
rect 46199 215 46213 229
rect 47615 215 47629 229
rect 48191 215 48205 229
rect 48311 215 48325 229
rect 48527 215 48541 229
rect 54479 215 54493 229
rect 54575 215 54589 229
rect 57647 215 57661 229
rect 58367 215 58381 229
rect 58391 215 58405 229
rect 59087 215 59101 229
rect 59111 215 59125 229
rect 59423 215 59437 229
rect 2351 191 2365 205
rect 2543 191 2557 205
rect 2567 191 2581 205
rect 2687 191 2701 205
rect 2711 191 2725 205
rect 14231 191 14245 205
rect 14255 191 14269 205
rect 14375 191 14389 205
rect 14783 191 14797 205
rect 14855 191 14869 205
rect 14879 191 14893 205
rect 21767 191 21781 205
rect 23951 191 23965 205
rect 24791 191 24805 205
rect 31295 191 31309 205
rect 38015 191 38029 205
rect 46655 191 46669 205
rect 46679 191 46693 205
rect 48551 191 48565 205
rect 48575 191 48589 205
rect 48743 191 48757 205
rect 48767 191 48781 205
rect 48815 191 48829 205
rect 50999 191 51013 205
rect 52127 191 52141 205
rect 53879 191 53893 205
rect 53903 191 53917 205
rect 54455 191 54469 205
rect 55223 191 55237 205
rect 57311 191 57325 205
rect 57335 191 57349 205
rect 57623 191 57637 205
rect 58343 191 58357 205
rect 58703 191 58717 205
rect 58775 191 58789 205
rect 59327 191 59341 205
rect 59351 191 59365 205
rect 59471 191 59485 205
rect 59519 191 59533 205
rect 1751 167 1765 181
rect 3359 167 3373 181
rect 3383 167 3397 181
rect 4991 167 5005 181
rect 5039 167 5053 181
rect 8663 167 8677 181
rect 8687 167 8701 181
rect 8975 167 8989 181
rect 8999 167 9013 181
rect 11279 167 11293 181
rect 11399 167 11413 181
rect 11423 167 11437 181
rect 11495 167 11509 181
rect 15023 167 15037 181
rect 15071 167 15085 181
rect 18863 167 18877 181
rect 20711 167 20725 181
rect 20807 167 20821 181
rect 21287 167 21301 181
rect 21311 167 21325 181
rect 28511 167 28525 181
rect 42527 167 42541 181
rect 45479 167 45493 181
rect 46415 167 46429 181
rect 53207 167 53221 181
rect 53231 167 53245 181
rect 53975 167 53989 181
rect 53999 167 54013 181
rect 55919 167 55933 181
rect 55943 167 55957 181
rect 57239 167 57253 181
rect 59207 167 59221 181
rect 59231 167 59245 181
rect 59543 167 59557 181
rect 1703 143 1717 157
rect 3071 143 3085 157
rect 3119 143 3133 157
rect 3263 143 3277 157
rect 3287 143 3301 157
rect 3911 143 3925 157
rect 3935 143 3949 157
rect 6911 143 6925 157
rect 6935 143 6949 157
rect 44759 143 44773 157
rect 45023 143 45037 157
rect 54599 143 54613 157
rect 55247 143 55261 157
rect 55319 143 55333 157
rect 57143 143 57157 157
rect 57191 143 57205 157
rect 59591 143 59605 157
rect 59639 143 59653 157
rect 1127 95 1141 109
rect 1751 119 1765 133
rect 1775 119 1789 133
rect 1967 119 1981 133
rect 1991 119 2005 133
rect 2519 119 2533 133
rect 2543 119 2557 133
rect 2879 119 2893 133
rect 3071 119 3085 133
rect 4847 119 4861 133
rect 4919 119 4933 133
rect 10295 119 10309 133
rect 10343 119 10357 133
rect 13007 119 13021 133
rect 13055 119 13069 133
rect 21191 119 21205 133
rect 24407 119 24421 133
rect 24431 119 24445 133
rect 28895 119 28909 133
rect 29087 119 29101 133
rect 34103 119 34117 133
rect 34127 119 34141 133
rect 36071 119 36085 133
rect 38831 119 38845 133
rect 38855 119 38869 133
rect 52655 119 52669 133
rect 52679 119 52693 133
rect 54047 119 54061 133
rect 54071 119 54085 133
rect 57527 119 57541 133
rect 57863 119 57877 133
rect 57887 119 57901 133
rect 59447 119 59461 133
rect 59471 119 59485 133
rect 59663 119 59677 133
rect 1367 95 1381 109
rect 1703 95 1717 109
rect 1727 95 1741 109
rect 3959 95 3973 109
rect 3983 95 3997 109
rect 4727 95 4741 109
rect 4751 95 4765 109
rect 5495 95 5509 109
rect 6167 95 6181 109
rect 6191 95 6205 109
rect 14543 95 14557 109
rect 14567 95 14581 109
rect 20903 95 20917 109
rect 46343 95 46357 109
rect 46367 95 46381 109
rect 51359 95 51373 109
rect 51383 95 51397 109
rect 54287 95 54301 109
rect 54311 95 54325 109
rect 55439 95 55453 109
rect 57119 95 57133 109
rect 58679 95 58693 109
rect 58727 95 58741 109
rect 59711 95 59725 109
rect 59759 95 59773 109
rect 743 71 757 85
rect 4535 71 4549 85
rect 4559 71 4573 85
rect 18743 71 18757 85
rect 18767 71 18781 85
rect 25175 71 25189 85
rect 26303 71 26317 85
rect 27455 71 27469 85
rect 30839 71 30853 85
rect 32063 71 32077 85
rect 33311 71 33325 85
rect 33743 71 33757 85
rect 33839 71 33853 85
rect 34247 71 34261 85
rect 38639 71 38653 85
rect 38663 71 38677 85
rect 40751 71 40765 85
rect 40775 71 40789 85
rect 52079 71 52093 85
rect 52103 71 52117 85
rect 56903 71 56917 85
rect 58199 71 58213 85
rect 58223 71 58237 85
rect 58271 71 58285 85
rect 58919 71 58933 85
rect 58943 71 58957 85
rect 59279 71 59293 85
rect 59303 71 59317 85
rect 59639 71 59653 85
rect 59663 71 59677 85
rect 59807 71 59821 85
rect 59879 71 59893 85
rect 2375 47 2389 61
rect 2399 47 2413 61
rect 2615 47 2629 61
rect 2639 47 2653 61
rect 3023 47 3037 61
rect 3143 47 3157 61
rect 23519 47 23533 61
rect 23543 47 23557 61
rect 24143 47 24157 61
rect 24167 47 24181 61
rect 26783 47 26797 61
rect 27983 47 27997 61
rect 28007 47 28021 61
rect 42047 47 42061 61
rect 49679 47 49693 61
rect 53063 47 53077 61
rect 58535 47 58549 61
rect 58559 47 58573 61
rect 58583 47 58597 61
rect 59399 47 59413 61
rect 59423 47 59437 61
rect 59567 47 59581 61
rect 59591 47 59605 61
rect 1127 23 1141 37
rect 2735 23 2749 37
rect 12095 23 12109 37
rect 12119 23 12133 37
rect 12143 23 12157 37
rect 20447 23 20461 37
rect 20471 23 20485 37
rect 20495 23 20509 37
rect 59519 23 59533 37
rect 59543 23 59557 37
rect 59711 23 59725 37
rect 59879 23 59893 37
rect 119 -1 133 13
rect 527 -1 541 13
rect 1151 -1 1165 13
rect 2759 -1 2773 13
rect 12119 -1 12133 13
rect 12143 -1 12157 13
rect 12167 -1 12181 13
rect 20471 -1 20485 13
rect 20495 -1 20509 13
rect 20519 -1 20533 13
rect 28991 -1 29005 13
rect 34271 -1 34285 13
rect 37271 -1 37285 13
rect 49583 -1 49597 13
rect 54719 -1 54733 13
rect 55031 -1 55045 13
rect 55799 -1 55813 13
rect 55895 -1 55909 13
rect 57983 -1 57997 13
rect 59519 -1 59533 13
rect 59687 -1 59701 13
rect 59879 -1 59893 13
rect 59927 -1 59941 13
<< metal2 >>
rect 32256 31549 32268 31583
rect 32256 30757 32268 30791
rect 32256 29989 32268 30023
rect 32280 29989 32292 30023
rect 32256 29245 32268 29279
rect 32280 29245 32292 29279
rect 32304 29245 32316 29279
rect 32256 28285 32268 28319
rect 32280 28285 32292 28319
rect 32304 28285 32316 28319
rect 32328 28285 32340 28319
rect 32256 27541 32268 27575
rect 32280 27541 32292 27575
rect 32304 27541 32316 27575
rect 32328 27541 32340 27575
rect 32352 27541 32364 27575
rect 32256 27373 32268 27407
rect 32280 27373 32292 27407
rect 32304 27373 32316 27407
rect 32328 27373 32340 27407
rect 32352 27373 32364 27407
rect 32376 27373 32388 27407
rect 32256 17965 32268 17999
rect 32280 17965 32292 17999
rect 32304 17965 32316 17999
rect 32328 17965 32340 17999
rect 32352 17965 32364 17999
rect 32376 17965 32388 17999
rect 32400 17965 32412 17999
rect 32256 17773 32268 17807
rect 32280 17773 32292 17807
rect 32304 17773 32316 17807
rect 32328 17773 32340 17807
rect 32352 17773 32364 17807
rect 32376 17773 32388 17807
rect 32400 17773 32412 17807
rect 32424 17773 32436 17807
rect 32256 17533 32268 17567
rect 32280 17533 32292 17567
rect 32304 17533 32316 17567
rect 32328 17533 32340 17567
rect 32352 17533 32364 17567
rect 32376 17533 32388 17567
rect 32400 17533 32412 17567
rect 32424 17533 32436 17567
rect 32256 17293 32268 17327
rect 32280 17293 32292 17327
rect 32304 17293 32316 17327
rect 32328 17293 32340 17327
rect 32352 17293 32364 17327
rect 32376 17293 32388 17327
rect 32400 17293 32412 17327
rect 32424 17293 32436 17327
rect 32448 17293 32460 17327
rect 32856 17173 32868 17207
rect 32256 16813 32268 16847
rect 32280 16813 32292 16847
rect 32304 16813 32316 16847
rect 32328 16813 32340 16847
rect 32352 16813 32364 16847
rect 32376 16813 32388 16847
rect 32400 16813 32412 16847
rect 32424 16813 32436 16847
rect 32448 16813 32460 16847
rect 32472 16813 32484 16847
rect 32496 16813 32508 16847
rect 32256 16573 32268 16607
rect 32280 16573 32292 16607
rect 32304 16573 32316 16607
rect 32328 16573 32340 16607
rect 32352 16573 32364 16607
rect 32376 16573 32388 16607
rect 32400 16573 32412 16607
rect 32424 16573 32436 16607
rect 32448 16573 32460 16607
rect 32472 16573 32484 16607
rect 32496 16573 32508 16607
rect 32520 16573 32532 16607
rect 32256 16333 32268 16367
rect 32280 16333 32292 16367
rect 32304 16333 32316 16367
rect 32328 16333 32340 16367
rect 32352 16333 32364 16367
rect 32376 16333 32388 16367
rect 32400 16333 32412 16367
rect 32424 16333 32436 16367
rect 32448 16333 32460 16367
rect 32472 16333 32484 16367
rect 32520 16357 32532 16391
rect 32544 16357 32556 16391
rect 32256 16093 32268 16127
rect 32280 16093 32292 16127
rect 32304 16093 32316 16127
rect 32328 16093 32340 16127
rect 32352 16093 32364 16127
rect 32400 16117 32412 16151
rect 32424 16117 32436 16151
rect 32448 16117 32460 16151
rect 32472 16117 32484 16151
rect 32496 16117 32508 16151
rect 32520 16117 32532 16151
rect 32544 16117 32556 16151
rect 32568 16117 32580 16151
rect 32856 15493 32868 15527
rect 32904 15493 32916 15527
rect 32928 15493 32940 15527
rect 32952 15493 32964 15527
rect 32976 15493 32988 15527
rect 33000 15493 33012 15527
rect 33024 15493 33036 15527
rect 32760 14293 32772 14327
rect 32856 14293 32868 14327
rect 32904 14293 32916 14327
rect 32928 14293 32940 14327
rect 32952 14293 32964 14327
rect 32976 14293 32988 14327
rect 33000 14293 33012 14327
rect 33024 14293 33036 14327
rect 33048 14293 33060 14327
rect 33072 14293 33084 14327
rect 33096 14293 33108 14327
rect 33120 14293 33132 14327
rect 32856 14053 32868 14087
rect 32904 14053 32916 14087
rect 32928 14053 32940 14087
rect 32952 14053 32964 14087
rect 32976 14053 32988 14087
rect 33000 14053 33012 14087
rect 33024 14053 33036 14087
rect 33048 14053 33060 14087
rect 33072 14053 33084 14087
rect 33096 14053 33108 14087
rect 33120 14053 33132 14087
rect 32856 13573 32868 13607
rect 32904 13573 32916 13607
rect 32928 13573 32940 13607
rect 32952 13573 32964 13607
rect 32976 13573 32988 13607
rect 33000 13573 33012 13607
rect 33024 13573 33036 13607
rect 33048 13573 33060 13607
rect 33072 13573 33084 13607
rect 33096 13573 33108 13607
rect 33120 13573 33132 13607
rect 33144 13573 33156 13607
rect 41160 12853 41172 12887
rect 41160 12613 41172 12647
rect 41160 12373 41172 12407
rect 32808 12133 32820 12167
rect 32832 12133 32844 12167
rect 32856 12133 32868 12167
rect 32904 12133 32916 12167
rect 32928 12133 32940 12167
rect 32952 12133 32964 12167
rect 32976 12133 32988 12167
rect 33000 12133 33012 12167
rect 33024 12133 33036 12167
rect 33048 12133 33060 12167
rect 33072 12133 33084 12167
rect 33096 12133 33108 12167
rect 33120 12133 33132 12167
rect 33144 12133 33156 12167
rect 33168 12133 33180 12167
rect 33192 12133 33204 12167
rect 33240 12133 33252 12167
rect 33264 12133 33276 12167
rect 41160 12133 41172 12167
rect 41160 11893 41172 11927
rect 41160 11653 41172 11687
rect 32256 9829 32268 9863
rect 32280 9829 32292 9863
rect 32304 9829 32316 9863
rect 32328 9829 32340 9863
rect 32352 9829 32364 9863
rect 32376 9829 32388 9863
rect 32400 9829 32412 9863
rect 32424 9829 32436 9863
rect 32448 9829 32460 9863
rect 32472 9829 32484 9863
rect 32496 9829 32508 9863
rect 32544 9853 32556 9887
rect 32568 9853 32580 9887
rect 32592 9853 32604 9887
rect 32616 9157 32628 9191
rect 32256 9085 32268 9119
rect 32280 9085 32292 9119
rect 32304 9085 32316 9119
rect 32328 9085 32340 9119
rect 32352 9085 32364 9119
rect 32376 9085 32388 9119
rect 32400 9085 32412 9119
rect 32448 9109 32460 9143
rect 32472 9109 32484 9143
rect 32496 9109 32508 9143
rect 32520 9109 32532 9143
rect 32544 9109 32556 9143
rect 33240 8773 33252 8807
rect 33264 8773 33276 8807
rect 33288 8773 33300 8807
rect 33312 8773 33324 8807
rect 41160 8773 41172 8807
rect 32688 8701 32700 8735
rect 32712 8701 32724 8735
rect 32736 8701 32748 8735
rect 32760 8701 32772 8735
rect 32784 8701 32796 8735
rect 32808 8701 32820 8735
rect 32832 8701 32844 8735
rect 32856 8701 32868 8735
rect 31800 8173 31812 8207
rect 31824 8173 31836 8255
rect 31848 8173 31860 8303
rect 31872 8173 31884 8327
rect 31896 8173 31908 8351
rect 31920 8173 31932 8375
rect 31944 8173 31956 8399
rect 31968 8173 31980 8423
rect 31992 8173 32004 8447
rect 32016 8173 32028 8471
rect 32040 8173 32052 8495
rect 32064 8173 32076 8519
rect 32088 8173 32100 8543
rect 32112 8173 32124 8567
rect 32136 8173 32148 8591
rect 32160 8173 32172 8615
rect 32256 8173 32268 8687
rect 32280 8173 32292 8687
rect 32304 8173 32316 8687
rect 32328 8269 32340 8687
rect 32352 8581 32364 8687
rect 32328 8173 32340 8207
rect 32352 8173 32364 8231
rect 32376 8173 32388 8687
rect 32400 8173 32412 8687
rect 32424 8173 32436 8687
rect 32448 8173 32460 8687
rect 32472 8173 32484 8687
rect 32496 8245 32508 8687
rect 32520 8269 32532 8687
rect 32544 8317 32556 8687
rect 32568 8389 32580 8687
rect 32592 8533 32604 8687
rect 32616 8581 32628 8687
rect 32664 8581 32676 8615
rect 32688 8581 32700 8615
rect 32616 8389 32628 8519
rect 32664 8389 32676 8519
rect 32592 8317 32604 8375
rect 32568 8269 32580 8303
rect 32520 8173 32532 8207
rect 32544 8173 32556 8207
rect 32568 8173 32580 8231
rect 32616 8149 32628 8303
rect 32640 8269 32652 8375
rect 32640 8149 32652 8231
rect 32664 8149 32676 8255
rect 32688 8149 32700 8519
rect 32712 8149 32724 8615
rect 32736 8149 32748 8615
rect 32760 8149 32772 8615
rect 32784 8149 32796 8615
rect 32808 8149 32820 8615
rect 32832 8149 32844 8615
rect 32856 8221 32868 8615
rect 32880 8125 32892 8615
rect 32904 8317 32916 8615
rect 32928 8509 32940 8615
rect 32952 8389 32964 8615
rect 32928 8317 32940 8375
rect 32976 8317 32988 8615
rect 33000 8317 33012 8615
rect 33024 8437 33036 8615
rect 33048 8389 33060 8615
rect 33072 8581 33084 8615
rect 33096 8581 33108 8615
rect 33120 8581 33132 8615
rect 33144 8581 33156 8615
rect 33072 8389 33084 8495
rect 33120 8437 33132 8495
rect 33144 8437 33156 8495
rect 33168 8437 33180 8495
rect 33192 8437 33204 8495
rect 33216 8437 33228 8567
rect 33240 8461 33252 8495
rect 33024 8317 33036 8375
rect 33216 8317 33228 8351
rect 32952 8221 32964 8279
rect 32904 8173 32916 8207
rect 31776 6373 31788 6407
rect 31800 6373 31812 6407
rect 31824 6373 31836 6407
rect 31848 6373 31860 6407
rect 31872 6373 31884 6407
rect 31896 6373 31908 6407
rect 31920 6373 31932 6407
rect 31944 6373 31956 6407
rect 31968 6373 31980 6407
rect 31992 6373 32004 6407
rect 32016 6373 32028 6407
rect 32040 6373 32052 6407
rect 32064 6373 32076 6407
rect 32088 6373 32100 6407
rect 32112 6373 32124 6407
rect 32136 6373 32148 6407
rect 32160 6373 32172 6407
rect 32256 6373 32268 6407
rect 32280 6373 32292 6407
rect 32304 6373 32316 6407
rect 32328 6373 32340 6407
rect 32352 6373 32364 6407
rect 32376 6373 32388 6407
rect 32400 6373 32412 6407
rect 32424 6373 32436 6407
rect 32448 6373 32460 6407
rect 32472 6373 32484 6407
rect 32520 6373 32532 6407
rect 32544 6373 32556 6407
rect 32568 6373 32580 6407
rect 32592 6373 32604 6407
rect 32616 6373 32628 6407
rect 32640 6373 32652 6407
rect 32664 6373 32676 6407
rect 32688 6373 32700 6407
rect 32712 6373 32724 6407
rect 32736 6373 32748 6407
rect 32760 6373 32772 6407
rect 32784 6373 32796 6407
rect 32808 6373 32820 6407
rect 32832 6373 32844 6407
rect 32856 6373 32868 6407
rect 32880 6373 32892 6407
rect 32904 6373 32916 6407
rect 33216 6373 33228 6407
rect 41160 6373 41172 6407
rect 31752 6133 31764 6167
rect 31776 6133 31788 6167
rect 31800 6133 31812 6167
rect 31824 6133 31836 6167
rect 31848 6133 31860 6167
rect 31872 6133 31884 6167
rect 31896 6133 31908 6167
rect 31920 6133 31932 6167
rect 31944 6133 31956 6167
rect 31968 6133 31980 6167
rect 31992 6133 32004 6167
rect 32016 6133 32028 6167
rect 32040 6133 32052 6167
rect 32064 6133 32076 6167
rect 32088 6133 32100 6167
rect 32112 6133 32124 6167
rect 32136 6133 32148 6167
rect 32160 6133 32172 6167
rect 32256 6133 32268 6167
rect 32280 6133 32292 6167
rect 32304 6133 32316 6167
rect 32328 6133 32340 6167
rect 32352 6133 32364 6167
rect 32376 6133 32388 6167
rect 32400 6133 32412 6167
rect 32424 6133 32436 6167
rect 32448 6133 32460 6167
rect 32472 6133 32484 6167
rect 32520 6133 32532 6167
rect 32544 6133 32556 6167
rect 32568 6133 32580 6167
rect 32592 6133 32604 6167
rect 32616 6133 32628 6167
rect 32640 6133 32652 6167
rect 32664 6133 32676 6167
rect 32688 6133 32700 6167
rect 32712 6133 32724 6167
rect 32736 6133 32748 6167
rect 32760 6133 32772 6167
rect 32784 6133 32796 6167
rect 32808 6133 32820 6167
rect 32832 6133 32844 6167
rect 32856 6133 32868 6167
rect 32880 6133 32892 6167
rect 32904 6133 32916 6167
rect 33216 6133 33228 6167
rect 41160 6133 41172 6167
rect 41160 5893 41172 5927
rect 41160 5653 41172 5687
rect 31728 5413 31740 5447
rect 31752 5413 31764 5447
rect 31776 5413 31788 5447
rect 31800 5413 31812 5447
rect 31824 5413 31836 5447
rect 31848 5413 31860 5447
rect 31872 5413 31884 5447
rect 31896 5413 31908 5447
rect 31920 5413 31932 5447
rect 31944 5413 31956 5447
rect 31968 5413 31980 5447
rect 31992 5413 32004 5447
rect 32016 5413 32028 5447
rect 32040 5413 32052 5447
rect 32064 5413 32076 5447
rect 32088 5413 32100 5447
rect 32112 5413 32124 5447
rect 32136 5413 32148 5447
rect 32160 5413 32172 5447
rect 32256 5413 32268 5447
rect 32280 5413 32292 5447
rect 32304 5413 32316 5447
rect 32328 5413 32340 5447
rect 32352 5413 32364 5447
rect 32376 5413 32388 5447
rect 32400 5413 32412 5447
rect 32424 5413 32436 5447
rect 32448 5413 32460 5447
rect 32472 5413 32484 5447
rect 32520 5413 32532 5447
rect 32544 5413 32556 5447
rect 32568 5413 32580 5447
rect 32592 5413 32604 5447
rect 32616 5413 32628 5447
rect 32640 5413 32652 5447
rect 32664 5413 32676 5447
rect 32688 5413 32700 5447
rect 32712 5413 32724 5447
rect 32736 5413 32748 5447
rect 32760 5413 32772 5447
rect 32784 5413 32796 5447
rect 32808 5413 32820 5447
rect 32832 5413 32844 5447
rect 32856 5413 32868 5447
rect 32880 5413 32892 5447
rect 32904 5413 32916 5447
rect 33216 5413 33228 5447
rect 33336 5413 33348 5447
rect 33384 5413 33396 5447
rect 41160 5413 41172 5447
rect 2640 349 2652 383
rect 1704 109 1716 143
rect 1752 133 1764 167
rect 1968 133 1980 191
rect 120 -24 132 -1
rect 528 -24 540 -1
rect 744 -24 756 71
rect 1128 37 1140 95
rect 1152 -24 1164 -1
rect 1368 -24 1380 95
rect 1728 -24 1740 95
rect 1776 -24 1788 119
rect 1992 -24 2004 119
rect 2352 -24 2364 191
rect 2376 61 2388 239
rect 2520 133 2532 263
rect 2544 205 2556 287
rect 2568 229 2580 311
rect 2400 -24 2412 47
rect 2544 -24 2556 119
rect 2568 -24 2580 191
rect 2592 -24 2604 215
rect 2616 61 2628 335
rect 2640 -24 2652 47
rect 2664 -24 2676 407
rect 2712 325 2724 431
rect 2688 205 2700 311
rect 2688 -24 2700 191
rect 2712 -24 2724 191
rect 2736 37 2748 455
rect 2760 253 2772 479
rect 2760 -24 2772 -1
rect 2784 -24 2796 479
rect 2808 -24 2820 479
rect 2832 -24 2844 527
rect 2856 445 2868 575
rect 2856 -24 2868 287
rect 2880 133 2892 599
rect 2904 445 2916 623
rect 2928 589 2940 647
rect 2976 613 2988 671
rect 2904 -24 2916 287
rect 2928 -24 2940 407
rect 2952 -24 2964 575
rect 2976 -24 2988 407
rect 3000 277 3012 695
rect 3000 -24 3012 239
rect 3024 61 3036 719
rect 3048 -24 3060 599
rect 3072 157 3084 743
rect 3168 637 3180 767
rect 3192 685 3204 791
rect 3072 -24 3084 119
rect 3096 -24 3108 263
rect 3120 -24 3132 143
rect 3144 -24 3156 47
rect 3192 -24 3204 623
rect 3216 -24 3228 671
rect 3240 -24 3252 791
rect 3264 157 3276 791
rect 3288 -24 3300 143
rect 3312 -24 3324 815
rect 3336 -24 3348 719
rect 3360 181 3372 839
rect 3384 733 3396 863
rect 3384 -24 3396 167
rect 3408 -24 3420 695
rect 3432 -24 3444 695
rect 3456 -24 3468 863
rect 3552 637 3564 863
rect 3576 -24 3588 623
rect 3912 157 3924 887
rect 3936 -24 3948 143
rect 3960 109 3972 911
rect 4176 325 4188 935
rect 3984 -24 3996 95
rect 4200 -24 4212 311
rect 4536 85 4548 959
rect 4584 277 4596 983
rect 4680 805 4692 1007
rect 4704 709 4716 1031
rect 4560 -24 4572 71
rect 4608 -24 4620 263
rect 4728 109 4740 1055
rect 4752 517 4764 1079
rect 4776 589 4788 1103
rect 4800 541 4812 791
rect 4752 -24 4764 95
rect 4776 -24 4788 503
rect 4800 -24 4812 527
rect 4824 -24 4836 695
rect 4848 133 4860 1127
rect 4896 1045 4908 1151
rect 4920 997 4932 1175
rect 4872 -24 4884 575
rect 4896 -24 4908 527
rect 4944 421 4956 1031
rect 4920 -24 4932 119
rect 4944 -24 4956 407
rect 4968 -24 4980 983
rect 4992 181 5004 1199
rect 5040 997 5052 1223
rect 5016 -24 5028 407
rect 5040 -24 5052 167
rect 5064 -24 5076 983
rect 5088 -24 5100 959
rect 5112 325 5124 1247
rect 5136 -24 5148 1271
rect 5160 -24 5172 959
rect 5184 -24 5196 311
rect 5208 -24 5220 551
rect 5232 445 5244 1295
rect 5256 757 5268 1319
rect 5256 -24 5268 551
rect 5280 -24 5292 743
rect 5304 -24 5316 431
rect 5328 -24 5340 1319
rect 5352 613 5364 1319
rect 5376 781 5388 1343
rect 5400 949 5412 1367
rect 5376 -24 5388 599
rect 5400 -24 5412 767
rect 5424 -24 5436 935
rect 5448 709 5460 1391
rect 5472 1381 5484 1415
rect 5472 -24 5484 695
rect 5496 229 5508 1439
rect 5520 253 5532 1463
rect 5544 1165 5556 1487
rect 5496 -24 5508 95
rect 5520 -24 5532 215
rect 5544 -24 5556 239
rect 5568 -24 5580 1367
rect 5592 445 5604 1511
rect 5616 -24 5628 1151
rect 5640 637 5652 1535
rect 5664 1357 5676 1559
rect 5640 -24 5652 431
rect 5664 -24 5676 623
rect 5688 253 5700 1583
rect 5712 1045 5724 1607
rect 5712 -24 5724 239
rect 5736 -24 5748 1343
rect 5760 1333 5772 1631
rect 5760 -24 5772 1031
rect 5784 589 5796 1655
rect 5784 -24 5796 335
rect 5808 -24 5820 1319
rect 5832 493 5844 1679
rect 5856 -24 5868 575
rect 5880 -24 5892 479
rect 5928 -24 5940 1679
rect 5952 613 5964 1679
rect 5976 -24 5988 599
rect 6000 -24 6012 839
rect 6048 -24 6060 887
rect 6072 421 6084 1703
rect 6096 -24 6108 887
rect 6120 -24 6132 407
rect 6144 -24 6156 1703
rect 6168 109 6180 1703
rect 6192 -24 6204 95
rect 6216 -24 6228 407
rect 6240 -24 6252 1199
rect 6264 1117 6276 1727
rect 6288 -24 6300 1199
rect 6312 -24 6324 1103
rect 6360 -24 6372 1727
rect 6384 565 6396 1727
rect 6408 -24 6420 551
rect 6432 -24 6444 407
rect 6456 -24 6468 1727
rect 6552 1141 6564 1727
rect 6576 -24 6588 1127
rect 6912 157 6924 1751
rect 6960 1477 6972 1775
rect 6936 -24 6948 143
rect 6984 -24 6996 1463
rect 7176 661 7188 1799
rect 7200 -24 7212 647
rect 7584 229 7596 1823
rect 7728 757 7740 1847
rect 7608 -24 7620 215
rect 7752 -24 7764 743
rect 7776 -24 7788 407
rect 7800 -24 7812 1271
rect 7824 1141 7836 1871
rect 7848 -24 7860 1271
rect 7872 1213 7884 1895
rect 7896 1237 7908 1919
rect 7944 1429 7956 1943
rect 7872 709 7884 1127
rect 7872 -24 7884 695
rect 7896 -24 7908 1199
rect 7920 -24 7932 1223
rect 7944 -24 7956 695
rect 7968 373 7980 1967
rect 7992 -24 8004 1415
rect 8016 469 8028 1991
rect 8040 1549 8052 2015
rect 8064 1765 8076 2039
rect 8016 -24 8028 359
rect 8040 -24 8052 455
rect 8064 -24 8076 1535
rect 8088 589 8100 2063
rect 8112 973 8124 2087
rect 8112 -24 8124 575
rect 8136 373 8148 1751
rect 8136 -24 8148 359
rect 8160 -24 8172 959
rect 8184 589 8196 2111
rect 8208 421 8220 2135
rect 8184 -24 8196 359
rect 8232 -24 8244 575
rect 8256 -24 8268 407
rect 8280 -24 8292 1247
rect 8304 1189 8316 2159
rect 8328 -24 8340 1247
rect 8352 -24 8364 1175
rect 8400 -24 8412 2159
rect 8448 -24 8460 599
rect 8472 -24 8484 791
rect 8496 -24 8508 863
rect 8520 733 8532 2159
rect 8544 1861 8556 2183
rect 8568 2029 8580 2207
rect 8544 -24 8556 863
rect 8568 -24 8580 1847
rect 8592 -24 8604 2015
rect 8616 -24 8628 719
rect 8640 -24 8652 2207
rect 8664 181 8676 2207
rect 8688 325 8700 2231
rect 8688 -24 8700 167
rect 8712 -24 8724 311
rect 8736 -24 8748 2231
rect 8760 2101 8772 2231
rect 8784 -24 8796 2087
rect 8808 -24 8820 839
rect 8832 -24 8844 2231
rect 8880 -24 8892 2087
rect 8904 -24 8916 1991
rect 8928 -24 8940 2207
rect 8952 997 8964 2207
rect 8976 181 8988 983
rect 8976 -24 8988 167
rect 9000 -24 9012 167
rect 9024 -24 9036 2207
rect 9072 -24 9084 2087
rect 9096 -24 9108 383
rect 9120 -24 9132 2183
rect 9168 1525 9180 2183
rect 9168 -24 9180 983
rect 9192 -24 9204 1511
rect 9216 -24 9228 2183
rect 9264 -24 9276 2087
rect 9288 -24 9300 1967
rect 9312 -24 9324 2159
rect 9336 2077 9348 2159
rect 9360 997 9372 2063
rect 9360 -24 9372 983
rect 9384 -24 9396 983
rect 9408 -24 9420 1487
rect 9432 1165 9444 2183
rect 9456 685 9468 1487
rect 9456 -24 9468 671
rect 9480 -24 9492 1151
rect 9504 -24 9516 671
rect 9528 -24 9540 2183
rect 9552 1045 9564 2183
rect 9576 -24 9588 1031
rect 9624 -24 9636 1679
rect 9648 1477 9660 2207
rect 9672 325 9684 2231
rect 9696 1213 9708 2255
rect 9720 781 9732 1679
rect 9696 -24 9708 311
rect 9720 -24 9732 767
rect 9744 -24 9756 1463
rect 9768 1213 9780 2279
rect 9768 -24 9780 767
rect 9792 -24 9804 1175
rect 9816 397 9828 2303
rect 9840 2197 9852 2327
rect 9864 1573 9876 2351
rect 9840 -24 9852 1175
rect 9864 349 9876 383
rect 9864 -24 9876 335
rect 9888 -24 9900 2183
rect 9912 1261 9924 2375
rect 9936 973 9948 2399
rect 9960 1837 9972 2423
rect 9912 -24 9924 335
rect 9960 -24 9972 1559
rect 9984 -24 9996 1823
rect 10008 397 10020 1247
rect 10008 -24 10020 383
rect 10032 -24 10044 959
rect 10056 877 10068 2447
rect 10056 -24 10068 383
rect 10080 373 10092 2471
rect 10128 2293 10140 2495
rect 10104 -24 10116 863
rect 10128 -24 10140 359
rect 10152 -24 10164 2279
rect 10176 517 10188 2519
rect 10200 -24 10212 503
rect 10248 -24 10260 2519
rect 10272 589 10284 2519
rect 10296 133 10308 2543
rect 10320 -24 10332 575
rect 10344 -24 10356 119
rect 10392 -24 10404 2543
rect 10440 -24 10452 263
rect 10464 -24 10476 263
rect 10488 -24 10500 2519
rect 10512 1717 10524 2519
rect 10536 -24 10548 1703
rect 10584 -24 10596 2327
rect 10608 613 10620 2543
rect 10632 277 10644 2567
rect 10656 -24 10668 2327
rect 10680 1957 10692 2591
rect 10680 -24 10692 599
rect 10704 -24 10716 1943
rect 10728 -24 10740 263
rect 10752 -24 10764 1871
rect 10776 1429 10788 2615
rect 10824 2077 10836 2639
rect 10848 2389 10860 2663
rect 10800 -24 10812 1871
rect 10824 -24 10836 1415
rect 10848 -24 10860 2063
rect 10872 -24 10884 2375
rect 10896 -24 10908 2663
rect 10920 949 10932 2663
rect 10944 1405 10956 2687
rect 11016 2245 11028 2711
rect 11040 1933 11052 2735
rect 10944 -24 10956 935
rect 10968 -24 10980 1391
rect 10992 -24 11004 791
rect 11016 -24 11028 1031
rect 11064 -24 11076 2231
rect 11088 -24 11100 1919
rect 11112 -24 11124 1583
rect 11136 -24 11148 2759
rect 11160 -24 11172 2159
rect 11184 829 11196 2783
rect 11232 2749 11244 2807
rect 11208 -24 11220 2159
rect 11256 1861 11268 2831
rect 11232 -24 11244 815
rect 11256 -24 11268 647
rect 11280 181 11292 2855
rect 11304 -24 11316 2735
rect 11328 -24 11340 1847
rect 11352 1549 11364 2879
rect 11352 -24 11364 647
rect 11376 -24 11388 1535
rect 11400 709 11412 2903
rect 11424 181 11436 2927
rect 11448 829 11460 2951
rect 11400 -24 11412 167
rect 11448 -24 11460 695
rect 11472 -24 11484 815
rect 11520 373 11532 2975
rect 11568 1309 11580 2999
rect 11592 1549 11604 3023
rect 11616 1813 11628 3047
rect 11544 277 11556 359
rect 11496 -24 11508 167
rect 11544 -24 11556 263
rect 11568 -24 11580 263
rect 11592 -24 11604 1295
rect 11616 -24 11628 1535
rect 11640 -24 11652 1799
rect 11664 1717 11676 3071
rect 11688 1861 11700 3095
rect 11712 3085 11724 3119
rect 11688 -24 11700 1703
rect 11712 -24 11724 1847
rect 11736 1093 11748 3071
rect 11784 2485 11796 3143
rect 11808 1717 11820 3167
rect 11736 -24 11748 1079
rect 11760 805 11772 1079
rect 11760 -24 11772 791
rect 11784 -24 11796 791
rect 11832 -24 11844 2471
rect 11856 2437 11868 3191
rect 11880 2725 11892 3215
rect 11904 2533 11916 3239
rect 11856 1645 11868 1703
rect 11856 -24 11868 1631
rect 11880 -24 11892 2423
rect 11928 1717 11940 3263
rect 11904 1021 11916 1631
rect 11904 -24 11916 1007
rect 11928 -24 11940 1007
rect 11952 853 11964 3287
rect 11976 -24 11988 2711
rect 12000 1597 12012 3311
rect 12000 -24 12012 839
rect 12024 -24 12036 2519
rect 12048 1357 12060 3335
rect 12048 -24 12060 407
rect 12072 -24 12084 1703
rect 12096 37 12108 3359
rect 12120 37 12132 1583
rect 12144 37 12156 1343
rect 12168 517 12180 3383
rect 12120 -24 12132 -1
rect 12144 -24 12156 -1
rect 12168 -24 12180 -1
rect 12192 -24 12204 503
rect 12216 -24 12228 3383
rect 12240 1765 12252 3383
rect 12264 1909 12276 3407
rect 12264 -24 12276 1751
rect 12288 -24 12300 1895
rect 12312 -24 12324 3407
rect 12336 1045 12348 3407
rect 12360 3205 12372 3431
rect 12360 -24 12372 1031
rect 12384 -24 12396 3191
rect 12432 -24 12444 3431
rect 12480 -24 12492 1151
rect 12504 -24 12516 671
rect 12528 -24 12540 2543
rect 12552 1309 12564 3431
rect 12576 2101 12588 3455
rect 12624 2605 12636 3479
rect 12576 -24 12588 1295
rect 12600 -24 12612 2543
rect 12624 -24 12636 2087
rect 12648 -24 12660 2591
rect 12672 -24 12684 3119
rect 12696 877 12708 3503
rect 12720 -24 12732 3119
rect 12744 -24 12756 863
rect 12768 -24 12780 3503
rect 12792 541 12804 3503
rect 12816 2653 12828 3527
rect 12816 -24 12828 527
rect 12840 -24 12852 2639
rect 12864 -24 12876 3527
rect 12936 2845 12948 3527
rect 12912 -24 12924 1463
rect 12960 -24 12972 2831
rect 12984 589 12996 3551
rect 13008 133 13020 3575
rect 13032 -24 13044 575
rect 13056 -24 13068 119
rect 13104 -24 13116 3575
rect 13128 3397 13140 3575
rect 13152 -24 13164 3383
rect 13176 -24 13188 863
rect 13200 -24 13212 3575
rect 13272 1453 13284 3575
rect 13368 2653 13380 3599
rect 13392 3181 13404 3623
rect 13248 -24 13260 695
rect 13296 -24 13308 1439
rect 13368 -24 13380 239
rect 13392 -24 13404 2639
rect 13416 -24 13428 3167
rect 13440 325 13452 3647
rect 13464 1645 13476 3671
rect 13488 3469 13500 3695
rect 13464 -24 13476 311
rect 13488 -24 13500 1631
rect 13512 -24 13524 3455
rect 13536 -24 13548 3695
rect 13560 2029 13572 3695
rect 13584 3541 13596 3719
rect 13584 -24 13596 2015
rect 13608 -24 13620 3527
rect 13656 -24 13668 3719
rect 13680 2269 13692 3719
rect 13704 -24 13716 2255
rect 13752 -24 13764 3719
rect 13824 -24 13836 2303
rect 13872 1933 13884 3719
rect 14016 2269 14028 3743
rect 14160 3733 14172 3767
rect 13896 -24 13908 1919
rect 13968 -24 13980 551
rect 14040 -24 14052 2255
rect 14112 -24 14124 1919
rect 14184 -24 14196 3719
rect 14232 205 14244 3791
rect 14256 1165 14268 3815
rect 14256 -24 14268 191
rect 14280 -24 14292 1151
rect 14328 -24 14340 3815
rect 14376 1477 14388 3815
rect 14376 -24 14388 191
rect 14400 -24 14412 1463
rect 14424 -24 14436 3815
rect 14448 709 14460 3815
rect 14472 1045 14484 3839
rect 14472 -24 14484 695
rect 14496 -24 14508 1031
rect 14520 -24 14532 3839
rect 14544 109 14556 3839
rect 14568 1573 14580 3863
rect 14568 -24 14580 95
rect 14592 -24 14604 1559
rect 14616 -24 14628 3863
rect 14640 253 14652 3863
rect 14664 2125 14676 3887
rect 14664 -24 14676 239
rect 14688 -24 14700 2111
rect 14712 -24 14724 3887
rect 14736 2365 14748 3887
rect 14760 -24 14772 2351
rect 14784 -24 14796 191
rect 14808 -24 14820 3887
rect 14832 3829 14844 3887
rect 14856 205 14868 3815
rect 14856 -24 14868 191
rect 14880 -24 14892 191
rect 14904 -24 14916 3887
rect 14928 733 14940 3887
rect 14952 325 14964 719
rect 14952 -24 14964 311
rect 14976 -24 14988 311
rect 15000 -24 15012 2183
rect 15024 181 15036 3911
rect 15072 3253 15084 3935
rect 15048 -24 15060 2183
rect 15072 -24 15084 167
rect 15096 -24 15108 3239
rect 15120 -24 15132 3935
rect 15168 -24 15180 2255
rect 15240 -24 15252 1919
rect 15312 -24 15324 3935
rect 15360 1333 15372 3959
rect 15384 2581 15396 3983
rect 15384 -24 15396 1319
rect 15408 -24 15420 2567
rect 15432 -24 15444 1487
rect 15456 -24 15468 3983
rect 15504 -24 15516 2255
rect 15576 -24 15588 1919
rect 15624 325 15636 3983
rect 15840 3589 15852 4007
rect 15648 -24 15660 311
rect 15720 -24 15732 2255
rect 15792 -24 15804 1919
rect 15864 -24 15876 3575
rect 16056 2941 16068 4031
rect 15936 -24 15948 2255
rect 16008 -24 16020 1919
rect 16080 -24 16092 2927
rect 16272 2869 16284 4055
rect 16152 -24 16164 2255
rect 16224 -24 16236 1919
rect 16296 -24 16308 2855
rect 16488 2533 16500 4079
rect 16704 2965 16716 4103
rect 16368 -24 16380 2255
rect 16440 -24 16452 1919
rect 16512 -24 16524 2519
rect 16584 -24 16596 2255
rect 16656 -24 16668 1919
rect 16728 -24 16740 2951
rect 16800 -24 16812 2255
rect 16920 1933 16932 4127
rect 16872 -24 16884 1919
rect 16944 -24 16956 1919
rect 17016 -24 17028 2255
rect 17088 -24 17100 4127
rect 17136 3061 17148 4151
rect 17160 -24 17172 3047
rect 17232 -24 17244 2255
rect 17304 -24 17316 4127
rect 17352 2269 17364 4175
rect 17376 -24 17388 2255
rect 17448 -24 17460 4175
rect 17520 -24 17532 4127
rect 17568 2389 17580 4175
rect 17592 -24 17604 2375
rect 17664 -24 17676 1967
rect 17736 -24 17748 4127
rect 17808 -24 17820 3839
rect 17880 -24 17892 1991
rect 17952 -24 17964 4127
rect 18024 -24 18036 887
rect 18096 -24 18108 3287
rect 18168 -24 18180 4127
rect 18264 2365 18276 4199
rect 18288 1525 18300 4223
rect 18240 -24 18252 743
rect 18312 -24 18324 2351
rect 18336 1765 18348 4247
rect 18336 -24 18348 1511
rect 18360 -24 18372 1751
rect 18384 -24 18396 4247
rect 18408 1429 18420 4247
rect 18432 3589 18444 4271
rect 18456 3757 18468 4295
rect 18432 -24 18444 1415
rect 18456 -24 18468 3575
rect 18480 -24 18492 3743
rect 18504 -24 18516 4295
rect 18528 781 18540 4295
rect 18552 1885 18564 4319
rect 18552 -24 18564 767
rect 18576 -24 18588 1871
rect 18600 -24 18612 2159
rect 18624 2077 18636 4343
rect 18648 -24 18660 2159
rect 18672 -24 18684 2063
rect 18720 -24 18732 4343
rect 18744 85 18756 4343
rect 18768 2725 18780 4367
rect 18768 -24 18780 71
rect 18792 -24 18804 2711
rect 18816 -24 18828 4367
rect 18864 445 18876 4367
rect 18864 -24 18876 167
rect 18888 -24 18900 431
rect 18912 -24 18924 1343
rect 18936 1093 18948 4391
rect 18960 -24 18972 1343
rect 18984 -24 18996 1079
rect 19032 -24 19044 3767
rect 19056 757 19068 4415
rect 19080 3493 19092 4439
rect 19080 661 19092 743
rect 19080 -24 19092 647
rect 19104 -24 19116 3767
rect 19128 -24 19140 3479
rect 19152 589 19164 4463
rect 19176 -24 19188 647
rect 19200 -24 19212 575
rect 19224 -24 19236 4463
rect 19248 1933 19260 4463
rect 19272 1957 19284 4487
rect 19272 -24 19284 1919
rect 19296 -24 19308 1943
rect 19344 -24 19356 4487
rect 19368 2797 19380 4487
rect 19392 3661 19404 4511
rect 19392 -24 19404 2783
rect 19416 -24 19428 3647
rect 19464 -24 19476 4511
rect 19488 2437 19500 4511
rect 19512 -24 19524 2423
rect 19560 -24 19572 4511
rect 19608 3877 19620 4511
rect 19632 973 19644 3863
rect 19632 -24 19644 959
rect 19656 -24 19668 959
rect 19704 -24 19716 4511
rect 19800 1933 19812 4511
rect 19824 -24 19836 1919
rect 20208 1717 20220 4535
rect 20328 3613 20340 4559
rect 20352 2341 20364 4583
rect 20424 4405 20436 4607
rect 20184 -24 20196 1535
rect 20232 -24 20244 1703
rect 20376 1405 20388 3599
rect 20376 -24 20388 1391
rect 20400 949 20412 2327
rect 20400 -24 20412 935
rect 20424 -24 20436 1391
rect 20448 37 20460 4631
rect 20472 37 20484 4391
rect 20496 37 20508 935
rect 20472 -24 20484 -1
rect 20496 -24 20508 -1
rect 20520 -24 20532 -1
rect 20544 -24 20556 4631
rect 20568 3445 20580 4631
rect 20592 -24 20604 3431
rect 20640 -24 20652 4631
rect 20712 3109 20724 4631
rect 20712 -24 20724 167
rect 20736 -24 20748 3095
rect 20760 -24 20772 4631
rect 20808 541 20820 4631
rect 20808 -24 20820 167
rect 20832 -24 20844 527
rect 20856 -24 20868 4631
rect 20904 -24 20916 95
rect 20928 -24 20940 2711
rect 20952 -24 20964 2015
rect 20976 301 20988 4631
rect 21000 -24 21012 2015
rect 21024 -24 21036 287
rect 21048 -24 21060 863
rect 21072 469 21084 4655
rect 21096 -24 21108 863
rect 21120 -24 21132 455
rect 21144 -24 21156 4655
rect 21192 -24 21204 119
rect 21216 -24 21228 863
rect 21240 -24 21252 4631
rect 21264 1693 21276 4631
rect 21288 181 21300 1679
rect 21288 -24 21300 167
rect 21312 -24 21324 167
rect 21336 -24 21348 4631
rect 21384 -24 21396 2567
rect 21408 -24 21420 719
rect 21432 -24 21444 4607
rect 21456 349 21468 4607
rect 21480 3157 21492 4631
rect 21480 -24 21492 335
rect 21504 -24 21516 3143
rect 21528 -24 21540 695
rect 21552 613 21564 4655
rect 21576 4045 21588 4679
rect 21576 -24 21588 695
rect 21600 -24 21612 4031
rect 21624 1573 21636 4703
rect 21624 -24 21636 599
rect 21648 -24 21660 1559
rect 21672 -24 21684 4703
rect 21720 2557 21732 4703
rect 21720 -24 21732 1055
rect 21744 -24 21756 2543
rect 21768 -24 21780 191
rect 21792 -24 21804 4703
rect 21840 3829 21852 4703
rect 21840 -24 21852 935
rect 21864 -24 21876 3815
rect 21912 -24 21924 4703
rect 21936 3085 21948 4703
rect 21960 -24 21972 3071
rect 21984 -24 21996 407
rect 22032 -24 22044 4703
rect 22056 4141 22068 4703
rect 22080 -24 22092 4127
rect 22128 -24 22140 4703
rect 22176 2989 22188 4703
rect 22200 2197 22212 4727
rect 22200 -24 22212 1727
rect 22224 -24 22236 2975
rect 22248 2437 22260 4751
rect 22248 -24 22260 2183
rect 22272 -24 22284 2423
rect 22296 -24 22308 4751
rect 22320 1141 22332 4751
rect 22344 3229 22356 4775
rect 22344 -24 22356 1127
rect 22368 -24 22380 3215
rect 22392 -24 22404 1871
rect 22416 853 22428 4799
rect 22440 -24 22452 1871
rect 22464 -24 22476 839
rect 22488 -24 22500 2543
rect 22512 -24 22524 1487
rect 22536 -24 22548 4799
rect 22560 1645 22572 4799
rect 22584 -24 22596 1631
rect 22632 -24 22644 4799
rect 22680 3037 22692 4799
rect 22704 -24 22716 3023
rect 22728 -24 22740 2039
rect 22752 -24 22764 4079
rect 22776 3181 22788 4823
rect 22800 3445 22812 4847
rect 22800 -24 22812 3167
rect 22824 -24 22836 4079
rect 22848 -24 22860 3431
rect 22872 -24 22884 2423
rect 22896 -24 22908 4847
rect 22944 2029 22956 4847
rect 22944 -24 22956 935
rect 22968 -24 22980 2015
rect 22992 -24 23004 4751
rect 23016 253 23028 4871
rect 23040 -24 23052 4751
rect 23064 -24 23076 239
rect 23088 -24 23100 4871
rect 23112 517 23124 4871
rect 23136 949 23148 4895
rect 23160 4621 23172 4919
rect 23136 -24 23148 503
rect 23160 -24 23172 935
rect 23184 -24 23196 4607
rect 23208 -24 23220 527
rect 23232 -24 23244 3983
rect 23256 3781 23268 4943
rect 23280 2293 23292 4967
rect 23304 3853 23316 4991
rect 23280 -24 23292 719
rect 23304 -24 23316 3767
rect 23328 -24 23340 3983
rect 23352 -24 23364 3839
rect 23376 -24 23388 2279
rect 23400 613 23412 5015
rect 23424 -24 23436 599
rect 23472 -24 23484 479
rect 23520 61 23532 5039
rect 23544 757 23556 5063
rect 23544 -24 23556 47
rect 23568 -24 23580 743
rect 23592 -24 23604 527
rect 23616 -24 23628 5063
rect 23640 1021 23652 5063
rect 23688 3325 23700 5087
rect 23664 541 23676 1007
rect 23664 -24 23676 527
rect 23688 -24 23700 527
rect 23712 -24 23724 3311
rect 23736 -24 23748 5087
rect 23784 -24 23796 4727
rect 23808 2245 23820 5087
rect 23808 -24 23820 527
rect 23832 -24 23844 2231
rect 23856 -24 23868 5087
rect 23880 2077 23892 5087
rect 23904 4141 23916 5111
rect 23904 -24 23916 2063
rect 23928 -24 23940 4127
rect 23952 -24 23964 191
rect 23976 -24 23988 5111
rect 24000 2533 24012 5111
rect 24024 4381 24036 5135
rect 24048 4141 24060 4367
rect 24024 -24 24036 2519
rect 24048 -24 24060 4127
rect 24072 -24 24084 4127
rect 24096 -24 24108 5135
rect 24120 325 24132 5135
rect 24144 61 24156 311
rect 24144 -24 24156 47
rect 24168 -24 24180 47
rect 24192 -24 24204 2231
rect 24216 -24 24228 2735
rect 24240 1813 24252 5159
rect 24264 1933 24276 5183
rect 24264 -24 24276 1799
rect 24288 -24 24300 2735
rect 24312 -24 24324 1919
rect 24336 -24 24348 5183
rect 24360 637 24372 5183
rect 24384 973 24396 5207
rect 24384 -24 24396 623
rect 24408 133 24420 959
rect 24408 -24 24420 119
rect 24432 -24 24444 119
rect 24456 -24 24468 5207
rect 24480 1117 24492 5207
rect 24504 1525 24516 5231
rect 24528 1693 24540 5255
rect 24552 2173 24564 5279
rect 24504 -24 24516 1103
rect 24528 -24 24540 1511
rect 24552 -24 24564 1679
rect 24576 -24 24588 2159
rect 24600 -24 24612 5279
rect 24648 -24 24660 3359
rect 24696 -24 24708 5255
rect 24768 -24 24780 2543
rect 24792 -24 24804 191
rect 24816 -24 24828 5231
rect 24840 2581 24852 5231
rect 24864 -24 24876 2567
rect 24888 -24 24900 2063
rect 24936 -24 24948 5231
rect 24960 4861 24972 5231
rect 24984 2077 24996 4847
rect 24984 -24 24996 2063
rect 25008 -24 25020 2063
rect 25032 -24 25044 5231
rect 25080 -24 25092 2543
rect 25104 -24 25116 623
rect 25128 -24 25140 5207
rect 25176 3637 25188 5207
rect 25176 -24 25188 71
rect 25200 -24 25212 3623
rect 25224 -24 25236 5207
rect 25248 877 25260 5207
rect 25272 -24 25284 863
rect 25296 -24 25308 4847
rect 25344 -24 25356 5207
rect 25368 2725 25380 5207
rect 25392 -24 25404 2711
rect 25416 -24 25428 3455
rect 25440 -24 25452 5207
rect 25464 1309 25476 5207
rect 25488 -24 25500 1295
rect 25512 -24 25524 3623
rect 25536 -24 25548 5207
rect 25632 3613 25644 5207
rect 25656 -24 25668 3599
rect 26016 -24 26028 1895
rect 26064 -24 26076 839
rect 26208 -24 26220 743
rect 26232 -24 26244 3623
rect 26256 -24 26268 5207
rect 26304 1405 26316 5207
rect 26304 -24 26316 71
rect 26328 -24 26340 1391
rect 26352 -24 26364 1079
rect 26376 613 26388 5231
rect 26400 661 26412 5255
rect 26448 1645 26460 5279
rect 26400 -24 26412 599
rect 26424 -24 26436 1079
rect 26448 -24 26460 647
rect 26472 -24 26484 1631
rect 26496 -24 26508 5279
rect 26544 -24 26556 623
rect 26568 -24 26580 4847
rect 26592 -24 26604 5255
rect 26640 3661 26652 5255
rect 26640 -24 26652 2543
rect 26664 -24 26676 3647
rect 26712 -24 26724 5255
rect 26736 4765 26748 5255
rect 26760 -24 26772 4751
rect 26784 349 26796 5279
rect 26784 -24 26796 47
rect 26808 -24 26820 335
rect 26832 -24 26844 3575
rect 26856 1621 26868 5303
rect 26880 -24 26892 3575
rect 26904 -24 26916 1607
rect 26952 -24 26964 4511
rect 26976 3517 26988 5327
rect 27000 2533 27012 4511
rect 27000 -24 27012 2519
rect 27024 -24 27036 3503
rect 27048 -24 27060 2519
rect 27072 -24 27084 5327
rect 27120 -24 27132 4847
rect 27144 -24 27156 719
rect 27168 -24 27180 2063
rect 27192 -24 27204 5303
rect 27216 589 27228 5303
rect 27240 1141 27252 5327
rect 27240 -24 27252 575
rect 27264 -24 27276 1127
rect 27288 -24 27300 5327
rect 27312 829 27324 5327
rect 27336 -24 27348 815
rect 27360 -24 27372 1295
rect 27384 -24 27396 4127
rect 27408 -24 27420 5327
rect 27456 1597 27468 5327
rect 27456 -24 27468 71
rect 27480 -24 27492 1583
rect 27504 -24 27516 4559
rect 27528 2773 27540 5351
rect 27552 3349 27564 5375
rect 27552 -24 27564 2759
rect 27576 -24 27588 4559
rect 27600 4213 27612 5399
rect 27600 -24 27612 3335
rect 27624 -24 27636 4199
rect 27648 -24 27660 5399
rect 27696 -24 27708 3503
rect 27720 -24 27732 4511
rect 27744 -24 27756 5375
rect 27792 4909 27804 5375
rect 27792 -24 27804 743
rect 27816 -24 27828 4895
rect 27840 -24 27852 3359
rect 27864 3037 27876 5399
rect 27888 -24 27900 3359
rect 27912 -24 27924 3023
rect 27936 -24 27948 5399
rect 27960 1357 27972 5399
rect 27984 61 27996 1343
rect 27984 -24 27996 47
rect 28008 -24 28020 47
rect 28032 -24 28044 5399
rect 28080 3205 28092 5399
rect 28080 -24 28092 1343
rect 28104 -24 28116 3191
rect 28128 -24 28140 5399
rect 28176 -24 28188 743
rect 28200 -24 28212 335
rect 28248 -24 28260 5375
rect 28296 -24 28308 743
rect 28320 -24 28332 3191
rect 28344 -24 28356 5351
rect 28392 4957 28404 5351
rect 28392 -24 28404 743
rect 28416 -24 28428 4943
rect 28440 -24 28452 5351
rect 28488 -24 28500 527
rect 28512 -24 28524 167
rect 28536 -24 28548 5327
rect 28584 1861 28596 5327
rect 28584 -24 28596 527
rect 28608 -24 28620 1847
rect 28632 -24 28644 5327
rect 28680 3757 28692 5327
rect 28680 -24 28692 527
rect 28704 -24 28716 3743
rect 28728 -24 28740 5327
rect 28752 1429 28764 5327
rect 28776 -24 28788 1415
rect 28800 -24 28812 1055
rect 28824 -24 28836 5327
rect 28872 -24 28884 863
rect 28896 -24 28908 119
rect 28920 -24 28932 5303
rect 28968 -24 28980 527
rect 28992 -24 29004 -1
rect 29016 -24 29028 5279
rect 29064 -24 29076 455
rect 29088 -24 29100 119
rect 29112 -24 29124 5255
rect 29160 -24 29172 815
rect 29184 -24 29196 1295
rect 29208 -24 29220 2519
rect 29232 -24 29244 5231
rect 29256 4813 29268 5231
rect 29280 541 29292 4799
rect 29280 -24 29292 527
rect 29304 -24 29316 527
rect 29328 -24 29340 5231
rect 29424 5029 29436 5231
rect 29448 -24 29460 5015
rect 29976 2557 29988 5255
rect 30000 2797 30012 5279
rect 29856 -24 29868 767
rect 30000 -24 30012 2543
rect 30024 -24 30036 2783
rect 30072 -24 30084 5279
rect 30096 3085 30108 5279
rect 30120 1429 30132 3071
rect 30120 -24 30132 1415
rect 30144 -24 30156 1415
rect 30168 -24 30180 5279
rect 30216 1237 30228 5279
rect 30240 1405 30252 5303
rect 30216 -24 30228 695
rect 30240 -24 30252 1223
rect 30264 -24 30276 1391
rect 30288 -24 30300 5303
rect 30312 2989 30324 5303
rect 30336 -24 30348 2975
rect 30384 -24 30396 5303
rect 30432 3565 30444 5303
rect 30456 3709 30468 5327
rect 30456 -24 30468 3551
rect 30480 -24 30492 3695
rect 30528 -24 30540 5327
rect 30576 -24 30588 2999
rect 30600 -24 30612 1055
rect 30648 -24 30660 5303
rect 30672 3589 30684 5303
rect 30696 -24 30708 3575
rect 30720 -24 30732 1127
rect 30744 -24 30756 3455
rect 30768 -24 30780 5303
rect 30816 -24 30828 1847
rect 30840 -24 30852 71
rect 30864 -24 30876 2063
rect 30888 -24 30900 5279
rect 30936 4861 30948 5279
rect 30936 -24 30948 1847
rect 30960 -24 30972 4847
rect 31008 -24 31020 5279
rect 31056 -24 31068 959
rect 31080 -24 31092 1847
rect 31128 -24 31140 5255
rect 31152 4621 31164 5255
rect 31176 4405 31188 4607
rect 31176 -24 31188 4391
rect 31200 -24 31212 4391
rect 31224 -24 31236 4847
rect 31248 -24 31260 5255
rect 31296 -24 31308 191
rect 31320 -24 31332 1847
rect 31368 -24 31380 3623
rect 31392 2677 31404 5255
rect 31416 -24 31428 3623
rect 31440 3613 31452 5279
rect 31440 -24 31452 2663
rect 31464 -24 31476 3599
rect 31488 -24 31500 5279
rect 31512 2725 31524 5279
rect 31536 1861 31548 2711
rect 31536 -24 31548 1847
rect 31560 -24 31572 1847
rect 31584 -24 31596 5279
rect 31632 -24 31644 3311
rect 31656 -24 31668 4391
rect 31680 -24 31692 4847
rect 31704 -24 31716 5231
rect 31728 2293 31740 5231
rect 31752 2701 31764 5231
rect 31752 -24 31764 2279
rect 31776 -24 31788 2687
rect 31800 -24 31812 3431
rect 31824 2389 31836 5183
rect 31848 -24 31860 3431
rect 31872 -24 31884 2375
rect 31896 -24 31908 5087
rect 31920 2845 31932 5087
rect 31944 2869 31956 5087
rect 31968 3061 31980 5087
rect 31944 -24 31956 2831
rect 31968 -24 31980 2855
rect 31992 -24 32004 3047
rect 32016 -24 32028 5015
rect 32064 4693 32076 4991
rect 32112 4933 32124 4967
rect 32064 -24 32076 71
rect 32088 -24 32100 4679
rect 32112 -24 32124 4871
rect 32136 4021 32148 4967
rect 32160 4837 32172 4967
rect 32256 4933 32268 4967
rect 32280 4933 32292 4967
rect 32304 4933 32316 4967
rect 32328 4933 32340 4967
rect 32352 4933 32364 4967
rect 32376 4933 32388 4967
rect 32400 4933 32412 4967
rect 32424 4933 32436 4967
rect 32448 4933 32460 4967
rect 32472 4933 32484 4967
rect 59760 4933 59772 4967
rect 32184 4357 32196 4823
rect 32208 4693 32220 4727
rect 32208 4621 32220 4655
rect 32208 4525 32220 4559
rect 32208 4357 32220 4391
rect 32232 4261 32244 4823
rect 32208 4213 32220 4247
rect 32208 4093 32220 4127
rect 32160 -24 32172 4007
rect 32184 2245 32196 4079
rect 32208 3781 32220 3887
rect 32208 3661 32220 3695
rect 32208 3445 32220 3551
rect 32208 3157 32220 3311
rect 32208 3013 32220 3047
rect 32208 2701 32220 2735
rect 32208 2605 32220 2639
rect 32208 2413 32220 2495
rect 32208 2245 32220 2351
rect 32232 2149 32244 4103
rect 32256 2893 32268 4871
rect 32280 2917 32292 4871
rect 32304 3925 32316 4871
rect 32328 3973 32340 4871
rect 32352 4549 32364 4871
rect 32376 4645 32388 4871
rect 32376 4429 32388 4535
rect 32208 -24 32220 2135
rect 32280 -24 32292 2879
rect 32304 -24 32316 2903
rect 32328 -24 32340 3911
rect 32352 -24 32364 3959
rect 32376 -24 32388 2975
rect 32400 493 32412 4871
rect 32424 1213 32436 4871
rect 32448 2821 32460 4871
rect 32472 2005 32484 4871
rect 32496 4837 32508 4871
rect 32496 4645 32508 4703
rect 32496 4285 32508 4415
rect 32424 -24 32436 479
rect 32448 -24 32460 1199
rect 32496 -24 32508 3983
rect 32520 397 32532 4871
rect 32544 4549 32556 4871
rect 32544 4285 32556 4511
rect 32544 397 32556 4031
rect 32568 1453 32580 4871
rect 32592 2269 32604 4871
rect 32592 1789 32604 1991
rect 32544 -24 32556 383
rect 32568 -24 32580 695
rect 32592 -24 32604 1583
rect 32616 565 32628 4871
rect 32640 2989 32652 4871
rect 32664 3949 32676 4871
rect 32688 3733 32700 4871
rect 32640 2821 32652 2903
rect 32640 565 32652 2471
rect 32664 2005 32676 2903
rect 32664 1597 32676 1967
rect 32640 -24 32652 551
rect 32664 -24 32676 1439
rect 32688 -24 32700 3551
rect 32712 901 32724 4871
rect 32736 2989 32748 4871
rect 32760 4477 32772 4871
rect 32760 3805 32772 4031
rect 32760 3421 32772 3719
rect 32760 2485 32772 2903
rect 32736 1381 32748 2471
rect 32760 1789 32772 2447
rect 32736 -24 32748 887
rect 32760 -24 32772 1367
rect 32784 805 32796 4871
rect 32808 4429 32820 4871
rect 32832 4045 32844 4871
rect 32856 3949 32868 4871
rect 32880 4717 32892 4775
rect 32808 3733 32820 3935
rect 32832 3565 32844 3791
rect 32808 2989 32820 3551
rect 32808 997 32820 2951
rect 32832 997 32844 3527
rect 32856 997 32868 3911
rect 32880 2005 32892 4679
rect 32904 3805 32916 4895
rect 32904 2269 32916 3767
rect 32808 589 32820 959
rect 32832 805 32844 863
rect 32784 -24 32796 575
rect 32832 -24 32844 791
rect 32856 -24 32868 863
rect 32880 -24 32892 1967
rect 32904 -24 32916 2087
rect 32928 2005 32940 4871
rect 32952 4429 32964 4847
rect 32952 2101 32964 4391
rect 32976 2485 32988 4823
rect 33000 2917 33012 4775
rect 33024 4405 33036 4751
rect 32952 -24 32964 2087
rect 32976 -24 32988 2447
rect 33000 -24 33012 2519
rect 33024 -24 33036 4295
rect 33048 2989 33060 4727
rect 33216 4693 33228 4727
rect 33336 4693 33348 4727
rect 33384 4693 33396 4727
rect 41160 4693 41172 4727
rect 59040 4693 59052 4727
rect 59760 4693 59772 4727
rect 33072 3565 33084 4655
rect 33096 3565 33108 4631
rect 33120 3733 33132 4607
rect 33072 -24 33084 3407
rect 33144 1693 33156 4583
rect 33168 3805 33180 4511
rect 33192 3805 33204 4463
rect 41160 4453 41172 4487
rect 59040 4453 59052 4487
rect 59760 4453 59772 4487
rect 33216 3949 33228 4415
rect 33240 3949 33252 4391
rect 33264 4045 33276 4367
rect 33120 -24 33132 1679
rect 33192 -24 33204 2975
rect 33264 2965 33276 3983
rect 33216 -24 33228 431
rect 33240 -24 33252 1031
rect 33288 613 33300 4343
rect 33312 2965 33324 4295
rect 33336 2941 33348 4295
rect 33360 2941 33372 4271
rect 33384 3493 33396 4271
rect 33408 2917 33420 4247
rect 33432 3493 33444 4199
rect 33264 -24 33276 599
rect 33312 -24 33324 71
rect 33336 -24 33348 1871
rect 33384 -24 33396 2903
rect 33432 -24 33444 3119
rect 33456 -24 33468 4199
rect 33480 4069 33492 4247
rect 41160 4213 41172 4247
rect 59040 4213 59052 4247
rect 59760 4213 59772 4247
rect 33504 2701 33516 4199
rect 33528 4069 33540 4175
rect 33480 -24 33492 2687
rect 33528 -24 33540 1175
rect 33552 -24 33564 4175
rect 33600 3373 33612 4175
rect 33576 -24 33588 3359
rect 33696 3085 33708 4151
rect 33624 -24 33636 2855
rect 33672 -24 33684 3071
rect 33816 3061 33828 4127
rect 33744 -24 33756 71
rect 33768 -24 33780 527
rect 33792 -24 33804 3047
rect 33840 -24 33852 71
rect 33864 -24 33876 2975
rect 33936 757 33948 4103
rect 33912 -24 33924 743
rect 33960 -24 33972 4103
rect 34032 2557 34044 4103
rect 33984 -24 33996 1751
rect 34008 -24 34020 2543
rect 34056 -24 34068 4103
rect 34080 -24 34092 3455
rect 34128 133 34140 4103
rect 34104 -24 34116 119
rect 34152 -24 34164 4103
rect 34224 4045 34236 4103
rect 34176 -24 34188 1175
rect 34200 -24 34212 4031
rect 34344 1357 34356 4079
rect 34440 3037 34452 4055
rect 34248 -24 34260 71
rect 34272 -24 34284 -1
rect 34320 -24 34332 1343
rect 34368 -24 34380 575
rect 34392 -24 34404 2087
rect 34416 -24 34428 3023
rect 34464 -24 34476 4055
rect 34536 3517 34548 4055
rect 34488 -24 34500 1175
rect 34512 -24 34524 3503
rect 34632 1309 34644 4031
rect 34560 -24 34572 1175
rect 34608 -24 34620 1295
rect 34680 -24 34692 4031
rect 34704 -24 34716 719
rect 34728 -24 34740 4055
rect 34800 4021 34812 4055
rect 34752 -24 34764 2975
rect 34776 -24 34788 4007
rect 34824 -24 34836 4055
rect 34848 -24 34860 4079
rect 34896 3349 34908 4079
rect 34872 -24 34884 3335
rect 34920 -24 34932 4079
rect 34944 -24 34956 4031
rect 34992 3589 35004 4079
rect 34968 -24 34980 3575
rect 35016 -24 35028 4079
rect 35040 -24 35052 3143
rect 35088 2293 35100 4079
rect 35064 -24 35076 2279
rect 35112 -24 35124 4079
rect 35136 -24 35148 4103
rect 35208 3709 35220 4103
rect 35184 -24 35196 3695
rect 35232 -24 35244 4103
rect 35256 -24 35268 4127
rect 35328 2197 35340 4127
rect 35304 -24 35316 2183
rect 35352 -24 35364 4127
rect 35376 -24 35388 4151
rect 35400 -24 35412 4175
rect 35448 3421 35460 4175
rect 35424 -24 35436 3407
rect 35472 -24 35484 3503
rect 35568 3445 35580 4151
rect 35496 -24 35508 2687
rect 35544 -24 35556 3431
rect 35592 -24 35604 863
rect 35616 -24 35628 1895
rect 35664 1285 35676 4127
rect 35760 3325 35772 4103
rect 35640 -24 35652 1271
rect 35688 -24 35700 863
rect 35712 -24 35724 1967
rect 35736 -24 35748 3311
rect 35784 -24 35796 863
rect 35808 -24 35820 3767
rect 35856 2245 35868 4079
rect 35952 2869 35964 4055
rect 35832 -24 35844 2231
rect 35880 -24 35892 863
rect 35904 -24 35916 311
rect 35928 -24 35940 2855
rect 35976 -24 35988 4055
rect 36048 1813 36060 4055
rect 36144 2725 36156 4031
rect 36000 -24 36012 215
rect 36024 -24 36036 1799
rect 36072 -24 36084 119
rect 36120 -24 36132 2711
rect 36192 -24 36204 719
rect 36216 -24 36228 1703
rect 36264 1189 36276 4007
rect 36240 -24 36252 1175
rect 36288 -24 36300 4007
rect 36312 -24 36324 1127
rect 36360 421 36372 4007
rect 41160 3973 41172 4007
rect 59040 3973 59052 4007
rect 59760 3973 59772 4007
rect 36336 -24 36348 407
rect 36384 -24 36396 407
rect 36408 -24 36420 2783
rect 36456 1669 36468 3959
rect 36552 3133 36564 3935
rect 36432 -24 36444 1655
rect 36480 -24 36492 1295
rect 36528 -24 36540 3119
rect 36672 2557 36684 3911
rect 36600 -24 36612 863
rect 36648 -24 36660 2543
rect 36792 1837 36804 3887
rect 36888 2605 36900 3863
rect 36720 -24 36732 407
rect 36744 -24 36756 1415
rect 36768 -24 36780 1823
rect 36816 -24 36828 407
rect 36840 -24 36852 623
rect 36864 -24 36876 2591
rect 36912 -24 36924 3863
rect 36936 -24 36948 1127
rect 36960 -24 36972 2639
rect 37032 1525 37044 3863
rect 36984 -24 36996 1031
rect 37008 -24 37020 1511
rect 37056 -24 37068 3863
rect 37128 3397 37140 3863
rect 37080 -24 37092 839
rect 37104 -24 37116 3383
rect 37152 -24 37164 3863
rect 37224 2677 37236 3863
rect 37176 -24 37188 839
rect 37200 -24 37212 2663
rect 37248 -24 37260 1463
rect 37344 613 37356 3839
rect 37272 -24 37284 -1
rect 37320 -24 37332 599
rect 37368 -24 37380 2471
rect 37392 -24 37404 3839
rect 37464 397 37476 3839
rect 37440 -24 37452 383
rect 37488 -24 37500 3839
rect 37512 -24 37524 3767
rect 37584 1213 37596 3839
rect 37560 -24 37572 1199
rect 37608 -24 37620 1895
rect 37632 -24 37644 1847
rect 37680 1453 37692 3815
rect 37656 -24 37668 1439
rect 37704 -24 37716 2207
rect 37728 -24 37740 3815
rect 37776 1381 37788 3815
rect 37752 -24 37764 1367
rect 37824 781 37836 1247
rect 37800 -24 37812 767
rect 37824 -24 37836 767
rect 37848 -24 37860 2735
rect 37872 1261 37884 3791
rect 37896 -24 37908 2735
rect 37920 -24 37932 2711
rect 37968 661 37980 3767
rect 37944 -24 37956 647
rect 37992 -24 38004 2015
rect 38016 -24 38028 191
rect 38040 -24 38052 3143
rect 38088 1237 38100 3743
rect 38064 -24 38076 1223
rect 38112 -24 38124 3743
rect 38184 1741 38196 3743
rect 59760 3733 59772 3767
rect 38304 2341 38316 3719
rect 38160 -24 38172 1727
rect 38232 -24 38244 407
rect 38256 -24 38268 1895
rect 38280 -24 38292 2327
rect 38328 -24 38340 2711
rect 38424 2101 38436 3695
rect 38352 -24 38364 1871
rect 38400 -24 38412 2087
rect 38448 -24 38460 815
rect 38520 301 38532 3671
rect 38496 -24 38508 287
rect 38568 -24 38580 719
rect 38592 -24 38604 1535
rect 38664 85 38676 3647
rect 38760 2509 38772 3623
rect 38640 -24 38652 71
rect 38688 -24 38700 407
rect 38712 -24 38724 263
rect 38736 -24 38748 2495
rect 38784 -24 38796 2711
rect 38808 -24 38820 647
rect 38856 133 38868 3599
rect 38832 -24 38844 119
rect 38880 -24 38892 3599
rect 38904 -24 38916 3623
rect 38952 2461 38964 3623
rect 38928 -24 38940 2447
rect 38976 -24 38988 575
rect 39000 -24 39012 1415
rect 39048 1309 39060 3599
rect 39024 -24 39036 1295
rect 39072 -24 39084 1295
rect 39096 -24 39108 3455
rect 39168 877 39180 3575
rect 39144 -24 39156 863
rect 39192 -24 39204 3575
rect 39216 -24 39228 3599
rect 39264 3013 39276 3599
rect 39240 -24 39252 2999
rect 39288 -24 39300 3599
rect 39360 3061 39372 3599
rect 39456 3517 39468 3575
rect 39312 -24 39324 215
rect 39336 -24 39348 3047
rect 39384 -24 39396 575
rect 39408 -24 39420 839
rect 39432 -24 39444 3503
rect 39480 -24 39492 3575
rect 39504 -24 39516 3599
rect 39552 445 39564 3599
rect 39528 -24 39540 431
rect 39576 -24 39588 1703
rect 39600 -24 39612 3599
rect 39648 1093 39660 3599
rect 39624 -24 39636 1079
rect 39672 -24 39684 3599
rect 39696 -24 39708 3623
rect 39768 493 39780 3623
rect 39744 -24 39756 479
rect 39792 -24 39804 3623
rect 39816 -24 39828 2543
rect 39864 2101 39876 3623
rect 39840 -24 39852 2087
rect 39888 -24 39900 3623
rect 39960 2821 39972 3623
rect 39912 -24 39924 2639
rect 39936 -24 39948 2807
rect 40056 2293 40068 3599
rect 39984 -24 39996 1055
rect 40008 -24 40020 1511
rect 40032 -24 40044 2279
rect 40080 -24 40092 1511
rect 40152 877 40164 3575
rect 40104 -24 40116 647
rect 40128 -24 40140 863
rect 40176 -24 40188 3575
rect 40248 3325 40260 3575
rect 40200 -24 40212 839
rect 40224 -24 40236 3311
rect 40272 -24 40284 3575
rect 40344 2869 40356 3575
rect 40296 -24 40308 1247
rect 40320 -24 40332 2855
rect 40368 -24 40380 3575
rect 40392 -24 40404 3599
rect 40440 3541 40452 3599
rect 40416 -24 40428 3527
rect 40464 -24 40476 3599
rect 40488 -24 40500 3623
rect 40560 1741 40572 3623
rect 40512 -24 40524 359
rect 40536 -24 40548 1727
rect 40584 -24 40596 3623
rect 40656 3133 40668 3623
rect 40608 -24 40620 1967
rect 40632 -24 40644 3119
rect 40680 -24 40692 1751
rect 40704 -24 40716 1055
rect 40776 85 40788 3599
rect 40752 -24 40764 71
rect 40800 -24 40812 3599
rect 40872 2509 40884 3599
rect 40824 -24 40836 623
rect 40848 -24 40860 2495
rect 40896 -24 40908 3455
rect 40920 -24 40932 1031
rect 40992 829 41004 3575
rect 40968 -24 40980 815
rect 41016 -24 41028 3575
rect 41040 -24 41052 3599
rect 41088 1813 41100 3599
rect 41064 -24 41076 1799
rect 41112 -24 41124 767
rect 41160 -24 41172 3599
rect 41232 -24 41244 3599
rect 41304 1285 41316 3599
rect 41256 -24 41268 1055
rect 41280 -24 41292 1271
rect 41328 -24 41340 3599
rect 41400 2629 41412 3599
rect 41352 -24 41364 263
rect 41376 -24 41388 2615
rect 41424 -24 41436 2447
rect 41496 733 41508 3575
rect 41472 -24 41484 719
rect 41544 -24 41556 2615
rect 41616 2605 41628 3551
rect 41568 -24 41580 1127
rect 41592 -24 41604 2591
rect 41640 -24 41652 2207
rect 41664 -24 41676 3551
rect 41712 2173 41724 3551
rect 41688 -24 41700 2159
rect 41736 -24 41748 3551
rect 41808 2773 41820 3551
rect 41760 -24 41772 2063
rect 41784 -24 41796 2759
rect 41832 -24 41844 3551
rect 41856 -24 41868 3575
rect 41904 2485 41916 3575
rect 41880 -24 41892 2471
rect 42000 1381 42012 3551
rect 41928 -24 41940 935
rect 41952 -24 41964 1007
rect 41976 -24 41988 1367
rect 42024 -24 42036 3551
rect 42120 1213 42132 3551
rect 42048 -24 42060 47
rect 42096 -24 42108 1199
rect 42144 -24 42156 695
rect 42216 541 42228 3527
rect 42336 2437 42348 3503
rect 59040 3493 59052 3527
rect 59640 3493 59652 3527
rect 59760 3493 59772 3527
rect 42192 -24 42204 527
rect 42264 -24 42276 1271
rect 42312 -24 42324 2423
rect 42456 1237 42468 3479
rect 42384 -24 42396 431
rect 42432 -24 42444 1223
rect 42504 -24 42516 2543
rect 42528 -24 42540 167
rect 42552 -24 42564 2975
rect 42600 1645 42612 3455
rect 42576 -24 42588 1631
rect 42624 -24 42636 1751
rect 42696 421 42708 3431
rect 42816 2725 42828 3407
rect 42672 -24 42684 407
rect 42744 -24 42756 1079
rect 42792 -24 42804 2711
rect 42864 -24 42876 2615
rect 42936 2605 42948 3383
rect 42888 -24 42900 791
rect 42912 -24 42924 2591
rect 42960 -24 42972 2615
rect 43056 2005 43068 3359
rect 42984 -24 42996 1415
rect 43032 -24 43044 1991
rect 43152 1861 43164 3335
rect 43080 -24 43092 1511
rect 43128 -24 43140 1847
rect 43200 -24 43212 3335
rect 43272 781 43284 3335
rect 43224 -24 43236 215
rect 43248 -24 43260 767
rect 43296 -24 43308 2207
rect 43320 -24 43332 3335
rect 43368 2605 43380 3335
rect 43344 -24 43356 2591
rect 43392 -24 43404 3335
rect 43416 -24 43428 3359
rect 43464 2677 43476 3359
rect 43440 -24 43452 2663
rect 43488 -24 43500 2903
rect 43512 -24 43524 2903
rect 43560 2845 43572 3335
rect 43536 -24 43548 2831
rect 43584 -24 43596 1487
rect 43608 -24 43620 3335
rect 43656 1477 43668 3335
rect 43632 -24 43644 1463
rect 43680 -24 43692 2735
rect 43752 1189 43764 3311
rect 43872 2749 43884 3287
rect 43728 -24 43740 1175
rect 43800 -24 43812 2567
rect 43824 -24 43836 1343
rect 43848 -24 43860 2735
rect 43968 2245 43980 3263
rect 43896 -24 43908 1703
rect 43920 -24 43932 479
rect 43944 -24 43956 2231
rect 43992 -24 44004 3263
rect 44016 -24 44028 3287
rect 44064 2101 44076 3287
rect 44040 -24 44052 2087
rect 44088 -24 44100 791
rect 44112 -24 44124 455
rect 44136 -24 44148 2687
rect 44184 1789 44196 3263
rect 58920 3253 58932 3287
rect 59040 3253 59052 3287
rect 59640 3253 59652 3287
rect 59760 3253 59772 3287
rect 44352 2821 44364 3239
rect 44160 -24 44172 1775
rect 44232 -24 44244 1847
rect 44256 -24 44268 743
rect 44304 -24 44316 1535
rect 44328 -24 44340 2807
rect 44400 -24 44412 3239
rect 44472 3133 44484 3239
rect 44424 -24 44436 1847
rect 44448 -24 44460 3119
rect 44496 -24 44508 2615
rect 44568 2365 44580 3215
rect 44544 -24 44556 2351
rect 44616 -24 44628 2807
rect 44640 -24 44652 2975
rect 44712 397 44724 3191
rect 44808 1813 44820 3167
rect 44688 -24 44700 383
rect 44736 -24 44748 1415
rect 44760 -24 44772 143
rect 44784 -24 44796 1799
rect 44832 -24 44844 1439
rect 44856 -24 44868 1007
rect 44904 709 44916 3143
rect 44880 -24 44892 695
rect 44928 -24 44940 1871
rect 44952 -24 44964 2807
rect 45000 1645 45012 3119
rect 44976 -24 44988 1631
rect 45024 -24 45036 143
rect 45048 -24 45060 2807
rect 45120 1285 45132 3095
rect 45096 -24 45108 1271
rect 45144 -24 45156 1295
rect 45216 589 45228 3071
rect 45336 2413 45348 3047
rect 45192 -24 45204 575
rect 45264 -24 45276 719
rect 45312 -24 45324 2399
rect 45384 -24 45396 1439
rect 45408 -24 45420 2135
rect 45456 445 45468 3023
rect 59640 3013 59652 3047
rect 59760 3013 59772 3047
rect 45432 -24 45444 431
rect 45480 -24 45492 167
rect 45504 -24 45516 647
rect 45552 613 45564 2999
rect 45648 2413 45660 2975
rect 45528 -24 45540 599
rect 45576 -24 45588 767
rect 45624 -24 45636 2399
rect 45768 1693 45780 2951
rect 45696 -24 45708 455
rect 45720 -24 45732 1415
rect 45744 -24 45756 1679
rect 45792 -24 45804 1415
rect 45816 -24 45828 2951
rect 45864 445 45876 2951
rect 45840 -24 45852 431
rect 45888 -24 45900 2951
rect 45960 1813 45972 2951
rect 46056 2461 46068 2927
rect 45912 -24 45924 1415
rect 45936 -24 45948 1799
rect 45984 -24 45996 1319
rect 46008 -24 46020 1127
rect 46032 -24 46044 2447
rect 46080 -24 46092 2927
rect 46104 -24 46116 1127
rect 46152 973 46164 2927
rect 46248 1765 46260 2903
rect 46128 -24 46140 959
rect 46176 -24 46188 959
rect 46200 -24 46212 215
rect 46224 -24 46236 1751
rect 46272 -24 46284 455
rect 46296 -24 46308 1127
rect 46368 109 46380 2879
rect 46464 829 46476 2855
rect 46344 -24 46356 95
rect 46392 -24 46404 311
rect 46416 -24 46428 167
rect 46440 -24 46452 815
rect 46488 -24 46500 2855
rect 46560 2509 46572 2855
rect 46512 -24 46524 239
rect 46536 -24 46548 2495
rect 46584 -24 46596 1631
rect 46608 -24 46620 671
rect 46680 205 46692 2831
rect 46656 -24 46668 191
rect 46704 -24 46716 2831
rect 46728 -24 46740 1535
rect 46752 -24 46764 2639
rect 46824 2341 46836 2831
rect 46776 -24 46788 695
rect 46800 -24 46812 2327
rect 46848 -24 46860 2831
rect 46872 -24 46884 2855
rect 46896 -24 46908 2879
rect 46944 829 46956 2879
rect 46920 -24 46932 815
rect 46968 -24 46980 2567
rect 47064 2293 47076 2855
rect 46992 -24 47004 2015
rect 47040 -24 47052 2279
rect 47088 -24 47100 2855
rect 47112 -24 47124 1895
rect 47160 997 47172 2855
rect 47136 -24 47148 983
rect 47184 -24 47196 983
rect 47208 -24 47220 1871
rect 47256 1189 47268 2831
rect 47232 -24 47244 1175
rect 47280 -24 47292 2015
rect 47304 -24 47316 1967
rect 47376 541 47388 2807
rect 47472 1093 47484 2783
rect 47328 -24 47340 335
rect 47352 -24 47364 527
rect 47400 -24 47412 527
rect 47424 -24 47436 1031
rect 47448 -24 47460 1079
rect 47496 -24 47508 2783
rect 47520 -24 47532 2807
rect 47544 -24 47556 2831
rect 47592 1525 47604 2831
rect 47712 2269 47724 2807
rect 47568 -24 47580 1511
rect 47616 -24 47628 215
rect 47640 -24 47652 239
rect 47664 -24 47676 1055
rect 47688 -24 47700 2255
rect 47736 -24 47748 2807
rect 47832 1213 47844 2807
rect 47760 -24 47772 1031
rect 47808 -24 47820 1199
rect 47880 -24 47892 1871
rect 47904 -24 47916 647
rect 47952 -24 47964 2807
rect 48000 2605 48012 2807
rect 47976 -24 47988 2591
rect 48120 2125 48132 2783
rect 59640 2773 59652 2807
rect 59760 2773 59772 2807
rect 48048 -24 48060 551
rect 48096 -24 48108 2111
rect 48168 -24 48180 2231
rect 48264 1957 48276 2759
rect 48384 2629 48396 2735
rect 48192 -24 48204 215
rect 48240 -24 48252 1943
rect 48288 -24 48300 239
rect 48312 -24 48324 215
rect 48360 -24 48372 2615
rect 48408 -24 48420 2735
rect 48432 -24 48444 1871
rect 48480 1741 48492 2735
rect 48456 -24 48468 1727
rect 48504 -24 48516 239
rect 48528 -24 48540 215
rect 48576 205 48588 2711
rect 48552 -24 48564 191
rect 48600 -24 48612 2639
rect 48624 -24 48636 2543
rect 48672 901 48684 2687
rect 48648 -24 48660 887
rect 48696 -24 48708 839
rect 48720 -24 48732 2687
rect 48768 205 48780 2687
rect 48864 2389 48876 2663
rect 48744 -24 48756 191
rect 48792 -24 48804 1703
rect 48816 -24 48828 191
rect 48840 -24 48852 2375
rect 48888 -24 48900 1319
rect 48912 -24 48924 1535
rect 48960 1309 48972 2639
rect 48936 -24 48948 1295
rect 48984 -24 48996 263
rect 49008 -24 49020 1703
rect 49056 733 49068 2615
rect 49032 -24 49044 719
rect 49080 -24 49092 2615
rect 49152 1933 49164 2615
rect 49248 2197 49260 2591
rect 49104 -24 49116 1703
rect 49128 -24 49140 1919
rect 49176 -24 49188 1727
rect 49200 -24 49212 815
rect 49224 -24 49236 2183
rect 49272 -24 49284 2327
rect 49344 877 49356 2567
rect 49296 -24 49308 647
rect 49320 -24 49332 863
rect 49368 -24 49380 2255
rect 49392 -24 49404 2111
rect 49440 1477 49452 2543
rect 49416 -24 49428 1463
rect 49464 -24 49476 2087
rect 49536 1381 49548 2519
rect 49488 -24 49500 335
rect 49512 -24 49524 1367
rect 49560 -24 49572 1295
rect 49632 1237 49644 2495
rect 49728 1693 49740 2471
rect 49584 -24 49596 -1
rect 49608 -24 49620 1223
rect 49656 -24 49668 1295
rect 49680 -24 49692 47
rect 49704 -24 49716 1679
rect 49752 -24 49764 2231
rect 49848 781 49860 2447
rect 49776 -24 49788 263
rect 49824 -24 49836 767
rect 49872 -24 49884 1199
rect 49896 -24 49908 2087
rect 49968 949 49980 2423
rect 49944 -24 49956 935
rect 49992 -24 50004 2423
rect 50016 -24 50028 2447
rect 50064 2173 50076 2447
rect 50040 -24 50052 2159
rect 50088 -24 50100 2279
rect 50160 1957 50172 2423
rect 50112 -24 50124 1175
rect 50136 -24 50148 1943
rect 50184 -24 50196 1727
rect 50208 -24 50220 671
rect 50256 421 50268 2399
rect 50232 -24 50244 407
rect 50280 -24 50292 287
rect 50304 -24 50316 1895
rect 50352 1837 50364 2375
rect 50328 -24 50340 1823
rect 50448 -24 50460 935
rect 50832 613 50844 2351
rect 50880 1765 50892 2327
rect 50808 -24 50820 599
rect 50856 -24 50868 1751
rect 51000 -24 51012 191
rect 51024 -24 51036 2327
rect 51072 1285 51084 2327
rect 51168 2005 51180 2303
rect 51048 -24 51060 1271
rect 51096 -24 51108 455
rect 51120 -24 51132 839
rect 51144 -24 51156 1991
rect 51192 -24 51204 1607
rect 51216 -24 51228 2303
rect 51264 1837 51276 2303
rect 59520 2293 59532 2327
rect 59640 2293 59652 2327
rect 59760 2293 59772 2327
rect 59880 2293 59892 2327
rect 51240 -24 51252 1823
rect 51288 -24 51300 1463
rect 51312 -24 51324 1703
rect 51336 -24 51348 407
rect 51384 109 51396 2279
rect 51360 -24 51372 95
rect 51408 -24 51420 1607
rect 51432 -24 51444 1463
rect 51504 997 51516 2255
rect 51600 1141 51612 2231
rect 51480 -24 51492 983
rect 51528 -24 51540 263
rect 51576 -24 51588 1127
rect 51648 -24 51660 1871
rect 51672 -24 51684 2231
rect 51720 1789 51732 2231
rect 51696 -24 51708 1775
rect 51744 -24 51756 1967
rect 51768 -24 51780 1895
rect 51792 -24 51804 2207
rect 51864 1117 51876 2207
rect 51816 -24 51828 1007
rect 51840 -24 51852 1103
rect 51888 -24 51900 1703
rect 51912 -24 51924 2063
rect 51984 877 51996 2183
rect 51960 -24 51972 863
rect 52008 -24 52020 1463
rect 52032 -24 52044 1703
rect 52056 -24 52068 1247
rect 52104 85 52116 2159
rect 52200 541 52212 2135
rect 52320 973 52332 2111
rect 52440 1645 52452 2087
rect 52080 -24 52092 71
rect 52128 -24 52140 191
rect 52176 -24 52188 527
rect 52248 -24 52260 239
rect 52296 -24 52308 959
rect 52368 -24 52380 743
rect 52416 -24 52428 1631
rect 52488 -24 52500 431
rect 52560 325 52572 2063
rect 59400 2053 59412 2087
rect 59520 2053 59532 2087
rect 59640 2053 59652 2087
rect 59760 2053 59772 2087
rect 59880 2053 59892 2087
rect 52536 -24 52548 311
rect 52608 -24 52620 791
rect 52632 -24 52644 1535
rect 52680 133 52692 2039
rect 52656 -24 52668 119
rect 52704 -24 52716 623
rect 52728 -24 52740 791
rect 52800 565 52812 2015
rect 52896 1429 52908 1991
rect 52776 -24 52788 551
rect 52824 -24 52836 1079
rect 52872 -24 52884 1415
rect 52944 -24 52956 1631
rect 53016 1453 53028 1967
rect 53136 1573 53148 1943
rect 52992 -24 53004 1439
rect 53064 -24 53076 47
rect 53088 -24 53100 407
rect 53112 -24 53124 1559
rect 53160 -24 53172 1391
rect 53232 181 53244 1919
rect 53208 -24 53220 167
rect 53280 -24 53292 407
rect 53304 -24 53316 1007
rect 53328 -24 53340 1031
rect 53376 493 53388 1895
rect 53472 1237 53484 1871
rect 53352 -24 53364 479
rect 53400 -24 53412 455
rect 53448 -24 53460 1223
rect 53592 1093 53604 1847
rect 53544 853 53556 1055
rect 53520 -24 53532 839
rect 53544 -24 53556 839
rect 53568 -24 53580 1055
rect 53616 -24 53628 1583
rect 53640 1093 53652 1823
rect 53664 1597 53676 1799
rect 53640 -24 53652 911
rect 53664 -24 53676 1175
rect 53688 925 53700 1775
rect 53712 1189 53724 1751
rect 53712 -24 53724 863
rect 53784 709 53796 1727
rect 53760 -24 53772 695
rect 53832 -24 53844 551
rect 53856 -24 53868 1007
rect 53904 205 53916 1703
rect 53880 -24 53892 191
rect 53928 -24 53940 359
rect 54000 181 54012 1679
rect 54096 493 54108 1655
rect 53976 -24 53988 167
rect 54072 133 54084 479
rect 54120 277 54132 1631
rect 54048 -24 54060 119
rect 54072 -24 54084 119
rect 54096 -24 54108 263
rect 54144 -24 54156 1151
rect 54216 997 54228 1607
rect 54264 1429 54276 1583
rect 54168 -24 54180 671
rect 54192 -24 54204 983
rect 54240 -24 54252 1415
rect 54288 589 54300 1559
rect 54264 -24 54276 575
rect 54312 109 54324 1535
rect 54288 -24 54300 95
rect 54336 -24 54348 1415
rect 54408 301 54420 1511
rect 54552 469 54564 1487
rect 54672 1333 54684 1463
rect 54384 -24 54396 287
rect 54456 -24 54468 191
rect 54480 -24 54492 215
rect 54528 -24 54540 455
rect 54576 -24 54588 215
rect 54600 -24 54612 143
rect 54648 -24 54660 1319
rect 54792 1189 54804 1439
rect 54696 -24 54708 1007
rect 54720 -24 54732 -1
rect 54768 -24 54780 1175
rect 54816 -24 54828 1319
rect 54840 -24 54852 647
rect 54888 445 54900 1415
rect 54864 -24 54876 431
rect 54912 -24 54924 1319
rect 54984 517 54996 1391
rect 54936 -24 54948 407
rect 54960 -24 54972 503
rect 55008 -24 55020 1223
rect 55080 1213 55092 1367
rect 55032 -24 55044 -1
rect 55056 -24 55068 1199
rect 55104 -24 55116 1199
rect 55152 -24 55164 1343
rect 55296 1141 55308 1319
rect 55224 -24 55236 191
rect 55248 -24 55260 143
rect 55272 -24 55284 1127
rect 55320 -24 55332 143
rect 55344 -24 55356 1223
rect 55392 -24 55404 1295
rect 55440 -24 55452 95
rect 55464 -24 55476 1127
rect 55536 709 55548 1271
rect 55512 -24 55524 695
rect 55560 -24 55572 911
rect 55632 397 55644 1247
rect 55608 -24 55620 383
rect 55680 -24 55692 551
rect 55704 -24 55716 527
rect 55752 517 55764 1223
rect 55728 -24 55740 503
rect 55776 -24 55788 1175
rect 55848 277 55860 1199
rect 55800 -24 55812 -1
rect 55824 -24 55836 263
rect 55872 -24 55884 1127
rect 55944 181 55956 1175
rect 55896 -24 55908 -1
rect 55920 -24 55932 167
rect 56040 -24 56052 1175
rect 56472 949 56484 1175
rect 56448 -24 56460 935
rect 56664 829 56676 1151
rect 56640 733 56652 815
rect 56688 781 56700 1127
rect 56592 -24 56604 671
rect 56616 -24 56628 719
rect 56640 -24 56652 719
rect 56664 -24 56676 767
rect 56712 -24 56724 1055
rect 56784 973 56796 1103
rect 56736 -24 56748 719
rect 56760 -24 56772 959
rect 56880 757 56892 1079
rect 56808 -24 56820 455
rect 56832 -24 56844 719
rect 56856 -24 56868 743
rect 56976 349 56988 1055
rect 57096 589 57108 1031
rect 56904 -24 56916 71
rect 56952 -24 56964 335
rect 57024 -24 57036 503
rect 57048 -24 57060 527
rect 57072 -24 57084 575
rect 57120 -24 57132 95
rect 57144 -24 57156 143
rect 57168 -24 57180 239
rect 57192 157 57204 1007
rect 57216 253 57228 959
rect 57288 493 57300 959
rect 57216 -24 57228 239
rect 57240 -24 57252 167
rect 57264 -24 57276 479
rect 57336 205 57348 239
rect 57312 -24 57324 191
rect 57336 -24 57348 191
rect 57360 -24 57372 599
rect 57384 253 57396 935
rect 57408 613 57420 911
rect 57408 -24 57420 527
rect 57432 -24 57444 647
rect 57480 613 57492 887
rect 57456 -24 57468 599
rect 57504 -24 57516 839
rect 57600 805 57612 863
rect 57528 -24 57540 119
rect 57576 -24 57588 791
rect 57696 373 57708 839
rect 57624 -24 57636 191
rect 57648 -24 57660 215
rect 57672 -24 57684 359
rect 57720 -24 57732 719
rect 57744 -24 57756 671
rect 57816 325 57828 815
rect 57864 373 57876 791
rect 57792 -24 57804 311
rect 57840 -24 57852 359
rect 57888 133 57900 767
rect 57936 637 57948 743
rect 57864 -24 57876 119
rect 57912 -24 57924 623
rect 57960 -24 57972 527
rect 57984 -24 57996 -1
rect 58008 -24 58020 695
rect 58056 -24 58068 647
rect 58080 -24 58092 383
rect 58128 277 58140 695
rect 58104 -24 58116 263
rect 58152 -24 58164 527
rect 58176 -24 58188 575
rect 58224 85 58236 671
rect 58200 -24 58212 71
rect 58248 -24 58260 383
rect 58320 301 58332 647
rect 58272 -24 58284 71
rect 58296 -24 58308 287
rect 58392 229 58404 623
rect 58440 445 58452 599
rect 58344 -24 58356 191
rect 58368 -24 58380 215
rect 58416 -24 58428 431
rect 58464 -24 58476 575
rect 58488 -24 58500 527
rect 58560 61 58572 575
rect 58656 373 58668 551
rect 58536 -24 58548 47
rect 58584 -24 58596 47
rect 58608 -24 58620 287
rect 58632 -24 58644 359
rect 58680 -24 58692 95
rect 58704 -24 58716 191
rect 58728 109 58740 527
rect 58752 -24 58764 479
rect 58776 205 58788 479
rect 58800 397 58812 479
rect 58824 397 58836 455
rect 58872 397 58884 431
rect 58800 -24 58812 383
rect 58848 -24 58860 383
rect 58920 85 58932 431
rect 58944 85 58956 407
rect 58992 349 59004 383
rect 59040 349 59052 383
rect 58920 -24 58932 71
rect 58968 -24 58980 335
rect 59040 -24 59052 335
rect 59112 229 59124 335
rect 59160 301 59172 335
rect 59088 -24 59100 215
rect 59160 -24 59172 287
rect 59232 181 59244 287
rect 59208 -24 59220 167
rect 59280 85 59292 287
rect 59304 85 59316 263
rect 59352 205 59364 239
rect 59280 -24 59292 71
rect 59328 -24 59340 191
rect 59400 61 59412 239
rect 59424 61 59436 215
rect 59472 133 59484 191
rect 59400 -24 59412 47
rect 59448 -24 59460 119
rect 59520 37 59532 191
rect 59544 37 59556 167
rect 59592 61 59604 143
rect 59640 85 59652 143
rect 59664 85 59676 119
rect 59520 -24 59532 -1
rect 59568 -24 59580 47
rect 59640 -24 59652 71
rect 59712 37 59724 95
rect 59688 -24 59700 -1
rect 59760 -24 59772 95
rect 59808 -24 59820 71
rect 59880 37 59892 71
rect 59880 -24 59892 -1
rect 59928 -24 59940 -1
use scandtype StatusReg_reg_0
timestamp 1386241841
transform 1 0 24 0 1 -823
box 0 0 624 799
use scandtype StatusReg_reg_1
timestamp 1386241841
transform 1 0 648 0 1 -823
box 0 0 624 799
use scandtype StatusReg_reg_2
timestamp 1386241841
transform 1 0 1272 0 1 -823
box 0 0 624 799
use scandtype StatusReg_reg_3
timestamp 1386241841
transform 1 0 1896 0 1 -823
box 0 0 624 799
use nand2 g11910
timestamp 1386234792
transform 1 0 2520 0 1 -823
box 0 0 96 799
use nand3 g11904
timestamp 1386234893
transform 1 0 2616 0 1 -823
box 0 0 120 799
use nand4 g11889
timestamp 1386234936
transform 1 0 2736 0 1 -823
box 0 0 144 799
use nand4 g11898
timestamp 1386234936
transform 1 0 2880 0 1 -823
box 0 0 144 799
use nand4 g11888
timestamp 1386234936
transform 1 0 3024 0 1 -823
box 0 0 144 799
use nand2 g11922
timestamp 1386234792
transform 1 0 3168 0 1 -823
box 0 0 96 799
use nand2 g11930
timestamp 1386234792
transform 1 0 3264 0 1 -823
box 0 0 96 799
use nand3 g11905
timestamp 1386234893
transform 1 0 3360 0 1 -823
box 0 0 120 799
use scandtype stateSub_reg_0
timestamp 1386241841
transform 1 0 3480 0 1 -823
box 0 0 624 799
use scandtype InISR_reg
timestamp 1386241841
transform 1 0 4104 0 1 -823
box 0 0 624 799
use nand3 g11909
timestamp 1386234893
transform 1 0 4728 0 1 -823
box 0 0 120 799
use nand4 g11925
timestamp 1386234936
transform 1 0 4848 0 1 -823
box 0 0 144 799
use nand3 g11902
timestamp 1386234893
transform 1 0 4992 0 1 -823
box 0 0 120 799
use nand3 g11900
timestamp 1386234893
transform 1 0 5112 0 1 -823
box 0 0 120 799
use nand3 g11903
timestamp 1386234893
transform 1 0 5232 0 1 -823
box 0 0 120 799
use nand2 g11957
timestamp 1386234792
transform 1 0 5352 0 1 -823
box 0 0 96 799
use nand4 g11906
timestamp 1386234936
transform 1 0 5448 0 1 -823
box 0 0 144 799
use nand2 g11921
timestamp 1386234792
transform 1 0 5592 0 1 -823
box 0 0 96 799
use nand4 g11911
timestamp 1386234936
transform 1 0 5688 0 1 -823
box 0 0 144 799
use nor2 g11907
timestamp 1386235306
transform 1 0 5832 0 1 -823
box 0 0 120 799
use nor2 g11931
timestamp 1386235306
transform 1 0 5952 0 1 -823
box 0 0 120 799
use nand2 g11914
timestamp 1386234792
transform 1 0 6072 0 1 -823
box 0 0 96 799
use nand2 g11916
timestamp 1386234792
transform 1 0 6168 0 1 -823
box 0 0 96 799
use and2 g11939
timestamp 1386234845
transform 1 0 6264 0 1 -823
box 0 0 120 799
use nand2 g11915
timestamp 1386234792
transform 1 0 6384 0 1 -823
box 0 0 96 799
use scandtype state_reg_0
timestamp 1386241841
transform 1 0 6480 0 1 -823
box 0 0 624 799
use scandtype state_reg_1
timestamp 1386241841
transform 1 0 7104 0 1 -823
box 0 0 624 799
use nand2 g11913
timestamp 1386234792
transform 1 0 7728 0 1 -823
box 0 0 96 799
use nand4 g11942
timestamp 1386234936
transform 1 0 7824 0 1 -823
box 0 0 144 799
use nand3 g11973
timestamp 1386234893
transform 1 0 7968 0 1 -823
box 0 0 120 799
use nand3 g11947
timestamp 1386234893
transform 1 0 8088 0 1 -823
box 0 0 120 799
use nand2 g11943
timestamp 1386234792
transform 1 0 8208 0 1 -823
box 0 0 96 799
use nor2 g11894
timestamp 1386235306
transform 1 0 8304 0 1 -823
box 0 0 120 799
use nand2 g11945
timestamp 1386234792
transform 1 0 8424 0 1 -823
box 0 0 96 799
use nand4 g11946
timestamp 1386234936
transform 1 0 8520 0 1 -823
box 0 0 144 799
use nand2 g11968
timestamp 1386234792
transform 1 0 8664 0 1 -823
box 0 0 96 799
use nand2 g11926
timestamp 1386234792
transform 1 0 8760 0 1 -823
box 0 0 96 799
use nand2 g11927
timestamp 1386234792
transform 1 0 8856 0 1 -823
box 0 0 96 799
use nand2 g11970
timestamp 1386234792
transform 1 0 8952 0 1 -823
box 0 0 96 799
use nand2 g11928
timestamp 1386234792
transform 1 0 9048 0 1 -823
box 0 0 96 799
use nand2 g11971
timestamp 1386234792
transform 1 0 9144 0 1 -823
box 0 0 96 799
use nand2 g11929
timestamp 1386234792
transform 1 0 9240 0 1 -823
box 0 0 96 799
use nand2 g11972
timestamp 1386234792
transform 1 0 9336 0 1 -823
box 0 0 96 799
use nand3 g11932
timestamp 1386234893
transform 1 0 9432 0 1 -823
box 0 0 120 799
use inv g11992
timestamp 1386238110
transform 1 0 9552 0 1 -823
box 0 0 120 799
use nand4 g11923
timestamp 1386234936
transform 1 0 9672 0 1 -823
box 0 0 144 799
use nand3 g11912
timestamp 1386234893
transform 1 0 9816 0 1 -823
box 0 0 120 799
use nand4 g11901
timestamp 1386234936
transform 1 0 9936 0 1 -823
box 0 0 144 799
use nand2 g11962
timestamp 1386234792
transform 1 0 10080 0 1 -823
box 0 0 96 799
use inv g11952
timestamp 1386238110
transform 1 0 10176 0 1 -823
box 0 0 120 799
use nor2 g11955
timestamp 1386235306
transform 1 0 10296 0 1 -823
box 0 0 120 799
use nand2 g11967
timestamp 1386234792
transform 1 0 10416 0 1 -823
box 0 0 96 799
use inv g11976
timestamp 1386238110
transform 1 0 10512 0 1 -823
box 0 0 120 799
use nand4 g11908
timestamp 1386234936
transform 1 0 10632 0 1 -823
box 0 0 144 799
use nand4 g11896
timestamp 1386234936
transform 1 0 10776 0 1 -823
box 0 0 144 799
use nand3 g11993
timestamp 1386234893
transform 1 0 10920 0 1 -823
box 0 0 120 799
use nand4 g11917
timestamp 1386234936
transform 1 0 11040 0 1 -823
box 0 0 144 799
use nand2 g11941
timestamp 1386234792
transform 1 0 11184 0 1 -823
box 0 0 96 799
use nand4 g11948
timestamp 1386234936
transform 1 0 11280 0 1 -823
box 0 0 144 799
use nand2 g11964
timestamp 1386234792
transform 1 0 11424 0 1 -823
box 0 0 96 799
use nand4 g11899
timestamp 1386234936
transform 1 0 11520 0 1 -823
box 0 0 144 799
use nand4 g11974
timestamp 1386234936
transform 1 0 11664 0 1 -823
box 0 0 144 799
use nand4 g11897
timestamp 1386234936
transform 1 0 11808 0 1 -823
box 0 0 144 799
use nand4 g11951
timestamp 1386234936
transform 1 0 11952 0 1 -823
box 0 0 144 799
use nand4 g11953
timestamp 1386234936
transform 1 0 12096 0 1 -823
box 0 0 144 799
use nand2 g11954
timestamp 1386234792
transform 1 0 12240 0 1 -823
box 0 0 96 799
use and2 g11958
timestamp 1386234845
transform 1 0 12336 0 1 -823
box 0 0 120 799
use nand2 g11963
timestamp 1386234792
transform 1 0 12456 0 1 -823
box 0 0 96 799
use nand4 g11977
timestamp 1386234936
transform 1 0 12552 0 1 -823
box 0 0 144 799
use nand2 g11983
timestamp 1386234792
transform 1 0 12696 0 1 -823
box 0 0 96 799
use nand2 g11984
timestamp 1386234792
transform 1 0 12792 0 1 -823
box 0 0 96 799
use inv g11985
timestamp 1386238110
transform 1 0 12888 0 1 -823
box 0 0 120 799
use and2 g11988
timestamp 1386234845
transform 1 0 13008 0 1 -823
box 0 0 120 799
use nand2 g11990
timestamp 1386234792
transform 1 0 13128 0 1 -823
box 0 0 96 799
use inv g11995
timestamp 1386238110
transform 1 0 13224 0 1 -823
box 0 0 120 799
use nand2 g11960
timestamp 1386234792
transform 1 0 13344 0 1 -823
box 0 0 96 799
use nand3 g11944
timestamp 1386234893
transform 1 0 13440 0 1 -823
box 0 0 120 799
use and2 g12002
timestamp 1386234845
transform 1 0 13560 0 1 -823
box 0 0 120 799
use inv g12006
timestamp 1386238110
transform 1 0 13680 0 1 -823
box 0 0 120 799
use trisbuf g746
timestamp 1386237216
transform 1 0 13800 0 1 -823
box 0 0 216 799
use trisbuf g738
timestamp 1386237216
transform 1 0 14016 0 1 -823
box 0 0 216 799
use and2 g11981
timestamp 1386234845
transform 1 0 14232 0 1 -823
box 0 0 120 799
use nand2 g11986
timestamp 1386234792
transform 1 0 14352 0 1 -823
box 0 0 96 799
use nand2 g11987
timestamp 1386234792
transform 1 0 14448 0 1 -823
box 0 0 96 799
use nand2 g11937
timestamp 1386234792
transform 1 0 14544 0 1 -823
box 0 0 96 799
use nand2 g11991
timestamp 1386234792
transform 1 0 14640 0 1 -823
box 0 0 96 799
use nand2 g11938
timestamp 1386234792
transform 1 0 14736 0 1 -823
box 0 0 96 799
use nand2 g11996
timestamp 1386234792
transform 1 0 14832 0 1 -823
box 0 0 96 799
use nand2 g11940
timestamp 1386234792
transform 1 0 14928 0 1 -823
box 0 0 96 799
use nand3 g11999
timestamp 1386234893
transform 1 0 15024 0 1 -823
box 0 0 120 799
use trisbuf g742
timestamp 1386237216
transform 1 0 15144 0 1 -823
box 0 0 216 799
use nand3 g12000
timestamp 1386234893
transform 1 0 15360 0 1 -823
box 0 0 120 799
use trisbuf g1
timestamp 1386237216
transform 1 0 15480 0 1 -823
box 0 0 216 799
use trisbuf g734
timestamp 1386237216
transform 1 0 15696 0 1 -823
box 0 0 216 799
use trisbuf g735
timestamp 1386237216
transform 1 0 15912 0 1 -823
box 0 0 216 799
use trisbuf g736
timestamp 1386237216
transform 1 0 16128 0 1 -823
box 0 0 216 799
use trisbuf g737
timestamp 1386237216
transform 1 0 16344 0 1 -823
box 0 0 216 799
use trisbuf g739
timestamp 1386237216
transform 1 0 16560 0 1 -823
box 0 0 216 799
use trisbuf g740
timestamp 1386237216
transform 1 0 16776 0 1 -823
box 0 0 216 799
use trisbuf g741
timestamp 1386237216
transform 1 0 16992 0 1 -823
box 0 0 216 799
use trisbuf g743
timestamp 1386237216
transform 1 0 17208 0 1 -823
box 0 0 216 799
use trisbuf g744
timestamp 1386237216
transform 1 0 17424 0 1 -823
box 0 0 216 799
use trisbuf g745
timestamp 1386237216
transform 1 0 17640 0 1 -823
box 0 0 216 799
use trisbuf g747
timestamp 1386237216
transform 1 0 17856 0 1 -823
box 0 0 216 799
use trisbuf g748
timestamp 1386237216
transform 1 0 18072 0 1 -823
box 0 0 216 799
use nand3 g12004
timestamp 1386234893
transform 1 0 18288 0 1 -823
box 0 0 120 799
use nand3 g12007
timestamp 1386234893
transform 1 0 18408 0 1 -823
box 0 0 120 799
use nand2 g11961
timestamp 1386234792
transform 1 0 18528 0 1 -823
box 0 0 96 799
use nor2 g11924
timestamp 1386235306
transform 1 0 18624 0 1 -823
box 0 0 120 799
use nand2 g12035
timestamp 1386234792
transform 1 0 18744 0 1 -823
box 0 0 96 799
use nand2 g12036
timestamp 1386234792
transform 1 0 18840 0 1 -823
box 0 0 96 799
use and2 g11969
timestamp 1386234845
transform 1 0 18936 0 1 -823
box 0 0 120 799
use nand2 g11997
timestamp 1386234792
transform 1 0 19056 0 1 -823
box 0 0 96 799
use nand2 g12043
timestamp 1386234792
transform 1 0 19152 0 1 -823
box 0 0 96 799
use nor2 g11933
timestamp 1386235306
transform 1 0 19248 0 1 -823
box 0 0 120 799
use nor2 g11982
timestamp 1386235306
transform 1 0 19368 0 1 -823
box 0 0 120 799
use inv g11935
timestamp 1386238110
transform 1 0 19488 0 1 -823
box 0 0 120 799
use and2 g11994
timestamp 1386234845
transform 1 0 19608 0 1 -823
box 0 0 120 799
use scandtype stateSub_reg_2
timestamp 1386241841
transform 1 0 19728 0 1 -823
box 0 0 624 799
use nand2 g12020
timestamp 1386234792
transform 1 0 20352 0 1 -823
box 0 0 96 799
use nand3 g12005
timestamp 1386234893
transform 1 0 20448 0 1 -823
box 0 0 120 799
use inv g11949
timestamp 1386238110
transform 1 0 20568 0 1 -823
box 0 0 120 799
use nand2 g12014
timestamp 1386234792
transform 1 0 20688 0 1 -823
box 0 0 96 799
use nand2 g12015
timestamp 1386234792
transform 1 0 20784 0 1 -823
box 0 0 96 799
use nand2 g12017
timestamp 1386234792
transform 1 0 20880 0 1 -823
box 0 0 96 799
use nand2 g12018
timestamp 1386234792
transform 1 0 20976 0 1 -823
box 0 0 96 799
use nand2 g12022
timestamp 1386234792
transform 1 0 21072 0 1 -823
box 0 0 96 799
use nand2 g12025
timestamp 1386234792
transform 1 0 21168 0 1 -823
box 0 0 96 799
use nand2 g12027
timestamp 1386234792
transform 1 0 21264 0 1 -823
box 0 0 96 799
use nand2 g12028
timestamp 1386234792
transform 1 0 21360 0 1 -823
box 0 0 96 799
use nand2 g12030
timestamp 1386234792
transform 1 0 21456 0 1 -823
box 0 0 96 799
use nand4 g11966
timestamp 1386234936
transform 1 0 21552 0 1 -823
box 0 0 144 799
use nand3 g12032
timestamp 1386234893
transform 1 0 21696 0 1 -823
box 0 0 120 799
use and2 g12038
timestamp 1386234845
transform 1 0 21816 0 1 -823
box 0 0 120 799
use and2 g12040
timestamp 1386234845
transform 1 0 21936 0 1 -823
box 0 0 120 799
use inv g12044
timestamp 1386238110
transform 1 0 22056 0 1 -823
box 0 0 120 799
use nand4 g11936
timestamp 1386234936
transform 1 0 22176 0 1 -823
box 0 0 144 799
use nand2 g11989
timestamp 1386234792
transform 1 0 22320 0 1 -823
box 0 0 96 799
use nand4 g11998
timestamp 1386234936
transform 1 0 22416 0 1 -823
box 0 0 144 799
use inv g12008
timestamp 1386238110
transform 1 0 22560 0 1 -823
box 0 0 120 799
use nand2 g12010
timestamp 1386234792
transform 1 0 22680 0 1 -823
box 0 0 96 799
use nand4 g11950
timestamp 1386234936
transform 1 0 22776 0 1 -823
box 0 0 144 799
use nand2 g12013
timestamp 1386234792
transform 1 0 22920 0 1 -823
box 0 0 96 799
use nand2 g12019
timestamp 1386234792
transform 1 0 23016 0 1 -823
box 0 0 96 799
use nand4 g11965
timestamp 1386234936
transform 1 0 23112 0 1 -823
box 0 0 144 799
use nand4 g11959
timestamp 1386234936
transform 1 0 23256 0 1 -823
box 0 0 144 799
use inv g12100
timestamp 1386238110
transform 1 0 23400 0 1 -823
box 0 0 120 799
use nand3 g12033
timestamp 1386234893
transform 1 0 23520 0 1 -823
box 0 0 120 799
use nand3 g12037
timestamp 1386234893
transform 1 0 23640 0 1 -823
box 0 0 120 799
use nand3 g12042
timestamp 1386234893
transform 1 0 23760 0 1 -823
box 0 0 120 799
use nand3 g12045
timestamp 1386234893
transform 1 0 23880 0 1 -823
box 0 0 120 799
use nand3 g12046
timestamp 1386234893
transform 1 0 24000 0 1 -823
box 0 0 120 799
use nand3 g12047
timestamp 1386234893
transform 1 0 24120 0 1 -823
box 0 0 120 799
use nand3 g12048
timestamp 1386234893
transform 1 0 24240 0 1 -823
box 0 0 120 799
use nand3 g12049
timestamp 1386234893
transform 1 0 24360 0 1 -823
box 0 0 120 799
use nand4 g11934
timestamp 1386234936
transform 1 0 24480 0 1 -823
box 0 0 144 799
use inv g12062
timestamp 1386238110
transform 1 0 24624 0 1 -823
box 0 0 120 799
use nand2 g12068
timestamp 1386234792
transform 1 0 24744 0 1 -823
box 0 0 96 799
use and2 g12069
timestamp 1386234845
transform 1 0 24840 0 1 -823
box 0 0 120 799
use nand2 g12070
timestamp 1386234792
transform 1 0 24960 0 1 -823
box 0 0 96 799
use nand2 g12073
timestamp 1386234792
transform 1 0 25056 0 1 -823
box 0 0 96 799
use nand2 g12080
timestamp 1386234792
transform 1 0 25152 0 1 -823
box 0 0 96 799
use and2 g12085
timestamp 1386234845
transform 1 0 25248 0 1 -823
box 0 0 120 799
use nand2 g12087
timestamp 1386234792
transform 1 0 25368 0 1 -823
box 0 0 96 799
use nand2 g12088
timestamp 1386234792
transform 1 0 25464 0 1 -823
box 0 0 96 799
use scandtype stateSub_reg_1
timestamp 1386241841
transform 1 0 25560 0 1 -823
box 0 0 624 799
use nand2 g12090
timestamp 1386234792
transform 1 0 26184 0 1 -823
box 0 0 96 799
use nand2 g12001
timestamp 1386234792
transform 1 0 26280 0 1 -823
box 0 0 96 799
use nand4 g12009
timestamp 1386234936
transform 1 0 26376 0 1 -823
box 0 0 144 799
use nand2 g12091
timestamp 1386234792
transform 1 0 26520 0 1 -823
box 0 0 96 799
use and2 g12012
timestamp 1386234845
transform 1 0 26616 0 1 -823
box 0 0 120 799
use nand3 g12021
timestamp 1386234893
transform 1 0 26736 0 1 -823
box 0 0 120 799
use and2 g11956
timestamp 1386234845
transform 1 0 26856 0 1 -823
box 0 0 120 799
use nand3 g12024
timestamp 1386234893
transform 1 0 26976 0 1 -823
box 0 0 120 799
use nand3 g12029
timestamp 1386234893
transform 1 0 27096 0 1 -823
box 0 0 120 799
use nand2 g12031
timestamp 1386234792
transform 1 0 27216 0 1 -823
box 0 0 96 799
use nand3 g12099
timestamp 1386234893
transform 1 0 27312 0 1 -823
box 0 0 120 799
use nand2 g12041
timestamp 1386234792
transform 1 0 27432 0 1 -823
box 0 0 96 799
use nand4 g11975
timestamp 1386234936
transform 1 0 27528 0 1 -823
box 0 0 144 799
use nand2 g12098
timestamp 1386234792
transform 1 0 27672 0 1 -823
box 0 0 96 799
use nand2 g12063
timestamp 1386234792
transform 1 0 27768 0 1 -823
box 0 0 96 799
use nand2 g12065
timestamp 1386234792
transform 1 0 27864 0 1 -823
box 0 0 96 799
use nand2 g12066
timestamp 1386234792
transform 1 0 27960 0 1 -823
box 0 0 96 799
use nand2 g12067
timestamp 1386234792
transform 1 0 28056 0 1 -823
box 0 0 96 799
use and2 g12097
timestamp 1386234845
transform 1 0 28152 0 1 -823
box 0 0 120 799
use nand2 g12074
timestamp 1386234792
transform 1 0 28272 0 1 -823
box 0 0 96 799
use nand2 g12075
timestamp 1386234792
transform 1 0 28368 0 1 -823
box 0 0 96 799
use nand2 g12076
timestamp 1386234792
transform 1 0 28464 0 1 -823
box 0 0 96 799
use nand2 g12077
timestamp 1386234792
transform 1 0 28560 0 1 -823
box 0 0 96 799
use nand2 g12078
timestamp 1386234792
transform 1 0 28656 0 1 -823
box 0 0 96 799
use nand2 g12081
timestamp 1386234792
transform 1 0 28752 0 1 -823
box 0 0 96 799
use nand2 g12082
timestamp 1386234792
transform 1 0 28848 0 1 -823
box 0 0 96 799
use nand2 g12084
timestamp 1386234792
transform 1 0 28944 0 1 -823
box 0 0 96 799
use nand2 g12086
timestamp 1386234792
transform 1 0 29040 0 1 -823
box 0 0 96 799
use nand3 g12101
timestamp 1386234893
transform 1 0 29136 0 1 -823
box 0 0 120 799
use nand2 g12089
timestamp 1386234792
transform 1 0 29256 0 1 -823
box 0 0 96 799
use scandtype IntReq_reg
timestamp 1386241841
transform 1 0 29352 0 1 -823
box 0 0 624 799
use and2 g12092
timestamp 1386234845
transform 1 0 29976 0 1 -823
box 0 0 120 799
use nand2 g12096
timestamp 1386234792
transform 1 0 30096 0 1 -823
box 0 0 96 799
use nand3 g12053
timestamp 1386234893
transform 1 0 30192 0 1 -823
box 0 0 120 799
use inv g12054
timestamp 1386238110
transform 1 0 30312 0 1 -823
box 0 0 120 799
use nor2 g12056
timestamp 1386235306
transform 1 0 30432 0 1 -823
box 0 0 120 799
use nor2 g12058
timestamp 1386235306
transform 1 0 30552 0 1 -823
box 0 0 120 799
use nand3 g12003
timestamp 1386234893
transform 1 0 30672 0 1 -823
box 0 0 120 799
use nand3 g12105
timestamp 1386234893
transform 1 0 30792 0 1 -823
box 0 0 120 799
use and2 g12120
timestamp 1386234845
transform 1 0 30912 0 1 -823
box 0 0 120 799
use and2 g12121
timestamp 1386234845
transform 1 0 31032 0 1 -823
box 0 0 120 799
use nand3 g12011
timestamp 1386234893
transform 1 0 31152 0 1 -823
box 0 0 120 799
use and2 g12130
timestamp 1386234845
transform 1 0 31272 0 1 -823
box 0 0 120 799
use nand3 g12016
timestamp 1386234893
transform 1 0 31392 0 1 -823
box 0 0 120 799
use nand2 g12139
timestamp 1386234792
transform 1 0 31512 0 1 -823
box 0 0 96 799
use nand3 g12023
timestamp 1386234893
transform 1 0 31608 0 1 -823
box 0 0 120 799
use nand2 g12026
timestamp 1386234792
transform 1 0 31728 0 1 -823
box 0 0 96 799
use nand2 g12034
timestamp 1386234792
transform 1 0 31824 0 1 -823
box 0 0 96 799
use nand3 g12039
timestamp 1386234893
transform 1 0 31920 0 1 -823
box 0 0 120 799
use nand2 g12094
timestamp 1386234792
transform 1 0 32040 0 1 -823
box 0 0 96 799
use inv g12051
timestamp 1386238110
transform 1 0 32136 0 1 -823
box 0 0 120 799
use nand4 g12055
timestamp 1386234936
transform 1 0 32256 0 1 -823
box 0 0 144 799
use nor2 g12057
timestamp 1386235306
transform 1 0 32400 0 1 -823
box 0 0 120 799
use nand2 g12060
timestamp 1386234792
transform 1 0 32520 0 1 -823
box 0 0 96 799
use nand2 g12061
timestamp 1386234792
transform 1 0 32616 0 1 -823
box 0 0 96 799
use nand2 g12064
timestamp 1386234792
transform 1 0 32712 0 1 -823
box 0 0 96 799
use nand3 g12083
timestamp 1386234893
transform 1 0 32808 0 1 -823
box 0 0 120 799
use nand3 g12102
timestamp 1386234893
transform 1 0 32928 0 1 -823
box 0 0 120 799
use inv g12103
timestamp 1386238110
transform 1 0 33048 0 1 -823
box 0 0 120 799
use nand3 g12106
timestamp 1386234893
transform 1 0 33168 0 1 -823
box 0 0 120 799
use and2 g12117
timestamp 1386234845
transform 1 0 33288 0 1 -823
box 0 0 120 799
use nand2 g12118
timestamp 1386234792
transform 1 0 33408 0 1 -823
box 0 0 96 799
use nand2 g12123
timestamp 1386234792
transform 1 0 33504 0 1 -823
box 0 0 96 799
use inv g12124
timestamp 1386238110
transform 1 0 33600 0 1 -823
box 0 0 120 799
use nand2 g12128
timestamp 1386234792
transform 1 0 33720 0 1 -823
box 0 0 96 799
use and2 g12129
timestamp 1386234845
transform 1 0 33816 0 1 -823
box 0 0 120 799
use nand2 g12132
timestamp 1386234792
transform 1 0 33936 0 1 -823
box 0 0 96 799
use nand2 g12135
timestamp 1386234792
transform 1 0 34032 0 1 -823
box 0 0 96 799
use nand2 g12136
timestamp 1386234792
transform 1 0 34128 0 1 -823
box 0 0 96 799
use and2 g12138
timestamp 1386234845
transform 1 0 34224 0 1 -823
box 0 0 120 799
use nand2 g12143
timestamp 1386234792
transform 1 0 34344 0 1 -823
box 0 0 96 799
use nand2 g12147
timestamp 1386234792
transform 1 0 34440 0 1 -823
box 0 0 96 799
use inv g12179
timestamp 1386238110
transform 1 0 34536 0 1 -823
box 0 0 120 799
use nand4 g12052
timestamp 1386234936
transform 1 0 34656 0 1 -823
box 0 0 144 799
use nand2 g12059
timestamp 1386234792
transform 1 0 34800 0 1 -823
box 0 0 96 799
use nand2 g12071
timestamp 1386234792
transform 1 0 34896 0 1 -823
box 0 0 96 799
use nand2 g12072
timestamp 1386234792
transform 1 0 34992 0 1 -823
box 0 0 96 799
use and2 g12079
timestamp 1386234845
transform 1 0 35088 0 1 -823
box 0 0 120 799
use and2 g12095
timestamp 1386234845
transform 1 0 35208 0 1 -823
box 0 0 120 799
use nand3 g12104
timestamp 1386234893
transform 1 0 35328 0 1 -823
box 0 0 120 799
use nor2 g12107
timestamp 1386235306
transform 1 0 35448 0 1 -823
box 0 0 120 799
use nand2 g12113
timestamp 1386234792
transform 1 0 35568 0 1 -823
box 0 0 96 799
use nand2 g12115
timestamp 1386234792
transform 1 0 35664 0 1 -823
box 0 0 96 799
use nand2 g12119
timestamp 1386234792
transform 1 0 35760 0 1 -823
box 0 0 96 799
use nand2 g12125
timestamp 1386234792
transform 1 0 35856 0 1 -823
box 0 0 96 799
use nand2 g12126
timestamp 1386234792
transform 1 0 35952 0 1 -823
box 0 0 96 799
use inv g12174
timestamp 1386238110
transform 1 0 36048 0 1 -823
box 0 0 120 799
use nand2 g12180
timestamp 1386234792
transform 1 0 36168 0 1 -823
box 0 0 96 799
use nand2 g12182
timestamp 1386234792
transform 1 0 36264 0 1 -823
box 0 0 96 799
use nand2 g12183
timestamp 1386234792
transform 1 0 36360 0 1 -823
box 0 0 96 799
use inv g12184
timestamp 1386238110
transform 1 0 36456 0 1 -823
box 0 0 120 799
use inv g12187
timestamp 1386238110
transform 1 0 36576 0 1 -823
box 0 0 120 799
use nand2 g12192
timestamp 1386234792
transform 1 0 36696 0 1 -823
box 0 0 96 799
use nand2 g12194
timestamp 1386234792
transform 1 0 36792 0 1 -823
box 0 0 96 799
use nand4 g12050
timestamp 1386234936
transform 1 0 36888 0 1 -823
box 0 0 144 799
use nand2 g12093
timestamp 1386234792
transform 1 0 37032 0 1 -823
box 0 0 96 799
use nand2 g12108
timestamp 1386234792
transform 1 0 37128 0 1 -823
box 0 0 96 799
use nor2 g12110
timestamp 1386235306
transform 1 0 37224 0 1 -823
box 0 0 120 799
use nor2 g12111
timestamp 1386235306
transform 1 0 37344 0 1 -823
box 0 0 120 799
use nor2 g12112
timestamp 1386235306
transform 1 0 37464 0 1 -823
box 0 0 120 799
use nand2 g12114
timestamp 1386234792
transform 1 0 37584 0 1 -823
box 0 0 96 799
use nand2 g12134
timestamp 1386234792
transform 1 0 37680 0 1 -823
box 0 0 96 799
use nand2 g12141
timestamp 1386234792
transform 1 0 37776 0 1 -823
box 0 0 96 799
use nand2 g12144
timestamp 1386234792
transform 1 0 37872 0 1 -823
box 0 0 96 799
use nand3 g12146
timestamp 1386234893
transform 1 0 37968 0 1 -823
box 0 0 120 799
use inv g12148
timestamp 1386238110
transform 1 0 38088 0 1 -823
box 0 0 120 799
use nand2 g12161
timestamp 1386234792
transform 1 0 38208 0 1 -823
box 0 0 96 799
use and2 g12162
timestamp 1386234845
transform 1 0 38304 0 1 -823
box 0 0 120 799
use inv g12163
timestamp 1386238110
transform 1 0 38424 0 1 -823
box 0 0 120 799
use and2 g12165
timestamp 1386234845
transform 1 0 38544 0 1 -823
box 0 0 120 799
use nand2 g12173
timestamp 1386234792
transform 1 0 38664 0 1 -823
box 0 0 96 799
use nand2 g12175
timestamp 1386234792
transform 1 0 38760 0 1 -823
box 0 0 96 799
use nand2 g12181
timestamp 1386234792
transform 1 0 38856 0 1 -823
box 0 0 96 799
use nand2 g12185
timestamp 1386234792
transform 1 0 38952 0 1 -823
box 0 0 96 799
use nor2 g12188
timestamp 1386235306
transform 1 0 39048 0 1 -823
box 0 0 120 799
use nand2 g12191
timestamp 1386234792
transform 1 0 39168 0 1 -823
box 0 0 96 799
use nand2 g12199
timestamp 1386234792
transform 1 0 39264 0 1 -823
box 0 0 96 799
use nand2 g12201
timestamp 1386234792
transform 1 0 39360 0 1 -823
box 0 0 96 799
use nand2 g12202
timestamp 1386234792
transform 1 0 39456 0 1 -823
box 0 0 96 799
use nand2 g12203
timestamp 1386234792
transform 1 0 39552 0 1 -823
box 0 0 96 799
use nor2 g12109
timestamp 1386235306
transform 1 0 39648 0 1 -823
box 0 0 120 799
use nand2 g12116
timestamp 1386234792
transform 1 0 39768 0 1 -823
box 0 0 96 799
use nand2 g12122
timestamp 1386234792
transform 1 0 39864 0 1 -823
box 0 0 96 799
use nand2 g12131
timestamp 1386234792
transform 1 0 39960 0 1 -823
box 0 0 96 799
use nand2 g12137
timestamp 1386234792
transform 1 0 40056 0 1 -823
box 0 0 96 799
use nand2 g12140
timestamp 1386234792
transform 1 0 40152 0 1 -823
box 0 0 96 799
use nand2 g12142
timestamp 1386234792
transform 1 0 40248 0 1 -823
box 0 0 96 799
use nand2 g12145
timestamp 1386234792
transform 1 0 40344 0 1 -823
box 0 0 96 799
use nand3 g12149
timestamp 1386234893
transform 1 0 40440 0 1 -823
box 0 0 120 799
use nand2 g12153
timestamp 1386234792
transform 1 0 40560 0 1 -823
box 0 0 96 799
use nor2 g12155
timestamp 1386235306
transform 1 0 40656 0 1 -823
box 0 0 120 799
use nand2 g12160
timestamp 1386234792
transform 1 0 40776 0 1 -823
box 0 0 96 799
use nor2 g12164
timestamp 1386235306
transform 1 0 40872 0 1 -823
box 0 0 120 799
use nand2 g12166
timestamp 1386234792
transform 1 0 40992 0 1 -823
box 0 0 96 799
use inv g12167
timestamp 1386238110
transform 1 0 41088 0 1 -823
box 0 0 120 799
use nand2 g12169
timestamp 1386234792
transform 1 0 41208 0 1 -823
box 0 0 96 799
use nand2 g12178
timestamp 1386234792
transform 1 0 41304 0 1 -823
box 0 0 96 799
use inv g12254
timestamp 1386238110
transform 1 0 41400 0 1 -823
box 0 0 120 799
use nand2 g12190
timestamp 1386234792
transform 1 0 41520 0 1 -823
box 0 0 96 799
use nand2 g12195
timestamp 1386234792
transform 1 0 41616 0 1 -823
box 0 0 96 799
use nand2 g12196
timestamp 1386234792
transform 1 0 41712 0 1 -823
box 0 0 96 799
use nand2 g12197
timestamp 1386234792
transform 1 0 41808 0 1 -823
box 0 0 96 799
use nand2 g12200
timestamp 1386234792
transform 1 0 41904 0 1 -823
box 0 0 96 799
use nor2 g12206
timestamp 1386235306
transform 1 0 42000 0 1 -823
box 0 0 120 799
use inv g12222
timestamp 1386238110
transform 1 0 42120 0 1 -823
box 0 0 120 799
use inv g12227
timestamp 1386238110
transform 1 0 42240 0 1 -823
box 0 0 120 799
use inv g12243
timestamp 1386238110
transform 1 0 42360 0 1 -823
box 0 0 120 799
use nand3 g12256
timestamp 1386234893
transform 1 0 42480 0 1 -823
box 0 0 120 799
use inv g12258
timestamp 1386238110
transform 1 0 42600 0 1 -823
box 0 0 120 799
use inv g12261
timestamp 1386238110
transform 1 0 42720 0 1 -823
box 0 0 120 799
use nand2 g12189
timestamp 1386234792
transform 1 0 42840 0 1 -823
box 0 0 96 799
use and2 g12186
timestamp 1386234845
transform 1 0 42936 0 1 -823
box 0 0 120 799
use inv g12170
timestamp 1386238110
transform 1 0 43056 0 1 -823
box 0 0 120 799
use nand2 g12168
timestamp 1386234792
transform 1 0 43176 0 1 -823
box 0 0 96 799
use nand2 g12133
timestamp 1386234792
transform 1 0 43272 0 1 -823
box 0 0 96 799
use nand2 g12150
timestamp 1386234792
transform 1 0 43368 0 1 -823
box 0 0 96 799
use nand2 g12151
timestamp 1386234792
transform 1 0 43464 0 1 -823
box 0 0 96 799
use nand2 g12154
timestamp 1386234792
transform 1 0 43560 0 1 -823
box 0 0 96 799
use inv g12176
timestamp 1386238110
transform 1 0 43656 0 1 -823
box 0 0 120 799
use nand2 g12177
timestamp 1386234792
transform 1 0 43776 0 1 -823
box 0 0 96 799
use nand2 g12193
timestamp 1386234792
transform 1 0 43872 0 1 -823
box 0 0 96 799
use nand2 g12204
timestamp 1386234792
transform 1 0 43968 0 1 -823
box 0 0 96 799
use nand3 g12205
timestamp 1386234893
transform 1 0 44064 0 1 -823
box 0 0 120 799
use mux2 g12207
timestamp 1386235218
transform 1 0 44184 0 1 -823
box 0 0 192 799
use nand2 g12213
timestamp 1386234792
transform 1 0 44376 0 1 -823
box 0 0 96 799
use inv g12215
timestamp 1386238110
transform 1 0 44472 0 1 -823
box 0 0 120 799
use nor2 g12218
timestamp 1386235306
transform 1 0 44592 0 1 -823
box 0 0 120 799
use nand2 g12221
timestamp 1386234792
transform 1 0 44712 0 1 -823
box 0 0 96 799
use nand2 g12223
timestamp 1386234792
transform 1 0 44808 0 1 -823
box 0 0 96 799
use nand2 g12226
timestamp 1386234792
transform 1 0 44904 0 1 -823
box 0 0 96 799
use nor2 g12228
timestamp 1386235306
transform 1 0 45000 0 1 -823
box 0 0 120 799
use inv g12231
timestamp 1386238110
transform 1 0 45120 0 1 -823
box 0 0 120 799
use inv g12233
timestamp 1386238110
transform 1 0 45240 0 1 -823
box 0 0 120 799
use nand2 g12244
timestamp 1386234792
transform 1 0 45360 0 1 -823
box 0 0 96 799
use nand2 g12248
timestamp 1386234792
transform 1 0 45456 0 1 -823
box 0 0 96 799
use inv g12249
timestamp 1386238110
transform 1 0 45552 0 1 -823
box 0 0 120 799
use nand2 g12251
timestamp 1386234792
transform 1 0 45672 0 1 -823
box 0 0 96 799
use nand2 g12252
timestamp 1386234792
transform 1 0 45768 0 1 -823
box 0 0 96 799
use nand2 g12253
timestamp 1386234792
transform 1 0 45864 0 1 -823
box 0 0 96 799
use nand2 g12255
timestamp 1386234792
transform 1 0 45960 0 1 -823
box 0 0 96 799
use nand2 g12257
timestamp 1386234792
transform 1 0 46056 0 1 -823
box 0 0 96 799
use nand2 g12259
timestamp 1386234792
transform 1 0 46152 0 1 -823
box 0 0 96 799
use and2 g12263
timestamp 1386234845
transform 1 0 46248 0 1 -823
box 0 0 120 799
use nand2 g12269
timestamp 1386234792
transform 1 0 46368 0 1 -823
box 0 0 96 799
use nand2 g12217
timestamp 1386234792
transform 1 0 46464 0 1 -823
box 0 0 96 799
use and2 g12237
timestamp 1386234845
transform 1 0 46560 0 1 -823
box 0 0 120 799
use nand4 g12127
timestamp 1386234936
transform 1 0 46680 0 1 -823
box 0 0 144 799
use nand3 g12152
timestamp 1386234893
transform 1 0 46824 0 1 -823
box 0 0 120 799
use and2 g12156
timestamp 1386234845
transform 1 0 46944 0 1 -823
box 0 0 120 799
use nand2 g12157
timestamp 1386234792
transform 1 0 47064 0 1 -823
box 0 0 96 799
use nand2 g12158
timestamp 1386234792
transform 1 0 47160 0 1 -823
box 0 0 96 799
use nand3 g12159
timestamp 1386234893
transform 1 0 47256 0 1 -823
box 0 0 120 799
use nand2 g12262
timestamp 1386234792
transform 1 0 47376 0 1 -823
box 0 0 96 799
use nand3 g12171
timestamp 1386234893
transform 1 0 47472 0 1 -823
box 0 0 120 799
use nand3 g12172
timestamp 1386234893
transform 1 0 47592 0 1 -823
box 0 0 120 799
use and2 g12266
timestamp 1386234845
transform 1 0 47712 0 1 -823
box 0 0 120 799
use mux2 g12208
timestamp 1386235218
transform 1 0 47832 0 1 -823
box 0 0 192 799
use inv g12270
timestamp 1386238110
transform 1 0 48024 0 1 -823
box 0 0 120 799
use nor2 g12214
timestamp 1386235306
transform 1 0 48144 0 1 -823
box 0 0 120 799
use nor2 g12216
timestamp 1386235306
transform 1 0 48264 0 1 -823
box 0 0 120 799
use nand2 g12220
timestamp 1386234792
transform 1 0 48384 0 1 -823
box 0 0 96 799
use nand2 g12224
timestamp 1386234792
transform 1 0 48480 0 1 -823
box 0 0 96 799
use nand2 g12225
timestamp 1386234792
transform 1 0 48576 0 1 -823
box 0 0 96 799
use nand2 g12229
timestamp 1386234792
transform 1 0 48672 0 1 -823
box 0 0 96 799
use nand2 g12230
timestamp 1386234792
transform 1 0 48768 0 1 -823
box 0 0 96 799
use nand2 g12232
timestamp 1386234792
transform 1 0 48864 0 1 -823
box 0 0 96 799
use nand2 g12234
timestamp 1386234792
transform 1 0 48960 0 1 -823
box 0 0 96 799
use nand2 g12236
timestamp 1386234792
transform 1 0 49056 0 1 -823
box 0 0 96 799
use nand2 g12239
timestamp 1386234792
transform 1 0 49152 0 1 -823
box 0 0 96 799
use nand2 g12240
timestamp 1386234792
transform 1 0 49248 0 1 -823
box 0 0 96 799
use nand2 g12277
timestamp 1386234792
transform 1 0 49344 0 1 -823
box 0 0 96 799
use nand2 g12245
timestamp 1386234792
transform 1 0 49440 0 1 -823
box 0 0 96 799
use nand2 g12246
timestamp 1386234792
transform 1 0 49536 0 1 -823
box 0 0 96 799
use nand2 g12247
timestamp 1386234792
transform 1 0 49632 0 1 -823
box 0 0 96 799
use nor2 g12250
timestamp 1386235306
transform 1 0 49728 0 1 -823
box 0 0 120 799
use and2 g12265
timestamp 1386234845
transform 1 0 49848 0 1 -823
box 0 0 120 799
use nand2 g12268
timestamp 1386234792
transform 1 0 49968 0 1 -823
box 0 0 96 799
use nand2 g12276
timestamp 1386234792
transform 1 0 50064 0 1 -823
box 0 0 96 799
use nand2 g12238
timestamp 1386234792
transform 1 0 50160 0 1 -823
box 0 0 96 799
use nand2 g12212
timestamp 1386234792
transform 1 0 50256 0 1 -823
box 0 0 96 799
use scandtype IRQ2_reg
timestamp 1386241841
transform 1 0 50352 0 1 -823
box 0 0 624 799
use nand2 g12275
timestamp 1386234792
transform 1 0 50976 0 1 -823
box 0 0 96 799
use nand2 g12260
timestamp 1386234792
transform 1 0 51072 0 1 -823
box 0 0 96 799
use nand2 g12209
timestamp 1386234792
transform 1 0 51168 0 1 -823
box 0 0 96 799
use nand3 g12242
timestamp 1386234893
transform 1 0 51264 0 1 -823
box 0 0 120 799
use and2 g12219
timestamp 1386234845
transform 1 0 51384 0 1 -823
box 0 0 120 799
use inv g12284
timestamp 1386238110
transform 1 0 51504 0 1 -823
box 0 0 120 799
use nand2 g12241
timestamp 1386234792
transform 1 0 51624 0 1 -823
box 0 0 96 799
use nand4 g12198
timestamp 1386234936
transform 1 0 51720 0 1 -823
box 0 0 144 799
use and2 g12264
timestamp 1386234845
transform 1 0 51864 0 1 -823
box 0 0 120 799
use nand3 g12274
timestamp 1386234893
transform 1 0 51984 0 1 -823
box 0 0 120 799
use inv g12288
timestamp 1386238110
transform 1 0 52104 0 1 -823
box 0 0 120 799
use inv g12290
timestamp 1386238110
transform 1 0 52224 0 1 -823
box 0 0 120 799
use inv g12293
timestamp 1386238110
transform 1 0 52344 0 1 -823
box 0 0 120 799
use inv g12307
timestamp 1386238110
transform 1 0 52464 0 1 -823
box 0 0 120 799
use nand2 g12235
timestamp 1386234792
transform 1 0 52584 0 1 -823
box 0 0 96 799
use nor2 g12271
timestamp 1386235306
transform 1 0 52680 0 1 -823
box 0 0 120 799
use inv g12324
timestamp 1386238110
transform 1 0 52800 0 1 -823
box 0 0 120 799
use inv g12304
timestamp 1386238110
transform 1 0 52920 0 1 -823
box 0 0 120 799
use nand2 g12267
timestamp 1386234792
transform 1 0 53040 0 1 -823
box 0 0 96 799
use inv g12299
timestamp 1386238110
transform 1 0 53136 0 1 -823
box 0 0 120 799
use nand3 g12273
timestamp 1386234893
transform 1 0 53256 0 1 -823
box 0 0 120 799
use inv g12286
timestamp 1386238110
transform 1 0 53376 0 1 -823
box 0 0 120 799
use nand2 g12325
timestamp 1386234792
transform 1 0 53496 0 1 -823
box 0 0 96 799
use nand2 g12281
timestamp 1386234792
transform 1 0 53592 0 1 -823
box 0 0 96 799
use inv g12317
timestamp 1386238110
transform 1 0 53688 0 1 -823
box 0 0 120 799
use nand2 g12289
timestamp 1386234792
transform 1 0 53808 0 1 -823
box 0 0 96 799
use inv g12315
timestamp 1386238110
transform 1 0 53904 0 1 -823
box 0 0 120 799
use nand2 g12285
timestamp 1386234792
transform 1 0 54024 0 1 -823
box 0 0 96 799
use nand2 g12295
timestamp 1386234792
transform 1 0 54120 0 1 -823
box 0 0 96 799
use nand2 g12280
timestamp 1386234792
transform 1 0 54216 0 1 -823
box 0 0 96 799
use inv g12282
timestamp 1386238110
transform 1 0 54312 0 1 -823
box 0 0 120 799
use nor2 g12287
timestamp 1386235306
transform 1 0 54432 0 1 -823
box 0 0 120 799
use nor2 g12297
timestamp 1386235306
transform 1 0 54552 0 1 -823
box 0 0 120 799
use and2 g12302
timestamp 1386234845
transform 1 0 54672 0 1 -823
box 0 0 120 799
use nand2 g12308
timestamp 1386234792
transform 1 0 54792 0 1 -823
box 0 0 96 799
use nand2 g12309
timestamp 1386234792
transform 1 0 54888 0 1 -823
box 0 0 96 799
use nand2 g12312
timestamp 1386234792
transform 1 0 54984 0 1 -823
box 0 0 96 799
use inv g12322
timestamp 1386238110
transform 1 0 55080 0 1 -823
box 0 0 120 799
use nand2 g12310
timestamp 1386234792
transform 1 0 55200 0 1 -823
box 0 0 96 799
use nor2 g12330
timestamp 1386235306
transform 1 0 55296 0 1 -823
box 0 0 120 799
use nor2 g12329
timestamp 1386235306
transform 1 0 55416 0 1 -823
box 0 0 120 799
use inv g12327
timestamp 1386238110
transform 1 0 55536 0 1 -823
box 0 0 120 799
use nand2 g12300
timestamp 1386234792
transform 1 0 55656 0 1 -823
box 0 0 96 799
use nand2 g12305
timestamp 1386234792
transform 1 0 55752 0 1 -823
box 0 0 96 799
use nand2 g12303
timestamp 1386234792
transform 1 0 55848 0 1 -823
box 0 0 96 799
use scandtype IRQ1_reg
timestamp 1386241841
transform 1 0 55944 0 1 -823
box 0 0 624 799
use nand3 g12272
timestamp 1386234893
transform 1 0 56568 0 1 -823
box 0 0 120 799
use nand2 g12296
timestamp 1386234792
transform 1 0 56688 0 1 -823
box 0 0 96 799
use nand2 g12294
timestamp 1386234792
transform 1 0 56784 0 1 -823
box 0 0 96 799
use inv g12320
timestamp 1386238110
transform 1 0 56880 0 1 -823
box 0 0 120 799
use nand2 g12306
timestamp 1386234792
transform 1 0 57000 0 1 -823
box 0 0 96 799
use nand2 g12291
timestamp 1386234792
transform 1 0 57096 0 1 -823
box 0 0 96 799
use nand2 g12313
timestamp 1386234792
transform 1 0 57192 0 1 -823
box 0 0 96 799
use nand2 g12319
timestamp 1386234792
transform 1 0 57288 0 1 -823
box 0 0 96 799
use nand2 g12328
timestamp 1386234792
transform 1 0 57384 0 1 -823
box 0 0 96 799
use nor2 g12298
timestamp 1386235306
transform 1 0 57480 0 1 -823
box 0 0 120 799
use nand2 g12316
timestamp 1386234792
transform 1 0 57600 0 1 -823
box 0 0 96 799
use nor2 g12279
timestamp 1386235306
transform 1 0 57696 0 1 -823
box 0 0 120 799
use and2 g12301
timestamp 1386234845
transform 1 0 57816 0 1 -823
box 0 0 120 799
use nand2 g12314
timestamp 1386234792
transform 1 0 57936 0 1 -823
box 0 0 96 799
use nand2 g12323
timestamp 1386234792
transform 1 0 58032 0 1 -823
box 0 0 96 799
use nand2 g12321
timestamp 1386234792
transform 1 0 58128 0 1 -823
box 0 0 96 799
use nand2 g12326
timestamp 1386234792
transform 1 0 58224 0 1 -823
box 0 0 96 799
use nor2 g12283
timestamp 1386235306
transform 1 0 58320 0 1 -823
box 0 0 120 799
use nor2 g12292
timestamp 1386235306
transform 1 0 58440 0 1 -823
box 0 0 120 799
use nand2 g12318
timestamp 1386234792
transform 1 0 58560 0 1 -823
box 0 0 96 799
use and2 g12311
timestamp 1386234845
transform 1 0 58656 0 1 -823
box 0 0 120 799
use inv g12335
timestamp 1386238110
transform 1 0 58776 0 1 -823
box 0 0 120 799
use inv g12346
timestamp 1386238110
transform 1 0 58896 0 1 -823
box 0 0 120 799
use inv g12347
timestamp 1386238110
transform 1 0 59016 0 1 -823
box 0 0 120 799
use inv g12337
timestamp 1386238110
transform 1 0 59136 0 1 -823
box 0 0 120 799
use inv g12345
timestamp 1386238110
transform 1 0 59256 0 1 -823
box 0 0 120 799
use inv g12340
timestamp 1386238110
transform 1 0 59376 0 1 -823
box 0 0 120 799
use inv g12339
timestamp 1386238110
transform 1 0 59496 0 1 -823
box 0 0 120 799
use inv g12334
timestamp 1386238110
transform 1 0 59616 0 1 -823
box 0 0 120 799
use inv g12341
timestamp 1386238110
transform 1 0 59736 0 1 -823
box 0 0 120 799
use inv g12342
timestamp 1386238110
transform 1 0 59856 0 1 -823
box 0 0 120 799
<< labels >>
rlabel metal1 32221 17972 32221 17982 3 Op1Sel
rlabel metal1 32221 9092 32221 9102 3 AluEn
rlabel metal1 32221 29252 32221 29262 3 LrEn
rlabel metal1 32221 29996 32221 30006 3 LrWe
rlabel metal1 32221 28292 32221 28302 3 PcWe
rlabel metal1 32221 27548 32221 27558 3 PcEn
rlabel metal1 32221 31556 32221 31566 3 IrWe
rlabel metal1 32221 27380 32221 27390 3 WdSel
rlabel metal1 32221 30764 32221 30774 3 ImmSel
rlabel metal1 32221 31748 32221 31758 3 MemEn
rlabel metal1 32221 16104 32221 16114 3 nWE
rlabel metal1 32221 16344 32221 16354 3 nOE
rlabel metal1 32221 16584 32221 16594 3 nME
rlabel metal1 32221 16824 32221 16834 3 ENB
rlabel metal1 32221 8664 32221 8674 3 ALE
rlabel metal1 32221 17304 32221 17314 3 CFlag
rlabel metal1 32221 9836 32221 9846 3 AluWe
rlabel metal1 32221 17540 32221 17550 3 Op2Sel[1]
rlabel metal1 32221 17780 32221 17790 3 Op2Sel[0]
rlabel metal1 66735 2072 66735 2082 5 OpcodeCondIn[7]
rlabel metal1 66735 2312 66735 2322 5 OpcodeCondIn[6]
rlabel metal1 66735 2552 66735 2562 5 OpcodeCondIn[5]
rlabel metal1 66735 2792 66735 2802 5 OpcodeCondIn[4]
rlabel metal1 66735 3032 66735 3042 5 OpcodeCondIn[3]
rlabel metal1 66735 3272 66735 3282 5 OpcodeCondIn[2]
rlabel metal1 66735 3512 66735 3522 5 OpcodeCondIn[1]
rlabel metal1 66735 3752 66735 3762 5 OpcodeCondIn[0]
rlabel metal1 66735 3992 66735 4002 5 Flags[3]
rlabel metal1 66735 4232 66735 4242 5 Flags[2]
rlabel metal1 66735 4472 66735 4482 5 Flags[1]
rlabel metal1 66735 4712 66735 4722 5 Flags[0]
rlabel metal1 66735 4952 66735 4962 5 nWait
rlabel metal1 66735 5192 66735 5202 5 nIRQ
rlabel metal1 66735 5432 66735 5442 5 AluOp[4]
rlabel metal1 66735 5672 66735 5682 5 AluOp[3]
rlabel metal1 66735 5912 66735 5922 5 AluOp[2]
rlabel metal1 66735 6152 66735 6162 5 AluOp[1]
rlabel metal1 66735 6392 66735 6402 5 AluOp[0]
rlabel metal1 66735 8792 66735 8802 5 RegWe
rlabel metal1 66735 23380 66735 23390 5 LrSel
rlabel metal1 66735 11672 66735 11682 5 Rs1Sel[1]
rlabel metal1 66735 11912 66735 11922 5 Rs1Sel[0]
rlabel metal1 66735 12152 66735 12162 5 RwSel[1]
rlabel metal1 66735 12392 66735 12402 5 RwSel[0]
rlabel metal1 66735 12632 66735 12642 5 AluOR[1]
rlabel metal1 66735 12872 66735 12882 5 AluOR[0]
rlabel metal1 66735 13112 66735 13122 5 PcSel[2]
rlabel metal1 66735 13352 66735 13362 5 PcSel[1]
rlabel metal1 66735 13592 66735 13602 5 PcSel[0]
rlabel metal1 66735 13832 66735 13842 5 SysBus[15]
rlabel metal1 66735 14072 66735 14082 5 SysBus[14]
rlabel metal1 66735 14312 66735 14322 5 SysBus[13]
rlabel metal1 66735 14552 66735 14562 5 SysBus[12]
rlabel metal1 66735 14792 66735 14802 5 SysBus[11]
rlabel metal1 66735 15032 66735 15042 5 SysBus[10]
rlabel metal1 66735 15272 66735 15282 5 SysBus[9]
rlabel metal1 66735 15512 66735 15522 5 SysBus[8]
rlabel metal1 66735 15752 66735 15762 5 SysBus[7]
rlabel metal1 66735 15992 66735 16002 5 SysBus[6]
rlabel metal1 66735 16232 66735 16242 5 SysBus[5]
rlabel metal1 66735 16472 66735 16482 5 SysBus[4]
rlabel metal1 66735 16712 66735 16722 5 SysBus[3]
rlabel metal1 66735 16952 66735 16962 5 SysBus[2]
rlabel metal1 66735 17192 66735 17202 5 SysBus[1]
rlabel metal1 66735 17432 66735 17442 5 SysBus[0]
<< end >>
