magic
tech c035u
timestamp 1394833348
<< checkpaint >>
rect 11921 22313 18638 22806
rect 5561 19679 18638 22313
rect 5561 18095 17377 19679
<< metal1 >>
rect 433 22062 13243 22072
rect 13257 22062 23764 22072
rect 456 22038 13436 22048
rect 13450 22038 23764 22048
rect 479 22014 13628 22024
rect 13642 22014 23764 22024
rect 502 21990 13820 22000
rect 13834 21990 23764 22000
rect 525 21966 14012 21976
rect 14026 21966 23764 21976
rect 548 21942 4340 21952
rect 4354 21942 23764 21952
rect 571 21918 4772 21928
rect 4786 21918 23764 21928
rect 594 21894 5204 21904
rect 5218 21894 23764 21904
rect 617 21870 4388 21880
rect 4402 21870 23764 21880
rect 640 21846 4820 21856
rect 4834 21846 23764 21856
rect 663 21822 5252 21832
rect 5266 21822 23764 21832
rect 686 21798 7340 21808
rect 7354 21798 23764 21808
rect 709 21774 7316 21784
rect 7330 21774 22772 21784
rect 22786 21774 23764 21784
rect 732 21750 7292 21760
rect 7306 21750 22964 21760
rect 22978 21750 23764 21760
rect 755 21726 23084 21736
rect 23098 21726 23764 21736
rect 778 21702 23204 21712
rect 23218 21702 23764 21712
rect 23997 18891 24189 18901
rect 3514 18780 3525 18790
rect -48 17893 419 17903
rect 433 17893 784 17903
rect -48 17861 784 17871
rect -48 17827 784 17837
rect 3477 17827 3525 17837
rect 23997 17827 24189 17837
rect 3477 17805 3525 17815
rect 23997 17715 24189 17725
rect 3514 17604 3525 17614
rect -48 16717 442 16727
rect 456 16717 784 16727
rect -48 16685 784 16695
rect -48 16651 784 16661
rect 3477 16651 3525 16661
rect 23997 16651 24189 16661
rect 3477 16629 3525 16639
rect 23997 16539 24189 16549
rect 3514 16428 3525 16438
rect -48 15541 465 15551
rect 479 15541 784 15551
rect -48 15509 784 15519
rect -48 15475 784 15485
rect 3477 15475 3525 15485
rect 23997 15475 24189 15485
rect 3477 15453 3525 15463
rect 23997 15363 24189 15373
rect 3514 15252 3525 15262
rect -48 14365 488 14375
rect 502 14365 784 14375
rect -48 14333 784 14343
rect -48 14299 784 14309
rect 3477 14299 3525 14309
rect 23997 14299 24189 14309
rect 3477 14277 3525 14287
rect 23997 14187 24189 14197
rect 3514 14076 3525 14086
rect -48 13189 511 13199
rect 525 13189 784 13199
rect -48 13157 784 13167
rect -48 13123 784 13133
rect 3477 13123 3525 13133
rect 23997 13123 24189 13133
rect 3477 13101 3525 13111
rect 23997 13011 24189 13021
rect 3514 12900 3525 12910
rect -48 12013 534 12023
rect 548 12013 784 12023
rect -48 11981 784 11991
rect -48 11947 784 11957
rect 3477 11947 3525 11957
rect 23997 11947 24189 11957
rect 3477 11925 3525 11935
rect 23997 11835 24189 11845
rect 3514 11724 3525 11734
rect -48 10837 557 10847
rect 571 10837 784 10847
rect -48 10805 784 10815
rect -48 10771 784 10781
rect 3477 10771 3525 10781
rect 23997 10771 24189 10781
rect 3477 10749 3525 10759
rect 23997 10659 24189 10669
rect 3514 10548 3525 10558
rect -48 9661 580 9671
rect 594 9661 784 9671
rect -48 9629 784 9639
rect -48 9595 784 9605
rect 3477 9595 3525 9605
rect 23997 9595 24189 9605
rect 3477 9573 3525 9583
rect 23997 9483 24189 9493
rect 3514 9372 3525 9382
rect -48 8485 603 8495
rect 617 8485 784 8495
rect -48 8453 784 8463
rect -48 8419 784 8429
rect 3477 8419 3525 8429
rect 23997 8419 24189 8429
rect 3477 8397 3525 8407
rect 23997 8307 24189 8317
rect 3514 8196 3525 8206
rect -48 7309 626 7319
rect 640 7309 784 7319
rect -48 7277 784 7287
rect -48 7243 784 7253
rect 3477 7243 3525 7253
rect 23997 7243 24189 7253
rect 3477 7221 3525 7231
rect 23997 7131 24189 7141
rect 3514 7020 3525 7030
rect -48 6133 649 6143
rect 663 6133 784 6143
rect -48 6101 784 6111
rect -48 6067 784 6077
rect 3477 6067 3525 6077
rect 23997 6067 24189 6077
rect 3477 6045 3525 6055
rect 23997 5955 24189 5965
rect 3514 5844 3525 5854
rect -48 4957 672 4967
rect 686 4957 784 4967
rect -48 4925 784 4935
rect -48 4891 784 4901
rect 3477 4891 3525 4901
rect 23997 4891 24189 4901
rect 3477 4869 3525 4879
rect 23997 4779 24189 4789
rect 3514 4668 3525 4678
rect -48 3781 695 3791
rect 709 3781 784 3791
rect -48 3749 784 3759
rect -48 3715 784 3725
rect 3477 3715 3525 3725
rect 23997 3715 24189 3725
rect 3477 3693 3525 3703
rect 23997 3603 24189 3613
rect 3514 3492 3525 3502
rect -48 2605 718 2615
rect 732 2605 784 2615
rect -48 2573 784 2583
rect -48 2539 784 2549
rect 3477 2539 3525 2549
rect 23997 2539 24189 2549
rect 3477 2517 3525 2527
rect 23997 2427 24189 2437
rect 3514 2316 3525 2326
rect -48 1429 741 1439
rect 755 1429 784 1439
rect -48 1397 784 1407
rect -48 1363 784 1373
rect 3477 1363 3525 1373
rect 23997 1363 24189 1373
rect 3477 1341 3525 1351
rect 23997 1251 24189 1261
rect 3514 1140 3525 1150
rect -48 253 764 263
rect 778 253 784 263
rect -48 221 784 231
rect -48 187 784 197
rect 3477 187 3525 197
rect 23997 187 24189 197
rect 3477 165 3525 175
rect 2474 72 17684 82
rect 17698 72 20348 82
rect 20362 72 20395 82
rect 20409 72 20444 82
rect 20458 72 20492 82
rect 20506 72 20540 82
rect 20554 72 20588 82
rect 20602 72 20636 82
rect 20650 72 20684 82
rect 20698 72 20996 82
rect 21010 72 21044 82
rect 21058 72 21091 82
rect 21105 72 21140 82
rect 21154 72 21452 82
rect 21466 72 21500 82
rect 21514 72 21884 82
rect 21898 72 25245 82
rect 989 51 3740 61
<< m2contact >>
rect 419 22060 433 22074
rect 13243 22061 13257 22075
rect 442 22036 456 22050
rect 13436 22036 13450 22050
rect 465 22012 479 22026
rect 13628 22012 13642 22026
rect 488 21988 502 22002
rect 13820 21988 13834 22002
rect 511 21964 525 21978
rect 14012 21964 14026 21979
rect 534 21940 548 21954
rect 4340 21940 4354 21954
rect 557 21916 571 21930
rect 4772 21916 4786 21930
rect 580 21892 594 21906
rect 5204 21892 5218 21906
rect 603 21868 617 21882
rect 4388 21868 4402 21882
rect 626 21844 640 21858
rect 4820 21844 4834 21858
rect 649 21820 663 21834
rect 5252 21820 5266 21834
rect 672 21796 686 21810
rect 7340 21796 7354 21810
rect 695 21772 709 21786
rect 7316 21772 7330 21786
rect 22772 21772 22786 21786
rect 718 21748 732 21762
rect 7292 21748 7306 21762
rect 22964 21747 22978 21761
rect 741 21724 755 21738
rect 23084 21724 23098 21738
rect 764 21700 778 21714
rect 23204 21700 23218 21714
rect 3500 18778 3514 18792
rect 419 17891 433 17905
rect 3500 17602 3514 17616
rect 442 16715 456 16729
rect 3500 16426 3514 16440
rect 465 15539 479 15553
rect 3500 15250 3514 15264
rect 488 14363 502 14377
rect 3500 14074 3514 14088
rect 511 13187 525 13201
rect 3500 12898 3514 12912
rect 534 12011 548 12025
rect 3500 11722 3514 11736
rect 557 10835 571 10849
rect 3500 10546 3514 10560
rect 580 9659 594 9673
rect 3500 9370 3514 9384
rect 603 8483 617 8497
rect 3500 8194 3514 8208
rect 626 7307 640 7321
rect 3500 7018 3514 7032
rect 649 6131 663 6145
rect 3500 5842 3514 5856
rect 672 4955 686 4969
rect 3500 4666 3514 4680
rect 695 3779 709 3793
rect 3500 3490 3514 3504
rect 718 2603 732 2617
rect 3500 2314 3514 2328
rect 741 1427 755 1441
rect 3500 1138 3514 1152
rect 764 251 778 265
rect 17684 70 17698 84
rect 20348 70 20362 84
rect 20395 70 20409 84
rect 20444 70 20458 84
rect 20492 70 20506 84
rect 20540 70 20554 84
rect 20588 70 20602 84
rect 20636 70 20650 84
rect 20684 70 20698 84
rect 20996 70 21010 84
rect 21044 70 21058 84
rect 21091 70 21105 84
rect 21140 70 21154 84
rect 21452 70 21466 84
rect 21500 70 21514 84
rect 21884 70 21898 84
rect 25245 70 25259 84
rect 975 49 989 63
rect 3740 48 3754 62
<< metal2 >>
rect 420 17905 432 22060
rect 443 16729 455 22036
rect 466 15553 478 22012
rect 489 14377 501 21988
rect 512 13201 524 21964
rect 535 12025 547 21940
rect 558 10849 570 21916
rect 581 9673 593 21892
rect 604 8497 616 21868
rect 627 7321 639 21844
rect 650 6145 662 21820
rect 673 4969 685 21796
rect 696 3793 708 21772
rect 719 2617 731 21748
rect 742 1441 754 21724
rect 765 265 777 21700
rect 789 21691 989 22218
rect 1005 21691 1017 22218
rect 1029 21691 1041 22218
rect 1053 21691 1065 22218
rect 1077 21691 1089 22218
rect 4317 21691 4329 22218
rect 4341 21691 4353 21940
rect 4389 21691 4401 21868
rect 4557 21691 4569 22218
rect 4773 21691 4785 21916
rect 4821 21691 4833 21844
rect 5205 21691 5217 21892
rect 5253 21691 5265 21820
rect 5613 21691 5625 22218
rect 5853 21691 5865 22218
rect 6983 21691 6995 22218
rect 7293 21691 7305 21748
rect 7317 21691 7329 21772
rect 7341 21691 7353 21796
rect 13221 21691 13233 22218
rect 13245 21691 13257 22061
rect 13437 21691 13449 22036
rect 13485 21691 13497 22218
rect 13629 21691 13641 22012
rect 13821 21691 13833 21988
rect 14013 21691 14025 21964
rect 14205 21691 14217 22218
rect 17757 21691 17769 22218
rect 17949 21691 17961 22218
rect 18021 21691 18033 22218
rect 18117 21691 18129 22218
rect 22773 21691 22785 21772
rect 22965 21691 22977 21747
rect 23085 21691 23097 21724
rect 23205 21691 23217 21700
rect 25244 21691 25444 22218
rect 24045 18885 24057 18908
rect 3501 18708 3513 18778
rect 24045 17709 24057 17843
rect 3501 17532 3513 17602
rect 24045 16533 24057 16667
rect 3501 16356 3513 16426
rect 24045 15357 24057 15491
rect 3501 15180 3513 15250
rect 24045 14181 24057 14315
rect 3501 14004 3513 14074
rect 24045 13005 24057 13139
rect 3501 12828 3513 12898
rect 24045 11829 24057 11963
rect 3501 11652 3513 11722
rect 24045 10653 24057 10787
rect 3501 10476 3513 10546
rect 24045 9477 24057 9611
rect 3501 9300 3513 9370
rect 24045 8301 24057 8435
rect 3501 8124 3513 8194
rect 24045 7125 24057 7259
rect 3501 6948 3513 7018
rect 24045 5949 24057 6083
rect 3501 5772 3513 5842
rect 24045 4773 24057 4907
rect 3501 4596 3513 4666
rect 24045 3597 24057 3731
rect 3501 3420 3513 3490
rect 24045 2421 24057 2555
rect 3501 2244 3513 2314
rect 24045 1245 24057 1379
rect 3501 1068 3513 1138
rect 789 63 989 92
rect 789 49 975 63
rect 789 0 989 49
rect 1005 0 1017 92
rect 1029 0 1041 92
rect 1053 0 1065 92
rect 1077 0 1089 92
rect 2349 0 2361 92
rect 2541 0 2553 92
rect 3333 0 3345 92
rect 3741 62 3753 92
rect 3885 0 3897 92
rect 4101 0 4113 92
rect 4845 0 4857 92
rect 5013 0 5025 92
rect 5397 0 5409 92
rect 5589 0 5601 103
rect 24045 92 24057 203
rect 5805 0 5817 92
rect 6549 0 6561 92
rect 6717 0 6729 92
rect 16125 0 16137 92
rect 16317 0 16329 92
rect 16557 0 16569 92
rect 17205 86 17217 92
rect 17397 86 17409 92
rect 17205 74 17409 86
rect 17685 84 17697 92
rect 20349 84 20361 92
rect 20397 84 20409 92
rect 20445 84 20457 92
rect 20493 84 20505 92
rect 20541 84 20553 92
rect 20589 84 20601 92
rect 20637 84 20649 92
rect 20685 84 20697 92
rect 20997 84 21009 92
rect 21045 84 21057 92
rect 21093 84 21105 92
rect 21141 84 21153 92
rect 21453 84 21465 92
rect 21501 84 21513 92
rect 21885 84 21897 92
rect 24261 0 24273 92
rect 25005 0 25017 92
rect 25245 84 25445 92
rect 25259 70 25445 84
rect 25245 0 25445 70
use slice17  slice17_0
timestamp 1394833348
transform 1 0 837 0 1 18908
box -48 0 24608 2783
use leftbuf_slice  leftbuf_slice_0
array 0 0 1685 0 15 1176
timestamp 1394551156
transform 1 0 784 0 1 98
box 0 -6 1685 1170
use IrAA  IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 2469 0 1 9611
box 0 -111 1008 1065
use tielow  tielow_0
timestamp 1386086605
transform 1 0 3477 0 1 17909
box 0 0 48 799
use tielow  tielow_1
timestamp 1386086605
transform 1 0 3477 0 1 16733
box 0 0 48 799
use tielow  tielow_2
timestamp 1386086605
transform 1 0 3477 0 1 15557
box 0 0 48 799
use tielow  tielow_3
timestamp 1386086605
transform 1 0 3477 0 1 14381
box 0 0 48 799
use tielow  tielow_4
timestamp 1386086605
transform 1 0 3477 0 1 13205
box 0 0 48 799
use tielow  tielow_5
timestamp 1386086605
transform 1 0 3477 0 1 12029
box 0 0 48 799
use tielow  tielow_6
timestamp 1386086605
transform 1 0 3477 0 1 10853
box 0 0 48 799
use tielow  tielow_7
timestamp 1386086605
transform 1 0 3477 0 1 9677
box 0 0 48 799
use IrBA  IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 2469 0 1 6083
box 0 -111 1008 1065
use tielow  tielow_8
timestamp 1386086605
transform 1 0 3477 0 1 8501
box 0 0 48 799
use tielow  tielow_9
timestamp 1386086605
transform 1 0 3477 0 1 7325
box 0 0 48 799
use tielow  tielow_10
timestamp 1386086605
transform 1 0 3477 0 1 6149
box 0 0 48 799
use IrBB  IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 2469 0 1 204
box 0 -112 1008 1064
use tiehigh  tiehigh_0
timestamp 1386086759
transform 1 0 3477 0 1 4973
box 0 0 48 799
use tielow  tielow_12
timestamp 1386086605
transform 1 0 3477 0 1 3797
box 0 0 48 799
use tielow  tielow_13
timestamp 1386086605
transform 1 0 3477 0 1 2621
box 0 0 48 799
use tielow  tielow_14
timestamp 1386086605
transform 1 0 3477 0 1 1445
box 0 0 48 799
use tielow  tielow_15
timestamp 1386086605
transform 1 0 3477 0 1 269
box 0 0 48 799
use Datapath_slice  Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394725603
transform 1 0 3525 0 1 92
box 0 0 20472 1176
use LLIcell_U  LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1394560148
transform 1 0 23997 0 1 9611
box 0 0 192 1042
use LLIcell_L  LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23997 0 1 203
box 0 0 192 1042
use Datapath_end  Datapath_end_0
array 0 0 1256 0 15 1176
timestamp 1394720841
transform 1 0 24189 0 1 92
box 0 0 1256 1176
<< labels >>
rlabel metal2 3885 0 3897 0 1 LrSel
rlabel metal2 4101 0 4113 0 1 LrWe
rlabel metal2 4845 0 4857 0 1 LrEn
rlabel metal2 5013 0 5025 0 1 PcSel[0]
rlabel metal2 5397 0 5409 0 1 PcSel[1]
rlabel metal1 24093 1257 24093 1257 1 Aluout[0]
rlabel metal2 24261 0 24273 0 1 AluWe
rlabel metal2 25005 0 25017 0 1 AluEn
rlabel metal2 25245 0 25445 0 1 GND!
rlabel metal2 22779 21767 22779 21767 1 Ir[3]
rlabel metal2 22970 21742 22970 21742 1 Ir[2]
rlabel metal2 23090 21717 23090 21717 1 Ir[1]
rlabel metal2 23211 21695 23211 21695 1 Ir[0]
rlabel metal2 17757 22218 17769 22218 5 Flags[2]
rlabel metal2 17949 22218 17961 22218 5 Flags[1]
rlabel metal2 18021 22218 18033 22218 5 Flags[3]
rlabel metal2 18117 22218 18129 22218 5 Flags[0]
rlabel metal2 25244 22218 25444 22218 1 GND!
rlabel metal1 -48 187 -48 197 3 SysBus[0]
rlabel metal1 -48 1363 -48 1373 3 SysBus[1]
rlabel metal1 -48 2539 -48 2549 3 SysBus[2]
rlabel metal1 -48 3715 -48 3725 3 SysBus[3]
rlabel metal1 -48 4891 -48 4901 3 SysBus[4]
rlabel metal1 -48 6067 -48 6077 3 SysBus[5]
rlabel metal1 -48 7243 -48 7253 3 SysBus[6]
rlabel metal1 -48 8419 -48 8429 3 SysBus[7]
rlabel metal1 -48 9595 -48 9605 3 SysBus[8]
rlabel metal1 -48 10771 -48 10781 3 SysBus[9]
rlabel metal1 -48 11947 -48 11957 3 SysBus[10]
rlabel metal1 -48 13123 -48 13133 3 SysBus[11]
rlabel metal1 -48 14299 -48 14309 3 SysBus[12]
rlabel metal1 -48 15475 -48 15485 3 SysBus[13]
rlabel metal1 -48 16651 -48 16661 3 SysBus[14]
rlabel metal1 -48 17827 -48 17837 3 SysBus[15]
rlabel metal1 -48 253 -48 263 3 Ir[0]
rlabel metal1 -48 1429 -48 1439 3 Ir[1]
rlabel metal1 -48 2605 -48 2615 3 Ir[2]
rlabel metal1 -48 3781 -48 3791 3 Ir[3]
rlabel metal1 -48 4957 -48 4967 3 Ir[4]
rlabel metal1 -48 6133 -48 6143 3 Ir[5]
rlabel metal1 -48 7309 -48 7319 3 Ir[6]
rlabel metal1 -48 8485 -48 8495 3 Ir[7]
rlabel metal1 -48 9661 -48 9671 3 Ir[8]
rlabel metal1 -48 10837 -48 10847 3 Ir[9]
rlabel metal1 -48 12013 -48 12023 3 Ir[10]
rlabel metal1 -48 13189 -48 13199 3 Ir[11]
rlabel metal1 -48 14365 -48 14375 3 Ir[12]
rlabel metal1 -48 15541 -48 15551 3 Ir[13]
rlabel metal1 -48 16717 -48 16727 3 Ir[14]
rlabel metal1 -48 17893 -48 17903 3 Ir[15]
rlabel metal2 789 0 989 0 1 Vdd!
rlabel metal2 1005 0 1017 0 1 SDI
rlabel metal2 1029 0 1041 0 1 Test
rlabel metal2 1053 0 1065 0 1 Clock
rlabel metal2 1077 0 1089 0 1 nReset
rlabel metal2 3333 0 3345 0 1 ImmSel
rlabel metal2 2541 0 2553 0 1 IrWe
rlabel metal1 -48 221 -48 231 3 DataIn[0]
rlabel metal1 -48 17861 -48 17871 3 DataIn[15]
rlabel metal1 -48 16685 -48 16695 3 DataIn[14]
rlabel metal1 -48 15509 -48 15519 3 DataIn[13]
rlabel metal1 -48 14333 -48 14343 3 DataIn[12]
rlabel metal1 -48 13157 -48 13167 3 DataIn[11]
rlabel metal1 -48 11981 -48 11991 3 DataIn[10]
rlabel metal1 -48 10805 -48 10815 3 DataIn[9]
rlabel metal1 -48 9629 -48 9639 3 DataIn[8]
rlabel metal1 -48 8453 -48 8463 3 DataIn[7]
rlabel metal1 -48 7277 -48 7287 3 DataIn[6]
rlabel metal1 -48 6101 -48 6111 3 DataIn[5]
rlabel metal1 -48 4925 -48 4935 3 DataIn[4]
rlabel metal1 -48 3749 -48 3759 3 DataIn[3]
rlabel metal1 -48 2573 -48 2583 3 DataIn[2]
rlabel metal1 -48 1397 -48 1407 3 DataIn[1]
rlabel metal2 2349 0 2361 0 1 MemEn
rlabel metal2 702 21769 702 21769 1 Ir[3]
rlabel metal2 679 21770 679 21770 1 Ir[4]
rlabel metal2 656 21769 656 21769 1 Ir[5]
rlabel metal2 633 21768 633 21768 1 Ir[6]
rlabel metal2 610 21767 610 21767 1 Ir[7]
rlabel metal2 587 21765 587 21765 1 Ir[8]
rlabel metal2 564 21765 564 21765 1 Ir[9]
rlabel metal2 541 21764 541 21764 1 Ir[10]
rlabel metal2 518 21765 518 21765 1 Ir[11]
rlabel metal2 495 21765 495 21765 1 Ir[12]
rlabel metal2 472 21764 472 21764 1 Ir[13]
rlabel metal2 449 21764 449 21764 1 Ir[14]
rlabel metal2 425 21765 425 21765 1 Ir[15]
rlabel metal2 1029 22218 1041 22218 1 Test
rlabel metal2 1053 22218 1065 22218 1 Clock
rlabel metal2 1077 22218 1089 22218 1 nReset
rlabel metal2 789 22218 989 22218 5 Vdd!
rlabel metal2 1005 22218 1017 22218 5 SDO
rlabel metal2 5805 0 5817 0 1 PcWe
rlabel metal2 5589 0 5601 0 1 PcSel[2]
rlabel metal2 6549 0 6561 0 1 PcEn
rlabel metal2 6717 0 6729 0 1 WdSel
rlabel metal2 6983 22218 6995 22218 5 RegWe
rlabel metal2 7297 21740 7297 21740 1 Ir[2]
rlabel metal2 7323 21764 7323 21764 1 Ir[3]
rlabel metal2 7346 21788 7346 21788 1 Ir[4]
rlabel metal2 4557 22218 4569 22218 5 Rs1Sel[1]
rlabel metal1 4798 21947 4798 21947 1 Ir[10]
rlabel metal2 5613 22218 5625 22218 5 RwSel[0]
rlabel metal2 5853 22218 5865 22218 5 RwSel[1]
rlabel metal2 4778 21908 4778 21908 1 Ir[9]
rlabel metal2 4827 21837 4827 21837 1 Ir[6]
rlabel metal2 5210 21885 5210 21885 1 Ir[8]
rlabel metal2 5260 21814 5260 21814 1 Ir[5]
rlabel metal2 4317 22218 4329 22218 5 Rs1Sel[0]
rlabel metal2 4346 21933 4346 21933 1 Ir[10]
rlabel metal2 4395 21860 4395 21860 1 Ir[7]
rlabel metal2 16125 0 16137 0 1 Op1Sel
rlabel metal2 16317 0 16329 0 1 Op2Sel[0]
rlabel metal2 16557 0 16569 0 1 Op2Sel[1]
rlabel metal2 14205 22218 14217 22218 5 CFlag
rlabel metal2 13250 22054 13250 22054 1 Ir[15]
rlabel metal2 13441 22029 13441 22029 1 Ir[14]
rlabel metal2 14019 21957 14019 21957 1 Ir[11]
rlabel metal2 13827 21982 13827 21982 1 Ir[12]
rlabel metal2 13634 22006 13634 22006 1 Ir[13]
rlabel metal2 13221 22218 13233 22218 5 AluOR[1]
rlabel metal2 13485 22218 13497 22218 5 AluOR[0]
<< end >>
