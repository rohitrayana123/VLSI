magic
tech c035u
timestamp 1394128665
<< metal1 >>
rect 4405 1025 5927 1035
rect 3997 1003 5519 1013
rect 3541 981 5063 991
rect 5102 980 5495 990
rect 5509 980 5903 990
rect 5917 981 6263 991
rect 3517 958 3959 968
rect 3973 958 4367 968
rect 4381 958 4727 968
rect 4765 959 6287 969
rect 397 936 599 946
rect 661 938 791 948
rect 3589 936 3791 946
rect 4045 936 4199 946
rect 4453 936 4559 946
rect 5125 936 5327 946
rect 5581 936 5735 946
rect 5989 937 6095 947
rect 6349 936 6407 946
rect 229 914 527 924
rect 637 914 647 924
rect 733 913 863 923
rect 877 914 1007 924
rect 1309 914 1343 924
rect 1645 914 1703 924
rect 2053 914 2111 924
rect 2389 914 2447 924
rect 2725 914 2759 924
rect 3061 914 3095 924
rect 3637 914 3647 924
rect 3685 914 3695 924
rect 3733 914 3743 924
rect 4093 914 4103 924
rect 4141 914 4151 924
rect 4501 914 4511 924
rect 4813 917 4871 927
rect 5053 914 5087 924
rect 5149 914 5159 924
rect 5197 914 5207 924
rect 5245 914 5255 924
rect 5293 914 5399 924
rect 5605 914 5615 924
rect 5653 914 5663 924
rect 5701 914 5807 924
rect 6013 915 6023 925
rect 6061 914 6167 924
rect 6373 914 6479 924
rect 0 892 263 902
rect 277 892 1247 902
rect 1261 892 1583 902
rect 1597 892 1943 902
rect 1957 892 2687 902
rect 2701 892 2999 902
rect 3013 892 3407 902
rect 3421 892 6768 902
rect 0 870 143 880
rect 157 870 1223 880
rect 1237 870 1559 880
rect 1573 870 1919 880
rect 1933 870 2327 880
rect 2341 870 2663 880
rect 2677 870 2975 880
rect 2989 870 3287 880
rect 3301 870 3359 880
rect 3445 870 3599 880
rect 3613 870 3815 880
rect 3901 870 4055 880
rect 4069 870 4223 880
rect 4309 870 4463 880
rect 4477 870 4583 880
rect 4669 870 4895 880
rect 4981 870 5351 880
rect 5437 870 5759 880
rect 5846 870 6119 880
rect 6205 870 6431 880
rect 6517 870 6575 880
rect 85 51 167 61
rect 901 44 935 54
rect 1165 51 1487 61
rect 1501 51 1847 61
rect 1861 51 2255 61
rect 2269 51 2591 61
rect 2605 51 2903 61
rect 2917 51 3239 61
rect 3253 51 6719 61
rect 6733 51 6768 61
rect 3613 29 3623 39
rect 3661 29 3671 39
rect 3709 29 3719 39
rect 3757 29 3863 39
rect 4069 29 4079 39
rect 4117 29 4127 39
rect 4165 29 4271 39
rect 4477 29 4487 39
rect 4525 29 4631 39
rect 4909 29 4943 39
rect 5053 29 5088 39
rect 5173 29 5183 39
rect 5221 29 5231 39
rect 5269 29 5279 39
rect 5629 29 5639 39
rect 5677 29 5687 39
rect 6037 29 6047 39
rect 6373 29 6431 39
rect 5149 7 5351 17
rect 5605 7 5759 17
rect 6013 7 6119 17
<< m2contact >>
rect 4391 1023 4405 1037
rect 5927 1023 5941 1037
rect 3983 1001 3997 1015
rect 5519 1001 5533 1015
rect 3527 978 3541 992
rect 5063 979 5077 993
rect 5088 979 5102 993
rect 5495 979 5509 993
rect 5903 979 5917 993
rect 6263 979 6277 993
rect 3503 956 3517 970
rect 3959 956 3973 970
rect 4367 956 4381 970
rect 4727 956 4741 970
rect 4751 956 4765 970
rect 6287 957 6301 971
rect 383 935 397 949
rect 599 934 613 948
rect 647 936 661 950
rect 791 936 805 950
rect 3575 934 3589 948
rect 3791 934 3805 948
rect 4031 934 4045 948
rect 4199 934 4213 948
rect 4439 934 4453 948
rect 4559 934 4573 948
rect 5111 934 5125 948
rect 5327 934 5341 948
rect 5567 934 5581 948
rect 5735 934 5749 948
rect 5975 935 5989 949
rect 6095 935 6109 949
rect 6335 934 6349 948
rect 6407 934 6421 948
rect 215 912 229 926
rect 527 912 541 926
rect 623 912 637 926
rect 647 912 661 926
rect 719 912 733 926
rect 863 912 877 926
rect 1007 912 1021 926
rect 1295 912 1309 926
rect 1343 912 1357 926
rect 1631 912 1645 926
rect 1703 912 1717 926
rect 2039 912 2053 926
rect 2111 912 2125 926
rect 2375 912 2389 926
rect 2447 912 2461 926
rect 2711 912 2725 926
rect 2759 912 2773 926
rect 3047 912 3061 926
rect 3095 912 3109 926
rect 3623 912 3637 926
rect 3647 912 3661 926
rect 3671 912 3685 926
rect 3695 912 3709 926
rect 3719 912 3733 926
rect 3743 912 3757 926
rect 4079 912 4093 926
rect 4103 912 4117 926
rect 4127 912 4141 926
rect 4151 912 4165 926
rect 4487 912 4501 926
rect 4511 912 4525 926
rect 4799 916 4813 930
rect 4871 916 4885 930
rect 5039 912 5053 926
rect 5087 912 5101 926
rect 5135 912 5149 926
rect 5159 912 5173 926
rect 5183 912 5197 926
rect 5207 912 5221 926
rect 5231 912 5245 926
rect 5255 912 5269 926
rect 5279 912 5293 926
rect 5399 912 5413 926
rect 5591 912 5605 926
rect 5615 912 5629 926
rect 5639 912 5653 926
rect 5663 912 5677 926
rect 5687 912 5701 926
rect 5807 912 5821 926
rect 5999 913 6013 927
rect 6023 913 6037 927
rect 6047 913 6061 927
rect 6167 912 6181 926
rect 6359 912 6373 926
rect 6479 912 6493 926
rect 263 890 277 904
rect 1247 890 1261 904
rect 1583 890 1597 904
rect 1943 890 1957 904
rect 2687 890 2701 904
rect 2999 890 3013 904
rect 3407 890 3421 904
rect 143 868 157 882
rect 1223 868 1237 882
rect 1559 868 1573 882
rect 1919 868 1933 882
rect 2327 868 2341 882
rect 2663 868 2677 882
rect 2975 868 2989 882
rect 3287 868 3301 882
rect 3359 868 3373 882
rect 3431 868 3445 882
rect 3599 868 3613 882
rect 3815 868 3829 882
rect 3887 868 3901 882
rect 4055 868 4069 882
rect 4223 868 4237 882
rect 4295 868 4309 882
rect 4463 868 4477 882
rect 4583 868 4597 882
rect 4655 868 4669 882
rect 4895 868 4909 882
rect 4967 868 4981 882
rect 5351 868 5365 882
rect 5423 868 5437 882
rect 5759 868 5773 882
rect 5832 868 5846 882
rect 6119 868 6133 882
rect 6191 868 6205 882
rect 6431 868 6445 882
rect 6503 868 6517 882
rect 6575 868 6589 882
rect 71 49 85 63
rect 167 49 181 63
rect 887 42 901 56
rect 935 42 949 56
rect 1151 49 1165 63
rect 1487 49 1501 63
rect 1847 49 1861 63
rect 2255 49 2269 63
rect 2591 49 2605 63
rect 2903 49 2917 63
rect 3239 49 3253 63
rect 6719 49 6733 63
rect 3599 27 3613 41
rect 3623 27 3637 41
rect 3647 27 3661 41
rect 3671 27 3685 41
rect 3695 27 3709 41
rect 3719 27 3733 41
rect 3743 27 3757 41
rect 3863 27 3877 41
rect 4055 27 4069 41
rect 4079 27 4093 41
rect 4103 27 4117 41
rect 4127 27 4141 41
rect 4151 27 4165 41
rect 4271 27 4285 41
rect 4463 27 4477 41
rect 4487 27 4501 41
rect 4511 27 4525 41
rect 4631 27 4645 41
rect 4895 27 4909 41
rect 4943 27 4957 41
rect 5039 27 5053 41
rect 5088 27 5102 41
rect 5159 27 5173 41
rect 5183 27 5197 41
rect 5207 27 5221 41
rect 5231 27 5245 41
rect 5255 27 5269 41
rect 5279 27 5293 41
rect 5615 27 5629 41
rect 5639 27 5653 41
rect 5663 27 5677 41
rect 5687 27 5701 41
rect 6023 27 6037 41
rect 6047 27 6061 41
rect 6359 27 6373 41
rect 6431 27 6445 41
rect 5135 5 5149 19
rect 5351 5 5365 19
rect 5591 5 5605 19
rect 5759 5 5773 19
rect 5999 5 6013 19
rect 6119 5 6133 19
<< metal2 >>
rect 24 865 36 1042
rect 144 865 156 868
rect 216 865 228 912
rect 264 865 276 890
rect 288 865 300 1042
rect 384 865 396 935
rect 456 865 468 1042
rect 528 865 540 912
rect 600 865 612 934
rect 624 926 636 1042
rect 648 950 660 1042
rect 720 926 732 1042
rect 648 865 660 912
rect 720 865 732 912
rect 792 865 804 936
rect 864 865 876 912
rect 936 865 948 1042
rect 1008 865 1020 912
rect 1080 865 1092 1042
rect 1224 865 1236 868
rect 1248 865 1260 890
rect 1296 865 1308 912
rect 1344 865 1356 912
rect 1416 865 1428 1042
rect 1560 865 1572 868
rect 1584 865 1596 890
rect 1632 865 1644 912
rect 1704 865 1716 912
rect 1776 865 1788 1042
rect 1920 865 1932 868
rect 1944 865 1956 890
rect 2040 865 2052 912
rect 2112 865 2124 912
rect 2184 865 2196 1042
rect 2328 865 2340 868
rect 2376 865 2388 912
rect 2448 865 2460 912
rect 2520 865 2532 1042
rect 2664 865 2676 868
rect 2688 865 2700 890
rect 2712 865 2724 912
rect 2760 865 2772 912
rect 2832 865 2844 1042
rect 2976 865 2988 868
rect 3000 865 3012 890
rect 3048 865 3060 912
rect 3096 865 3108 912
rect 3168 865 3180 1042
rect 3288 882 3300 1042
rect 3336 865 3348 1042
rect 3504 970 3516 1042
rect 3360 865 3372 868
rect 3408 865 3420 890
rect 3432 865 3444 868
rect 3504 865 3516 956
rect 3528 865 3540 978
rect 3576 865 3588 934
rect 3600 882 3612 1042
rect 3648 926 3660 1042
rect 3696 926 3708 1042
rect 3744 926 3756 1042
rect 3624 865 3636 912
rect 3672 865 3684 912
rect 3720 865 3732 912
rect 3792 865 3804 934
rect 3816 865 3828 868
rect 3888 865 3900 868
rect 3960 865 3972 956
rect 3984 865 3996 1001
rect 4032 865 4044 934
rect 4056 882 4068 1042
rect 4104 926 4116 1042
rect 4152 926 4164 1042
rect 4080 865 4092 912
rect 4128 865 4140 912
rect 4200 865 4212 934
rect 4224 865 4236 868
rect 4296 865 4308 868
rect 4368 865 4380 956
rect 4392 865 4404 1023
rect 4440 865 4452 934
rect 4464 882 4476 1042
rect 4512 926 4524 1042
rect 4488 865 4500 912
rect 4560 865 4572 934
rect 4584 865 4596 868
rect 4656 865 4668 868
rect 4728 865 4740 956
rect 4752 865 4764 956
rect 4800 865 4812 916
rect 4872 865 4884 916
rect 4896 882 4908 1042
rect 5064 993 5076 1042
rect 5089 993 5101 1042
rect 4896 865 4908 868
rect 4968 865 4980 868
rect 5040 865 5052 912
rect 5064 865 5076 979
rect 5089 926 5101 979
rect 5112 865 5124 934
rect 5136 926 5148 1042
rect 5184 926 5196 1042
rect 5232 926 5244 1042
rect 5280 926 5292 1042
rect 5520 1015 5532 1042
rect 5160 865 5172 912
rect 5208 865 5220 912
rect 5256 865 5268 912
rect 5328 865 5340 934
rect 5352 865 5364 868
rect 5400 865 5412 912
rect 5424 865 5436 868
rect 5496 865 5508 979
rect 5520 865 5532 1001
rect 5568 865 5580 934
rect 5592 926 5604 1042
rect 5640 926 5652 1042
rect 5688 926 5700 1042
rect 5928 1037 5940 1042
rect 5616 865 5628 912
rect 5664 865 5676 912
rect 5736 865 5748 934
rect 5760 865 5772 868
rect 5808 865 5820 912
rect 5832 865 5844 868
rect 5904 865 5916 979
rect 5928 865 5940 1023
rect 5976 865 5988 935
rect 6000 927 6012 1042
rect 6048 927 6060 1042
rect 6024 865 6036 913
rect 6096 865 6108 935
rect 6120 865 6132 868
rect 6168 865 6180 912
rect 6192 865 6204 868
rect 6264 865 6276 979
rect 6288 971 6300 1042
rect 6288 865 6300 957
rect 6336 865 6348 934
rect 6360 926 6372 1042
rect 6408 865 6420 934
rect 6432 865 6444 868
rect 6480 865 6492 912
rect 6504 865 6516 868
rect 6576 865 6588 868
rect 6648 865 6660 1042
rect 24 0 36 66
rect 72 63 84 66
rect 168 63 180 66
rect 288 0 300 66
rect 456 0 468 66
rect 648 0 660 66
rect 888 56 900 66
rect 936 0 948 42
rect 1080 0 1092 66
rect 1152 63 1164 66
rect 1416 0 1428 66
rect 1488 63 1500 66
rect 1776 0 1788 66
rect 1848 63 1860 66
rect 2184 0 2196 66
rect 2256 63 2268 66
rect 2520 0 2532 66
rect 2592 63 2604 66
rect 2832 0 2844 66
rect 2904 63 2916 66
rect 3168 0 3180 66
rect 3240 63 3252 66
rect 3336 0 3348 66
rect 3504 0 3516 66
rect 3624 41 3636 66
rect 3672 41 3684 66
rect 3720 41 3732 66
rect 3864 41 3876 66
rect 4080 41 4092 66
rect 4128 41 4140 66
rect 4272 41 4284 66
rect 4488 41 4500 66
rect 4632 41 4644 66
rect 4944 41 4956 66
rect 5040 41 5052 66
rect 3600 0 3612 27
rect 3648 0 3660 27
rect 3696 0 3708 27
rect 3744 0 3756 27
rect 4056 0 4068 27
rect 4104 0 4116 27
rect 4152 0 4164 27
rect 4464 0 4476 27
rect 4512 0 4524 27
rect 4896 0 4908 27
rect 5064 0 5076 66
rect 5160 41 5172 66
rect 5208 41 5220 66
rect 5256 41 5268 66
rect 5089 0 5101 27
rect 5136 0 5148 5
rect 5184 0 5196 27
rect 5232 0 5244 27
rect 5280 0 5292 27
rect 5352 19 5364 66
rect 5520 0 5532 66
rect 5616 41 5628 66
rect 5664 41 5676 66
rect 5592 0 5604 5
rect 5640 0 5652 27
rect 5688 0 5700 27
rect 5760 19 5772 66
rect 5928 0 5940 66
rect 6024 41 6036 66
rect 6000 0 6012 5
rect 6048 0 6060 27
rect 6120 19 6132 66
rect 6288 0 6300 66
rect 6432 41 6444 66
rect 6360 0 6372 27
rect 6648 0 6660 66
rect 6720 63 6732 66
use inv inv_1
timestamp 1386238110
transform 1 0 0 0 1 66
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 120 0 1 66
box 0 0 120 799
use xor2 xor2_0
timestamp 1386237344
transform 1 0 240 0 1 66
box 0 0 192 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 432 0 1 66
box 0 0 48 799
use fulladder fulladder_0
timestamp 1386234928
transform 1 0 480 0 1 66
box 0 0 360 799
use or2 or2_0
timestamp 1386235472
transform 1 0 840 0 1 66
box 0 0 144 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 984 0 1 66
box 0 0 216 799
use and2 and2_1
timestamp 1386234845
transform 1 0 1200 0 1 66
box 0 0 120 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 1320 0 1 66
box 0 0 216 799
use or2 or2_1
timestamp 1386235472
transform 1 0 1536 0 1 66
box 0 0 144 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1680 0 1 66
box 0 0 216 799
use xor2 xor2_1
timestamp 1386237344
transform 1 0 1896 0 1 66
box 0 0 192 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2088 0 1 66
box 0 0 216 799
use inv inv_0
timestamp 1386238110
transform 1 0 2304 0 1 66
box 0 0 120 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 2424 0 1 66
box 0 0 216 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 2640 0 1 66
box 0 0 96 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 2736 0 1 66
box 0 0 216 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 2952 0 1 66
box 0 0 120 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 3072 0 1 66
box 0 0 216 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 3288 0 1 66
box 0 0 192 799
use and2 and2_2
timestamp 1386234845
transform 1 0 3480 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 3600 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_2
timestamp 1386086759
transform 1 0 3648 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_3
timestamp 1386086759
transform 1 0 3696 0 1 66
box 0 0 48 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 3744 0 1 66
box 0 0 192 799
use and2 and2_3
timestamp 1386234845
transform 1 0 3936 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_7
timestamp 1386086759
transform 1 0 4056 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_10
timestamp 1386086759
transform 1 0 4104 0 1 66
box 0 0 48 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4152 0 1 66
box 0 0 192 799
use and2 and2_4
timestamp 1386234845
transform 1 0 4344 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_9
timestamp 1386086759
transform 1 0 4464 0 1 66
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 4512 0 1 66
box 0 0 192 799
use and2 and2_5
timestamp 1386234845
transform 1 0 4704 0 1 66
box 0 0 120 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 4824 0 1 66
box 0 0 192 799
use and2 and2_6
timestamp 1386234845
transform 1 0 5016 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_4
timestamp 1386086759
transform 1 0 5136 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_5
timestamp 1386086759
transform 1 0 5184 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_6
timestamp 1386086759
transform 1 0 5232 0 1 66
box 0 0 48 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 5280 0 1 66
box 0 0 192 799
use and2 and2_7
timestamp 1386234845
transform 1 0 5472 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_11
timestamp 1386086759
transform 1 0 5592 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_12
timestamp 1386086759
transform 1 0 5640 0 1 66
box 0 0 48 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 5688 0 1 66
box 0 0 192 799
use and2 and2_8
timestamp 1386234845
transform 1 0 5880 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_15
timestamp 1386086759
transform 1 0 6000 0 1 66
box 0 0 48 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 6048 0 1 66
box 0 0 192 799
use and2 and2_9
timestamp 1386234845
transform 1 0 6240 0 1 66
box 0 0 120 799
use mux2 mux2_8
timestamp 1386235218
transform 1 0 6360 0 1 66
box 0 0 192 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 6552 0 1 66
box 0 0 216 799
<< labels >>
rlabel metal2 648 0 660 0 1 CIn_Slice
rlabel metal2 624 1042 636 1042 5 CIn_Slice
rlabel metal2 936 0 948 0 1 nZ_prev
rlabel metal1 6768 51 6768 61 7 ALUOut
rlabel metal2 6288 0 6300 0 1 Sh1
rlabel metal2 5928 0 5940 0 1 Sh2
rlabel metal2 5520 0 5532 0 1 Sh4
rlabel metal2 5064 0 5076 0 1 Sh8
rlabel metal2 288 0 300 0 1 SUB
rlabel metal2 3336 0 3348 0 1 ShB
rlabel metal2 6648 0 6660 0 1 ShOut
rlabel metal2 5089 0 5101 0 1 ShR
rlabel metal2 3504 0 3516 0 1 ShL
rlabel metal2 3168 0 3180 0 1 NOR
rlabel metal2 2832 0 2844 0 1 NAND
rlabel metal2 2520 0 2532 0 1 NOT
rlabel metal2 2184 0 2196 0 1 XOR
rlabel metal2 1776 0 1788 0 1 OR
rlabel metal2 1416 0 1428 0 1 AND
rlabel metal2 456 0 468 0 1 CIn
rlabel metal2 1080 0 1092 0 1 FAOut
rlabel metal2 3504 1042 3516 1042 5 ShL
rlabel metal2 5089 1042 5101 1042 5 ShR
rlabel metal2 4464 1042 4476 1042 5 Sh2A_L
rlabel metal2 4512 1042 4524 1042 5 Sh2B_L
rlabel metal2 3600 1042 3612 1042 5 Sh8A_L
rlabel metal2 3648 1042 3660 1042 5 Sh8B_L
rlabel metal2 3696 1042 3708 1042 5 Sh8C_L
rlabel metal2 3744 1042 3756 1042 5 Sh8D_L
rlabel metal2 4056 1042 4068 1042 5 Sh4A_L
rlabel metal2 4104 1042 4116 1042 5 Sh4B_L
rlabel metal2 4152 1042 4164 1042 5 Sh4C_L
rlabel metal2 5136 1042 5148 1042 5 Sh8A_R
rlabel metal2 5184 1042 5196 1042 5 Sh8B_R
rlabel metal2 5232 1042 5244 1042 5 Sh8C_R
rlabel metal2 5592 1042 5604 1042 5 Sh4A_R
rlabel metal2 5640 1042 5652 1042 5 Sh4B_R
rlabel metal2 5688 1042 5700 1042 5 Sh4C_R
rlabel metal2 6000 1042 6012 1042 5 Sh2A_R
rlabel metal2 6048 1042 6060 1042 5 Sh2B_R
rlabel metal2 6648 1042 6660 1042 5 ShOut
rlabel metal2 5280 1042 5292 1042 5 Sh8D_R
rlabel metal2 5064 1042 5076 1042 5 Sh8
rlabel metal2 5520 1042 5532 1042 5 Sh4
rlabel metal2 5928 1042 5940 1042 5 Sh2
rlabel metal2 6288 1042 6300 1042 5 Sh1
rlabel metal2 1080 1042 1092 1042 5 FAOut
rlabel metal2 936 1042 948 1042 5 nZ
rlabel metal2 288 1042 300 1042 5 SUB
rlabel metal2 1416 1042 1428 1042 5 AND
rlabel metal2 1776 1042 1788 1042 5 OR
rlabel metal2 2184 1042 2196 1042 5 XOR
rlabel metal2 2520 1042 2532 1042 5 NOT
rlabel metal2 2832 1042 2844 1042 5 NAND
rlabel metal2 3168 1042 3180 1042 5 NOR
rlabel metal2 3336 1042 3348 1042 5 ShB
rlabel metal2 648 1042 660 1042 5 COut
rlabel metal2 720 1042 732 1042 5 Sum
rlabel metal2 456 1042 468 1042 5 CIn
rlabel metal2 3288 1042 3300 1042 5 A
rlabel metal2 4464 0 4476 0 1 Sh2B_L
rlabel metal2 4512 0 4524 0 1 Sh2C_L
rlabel metal2 3600 0 3612 0 1 Sh8B_L
rlabel metal2 3648 0 3660 0 1 Sh8C_L
rlabel metal2 3696 0 3708 0 1 Sh8D_L
rlabel metal2 3744 0 3756 0 1 Sh8E_L
rlabel metal2 4056 0 4068 0 1 Sh4B_L
rlabel metal2 4104 0 4116 0 1 Sh4C_L
rlabel metal2 4152 0 4164 0 1 Sh4D_L
rlabel metal2 5280 0 5292 0 1 Sh8C_R
rlabel metal2 5232 0 5244 0 1 Sh8B_R
rlabel metal2 5184 0 5196 0 1 Sh8A_R
rlabel metal2 5136 0 5148 0 1 Sh8Z_R
rlabel metal2 5688 0 5700 0 1 Sh4B_R
rlabel metal2 5640 0 5652 0 1 Sh4A_R
rlabel metal2 5592 0 5604 0 1 Sh4Z_R
rlabel metal2 6000 0 6012 0 1 Sh2Z_R
rlabel metal2 6048 0 6060 0 1 Sh2A_R
rlabel metal2 4896 0 4908 0 1 Sh1_L_In
rlabel metal2 4896 1042 4908 1042 5 Sh1_L_Out
rlabel metal2 6360 0 6372 0 1 Sh1_R_Out
rlabel metal2 6360 1042 6372 1042 5 Sh1_R_In
rlabel metal1 509 917 509 917 1 FA_1
rlabel metal1 586 941 586 941 1 FA_2
rlabel metal2 24 0 36 0 1 ZeroA
rlabel metal2 24 1042 36 1042 5 ZeroA
rlabel metal1 6768 892 6768 902 7 B
rlabel metal1 0 892 0 902 3 B
rlabel metal1 0 870 0 880 3 A
<< end >>
