../../../Design/Implementation/verilog/behavioural/options.sv