magic
tech c035u
timestamp 1394209539
use slice17 slice17_0
timestamp 1394209539
transform 1 0 50 0 1 8600
box 0 0 9108 1618
use regBlock_slice regBlock_slice_0
array 0 0 9385 0 7 1075
timestamp 1394121372
transform 1 0 0 0 1 0
box 0 0 9385 1075
<< end >>
