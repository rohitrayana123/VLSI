magic
tech c035u
timestamp 1396383839
<< checkpaint >>
rect 0 0 26708 21542
rect 20800 -1300 26708 0
<< metal1 >>
rect 14 20182 14577 20192
rect 37 20158 14770 20168
rect 60 20134 14962 20144
rect 83 20110 15154 20120
rect 106 20086 15346 20096
rect 129 20062 4161 20072
rect 152 20038 4593 20048
rect 175 20014 4977 20024
rect 198 19990 4209 20000
rect 221 19966 4641 19976
rect 244 19942 5025 19952
rect 267 19918 7165 19928
rect 290 19894 7141 19904
rect 7155 19894 22353 19904
rect 313 19870 7117 19880
rect 7131 19870 22545 19880
rect 336 19846 22665 19856
rect 359 19822 22785 19832
rect 3095 18363 3106 18373
rect 14 17476 365 17486
rect 3058 17409 3106 17419
rect 25391 17409 25408 17419
rect 3058 17387 3106 17397
rect 3058 17365 3106 17375
rect 25391 17365 25408 17375
rect 3095 17209 3106 17219
rect 37 16322 365 16332
rect 3058 16255 3106 16265
rect 25391 16255 25408 16265
rect 3058 16233 3106 16243
rect 3058 16211 3106 16221
rect 25391 16211 25408 16221
rect 3095 16055 3106 16065
rect 60 15168 365 15178
rect 3058 15101 3106 15111
rect 25391 15101 25408 15111
rect 3058 15079 3106 15089
rect 3058 15057 3106 15067
rect 25391 15057 25408 15067
rect 3095 14901 3106 14911
rect 83 14014 365 14024
rect 3058 13947 3106 13957
rect 25391 13947 25408 13957
rect 3058 13925 3106 13935
rect 3058 13903 3106 13913
rect 25391 13903 25408 13913
rect 3095 13747 3106 13757
rect 106 12860 365 12870
rect 3058 12793 3106 12803
rect 25391 12793 25408 12803
rect 3058 12771 3106 12781
rect 3058 12749 3106 12759
rect 25391 12749 25408 12759
rect 3095 12593 3106 12603
rect 129 11706 365 11716
rect 3058 11639 3106 11649
rect 25391 11639 25408 11649
rect 3058 11617 3106 11627
rect 3058 11595 3106 11605
rect 25391 11595 25408 11605
rect 3095 11439 3106 11449
rect 152 10552 365 10562
rect 3058 10485 3106 10495
rect 25391 10485 25408 10495
rect 3058 10463 3106 10473
rect 3058 10441 3106 10451
rect 25391 10441 25408 10451
rect 3095 10285 3106 10295
rect 175 9398 365 9408
rect 3058 9331 3106 9341
rect 25391 9331 25408 9341
rect 3058 9309 3106 9319
rect 3058 9287 3106 9297
rect 25391 9287 25408 9297
rect 3095 9131 3106 9141
rect 198 8244 365 8254
rect 3058 8177 3106 8187
rect 25391 8177 25408 8187
rect 3058 8155 3106 8165
rect 3058 8133 3106 8143
rect 25391 8133 25408 8143
rect 3095 7977 3106 7987
rect 221 7090 365 7100
rect 3058 7023 3106 7033
rect 25391 7023 25408 7033
rect 3058 7001 3106 7011
rect 3058 6979 3106 6989
rect 25391 6979 25408 6989
rect 3095 6823 3106 6833
rect 244 5936 365 5946
rect 3058 5869 3106 5879
rect 25391 5869 25408 5879
rect 3058 5847 3106 5857
rect 3058 5825 3106 5835
rect 25391 5825 25408 5835
rect 3095 5669 3106 5679
rect 267 4782 365 4792
rect 3058 4715 3106 4725
rect 25391 4715 25408 4725
rect 3058 4693 3106 4703
rect 3058 4671 3106 4681
rect 25391 4671 25408 4681
rect 3095 4515 3106 4525
rect 290 3628 365 3638
rect 3058 3561 3106 3571
rect 25391 3561 25408 3571
rect 3058 3539 3106 3549
rect 3058 3517 3106 3527
rect 25391 3517 25408 3527
rect 3095 3361 3106 3371
rect 313 2474 365 2484
rect 3058 2407 3106 2417
rect 25391 2407 25408 2417
rect 3058 2385 3106 2395
rect 3058 2363 3106 2373
rect 25391 2363 25408 2373
rect 3095 2207 3106 2217
rect 336 1320 365 1330
rect 3058 1253 3106 1263
rect 25391 1253 25408 1263
rect 3058 1231 3106 1241
rect 3058 1209 3106 1219
rect 25391 1209 25408 1219
rect 3095 1053 3106 1063
rect 359 166 365 176
rect 3058 99 3106 109
rect 25391 99 25408 109
rect 3058 77 3106 87
rect 3058 55 3106 65
rect 25391 55 25408 65
rect 570 8 3321 18
rect 17279 7 19929 17
rect 19943 7 19976 17
rect 19990 7 20025 17
rect 20039 7 20073 17
rect 20087 7 20121 17
rect 20135 7 20169 17
rect 20183 7 20217 17
rect 20231 7 20265 17
rect 20279 7 20577 17
rect 20591 7 20625 17
rect 20639 7 20672 17
rect 20686 7 20721 17
rect 20735 7 21033 17
rect 21047 7 21081 17
rect 21095 7 21465 17
rect 21479 7 25186 17
<< m2contact >>
rect 0 20180 14 20194
rect 14577 20181 14591 20195
rect 23 20156 37 20170
rect 14770 20156 14784 20170
rect 46 20132 60 20146
rect 14962 20132 14976 20146
rect 69 20108 83 20122
rect 15154 20108 15168 20122
rect 92 20084 106 20098
rect 15346 20084 15360 20099
rect 115 20060 129 20074
rect 4161 20060 4175 20074
rect 138 20036 152 20050
rect 4593 20036 4607 20050
rect 161 20012 175 20026
rect 4977 20012 4991 20026
rect 184 19988 198 20002
rect 4209 19988 4223 20002
rect 207 19964 221 19978
rect 4641 19964 4655 19978
rect 230 19940 244 19954
rect 5025 19940 5039 19954
rect 253 19916 267 19930
rect 7165 19916 7179 19930
rect 276 19892 290 19906
rect 7141 19892 7155 19906
rect 22353 19892 22367 19906
rect 299 19868 313 19882
rect 7117 19868 7131 19882
rect 22545 19867 22559 19881
rect 322 19844 336 19858
rect 22665 19844 22679 19858
rect 345 19820 359 19834
rect 22785 19820 22799 19834
rect 3081 18361 3095 18375
rect 0 17474 14 17488
rect 3081 17207 3095 17221
rect 23 16320 37 16334
rect 3081 16053 3095 16067
rect 46 15166 60 15180
rect 3081 14899 3095 14913
rect 69 14012 83 14026
rect 3081 13745 3095 13759
rect 92 12858 106 12872
rect 3081 12591 3095 12605
rect 115 11704 129 11718
rect 3081 11437 3095 11451
rect 138 10550 152 10564
rect 3081 10283 3095 10297
rect 161 9396 175 9410
rect 3081 9129 3095 9143
rect 184 8242 198 8256
rect 3081 7975 3095 7989
rect 207 7088 221 7102
rect 3081 6821 3095 6835
rect 230 5934 244 5948
rect 3081 5667 3095 5681
rect 253 4780 267 4794
rect 3081 4513 3095 4527
rect 276 3626 290 3640
rect 3081 3359 3095 3373
rect 299 2472 313 2486
rect 3081 2205 3095 2219
rect 322 1318 336 1332
rect 3081 1051 3095 1065
rect 345 164 359 178
rect 556 6 570 20
rect 3321 5 3335 19
rect 17265 5 17279 19
rect 19929 5 19943 19
rect 19976 5 19990 19
rect 20025 5 20039 19
rect 20073 5 20087 19
rect 20121 5 20135 19
rect 20169 5 20183 19
rect 20217 5 20231 19
rect 20265 5 20279 19
rect 20577 5 20591 19
rect 20625 5 20639 19
rect 20672 5 20686 19
rect 20721 5 20735 19
rect 21033 5 21047 19
rect 21081 5 21095 19
rect 21465 5 21479 19
rect 25186 5 25200 19
<< metal2 >>
rect 1 17488 13 20180
rect 1 0 13 17474
rect 24 16334 36 20156
rect 24 0 36 16320
rect 47 15180 59 20132
rect 47 0 59 15166
rect 70 14026 82 20108
rect 70 0 82 14012
rect 93 12872 105 20084
rect 93 0 105 12858
rect 116 11718 128 20060
rect 116 0 128 11704
rect 139 10564 151 20036
rect 139 0 151 10550
rect 162 9410 174 20012
rect 162 0 174 9396
rect 185 8256 197 19988
rect 185 0 197 8242
rect 208 7102 220 19964
rect 208 0 220 7088
rect 231 5948 243 19940
rect 231 0 243 5934
rect 254 4794 266 19916
rect 254 0 266 4780
rect 277 3640 289 19892
rect 277 0 289 3626
rect 300 2486 312 19868
rect 300 0 312 2472
rect 323 1332 335 19844
rect 323 0 335 1318
rect 346 178 358 19820
rect 370 19812 570 20197
rect 586 19812 598 20197
rect 610 19812 622 20197
rect 634 19812 646 20197
rect 658 19812 670 20197
rect 4138 19812 4150 20197
rect 4162 19812 4174 20060
rect 4210 19812 4222 19988
rect 4378 19812 4390 20197
rect 4594 19812 4606 20036
rect 4642 19812 4654 19964
rect 4978 19812 4990 20012
rect 5026 19812 5038 19940
rect 5338 19812 5350 20197
rect 5530 19812 5542 20197
rect 6564 19812 6576 20197
rect 7118 19812 7130 19868
rect 7142 19812 7154 19892
rect 7166 19812 7178 19916
rect 14555 19812 14567 20197
rect 14579 19812 14591 20181
rect 14771 19812 14783 20156
rect 14819 19812 14831 20197
rect 14963 19812 14975 20132
rect 15155 19812 15167 20108
rect 15347 19812 15359 20084
rect 15539 19812 15551 20197
rect 17338 19812 17350 20197
rect 17530 19812 17542 20197
rect 17602 19812 17614 20197
rect 17698 19812 17710 20197
rect 22354 19812 22366 19892
rect 22546 19812 22558 19867
rect 22666 19812 22678 19844
rect 22786 19812 22798 19820
rect 25186 19812 25386 20197
rect 3082 18291 3094 18361
rect 3082 17137 3094 17207
rect 3082 15983 3094 16053
rect 3082 14829 3094 14899
rect 3082 13675 3094 13745
rect 3082 12521 3094 12591
rect 3082 11367 3094 11437
rect 3082 10213 3094 10283
rect 3082 9059 3094 9129
rect 3082 7905 3094 7975
rect 3082 6751 3094 6821
rect 3082 5597 3094 5667
rect 3082 4443 3094 4513
rect 3082 3289 3094 3359
rect 3082 2135 3094 2205
rect 3082 981 3094 1051
rect 346 0 358 164
rect 370 20 570 27
rect 370 6 556 20
rect 370 0 570 6
rect 586 0 598 27
rect 610 0 622 27
rect 634 0 646 27
rect 658 0 670 27
rect 1930 0 1942 27
rect 2122 0 2134 27
rect 2914 0 2926 27
rect 3322 19 3334 27
rect 3466 0 3478 27
rect 3682 0 3694 27
rect 4426 0 4438 27
rect 4594 0 4606 27
rect 4978 0 4990 27
rect 5170 0 5182 27
rect 5386 0 5398 27
rect 6130 0 6142 27
rect 6298 0 6310 27
rect 15706 0 15718 27
rect 15898 0 15910 27
rect 16138 0 16150 27
rect 16786 21 16798 27
rect 16978 21 16990 27
rect 16786 9 16990 21
rect 17266 19 17278 27
rect 19930 19 19942 27
rect 19978 19 19990 27
rect 20026 19 20038 27
rect 20074 19 20086 27
rect 20122 19 20134 27
rect 20170 19 20182 27
rect 20218 19 20230 27
rect 20266 19 20278 27
rect 20578 19 20590 27
rect 20626 19 20638 27
rect 20674 19 20686 27
rect 20722 19 20734 27
rect 21034 19 21046 27
rect 21082 19 21094 27
rect 21466 19 21478 27
rect 23842 0 23854 27
rect 24586 0 24598 27
rect 24730 0 24742 27
rect 24778 0 24790 27
rect 24826 0 24838 27
rect 24874 0 24886 27
rect 24946 0 24958 27
rect 25186 19 25386 27
rect 25200 5 25386 19
rect 25186 0 25386 5
use slice17 slice17_0
timestamp 1395569125
transform 1 0 370 0 1 18491
box 0 0 25016 1321
use leftbuf_slice leftbuf_slice_15
timestamp 1396382297
transform 1 0 365 0 1 17337
box 0 0 1685 1154
use IrAA IrAA_7
timestamp 1396382230
transform 1 0 2050 0 1 17337
box 0 0 1008 1154
use tielow tielow_0
timestamp 1386086605
transform 1 0 3058 0 1 17492
box 0 0 48 799
use leftbuf_slice leftbuf_slice_14
timestamp 1396382297
transform 1 0 365 0 1 16183
box 0 0 1685 1154
use IrAA IrAA_6
timestamp 1396382230
transform 1 0 2050 0 1 16183
box 0 0 1008 1154
use Datapath_slice Datapath_slice_15
timestamp 1396308628
transform 1 0 3106 0 1 17337
box 0 0 20472 1154
use LLIcell_U LLIcell_U_7
timestamp 1396314228
transform 1 0 23578 0 1 17337
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_11
timestamp 1396310136
transform 1 0 23770 0 1 17337
box 0 0 1621 1154
use tielow tielow_1
timestamp 1386086605
transform 1 0 3058 0 1 16338
box 0 0 48 799
use leftbuf_slice leftbuf_slice_13
timestamp 1396382297
transform 1 0 365 0 1 15029
box 0 0 1685 1154
use IrAA IrAA_5
timestamp 1396382230
transform 1 0 2050 0 1 15029
box 0 0 1008 1154
use Datapath_slice Datapath_slice_14
timestamp 1396308628
transform 1 0 3106 0 1 16183
box 0 0 20472 1154
use LLIcell_U LLIcell_U_6
timestamp 1396314228
transform 1 0 23578 0 1 16183
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_10
timestamp 1396310136
transform 1 0 23770 0 1 16183
box 0 0 1621 1154
use tielow tielow_2
timestamp 1386086605
transform 1 0 3058 0 1 15184
box 0 0 48 799
use leftbuf_slice leftbuf_slice_12
timestamp 1396382297
transform 1 0 365 0 1 13875
box 0 0 1685 1154
use IrAA IrAA_4
timestamp 1396382230
transform 1 0 2050 0 1 13875
box 0 0 1008 1154
use Datapath_slice Datapath_slice_13
timestamp 1396308628
transform 1 0 3106 0 1 15029
box 0 0 20472 1154
use LLIcell_U LLIcell_U_5
timestamp 1396314228
transform 1 0 23578 0 1 15029
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_9
timestamp 1396310136
transform 1 0 23770 0 1 15029
box 0 0 1621 1154
use tielow tielow_3
timestamp 1386086605
transform 1 0 3058 0 1 14030
box 0 0 48 799
use leftbuf_slice leftbuf_slice_11
timestamp 1396382297
transform 1 0 365 0 1 12721
box 0 0 1685 1154
use IrAA IrAA_3
timestamp 1396382230
transform 1 0 2050 0 1 12721
box 0 0 1008 1154
use Datapath_slice Datapath_slice_12
timestamp 1396308628
transform 1 0 3106 0 1 13875
box 0 0 20472 1154
use LLIcell_U LLIcell_U_4
timestamp 1396314228
transform 1 0 23578 0 1 13875
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_8
timestamp 1396310136
transform 1 0 23770 0 1 13875
box 0 0 1621 1154
use tielow tielow_4
timestamp 1386086605
transform 1 0 3058 0 1 12876
box 0 0 48 799
use leftbuf_slice leftbuf_slice_10
timestamp 1396382297
transform 1 0 365 0 1 11567
box 0 0 1685 1154
use IrAA IrAA_2
timestamp 1396382230
transform 1 0 2050 0 1 11567
box 0 0 1008 1154
use Datapath_slice Datapath_slice_11
timestamp 1396308628
transform 1 0 3106 0 1 12721
box 0 0 20472 1154
use LLIcell_U LLIcell_U_3
timestamp 1396314228
transform 1 0 23578 0 1 12721
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_7
timestamp 1396310136
transform 1 0 23770 0 1 12721
box 0 0 1621 1154
use tielow tielow_5
timestamp 1386086605
transform 1 0 3058 0 1 11722
box 0 0 48 799
use leftbuf_slice leftbuf_slice_9
timestamp 1396382297
transform 1 0 365 0 1 10413
box 0 0 1685 1154
use IrAA IrAA_1
timestamp 1396382230
transform 1 0 2050 0 1 10413
box 0 0 1008 1154
use Datapath_slice Datapath_slice_10
timestamp 1396308628
transform 1 0 3106 0 1 11567
box 0 0 20472 1154
use LLIcell_U LLIcell_U_2
timestamp 1396314228
transform 1 0 23578 0 1 11567
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_6
timestamp 1396310136
transform 1 0 23770 0 1 11567
box 0 0 1621 1154
use tielow tielow_6
timestamp 1386086605
transform 1 0 3058 0 1 10568
box 0 0 48 799
use leftbuf_slice leftbuf_slice_8
timestamp 1396382297
transform 1 0 365 0 1 9259
box 0 0 1685 1154
use IrAA IrAA_0
timestamp 1396382230
transform 1 0 2050 0 1 9259
box 0 0 1008 1154
use Datapath_slice Datapath_slice_9
timestamp 1396308628
transform 1 0 3106 0 1 10413
box 0 0 20472 1154
use LLIcell_U LLIcell_U_1
timestamp 1396314228
transform 1 0 23578 0 1 10413
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_5
timestamp 1396310136
transform 1 0 23770 0 1 10413
box 0 0 1621 1154
use tielow tielow_7
timestamp 1386086605
transform 1 0 3058 0 1 9414
box 0 0 48 799
use leftbuf_slice leftbuf_slice_7
timestamp 1396382297
transform 1 0 365 0 1 8105
box 0 0 1685 1154
use IrBA IrBA_2
timestamp 1396382245
transform 1 0 2050 0 1 8105
box 0 0 1008 1154
use Datapath_slice Datapath_slice_8
timestamp 1396308628
transform 1 0 3106 0 1 9259
box 0 0 20472 1154
use LLIcell_U LLIcell_U_0
timestamp 1396314228
transform 1 0 23578 0 1 9259
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_4
timestamp 1396310136
transform 1 0 23770 0 1 9259
box 0 0 1621 1154
use tielow tielow_8
timestamp 1386086605
transform 1 0 3058 0 1 8260
box 0 0 48 799
use leftbuf_slice leftbuf_slice_6
timestamp 1396382297
transform 1 0 365 0 1 6951
box 0 0 1685 1154
use IrBA IrBA_1
timestamp 1396382245
transform 1 0 2050 0 1 6951
box 0 0 1008 1154
use Datapath_slice Datapath_slice_7
timestamp 1396308628
transform 1 0 3106 0 1 8105
box 0 0 20472 1154
use LLIcell_L LLIcell_L_7
timestamp 1396313505
transform 1 0 23578 0 1 8105
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_3
timestamp 1396310136
transform 1 0 23770 0 1 8105
box 0 0 1621 1154
use tielow tielow_9
timestamp 1386086605
transform 1 0 3058 0 1 7106
box 0 0 48 799
use leftbuf_slice leftbuf_slice_5
timestamp 1396382297
transform 1 0 365 0 1 5797
box 0 0 1685 1154
use IrBA IrBA_0
timestamp 1396382245
transform 1 0 2050 0 1 5797
box 0 0 1008 1154
use Datapath_slice Datapath_slice_6
timestamp 1396308628
transform 1 0 3106 0 1 6951
box 0 0 20472 1154
use LLIcell_L LLIcell_L_6
timestamp 1396313505
transform 1 0 23578 0 1 6951
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_2
timestamp 1396310136
transform 1 0 23770 0 1 6951
box 0 0 1621 1154
use tielow tielow_10
timestamp 1386086605
transform 1 0 3058 0 1 5952
box 0 0 48 799
use leftbuf_slice leftbuf_slice_4
timestamp 1396382297
transform 1 0 365 0 1 4643
box 0 0 1685 1154
use IrBB IrBB_4
timestamp 1396382275
transform 1 0 2050 0 1 4643
box 0 0 1008 1154
use Datapath_slice Datapath_slice_5
timestamp 1396308628
transform 1 0 3106 0 1 5797
box 0 0 20472 1154
use LLIcell_L LLIcell_L_5
timestamp 1396313505
transform 1 0 23578 0 1 5797
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_1
timestamp 1396310136
transform 1 0 23770 0 1 5797
box 0 0 1621 1154
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 3058 0 1 4798
box 0 0 48 799
use leftbuf_slice leftbuf_slice_3
timestamp 1396382297
transform 1 0 365 0 1 3489
box 0 0 1685 1154
use IrBB IrBB_3
timestamp 1396382275
transform 1 0 2050 0 1 3489
box 0 0 1008 1154
use Datapath_slice Datapath_slice_4
timestamp 1396308628
transform 1 0 3106 0 1 4643
box 0 0 20472 1154
use LLIcell_L LLIcell_L_4
timestamp 1396313505
transform 1 0 23578 0 1 4643
box 0 0 192 1154
use Datapath_end_high Datapath_end_high_0
timestamp 1396310136
transform 1 0 23770 0 1 4643
box 0 0 1621 1154
use tielow tielow_12
timestamp 1386086605
transform 1 0 3058 0 1 3644
box 0 0 48 799
use leftbuf_slice leftbuf_slice_2
timestamp 1396382297
transform 1 0 365 0 1 2335
box 0 0 1685 1154
use IrBB IrBB_2
timestamp 1396382275
transform 1 0 2050 0 1 2335
box 0 0 1008 1154
use Datapath_slice Datapath_slice_3
timestamp 1396308628
transform 1 0 3106 0 1 3489
box 0 0 20472 1154
use LLIcell_L LLIcell_L_3
timestamp 1396313505
transform 1 0 23578 0 1 3489
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_3
timestamp 1396310181
transform 1 0 23770 0 1 3467
box 0 22 1621 1176
use tielow tielow_13
timestamp 1386086605
transform 1 0 3058 0 1 2490
box 0 0 48 799
use leftbuf_slice leftbuf_slice_1
timestamp 1396382297
transform 1 0 365 0 1 1181
box 0 0 1685 1154
use IrBB IrBB_1
timestamp 1396382275
transform 1 0 2050 0 1 1181
box 0 0 1008 1154
use Datapath_slice Datapath_slice_2
timestamp 1396308628
transform 1 0 3106 0 1 2335
box 0 0 20472 1154
use LLIcell_L LLIcell_L_2
timestamp 1396313505
transform 1 0 23578 0 1 2335
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_2
timestamp 1396310181
transform 1 0 23770 0 1 2313
box 0 22 1621 1176
use tielow tielow_14
timestamp 1386086605
transform 1 0 3058 0 1 1336
box 0 0 48 799
use leftbuf_slice leftbuf_slice_0
timestamp 1396382297
transform 1 0 365 0 1 27
box 0 0 1685 1154
use IrBB IrBB_0
timestamp 1396382275
transform 1 0 2050 0 1 27
box 0 0 1008 1154
use Datapath_slice Datapath_slice_1
timestamp 1396308628
transform 1 0 3106 0 1 1181
box 0 0 20472 1154
use LLIcell_L LLIcell_L_1
timestamp 1396313505
transform 1 0 23578 0 1 1181
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_1
timestamp 1396310181
transform 1 0 23770 0 1 1159
box 0 22 1621 1176
use tielow tielow_15
timestamp 1386086605
transform 1 0 3058 0 1 182
box 0 0 48 799
use Datapath_slice Datapath_slice_0
timestamp 1396308628
transform 1 0 3106 0 1 27
box 0 0 20472 1154
use LLIcell_L LLIcell_L_0
timestamp 1396313505
transform 1 0 23578 0 1 27
box 0 0 192 1154
use Datapath_end_low Datapath_end_low_0
timestamp 1396310181
transform 1 0 23770 0 1 5
box 0 22 1621 1176
<< labels >>
rlabel metal2 6 19885 6 19885 1 Ir[15]
rlabel metal2 30 19884 30 19884 1 Ir[14]
rlabel metal2 53 19884 53 19884 1 Ir[13]
rlabel metal2 76 19885 76 19885 1 Ir[12]
rlabel metal2 99 19885 99 19885 1 Ir[11]
rlabel metal2 122 19884 122 19884 1 Ir[10]
rlabel metal2 145 19885 145 19885 1 Ir[9]
rlabel metal2 168 19885 168 19885 1 Ir[8]
rlabel metal2 191 19887 191 19887 1 Ir[7]
rlabel metal2 214 19888 214 19888 1 Ir[6]
rlabel metal2 237 19889 237 19889 1 Ir[5]
rlabel metal2 260 19890 260 19890 1 Ir[4]
rlabel metal2 283 19889 283 19889 1 Ir[3]
rlabel metal2 22792 19815 22792 19815 1 Ir[0]
rlabel metal2 22671 19837 22671 19837 1 Ir[1]
rlabel metal2 22551 19862 22551 19862 1 Ir[2]
rlabel metal2 22360 19887 22360 19887 1 Ir[3]
rlabel metal2 14968 20126 14968 20126 1 Ir[13]
rlabel metal2 15161 20102 15161 20102 1 Ir[12]
rlabel metal2 15353 20077 15353 20077 1 Ir[11]
rlabel metal2 14775 20149 14775 20149 1 Ir[14]
rlabel metal2 14584 20174 14584 20174 1 Ir[15]
rlabel metal2 7122 19860 7122 19860 1 Ir[2]
rlabel metal2 7148 19884 7148 19884 1 Ir[3]
rlabel metal2 7171 19908 7171 19908 1 Ir[4]
rlabel metal2 4216 19980 4216 19980 1 Ir[7]
rlabel metal2 4167 20053 4167 20053 1 Ir[10]
rlabel metal2 4648 19957 4648 19957 1 Ir[6]
rlabel metal2 4599 20028 4599 20028 1 Ir[9]
rlabel metal2 4983 20005 4983 20005 1 Ir[8]
rlabel metal2 5033 19934 5033 19934 1 Ir[5]
rlabel metal2 6564 20197 6576 20197 5 RegWe
rlabel metal2 586 20197 598 20197 5 SDO
rlabel metal2 370 20197 570 20197 5 Vdd!
rlabel metal2 658 20197 670 20197 1 nReset
rlabel metal2 634 20197 646 20197 1 Clock
rlabel metal2 610 20197 622 20197 1 Test
rlabel metal2 17698 20197 17710 20197 5 Flags[0]
rlabel metal2 17602 20197 17614 20197 5 Flags[3]
rlabel metal2 17530 20197 17542 20197 5 Flags[1]
rlabel metal2 17338 20197 17350 20197 5 Flags[2]
rlabel metal2 14819 20197 14831 20197 5 AluOR[0]
rlabel metal2 14555 20197 14567 20197 5 AluOR[1]
rlabel metal2 15539 20197 15551 20197 5 CFlag
rlabel metal2 4138 20197 4150 20197 5 Rs1Sel[0]
rlabel metal2 4378 20197 4390 20197 5 Rs1Sel[1]
rlabel metal2 5338 20197 5350 20197 5 RwSel[0]
rlabel metal2 5530 20197 5542 20197 5 RwSel[1]
rlabel metal2 25186 20197 25386 20197 1 GND!
rlabel metal1 25408 1209 25408 1219 7 DataIn[1]
rlabel metal1 25408 1253 25408 1263 7 DataOut[1]
rlabel metal1 25408 2363 25408 2373 7 DataIn[2]
rlabel metal1 25408 2407 25408 2417 7 DataOut[2]
rlabel metal1 25408 3517 25408 3527 7 DataIn[3]
rlabel metal1 25408 3561 25408 3571 7 DataOut[3]
rlabel metal1 25408 4671 25408 4681 7 DataIn[4]
rlabel metal1 25408 4715 25408 4725 7 DataOut[4]
rlabel metal1 25408 5825 25408 5835 7 DataIn[5]
rlabel metal1 25408 5869 25408 5879 7 DataOut[5]
rlabel metal1 25408 6979 25408 6989 7 DataIn[6]
rlabel metal1 25408 7023 25408 7033 7 DataOut[6]
rlabel metal1 25408 8133 25408 8143 7 DataIn[7]
rlabel metal1 25408 8177 25408 8187 7 DataOut[7]
rlabel metal1 25408 9287 25408 9297 7 DataIn[8]
rlabel metal1 25408 9331 25408 9341 7 DataOut[8]
rlabel metal1 25408 10441 25408 10451 7 DataIn[9]
rlabel metal1 25408 10485 25408 10495 7 DataOut[9]
rlabel metal1 25408 11595 25408 11605 7 DataIn[10]
rlabel metal1 25408 11639 25408 11649 7 DataOut[10]
rlabel metal1 25408 12749 25408 12759 7 DataIn[11]
rlabel metal1 25408 12793 25408 12803 7 DataOut[11]
rlabel metal1 25408 13903 25408 13913 7 DataIn[12]
rlabel metal1 25408 13947 25408 13957 7 DataOut[12]
rlabel metal1 25408 15057 25408 15067 7 DataIn[13]
rlabel metal1 25408 15101 25408 15111 7 DataOut[13]
rlabel metal1 25408 16211 25408 16221 7 DataIn[14]
rlabel metal1 25408 16255 25408 16265 7 DataOut[14]
rlabel metal1 25408 17365 25408 17375 7 DataIn[15]
rlabel metal1 25408 17409 25408 17419 7 DataOut[15]
rlabel metal1 25408 99 25408 109 7 DataOut[0]
rlabel metal1 25408 55 25408 65 7 DataIn[0]
rlabel metal2 1 0 13 0 1 Ir[15]
rlabel metal2 24 0 36 0 1 Ir[14]
rlabel metal2 47 0 59 0 1 Ir[13]
rlabel metal2 70 0 82 0 1 Ir[12]
rlabel metal2 93 0 105 0 1 Ir[11]
rlabel metal2 116 0 128 0 1 Ir[10]
rlabel metal2 139 0 151 0 1 Ir[9]
rlabel metal2 162 0 174 0 1 Ir[8]
rlabel metal2 185 0 197 0 1 Ir[7]
rlabel metal2 208 0 220 0 1 Ir[6]
rlabel metal2 231 0 243 0 1 Ir[5]
rlabel metal2 254 0 266 0 1 Ir[4]
rlabel metal2 277 0 289 0 1 Ir[3]
rlabel metal2 300 0 312 0 1 Ir[2]
rlabel metal2 323 0 335 0 1 Ir[1]
rlabel metal2 346 0 358 0 1 Ir[0]
rlabel metal2 3466 0 3478 0 1 LrSel
rlabel metal2 3682 0 3694 0 1 LrWe
rlabel metal2 2914 0 2926 0 1 ImmSel
rlabel metal2 2122 0 2134 0 1 IrWe
rlabel metal2 1930 0 1942 0 1 MemEn
rlabel metal2 24874 0 24886 0 1 StatusReg[0]
rlabel metal2 24826 0 24838 0 1 StatusReg[1]
rlabel metal2 24778 0 24790 0 1 StatusReg[2]
rlabel metal2 24730 0 24742 0 1 StatusReg[3]
rlabel metal2 24946 0 24958 0 1 StatusRegEn
rlabel metal2 25186 0 25386 0 1 GND!
rlabel metal2 16138 0 16150 0 1 Op2Sel[1]
rlabel metal2 15898 0 15910 0 1 Op2Sel[0]
rlabel metal2 15706 0 15718 0 1 Op1Sel
rlabel metal2 6298 0 6310 0 1 WdSel
rlabel metal2 6130 0 6142 0 1 PcEn
rlabel metal2 5170 0 5182 0 1 PcSel[2]
rlabel metal2 5386 0 5398 0 1 PcWe
rlabel metal2 658 0 670 0 1 nReset
rlabel metal2 634 0 646 0 1 Clock
rlabel metal2 610 0 622 0 1 Test
rlabel metal2 586 0 598 0 1 SDI
rlabel metal2 370 0 570 0 1 Vdd!
rlabel metal2 24586 0 24598 0 1 AluEn
rlabel metal2 23842 0 23854 0 1 AluWe
rlabel metal2 4978 0 4990 0 1 PcSel[1]
rlabel metal2 4594 0 4606 0 1 PcSel[0]
rlabel metal2 4426 0 4438 0 1 LrEn
<< end >>
