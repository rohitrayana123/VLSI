magic
tech c035u
timestamp 1394559066
<< glass >>
rect 168 375 768 1174
rect 1680 375 2688 1174
rect 3840 375 4896 1174
rect 5136 375 5640 1174
rect 5760 375 6264 1174
rect 6480 375 6840 1174
rect 7128 375 7176 1174
<< metal1 >>
rect 3709 1442 4751 1452
rect 3589 1420 4655 1430
rect 3349 1398 4463 1408
rect 3109 1377 4271 1387
rect 2989 1355 4175 1365
rect 3829 1333 4079 1343
rect 4093 1333 4847 1343
rect 3469 1311 3983 1321
rect 3997 1311 4559 1321
rect 1933 1289 1967 1299
rect 2197 1289 2471 1299
rect 3229 1289 3887 1299
rect 3901 1289 4367 1299
rect 4597 1289 6407 1299
rect 685 1267 3071 1277
rect 3085 1267 3311 1277
rect 3325 1267 3551 1277
rect 3565 1267 3791 1277
rect 3805 1267 4967 1277
rect 4981 1267 5303 1277
rect 565 1245 3167 1255
rect 3181 1245 3287 1255
rect 3301 1245 3647 1255
rect 3661 1245 3767 1255
rect 3781 1245 4943 1255
rect 4957 1245 5183 1255
rect 5197 1245 5279 1255
rect 5293 1245 5927 1255
rect 5941 1245 6911 1255
rect 445 1223 1727 1233
rect 1741 1223 3383 1233
rect 3397 1223 3503 1233
rect 3517 1223 3623 1233
rect 3637 1223 3743 1233
rect 3757 1223 6887 1233
rect 7117 1223 7223 1233
rect 325 1201 2831 1211
rect 2845 1201 4919 1211
rect 5005 1201 5038 1211
rect 5365 1201 5423 1211
rect 5869 1201 6047 1211
rect 6109 1201 6143 1211
rect 6253 1201 6287 1211
rect 6301 1201 6503 1211
rect 6517 1201 6623 1211
rect 6637 1201 6743 1211
rect 6973 1201 7199 1211
rect 205 1179 1703 1189
rect 1717 1179 2711 1189
rect 2725 1179 2807 1189
rect 2821 1179 5063 1189
rect 5245 1179 5399 1189
rect 5485 1179 5519 1189
rect 5989 1179 6023 1189
rect 6037 1179 7247 1189
rect 7309 1179 7343 1189
rect 0 1096 168 1121
rect 7440 1096 7602 1121
rect 0 451 168 476
rect 7440 451 7602 476
rect 253 360 5543 370
rect 5557 360 6167 370
rect 6181 360 7367 370
rect 373 338 2735 348
rect 2749 338 5159 348
rect 5173 338 6191 348
rect 6205 338 6863 348
rect 6877 338 7007 348
rect 7165 338 7583 348
rect 493 316 1751 326
rect 1765 316 2903 326
rect 2917 316 3023 326
rect 3037 316 3143 326
rect 3157 316 3263 326
rect 3277 316 5567 326
rect 5581 316 5783 326
rect 5797 316 5903 326
rect 5917 316 7031 326
rect 7189 316 7415 326
rect 613 294 2927 304
rect 2941 294 3047 304
rect 3061 294 3407 304
rect 3421 294 3527 304
rect 3565 294 4103 304
rect 4165 294 4247 304
rect 4261 294 4343 304
rect 4357 294 4439 304
rect 4453 294 4535 304
rect 4549 294 4631 304
rect 4645 294 4727 304
rect 4741 294 4823 304
rect 5390 294 5615 304
rect 6349 294 6383 304
rect 733 272 2951 282
rect 2965 272 3191 282
rect 3205 272 3431 282
rect 3445 272 3671 282
rect 3685 272 5807 282
rect 5821 272 7055 282
rect 349 250 1991 260
rect 2005 250 2351 260
rect 2869 249 3863 259
rect 3877 249 3959 259
rect 3973 249 4055 259
rect 5365 250 6455 260
rect 1813 228 1871 238
rect 2773 227 4151 237
rect 4353 228 4487 238
rect 6013 228 6575 238
rect 85 205 3911 215
rect 4021 205 5687 215
rect 6469 206 6695 216
rect 517 183 2087 193
rect 2245 183 4339 193
rect 4693 183 7343 193
rect 685 161 2159 171
rect 2893 161 4775 171
rect 709 139 2375 149
rect 3229 139 4871 149
rect 781 117 2543 127
rect 3349 117 5663 127
rect 997 95 2591 105
rect 3397 95 4583 105
rect 1141 73 5111 83
rect 1477 51 4199 61
rect 1837 29 4295 39
rect 2581 7 4391 17
<< m2contact >>
rect 3695 1440 3709 1454
rect 4751 1440 4765 1454
rect 3575 1418 3589 1432
rect 4655 1418 4669 1432
rect 3335 1397 3349 1411
rect 4463 1396 4477 1410
rect 3095 1375 3109 1389
rect 4271 1374 4285 1388
rect 2975 1353 2989 1367
rect 4175 1353 4189 1367
rect 3815 1331 3829 1345
rect 4079 1331 4093 1345
rect 4847 1331 4861 1345
rect 3455 1309 3469 1323
rect 3983 1309 3997 1323
rect 4559 1309 4573 1323
rect 1919 1287 1933 1301
rect 1967 1287 1981 1301
rect 2183 1287 2197 1301
rect 2471 1287 2485 1301
rect 3215 1287 3229 1301
rect 3887 1287 3901 1301
rect 4367 1287 4381 1301
rect 4583 1287 4597 1301
rect 6407 1287 6421 1301
rect 671 1265 685 1279
rect 3071 1265 3085 1279
rect 3311 1265 3325 1279
rect 3551 1265 3565 1279
rect 3791 1265 3805 1279
rect 4967 1265 4981 1279
rect 5303 1265 5317 1279
rect 551 1243 565 1257
rect 3167 1243 3181 1257
rect 3287 1243 3301 1257
rect 3647 1243 3661 1257
rect 3767 1243 3781 1257
rect 4943 1243 4957 1257
rect 5183 1243 5197 1257
rect 5279 1243 5293 1257
rect 5927 1243 5941 1257
rect 6911 1243 6925 1257
rect 431 1221 445 1235
rect 1727 1221 1741 1235
rect 3383 1221 3397 1235
rect 3503 1221 3517 1235
rect 3623 1221 3637 1235
rect 3743 1221 3757 1235
rect 6887 1221 6901 1235
rect 7103 1221 7117 1235
rect 7223 1221 7237 1235
rect 311 1199 325 1213
rect 2831 1199 2845 1213
rect 4919 1199 4933 1213
rect 4991 1199 5005 1213
rect 5038 1199 5052 1213
rect 5351 1199 5365 1213
rect 5423 1199 5437 1213
rect 5855 1199 5869 1213
rect 6047 1199 6061 1213
rect 6095 1199 6109 1213
rect 6143 1199 6157 1213
rect 6239 1199 6253 1213
rect 6287 1199 6301 1213
rect 6503 1199 6517 1213
rect 6623 1199 6637 1213
rect 6743 1199 6757 1213
rect 6959 1199 6973 1213
rect 7199 1199 7213 1213
rect 191 1177 205 1191
rect 1703 1177 1717 1191
rect 2711 1177 2725 1191
rect 2807 1177 2821 1191
rect 5063 1177 5077 1191
rect 5231 1177 5245 1191
rect 5399 1177 5413 1191
rect 5471 1177 5485 1191
rect 5519 1177 5533 1191
rect 5975 1177 5989 1191
rect 6023 1177 6037 1191
rect 7247 1177 7261 1191
rect 7295 1177 7309 1191
rect 7343 1177 7357 1191
rect 239 358 253 372
rect 5543 358 5557 372
rect 6167 358 6181 372
rect 7367 358 7381 372
rect 359 336 373 350
rect 2735 336 2749 350
rect 5159 336 5173 350
rect 6191 336 6205 350
rect 6863 336 6877 350
rect 7007 336 7021 350
rect 7151 336 7165 350
rect 7583 336 7597 350
rect 479 314 493 328
rect 1751 314 1765 328
rect 2903 314 2917 328
rect 3023 314 3037 328
rect 3143 314 3157 328
rect 3263 314 3277 328
rect 5567 314 5581 328
rect 5783 314 5797 328
rect 5903 314 5917 328
rect 7031 314 7045 328
rect 7175 314 7189 328
rect 7415 314 7429 328
rect 599 292 613 306
rect 2927 292 2941 306
rect 3047 292 3061 306
rect 3407 292 3421 306
rect 3527 292 3541 306
rect 3551 292 3565 306
rect 4103 292 4117 306
rect 4151 292 4165 306
rect 4247 292 4261 306
rect 4343 292 4357 306
rect 4439 292 4453 306
rect 4535 292 4549 306
rect 4631 292 4645 306
rect 4727 292 4741 306
rect 4823 292 4837 306
rect 5376 292 5390 306
rect 5615 292 5629 306
rect 6335 292 6349 306
rect 6383 292 6397 306
rect 719 270 733 284
rect 2951 270 2965 284
rect 3191 270 3205 284
rect 3431 270 3445 284
rect 3671 270 3685 284
rect 5807 270 5821 284
rect 7055 269 7069 283
rect 335 248 349 262
rect 1991 248 2005 262
rect 2351 248 2365 262
rect 2855 247 2869 261
rect 3863 247 3877 261
rect 3959 247 3973 261
rect 4055 247 4069 261
rect 5351 248 5365 262
rect 6455 248 6469 262
rect 1799 226 1813 240
rect 1871 226 1885 240
rect 2759 225 2773 239
rect 4151 225 4165 239
rect 4339 226 4353 240
rect 4487 226 4501 240
rect 5999 226 6013 240
rect 6575 226 6589 240
rect 71 203 85 217
rect 3911 203 3925 217
rect 4007 203 4021 217
rect 5687 203 5701 217
rect 6455 204 6469 218
rect 6695 204 6709 218
rect 503 181 517 195
rect 2087 181 2101 195
rect 2231 181 2245 195
rect 4339 181 4353 195
rect 4679 181 4693 195
rect 7343 181 7357 195
rect 671 159 685 173
rect 2159 159 2173 173
rect 2879 159 2893 173
rect 4775 159 4789 173
rect 695 137 709 151
rect 2375 137 2389 151
rect 3215 137 3229 151
rect 4871 137 4885 151
rect 767 115 781 129
rect 2543 115 2557 129
rect 3335 115 3349 129
rect 5663 115 5677 129
rect 983 93 997 107
rect 2591 93 2605 107
rect 3383 93 3397 107
rect 4583 93 4597 107
rect 1127 71 1141 85
rect 5111 71 5125 85
rect 1463 49 1477 63
rect 4199 49 4213 63
rect 1823 27 1837 41
rect 4295 27 4309 41
rect 2567 5 2581 19
rect 4391 5 4405 19
<< metal2 >>
rect 192 1191 204 1659
rect 312 1213 324 1659
rect 432 1235 444 1659
rect 552 1257 564 1659
rect 672 1279 684 1659
rect 192 1174 204 1177
rect 312 1174 324 1199
rect 432 1174 444 1221
rect 552 1174 564 1243
rect 672 1174 684 1265
rect 1704 1174 1716 1177
rect 1728 1174 1740 1221
rect 1848 1174 1860 1659
rect 1920 1174 1932 1287
rect 1968 1174 1980 1287
rect 2184 1174 2196 1287
rect 2280 1174 2292 1659
rect 2472 1301 2484 1659
rect 2472 1174 2484 1287
rect 2544 1174 2556 1659
rect 2640 1174 2652 1659
rect 2712 1174 2724 1177
rect 2808 1174 2820 1177
rect 2832 1174 2844 1199
rect 2976 1174 2988 1353
rect 3072 1174 3084 1265
rect 3096 1174 3108 1375
rect 3168 1174 3180 1243
rect 3216 1174 3228 1287
rect 3288 1174 3300 1243
rect 3312 1174 3324 1265
rect 3336 1174 3348 1397
rect 3384 1174 3396 1221
rect 3456 1174 3468 1309
rect 3504 1174 3516 1221
rect 3552 1174 3564 1265
rect 3576 1174 3588 1418
rect 3624 1174 3636 1221
rect 3648 1174 3660 1243
rect 3696 1174 3708 1440
rect 3744 1174 3756 1221
rect 3768 1174 3780 1243
rect 3792 1174 3804 1265
rect 3816 1174 3828 1331
rect 3888 1174 3900 1287
rect 3984 1174 3996 1309
rect 4080 1174 4092 1331
rect 4176 1174 4188 1353
rect 4272 1174 4284 1374
rect 4368 1174 4380 1287
rect 4464 1174 4476 1396
rect 4560 1174 4572 1309
rect 4584 1174 4596 1287
rect 4656 1174 4668 1418
rect 4752 1174 4764 1440
rect 4848 1174 4860 1331
rect 4920 1174 4932 1199
rect 4944 1174 4956 1243
rect 4968 1174 4980 1265
rect 4992 1174 5004 1199
rect 5040 1174 5052 1199
rect 5064 1174 5076 1177
rect 5184 1174 5196 1243
rect 5232 1174 5244 1177
rect 5280 1174 5292 1243
rect 5304 1174 5316 1265
rect 5352 1174 5364 1199
rect 5400 1174 5412 1177
rect 5424 1174 5436 1199
rect 5472 1174 5484 1177
rect 5520 1174 5532 1177
rect 5856 1174 5868 1199
rect 5928 1174 5940 1243
rect 5976 1174 5988 1177
rect 6024 1174 6036 1177
rect 6048 1174 6060 1199
rect 6096 1174 6108 1199
rect 6144 1174 6156 1199
rect 6240 1174 6252 1199
rect 6288 1174 6300 1199
rect 6312 1174 6324 1659
rect 6408 1174 6420 1287
rect 6504 1174 6516 1199
rect 6528 1174 6540 1659
rect 6624 1174 6636 1199
rect 6648 1174 6660 1659
rect 6744 1174 6756 1199
rect 6768 1174 6780 1659
rect 6888 1174 6900 1221
rect 6912 1174 6924 1243
rect 6960 1174 6972 1199
rect 7104 1174 7116 1221
rect 7152 1174 7164 1659
rect 7200 1174 7212 1199
rect 7224 1174 7236 1221
rect 7248 1174 7260 1177
rect 7296 1174 7308 1177
rect 7344 1174 7356 1177
rect 240 372 252 375
rect 360 350 372 375
rect 480 328 492 375
rect 600 306 612 375
rect 720 284 732 375
rect 1752 328 1764 375
rect 72 -200 84 203
rect 336 -200 348 248
rect 1800 240 1812 375
rect 1872 240 1884 375
rect 1992 262 2004 375
rect 2088 195 2100 375
rect 504 -200 516 181
rect 2160 173 2172 375
rect 2352 262 2364 375
rect 672 -200 684 159
rect 696 -200 708 137
rect 768 -200 780 115
rect 984 -200 996 93
rect 1128 -200 1140 71
rect 1464 -200 1476 49
rect 1824 -200 1836 27
rect 2232 -200 2244 181
rect 2376 151 2388 375
rect 2544 129 2556 375
rect 2592 107 2604 375
rect 2736 350 2748 375
rect 2760 239 2772 375
rect 2856 261 2868 375
rect 2904 328 2916 375
rect 2928 306 2940 375
rect 2952 284 2964 375
rect 3024 328 3036 375
rect 3048 306 3060 375
rect 3144 328 3156 375
rect 3192 284 3204 375
rect 3264 328 3276 375
rect 3408 306 3420 375
rect 3432 284 3444 375
rect 3528 306 3540 375
rect 2568 -200 2580 5
rect 2880 -200 2892 159
rect 3216 -200 3228 137
rect 3336 -200 3348 115
rect 3384 -200 3396 93
rect 3552 -200 3564 292
rect 3672 284 3684 375
rect 3864 261 3876 375
rect 3912 217 3924 375
rect 3960 261 3972 375
rect 4008 217 4020 375
rect 4056 261 4068 375
rect 4104 306 4116 375
rect 4152 306 4164 375
rect 4152 239 4164 292
rect 4200 63 4212 375
rect 4248 306 4260 375
rect 4296 41 4308 375
rect 4344 306 4356 375
rect 4340 195 4352 226
rect 4392 19 4404 375
rect 4440 306 4452 375
rect 4488 240 4500 375
rect 4536 306 4548 375
rect 4584 107 4596 375
rect 4632 306 4644 375
rect 4680 195 4692 375
rect 4728 306 4740 375
rect 4776 173 4788 375
rect 4824 306 4836 375
rect 4872 151 4884 375
rect 5112 85 5124 375
rect 5160 350 5172 375
rect 5544 372 5556 375
rect 5568 328 5580 375
rect 5616 306 5628 375
rect 5352 -200 5364 248
rect 5377 -200 5389 292
rect 5664 129 5676 375
rect 5688 217 5700 375
rect 5736 -200 5748 375
rect 5784 328 5796 375
rect 5808 284 5820 375
rect 5904 328 5916 375
rect 6168 372 6180 375
rect 6192 350 6204 375
rect 6336 306 6348 375
rect 6384 306 6396 375
rect 6456 262 6468 375
rect 6576 240 6588 375
rect 6000 -200 6012 226
rect 6696 218 6708 375
rect 6456 -200 6468 204
rect 6816 -200 6828 375
rect 6864 350 6876 375
rect 7008 350 7020 375
rect 7032 328 7044 375
rect 7056 283 7068 375
rect 7152 350 7164 375
rect 7368 372 7380 375
rect 7416 328 7428 375
rect 7176 -200 7188 314
rect 7344 -200 7356 181
rect 7584 -200 7596 336
use inv inv_0
timestamp 1386238110
transform 1 0 168 0 1 375
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 288 0 1 375
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 408 0 1 375
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 528 0 1 375
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 648 0 1 375
box 0 0 120 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 1680 0 1 375
box 0 0 144 799
use and2 and2_4
timestamp 1386234845
transform 1 0 1824 0 1 375
box 0 0 120 799
use xor2 xor2_3
timestamp 1386237344
transform 1 0 1944 0 1 375
box 0 0 192 799
use xor2 xor2_4
timestamp 1386237344
transform 1 0 2136 0 1 375
box 0 0 192 799
use xor2 xor2_5
timestamp 1386237344
transform 1 0 2328 0 1 375
box 0 0 192 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 2520 0 1 375
box 0 0 48 799
use inv inv_6
timestamp 1386238110
transform 1 0 2568 0 1 375
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 2688 0 1 375
box 0 0 96 799
use nand2 nand2_3
timestamp 1386234792
transform 1 0 2784 0 1 375
box 0 0 96 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 2880 0 1 375
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 3000 0 1 375
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 3120 0 1 375
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 3240 0 1 375
box 0 0 120 799
use nand3 nand3_8
timestamp 1386234893
transform 1 0 3360 0 1 375
box 0 0 120 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 3480 0 1 375
box 0 0 120 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 3600 0 1 375
box 0 0 120 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 3720 0 1 375
box 0 0 120 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 3840 0 1 375
box 0 0 96 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 3936 0 1 375
box 0 0 96 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 4032 0 1 375
box 0 0 96 799
use nand2 nand2_7
timestamp 1386234792
transform 1 0 4128 0 1 375
box 0 0 96 799
use nand2 nand2_8
timestamp 1386234792
transform 1 0 4224 0 1 375
box 0 0 96 799
use nand2 nand2_9
timestamp 1386234792
transform 1 0 4320 0 1 375
box 0 0 96 799
use nand2 nand2_10
timestamp 1386234792
transform 1 0 4416 0 1 375
box 0 0 96 799
use nand2 nand2_11
timestamp 1386234792
transform 1 0 4512 0 1 375
box 0 0 96 799
use nand2 nand2_12
timestamp 1386234792
transform 1 0 4608 0 1 375
box 0 0 96 799
use nand2 nand2_13
timestamp 1386234792
transform 1 0 4704 0 1 375
box 0 0 96 799
use nand2 nand2_14
timestamp 1386234792
transform 1 0 4800 0 1 375
box 0 0 96 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 4896 0 1 375
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 5016 0 1 375
box 0 0 120 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 5136 0 1 375
box 0 0 120 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 5256 0 1 375
box 0 0 120 799
use nor2 nor2_6
timestamp 1386235306
transform 1 0 5376 0 1 375
box 0 0 120 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 5496 0 1 375
box 0 0 144 799
use and2 and2_3
timestamp 1386234845
transform 1 0 5640 0 1 375
box 0 0 120 799
use nor2 nor2_7
timestamp 1386235306
transform 1 0 5760 0 1 375
box 0 0 120 799
use nor2 nor2_8
timestamp 1386235306
transform 1 0 5880 0 1 375
box 0 0 120 799
use nor2 nor2_9
timestamp 1386235306
transform 1 0 6000 0 1 375
box 0 0 120 799
use nor3 nor3_2
timestamp 1386235396
transform 1 0 6120 0 1 375
box 0 0 144 799
use nand2 nand2_15
timestamp 1386234792
transform 1 0 6264 0 1 375
box 0 0 96 799
use nor2 nor2_10
timestamp 1386235306
transform 1 0 6360 0 1 375
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 6480 0 1 375
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 6600 0 1 375
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 6720 0 1 375
box 0 0 120 799
use nor3 nor3_3
timestamp 1386235396
transform 1 0 6840 0 1 375
box 0 0 144 799
use nor3 nor3_4
timestamp 1386235396
transform 1 0 6984 0 1 375
box 0 0 144 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 7128 0 1 375
box 0 0 48 799
use nor3 nor3_5
timestamp 1386235396
transform 1 0 7176 0 1 375
box 0 0 144 799
use nor2 nor2_11
timestamp 1386235306
transform 1 0 7320 0 1 375
box 0 0 120 799
<< labels >>
rlabel metal1 504 322 504 322 1 nC
rlabel metal1 747 275 747 275 1 nE
rlabel metal1 272 364 272 364 1 nA
rlabel metal1 378 342 378 342 1 nB
rlabel metal1 627 297 627 297 1 nD
rlabel metal2 6245 1176 6245 1176 1 N
rlabel metal1 5502 209 5502 209 1 ShSign
rlabel metal1 0 1096 0 1121 3 Vdd!
rlabel metal1 0 451 0 476 3 GND!
rlabel metal1 7602 1096 7602 1121 7 Vdd!
rlabel metal1 7602 451 7602 476 7 GND!
rlabel metal1 1837 232 1837 232 1 UseC
rlabel metal2 5736 -200 5748 -200 1 ShInBit
rlabel metal2 2880 -200 2892 -200 1 NAND
rlabel metal2 336 -200 348 -200 1 SUB
rlabel metal2 504 -200 516 -200 1 CIn_slice
rlabel metal2 672 -200 684 -200 1 LastCIn
rlabel metal2 696 -200 708 -200 1 COut
rlabel metal2 984 -200 996 -200 1 nZ
rlabel metal2 1128 -200 1140 -200 1 FAOut
rlabel metal2 1464 -200 1476 -200 1 AND
rlabel metal2 1824 -200 1836 -200 1 OR
rlabel metal2 2232 -200 2244 -200 1 XOR
rlabel metal2 2568 -200 2580 -200 1 NOT
rlabel metal2 3552 -200 3564 -200 1 ShL
rlabel metal2 3336 -200 3348 -200 1 ASign
rlabel metal2 3384 -200 3396 -200 1 ShB
rlabel metal2 3216 -200 3228 -200 1 NOR
rlabel metal2 768 -200 780 -200 1 N
rlabel metal2 72 -200 84 -200 1 ZeroA
rlabel metal2 5352 -200 5364 -200 1 Sh8
rlabel metal2 6000 -200 6012 -200 1 Sh4
rlabel metal2 6816 -200 6828 -200 1 Sh1
rlabel metal2 5377 -200 5389 -200 1 ShR
rlabel metal2 6456 -200 6468 -200 1 Sh2
rlabel metal2 7176 -200 7188 -200 1 ShOut
rlabel metal2 7344 -200 7356 -200 1 LLI
rlabel metal2 7584 -200 7596 -200 1 OutEn
rlabel metal2 192 1659 204 1659 5 OpCode[4]
rlabel metal2 312 1659 324 1659 5 OpCode[3]
rlabel metal2 432 1659 444 1659 5 OpCode[2]
rlabel metal2 552 1659 564 1659 5 OpCode[1]
rlabel metal2 672 1659 684 1659 5 OpCode[0]
rlabel metal2 2640 1659 2652 1659 5 Z
rlabel metal2 2544 1659 2556 1659 5 N
rlabel metal2 2280 1659 2292 1659 5 V
rlabel metal2 1848 1659 1860 1659 5 Cin
rlabel metal2 2472 1659 2484 1659 5 C
rlabel metal2 6768 1659 6780 1659 5 imm4[0]
rlabel metal2 6648 1659 6660 1659 5 imm4[1]
rlabel metal2 6528 1659 6540 1659 5 imm4[2]
rlabel metal2 6312 1659 6324 1659 5 imm4[3]
rlabel metal2 7152 1659 7164 1659 5 OutEn
<< end >>
