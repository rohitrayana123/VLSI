magic
tech c035u
timestamp 1393852311
<< metal1 >>
rect 4285 1025 5807 1035
rect 3877 1003 5399 1013
rect 3421 981 4943 991
rect 4982 980 5375 990
rect 5389 980 5783 990
rect 5797 981 6143 991
rect 3397 958 3839 968
rect 3853 958 4247 968
rect 4261 958 4607 968
rect 4645 959 6167 969
rect 61 936 196 946
rect 277 936 479 946
rect 541 938 671 948
rect 3469 936 3671 946
rect 3925 936 4079 946
rect 4333 936 4439 946
rect 5005 936 5207 946
rect 5461 936 5615 946
rect 5869 937 5975 947
rect 6229 936 6287 946
rect 109 914 406 924
rect 517 914 527 924
rect 613 913 743 923
rect 757 914 887 924
rect 1189 914 1223 924
rect 1525 914 1583 924
rect 1933 914 1991 924
rect 2269 914 2327 924
rect 2605 914 2639 924
rect 2941 914 2975 924
rect 3517 914 3527 924
rect 3565 914 3575 924
rect 3613 914 3623 924
rect 3973 914 3983 924
rect 4021 914 4031 924
rect 4381 914 4391 924
rect 4693 917 4751 927
rect 4933 914 4967 924
rect 5029 914 5039 924
rect 5077 914 5087 924
rect 5125 914 5135 924
rect 5173 914 5279 924
rect 5485 914 5495 924
rect 5533 914 5543 924
rect 5581 914 5687 924
rect 5893 915 5903 925
rect 5941 914 6047 924
rect 6253 914 6359 924
rect 0 892 143 902
rect 157 892 1127 902
rect 1141 892 1463 902
rect 1477 892 1823 902
rect 1837 892 2567 902
rect 2581 892 2879 902
rect 2893 892 3287 902
rect 3301 892 6648 902
rect 0 870 23 880
rect 37 870 1103 880
rect 1117 870 1439 880
rect 1453 870 1799 880
rect 1813 870 2207 880
rect 2221 870 2543 880
rect 2557 870 2855 880
rect 2869 870 3167 880
rect 3181 870 3239 880
rect 3325 870 3479 880
rect 3493 870 3695 880
rect 3781 870 3935 880
rect 3949 870 4103 880
rect 4189 870 4343 880
rect 4357 870 4463 880
rect 4549 870 4775 880
rect 4861 870 5231 880
rect 5317 870 5639 880
rect 5726 870 5999 880
rect 6085 870 6311 880
rect 6397 870 6455 880
rect 61 51 196 61
rect 781 51 815 61
rect 1045 51 1367 61
rect 1381 51 1727 61
rect 1741 51 2135 61
rect 2149 51 2471 61
rect 2485 51 2783 61
rect 2797 51 3119 61
rect 3133 51 6599 61
rect 6613 51 6648 61
rect 3493 29 3503 39
rect 3541 29 3551 39
rect 3589 29 3599 39
rect 3637 29 3743 39
rect 3949 29 3959 39
rect 3997 29 4007 39
rect 4045 29 4151 39
rect 4357 29 4367 39
rect 4405 29 4511 39
rect 4789 29 4823 39
rect 4933 29 4968 39
rect 5053 29 5063 39
rect 5101 29 5111 39
rect 5149 29 5159 39
rect 5509 29 5519 39
rect 5557 29 5567 39
rect 5917 29 5927 39
rect 6253 29 6311 39
rect 5029 7 5231 17
rect 5485 7 5639 17
rect 5893 7 5999 17
<< m2contact >>
rect 4271 1023 4285 1037
rect 5807 1023 5821 1037
rect 3863 1001 3877 1015
rect 5399 1001 5413 1015
rect 3407 978 3421 992
rect 4943 979 4957 993
rect 4968 979 4982 993
rect 5375 979 5389 993
rect 5783 979 5797 993
rect 6143 979 6157 993
rect 3383 956 3397 970
rect 3839 956 3853 970
rect 4247 956 4261 970
rect 4607 956 4621 970
rect 4631 956 4645 970
rect 6167 957 6181 971
rect 47 934 61 948
rect 196 934 210 948
rect 263 935 277 949
rect 479 934 493 948
rect 527 936 541 950
rect 671 936 685 950
rect 3455 934 3469 948
rect 3671 934 3685 948
rect 3911 934 3925 948
rect 4079 934 4093 948
rect 4319 934 4333 948
rect 4439 934 4453 948
rect 4991 934 5005 948
rect 5207 934 5221 948
rect 5447 934 5461 948
rect 5615 934 5629 948
rect 5855 935 5869 949
rect 5975 935 5989 949
rect 6215 934 6229 948
rect 6287 934 6301 948
rect 95 912 109 926
rect 406 912 420 926
rect 503 912 517 926
rect 527 912 541 926
rect 599 912 613 926
rect 743 912 757 926
rect 887 912 901 926
rect 1175 912 1189 926
rect 1223 912 1237 926
rect 1511 912 1525 926
rect 1583 912 1597 926
rect 1919 912 1933 926
rect 1991 912 2005 926
rect 2255 912 2269 926
rect 2327 912 2341 926
rect 2591 912 2605 926
rect 2639 912 2653 926
rect 2927 912 2941 926
rect 2975 912 2989 926
rect 3503 912 3517 926
rect 3527 912 3541 926
rect 3551 912 3565 926
rect 3575 912 3589 926
rect 3599 912 3613 926
rect 3623 912 3637 926
rect 3959 912 3973 926
rect 3983 912 3997 926
rect 4007 912 4021 926
rect 4031 912 4045 926
rect 4367 912 4381 926
rect 4391 912 4405 926
rect 4679 916 4693 930
rect 4751 916 4765 930
rect 4919 912 4933 926
rect 4967 912 4981 926
rect 5015 912 5029 926
rect 5039 912 5053 926
rect 5063 912 5077 926
rect 5087 912 5101 926
rect 5111 912 5125 926
rect 5135 912 5149 926
rect 5159 912 5173 926
rect 5279 912 5293 926
rect 5471 912 5485 926
rect 5495 912 5509 926
rect 5519 912 5533 926
rect 5543 912 5557 926
rect 5567 912 5581 926
rect 5687 912 5701 926
rect 5879 913 5893 927
rect 5903 913 5917 927
rect 5927 913 5941 927
rect 6047 912 6061 926
rect 6239 912 6253 926
rect 6359 912 6373 926
rect 143 890 157 904
rect 1127 890 1141 904
rect 1463 890 1477 904
rect 1823 890 1837 904
rect 2567 890 2581 904
rect 2879 890 2893 904
rect 3287 890 3301 904
rect 23 868 37 882
rect 1103 868 1117 882
rect 1439 868 1453 882
rect 1799 868 1813 882
rect 2207 868 2221 882
rect 2543 868 2557 882
rect 2855 868 2869 882
rect 3167 868 3181 882
rect 3239 868 3253 882
rect 3311 868 3325 882
rect 3479 868 3493 882
rect 3695 868 3709 882
rect 3767 868 3781 882
rect 3935 868 3949 882
rect 4103 868 4117 882
rect 4175 868 4189 882
rect 4343 868 4357 882
rect 4463 868 4477 882
rect 4535 868 4549 882
rect 4775 868 4789 882
rect 4847 868 4861 882
rect 5231 868 5245 882
rect 5303 868 5317 882
rect 5639 868 5653 882
rect 5712 868 5726 882
rect 5999 868 6013 882
rect 6071 868 6085 882
rect 6311 868 6325 882
rect 6383 868 6397 882
rect 6455 868 6469 882
rect 47 49 61 63
rect 196 49 210 63
rect 767 49 781 63
rect 815 49 829 63
rect 1031 49 1045 63
rect 1367 49 1381 63
rect 1727 49 1741 63
rect 2135 49 2149 63
rect 2471 49 2485 63
rect 2783 49 2797 63
rect 3119 49 3133 63
rect 6599 49 6613 63
rect 3479 27 3493 41
rect 3503 27 3517 41
rect 3527 27 3541 41
rect 3551 27 3565 41
rect 3575 27 3589 41
rect 3599 27 3613 41
rect 3623 27 3637 41
rect 3743 27 3757 41
rect 3935 27 3949 41
rect 3959 27 3973 41
rect 3983 27 3997 41
rect 4007 27 4021 41
rect 4031 27 4045 41
rect 4151 27 4165 41
rect 4343 27 4357 41
rect 4367 27 4381 41
rect 4391 27 4405 41
rect 4511 27 4525 41
rect 4775 27 4789 41
rect 4823 27 4837 41
rect 4919 27 4933 41
rect 4968 27 4982 41
rect 5039 27 5053 41
rect 5063 27 5077 41
rect 5087 27 5101 41
rect 5111 27 5125 41
rect 5135 27 5149 41
rect 5159 27 5173 41
rect 5495 27 5509 41
rect 5519 27 5533 41
rect 5543 27 5557 41
rect 5567 27 5581 41
rect 5903 27 5917 41
rect 5927 27 5941 41
rect 6239 27 6253 41
rect 6311 27 6325 41
rect 5015 5 5029 19
rect 5231 5 5245 19
rect 5471 5 5485 19
rect 5639 5 5653 19
rect 5879 5 5893 19
rect 5999 5 6013 19
<< metal2 >>
rect 24 865 36 868
rect 48 865 60 934
rect 96 865 108 912
rect 144 865 156 890
rect 168 865 180 1042
rect 197 948 209 1042
rect 264 865 276 935
rect 336 865 348 1042
rect 408 865 420 912
rect 480 865 492 934
rect 504 926 516 1042
rect 528 950 540 1042
rect 600 926 612 1042
rect 528 865 540 912
rect 600 865 612 912
rect 672 865 684 936
rect 744 865 756 912
rect 816 865 828 1042
rect 888 865 900 912
rect 960 865 972 1042
rect 1104 865 1116 868
rect 1128 865 1140 890
rect 1176 865 1188 912
rect 1224 865 1236 912
rect 1296 865 1308 1042
rect 1440 865 1452 868
rect 1464 865 1476 890
rect 1512 865 1524 912
rect 1584 865 1596 912
rect 1656 865 1668 1042
rect 1800 865 1812 868
rect 1824 865 1836 890
rect 1920 865 1932 912
rect 1992 865 2004 912
rect 2064 865 2076 1042
rect 2208 865 2220 868
rect 2256 865 2268 912
rect 2328 865 2340 912
rect 2400 865 2412 1042
rect 2544 865 2556 868
rect 2568 865 2580 890
rect 2592 865 2604 912
rect 2640 865 2652 912
rect 2712 865 2724 1042
rect 2856 865 2868 868
rect 2880 865 2892 890
rect 2928 865 2940 912
rect 2976 865 2988 912
rect 3048 865 3060 1042
rect 3168 882 3180 1042
rect 3216 865 3228 1042
rect 3384 970 3396 1042
rect 3240 865 3252 868
rect 3288 865 3300 890
rect 3312 865 3324 868
rect 3384 865 3396 956
rect 3408 865 3420 978
rect 3456 865 3468 934
rect 3480 882 3492 1042
rect 3528 926 3540 1042
rect 3576 926 3588 1042
rect 3624 926 3636 1042
rect 3504 865 3516 912
rect 3552 865 3564 912
rect 3600 865 3612 912
rect 3672 865 3684 934
rect 3696 865 3708 868
rect 3768 865 3780 868
rect 3840 865 3852 956
rect 3864 865 3876 1001
rect 3912 865 3924 934
rect 3936 882 3948 1042
rect 3984 926 3996 1042
rect 4032 926 4044 1042
rect 3960 865 3972 912
rect 4008 865 4020 912
rect 4080 865 4092 934
rect 4104 865 4116 868
rect 4176 865 4188 868
rect 4248 865 4260 956
rect 4272 865 4284 1023
rect 4320 865 4332 934
rect 4344 882 4356 1042
rect 4392 926 4404 1042
rect 4368 865 4380 912
rect 4440 865 4452 934
rect 4464 865 4476 868
rect 4536 865 4548 868
rect 4608 865 4620 956
rect 4632 865 4644 956
rect 4680 865 4692 916
rect 4752 865 4764 916
rect 4776 882 4788 1042
rect 4944 993 4956 1042
rect 4969 993 4981 1042
rect 4776 865 4788 868
rect 4848 865 4860 868
rect 4920 865 4932 912
rect 4944 865 4956 979
rect 4969 926 4981 979
rect 4992 865 5004 934
rect 5016 926 5028 1042
rect 5064 926 5076 1042
rect 5112 926 5124 1042
rect 5160 926 5172 1042
rect 5400 1015 5412 1042
rect 5040 865 5052 912
rect 5088 865 5100 912
rect 5136 865 5148 912
rect 5208 865 5220 934
rect 5232 865 5244 868
rect 5280 865 5292 912
rect 5304 865 5316 868
rect 5376 865 5388 979
rect 5400 865 5412 1001
rect 5448 865 5460 934
rect 5472 926 5484 1042
rect 5520 926 5532 1042
rect 5568 926 5580 1042
rect 5808 1037 5820 1042
rect 5496 865 5508 912
rect 5544 865 5556 912
rect 5616 865 5628 934
rect 5640 865 5652 868
rect 5688 865 5700 912
rect 5712 865 5724 868
rect 5784 865 5796 979
rect 5808 865 5820 1023
rect 5856 865 5868 935
rect 5880 927 5892 1042
rect 5928 927 5940 1042
rect 5904 865 5916 913
rect 5976 865 5988 935
rect 6000 865 6012 868
rect 6048 865 6060 912
rect 6072 865 6084 868
rect 6144 865 6156 979
rect 6168 971 6180 1042
rect 6168 865 6180 957
rect 6216 865 6228 934
rect 6240 926 6252 1042
rect 6288 865 6300 934
rect 6312 865 6324 868
rect 6360 865 6372 912
rect 6384 865 6396 868
rect 6456 865 6468 868
rect 6528 865 6540 1042
rect 48 63 60 66
rect 168 0 180 66
rect 197 0 209 49
rect 336 0 348 66
rect 528 0 540 66
rect 768 63 780 66
rect 816 63 828 66
rect 816 0 828 49
rect 960 0 972 66
rect 1032 63 1044 66
rect 1296 0 1308 66
rect 1368 63 1380 66
rect 1656 0 1668 66
rect 1728 63 1740 66
rect 2064 0 2076 66
rect 2136 63 2148 66
rect 2400 0 2412 66
rect 2472 63 2484 66
rect 2712 0 2724 66
rect 2784 63 2796 66
rect 3048 0 3060 66
rect 3120 63 3132 66
rect 3216 0 3228 66
rect 3384 0 3396 66
rect 3504 41 3516 66
rect 3552 41 3564 66
rect 3600 41 3612 66
rect 3744 41 3756 66
rect 3960 41 3972 66
rect 4008 41 4020 66
rect 4152 41 4164 66
rect 4368 41 4380 66
rect 4512 41 4524 66
rect 4824 41 4836 66
rect 4920 41 4932 66
rect 3480 0 3492 27
rect 3528 0 3540 27
rect 3576 0 3588 27
rect 3624 0 3636 27
rect 3936 0 3948 27
rect 3984 0 3996 27
rect 4032 0 4044 27
rect 4344 0 4356 27
rect 4392 0 4404 27
rect 4776 0 4788 27
rect 4944 0 4956 66
rect 5040 41 5052 66
rect 5088 41 5100 66
rect 5136 41 5148 66
rect 4969 0 4981 27
rect 5016 0 5028 5
rect 5064 0 5076 27
rect 5112 0 5124 27
rect 5160 0 5172 27
rect 5232 19 5244 66
rect 5400 0 5412 66
rect 5496 41 5508 66
rect 5544 41 5556 66
rect 5472 0 5484 5
rect 5520 0 5532 27
rect 5568 0 5580 27
rect 5640 19 5652 66
rect 5808 0 5820 66
rect 5904 41 5916 66
rect 5880 0 5892 5
rect 5928 0 5940 27
rect 6000 19 6012 66
rect 6168 0 6180 66
rect 6312 41 6324 66
rect 6240 0 6252 27
rect 6528 0 6540 66
rect 6600 63 6612 66
use and2 and2_0
timestamp 1386234845
transform 1 0 0 0 1 66
box 0 0 120 799
use xor2 xor2_0
timestamp 1386237344
transform 1 0 120 0 1 66
box 0 0 192 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 312 0 1 66
box 0 0 48 799
use fulladder fulladder_0
timestamp 1386234928
transform 1 0 360 0 1 66
box 0 0 360 799
use or2 or2_0
timestamp 1386235472
transform 1 0 720 0 1 66
box 0 0 144 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 864 0 1 66
box 0 0 216 799
use and2 and2_1
timestamp 1386234845
transform 1 0 1080 0 1 66
box 0 0 120 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 1200 0 1 66
box 0 0 216 799
use or2 or2_1
timestamp 1386235472
transform 1 0 1416 0 1 66
box 0 0 144 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1560 0 1 66
box 0 0 216 799
use xor2 xor2_1
timestamp 1386237344
transform 1 0 1776 0 1 66
box 0 0 192 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 1968 0 1 66
box 0 0 216 799
use inv inv_0
timestamp 1386238110
transform 1 0 2184 0 1 66
box 0 0 120 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 2304 0 1 66
box 0 0 216 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 2520 0 1 66
box 0 0 96 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 2616 0 1 66
box 0 0 216 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 2832 0 1 66
box 0 0 120 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 2952 0 1 66
box 0 0 216 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 3168 0 1 66
box 0 0 192 799
use and2 and2_2
timestamp 1386234845
transform 1 0 3360 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 3480 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_2
timestamp 1386086759
transform 1 0 3528 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_3
timestamp 1386086759
transform 1 0 3576 0 1 66
box 0 0 48 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 3624 0 1 66
box 0 0 192 799
use and2 and2_3
timestamp 1386234845
transform 1 0 3816 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_7
timestamp 1386086759
transform 1 0 3936 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_10
timestamp 1386086759
transform 1 0 3984 0 1 66
box 0 0 48 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4032 0 1 66
box 0 0 192 799
use and2 and2_4
timestamp 1386234845
transform 1 0 4224 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_9
timestamp 1386086759
transform 1 0 4344 0 1 66
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 4392 0 1 66
box 0 0 192 799
use and2 and2_5
timestamp 1386234845
transform 1 0 4584 0 1 66
box 0 0 120 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 4704 0 1 66
box 0 0 192 799
use and2 and2_6
timestamp 1386234845
transform 1 0 4896 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_4
timestamp 1386086759
transform 1 0 5016 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_5
timestamp 1386086759
transform 1 0 5064 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_6
timestamp 1386086759
transform 1 0 5112 0 1 66
box 0 0 48 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 5160 0 1 66
box 0 0 192 799
use and2 and2_7
timestamp 1386234845
transform 1 0 5352 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_11
timestamp 1386086759
transform 1 0 5472 0 1 66
box 0 0 48 799
use rowcrosser rowcrosser_12
timestamp 1386086759
transform 1 0 5520 0 1 66
box 0 0 48 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 5568 0 1 66
box 0 0 192 799
use and2 and2_8
timestamp 1386234845
transform 1 0 5760 0 1 66
box 0 0 120 799
use rowcrosser rowcrosser_15
timestamp 1386086759
transform 1 0 5880 0 1 66
box 0 0 48 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 5928 0 1 66
box 0 0 192 799
use and2 and2_9
timestamp 1386234845
transform 1 0 6120 0 1 66
box 0 0 120 799
use mux2 mux2_8
timestamp 1386235218
transform 1 0 6240 0 1 66
box 0 0 192 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 6432 0 1 66
box 0 0 216 799
<< labels >>
rlabel metal1 0 870 0 880 3 A
rlabel metal1 0 892 0 902 3 B
rlabel metal1 6648 51 6648 61 7 ALUOut
rlabel metal2 6168 0 6180 0 1 Sh1
rlabel metal2 5808 0 5820 0 1 Sh2
rlabel metal2 5400 0 5412 0 1 Sh4
rlabel metal2 4944 0 4956 0 1 Sh8
rlabel metal2 197 0 209 0 1 ZeroA
rlabel metal2 168 0 180 0 1 SUB
rlabel metal2 816 0 828 0 1 nZ
rlabel metal2 3216 0 3228 0 1 ShB
rlabel metal2 6528 0 6540 0 1 ShOut
rlabel metal2 6240 0 6252 0 1 Sh1A_R
rlabel metal2 5928 0 5940 0 1 Sh2B_R
rlabel metal2 5880 0 5892 0 1 Sh2A_R
rlabel metal2 5568 0 5580 0 1 Sh4C_R
rlabel metal2 5520 0 5532 0 1 Sh4B_R
rlabel metal2 5472 0 5484 0 1 Sh4A_R
rlabel metal2 5160 0 5172 0 1 Sh8D_R
rlabel metal2 5112 0 5124 0 1 Sh8C_R
rlabel metal2 5064 0 5076 0 1 Sh8B_R
rlabel metal2 5016 0 5028 0 1 Sh8A_R
rlabel metal2 4969 0 4981 0 1 ShR
rlabel metal2 4776 0 4788 0 1 Sh1A_L
rlabel metal2 4392 0 4404 0 1 Sh2B_L
rlabel metal2 4344 0 4356 0 1 Sh2A_L
rlabel metal2 4032 0 4044 0 1 Sh4C_L
rlabel metal2 3984 0 3996 0 1 Sh4B_L
rlabel metal2 3936 0 3948 0 1 Sh4A_L
rlabel metal2 3624 0 3636 0 1 Sh8D_L
rlabel metal2 3576 0 3588 0 1 Sh8C_L
rlabel metal2 3528 0 3540 0 1 Sh8B_L
rlabel metal2 3480 0 3492 0 1 Sh8A_L
rlabel metal2 3384 0 3396 0 1 ShL
rlabel metal2 3048 0 3060 0 1 NOR
rlabel metal2 2712 0 2724 0 1 NAND
rlabel metal2 2400 0 2412 0 1 NOT
rlabel metal2 2064 0 2076 0 1 XOR
rlabel metal2 1656 0 1668 0 1 OR
rlabel metal2 1296 0 1308 0 1 AND
rlabel metal2 528 0 540 0 1 CIn_slice
rlabel metal2 336 0 348 0 1 CIn
rlabel metal2 960 0 972 0 1 FAOut
rlabel metal1 6648 892 6648 902 7 B
rlabel metal2 3384 1042 3396 1042 5 ShL
rlabel metal2 4969 1042 4981 1042 5 ShR
rlabel metal2 4344 1042 4356 1042 5 Sh2A_L
rlabel metal2 4392 1042 4404 1042 5 Sh2B_L
rlabel metal2 4776 1042 4788 1042 5 Sh1A_L
rlabel metal2 3480 1042 3492 1042 5 Sh8A_L
rlabel metal2 3528 1042 3540 1042 5 Sh8B_L
rlabel metal2 3576 1042 3588 1042 5 Sh8C_L
rlabel metal2 3624 1042 3636 1042 5 Sh8D_L
rlabel metal2 3936 1042 3948 1042 5 Sh4A_L
rlabel metal2 3984 1042 3996 1042 5 Sh4B_L
rlabel metal2 4032 1042 4044 1042 5 Sh4C_L
rlabel metal2 5016 1042 5028 1042 5 Sh8A_R
rlabel metal2 5064 1042 5076 1042 5 Sh8B_R
rlabel metal2 5112 1042 5124 1042 5 Sh8C_R
rlabel metal2 5472 1042 5484 1042 5 Sh4A_R
rlabel metal2 5520 1042 5532 1042 5 Sh4B_R
rlabel metal2 5568 1042 5580 1042 5 Sh4C_R
rlabel metal2 5880 1042 5892 1042 5 Sh2A_R
rlabel metal2 5928 1042 5940 1042 5 Sh2B_R
rlabel metal2 6240 1042 6252 1042 5 Sh1A_R
rlabel metal2 6528 1042 6540 1042 5 ShOut
rlabel metal2 5160 1042 5172 1042 5 Sh8D_R
rlabel metal2 4944 1042 4956 1042 5 Sh8
rlabel metal2 5400 1042 5412 1042 5 Sh4
rlabel metal2 5808 1042 5820 1042 5 Sh2
rlabel metal2 6168 1042 6180 1042 5 Sh1
rlabel metal2 960 1042 972 1042 5 FAOut
rlabel metal2 816 1042 828 1042 5 nZ
rlabel metal2 168 1042 180 1042 5 SUB
rlabel metal2 197 1042 209 1042 5 ZeroA
rlabel metal2 1296 1042 1308 1042 5 AND
rlabel metal2 1656 1042 1668 1042 5 OR
rlabel metal2 2064 1042 2076 1042 5 XOR
rlabel metal2 2400 1042 2412 1042 5 NOT
rlabel metal2 2712 1042 2724 1042 5 NAND
rlabel metal2 3048 1042 3060 1042 5 NOR
rlabel metal2 3216 1042 3228 1042 5 ShB
rlabel metal2 504 1042 516 1042 5 LastCIn
rlabel metal2 528 1042 540 1042 5 COut
rlabel metal2 600 1042 612 1042 5 Sum
rlabel metal2 3168 1042 3180 1042 5 ASign
rlabel metal2 336 1042 348 1042 5 CIn
<< end >>
