../../../Design/Implementation/verilog/behavioural/alu.sv