magic
tech c035u
timestamp 1394232814
<< metal1 >>
rect 172 951 2533 961
rect 1227 928 1669 938
rect 55 899 181 909
rect 387 903 1621 913
rect 387 878 493 888
rect 579 873 637 883
rect 1708 868 1812 878
rect 1899 873 1957 883
rect 2547 863 2677 873
rect 0 835 110 845
rect 2870 835 2935 845
rect 0 788 42 799
rect 56 788 110 799
rect 0 774 110 788
rect 2870 774 2935 799
rect 0 129 110 154
rect 2870 129 2935 154
rect 0 106 110 116
rect 2870 106 2935 116
rect 0 83 110 93
rect 2870 83 2935 93
rect 0 60 110 70
rect 2870 60 2935 70
rect 0 2 541 12
rect 555 2 1500 12
rect 1516 2 2820 12
rect 2836 2 2935 12
<< m2contact >>
rect 158 949 172 963
rect 2533 949 2548 963
rect 1213 927 1227 941
rect 1669 927 1683 941
rect 41 898 55 912
rect 181 898 195 912
rect 373 903 387 917
rect 1621 901 1635 915
rect 373 877 387 891
rect 493 876 507 890
rect 565 872 579 886
rect 637 871 651 885
rect 1693 866 1708 880
rect 1812 867 1827 881
rect 1885 872 1899 886
rect 1957 871 1971 885
rect 2532 861 2547 875
rect 2677 862 2691 876
rect 42 788 56 802
rect 541 1 555 15
rect 1500 1 1516 15
rect 2820 0 2836 14
<< metal2 >>
rect 42 802 54 898
rect 158 852 170 949
rect 182 852 194 898
rect 374 891 386 903
rect 374 852 386 877
rect 470 852 482 978
rect 494 852 506 876
rect 566 852 578 872
rect 638 852 650 871
rect 686 852 698 978
rect 1214 883 1226 927
rect 1214 871 1370 883
rect 1214 852 1226 871
rect 1358 852 1370 871
rect 1430 852 1442 978
rect 1598 852 1610 978
rect 1622 852 1634 901
rect 1670 852 1682 927
rect 1694 852 1706 866
rect 1790 852 1802 978
rect 1814 852 1826 867
rect 1862 852 1874 978
rect 1886 852 1898 872
rect 1958 852 1970 871
rect 2006 852 2018 978
rect 2534 875 2546 949
rect 2534 852 2546 861
rect 2678 852 2690 862
rect 2750 852 2762 978
rect 542 15 554 53
rect 1502 15 1514 53
rect 2822 14 2834 53
use halfadder halfadder_0
timestamp 1386235204
transform 1 0 110 0 1 53
box 0 0 312 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 422 0 1 53
box 0 0 192 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 614 0 1 53
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 1334 0 1 53
box 0 0 216 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 1550 0 1 53
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 1742 0 1 53
box 0 0 192 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 1934 0 1 53
box 0 0 720 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 2654 0 1 53
box 0 0 216 799
<< labels >>
rlabel metal1 2935 774 2935 799 7 Vdd!
rlabel metal1 2935 835 2935 845 7 ScanReturn
rlabel metal1 2935 129 2935 154 7 GND!
rlabel metal1 2935 60 2935 70 7 nReset
rlabel metal1 2935 83 2935 93 7 Test
rlabel metal1 2935 106 2935 116 7 Clock
rlabel metal1 0 774 0 799 3 Vdd!
rlabel metal1 0 835 0 845 3 ScanReturn
rlabel metal1 0 60 0 70 3 nReset
rlabel metal1 0 83 0 93 3 Test
rlabel metal1 0 106 0 116 3 Clock
rlabel metal1 0 129 0 154 3 GND!
rlabel metal2 2750 978 2762 978 1 PcEn
rlabel metal2 2006 978 2018 978 1 PcWe
rlabel metal2 1862 978 1874 978 1 ALU
rlabel metal2 1790 978 1802 978 1 PcSel[1]
rlabel metal2 1598 978 1610 978 1 PcSel[0]
rlabel metal2 1430 978 1442 978 1 LrEn
rlabel metal2 686 978 698 978 1 LrWe
rlabel metal2 470 978 482 978 1 LrSel
rlabel metal1 0 2 0 12 3 DataBus
rlabel metal1 2935 2 2935 12 7 DataBus
<< end >>
