magic
tech c035u
timestamp 1394111260
<< metal1 >>
rect 0 920 81 930
rect 95 920 201 930
rect 215 920 441 930
rect 455 920 777 930
rect 791 920 1017 930
rect 1031 920 1137 930
rect 1151 920 1353 930
rect 1367 920 1689 930
rect 0 898 57 908
rect 71 898 177 908
rect 191 898 561 908
rect 575 898 681 908
rect 695 898 897 908
rect 911 898 1233 908
rect 1247 898 1329 908
rect 1343 898 1569 908
rect 1583 898 1703 908
rect 0 875 33 885
rect 47 875 321 885
rect 335 875 417 885
rect 431 875 657 885
rect 671 875 873 885
rect 887 875 1113 885
rect 1127 875 1449 885
rect 1463 875 1545 885
rect 1559 875 1703 885
rect 0 827 10 837
rect 0 804 10 814
rect 0 766 10 791
rect 0 98 10 108
rect 0 75 10 85
rect 0 52 10 62
<< m2contact >>
rect 81 918 95 932
rect 201 918 215 932
rect 441 918 455 932
rect 777 918 791 932
rect 1017 918 1031 932
rect 1137 918 1151 932
rect 1353 918 1367 932
rect 1689 918 1703 932
rect 57 896 71 910
rect 177 896 191 910
rect 561 896 575 910
rect 681 896 695 910
rect 897 896 911 910
rect 1233 896 1247 910
rect 1329 896 1343 910
rect 1569 896 1583 910
rect 33 873 47 887
rect 321 873 335 887
rect 417 873 431 887
rect 657 873 671 887
rect 873 873 887 887
rect 1113 873 1127 887
rect 1449 873 1463 887
rect 1545 873 1559 887
<< metal2 >>
rect 34 844 46 873
rect 58 844 70 896
rect 82 844 94 918
rect 178 844 190 896
rect 202 844 214 918
rect 322 844 334 873
rect 418 844 430 873
rect 442 844 454 918
rect 562 844 574 896
rect 658 844 670 873
rect 682 844 694 896
rect 778 844 790 918
rect 874 844 886 873
rect 898 844 910 896
rect 1018 844 1030 918
rect 1114 844 1126 873
rect 1138 844 1150 918
rect 1234 844 1246 896
rect 1330 844 1342 896
rect 1354 844 1366 918
rect 1450 844 1462 873
rect 1546 844 1558 873
rect 1570 844 1582 896
rect 1690 844 1702 918
rect 130 0 142 45
rect 250 33 310 45
rect 370 0 382 45
rect 490 33 550 45
rect 610 0 622 45
rect 706 33 766 45
rect 826 0 838 45
rect 946 33 1006 45
rect 1066 0 1078 45
rect 1162 33 1222 45
rect 1282 0 1294 45
rect 1378 33 1438 45
rect 1498 0 1510 45
rect 1618 33 1678 45
rect 1738 0 1750 45
use nor3 nor3_0
timestamp 1386235396
transform 1 0 10 0 1 45
box 0 0 144 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 154 0 1 45
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 274 0 1 45
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 394 0 1 45
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 514 0 1 45
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 634 0 1 45
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 730 0 1 45
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 850 0 1 45
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 970 0 1 45
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1090 0 1 45
box 0 0 96 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 1186 0 1 45
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 1306 0 1 45
box 0 0 96 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 1402 0 1 45
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 1522 0 1 45
box 0 0 120 799
use and2 and2_4
timestamp 1386234845
transform 1 0 1642 0 1 45
box 0 0 120 799
<< labels >>
rlabel metal2 130 0 142 0 1 Out[0]
rlabel metal2 370 0 382 0 1 Out[1]
rlabel metal2 610 0 622 0 1 Out[2]
rlabel metal2 826 0 838 0 1 Out[3]
rlabel metal2 1066 0 1078 0 1 Out[4]
rlabel metal2 1282 0 1294 0 1 Out[5]
rlabel metal2 1498 0 1510 0 1 Out[6]
rlabel metal2 1738 0 1750 0 1 Out[7]
rlabel metal1 0 875 0 885 3 In[0]
rlabel metal1 0 898 0 908 3 In[1]
rlabel metal1 0 920 0 930 4 In[2]
rlabel metal1 0 827 0 837 3 ScanReturn
rlabel metal1 0 804 0 814 3 Scan
rlabel metal1 0 766 0 791 3 Vdd!
rlabel metal1 0 52 0 62 3 nReset
rlabel metal1 0 75 0 85 3 Test
rlabel metal1 0 98 0 108 3 Clock
<< end >>
