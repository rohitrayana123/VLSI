../../../Design/Implementation/verilog/behavioural/cpu_core.sv