magic
tech c035u
timestamp 1396693766
<< metal1 >>
rect 21120 39730 21130 39773
rect 21168 39730 21178 39773
rect 21120 39720 21178 39730
rect 21120 39536 21130 39720
rect 21170 38937 21180 39561
rect 20306 38927 21180 38937
rect 20207 38832 20266 38842
rect 20256 38818 20266 38832
rect 20256 38808 20279 38818
rect 20306 38790 20316 38927
rect 20207 38780 20316 38790
rect 20280 34837 20290 38755
rect 20207 34776 20255 34786
rect 20306 34748 20316 38780
rect 20206 34738 20316 34748
rect 20256 30781 20266 34703
rect 20280 30781 20290 34703
rect 20306 30781 20316 34738
rect 21216 30781 21226 39773
rect 24545 39757 24559 39773
rect 24600 39730 24610 39773
rect 28071 39756 28081 39773
rect 21480 39720 24610 39730
rect 21480 39706 21490 39720
rect 28128 39730 28138 39773
rect 28199 39742 31546 39752
rect 31584 39730 31594 39773
rect 31632 39757 31642 39773
rect 31776 39757 31786 39773
rect 38640 39730 38650 39773
rect 38688 39757 38698 39773
rect 38832 39757 38842 39773
rect 42168 39730 42178 39773
rect 42216 39757 42226 39773
rect 42360 39757 42370 39773
rect 45696 39730 45706 39773
rect 45744 39757 45754 39773
rect 45888 39757 45898 39773
rect 47338 39752 47506 39753
rect 46812 39743 47506 39752
rect 46812 39742 47352 39743
rect 46812 39730 46822 39742
rect 28117 39720 28138 39730
rect 28152 39720 46823 39730
rect 46848 39720 47459 39730
rect 21456 39696 21490 39706
rect 21456 39658 21466 39696
rect 28152 39706 28162 39720
rect 21517 39696 28162 39706
rect 46848 39706 46858 39720
rect 31645 39696 46858 39706
rect 46872 39696 47436 39706
rect 21480 39672 28103 39682
rect 21480 39661 21490 39672
rect 21432 39648 21466 39658
rect 21432 39325 21442 39648
rect 21480 39301 21490 39599
rect 21504 39274 21514 39599
rect 31776 39589 31786 39672
rect 46872 39682 46882 39696
rect 38845 39672 46882 39682
rect 31822 39649 38660 39659
rect 38650 39609 38660 39649
rect 38688 39634 38698 39671
rect 45901 39648 47338 39658
rect 38688 39624 47314 39634
rect 38650 39599 46725 39609
rect 21614 39566 24545 39576
rect 27888 39552 47219 39562
rect 27888 39469 27898 39552
rect 45757 39528 46961 39538
rect 47209 39537 47219 39552
rect 31776 39469 31786 39527
rect 38869 39504 47183 39514
rect 38664 39480 47231 39490
rect 38664 39469 38674 39480
rect 39037 39456 46991 39466
rect 47304 39445 47314 39624
rect 21456 39264 21514 39274
rect 25464 39432 47279 39442
rect 21456 39253 21466 39264
rect 21384 39168 22138 39178
rect 21384 30754 21394 39168
rect 22128 39157 22138 39168
rect 25464 39157 25474 39432
rect 26856 39408 47135 39418
rect 26856 39373 26866 39408
rect 47328 39408 47338 39648
rect 36144 39384 47063 39394
rect 36144 39373 36154 39384
rect 36877 39360 47255 39370
rect 26664 39336 47015 39346
rect 26664 39277 26674 39336
rect 35880 39312 47122 39322
rect 26856 39277 26866 39311
rect 27888 39277 27898 39311
rect 31776 39277 31786 39311
rect 35880 39277 35890 39312
rect 47112 39301 47122 39312
rect 47317 39312 47399 39322
rect 38928 39288 47087 39298
rect 38928 39277 38938 39288
rect 47426 39288 47436 39696
rect 42373 39264 45743 39274
rect 45781 39264 47314 39274
rect 47304 39253 47314 39264
rect 47449 39261 47459 39720
rect 25704 39240 47159 39250
rect 25704 39157 25714 39240
rect 31789 39216 47482 39226
rect 26664 39157 26674 39215
rect 26856 39157 26866 39215
rect 27888 39157 27898 39215
rect 42229 39192 46882 39202
rect 46872 39178 46882 39192
rect 46975 39192 47386 39202
rect 46872 39168 47362 39178
rect 20207 30744 21394 30754
rect 20207 30696 20303 30706
rect 20256 26916 20266 30671
rect 20280 26943 20290 30671
rect 21216 26919 21226 30719
rect 20256 26906 20314 26916
rect 20207 22800 20266 22810
rect 20256 18805 20266 22800
rect 20280 19618 20290 26857
rect 20304 19645 20314 26906
rect 21216 19645 21226 26857
rect 21432 19669 21442 39143
rect 21456 19669 21466 39143
rect 21480 19642 21490 39143
rect 46992 36469 47002 39143
rect 47016 36469 47026 39143
rect 47064 36469 47074 39143
rect 47088 36469 47098 39143
rect 47112 36469 47122 39143
rect 47136 36469 47146 39143
rect 47160 36469 47170 39143
rect 47184 36469 47194 39143
rect 47208 36469 47218 39143
rect 47232 36469 47242 39143
rect 47256 36469 47266 39143
rect 47280 36469 47290 39143
rect 47304 36469 47314 39143
rect 47328 36469 47338 39143
rect 47352 36469 47362 39168
rect 47376 36469 47386 39192
rect 47400 36469 47410 39191
rect 47424 36469 47434 39191
rect 47448 36469 47458 39191
rect 47472 36442 47482 39216
rect 47496 39034 47506 39743
rect 47496 39024 50307 39034
rect 50256 39013 50266 39024
rect 50232 38976 50307 38986
rect 50232 38893 50242 38976
rect 50256 38866 50266 38951
rect 46968 36440 47482 36442
rect 46943 36432 47482 36440
rect 50208 38856 50266 38866
rect 46943 36430 46978 36432
rect 46943 36370 46978 36374
rect 47448 36370 47458 36407
rect 46943 36364 47458 36370
rect 46968 36360 47458 36364
rect 46992 35365 47002 36335
rect 47016 35365 47026 36335
rect 47064 35365 47074 36335
rect 47088 35365 47098 36335
rect 47112 35365 47122 36335
rect 47136 35365 47146 36335
rect 47160 35365 47170 36335
rect 47184 35365 47194 36335
rect 47208 35365 47218 36335
rect 47232 35365 47242 36335
rect 47256 35365 47266 36335
rect 47280 35365 47290 36335
rect 47304 35365 47314 36335
rect 47328 35365 47338 36335
rect 47352 35365 47362 36335
rect 47376 35365 47386 36335
rect 47400 35365 47410 36335
rect 47424 35338 47434 36335
rect 46968 35329 47434 35338
rect 46943 35328 47434 35329
rect 46943 35319 46978 35328
rect 47400 35266 47410 35303
rect 46968 35263 47410 35266
rect 46943 35256 47410 35263
rect 46943 35253 46978 35256
rect 46992 34237 47002 35231
rect 47016 34237 47026 35231
rect 47064 34237 47074 35231
rect 47088 34237 47098 35231
rect 47112 34237 47122 35231
rect 47136 34237 47146 35231
rect 47160 34237 47170 35231
rect 47184 34237 47194 35231
rect 47208 34237 47218 35231
rect 47232 34237 47242 35231
rect 47256 34237 47266 35231
rect 47280 34237 47290 35231
rect 47304 34237 47314 35231
rect 47328 34237 47338 35231
rect 47352 34237 47362 35231
rect 46943 34210 46978 34218
rect 47376 34210 47386 35231
rect 50208 35005 50218 38856
rect 50256 38832 50307 38842
rect 50232 35029 50242 38831
rect 50256 35029 50266 38832
rect 50221 34992 50307 35002
rect 50184 34968 50231 34978
rect 50184 34861 50194 34968
rect 50232 34944 50307 34954
rect 50208 34861 50218 34943
rect 50232 34861 50242 34944
rect 50256 34834 50266 34919
rect 46943 34208 47386 34210
rect 46968 34200 47386 34208
rect 50160 34824 50266 34834
rect 46943 34142 46978 34152
rect 46968 34138 46978 34142
rect 47352 34138 47362 34175
rect 46968 34128 47362 34138
rect 46992 33133 47002 34103
rect 47016 33133 47026 34103
rect 47064 33133 47074 34103
rect 47088 33133 47098 34103
rect 47112 33133 47122 34103
rect 47136 33133 47146 34103
rect 47160 33133 47170 34103
rect 47184 33133 47194 34103
rect 47208 33133 47218 34103
rect 47232 33133 47242 34103
rect 47256 33133 47266 34103
rect 47280 33133 47290 34103
rect 47304 33133 47314 34103
rect 46943 33106 46978 33107
rect 47328 33106 47338 34103
rect 46943 33097 47338 33106
rect 46968 33096 47338 33097
rect 46943 33034 46978 33041
rect 47304 33034 47314 33071
rect 46943 33031 47314 33034
rect 46968 33024 47314 33031
rect 46992 32029 47002 32999
rect 47016 32029 47026 32999
rect 47064 32029 47074 32999
rect 47088 32029 47098 32999
rect 47112 32029 47122 32999
rect 47136 32029 47146 32999
rect 47160 32029 47170 32999
rect 47184 32029 47194 32999
rect 47208 32029 47218 32999
rect 47232 32029 47242 32999
rect 47256 32029 47266 32999
rect 47280 32029 47290 32999
rect 50160 32002 50170 34824
rect 50256 34800 50307 34810
rect 46968 31996 50170 32002
rect 46943 31992 50170 31996
rect 46943 31986 46978 31992
rect 50184 31930 50194 34799
rect 46943 31920 50194 31930
rect 46992 30901 47002 31895
rect 47016 30901 47026 31895
rect 47064 30901 47074 31895
rect 47088 30901 47098 31895
rect 47112 30901 47122 31895
rect 47136 30901 47146 31895
rect 47160 30901 47170 31895
rect 47184 30901 47194 31895
rect 47208 30901 47218 31895
rect 47232 30901 47242 31895
rect 47256 30901 47266 31895
rect 47280 30901 47290 31895
rect 50208 30970 50218 34799
rect 50232 30997 50242 34799
rect 50256 30997 50266 34800
rect 50208 30960 50307 30970
rect 50208 30936 50255 30946
rect 46943 30875 46978 30885
rect 46968 30874 46978 30875
rect 50208 30874 50218 30936
rect 50256 30912 50307 30922
rect 46968 30864 50218 30874
rect 50232 30826 50242 30911
rect 46968 30819 50242 30826
rect 46943 30816 50242 30819
rect 46943 30809 46978 30816
rect 50256 30805 50266 30912
rect 46992 29797 47002 30791
rect 47016 29797 47026 30791
rect 47064 29797 47074 30791
rect 47088 29797 47098 30791
rect 47112 29797 47122 30791
rect 47136 29797 47146 30791
rect 47160 29797 47170 30791
rect 47184 29797 47194 30791
rect 47208 29797 47218 30791
rect 47232 29797 47242 30791
rect 47256 29797 47266 30791
rect 47280 29797 47290 30791
rect 50232 30768 50307 30778
rect 46943 29770 46978 29774
rect 50232 29770 50242 30768
rect 46943 29764 50242 29770
rect 46968 29760 50242 29764
rect 46943 29698 46978 29708
rect 50256 29698 50266 30743
rect 46968 29688 50266 29698
rect 46992 28693 47002 29663
rect 47016 28693 47026 29663
rect 47064 28693 47074 29663
rect 47088 28693 47098 29663
rect 47112 28693 47122 29663
rect 47136 28693 47146 29663
rect 47160 28693 47170 29663
rect 47184 28693 47194 29663
rect 47208 28690 47218 29663
rect 47232 28717 47242 29663
rect 47256 28717 47266 29663
rect 47280 28717 47290 29663
rect 47208 28680 47314 28690
rect 46968 28663 47218 28666
rect 46943 28656 47218 28663
rect 46943 28653 46978 28656
rect 47208 28645 47218 28656
rect 47304 28645 47314 28680
rect 47064 28618 47074 28631
rect 47064 28608 47338 28618
rect 46943 28594 46978 28597
rect 46943 28587 47074 28594
rect 46968 28584 47074 28587
rect 46992 27565 47002 28559
rect 47016 27565 47026 28559
rect 46943 27542 46978 27552
rect 47064 27562 47074 28584
rect 47088 27589 47098 28583
rect 47112 27589 47122 28583
rect 47136 27589 47146 28583
rect 47160 27589 47170 28583
rect 47184 27589 47194 28583
rect 47208 27589 47218 28583
rect 47232 27589 47242 28583
rect 47256 27589 47266 28583
rect 47280 27589 47290 28583
rect 47304 27589 47314 28583
rect 47328 27589 47338 28608
rect 47064 27552 47362 27562
rect 46968 27538 46978 27542
rect 47352 27541 47362 27552
rect 46968 27528 47063 27538
rect 46968 27486 47050 27490
rect 46943 27480 47050 27486
rect 46943 27476 46978 27480
rect 46992 26461 47002 27455
rect 47016 26461 47026 27455
rect 47040 26461 47050 27480
rect 47064 26461 47074 27479
rect 47088 26461 47098 27479
rect 47112 26458 47122 27479
rect 47136 26485 47146 27479
rect 47160 26485 47170 27479
rect 47184 26485 47194 27479
rect 47208 26485 47218 27479
rect 47232 26485 47242 27479
rect 47256 26485 47266 27479
rect 47280 26485 47290 27479
rect 47304 26485 47314 27479
rect 47328 26485 47338 27479
rect 47352 26485 47362 27479
rect 47112 26448 47386 26458
rect 46943 26434 46978 26441
rect 46943 26431 47122 26434
rect 46968 26424 47122 26431
rect 47112 26413 47122 26424
rect 47376 26413 47386 26448
rect 47016 26386 47026 26399
rect 47016 26376 47410 26386
rect 46943 26365 46978 26375
rect 46968 26362 46978 26365
rect 46968 26352 47026 26362
rect 46992 25357 47002 26327
rect 47016 25357 47026 26352
rect 47040 25357 47050 26351
rect 47064 25357 47074 26351
rect 47088 25357 47098 26351
rect 47112 25357 47122 26351
rect 47136 25357 47146 26351
rect 47160 25357 47170 26351
rect 47184 25354 47194 26351
rect 47208 25381 47218 26351
rect 47232 25381 47242 26351
rect 47256 25381 47266 26351
rect 47280 25381 47290 26351
rect 47304 25381 47314 26351
rect 47328 25381 47338 26351
rect 47352 25381 47362 26351
rect 47376 25381 47386 26351
rect 47400 25381 47410 26376
rect 47184 25344 47434 25354
rect 46943 25320 47194 25330
rect 47184 25309 47194 25320
rect 47424 25309 47434 25344
rect 47088 25282 47098 25295
rect 47088 25272 47458 25282
rect 46943 25258 46978 25264
rect 46943 25254 47098 25258
rect 46968 25248 47098 25254
rect 46992 24250 47002 25223
rect 47016 24277 47026 25223
rect 47040 24277 47050 25223
rect 47064 24277 47074 25223
rect 47088 24277 47098 25248
rect 47112 24277 47122 25247
rect 47136 24277 47146 25247
rect 47160 24277 47170 25247
rect 47184 24277 47194 25247
rect 47208 24277 47218 25247
rect 47232 24277 47242 25247
rect 47256 24277 47266 25247
rect 47280 24277 47290 25247
rect 47304 24277 47314 25247
rect 47328 24277 47338 25247
rect 47352 24277 47362 25247
rect 47376 24277 47386 25247
rect 47400 24277 47410 25247
rect 47424 24277 47434 25247
rect 47448 24277 47458 25272
rect 46992 24240 47482 24250
rect 46968 24219 47002 24226
rect 46943 24216 47002 24219
rect 46943 24209 46978 24216
rect 46992 24181 47002 24216
rect 47016 24181 47026 24215
rect 47040 24181 47050 24215
rect 47064 24181 47074 24215
rect 47088 24181 47098 24215
rect 47112 24181 47122 24215
rect 47136 24181 47146 24215
rect 47160 24178 47170 24215
rect 47472 24205 47482 24240
rect 47160 24168 47506 24178
rect 46968 24153 47170 24154
rect 46943 24144 47170 24153
rect 46943 24143 46978 24144
rect 46992 23125 47002 24119
rect 47016 23125 47026 24119
rect 47040 23125 47050 24119
rect 47064 23125 47074 24119
rect 47088 23125 47098 24119
rect 47112 23125 47122 24119
rect 47136 23122 47146 24119
rect 47160 23149 47170 24144
rect 47184 23149 47194 24143
rect 47208 23149 47218 24143
rect 47232 23149 47242 24143
rect 47256 23149 47266 24143
rect 47280 23149 47290 24143
rect 47304 23149 47314 24143
rect 47328 23149 47338 24143
rect 47352 23149 47362 24143
rect 47376 23149 47386 24143
rect 47400 23149 47410 24143
rect 47424 23149 47434 24143
rect 47448 23149 47458 24143
rect 47472 23149 47482 24143
rect 47496 23149 47506 24168
rect 47136 23112 47530 23122
rect 46943 23098 46978 23108
rect 47520 23101 47530 23112
rect 46968 23088 47146 23098
rect 47136 23077 47146 23088
rect 47376 23074 47386 23087
rect 47376 23064 47554 23074
rect 46968 23042 47386 23050
rect 46943 23040 47386 23042
rect 46943 23032 46978 23040
rect 46992 22021 47002 23015
rect 47016 22021 47026 23015
rect 47040 22021 47050 23015
rect 47064 22021 47074 23015
rect 47088 22021 47098 23015
rect 47112 22021 47122 23015
rect 47136 22021 47146 23015
rect 47160 22021 47170 23015
rect 47184 22021 47194 23015
rect 47208 22021 47218 23015
rect 47232 22021 47242 23015
rect 47256 22018 47266 23015
rect 47280 22045 47290 23015
rect 47304 22045 47314 23015
rect 47328 22045 47338 23015
rect 47352 22045 47362 23015
rect 47376 22045 47386 23040
rect 47400 22045 47410 23039
rect 47424 22045 47434 23039
rect 47448 22045 47458 23039
rect 47472 22045 47482 23039
rect 47496 22045 47506 23039
rect 47520 22045 47530 23039
rect 47544 22045 47554 23064
rect 47256 22008 47578 22018
rect 46943 21994 46978 21997
rect 46943 21987 47266 21994
rect 46968 21984 47266 21987
rect 47256 21973 47266 21984
rect 47568 21973 47578 22008
rect 47088 21946 47098 21959
rect 47088 21936 47602 21946
rect 46943 21922 46978 21931
rect 46943 21921 47098 21922
rect 46968 21912 47098 21921
rect 46992 20917 47002 21887
rect 47016 20917 47026 21887
rect 47040 20917 47050 21887
rect 47064 20917 47074 21887
rect 47088 20917 47098 21912
rect 47112 20917 47122 21911
rect 47136 20917 47146 21911
rect 47160 20917 47170 21911
rect 47184 20917 47194 21911
rect 47208 20917 47218 21911
rect 47232 20917 47242 21911
rect 47256 20917 47266 21911
rect 47280 20917 47290 21911
rect 47304 20917 47314 21911
rect 47328 20917 47338 21911
rect 47352 20917 47362 21911
rect 47376 20917 47386 21911
rect 47400 20917 47410 21911
rect 47424 20917 47434 21911
rect 47448 20917 47458 21911
rect 47472 20917 47482 21911
rect 47496 20917 47506 21911
rect 47520 20917 47530 21911
rect 47544 20914 47554 21911
rect 47568 20941 47578 21911
rect 47592 20941 47602 21936
rect 47544 20904 47626 20914
rect 46968 20886 47554 20890
rect 46943 20880 47554 20886
rect 46943 20876 46978 20880
rect 47544 20869 47554 20880
rect 47616 20869 47626 20904
rect 46992 20842 47002 20855
rect 46992 20832 47650 20842
rect 46943 20818 46978 20820
rect 46943 20810 47002 20818
rect 46968 20808 47002 20810
rect 46992 19789 47002 20808
rect 47016 19789 47026 20807
rect 47040 19789 47050 20807
rect 47064 19789 47074 20807
rect 47088 19789 47098 20807
rect 47112 19786 47122 20807
rect 47136 19813 47146 20807
rect 47160 19813 47170 20807
rect 47184 19813 47194 20807
rect 47208 19813 47218 20807
rect 47232 19813 47242 20807
rect 47256 19813 47266 20807
rect 47280 19813 47290 20807
rect 47304 19813 47314 20807
rect 47328 19813 47338 20807
rect 47352 19813 47362 20807
rect 47376 19813 47386 20807
rect 47400 19813 47410 20807
rect 47424 19813 47434 20807
rect 47448 19813 47458 20807
rect 47472 19813 47482 20807
rect 47496 19813 47506 20807
rect 47520 19813 47530 20807
rect 47544 19813 47554 20807
rect 47568 19813 47578 20807
rect 47592 19813 47602 20807
rect 47616 19813 47626 20807
rect 47640 19813 47650 20832
rect 47112 19776 47674 19786
rect 46943 19765 46978 19775
rect 47664 19765 47674 19776
rect 46968 19762 46978 19765
rect 46968 19752 47122 19762
rect 47112 19741 47122 19752
rect 47256 19738 47266 19751
rect 47256 19728 47698 19738
rect 46968 19709 47266 19714
rect 46943 19704 47266 19709
rect 46943 19699 46978 19704
rect 21397 19632 21490 19642
rect 20280 19608 21490 19618
rect 20207 18768 20290 18778
rect 20256 14749 20266 18743
rect 20280 18442 20290 18768
rect 20304 18469 20314 19583
rect 21216 18469 21226 19583
rect 21384 18469 21394 19583
rect 21432 18469 21442 19583
rect 21456 18469 21466 19583
rect 21480 18469 21490 19608
rect 21534 19599 21544 19607
rect 21528 19589 21544 19599
rect 21582 19594 21592 19607
rect 23448 19594 23458 19607
rect 21528 18562 21538 19589
rect 21582 19584 23434 19594
rect 23448 19584 27599 19594
rect 21552 19567 21558 19579
rect 21552 18589 21562 19567
rect 23424 19570 23434 19584
rect 27624 19594 27634 19607
rect 27624 19584 37439 19594
rect 37464 19594 37474 19607
rect 37464 19584 41242 19594
rect 23424 19560 24226 19570
rect 21604 19544 21614 19559
rect 21600 19534 21614 19544
rect 21651 19546 21661 19559
rect 24216 19546 24226 19560
rect 24253 19560 26687 19570
rect 26725 19560 37199 19570
rect 37237 19560 40444 19570
rect 21651 19536 24202 19546
rect 24216 19536 27431 19546
rect 21600 18610 21610 19534
rect 21624 19518 21627 19529
rect 21624 18637 21634 19518
rect 24192 19522 24202 19536
rect 27469 19536 37018 19546
rect 24192 19512 24778 19522
rect 21672 18637 21682 19511
rect 24768 19498 24778 19512
rect 24805 19512 26471 19522
rect 37008 19522 37018 19536
rect 37045 19536 40420 19546
rect 26509 19512 36423 19522
rect 37008 19512 39490 19522
rect 24768 19488 24994 19498
rect 21696 18637 21706 19487
rect 24984 19474 24994 19488
rect 25021 19488 26279 19498
rect 26317 19488 36399 19498
rect 24984 19464 25738 19474
rect 25728 19450 25738 19464
rect 25765 19464 25906 19474
rect 25896 19450 25906 19464
rect 25933 19464 34810 19474
rect 25728 19440 25810 19450
rect 25896 19440 33994 19450
rect 25800 18637 25810 19440
rect 26293 19416 33970 19426
rect 26485 19392 33154 19402
rect 26701 19368 32050 19378
rect 27445 19344 27466 19354
rect 21600 18600 27034 18610
rect 27024 18589 27034 18600
rect 27456 18589 27466 19344
rect 27613 19344 31162 19354
rect 21528 18552 29794 18562
rect 21685 18528 24994 18538
rect 21552 18469 21562 18527
rect 21624 18490 21634 18527
rect 24984 18517 24994 18528
rect 21733 18504 22168 18514
rect 21624 18480 25834 18490
rect 21709 18456 24178 18466
rect 24168 18445 24178 18456
rect 25824 18445 25834 18480
rect 27024 18445 27034 18527
rect 27456 18445 27466 18527
rect 20280 18432 22144 18442
rect 21565 18408 29074 18418
rect 20304 14749 20314 18407
rect 21216 14749 21226 18407
rect 21384 18197 21394 18407
rect 21432 18229 21442 18407
rect 21456 18229 21466 18407
rect 21480 18229 21490 18407
rect 29064 18397 29074 18408
rect 29784 18397 29794 18552
rect 31152 18445 31162 19344
rect 32040 18445 32050 19368
rect 33144 18445 33154 19392
rect 33960 18445 33970 19416
rect 33984 18445 33994 19440
rect 34800 18445 34810 19464
rect 36389 18445 36399 19488
rect 36413 18445 36423 19512
rect 37213 19488 37234 19498
rect 37224 18445 37234 19488
rect 37453 19488 38026 19498
rect 38016 18445 38026 19488
rect 39480 18445 39490 19512
rect 40410 18445 40420 19536
rect 40434 18445 40444 19560
rect 41232 18445 41242 19584
rect 45168 18514 45178 19607
rect 44437 18504 45178 18514
rect 45912 18514 45922 19607
rect 46128 18514 46138 19607
rect 45253 18504 45922 18514
rect 46032 18504 46138 18514
rect 46032 18490 46042 18504
rect 43645 18480 46042 18490
rect 46272 18490 46282 19607
rect 46069 18480 46282 18490
rect 43525 18456 45239 18466
rect 46320 18466 46330 19607
rect 45277 18456 46330 18466
rect 42829 18432 44423 18442
rect 46368 18442 46378 19607
rect 44461 18432 46378 18442
rect 30264 18408 43631 18418
rect 30264 18397 30274 18408
rect 46416 18418 46426 19607
rect 46488 19594 46498 19607
rect 46488 19584 46690 19594
rect 46680 19042 46690 19584
rect 46680 19032 46882 19042
rect 43656 18408 46426 18418
rect 43656 18397 43666 18408
rect 46872 18397 46882 19032
rect 46992 18418 47002 19679
rect 47016 18442 47026 19679
rect 47040 18466 47050 19679
rect 47064 18490 47074 19679
rect 47088 18514 47098 19679
rect 47112 18538 47122 19679
rect 47136 18562 47146 19679
rect 47160 18586 47170 19679
rect 47184 18610 47194 19679
rect 47208 18634 47218 19679
rect 47232 18658 47242 19679
rect 47256 18682 47266 19704
rect 47280 18706 47290 19703
rect 47304 18730 47314 19703
rect 47328 18754 47338 19703
rect 47352 18778 47362 19703
rect 47376 18802 47386 19703
rect 47400 18826 47410 19703
rect 47424 18850 47434 19703
rect 47448 18874 47458 19703
rect 47472 18898 47482 19703
rect 47496 18922 47506 19703
rect 47520 18946 47530 19703
rect 47544 18970 47554 19703
rect 47568 18994 47578 19703
rect 47592 19018 47602 19703
rect 47616 19042 47626 19703
rect 47640 19066 47650 19703
rect 47664 19330 47674 19703
rect 47688 19354 47698 19728
rect 47688 19344 48191 19354
rect 47664 19320 48226 19330
rect 48192 19090 48202 19295
rect 48216 19114 48226 19320
rect 48216 19104 48359 19114
rect 48192 19080 48383 19090
rect 47640 19056 48407 19066
rect 47616 19032 48431 19042
rect 47592 19008 48455 19018
rect 47568 18984 48479 18994
rect 47544 18960 48503 18970
rect 47520 18936 48527 18946
rect 47496 18912 48551 18922
rect 47472 18888 48575 18898
rect 47448 18864 48599 18874
rect 47424 18840 48623 18850
rect 47400 18816 48647 18826
rect 50256 18816 50307 18826
rect 50256 18805 50266 18816
rect 47376 18792 48671 18802
rect 47352 18768 50307 18778
rect 47328 18744 48695 18754
rect 47304 18720 48719 18730
rect 47280 18696 48743 18706
rect 47256 18672 48767 18682
rect 50256 18661 50266 18743
rect 47232 18648 48839 18658
rect 47208 18624 50307 18634
rect 47184 18600 48863 18610
rect 47160 18576 48887 18586
rect 47136 18552 48911 18562
rect 47112 18528 48935 18538
rect 47088 18504 48983 18514
rect 47064 18480 50111 18490
rect 47040 18456 50159 18466
rect 47016 18432 50207 18442
rect 50256 18418 50266 18599
rect 46992 18408 48802 18418
rect 21720 18229 21730 18383
rect 21384 18187 21743 18197
rect 48360 18177 48370 18383
rect 48384 18177 48394 18383
rect 48408 18177 48418 18383
rect 48432 18177 48442 18383
rect 48456 18177 48466 18383
rect 21445 18163 21743 18173
rect 48480 18150 48490 18383
rect 48504 18153 48514 18383
rect 48528 18153 48538 18383
rect 48552 18153 48562 18383
rect 48576 18153 48586 18383
rect 48344 18140 48490 18150
rect 21456 14749 21466 18138
rect 21480 14749 21490 18138
rect 21720 14722 21730 18138
rect 48600 18126 48610 18383
rect 48624 18129 48634 18383
rect 48648 18129 48658 18383
rect 48672 18129 48682 18383
rect 48696 18129 48706 18383
rect 48720 18129 48730 18383
rect 48744 18129 48754 18383
rect 48768 18129 48778 18383
rect 48792 18129 48802 18408
rect 48816 18408 50266 18418
rect 48816 18129 48826 18408
rect 48344 18116 48610 18126
rect 48840 18102 48850 18383
rect 48344 18092 48850 18102
rect 48344 18068 48623 18078
rect 48344 18044 48575 18054
rect 20207 14712 21730 14722
rect 20256 10717 20266 14687
rect 20207 10680 20290 10690
rect 20256 10186 20266 10655
rect 20280 10234 20290 10680
rect 20304 10363 20314 14687
rect 21216 13980 21226 14687
rect 21456 14007 21466 14687
rect 21480 14007 21490 14687
rect 48360 14629 48370 18019
rect 48384 14629 48394 18019
rect 48408 14629 48418 18019
rect 48432 14629 48442 18019
rect 48456 14629 48466 18019
rect 48504 14629 48514 18019
rect 48528 14629 48538 18019
rect 48552 14629 48562 18019
rect 48648 14629 48658 18067
rect 48672 14629 48682 18067
rect 48696 14629 48706 18067
rect 48720 14629 48730 18067
rect 48744 14602 48754 18067
rect 48349 14592 48754 14602
rect 21216 13970 21743 13980
rect 21493 13946 21743 13956
rect 21456 10390 21466 13943
rect 48360 13213 48370 14567
rect 48384 13213 48394 14567
rect 48408 13213 48418 14567
rect 48432 13213 48442 14567
rect 48456 13213 48466 14567
rect 48504 13213 48514 14567
rect 48528 13213 48538 14567
rect 48552 13186 48562 14567
rect 48349 13176 48562 13186
rect 48360 12949 48370 13151
rect 48384 12949 48394 13151
rect 48408 12949 48418 13151
rect 48432 12949 48442 13151
rect 48456 12949 48466 13151
rect 48504 12949 48514 13151
rect 48528 12949 48538 13151
rect 48648 12922 48658 14567
rect 48349 12912 48658 12922
rect 48360 12613 48370 12887
rect 48384 12613 48394 12887
rect 48408 12613 48418 12887
rect 48432 12613 48442 12887
rect 48456 12613 48466 12887
rect 48504 12613 48514 12887
rect 48528 12586 48538 12887
rect 48349 12576 48538 12586
rect 48360 10813 48370 12551
rect 48384 10813 48394 12551
rect 48408 10813 48418 12551
rect 48432 10813 48442 12551
rect 48456 10813 48466 12551
rect 48504 10813 48514 12551
rect 48672 10813 48682 14567
rect 48696 10813 48706 14567
rect 48720 10786 48730 14567
rect 48349 10776 48730 10786
rect 48360 10546 48370 10751
rect 48384 10573 48394 10751
rect 48408 10573 48418 10751
rect 48432 10573 48442 10751
rect 48456 10573 48466 10751
rect 48504 10573 48514 10751
rect 48672 10573 48682 10751
rect 48696 10573 48706 10751
rect 48768 10573 48778 18067
rect 48792 10573 48802 18067
rect 48816 10738 48826 18067
rect 48864 10765 48874 18383
rect 48888 10765 48898 18383
rect 48912 10765 48922 18383
rect 48936 10765 48946 18383
rect 48984 10765 48994 18383
rect 50112 14602 50122 18383
rect 50160 14746 50170 18383
rect 50208 14773 50218 18383
rect 50256 14794 50266 18408
rect 50256 14784 50307 14794
rect 50160 14736 50307 14746
rect 50208 14629 50218 14711
rect 50112 14592 50307 14602
rect 50208 10765 50218 14567
rect 48816 10728 50307 10738
rect 50256 10717 50266 10728
rect 48864 10573 48874 10703
rect 48888 10573 48898 10703
rect 48912 10573 48922 10703
rect 48936 10573 48946 10703
rect 48984 10573 48994 10703
rect 50208 10690 50218 10703
rect 50208 10680 50307 10690
rect 50256 10573 50266 10655
rect 48360 10536 50307 10546
rect 48384 10391 48394 10511
rect 48408 10391 48418 10511
rect 48432 10391 48442 10511
rect 48456 10391 48466 10511
rect 48504 10391 48514 10511
rect 48672 10391 48682 10511
rect 20304 10353 21743 10363
rect 48696 10363 48706 10511
rect 48349 10353 48706 10363
rect 21720 10329 21743 10339
rect 21720 10261 21730 10329
rect 48349 10329 48431 10339
rect 48768 10333 48778 10511
rect 48792 10333 48802 10511
rect 48864 10333 48874 10511
rect 48888 10333 48898 10511
rect 48912 10333 48922 10511
rect 48936 10333 48946 10511
rect 48984 10333 48994 10511
rect 50256 10306 50266 10511
rect 48349 10296 50266 10306
rect 22200 10234 22210 10247
rect 48360 10258 48370 10296
rect 45997 10248 48370 10258
rect 20280 10224 22210 10234
rect 24744 10224 29447 10234
rect 22032 10200 22127 10210
rect 22032 10186 22042 10200
rect 20256 10176 22042 10186
rect 21456 9874 21466 10151
rect 21720 9901 21730 10151
rect 24744 9949 24754 10224
rect 29485 10224 35567 10234
rect 35605 10224 41543 10234
rect 41581 10224 41687 10234
rect 48408 10234 48418 10271
rect 48456 10237 48466 10271
rect 42253 10224 48418 10234
rect 48504 10210 48514 10271
rect 48792 10261 48802 10271
rect 28128 10200 48514 10210
rect 48524 10251 48802 10261
rect 28128 9949 28138 10200
rect 28272 10176 29471 10186
rect 28272 9949 28282 10176
rect 31800 10176 35591 10186
rect 31800 10165 31810 10176
rect 38869 10176 41567 10186
rect 45925 10176 48455 10186
rect 48524 10162 48534 10251
rect 35581 10152 48534 10162
rect 29448 10042 29458 10151
rect 31656 10128 48383 10138
rect 31656 10069 31666 10128
rect 48558 10115 48568 10195
rect 47848 10105 48568 10115
rect 31800 10069 31810 10103
rect 38856 10069 38866 10103
rect 41544 10069 41554 10103
rect 41688 10090 41698 10103
rect 48672 10090 48682 10218
rect 41688 10080 48682 10090
rect 48768 10042 48778 10218
rect 29448 10032 48778 10042
rect 31656 9949 31666 10007
rect 31800 9949 31810 10007
rect 38856 9973 38866 10007
rect 41544 9994 41554 10007
rect 41544 9984 47835 9994
rect 48912 9946 48922 10271
rect 38725 9936 48922 9946
rect 48936 9922 48946 10271
rect 48984 10210 48994 10271
rect 24600 9912 48946 9922
rect 21456 9864 21778 9874
rect 21096 9840 21719 9850
rect 21096 9826 21106 9840
rect 21072 9816 21106 9826
rect 21072 9759 21082 9816
rect 21768 9826 21778 9864
rect 24600 9853 24610 9912
rect 45960 9888 46031 9898
rect 24744 9853 24754 9887
rect 28128 9853 28138 9887
rect 28272 9853 28282 9887
rect 31656 9853 31666 9887
rect 31800 9853 31810 9887
rect 38712 9853 38722 9887
rect 38856 9853 38866 9887
rect 42240 9853 42250 9887
rect 45960 9874 45970 9888
rect 45781 9864 45970 9874
rect 42397 9840 46018 9850
rect 21143 9816 21191 9826
rect 21768 9816 45983 9826
rect 21132 9759 21142 9815
rect 21181 9759 21191 9816
rect 24600 9759 24610 9791
rect 24744 9759 24754 9791
rect 24792 9759 24802 9816
rect 28128 9759 28138 9791
rect 28272 9759 28282 9791
rect 28320 9759 28330 9816
rect 31656 9759 31666 9791
rect 31800 9759 31810 9791
rect 31848 9759 31858 9816
rect 38712 9759 38722 9791
rect 38856 9759 38866 9791
rect 38904 9759 38914 9816
rect 42240 9759 42250 9791
rect 42384 9759 42394 9791
rect 42432 9759 42442 9816
rect 45768 9759 45778 9791
rect 45912 9759 45922 9791
rect 45960 9759 45970 9816
rect 46008 9826 46018 9840
rect 49010 9850 49020 10225
rect 46045 9840 49020 9850
rect 49038 9826 49048 10248
rect 46008 9816 49048 9826
<< m2contact >>
rect 21168 39561 21182 39575
rect 21118 39522 21132 39536
rect 20279 38807 20293 38821
rect 20279 38755 20293 38769
rect 20279 34823 20293 34837
rect 20255 34774 20269 34788
rect 20255 34703 20269 34717
rect 20279 34703 20293 34717
rect 24545 39743 24559 39757
rect 28070 39742 28084 39756
rect 28103 39719 28117 39733
rect 28185 39742 28199 39756
rect 31546 39740 31560 39754
rect 31631 39743 31645 39757
rect 31775 39743 31789 39757
rect 38687 39743 38701 39757
rect 38831 39743 38845 39757
rect 42215 39743 42229 39757
rect 42359 39743 42373 39757
rect 45743 39743 45757 39757
rect 45887 39743 45901 39757
rect 21503 39695 21517 39709
rect 31631 39695 31645 39709
rect 28103 39671 28117 39685
rect 31775 39672 31789 39686
rect 21479 39647 21493 39661
rect 21479 39599 21493 39613
rect 21503 39599 21517 39613
rect 21431 39311 21445 39325
rect 21479 39287 21493 39301
rect 38687 39671 38701 39685
rect 38831 39671 38845 39685
rect 31808 39649 31822 39663
rect 45887 39647 45901 39661
rect 46725 39597 46739 39611
rect 21600 39562 21614 39576
rect 24545 39564 24559 39578
rect 31775 39575 31789 39589
rect 31775 39527 31789 39541
rect 45743 39527 45757 39541
rect 46961 39527 46975 39541
rect 47207 39523 47221 39537
rect 38855 39503 38869 39517
rect 47183 39503 47197 39517
rect 47231 39479 47245 39493
rect 27887 39455 27901 39469
rect 31775 39455 31789 39469
rect 38663 39455 38677 39469
rect 39023 39455 39037 39469
rect 46991 39455 47005 39469
rect 21455 39239 21469 39253
rect 20255 30767 20269 30781
rect 20279 30767 20293 30781
rect 20303 30767 20317 30781
rect 21215 30767 21229 30781
rect 47279 39431 47293 39445
rect 47303 39431 47317 39445
rect 47135 39407 47149 39421
rect 47063 39383 47077 39397
rect 47327 39394 47341 39408
rect 26855 39359 26869 39373
rect 36143 39359 36157 39373
rect 36863 39359 36877 39373
rect 47255 39359 47269 39373
rect 47015 39335 47029 39349
rect 26855 39311 26869 39325
rect 27887 39311 27901 39325
rect 31775 39311 31789 39325
rect 47303 39311 47317 39325
rect 47399 39311 47413 39325
rect 47087 39287 47101 39301
rect 47111 39287 47125 39301
rect 26663 39263 26677 39277
rect 26855 39263 26869 39277
rect 27887 39263 27901 39277
rect 31775 39263 31789 39277
rect 35879 39263 35893 39277
rect 38927 39263 38941 39277
rect 42359 39263 42373 39277
rect 45743 39263 45757 39277
rect 45767 39263 45781 39277
rect 47423 39274 47437 39288
rect 47159 39239 47173 39253
rect 47303 39239 47317 39253
rect 47447 39247 47461 39261
rect 26663 39215 26677 39229
rect 26855 39215 26869 39229
rect 27887 39215 27901 39229
rect 31775 39215 31789 39229
rect 42215 39191 42229 39205
rect 46961 39191 46975 39205
rect 21431 39143 21445 39157
rect 21455 39143 21469 39157
rect 21479 39143 21493 39157
rect 22127 39143 22141 39157
rect 25463 39143 25477 39157
rect 25703 39143 25717 39157
rect 26663 39143 26677 39157
rect 26855 39143 26869 39157
rect 27887 39143 27901 39157
rect 46991 39143 47005 39157
rect 47015 39143 47029 39157
rect 47063 39143 47077 39157
rect 47087 39143 47101 39157
rect 47111 39143 47125 39157
rect 47135 39143 47149 39157
rect 47159 39143 47173 39157
rect 47183 39143 47197 39157
rect 47207 39143 47221 39157
rect 47231 39143 47245 39157
rect 47255 39143 47269 39157
rect 47279 39143 47293 39157
rect 47303 39143 47317 39157
rect 47327 39143 47341 39157
rect 21215 30719 21229 30733
rect 20303 30694 20317 30708
rect 20255 30671 20269 30685
rect 20279 30671 20293 30685
rect 20279 26929 20293 26943
rect 20279 26857 20293 26871
rect 21215 26905 21229 26919
rect 21215 26857 21229 26871
rect 21431 19655 21445 19669
rect 21455 19655 21469 19669
rect 20303 19631 20317 19645
rect 21215 19631 21229 19645
rect 21383 19631 21397 19645
rect 47399 39191 47413 39205
rect 47423 39191 47437 39205
rect 47447 39191 47461 39205
rect 46991 36455 47005 36469
rect 47015 36455 47029 36469
rect 47063 36455 47077 36469
rect 47087 36455 47101 36469
rect 47111 36455 47125 36469
rect 47135 36455 47149 36469
rect 47159 36455 47173 36469
rect 47183 36455 47197 36469
rect 47207 36455 47221 36469
rect 47231 36455 47245 36469
rect 47255 36455 47269 36469
rect 47279 36455 47293 36469
rect 47303 36455 47317 36469
rect 47327 36455 47341 36469
rect 47351 36455 47365 36469
rect 47375 36455 47389 36469
rect 47399 36455 47413 36469
rect 47423 36455 47437 36469
rect 47447 36455 47461 36469
rect 50255 38999 50269 39013
rect 50255 38951 50269 38965
rect 50231 38879 50245 38893
rect 47447 36407 47461 36421
rect 46991 36335 47005 36349
rect 47015 36335 47029 36349
rect 47063 36335 47077 36349
rect 47087 36335 47101 36349
rect 47111 36335 47125 36349
rect 47135 36335 47149 36349
rect 47159 36335 47173 36349
rect 47183 36335 47197 36349
rect 47207 36335 47221 36349
rect 47231 36335 47245 36349
rect 47255 36335 47269 36349
rect 47279 36335 47293 36349
rect 47303 36335 47317 36349
rect 47327 36335 47341 36349
rect 47351 36335 47365 36349
rect 47375 36335 47389 36349
rect 47399 36335 47413 36349
rect 47423 36335 47437 36349
rect 46991 35351 47005 35365
rect 47015 35351 47029 35365
rect 47063 35351 47077 35365
rect 47087 35351 47101 35365
rect 47111 35351 47125 35365
rect 47135 35351 47149 35365
rect 47159 35351 47173 35365
rect 47183 35351 47197 35365
rect 47207 35351 47221 35365
rect 47231 35351 47245 35365
rect 47255 35351 47269 35365
rect 47279 35351 47293 35365
rect 47303 35351 47317 35365
rect 47327 35351 47341 35365
rect 47351 35351 47365 35365
rect 47375 35351 47389 35365
rect 47399 35351 47413 35365
rect 47399 35303 47413 35317
rect 46991 35231 47005 35245
rect 47015 35231 47029 35245
rect 47063 35231 47077 35245
rect 47087 35231 47101 35245
rect 47111 35231 47125 35245
rect 47135 35231 47149 35245
rect 47159 35231 47173 35245
rect 47183 35231 47197 35245
rect 47207 35231 47221 35245
rect 47231 35231 47245 35245
rect 47255 35231 47269 35245
rect 47279 35231 47293 35245
rect 47303 35231 47317 35245
rect 47327 35231 47341 35245
rect 47351 35231 47365 35245
rect 47375 35231 47389 35245
rect 46991 34223 47005 34237
rect 47015 34223 47029 34237
rect 47063 34223 47077 34237
rect 47087 34223 47101 34237
rect 47111 34223 47125 34237
rect 47135 34223 47149 34237
rect 47159 34223 47173 34237
rect 47183 34223 47197 34237
rect 47207 34223 47221 34237
rect 47231 34223 47245 34237
rect 47255 34223 47269 34237
rect 47279 34223 47293 34237
rect 47303 34223 47317 34237
rect 47327 34223 47341 34237
rect 47351 34223 47365 34237
rect 50231 38831 50245 38845
rect 50231 35015 50245 35029
rect 50255 35015 50269 35029
rect 50207 34991 50221 35005
rect 50231 34967 50245 34981
rect 50207 34943 50221 34957
rect 50255 34919 50269 34933
rect 50183 34847 50197 34861
rect 50207 34847 50221 34861
rect 50231 34847 50245 34861
rect 47351 34175 47365 34189
rect 46991 34103 47005 34117
rect 47015 34103 47029 34117
rect 47063 34103 47077 34117
rect 47087 34103 47101 34117
rect 47111 34103 47125 34117
rect 47135 34103 47149 34117
rect 47159 34103 47173 34117
rect 47183 34103 47197 34117
rect 47207 34103 47221 34117
rect 47231 34103 47245 34117
rect 47255 34103 47269 34117
rect 47279 34103 47293 34117
rect 47303 34103 47317 34117
rect 47327 34103 47341 34117
rect 46991 33119 47005 33133
rect 47015 33119 47029 33133
rect 47063 33119 47077 33133
rect 47087 33119 47101 33133
rect 47111 33119 47125 33133
rect 47135 33119 47149 33133
rect 47159 33119 47173 33133
rect 47183 33119 47197 33133
rect 47207 33119 47221 33133
rect 47231 33119 47245 33133
rect 47255 33119 47269 33133
rect 47279 33119 47293 33133
rect 47303 33119 47317 33133
rect 47303 33071 47317 33085
rect 46991 32999 47005 33013
rect 47015 32999 47029 33013
rect 47063 32999 47077 33013
rect 47087 32999 47101 33013
rect 47111 32999 47125 33013
rect 47135 32999 47149 33013
rect 47159 32999 47173 33013
rect 47183 32999 47197 33013
rect 47207 32999 47221 33013
rect 47231 32999 47245 33013
rect 47255 32999 47269 33013
rect 47279 32999 47293 33013
rect 46991 32015 47005 32029
rect 47015 32015 47029 32029
rect 47063 32015 47077 32029
rect 47087 32015 47101 32029
rect 47111 32015 47125 32029
rect 47135 32015 47149 32029
rect 47159 32015 47173 32029
rect 47183 32015 47197 32029
rect 47207 32015 47221 32029
rect 47231 32015 47245 32029
rect 47255 32015 47269 32029
rect 47279 32015 47293 32029
rect 50183 34799 50197 34813
rect 50207 34799 50221 34813
rect 50231 34799 50245 34813
rect 46991 31895 47005 31909
rect 47015 31895 47029 31909
rect 47063 31895 47077 31909
rect 47087 31895 47101 31909
rect 47111 31895 47125 31909
rect 47135 31895 47149 31909
rect 47159 31895 47173 31909
rect 47183 31895 47197 31909
rect 47207 31895 47221 31909
rect 47231 31895 47245 31909
rect 47255 31895 47269 31909
rect 47279 31895 47293 31909
rect 50231 30983 50245 30997
rect 50255 30983 50269 30997
rect 46991 30887 47005 30901
rect 47015 30887 47029 30901
rect 47063 30887 47077 30901
rect 47087 30887 47101 30901
rect 47111 30887 47125 30901
rect 47135 30887 47149 30901
rect 47159 30887 47173 30901
rect 47183 30887 47197 30901
rect 47207 30887 47221 30901
rect 47231 30887 47245 30901
rect 47255 30887 47269 30901
rect 47279 30887 47293 30901
rect 50255 30935 50269 30949
rect 50231 30911 50245 30925
rect 46991 30791 47005 30805
rect 47015 30791 47029 30805
rect 47063 30791 47077 30805
rect 47087 30791 47101 30805
rect 47111 30791 47125 30805
rect 47135 30791 47149 30805
rect 47159 30791 47173 30805
rect 47183 30791 47197 30805
rect 47207 30791 47221 30805
rect 47231 30791 47245 30805
rect 47255 30791 47269 30805
rect 47279 30791 47293 30805
rect 50255 30791 50269 30805
rect 46991 29783 47005 29797
rect 47015 29783 47029 29797
rect 47063 29783 47077 29797
rect 47087 29783 47101 29797
rect 47111 29783 47125 29797
rect 47135 29783 47149 29797
rect 47159 29783 47173 29797
rect 47183 29783 47197 29797
rect 47207 29783 47221 29797
rect 47231 29783 47245 29797
rect 47255 29783 47269 29797
rect 47279 29783 47293 29797
rect 50255 30743 50269 30757
rect 46991 29663 47005 29677
rect 47015 29663 47029 29677
rect 47063 29663 47077 29677
rect 47087 29663 47101 29677
rect 47111 29663 47125 29677
rect 47135 29663 47149 29677
rect 47159 29663 47173 29677
rect 47183 29663 47197 29677
rect 47207 29663 47221 29677
rect 47231 29663 47245 29677
rect 47255 29663 47269 29677
rect 47279 29663 47293 29677
rect 46991 28679 47005 28693
rect 47015 28679 47029 28693
rect 47063 28679 47077 28693
rect 47087 28679 47101 28693
rect 47111 28679 47125 28693
rect 47135 28679 47149 28693
rect 47159 28679 47173 28693
rect 47183 28679 47197 28693
rect 47231 28703 47245 28717
rect 47255 28703 47269 28717
rect 47279 28703 47293 28717
rect 47063 28631 47077 28645
rect 47207 28631 47221 28645
rect 47303 28631 47317 28645
rect 46991 28559 47005 28573
rect 47015 28559 47029 28573
rect 46991 27551 47005 27565
rect 47015 27551 47029 27565
rect 47087 28583 47101 28597
rect 47111 28583 47125 28597
rect 47135 28583 47149 28597
rect 47159 28583 47173 28597
rect 47183 28583 47197 28597
rect 47207 28583 47221 28597
rect 47231 28583 47245 28597
rect 47255 28583 47269 28597
rect 47279 28583 47293 28597
rect 47303 28583 47317 28597
rect 47087 27575 47101 27589
rect 47111 27575 47125 27589
rect 47135 27575 47149 27589
rect 47159 27575 47173 27589
rect 47183 27575 47197 27589
rect 47207 27575 47221 27589
rect 47231 27575 47245 27589
rect 47255 27575 47269 27589
rect 47279 27575 47293 27589
rect 47303 27575 47317 27589
rect 47327 27575 47341 27589
rect 47063 27527 47077 27541
rect 47351 27527 47365 27541
rect 46991 27455 47005 27469
rect 47015 27455 47029 27469
rect 47063 27479 47077 27493
rect 47087 27479 47101 27493
rect 47111 27479 47125 27493
rect 47135 27479 47149 27493
rect 47159 27479 47173 27493
rect 47183 27479 47197 27493
rect 47207 27479 47221 27493
rect 47231 27479 47245 27493
rect 47255 27479 47269 27493
rect 47279 27479 47293 27493
rect 47303 27479 47317 27493
rect 47327 27479 47341 27493
rect 47351 27479 47365 27493
rect 46991 26447 47005 26461
rect 47015 26447 47029 26461
rect 47039 26447 47053 26461
rect 47063 26447 47077 26461
rect 47087 26447 47101 26461
rect 47135 26471 47149 26485
rect 47159 26471 47173 26485
rect 47183 26471 47197 26485
rect 47207 26471 47221 26485
rect 47231 26471 47245 26485
rect 47255 26471 47269 26485
rect 47279 26471 47293 26485
rect 47303 26471 47317 26485
rect 47327 26471 47341 26485
rect 47351 26471 47365 26485
rect 47015 26399 47029 26413
rect 47111 26399 47125 26413
rect 47375 26399 47389 26413
rect 46991 26327 47005 26341
rect 47039 26351 47053 26365
rect 47063 26351 47077 26365
rect 47087 26351 47101 26365
rect 47111 26351 47125 26365
rect 47135 26351 47149 26365
rect 47159 26351 47173 26365
rect 47183 26351 47197 26365
rect 47207 26351 47221 26365
rect 47231 26351 47245 26365
rect 47255 26351 47269 26365
rect 47279 26351 47293 26365
rect 47303 26351 47317 26365
rect 47327 26351 47341 26365
rect 47351 26351 47365 26365
rect 47375 26351 47389 26365
rect 46991 25343 47005 25357
rect 47015 25343 47029 25357
rect 47039 25343 47053 25357
rect 47063 25343 47077 25357
rect 47087 25343 47101 25357
rect 47111 25343 47125 25357
rect 47135 25343 47149 25357
rect 47159 25343 47173 25357
rect 47207 25367 47221 25381
rect 47231 25367 47245 25381
rect 47255 25367 47269 25381
rect 47279 25367 47293 25381
rect 47303 25367 47317 25381
rect 47327 25367 47341 25381
rect 47351 25367 47365 25381
rect 47375 25367 47389 25381
rect 47399 25367 47413 25381
rect 47087 25295 47101 25309
rect 47183 25295 47197 25309
rect 47423 25295 47437 25309
rect 46991 25223 47005 25237
rect 47015 25223 47029 25237
rect 47039 25223 47053 25237
rect 47063 25223 47077 25237
rect 47111 25247 47125 25261
rect 47135 25247 47149 25261
rect 47159 25247 47173 25261
rect 47183 25247 47197 25261
rect 47207 25247 47221 25261
rect 47231 25247 47245 25261
rect 47255 25247 47269 25261
rect 47279 25247 47293 25261
rect 47303 25247 47317 25261
rect 47327 25247 47341 25261
rect 47351 25247 47365 25261
rect 47375 25247 47389 25261
rect 47399 25247 47413 25261
rect 47423 25247 47437 25261
rect 47015 24263 47029 24277
rect 47039 24263 47053 24277
rect 47063 24263 47077 24277
rect 47087 24263 47101 24277
rect 47111 24263 47125 24277
rect 47135 24263 47149 24277
rect 47159 24263 47173 24277
rect 47183 24263 47197 24277
rect 47207 24263 47221 24277
rect 47231 24263 47245 24277
rect 47255 24263 47269 24277
rect 47279 24263 47293 24277
rect 47303 24263 47317 24277
rect 47327 24263 47341 24277
rect 47351 24263 47365 24277
rect 47375 24263 47389 24277
rect 47399 24263 47413 24277
rect 47423 24263 47437 24277
rect 47447 24263 47461 24277
rect 47015 24215 47029 24229
rect 47039 24215 47053 24229
rect 47063 24215 47077 24229
rect 47087 24215 47101 24229
rect 47111 24215 47125 24229
rect 47135 24215 47149 24229
rect 47159 24215 47173 24229
rect 46991 24167 47005 24181
rect 47015 24167 47029 24181
rect 47039 24167 47053 24181
rect 47063 24167 47077 24181
rect 47087 24167 47101 24181
rect 47111 24167 47125 24181
rect 47135 24167 47149 24181
rect 47471 24191 47485 24205
rect 46991 24119 47005 24133
rect 47015 24119 47029 24133
rect 47039 24119 47053 24133
rect 47063 24119 47077 24133
rect 47087 24119 47101 24133
rect 47111 24119 47125 24133
rect 47135 24119 47149 24133
rect 46991 23111 47005 23125
rect 47015 23111 47029 23125
rect 47039 23111 47053 23125
rect 47063 23111 47077 23125
rect 47087 23111 47101 23125
rect 47111 23111 47125 23125
rect 47183 24143 47197 24157
rect 47207 24143 47221 24157
rect 47231 24143 47245 24157
rect 47255 24143 47269 24157
rect 47279 24143 47293 24157
rect 47303 24143 47317 24157
rect 47327 24143 47341 24157
rect 47351 24143 47365 24157
rect 47375 24143 47389 24157
rect 47399 24143 47413 24157
rect 47423 24143 47437 24157
rect 47447 24143 47461 24157
rect 47471 24143 47485 24157
rect 47159 23135 47173 23149
rect 47183 23135 47197 23149
rect 47207 23135 47221 23149
rect 47231 23135 47245 23149
rect 47255 23135 47269 23149
rect 47279 23135 47293 23149
rect 47303 23135 47317 23149
rect 47327 23135 47341 23149
rect 47351 23135 47365 23149
rect 47375 23135 47389 23149
rect 47399 23135 47413 23149
rect 47423 23135 47437 23149
rect 47447 23135 47461 23149
rect 47471 23135 47485 23149
rect 47495 23135 47509 23149
rect 47375 23087 47389 23101
rect 47519 23087 47533 23101
rect 47135 23063 47149 23077
rect 46991 23015 47005 23029
rect 47015 23015 47029 23029
rect 47039 23015 47053 23029
rect 47063 23015 47077 23029
rect 47087 23015 47101 23029
rect 47111 23015 47125 23029
rect 47135 23015 47149 23029
rect 47159 23015 47173 23029
rect 47183 23015 47197 23029
rect 47207 23015 47221 23029
rect 47231 23015 47245 23029
rect 47255 23015 47269 23029
rect 47279 23015 47293 23029
rect 47303 23015 47317 23029
rect 47327 23015 47341 23029
rect 47351 23015 47365 23029
rect 46991 22007 47005 22021
rect 47015 22007 47029 22021
rect 47039 22007 47053 22021
rect 47063 22007 47077 22021
rect 47087 22007 47101 22021
rect 47111 22007 47125 22021
rect 47135 22007 47149 22021
rect 47159 22007 47173 22021
rect 47183 22007 47197 22021
rect 47207 22007 47221 22021
rect 47231 22007 47245 22021
rect 47399 23039 47413 23053
rect 47423 23039 47437 23053
rect 47447 23039 47461 23053
rect 47471 23039 47485 23053
rect 47495 23039 47509 23053
rect 47519 23039 47533 23053
rect 47279 22031 47293 22045
rect 47303 22031 47317 22045
rect 47327 22031 47341 22045
rect 47351 22031 47365 22045
rect 47375 22031 47389 22045
rect 47399 22031 47413 22045
rect 47423 22031 47437 22045
rect 47447 22031 47461 22045
rect 47471 22031 47485 22045
rect 47495 22031 47509 22045
rect 47519 22031 47533 22045
rect 47543 22031 47557 22045
rect 47087 21959 47101 21973
rect 47255 21959 47269 21973
rect 47567 21959 47581 21973
rect 46991 21887 47005 21901
rect 47015 21887 47029 21901
rect 47039 21887 47053 21901
rect 47063 21887 47077 21901
rect 47111 21911 47125 21925
rect 47135 21911 47149 21925
rect 47159 21911 47173 21925
rect 47183 21911 47197 21925
rect 47207 21911 47221 21925
rect 47231 21911 47245 21925
rect 47255 21911 47269 21925
rect 47279 21911 47293 21925
rect 47303 21911 47317 21925
rect 47327 21911 47341 21925
rect 47351 21911 47365 21925
rect 47375 21911 47389 21925
rect 47399 21911 47413 21925
rect 47423 21911 47437 21925
rect 47447 21911 47461 21925
rect 47471 21911 47485 21925
rect 47495 21911 47509 21925
rect 47519 21911 47533 21925
rect 47543 21911 47557 21925
rect 47567 21911 47581 21925
rect 46991 20903 47005 20917
rect 47015 20903 47029 20917
rect 47039 20903 47053 20917
rect 47063 20903 47077 20917
rect 47087 20903 47101 20917
rect 47111 20903 47125 20917
rect 47135 20903 47149 20917
rect 47159 20903 47173 20917
rect 47183 20903 47197 20917
rect 47207 20903 47221 20917
rect 47231 20903 47245 20917
rect 47255 20903 47269 20917
rect 47279 20903 47293 20917
rect 47303 20903 47317 20917
rect 47327 20903 47341 20917
rect 47351 20903 47365 20917
rect 47375 20903 47389 20917
rect 47399 20903 47413 20917
rect 47423 20903 47437 20917
rect 47447 20903 47461 20917
rect 47471 20903 47485 20917
rect 47495 20903 47509 20917
rect 47519 20903 47533 20917
rect 47567 20927 47581 20941
rect 47591 20927 47605 20941
rect 46991 20855 47005 20869
rect 47543 20855 47557 20869
rect 47615 20855 47629 20869
rect 47015 20807 47029 20821
rect 47039 20807 47053 20821
rect 47063 20807 47077 20821
rect 47087 20807 47101 20821
rect 47111 20807 47125 20821
rect 47135 20807 47149 20821
rect 47159 20807 47173 20821
rect 47183 20807 47197 20821
rect 47207 20807 47221 20821
rect 47231 20807 47245 20821
rect 47255 20807 47269 20821
rect 47279 20807 47293 20821
rect 47303 20807 47317 20821
rect 47327 20807 47341 20821
rect 47351 20807 47365 20821
rect 47375 20807 47389 20821
rect 47399 20807 47413 20821
rect 47423 20807 47437 20821
rect 47447 20807 47461 20821
rect 47471 20807 47485 20821
rect 47495 20807 47509 20821
rect 47519 20807 47533 20821
rect 47543 20807 47557 20821
rect 47567 20807 47581 20821
rect 47591 20807 47605 20821
rect 47615 20807 47629 20821
rect 46991 19775 47005 19789
rect 47015 19775 47029 19789
rect 47039 19775 47053 19789
rect 47063 19775 47077 19789
rect 47087 19775 47101 19789
rect 47135 19799 47149 19813
rect 47159 19799 47173 19813
rect 47183 19799 47197 19813
rect 47207 19799 47221 19813
rect 47231 19799 47245 19813
rect 47255 19799 47269 19813
rect 47279 19799 47293 19813
rect 47303 19799 47317 19813
rect 47327 19799 47341 19813
rect 47351 19799 47365 19813
rect 47375 19799 47389 19813
rect 47399 19799 47413 19813
rect 47423 19799 47437 19813
rect 47447 19799 47461 19813
rect 47471 19799 47485 19813
rect 47495 19799 47509 19813
rect 47519 19799 47533 19813
rect 47543 19799 47557 19813
rect 47567 19799 47581 19813
rect 47591 19799 47605 19813
rect 47615 19799 47629 19813
rect 47639 19799 47653 19813
rect 47255 19751 47269 19765
rect 47663 19751 47677 19765
rect 47111 19727 47125 19741
rect 46991 19679 47005 19693
rect 47015 19679 47029 19693
rect 47039 19679 47053 19693
rect 47063 19679 47077 19693
rect 47087 19679 47101 19693
rect 47111 19679 47125 19693
rect 47135 19679 47149 19693
rect 47159 19679 47173 19693
rect 47183 19679 47197 19693
rect 47207 19679 47221 19693
rect 47231 19679 47245 19693
rect 20303 19583 20317 19597
rect 21215 19583 21229 19597
rect 21383 19583 21397 19597
rect 21431 19583 21445 19597
rect 21455 19583 21469 19597
rect 20255 18791 20269 18805
rect 20255 18743 20269 18757
rect 21534 19607 21548 19621
rect 21581 19607 21595 19621
rect 23447 19607 23461 19621
rect 27623 19607 27637 19621
rect 37463 19607 37477 19621
rect 45167 19607 45181 19621
rect 45911 19607 45925 19621
rect 46127 19607 46141 19621
rect 46271 19607 46285 19621
rect 46319 19607 46333 19621
rect 46367 19607 46381 19621
rect 46415 19607 46429 19621
rect 46487 19607 46501 19621
rect 21558 19567 21572 19581
rect 21603 19559 21617 19573
rect 21650 19559 21664 19573
rect 27599 19583 27613 19597
rect 37439 19583 37453 19597
rect 24239 19559 24253 19573
rect 26687 19559 26701 19573
rect 26711 19559 26725 19573
rect 37199 19559 37213 19573
rect 37223 19559 37237 19573
rect 21627 19518 21641 19532
rect 21672 19511 21686 19525
rect 27431 19535 27445 19549
rect 27455 19535 27469 19549
rect 21695 19487 21709 19501
rect 24791 19511 24805 19525
rect 26471 19511 26485 19525
rect 26495 19511 26509 19525
rect 37031 19535 37045 19549
rect 25007 19487 25021 19501
rect 26279 19487 26293 19501
rect 26303 19487 26317 19501
rect 25751 19463 25765 19477
rect 25919 19463 25933 19477
rect 26279 19415 26293 19429
rect 26471 19391 26485 19405
rect 26687 19367 26701 19381
rect 27431 19343 27445 19357
rect 21623 18623 21637 18637
rect 21671 18623 21685 18637
rect 21695 18623 21709 18637
rect 25799 18623 25813 18637
rect 27599 19343 27613 19357
rect 21551 18575 21565 18589
rect 27023 18575 27037 18589
rect 27455 18575 27469 18589
rect 21551 18527 21565 18541
rect 21623 18527 21637 18541
rect 21671 18527 21685 18541
rect 27023 18527 27037 18541
rect 27455 18527 27469 18541
rect 21719 18503 21733 18517
rect 22168 18503 22182 18517
rect 24983 18503 24997 18517
rect 20303 18455 20317 18469
rect 21215 18455 21229 18469
rect 21383 18455 21397 18469
rect 21431 18455 21445 18469
rect 21455 18455 21469 18469
rect 21479 18455 21493 18469
rect 21551 18455 21565 18469
rect 21695 18455 21709 18469
rect 22144 18431 22158 18445
rect 24167 18431 24181 18445
rect 25823 18431 25837 18445
rect 27023 18431 27037 18445
rect 27455 18431 27469 18445
rect 20303 18407 20317 18421
rect 21215 18407 21229 18421
rect 21383 18407 21397 18421
rect 21431 18407 21445 18421
rect 21455 18407 21469 18421
rect 21479 18407 21493 18421
rect 21551 18407 21565 18421
rect 37199 19487 37213 19501
rect 37439 19487 37453 19501
rect 44423 18503 44437 18517
rect 45239 18503 45253 18517
rect 43631 18479 43645 18493
rect 46055 18479 46069 18493
rect 43511 18455 43525 18469
rect 45239 18455 45253 18469
rect 45263 18455 45277 18469
rect 31151 18431 31165 18445
rect 32039 18431 32053 18445
rect 33143 18431 33157 18445
rect 33959 18431 33973 18445
rect 33983 18431 33997 18445
rect 34799 18431 34813 18445
rect 36388 18431 36402 18445
rect 36412 18431 36426 18445
rect 37223 18431 37237 18445
rect 38015 18431 38029 18445
rect 39479 18431 39493 18445
rect 40408 18431 40422 18445
rect 40432 18431 40446 18445
rect 41231 18431 41245 18445
rect 42815 18431 42829 18445
rect 44423 18431 44437 18445
rect 44447 18431 44461 18445
rect 43631 18407 43645 18421
rect 47279 19703 47293 19717
rect 47303 19703 47317 19717
rect 47327 19703 47341 19717
rect 47351 19703 47365 19717
rect 47375 19703 47389 19717
rect 47399 19703 47413 19717
rect 47423 19703 47437 19717
rect 47447 19703 47461 19717
rect 47471 19703 47485 19717
rect 47495 19703 47509 19717
rect 47519 19703 47533 19717
rect 47543 19703 47557 19717
rect 47567 19703 47581 19717
rect 47591 19703 47605 19717
rect 47615 19703 47629 19717
rect 47639 19703 47653 19717
rect 47663 19703 47677 19717
rect 48191 19343 48205 19357
rect 48191 19295 48205 19309
rect 48359 19103 48373 19117
rect 48383 19079 48397 19093
rect 48407 19055 48421 19069
rect 48431 19031 48445 19045
rect 48455 19007 48469 19021
rect 48479 18983 48493 18997
rect 48503 18959 48517 18973
rect 48527 18935 48541 18949
rect 48551 18911 48565 18925
rect 48575 18887 48589 18901
rect 48599 18863 48613 18877
rect 48623 18839 48637 18853
rect 48647 18815 48661 18829
rect 48671 18791 48685 18805
rect 50255 18791 50269 18805
rect 48695 18743 48709 18757
rect 50255 18743 50269 18757
rect 48719 18719 48733 18733
rect 48743 18695 48757 18709
rect 48767 18671 48781 18685
rect 48839 18647 48853 18661
rect 50255 18647 50269 18661
rect 48863 18599 48877 18613
rect 50255 18599 50269 18613
rect 48887 18575 48901 18589
rect 48911 18551 48925 18565
rect 48935 18527 48949 18541
rect 48983 18503 48997 18517
rect 50111 18479 50125 18493
rect 50159 18455 50173 18469
rect 50207 18431 50221 18445
rect 21719 18383 21733 18397
rect 29063 18383 29077 18397
rect 29783 18383 29797 18397
rect 30263 18383 30277 18397
rect 43655 18383 43669 18397
rect 46871 18383 46885 18397
rect 48359 18383 48373 18397
rect 48383 18383 48397 18397
rect 48407 18383 48421 18397
rect 48431 18383 48445 18397
rect 48455 18383 48469 18397
rect 48479 18383 48493 18397
rect 48503 18383 48517 18397
rect 48527 18383 48541 18397
rect 48551 18383 48565 18397
rect 48575 18383 48589 18397
rect 48599 18383 48613 18397
rect 48623 18383 48637 18397
rect 48647 18383 48661 18397
rect 48671 18383 48685 18397
rect 48695 18383 48709 18397
rect 48719 18383 48733 18397
rect 48743 18383 48757 18397
rect 48767 18383 48781 18397
rect 21431 18215 21445 18229
rect 21455 18215 21469 18229
rect 21479 18215 21493 18229
rect 21719 18215 21733 18229
rect 21743 18186 21757 18200
rect 21431 18162 21445 18176
rect 21743 18162 21757 18176
rect 48359 18163 48373 18177
rect 48383 18163 48397 18177
rect 48407 18163 48421 18177
rect 48431 18163 48445 18177
rect 48455 18163 48469 18177
rect 21455 18138 21469 18152
rect 21479 18138 21493 18152
rect 21719 18138 21733 18152
rect 48330 18138 48344 18152
rect 48503 18139 48517 18153
rect 48527 18139 48541 18153
rect 48551 18139 48565 18153
rect 48575 18139 48589 18153
rect 20255 14735 20269 14749
rect 20303 14735 20317 14749
rect 21215 14735 21229 14749
rect 21455 14735 21469 14749
rect 21479 14735 21493 14749
rect 48330 18114 48344 18128
rect 48839 18383 48853 18397
rect 48863 18383 48877 18397
rect 48887 18383 48901 18397
rect 48911 18383 48925 18397
rect 48935 18383 48949 18397
rect 48983 18383 48997 18397
rect 50111 18383 50125 18397
rect 50159 18383 50173 18397
rect 50207 18383 50221 18397
rect 48623 18115 48637 18129
rect 48647 18115 48661 18129
rect 48671 18115 48685 18129
rect 48695 18115 48709 18129
rect 48719 18115 48733 18129
rect 48743 18115 48757 18129
rect 48767 18115 48781 18129
rect 48791 18115 48805 18129
rect 48815 18115 48829 18129
rect 48330 18090 48344 18104
rect 48330 18066 48344 18080
rect 48623 18067 48637 18081
rect 48647 18067 48661 18081
rect 48671 18067 48685 18081
rect 48695 18067 48709 18081
rect 48719 18067 48733 18081
rect 48743 18067 48757 18081
rect 48767 18067 48781 18081
rect 48791 18067 48805 18081
rect 48815 18067 48829 18081
rect 48330 18042 48344 18056
rect 48575 18043 48589 18057
rect 48359 18019 48373 18033
rect 48383 18019 48397 18033
rect 48407 18019 48421 18033
rect 48431 18019 48445 18033
rect 48455 18019 48469 18033
rect 48503 18019 48517 18033
rect 48527 18019 48541 18033
rect 48551 18019 48565 18033
rect 20255 14687 20269 14701
rect 20303 14687 20317 14701
rect 21215 14687 21229 14701
rect 21455 14687 21469 14701
rect 21479 14687 21493 14701
rect 20255 10703 20269 10717
rect 20255 10655 20269 10669
rect 48359 14615 48373 14629
rect 48383 14615 48397 14629
rect 48407 14615 48421 14629
rect 48431 14615 48445 14629
rect 48455 14615 48469 14629
rect 48503 14615 48517 14629
rect 48527 14615 48541 14629
rect 48551 14615 48565 14629
rect 48647 14615 48661 14629
rect 48671 14615 48685 14629
rect 48695 14615 48709 14629
rect 48719 14615 48733 14629
rect 48335 14591 48349 14605
rect 48359 14567 48373 14581
rect 48383 14567 48397 14581
rect 48407 14567 48421 14581
rect 48431 14567 48445 14581
rect 48455 14567 48469 14581
rect 48503 14567 48517 14581
rect 48527 14567 48541 14581
rect 48551 14567 48565 14581
rect 48647 14567 48661 14581
rect 48671 14567 48685 14581
rect 48695 14567 48709 14581
rect 48719 14567 48733 14581
rect 21455 13993 21469 14007
rect 21479 13993 21493 14007
rect 21743 13969 21757 13983
rect 21455 13943 21469 13957
rect 21479 13943 21493 13957
rect 21743 13945 21757 13959
rect 48359 13199 48373 13213
rect 48383 13199 48397 13213
rect 48407 13199 48421 13213
rect 48431 13199 48445 13213
rect 48455 13199 48469 13213
rect 48503 13199 48517 13213
rect 48527 13199 48541 13213
rect 48335 13175 48349 13189
rect 48359 13151 48373 13165
rect 48383 13151 48397 13165
rect 48407 13151 48421 13165
rect 48431 13151 48445 13165
rect 48455 13151 48469 13165
rect 48503 13151 48517 13165
rect 48527 13151 48541 13165
rect 48359 12935 48373 12949
rect 48383 12935 48397 12949
rect 48407 12935 48421 12949
rect 48431 12935 48445 12949
rect 48455 12935 48469 12949
rect 48503 12935 48517 12949
rect 48527 12935 48541 12949
rect 48335 12911 48349 12925
rect 48359 12887 48373 12901
rect 48383 12887 48397 12901
rect 48407 12887 48421 12901
rect 48431 12887 48445 12901
rect 48455 12887 48469 12901
rect 48503 12887 48517 12901
rect 48527 12887 48541 12901
rect 48359 12599 48373 12613
rect 48383 12599 48397 12613
rect 48407 12599 48421 12613
rect 48431 12599 48445 12613
rect 48455 12599 48469 12613
rect 48503 12599 48517 12613
rect 48335 12575 48349 12589
rect 48359 12551 48373 12565
rect 48383 12551 48397 12565
rect 48407 12551 48421 12565
rect 48431 12551 48445 12565
rect 48455 12551 48469 12565
rect 48503 12551 48517 12565
rect 48359 10799 48373 10813
rect 48383 10799 48397 10813
rect 48407 10799 48421 10813
rect 48431 10799 48445 10813
rect 48455 10799 48469 10813
rect 48503 10799 48517 10813
rect 48671 10799 48685 10813
rect 48695 10799 48709 10813
rect 48335 10775 48349 10789
rect 48359 10751 48373 10765
rect 48383 10751 48397 10765
rect 48407 10751 48421 10765
rect 48431 10751 48445 10765
rect 48455 10751 48469 10765
rect 48503 10751 48517 10765
rect 48671 10751 48685 10765
rect 48695 10751 48709 10765
rect 50207 14759 50221 14773
rect 50207 14711 50221 14725
rect 50207 14615 50221 14629
rect 50207 14567 50221 14581
rect 48863 10751 48877 10765
rect 48887 10751 48901 10765
rect 48911 10751 48925 10765
rect 48935 10751 48949 10765
rect 48983 10751 48997 10765
rect 50207 10751 50221 10765
rect 48863 10703 48877 10717
rect 48887 10703 48901 10717
rect 48911 10703 48925 10717
rect 48935 10703 48949 10717
rect 48983 10703 48997 10717
rect 50207 10703 50221 10717
rect 50255 10703 50269 10717
rect 50255 10655 50269 10669
rect 48383 10559 48397 10573
rect 48407 10559 48421 10573
rect 48431 10559 48445 10573
rect 48455 10559 48469 10573
rect 48503 10559 48517 10573
rect 48671 10559 48685 10573
rect 48695 10559 48709 10573
rect 48767 10559 48781 10573
rect 48791 10559 48805 10573
rect 48863 10559 48877 10573
rect 48887 10559 48901 10573
rect 48911 10559 48925 10573
rect 48935 10559 48949 10573
rect 48983 10559 48997 10573
rect 50255 10559 50269 10573
rect 48383 10511 48397 10525
rect 48407 10511 48421 10525
rect 48431 10511 48445 10525
rect 48455 10511 48469 10525
rect 48503 10511 48517 10525
rect 48671 10511 48685 10525
rect 48695 10511 48709 10525
rect 48767 10511 48781 10525
rect 48791 10511 48805 10525
rect 48863 10511 48877 10525
rect 48887 10511 48901 10525
rect 48911 10511 48925 10525
rect 48935 10511 48949 10525
rect 48983 10511 48997 10525
rect 50255 10511 50269 10525
rect 21455 10376 21469 10390
rect 48383 10377 48397 10391
rect 48407 10377 48421 10391
rect 48431 10377 48445 10391
rect 48455 10377 48469 10391
rect 48503 10377 48517 10391
rect 48671 10377 48685 10391
rect 21743 10352 21757 10366
rect 48335 10352 48349 10366
rect 21743 10328 21757 10342
rect 48335 10328 48349 10342
rect 48431 10328 48445 10342
rect 48767 10319 48781 10333
rect 48791 10319 48805 10333
rect 48863 10319 48877 10333
rect 48887 10319 48901 10333
rect 48911 10319 48925 10333
rect 48935 10319 48949 10333
rect 48983 10319 48997 10333
rect 48335 10295 48349 10309
rect 21719 10247 21733 10261
rect 22199 10247 22213 10261
rect 45983 10246 45997 10260
rect 48407 10271 48421 10285
rect 48455 10271 48469 10285
rect 48503 10271 48517 10285
rect 48791 10271 48805 10285
rect 48911 10271 48925 10285
rect 48935 10271 48949 10285
rect 48983 10271 48997 10285
rect 22127 10199 22141 10213
rect 21455 10151 21469 10165
rect 21719 10151 21733 10165
rect 29447 10223 29461 10237
rect 29471 10223 29485 10237
rect 35567 10223 35581 10237
rect 35591 10223 35605 10237
rect 41543 10223 41557 10237
rect 41567 10223 41581 10237
rect 41687 10223 41701 10237
rect 42239 10223 42253 10237
rect 48455 10223 48469 10237
rect 29471 10175 29485 10189
rect 35591 10175 35605 10189
rect 38855 10175 38869 10189
rect 41567 10175 41581 10189
rect 45911 10175 45925 10189
rect 48455 10175 48469 10189
rect 29447 10151 29461 10165
rect 31799 10151 31813 10165
rect 35567 10151 35581 10165
rect 48671 10218 48685 10232
rect 48767 10218 48781 10232
rect 48554 10195 48568 10209
rect 48383 10127 48397 10141
rect 31799 10103 31813 10117
rect 38855 10103 38869 10117
rect 41543 10103 41557 10117
rect 41687 10103 41701 10117
rect 47834 10103 47848 10117
rect 31655 10055 31669 10069
rect 31799 10055 31813 10069
rect 38855 10055 38869 10069
rect 41543 10055 41557 10069
rect 31655 10007 31669 10021
rect 31799 10007 31813 10021
rect 38855 10007 38869 10021
rect 41543 10007 41557 10021
rect 47835 9984 47849 9998
rect 38855 9959 38869 9973
rect 24743 9935 24757 9949
rect 28127 9935 28141 9949
rect 28271 9935 28285 9949
rect 31655 9935 31669 9949
rect 31799 9935 31813 9949
rect 38711 9935 38725 9949
rect 49038 10248 49052 10262
rect 49010 10225 49024 10239
rect 48982 10196 48996 10210
rect 21719 9887 21733 9901
rect 21719 9839 21733 9853
rect 21129 9815 21143 9829
rect 24743 9887 24757 9901
rect 28127 9887 28141 9901
rect 28271 9887 28285 9901
rect 31655 9887 31669 9901
rect 31799 9887 31813 9901
rect 38711 9887 38725 9901
rect 38855 9887 38869 9901
rect 42239 9887 42253 9901
rect 45767 9863 45781 9877
rect 46031 9887 46045 9901
rect 24599 9839 24613 9853
rect 24743 9839 24757 9853
rect 28127 9839 28141 9853
rect 28271 9839 28285 9853
rect 31655 9839 31669 9853
rect 31799 9839 31813 9853
rect 38711 9839 38725 9853
rect 38855 9839 38869 9853
rect 42239 9839 42253 9853
rect 42383 9839 42397 9853
rect 24599 9791 24613 9805
rect 24743 9791 24757 9805
rect 28127 9791 28141 9805
rect 28271 9791 28285 9805
rect 31655 9791 31669 9805
rect 31799 9791 31813 9805
rect 38711 9791 38725 9805
rect 38855 9791 38869 9805
rect 42239 9791 42253 9805
rect 42383 9791 42397 9805
rect 45767 9791 45781 9805
rect 45911 9791 45925 9805
rect 45983 9815 45997 9829
rect 46031 9839 46045 9853
<< metal2 >>
rect 24559 39743 28070 39755
rect 21480 39613 21492 39647
rect 21504 39613 21516 39695
rect 24547 39578 24559 39743
rect 28084 39743 28185 39755
rect 28104 39685 28116 39719
rect 31546 39682 31558 39740
rect 31632 39709 31644 39743
rect 31776 39686 31788 39743
rect 31546 39670 31705 39682
rect 38688 39685 38700 39743
rect 38832 39685 38844 39743
rect 31693 39662 31705 39670
rect 31693 39650 31808 39662
rect 21182 39563 21600 39575
rect 20850 39536 22105 39547
rect 31776 39541 31788 39575
rect 20850 39522 21118 39536
rect 21132 39522 22105 39536
rect 20850 39347 22105 39522
rect 20280 38769 20292 38807
rect 20256 34717 20268 34774
rect 20280 34717 20292 34823
rect 20256 30685 20268 30767
rect 20280 30685 20292 30767
rect 20304 30708 20316 30767
rect 20850 27366 21050 39347
rect 21432 39157 21444 39311
rect 21456 39157 21468 39239
rect 21480 39157 21492 39287
rect 21905 39133 22105 39347
rect 26856 39325 26868 39359
rect 27888 39325 27900 39455
rect 31776 39325 31788 39455
rect 26664 39229 26676 39263
rect 26856 39229 26868 39263
rect 27888 39229 27900 39263
rect 31776 39229 31788 39263
rect 22121 39143 22127 39157
rect 25457 39143 25463 39157
rect 25697 39143 25703 39157
rect 26657 39143 26663 39157
rect 26849 39143 26855 39157
rect 27883 39143 27887 39157
rect 35880 39156 35892 39263
rect 36144 39156 36156 39359
rect 36864 39156 36876 39359
rect 38664 39156 38676 39455
rect 38856 39156 38868 39503
rect 38928 39156 38940 39263
rect 39024 39156 39036 39455
rect 42216 39205 42228 39743
rect 42360 39277 42372 39743
rect 45744 39588 45756 39743
rect 45888 39661 45900 39743
rect 46721 39611 47826 39764
rect 46721 39597 46725 39611
rect 46739 39597 47826 39611
rect 45744 39576 45780 39588
rect 45744 39277 45756 39527
rect 45768 39277 45780 39576
rect 46721 39564 47826 39597
rect 35874 39144 35892 39156
rect 36138 39144 36156 39156
rect 36858 39144 36876 39156
rect 38657 39144 38676 39156
rect 38849 39144 38868 39156
rect 38921 39144 38940 39156
rect 39017 39144 39036 39156
rect 22121 39133 22133 39143
rect 25457 39133 25469 39143
rect 25697 39133 25709 39143
rect 26657 39133 26669 39143
rect 26849 39133 26861 39143
rect 27883 39133 27895 39143
rect 35874 39133 35886 39144
rect 36138 39133 36150 39144
rect 36858 39133 36870 39144
rect 38657 39133 38669 39144
rect 38849 39133 38861 39144
rect 38921 39133 38933 39144
rect 39017 39133 39029 39144
rect 46721 39133 46921 39564
rect 46962 39205 46974 39527
rect 46992 39157 47004 39455
rect 47016 39157 47028 39335
rect 47064 39157 47076 39383
rect 47088 39157 47100 39287
rect 47112 39157 47124 39287
rect 47136 39157 47148 39407
rect 47160 39157 47172 39239
rect 47184 39157 47196 39503
rect 47208 39157 47220 39523
rect 47232 39157 47244 39479
rect 47256 39157 47268 39359
rect 47280 39157 47292 39431
rect 47304 39325 47316 39431
rect 47304 39157 47316 39239
rect 47328 39157 47340 39394
rect 47400 39205 47412 39311
rect 47424 39205 47436 39274
rect 47448 39205 47460 39247
rect 46992 36349 47004 36455
rect 47016 36349 47028 36455
rect 47064 36349 47076 36455
rect 47088 36349 47100 36455
rect 47112 36349 47124 36455
rect 47136 36349 47148 36455
rect 47160 36349 47172 36455
rect 47184 36349 47196 36455
rect 47208 36349 47220 36455
rect 47232 36349 47244 36455
rect 47256 36349 47268 36455
rect 47280 36349 47292 36455
rect 47304 36349 47316 36455
rect 47328 36349 47340 36455
rect 47352 36349 47364 36455
rect 47376 36349 47388 36455
rect 47400 36349 47412 36455
rect 47424 36349 47436 36455
rect 47448 36421 47460 36455
rect 46992 35245 47004 35351
rect 47016 35245 47028 35351
rect 47064 35245 47076 35351
rect 47088 35245 47100 35351
rect 47112 35245 47124 35351
rect 47136 35245 47148 35351
rect 47160 35245 47172 35351
rect 47184 35245 47196 35351
rect 47208 35245 47220 35351
rect 47232 35245 47244 35351
rect 47256 35245 47268 35351
rect 47280 35245 47292 35351
rect 47304 35245 47316 35351
rect 47328 35245 47340 35351
rect 47352 35245 47364 35351
rect 47376 35245 47388 35351
rect 47400 35317 47412 35351
rect 46992 34117 47004 34223
rect 47016 34117 47028 34223
rect 47064 34117 47076 34223
rect 47088 34117 47100 34223
rect 47112 34117 47124 34223
rect 47136 34117 47148 34223
rect 47160 34117 47172 34223
rect 47184 34117 47196 34223
rect 47208 34117 47220 34223
rect 47232 34117 47244 34223
rect 47256 34117 47268 34223
rect 47280 34117 47292 34223
rect 47304 34117 47316 34223
rect 47328 34117 47340 34223
rect 47352 34189 47364 34223
rect 46992 33013 47004 33119
rect 47016 33013 47028 33119
rect 47064 33013 47076 33119
rect 47088 33013 47100 33119
rect 47112 33013 47124 33119
rect 47136 33013 47148 33119
rect 47160 33013 47172 33119
rect 47184 33013 47196 33119
rect 47208 33013 47220 33119
rect 47232 33013 47244 33119
rect 47256 33013 47268 33119
rect 47280 33013 47292 33119
rect 47304 33085 47316 33119
rect 46992 31909 47004 32015
rect 47016 31909 47028 32015
rect 47064 31909 47076 32015
rect 47088 31909 47100 32015
rect 47112 31909 47124 32015
rect 47136 31909 47148 32015
rect 47160 31909 47172 32015
rect 47184 31909 47196 32015
rect 47208 31909 47220 32015
rect 47232 31909 47244 32015
rect 47256 31909 47268 32015
rect 47280 31909 47292 32015
rect 46992 30805 47004 30887
rect 47016 30805 47028 30887
rect 47064 30805 47076 30887
rect 47088 30805 47100 30887
rect 47112 30805 47124 30887
rect 47136 30805 47148 30887
rect 47160 30805 47172 30887
rect 47184 30805 47196 30887
rect 47208 30805 47220 30887
rect 47232 30805 47244 30887
rect 47256 30805 47268 30887
rect 47280 30805 47292 30887
rect 21216 30733 21228 30767
rect 46992 29677 47004 29783
rect 47016 29677 47028 29783
rect 47064 29677 47076 29783
rect 47088 29677 47100 29783
rect 47112 29677 47124 29783
rect 47136 29677 47148 29783
rect 47160 29677 47172 29783
rect 47184 29677 47196 29783
rect 47208 29677 47220 29783
rect 47232 29677 47244 29783
rect 47256 29677 47268 29783
rect 47280 29677 47292 29783
rect 46992 28573 47004 28679
rect 47016 28573 47028 28679
rect 47064 28645 47076 28679
rect 47088 28597 47100 28679
rect 47112 28597 47124 28679
rect 47136 28597 47148 28679
rect 47160 28597 47172 28679
rect 47184 28597 47196 28679
rect 47208 28597 47220 28631
rect 47232 28597 47244 28703
rect 47256 28597 47268 28703
rect 47280 28597 47292 28703
rect 47304 28597 47316 28631
rect 46992 27469 47004 27551
rect 47016 27469 47028 27551
rect 47064 27493 47076 27527
rect 47088 27493 47100 27575
rect 47112 27493 47124 27575
rect 47136 27493 47148 27575
rect 47160 27493 47172 27575
rect 47184 27493 47196 27575
rect 47208 27493 47220 27575
rect 47232 27493 47244 27575
rect 47256 27493 47268 27575
rect 47280 27493 47292 27575
rect 47304 27493 47316 27575
rect 47328 27493 47340 27575
rect 47352 27493 47364 27527
rect 20207 27166 21050 27366
rect 47626 27373 47826 39564
rect 50256 38965 50268 38999
rect 50232 38845 50244 38879
rect 50208 34957 50220 34991
rect 50232 34981 50244 35015
rect 50256 34933 50268 35015
rect 50184 34813 50196 34847
rect 50208 34813 50220 34847
rect 50232 34813 50244 34847
rect 50232 30925 50244 30983
rect 50256 30949 50268 30983
rect 50256 30757 50268 30791
rect 47626 27173 50307 27373
rect 20280 26871 20292 26929
rect 21216 26871 21228 26905
rect 20207 26210 21096 26810
rect 46992 26341 47004 26447
rect 47016 26413 47028 26447
rect 47040 26365 47052 26447
rect 47064 26365 47076 26447
rect 47088 26365 47100 26447
rect 47112 26365 47124 26399
rect 47136 26365 47148 26471
rect 47160 26365 47172 26471
rect 47184 26365 47196 26471
rect 47208 26365 47220 26471
rect 47232 26365 47244 26471
rect 47256 26365 47268 26471
rect 47280 26365 47292 26471
rect 47304 26365 47316 26471
rect 47328 26365 47340 26471
rect 47352 26365 47364 26471
rect 47376 26365 47388 26399
rect 20304 19597 20316 19631
rect 20496 19462 21096 26210
rect 48690 26194 50307 26794
rect 46992 25237 47004 25343
rect 47016 25237 47028 25343
rect 47040 25237 47052 25343
rect 47064 25237 47076 25343
rect 47088 25309 47100 25343
rect 47112 25261 47124 25343
rect 47136 25261 47148 25343
rect 47160 25261 47172 25343
rect 47184 25261 47196 25295
rect 47208 25261 47220 25367
rect 47232 25261 47244 25367
rect 47256 25261 47268 25367
rect 47280 25261 47292 25367
rect 47304 25261 47316 25367
rect 47328 25261 47340 25367
rect 47352 25261 47364 25367
rect 47376 25261 47388 25367
rect 47400 25261 47412 25367
rect 47424 25261 47436 25295
rect 47016 24229 47028 24263
rect 47040 24229 47052 24263
rect 47064 24229 47076 24263
rect 47088 24229 47100 24263
rect 47112 24229 47124 24263
rect 47136 24229 47148 24263
rect 47160 24229 47172 24263
rect 46992 24133 47004 24167
rect 47016 24133 47028 24167
rect 47040 24133 47052 24167
rect 47064 24133 47076 24167
rect 47088 24133 47100 24167
rect 47112 24133 47124 24167
rect 47136 24133 47148 24167
rect 47184 24157 47196 24263
rect 47208 24157 47220 24263
rect 47232 24157 47244 24263
rect 47256 24157 47268 24263
rect 47280 24157 47292 24263
rect 47304 24157 47316 24263
rect 47328 24157 47340 24263
rect 47352 24157 47364 24263
rect 47376 24157 47388 24263
rect 47400 24157 47412 24263
rect 47424 24157 47436 24263
rect 47448 24157 47460 24263
rect 47472 24157 47484 24191
rect 46992 23029 47004 23111
rect 47016 23029 47028 23111
rect 47040 23029 47052 23111
rect 47064 23029 47076 23111
rect 47088 23029 47100 23111
rect 47112 23029 47124 23111
rect 47136 23029 47148 23063
rect 47160 23029 47172 23135
rect 47184 23029 47196 23135
rect 47208 23029 47220 23135
rect 47232 23029 47244 23135
rect 47256 23029 47268 23135
rect 47280 23029 47292 23135
rect 47304 23029 47316 23135
rect 47328 23029 47340 23135
rect 47352 23029 47364 23135
rect 47376 23101 47388 23135
rect 47400 23053 47412 23135
rect 47424 23053 47436 23135
rect 47448 23053 47460 23135
rect 47472 23053 47484 23135
rect 47496 23053 47508 23135
rect 47520 23053 47532 23087
rect 46992 21901 47004 22007
rect 47016 21901 47028 22007
rect 47040 21901 47052 22007
rect 47064 21901 47076 22007
rect 47088 21973 47100 22007
rect 47112 21925 47124 22007
rect 47136 21925 47148 22007
rect 47160 21925 47172 22007
rect 47184 21925 47196 22007
rect 47208 21925 47220 22007
rect 47232 21925 47244 22007
rect 47256 21925 47268 21959
rect 47280 21925 47292 22031
rect 47304 21925 47316 22031
rect 47328 21925 47340 22031
rect 47352 21925 47364 22031
rect 47376 21925 47388 22031
rect 47400 21925 47412 22031
rect 47424 21925 47436 22031
rect 47448 21925 47460 22031
rect 47472 21925 47484 22031
rect 47496 21925 47508 22031
rect 47520 21925 47532 22031
rect 47544 21925 47556 22031
rect 47568 21925 47580 21959
rect 46992 20869 47004 20903
rect 47016 20821 47028 20903
rect 47040 20821 47052 20903
rect 47064 20821 47076 20903
rect 47088 20821 47100 20903
rect 47112 20821 47124 20903
rect 47136 20821 47148 20903
rect 47160 20821 47172 20903
rect 47184 20821 47196 20903
rect 47208 20821 47220 20903
rect 47232 20821 47244 20903
rect 47256 20821 47268 20903
rect 47280 20821 47292 20903
rect 47304 20821 47316 20903
rect 47328 20821 47340 20903
rect 47352 20821 47364 20903
rect 47376 20821 47388 20903
rect 47400 20821 47412 20903
rect 47424 20821 47436 20903
rect 47448 20821 47460 20903
rect 47472 20821 47484 20903
rect 47496 20821 47508 20903
rect 47520 20821 47532 20903
rect 47544 20821 47556 20855
rect 47568 20821 47580 20927
rect 47592 20821 47604 20927
rect 47616 20821 47628 20855
rect 48690 20047 49290 26194
rect 46992 19693 47004 19775
rect 47016 19693 47028 19775
rect 47040 19693 47052 19775
rect 47064 19693 47076 19775
rect 47088 19693 47100 19775
rect 47112 19693 47124 19727
rect 47136 19693 47148 19799
rect 47160 19693 47172 19799
rect 47184 19693 47196 19799
rect 47208 19693 47220 19799
rect 47232 19693 47244 19799
rect 47256 19765 47268 19799
rect 47280 19717 47292 19799
rect 47304 19717 47316 19799
rect 47328 19717 47340 19799
rect 47352 19717 47364 19799
rect 47376 19717 47388 19799
rect 47400 19717 47412 19799
rect 47424 19717 47436 19799
rect 47448 19717 47460 19799
rect 47472 19717 47484 19799
rect 47496 19717 47508 19799
rect 47520 19717 47532 19799
rect 47544 19717 47556 19799
rect 47568 19717 47580 19799
rect 47592 19717 47604 19799
rect 47616 19717 47628 19799
rect 47640 19717 47652 19799
rect 47664 19717 47676 19751
rect 21216 19597 21228 19631
rect 21384 19597 21396 19631
rect 21432 19597 21444 19655
rect 21456 19597 21468 19655
rect 47721 19647 49290 20047
rect 21536 19621 21548 19643
rect 21559 19581 21571 19643
rect 21582 19621 21594 19643
rect 21605 19573 21617 19643
rect 21628 19532 21640 19643
rect 21651 19573 21663 19643
rect 21674 19525 21686 19643
rect 21697 19501 21709 19643
rect 20496 19262 21357 19462
rect 21905 19262 22105 19643
rect 20496 18862 22105 19262
rect 20256 18757 20268 18791
rect 20304 18421 20316 18455
rect 20256 14701 20268 14735
rect 20304 14701 20316 14735
rect 20256 10669 20268 10703
rect 20759 10136 20959 18862
rect 21552 18541 21564 18575
rect 21624 18541 21636 18623
rect 21672 18541 21684 18623
rect 21696 18469 21708 18623
rect 21216 18421 21228 18455
rect 21384 18421 21396 18455
rect 21432 18421 21444 18455
rect 21456 18421 21468 18455
rect 21480 18421 21492 18455
rect 21552 18421 21564 18455
rect 21720 18397 21732 18503
rect 21905 18354 22105 18862
rect 22121 18353 22133 19644
rect 22145 18445 22157 19643
rect 22169 18517 22181 19643
rect 22145 18354 22157 18431
rect 22169 18354 22181 18503
rect 22193 18354 22205 19643
rect 23441 19621 23453 19643
rect 23441 19607 23447 19621
rect 24233 19620 24245 19643
rect 24785 19620 24797 19643
rect 25001 19620 25013 19643
rect 25745 19620 25757 19643
rect 25913 19620 25925 19643
rect 26297 19620 26309 19643
rect 26489 19620 26501 19643
rect 26705 19620 26717 19643
rect 27449 19620 27461 19643
rect 27617 19621 27629 19643
rect 24233 19608 24252 19620
rect 24785 19608 24804 19620
rect 25001 19608 25020 19620
rect 25745 19608 25764 19620
rect 25913 19608 25932 19620
rect 26297 19608 26316 19620
rect 26489 19608 26508 19620
rect 26705 19608 26724 19620
rect 27449 19608 27468 19620
rect 24240 19573 24252 19608
rect 24792 19525 24804 19608
rect 25008 19501 25020 19608
rect 25752 19477 25764 19608
rect 25920 19477 25932 19608
rect 26304 19501 26316 19608
rect 26496 19525 26508 19608
rect 26712 19573 26724 19608
rect 26280 19429 26292 19487
rect 26472 19405 26484 19511
rect 26688 19381 26700 19559
rect 27456 19549 27468 19608
rect 27617 19607 27623 19621
rect 37025 19620 37037 19643
rect 37217 19620 37229 19643
rect 37457 19621 37469 19643
rect 45161 19621 45173 19643
rect 45905 19621 45917 19643
rect 46121 19621 46133 19643
rect 46265 19621 46277 19643
rect 46313 19621 46325 19643
rect 46361 19621 46373 19643
rect 46409 19621 46421 19643
rect 46481 19621 46493 19643
rect 37025 19608 37044 19620
rect 37217 19608 37236 19620
rect 27432 19357 27444 19535
rect 27600 19357 27612 19583
rect 37032 19549 37044 19608
rect 37224 19573 37236 19608
rect 37457 19607 37463 19621
rect 45161 19607 45167 19621
rect 45905 19607 45911 19621
rect 46121 19607 46127 19621
rect 46265 19607 46271 19621
rect 46313 19607 46319 19621
rect 46361 19607 46367 19621
rect 46409 19607 46415 19621
rect 46481 19607 46487 19621
rect 37200 19501 37212 19559
rect 37440 19501 37452 19583
rect 46721 19496 46921 19643
rect 47721 19496 48121 19647
rect 46721 19096 48121 19496
rect 48192 19309 48204 19343
rect 24168 18396 24180 18431
rect 24984 18396 24996 18503
rect 25800 18396 25812 18623
rect 27024 18541 27036 18575
rect 27456 18541 27468 18575
rect 24161 18384 24180 18396
rect 24977 18384 24996 18396
rect 25793 18384 25812 18396
rect 25824 18396 25836 18431
rect 27024 18396 27036 18431
rect 27456 18396 27468 18431
rect 25824 18384 25841 18396
rect 27024 18384 27041 18396
rect 27456 18384 27473 18396
rect 24161 18354 24173 18384
rect 24977 18354 24989 18384
rect 25793 18354 25805 18384
rect 25829 18354 25841 18384
rect 27029 18354 27041 18384
rect 27461 18354 27473 18384
rect 29057 18383 29063 18397
rect 29797 18383 29801 18397
rect 30277 18383 30281 18397
rect 31152 18396 31164 18431
rect 32040 18396 32052 18431
rect 33144 18396 33156 18431
rect 33960 18396 33972 18431
rect 31152 18384 31169 18396
rect 32040 18384 32057 18396
rect 29057 18354 29069 18383
rect 29789 18354 29801 18383
rect 30269 18354 30281 18383
rect 31157 18354 31169 18384
rect 32045 18354 32057 18384
rect 33137 18384 33156 18396
rect 33953 18384 33972 18396
rect 33984 18396 33996 18431
rect 34800 18396 34812 18431
rect 33984 18384 34001 18396
rect 34800 18384 34817 18396
rect 33137 18354 33149 18384
rect 33953 18354 33965 18384
rect 33989 18354 34001 18384
rect 34805 18354 34817 18384
rect 36389 18354 36401 18431
rect 36413 18354 36425 18431
rect 37224 18396 37236 18431
rect 37217 18384 37236 18396
rect 38016 18396 38028 18431
rect 39480 18396 39492 18431
rect 38016 18384 38033 18396
rect 39480 18384 39497 18396
rect 37217 18354 37229 18384
rect 38021 18354 38033 18384
rect 39485 18354 39497 18384
rect 40409 18354 40421 18431
rect 40433 18354 40445 18431
rect 41232 18396 41244 18431
rect 42816 18396 42828 18431
rect 43512 18396 43524 18455
rect 43632 18421 43644 18479
rect 44424 18445 44436 18503
rect 45240 18469 45252 18503
rect 41232 18384 41249 18396
rect 42816 18384 42833 18396
rect 43512 18384 43529 18396
rect 41237 18354 41249 18384
rect 42821 18354 42833 18384
rect 43517 18354 43529 18384
rect 43649 18383 43655 18397
rect 44448 18396 44460 18431
rect 45264 18396 45276 18455
rect 44448 18384 44465 18396
rect 43649 18354 43661 18383
rect 44453 18354 44465 18384
rect 45257 18384 45276 18396
rect 46056 18396 46068 18479
rect 46056 18384 46073 18396
rect 45257 18354 45269 18384
rect 46061 18354 46073 18384
rect 46865 18383 46871 18397
rect 46865 18354 46877 18383
rect 47921 18354 48121 19096
rect 48360 18397 48372 19103
rect 48384 18397 48396 19079
rect 48408 18397 48420 19055
rect 48432 18397 48444 19031
rect 48456 18397 48468 19007
rect 48480 18397 48492 18983
rect 48504 18397 48516 18959
rect 48528 18397 48540 18935
rect 48552 18397 48564 18911
rect 48576 18397 48588 18887
rect 48600 18397 48612 18863
rect 48624 18397 48636 18839
rect 48648 18397 48660 18815
rect 48672 18397 48684 18791
rect 48696 18397 48708 18743
rect 48720 18397 48732 18719
rect 48744 18397 48756 18695
rect 48768 18397 48780 18671
rect 48840 18397 48852 18647
rect 48864 18397 48876 18599
rect 48888 18397 48900 18575
rect 48912 18397 48924 18551
rect 48936 18397 48948 18527
rect 48984 18397 48996 18503
rect 21432 18176 21444 18215
rect 21456 18152 21468 18215
rect 21480 18152 21492 18215
rect 21720 18152 21732 18215
rect 21757 18187 21782 18199
rect 21757 18163 21782 18175
rect 48303 18139 48330 18151
rect 48303 18115 48330 18127
rect 48303 18091 48330 18103
rect 48303 18067 48330 18079
rect 48303 18043 48330 18055
rect 48360 18033 48372 18163
rect 48384 18033 48396 18163
rect 48408 18033 48420 18163
rect 48432 18033 48444 18163
rect 48456 18033 48468 18163
rect 48504 18033 48516 18139
rect 48528 18033 48540 18139
rect 48552 18033 48564 18139
rect 48576 18057 48588 18139
rect 48624 18081 48636 18115
rect 48648 18081 48660 18115
rect 48672 18081 48684 18115
rect 48696 18081 48708 18115
rect 48720 18081 48732 18115
rect 48744 18081 48756 18115
rect 48768 18081 48780 18115
rect 48792 18081 48804 18115
rect 48816 18081 48828 18115
rect 21216 14701 21228 14735
rect 21456 14701 21468 14735
rect 21480 14701 21492 14735
rect 48303 14605 48349 14606
rect 48303 14594 48335 14605
rect 48360 14581 48372 14615
rect 48384 14581 48396 14615
rect 48408 14581 48420 14615
rect 48432 14581 48444 14615
rect 48456 14581 48468 14615
rect 48504 14581 48516 14615
rect 48528 14581 48540 14615
rect 48552 14581 48564 14615
rect 48648 14581 48660 14615
rect 48672 14581 48684 14615
rect 48696 14581 48708 14615
rect 48720 14581 48732 14615
rect 21456 13957 21468 13993
rect 21480 13957 21492 13993
rect 21757 13970 21782 13982
rect 21757 13946 21782 13958
rect 48303 13189 48349 13190
rect 48303 13178 48335 13189
rect 48360 13165 48372 13199
rect 48384 13165 48396 13199
rect 48408 13165 48420 13199
rect 48432 13165 48444 13199
rect 48456 13165 48468 13199
rect 48504 13165 48516 13199
rect 48528 13165 48540 13199
rect 48303 12925 48349 12926
rect 48303 12914 48335 12925
rect 48360 12901 48372 12935
rect 48384 12901 48396 12935
rect 48408 12901 48420 12935
rect 48432 12901 48444 12935
rect 48456 12901 48468 12935
rect 48504 12901 48516 12935
rect 48528 12901 48540 12935
rect 48303 12589 48349 12590
rect 48303 12578 48335 12589
rect 48360 12565 48372 12599
rect 48384 12565 48396 12599
rect 48408 12565 48420 12599
rect 48432 12565 48444 12599
rect 48456 12565 48468 12599
rect 48504 12565 48516 12599
rect 48303 10789 48349 10797
rect 48303 10785 48335 10789
rect 48360 10765 48372 10799
rect 48384 10765 48396 10799
rect 48408 10765 48420 10799
rect 48432 10765 48444 10799
rect 48456 10765 48468 10799
rect 48504 10765 48516 10799
rect 48672 10765 48684 10799
rect 48696 10765 48708 10799
rect 48864 10717 48876 10751
rect 48888 10717 48900 10751
rect 48912 10717 48924 10751
rect 48936 10717 48948 10751
rect 48984 10717 48996 10751
rect 48384 10525 48396 10559
rect 48408 10525 48420 10559
rect 48432 10525 48444 10559
rect 48456 10525 48468 10559
rect 48504 10525 48516 10559
rect 48672 10525 48684 10559
rect 48696 10525 48708 10559
rect 48768 10525 48780 10559
rect 48792 10525 48804 10559
rect 48864 10525 48876 10559
rect 48888 10525 48900 10559
rect 48912 10525 48924 10559
rect 48936 10525 48948 10559
rect 48984 10525 48996 10559
rect 21456 10165 21468 10376
rect 21757 10353 21782 10365
rect 48303 10353 48335 10365
rect 21757 10329 21782 10341
rect 48303 10329 48335 10341
rect 48303 10309 48349 10317
rect 48303 10305 48335 10309
rect 21720 10165 21732 10247
rect 21905 10136 22105 10294
rect 22121 10260 22133 10294
rect 22193 10261 22205 10294
rect 22121 10248 22140 10260
rect 22128 10213 22140 10248
rect 22193 10247 22199 10261
rect 29453 10260 29465 10294
rect 29448 10248 29465 10260
rect 35561 10260 35573 10294
rect 41549 10260 41561 10294
rect 35561 10248 35580 10260
rect 29448 10237 29460 10248
rect 35568 10237 35580 10248
rect 41544 10248 41561 10260
rect 41681 10260 41693 10294
rect 41681 10248 41700 10260
rect 41544 10237 41556 10248
rect 41688 10237 41700 10248
rect 29448 10165 29460 10223
rect 29472 10189 29484 10223
rect 35568 10165 35580 10223
rect 35592 10189 35604 10223
rect 20759 9936 22105 10136
rect 31800 10117 31812 10151
rect 38856 10117 38868 10175
rect 41544 10117 41556 10223
rect 41568 10189 41580 10223
rect 41688 10117 41700 10223
rect 31656 10021 31668 10055
rect 31800 10021 31812 10055
rect 38856 10021 38868 10055
rect 41544 10021 41556 10055
rect 21130 9829 21142 9936
rect 24744 9901 24756 9935
rect 28128 9901 28140 9935
rect 28272 9901 28284 9935
rect 31656 9901 31668 9935
rect 31800 9901 31812 9935
rect 38712 9901 38724 9935
rect 38856 9901 38868 9959
rect 42240 9901 42252 10223
rect 21720 9853 21732 9887
rect 24600 9805 24612 9839
rect 24744 9805 24756 9839
rect 28128 9805 28140 9839
rect 28272 9805 28284 9839
rect 31656 9805 31668 9839
rect 31800 9805 31812 9839
rect 38712 9805 38724 9839
rect 38856 9805 38868 9839
rect 42240 9805 42252 9839
rect 42384 9805 42396 9839
rect 45768 9805 45780 9863
rect 45912 9805 45924 10175
rect 45984 9829 45996 10246
rect 47836 9998 47848 10103
rect 47921 10083 48121 10294
rect 48384 10141 48396 10377
rect 48408 10285 48420 10377
rect 48432 10342 48444 10377
rect 48456 10285 48468 10377
rect 48504 10285 48516 10377
rect 48672 10232 48684 10377
rect 48768 10232 48780 10319
rect 48792 10285 48804 10319
rect 48864 10238 48876 10319
rect 48888 10261 48900 10319
rect 48912 10285 48924 10319
rect 48936 10285 48948 10319
rect 48984 10285 48996 10319
rect 48888 10249 49038 10261
rect 48456 10189 48468 10223
rect 48864 10226 49010 10238
rect 48568 10196 48982 10208
rect 49090 10083 49290 19647
rect 50256 18757 50268 18791
rect 50256 18613 50268 18647
rect 50112 18397 50124 18479
rect 50160 18397 50172 18455
rect 50208 18397 50220 18431
rect 50208 14725 50220 14759
rect 50208 14581 50220 14615
rect 50208 10717 50220 10751
rect 50256 10669 50268 10703
rect 50256 10525 50268 10559
rect 46032 9853 46044 9887
rect 47921 9883 49290 10083
<< metal4 >>
rect 20373 44585 21933 46145
rect 23899 44585 25459 46145
rect 27425 44585 28985 46145
rect 30951 44585 32511 46145
rect 34477 44585 36037 46145
rect 38003 44585 39563 46145
rect 41529 44585 43089 46145
rect 45055 44585 46615 46145
rect 48581 44585 50141 46145
rect 13835 38133 15395 39693
rect 55119 38133 56679 39693
rect 13835 34091 15395 35651
rect 55119 34091 56679 35651
rect 13835 30049 15395 31609
rect 55119 30049 56679 31609
rect 13835 26007 15395 27567
rect 55119 26007 56679 27567
rect 13835 21965 15395 23525
rect 55119 21965 56679 23525
rect 13835 17923 15395 19483
rect 55119 17923 56679 19483
rect 13835 13881 15395 15441
rect 55119 13881 56679 15441
rect 13835 9839 15395 11399
rect 55119 9839 56679 11399
rect 20373 3387 21933 4947
rect 23899 3387 25459 4947
rect 27425 3387 28985 4947
rect 30951 3387 32511 4947
rect 34477 3387 36037 4947
rect 38003 3387 39563 4947
rect 41529 3387 43089 4947
rect 45055 3387 46615 4947
rect 48581 3387 50141 4947
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 13757 -1 0 46223
box 0 0 6450 6450
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 20293 1 0 39773
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 22013 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 22099 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 22185 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 22271 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 22357 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 22443 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 22529 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 22615 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 22701 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 22787 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 22873 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 22959 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 23045 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 23131 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 23217 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 23303 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 23389 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 23475 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 23561 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 23647 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 23733 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 23819 1 0 39773
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 25539 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 25625 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 25711 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 25797 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 25883 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 25969 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 26055 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 26141 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 26227 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 26313 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 26399 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 26485 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 26571 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 26657 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 26743 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 26829 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 26915 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 27001 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 27087 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 27173 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 27259 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 27345 1 0 39773
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 29065 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 29151 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 29237 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 29323 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 29409 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 29495 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 29581 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 29667 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 29753 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 29839 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 29925 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 30011 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 0 -1 30097 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 0 -1 30183 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 0 -1 30269 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 0 -1 30355 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 0 -1 30441 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 0 -1 30527 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 0 -1 30613 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 0 -1 30699 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 0 -1 30785 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 0 -1 30871 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 32591 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 0 -1 32677 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 0 -1 32763 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 0 -1 32849 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 0 -1 32935 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 0 -1 33021 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 0 -1 33107 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 0 -1 33193 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 0 -1 33279 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 0 -1 33365 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 0 -1 33451 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 0 -1 33537 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 0 -1 33623 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 0 -1 33709 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 0 -1 33795 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 0 -1 33881 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 0 -1 33967 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 0 -1 34053 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 0 -1 34139 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 0 -1 34225 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 0 -1 34311 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 0 -1 34397 1 0 39773
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 36117 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 0 -1 36203 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 0 -1 36289 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 0 -1 36375 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 0 -1 36461 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 0 -1 36547 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 0 -1 36633 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 0 -1 36719 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 0 -1 36805 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 0 -1 36891 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 0 -1 36977 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 0 -1 37063 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 0 -1 37149 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 0 -1 37235 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 0 -1 37321 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 0 -1 37407 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 0 -1 37493 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 0 -1 37579 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 0 -1 37665 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 0 -1 37751 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 0 -1 37837 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 0 -1 37923 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 39643 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 0 -1 39729 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 0 -1 39815 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 0 -1 39901 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 0 -1 39987 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 0 -1 40073 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 0 -1 40159 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 0 -1 40245 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 0 -1 40331 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 0 -1 40417 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 0 -1 40503 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 0 -1 40589 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 0 -1 40675 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 0 -1 40761 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 0 -1 40847 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 0 -1 40933 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 0 -1 41019 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 0 -1 41105 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 0 -1 41191 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 0 -1 41277 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 0 -1 41363 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 0 -1 41449 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 43169 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 0 -1 43255 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 0 -1 43341 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 0 -1 43427 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 0 -1 43513 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 0 -1 43599 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 0 -1 43685 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 0 -1 43771 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 0 -1 43857 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 0 -1 43943 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 0 -1 44029 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 0 -1 44115 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 0 -1 44201 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 0 -1 44287 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 0 -1 44373 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 0 -1 44459 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 0 -1 44545 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 0 -1 44631 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 0 -1 44717 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 0 -1 44803 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 0 -1 44889 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 0 -1 44975 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 46695 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 0 -1 46781 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 0 -1 46867 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 0 -1 46953 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 0 -1 47039 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 0 -1 47125 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 0 -1 47211 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 0 -1 47297 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 0 -1 47383 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 0 -1 47469 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 0 -1 47555 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 0 -1 47641 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 0 -1 47727 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 0 -1 47813 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 0 -1 47899 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 0 -1 47985 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 0 -1 48071 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 0 -1 48157 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 0 -1 48243 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 0 -1 48329 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 0 -1 48415 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 0 -1 48501 1 0 39773
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 50221 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 0 -1 50307 1 0 39773
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 56757 0 -1 46223
box 0 0 6450 6450
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 20207 0 -1 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform -1 0 20207 0 -1 38053
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform -1 0 20207 0 -1 37967
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform -1 0 20207 0 -1 37881
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform -1 0 20207 0 -1 37795
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform -1 0 20207 0 -1 37709
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform -1 0 20207 0 -1 37623
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform -1 0 20207 0 -1 37537
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform -1 0 20207 0 -1 37451
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform -1 0 20207 0 -1 37365
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform -1 0 20207 0 -1 37279
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform -1 0 20207 0 -1 37193
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform -1 0 20207 0 -1 37107
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform -1 0 20207 0 -1 37021
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform -1 0 20207 0 -1 36935
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform -1 0 20207 0 -1 36849
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform -1 0 20207 0 -1 36763
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform -1 0 20207 0 -1 36677
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform -1 0 20207 0 -1 36591
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform -1 0 20207 0 -1 36505
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform -1 0 20207 0 -1 36419
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform -1 0 20207 0 -1 36333
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform -1 0 20207 0 -1 36247
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform -1 0 20207 0 -1 36161
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform -1 0 20207 0 -1 36075
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform -1 0 20207 0 -1 35989
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform -1 0 20207 0 -1 35903
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform -1 0 20207 0 -1 35817
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 20207 0 -1 35731
box 0 0 6450 1720
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform -1 0 20207 0 -1 34011
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform -1 0 20207 0 -1 33925
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform -1 0 20207 0 -1 33839
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform -1 0 20207 0 -1 33753
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform -1 0 20207 0 -1 33667
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform -1 0 20207 0 -1 33581
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform -1 0 20207 0 -1 33495
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform -1 0 20207 0 -1 33409
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform -1 0 20207 0 -1 33323
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform -1 0 20207 0 -1 33237
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform -1 0 20207 0 -1 33151
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform -1 0 20207 0 -1 33065
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform -1 0 20207 0 -1 32979
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform -1 0 20207 0 -1 32893
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform -1 0 20207 0 -1 32807
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform -1 0 20207 0 -1 32721
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform -1 0 20207 0 -1 32635
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform -1 0 20207 0 -1 32549
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform -1 0 20207 0 -1 32463
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform -1 0 20207 0 -1 32377
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform -1 0 20207 0 -1 32291
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform -1 0 20207 0 -1 32205
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform -1 0 20207 0 -1 32119
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform -1 0 20207 0 -1 32033
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform -1 0 20207 0 -1 31947
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform -1 0 20207 0 -1 31861
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform -1 0 20207 0 -1 31775
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 20207 0 -1 31689
box 0 0 6450 1720
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform -1 0 20207 0 -1 29969
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform -1 0 20207 0 -1 29883
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform -1 0 20207 0 -1 29797
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform -1 0 20207 0 -1 29711
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform -1 0 20207 0 -1 29625
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform -1 0 20207 0 -1 29539
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform -1 0 20207 0 -1 29453
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform -1 0 20207 0 -1 29367
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform -1 0 20207 0 -1 29281
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform -1 0 20207 0 -1 29195
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform -1 0 20207 0 -1 29109
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform -1 0 20207 0 -1 29023
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform -1 0 20207 0 -1 28937
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform -1 0 20207 0 -1 28851
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform -1 0 20207 0 -1 28765
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform -1 0 20207 0 -1 28679
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform -1 0 20207 0 -1 28593
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform -1 0 20207 0 -1 28507
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform -1 0 20207 0 -1 28421
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform -1 0 20207 0 -1 28335
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform -1 0 20207 0 -1 28249
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform -1 0 20207 0 -1 28163
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform -1 0 20207 0 -1 28077
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform -1 0 20207 0 -1 27991
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform -1 0 20207 0 -1 27905
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform -1 0 20207 0 -1 27819
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform -1 0 20207 0 -1 27733
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 20207 0 -1 27647
box 0 0 6450 1720
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform -1 0 20207 0 -1 25927
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform -1 0 20207 0 -1 25841
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform -1 0 20207 0 -1 25755
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform -1 0 20207 0 -1 25669
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform -1 0 20207 0 -1 25583
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform -1 0 20207 0 -1 25497
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform -1 0 20207 0 -1 25411
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform -1 0 20207 0 -1 25325
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform -1 0 20207 0 -1 25239
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform -1 0 20207 0 -1 25153
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform -1 0 20207 0 -1 25067
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform -1 0 20207 0 -1 24981
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform -1 0 20207 0 -1 24895
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform -1 0 20207 0 -1 24809
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform -1 0 20207 0 -1 24723
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform -1 0 20207 0 -1 24637
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform -1 0 20207 0 -1 24551
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform -1 0 20207 0 -1 24465
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform -1 0 20207 0 -1 24379
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform -1 0 20207 0 -1 24293
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform -1 0 20207 0 -1 24207
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform -1 0 20207 0 -1 24121
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform -1 0 20207 0 -1 24035
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform -1 0 20207 0 -1 23949
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform -1 0 20207 0 -1 23863
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform -1 0 20207 0 -1 23777
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform -1 0 20207 0 -1 23691
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 20207 0 -1 23605
box 0 0 6450 1720
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform -1 0 20207 0 -1 21885
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform -1 0 20207 0 -1 21799
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform -1 0 20207 0 -1 21713
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform -1 0 20207 0 -1 21627
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform -1 0 20207 0 -1 21541
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform -1 0 20207 0 -1 21455
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform -1 0 20207 0 -1 21369
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform -1 0 20207 0 -1 21283
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform -1 0 20207 0 -1 21197
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform -1 0 20207 0 -1 21111
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform -1 0 20207 0 -1 21025
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform -1 0 20207 0 -1 20939
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform -1 0 20207 0 -1 20853
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform -1 0 20207 0 -1 20767
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform -1 0 20207 0 -1 20681
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform -1 0 20207 0 -1 20595
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform -1 0 20207 0 -1 20509
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform -1 0 20207 0 -1 20423
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform -1 0 20207 0 -1 20337
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform -1 0 20207 0 -1 20251
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform -1 0 20207 0 -1 20165
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform -1 0 20207 0 -1 20079
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform -1 0 20207 0 -1 19993
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform -1 0 20207 0 -1 19907
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform -1 0 20207 0 -1 19821
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform -1 0 20207 0 -1 19735
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform -1 0 20207 0 -1 19649
box 0 0 6450 86
use datapath datapath_0
timestamp 1396540370
transform 1 0 21535 0 1 19643
box 0 0 25408 19490
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 50307 0 1 38053
box 0 0 6450 1720
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 50307 0 1 37967
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 50307 0 1 37881
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 50307 0 1 37795
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 50307 0 1 37709
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 50307 0 1 37623
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 50307 0 1 37537
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 50307 0 1 37451
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 50307 0 1 37365
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 50307 0 1 37279
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 50307 0 1 37193
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 50307 0 1 37107
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 50307 0 1 37021
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 50307 0 1 36935
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 50307 0 1 36849
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 50307 0 1 36763
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 50307 0 1 36677
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 50307 0 1 36591
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 50307 0 1 36505
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 50307 0 1 36419
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 50307 0 1 36333
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 50307 0 1 36247
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 50307 0 1 36161
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 50307 0 1 36075
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 50307 0 1 35989
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 50307 0 1 35903
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 50307 0 1 35817
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 50307 0 1 35731
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 50307 0 1 34011
box 0 0 6450 1720
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 50307 0 1 33925
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 50307 0 1 33839
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 50307 0 1 33753
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 50307 0 1 33667
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 50307 0 1 33581
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 50307 0 1 33495
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 50307 0 1 33409
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 50307 0 1 33323
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 50307 0 1 33237
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 50307 0 1 33151
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 50307 0 1 33065
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 50307 0 1 32979
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 50307 0 1 32893
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 50307 0 1 32807
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 50307 0 1 32721
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 50307 0 1 32635
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 50307 0 1 32549
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 50307 0 1 32463
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 50307 0 1 32377
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 50307 0 1 32291
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 50307 0 1 32205
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 50307 0 1 32119
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 50307 0 1 32033
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 50307 0 1 31947
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 50307 0 1 31861
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 50307 0 1 31775
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 50307 0 1 31689
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 50307 0 1 29969
box 0 0 6450 1720
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 50307 0 1 29883
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 50307 0 1 29797
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 50307 0 1 29711
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 50307 0 1 29625
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 50307 0 1 29539
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 50307 0 1 29453
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 50307 0 1 29367
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 50307 0 1 29281
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 50307 0 1 29195
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 50307 0 1 29109
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 50307 0 1 29023
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 50307 0 1 28937
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 50307 0 1 28851
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 50307 0 1 28765
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 50307 0 1 28679
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 50307 0 1 28593
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 50307 0 1 28507
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 50307 0 1 28421
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 50307 0 1 28335
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 50307 0 1 28249
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 50307 0 1 28163
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 50307 0 1 28077
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 50307 0 1 27991
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 50307 0 1 27905
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 50307 0 1 27819
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 50307 0 1 27733
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 50307 0 1 27647
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 50307 0 1 25927
box 0 0 6450 1720
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 50307 0 1 25841
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 50307 0 1 25755
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 50307 0 1 25669
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 50307 0 1 25583
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 50307 0 1 25497
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 50307 0 1 25411
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 50307 0 1 25325
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 50307 0 1 25239
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 50307 0 1 25153
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 50307 0 1 25067
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 50307 0 1 24981
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 50307 0 1 24895
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 50307 0 1 24809
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 50307 0 1 24723
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 50307 0 1 24637
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 50307 0 1 24551
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 50307 0 1 24465
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 50307 0 1 24379
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 50307 0 1 24293
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 50307 0 1 24207
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 50307 0 1 24121
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 50307 0 1 24035
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 50307 0 1 23949
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 50307 0 1 23863
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 50307 0 1 23777
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 50307 0 1 23691
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 50307 0 1 23605
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 50307 0 1 21885
box 0 0 6450 1720
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 50307 0 1 21799
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 50307 0 1 21713
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 50307 0 1 21627
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 50307 0 1 21541
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 50307 0 1 21455
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 50307 0 1 21369
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 50307 0 1 21283
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 50307 0 1 21197
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 50307 0 1 21111
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 50307 0 1 21025
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 50307 0 1 20939
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 50307 0 1 20853
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 50307 0 1 20767
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 50307 0 1 20681
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 50307 0 1 20595
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 50307 0 1 20509
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 50307 0 1 20423
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 50307 0 1 20337
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 50307 0 1 20251
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 50307 0 1 20165
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 50307 0 1 20079
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 50307 0 1 19993
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 50307 0 1 19907
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 1 0 50307 0 1 19821
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 1 0 50307 0 1 19735
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 1 0 50307 0 1 19649
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 20207 0 -1 19563
box 0 0 6450 1720
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 1 0 50307 0 1 19563
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform -1 0 20207 0 -1 17843
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform -1 0 20207 0 -1 17757
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform -1 0 20207 0 -1 17671
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform -1 0 20207 0 -1 17585
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform -1 0 20207 0 -1 17499
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform -1 0 20207 0 -1 17413
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform -1 0 20207 0 -1 17327
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform -1 0 20207 0 -1 17241
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform -1 0 20207 0 -1 17155
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform -1 0 20207 0 -1 17069
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform -1 0 20207 0 -1 16983
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform -1 0 20207 0 -1 16897
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform -1 0 20207 0 -1 16811
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform -1 0 20207 0 -1 16725
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform -1 0 20207 0 -1 16639
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform -1 0 20207 0 -1 16553
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform -1 0 20207 0 -1 16467
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform -1 0 20207 0 -1 16381
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform -1 0 20207 0 -1 16295
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform -1 0 20207 0 -1 16209
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform -1 0 20207 0 -1 16123
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform -1 0 20207 0 -1 16037
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform -1 0 20207 0 -1 15951
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform -1 0 20207 0 -1 15865
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform -1 0 20207 0 -1 15779
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform -1 0 20207 0 -1 15693
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform -1 0 20207 0 -1 15607
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 20207 0 -1 15521
box 0 0 6450 1720
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform -1 0 20207 0 -1 13801
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform -1 0 20207 0 -1 13715
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform -1 0 20207 0 -1 13629
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform -1 0 20207 0 -1 13543
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform -1 0 20207 0 -1 13457
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform -1 0 20207 0 -1 13371
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform -1 0 20207 0 -1 13285
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform -1 0 20207 0 -1 13199
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform -1 0 20207 0 -1 13113
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform -1 0 20207 0 -1 13027
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform -1 0 20207 0 -1 12941
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform -1 0 20207 0 -1 12855
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 20207 0 -1 12769
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 20207 0 -1 12683
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 20207 0 -1 12597
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 20207 0 -1 12511
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 20207 0 -1 12425
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 20207 0 -1 12339
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 20207 0 -1 12253
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 20207 0 -1 12167
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 20207 0 -1 12081
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 20207 0 -1 11995
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 20207 0 -1 11909
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 20207 0 -1 11823
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 20207 0 -1 11737
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 20207 0 -1 11651
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 20207 0 -1 11565
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 20207 0 -1 11479
box 0 0 6450 1720
use control control_0
timestamp 1395929462
transform 1 0 21782 0 1 10294
box 0 0 26521 8060
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 50307 0 1 17843
box 0 0 6450 1720
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 1 0 50307 0 1 17757
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 1 0 50307 0 1 17671
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 1 0 50307 0 1 17585
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 1 0 50307 0 1 17499
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 1 0 50307 0 1 17413
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 1 0 50307 0 1 17327
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 1 0 50307 0 1 17241
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 1 0 50307 0 1 17155
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 1 0 50307 0 1 17069
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 1 0 50307 0 1 16983
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 1 0 50307 0 1 16897
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 1 0 50307 0 1 16811
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 1 0 50307 0 1 16725
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 1 0 50307 0 1 16639
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 1 0 50307 0 1 16553
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 1 0 50307 0 1 16467
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 1 0 50307 0 1 16381
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 1 0 50307 0 1 16295
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 1 0 50307 0 1 16209
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 1 0 50307 0 1 16123
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 1 0 50307 0 1 16037
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 1 0 50307 0 1 15951
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 1 0 50307 0 1 15865
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 1 0 50307 0 1 15779
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 1 0 50307 0 1 15693
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 1 0 50307 0 1 15607
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 1 0 50307 0 1 15521
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 50307 0 1 13801
box 0 0 6450 1720
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 1 0 50307 0 1 13715
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 1 0 50307 0 1 13629
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 1 0 50307 0 1 13543
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 1 0 50307 0 1 13457
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 1 0 50307 0 1 13371
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 1 0 50307 0 1 13285
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 1 0 50307 0 1 13199
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 1 0 50307 0 1 13113
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 1 0 50307 0 1 13027
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 1 0 50307 0 1 12941
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 1 0 50307 0 1 12855
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 1 0 50307 0 1 12769
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 1 0 50307 0 1 12683
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 1 0 50307 0 1 12597
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 1 0 50307 0 1 12511
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 1 0 50307 0 1 12425
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 1 0 50307 0 1 12339
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 1 0 50307 0 1 12253
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 1 0 50307 0 1 12167
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 1 0 50307 0 1 12081
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 1 0 50307 0 1 11995
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 1 0 50307 0 1 11909
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 1 0 50307 0 1 11823
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 1 0 50307 0 1 11737
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 1 0 50307 0 1 11651
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 1 0 50307 0 1 11565
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 1 0 50307 0 1 11479
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 50307 0 1 9759
box 0 0 6450 1720
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 13757 0 1 3309
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 20207 -1 0 9759
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 20293 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 22013 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 22099 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 22185 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 22271 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 22357 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 22443 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 22529 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 22615 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 22701 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 22787 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 22873 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 22959 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 23045 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 23131 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 23217 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 23303 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 23389 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 23475 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 23561 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 23647 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 23733 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 23819 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 25539 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 25625 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 25711 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 25797 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 25883 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 25969 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 26055 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 26141 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 26227 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 26313 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 26399 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 26485 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 26571 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 26657 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 26743 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 26829 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 26915 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 27001 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 27087 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 27173 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 27259 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 27345 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 29065 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 29151 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 29237 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 29323 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 29409 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 29495 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 29581 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 29667 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 29753 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 29839 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 29925 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 30011 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 30097 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 30183 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 30269 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 30355 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 30441 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 30527 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 30613 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 30699 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 30785 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 30871 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 32591 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 32677 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 32763 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 32849 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 32935 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 33021 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 33107 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 33193 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 33279 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 33365 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 33451 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 33537 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 33623 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 33709 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 33795 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 33881 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 33967 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 34053 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 34139 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 34225 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 34311 -1 0 9759
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 34397 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 36117 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 36203 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 36289 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 36375 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 36461 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 36547 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 36633 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 36719 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 36805 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 36891 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 36977 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 37063 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 37149 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 37235 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 37321 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 37407 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 37493 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 37579 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 37665 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 37751 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 37837 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 37923 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 39643 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 39729 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 39815 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 39901 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 39987 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 40073 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 40159 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 40245 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 40331 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 40417 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 40503 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 40589 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 40675 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 40761 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 40847 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 40933 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 41019 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 41105 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 41191 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 41277 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 41363 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 41449 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 43169 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 43255 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 43341 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 43427 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 43513 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 43599 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 43685 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 43771 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 43857 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 43943 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 44029 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 44115 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 44201 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 44287 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 44373 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 44459 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 44545 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 44631 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 44717 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 44803 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 44889 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 44975 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 46695 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 46781 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 46867 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 46953 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 47039 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 47125 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 47211 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 47297 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 47383 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 47469 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 47555 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 47641 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 47727 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 47813 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 47899 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 47985 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 48071 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 48157 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 48243 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 48329 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 48415 -1 0 9759
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 48501 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 50221 -1 0 9759
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 56757 1 0 3309
box 0 0 6450 6450
<< labels >>
rlabel metal4 20373 3387 21933 4947 0 nIRQ
rlabel metal4 23899 3387 25459 4947 0 Data[0]
rlabel metal4 27425 3387 28985 4947 0 Data[1]
rlabel metal4 30951 3387 32511 4947 0 Data[2]
rlabel metal4 34477 3387 36037 4947 0 vdde!
rlabel metal4 38003 3387 39563 4947 0 Data[3]
rlabel metal4 41529 3387 43089 4947 0 Data[4]
rlabel metal4 45055 3387 46615 4947 0 Data[5]
rlabel metal4 48581 3387 50141 4947 0 gnde!
rlabel metal4 55119 9839 56679 11399 0 Data[6]
rlabel metal4 55119 13881 56679 15441 0 Data[7]
rlabel metal4 55119 17923 56679 19483 0 Data[8]
rlabel metal4 55119 21965 56679 23525 0 gnde!
rlabel metal4 55119 26007 56679 27567 0 GND!
rlabel metal4 55119 30049 56679 31609 0 Data[9]
rlabel metal4 55119 34091 56679 35651 0 Data[10]
rlabel metal4 55119 38133 56679 39693 0 Data[11]
rlabel metal4 48581 44585 50141 46145 0 vdde!
rlabel metal4 45055 44585 46615 46145 0 Data[12]
rlabel metal4 41529 44585 43089 46145 0 Data[13]
rlabel metal4 38003 44585 39563 46145 0 Data[14]
rlabel metal4 34477 44585 36037 46145 0 gnde!
rlabel metal4 30951 44585 32511 46145 0 Data[15]
rlabel metal4 27425 44585 28985 46145 0 ALE
rlabel metal4 23899 44585 25459 46145 0 nME
rlabel metal4 20373 44585 21933 46145 0 nWait
rlabel metal4 13835 38133 15395 39693 0 nOE
rlabel metal4 13835 34091 15395 35651 0 RnW
rlabel metal4 13835 30049 15395 31609 0 SDO
rlabel metal4 13835 26007 15395 27567 0 Vdd!
rlabel metal4 13835 21965 15395 23525 0 SDI
rlabel metal4 13835 17923 15395 19483 0 Test
rlabel metal4 13835 13881 15395 15441 0 Clock
rlabel metal4 13835 9839 15395 11399 0 nReset
<< end >>
