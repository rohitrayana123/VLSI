magic
tech c035u
timestamp 1394564637
<< metal1 >>
rect 0 16478 35 16488
rect 2987 16478 3040 16488
rect 0 16455 35 16465
rect 2987 16455 3040 16465
rect 0 16417 35 16442
rect 2987 16417 3040 16442
rect 0 15772 35 15797
rect 2987 15772 3040 15797
rect 0 15749 35 15759
rect 2987 15749 3040 15759
rect 0 15726 35 15736
rect 2987 15726 3040 15736
rect 0 15703 35 15713
rect 2987 15703 3040 15713
rect 8 15436 35 15446
rect 2987 15436 3040 15446
rect 8 15413 35 15423
rect 2987 15413 3040 15423
rect 8 15375 35 15400
rect 2987 15375 3040 15400
rect 0 14730 35 14755
rect 2987 14730 3040 14755
rect 0 14707 35 14717
rect 2987 14707 3040 14717
rect 0 14684 35 14694
rect 2987 14684 3040 14694
rect 0 14661 35 14671
rect 2987 14661 3040 14671
rect 0 14394 35 14404
rect 2987 14394 3040 14404
rect 0 14371 35 14381
rect 2987 14371 3040 14381
rect 0 14333 35 14358
rect 2987 14333 3040 14358
rect 0 13688 35 13713
rect 2987 13688 3040 13713
rect 0 13665 35 13675
rect 2987 13665 3040 13675
rect 0 13642 35 13652
rect 2987 13642 3040 13652
rect 0 13619 35 13629
rect 2987 13619 3040 13629
rect 0 13352 35 13362
rect 2987 13352 3040 13362
rect 0 13329 35 13339
rect 2987 13329 3040 13339
rect 0 13291 35 13316
rect 2987 13291 3040 13316
rect 0 12646 35 12671
rect 2987 12646 3040 12671
rect 0 12623 35 12633
rect 2987 12623 3040 12633
rect 0 12600 35 12610
rect 2987 12600 3040 12610
rect 0 12577 35 12587
rect 2987 12577 3040 12587
rect 0 12310 35 12320
rect 2987 12310 3040 12320
rect 0 12287 35 12297
rect 2987 12287 3040 12297
rect 0 12249 35 12274
rect 2987 12249 3040 12274
rect 0 11604 35 11629
rect 2987 11604 3040 11629
rect 0 11581 35 11591
rect 2987 11581 3040 11591
rect 0 11558 35 11568
rect 2987 11558 3040 11568
rect 0 11535 35 11545
rect 2987 11535 3040 11545
rect 0 11268 35 11278
rect 2987 11268 3040 11278
rect 0 11245 35 11255
rect 2987 11245 3040 11255
rect 0 11207 35 11232
rect 2987 11207 3040 11232
rect 0 10562 35 10587
rect 2987 10562 3040 10587
rect 0 10539 35 10549
rect 2987 10539 3040 10549
rect 0 10516 35 10526
rect 2987 10516 3040 10526
rect 0 10493 35 10503
rect 2987 10493 3040 10503
rect 0 10226 35 10236
rect 2987 10226 3040 10236
rect 0 10203 35 10213
rect 2987 10203 3040 10213
rect 0 10165 35 10190
rect 2987 10165 3040 10190
rect 0 9520 35 9545
rect 2987 9520 3040 9545
rect 0 9497 35 9507
rect 2987 9497 3040 9507
rect 0 9474 35 9484
rect 2987 9474 3040 9484
rect 0 9451 35 9461
rect 2987 9451 3040 9461
rect 0 9184 35 9194
rect 2987 9184 3040 9194
rect 0 9161 35 9171
rect 2987 9161 3040 9171
rect 0 9123 35 9148
rect 2987 9123 3040 9148
rect 0 8478 35 8503
rect 2987 8478 3040 8503
rect 0 8455 35 8465
rect 2987 8455 3040 8465
rect 0 8432 35 8442
rect 2987 8432 3040 8442
rect 0 8409 35 8419
rect 2987 8409 3040 8419
rect 0 8142 35 8152
rect 2987 8142 3040 8152
rect 0 8119 35 8129
rect 2987 8119 3040 8129
rect 0 8081 35 8106
rect 2987 8081 3040 8106
rect 0 7436 35 7461
rect 2987 7436 3040 7461
rect 0 7413 35 7423
rect 2987 7413 3040 7423
rect 0 7390 35 7400
rect 2987 7390 3040 7400
rect 0 7367 35 7377
rect 2987 7367 3040 7377
rect 0 7100 35 7110
rect 2987 7100 3040 7110
rect 0 7077 35 7087
rect 2987 7077 3040 7087
rect 0 7039 35 7064
rect 2987 7039 3040 7064
rect 0 6394 35 6419
rect 2987 6394 3040 6419
rect 0 6371 35 6381
rect 2987 6371 3040 6381
rect 0 6348 35 6358
rect 2987 6348 3040 6358
rect 0 6325 35 6335
rect 2987 6325 3040 6335
rect 0 6058 35 6068
rect 2987 6058 3040 6068
rect 0 6035 35 6045
rect 2987 6035 3040 6045
rect 0 5997 35 6022
rect 2987 5997 3040 6022
rect 0 5352 35 5377
rect 2987 5352 3040 5377
rect 0 5329 35 5339
rect 2987 5329 3040 5339
rect 0 5306 35 5316
rect 2987 5306 3040 5316
rect 0 5283 35 5293
rect 2987 5283 3040 5293
rect 0 5016 35 5026
rect 2987 5016 3040 5026
rect 0 4993 35 5003
rect 2987 4993 3040 5003
rect 0 4955 35 4980
rect 2987 4955 3040 4980
rect 0 4310 35 4335
rect 2987 4310 3040 4335
rect 0 4287 35 4297
rect 2987 4287 3040 4297
rect 0 4264 35 4274
rect 2987 4264 3040 4274
rect 0 4241 35 4251
rect 2987 4241 3040 4251
rect 0 3974 35 3984
rect 2987 3974 3040 3984
rect 0 3951 35 3961
rect 2987 3951 3040 3961
rect 0 3913 35 3938
rect 2987 3913 3040 3938
rect 0 3268 35 3293
rect 2987 3268 3040 3293
rect 0 3245 35 3255
rect 2987 3245 3040 3255
rect 0 3222 35 3232
rect 2987 3222 3040 3232
rect 0 3199 35 3209
rect 2987 3199 3040 3209
rect 0 2932 35 2942
rect 2987 2932 3040 2942
rect 0 2909 35 2919
rect 2987 2909 3040 2919
rect 0 2871 35 2896
rect 2987 2871 3040 2896
rect 0 2226 35 2251
rect 2987 2226 3040 2251
rect 0 2203 35 2213
rect 2987 2203 3040 2213
rect 0 2180 35 2190
rect 2987 2180 3040 2190
rect 0 2157 35 2167
rect 2987 2157 3040 2167
rect 0 1890 35 1900
rect 2987 1890 3040 1900
rect 0 1867 35 1877
rect 2987 1867 3040 1877
rect 0 1829 35 1854
rect 2987 1829 3040 1854
rect 0 1184 35 1209
rect 2987 1184 3040 1209
rect 0 1161 35 1171
rect 2987 1161 3040 1171
rect 0 1138 35 1148
rect 2987 1138 3040 1148
rect 0 1115 35 1125
rect 2987 1115 3040 1125
rect 0 848 35 858
rect 2987 848 3040 858
rect 0 825 35 835
rect 2987 825 3040 835
rect 0 787 35 812
rect 2987 787 3040 812
rect 0 142 35 167
rect 2987 142 3040 167
rect 0 119 35 129
rect 2987 119 3040 129
rect 0 96 35 106
rect 2987 96 3040 106
rect 0 73 35 83
rect 2987 73 3040 83
<< metal2 >>
rect 395 16672 407 16872
rect 611 16672 623 16872
rect 1355 16672 1367 16872
rect 1523 16672 1535 16872
rect 1595 16672 1607 16872
rect 1907 16672 1919 16872
rect 2123 16672 2135 16872
rect 2867 16672 2879 16872
rect 2939 16672 2951 16872
use Pc_slice.mag Pc_slice.mag_15
timestamp 1394563293
transform 1 0 35 0 1 15630
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_14
timestamp 1394563293
transform 1 0 35 0 1 14588
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_13
timestamp 1394563293
transform 1 0 35 0 1 13546
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_12
timestamp 1394563293
transform 1 0 35 0 1 12504
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_11
timestamp 1394563293
transform 1 0 35 0 1 11462
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_10
timestamp 1394563293
transform 1 0 35 0 1 10420
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_9
timestamp 1394563293
transform 1 0 35 0 1 9378
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_8
timestamp 1394563293
transform 1 0 35 0 1 8336
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_7
timestamp 1394563293
transform 1 0 35 0 1 7294
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_6
timestamp 1394563293
transform 1 0 35 0 1 6252
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_5
timestamp 1394563293
transform 1 0 35 0 1 5210
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_4
timestamp 1394563293
transform 1 0 35 0 1 4168
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_3
timestamp 1394563293
transform 1 0 35 0 1 3126
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_2
timestamp 1394563293
transform 1 0 35 0 1 2084
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_1
timestamp 1394563293
transform 1 0 35 0 1 1042
box 0 0 2952 1042
use Pc_slice.mag Pc_slice.mag_0
timestamp 1394563293
transform 1 0 35 0 1 0
box 0 0 2952 1042
<< labels >>
rlabel metal1 8 15375 8 15400 3 Vdd!
rlabel metal1 8 15413 8 15423 3 Scan
rlabel metal1 8 15436 8 15446 3 ScanReturn
rlabel metal1 0 73 0 83 3 nReset
rlabel metal1 0 96 0 106 3 Test
rlabel metal1 0 119 0 129 3 Clock
rlabel metal1 0 142 0 167 3 GND!
rlabel metal1 0 1867 0 1877 3 Scan
rlabel metal1 0 1890 0 1900 3 ScanReturn
rlabel metal1 0 1829 0 1854 3 Vdd!
rlabel metal1 0 1184 0 1209 3 GND!
rlabel metal1 0 1115 0 1125 3 nReset
rlabel metal1 0 1138 0 1148 3 Test
rlabel metal1 0 1161 0 1171 3 Clock
rlabel metal1 0 848 0 858 3 ScanReturn
rlabel metal1 0 825 0 835 3 Scan
rlabel metal1 0 787 0 812 3 Vdd!
rlabel metal1 0 2157 0 2167 3 nReset
rlabel metal1 0 2180 0 2190 3 Test
rlabel metal1 0 2203 0 2213 3 Clock
rlabel metal1 0 2226 0 2251 3 GND!
rlabel metal1 0 2932 0 2942 3 ScanReturn
rlabel metal1 0 2909 0 2919 3 Scan
rlabel metal1 0 2871 0 2896 3 Vdd!
rlabel metal1 0 3268 0 3293 3 GND!
rlabel metal1 0 3222 0 3232 3 Test
rlabel metal1 0 3245 0 3255 3 Clock
rlabel metal1 0 3199 0 3209 3 nReset
rlabel metal1 0 3974 0 3984 3 ScanReturn
rlabel metal1 0 3951 0 3961 3 Scan
rlabel metal1 0 3913 0 3938 3 Vdd!
rlabel metal1 0 6058 0 6068 3 ScanReturn
rlabel metal1 0 6035 0 6045 3 Scan
rlabel metal1 0 5997 0 6022 3 Vdd!
rlabel metal1 0 6394 0 6419 3 GND!
rlabel metal1 0 6348 0 6358 3 Test
rlabel metal1 0 6371 0 6381 3 Clock
rlabel metal1 0 6325 0 6335 3 nReset
rlabel metal1 0 7100 0 7110 3 ScanReturn
rlabel metal1 0 7077 0 7087 3 Scan
rlabel metal1 0 7039 0 7064 3 Vdd!
rlabel metal1 0 7436 0 7461 3 GND!
rlabel metal1 0 7390 0 7400 3 Test
rlabel metal1 0 7413 0 7423 3 Clock
rlabel metal1 0 7367 0 7377 3 nReset
rlabel metal1 0 9123 0 9148 3 Vdd!
rlabel metal1 0 9161 0 9171 3 Scan
rlabel metal1 0 9184 0 9194 3 ScanReturn
rlabel metal1 0 9520 0 9545 3 GND!
rlabel metal1 0 9451 0 9461 3 nReset
rlabel metal1 0 9474 0 9484 3 Test
rlabel metal1 0 9497 0 9507 3 Clock
rlabel metal1 0 10226 0 10236 3 ScanReturn
rlabel metal1 0 10203 0 10213 3 Scan
rlabel metal1 0 10165 0 10190 3 Vdd!
rlabel metal1 0 10562 0 10587 3 GND!
rlabel metal1 0 10539 0 10549 3 Clock
rlabel metal1 0 10516 0 10526 3 Test
rlabel metal1 0 10493 0 10503 3 nReset
rlabel metal1 0 11268 0 11278 3 ScanReturn
rlabel metal1 0 11245 0 11255 3 Scan
rlabel metal1 0 11207 0 11232 3 Vdd!
rlabel metal1 0 11604 0 11629 3 GND!
rlabel metal1 0 11558 0 11568 3 Test
rlabel metal1 0 11581 0 11591 3 Clock
rlabel metal1 0 11535 0 11545 3 nReset
rlabel metal1 0 12249 0 12274 3 Vdd!
rlabel metal1 0 15772 0 15797 3 GND!
rlabel metal1 0 15703 0 15713 3 nReset
rlabel metal1 0 15726 0 15736 3 Test
rlabel metal1 0 15749 0 15759 3 Clock
rlabel metal1 0 8478 0 8503 3 GND!
rlabel metal1 0 8432 0 8442 3 Test
rlabel metal1 0 8455 0 8465 3 Clock
rlabel metal1 0 8409 0 8419 3 nReset
rlabel metal1 0 4310 0 4335 3 GND!
rlabel metal1 0 4264 0 4274 3 Test
rlabel metal1 0 4287 0 4297 3 Clock
rlabel metal1 0 4241 0 4251 3 nReset
rlabel metal1 0 4955 0 4980 3 Vdd!
rlabel metal1 0 4993 0 5003 3 Scan
rlabel metal1 0 5016 0 5026 3 ScanReturn
rlabel metal1 0 5352 0 5377 3 GND!
rlabel metal1 0 5306 0 5316 3 Test
rlabel metal1 0 5329 0 5339 3 Clock
rlabel metal1 0 5283 0 5293 3 nReset
rlabel metal1 0 12646 0 12671 3 GND!
rlabel metal1 0 12600 0 12610 3 Test
rlabel metal1 0 12623 0 12633 3 Clock
rlabel metal1 0 12577 0 12587 3 nReset
rlabel metal1 0 12287 0 12297 3 Scan
rlabel metal1 0 12310 0 12320 3 ScanReturn
rlabel metal1 0 14333 0 14358 3 Vdd!
rlabel metal1 0 14371 0 14381 3 Scan
rlabel metal1 0 14394 0 14404 3 ScanReturn
rlabel metal1 0 14661 0 14671 3 nReset
rlabel metal1 0 14684 0 14694 3 Test
rlabel metal1 0 14707 0 14717 3 Clock
rlabel metal1 0 14730 0 14755 3 GND!
rlabel metal1 0 13619 0 13629 3 nReset
rlabel metal1 0 13642 0 13652 3 Test
rlabel metal1 0 13665 0 13675 3 Clock
rlabel metal1 0 13688 0 13713 3 GND!
rlabel metal1 0 16478 0 16488 3 ScanReturn
rlabel metal1 0 16455 0 16465 3 Scan
rlabel metal1 0 16417 0 16442 3 Vdd!
rlabel metal1 0 13291 0 13316 3 Vdd!
rlabel metal1 0 13329 0 13339 3 Scan
rlabel metal1 0 13352 0 13362 3 ScanReturn
rlabel metal1 0 8142 0 8152 3 ScanReturn
rlabel metal1 0 8119 0 8129 3 Scan
rlabel metal1 0 8081 0 8106 3 Vdd!
rlabel metal1 3040 1115 3040 1125 7 nReset
rlabel metal1 3040 1138 3040 1148 7 Test
rlabel metal1 3040 1161 3040 1171 7 Clock
rlabel metal1 3040 1184 3040 1209 7 GND!
rlabel metal1 3040 73 3040 83 7 nReset
rlabel metal1 3040 96 3040 106 7 Test
rlabel metal1 3040 119 3040 129 7 Clock
rlabel metal1 3040 142 3040 167 7 GND!
rlabel metal1 3040 787 3040 812 7 Vdd!
rlabel metal1 3040 825 3040 835 7 Scan
rlabel metal1 3040 848 3040 858 7 ScanReturn
rlabel metal1 3040 1890 3040 1900 7 ScanReturn
rlabel metal1 3040 1867 3040 1877 7 Scan
rlabel metal1 3040 1829 3040 1854 7 Vdd!
rlabel metal1 3040 2226 3040 2251 7 GND!
rlabel metal1 3040 2203 3040 2213 7 Clock
rlabel metal1 3040 2180 3040 2190 7 Test
rlabel metal1 3040 2157 3040 2167 7 nReset
rlabel metal1 3040 3268 3040 3293 7 GND!
rlabel metal1 3040 3245 3040 3255 7 Clock
rlabel metal1 3040 3222 3040 3232 7 Test
rlabel metal1 3040 3199 3040 3209 7 nReset
rlabel metal1 3040 2932 3040 2942 7 ScanReturn
rlabel metal1 3040 2909 3040 2919 7 Scan
rlabel metal1 3040 2871 3040 2896 7 Vdd!
rlabel metal1 3040 4310 3040 4335 7 GND!
rlabel metal1 3040 4287 3040 4297 7 Clock
rlabel metal1 3040 4264 3040 4274 7 Test
rlabel metal1 3040 4241 3040 4251 7 nReset
rlabel metal1 3040 6058 3040 6068 7 ScanReturn
rlabel metal1 3040 6035 3040 6045 7 Scan
rlabel metal1 3040 5997 3040 6022 7 Vdd!
rlabel metal1 3040 6394 3040 6419 7 GND!
rlabel metal1 3040 6371 3040 6381 7 Clock
rlabel metal1 3040 6348 3040 6358 7 Test
rlabel metal1 3040 6325 3040 6335 7 nReset
rlabel metal1 3040 3974 3040 3984 7 ScanReturn
rlabel metal1 3040 3951 3040 3961 7 Scan
rlabel metal1 3040 3913 3040 3938 7 Vdd!
rlabel metal1 3040 7436 3040 7461 7 GND!
rlabel metal1 3040 7413 3040 7423 7 Clock
rlabel metal1 3040 7390 3040 7400 7 Test
rlabel metal1 3040 7367 3040 7377 7 nReset
rlabel metal1 3040 8119 3040 8129 7 Scan
rlabel metal1 3040 8081 3040 8106 7 Vdd!
rlabel metal1 3040 8142 3040 8152 7 ScanReturn
rlabel metal1 3040 7100 3040 7110 7 ScanReturn
rlabel metal1 3040 7077 3040 7087 7 Scan
rlabel metal1 3040 7039 3040 7064 7 Vdd!
rlabel metal1 3040 8478 3040 8503 7 GND!
rlabel metal1 3040 8455 3040 8465 7 Clock
rlabel metal1 3040 8432 3040 8442 7 Test
rlabel metal1 3040 8409 3040 8419 7 nReset
rlabel metal1 3040 9520 3040 9545 7 GND!
rlabel metal1 3040 9497 3040 9507 7 Clock
rlabel metal1 3040 9474 3040 9484 7 Test
rlabel metal1 3040 9451 3040 9461 7 nReset
rlabel metal1 3040 9184 3040 9194 7 ScanReturn
rlabel metal1 3040 9161 3040 9171 7 Scan
rlabel metal1 3040 9123 3040 9148 7 Vdd!
rlabel metal1 3040 10165 3040 10190 7 Vdd!
rlabel metal1 3040 10203 3040 10213 7 Scan
rlabel metal1 3040 10226 3040 10236 7 ScanReturn
rlabel metal1 3040 11604 3040 11629 7 GND!
rlabel metal1 3040 11581 3040 11591 7 Clock
rlabel metal1 3040 11558 3040 11568 7 Test
rlabel metal1 3040 11535 3040 11545 7 nReset
rlabel metal1 3040 12310 3040 12320 7 ScanReturn
rlabel metal1 3040 12287 3040 12297 7 Scan
rlabel metal1 3040 12249 3040 12274 7 Vdd!
rlabel metal1 3040 11268 3040 11278 7 ScanReturn
rlabel metal1 3040 11245 3040 11255 7 Scan
rlabel metal1 3040 11207 3040 11232 7 Vdd!
rlabel metal1 3040 10562 3040 10587 7 GND!
rlabel metal1 3040 10539 3040 10549 7 Clock
rlabel metal1 3040 10516 3040 10526 7 Test
rlabel metal1 3040 10493 3040 10503 7 nReset
rlabel metal1 3040 12646 3040 12671 7 GND!
rlabel metal1 3040 12623 3040 12633 7 Clock
rlabel metal1 3040 12600 3040 12610 7 Test
rlabel metal1 3040 12577 3040 12587 7 nReset
rlabel metal1 3040 13688 3040 13713 7 GND!
rlabel metal1 3040 13665 3040 13675 7 Clock
rlabel metal1 3040 13642 3040 13652 7 Test
rlabel metal1 3040 13619 3040 13629 7 nReset
rlabel metal1 3040 13352 3040 13362 7 ScanReturn
rlabel metal1 3040 13329 3040 13339 7 Scan
rlabel metal1 3040 13291 3040 13316 7 Vdd!
rlabel metal1 3040 15375 3040 15400 7 Vdd!
rlabel metal1 3040 15413 3040 15423 7 Scan
rlabel metal1 3040 15436 3040 15446 7 ScanReturn
rlabel metal1 3040 14661 3040 14671 7 nReset
rlabel metal1 3040 14684 3040 14694 7 Test
rlabel metal1 3040 14707 3040 14717 7 Clock
rlabel metal1 3040 14730 3040 14755 7 GND!
rlabel metal1 3040 14333 3040 14358 7 Vdd!
rlabel metal1 3040 14371 3040 14381 7 Scan
rlabel metal1 3040 14394 3040 14404 7 ScanReturn
rlabel metal1 3040 15703 3040 15713 7 nReset
rlabel metal1 3040 15726 3040 15736 7 Test
rlabel metal1 3040 15749 3040 15759 7 Clock
rlabel metal1 3040 15772 3040 15797 7 GND!
rlabel metal1 3040 16417 3040 16442 7 Vdd!
rlabel metal1 3040 16455 3040 16465 7 Scan
rlabel metal1 3040 16478 3040 16488 7 ScanReturn
rlabel metal1 3040 5016 3040 5026 7 ScanReturn
rlabel metal1 3040 4993 3040 5003 7 Scan
rlabel metal1 3040 4955 3040 4980 7 Vdd!
rlabel metal1 3040 5352 3040 5377 7 GND!
rlabel metal1 3040 5329 3040 5339 7 Clock
rlabel metal1 3040 5306 3040 5316 7 Test
rlabel metal1 3040 5283 3040 5293 7 nReset
rlabel metal2 395 16872 407 16872 5 LrSel
rlabel metal2 611 16872 623 16872 5 LrWe
rlabel metal2 1355 16872 1367 16872 5 LrEn
rlabel metal2 1523 16872 1535 16872 5 PcSel[0]
rlabel metal2 1595 16872 1607 16872 5 ALU
rlabel metal2 1907 16872 1919 16872 5 PcSel[1]
rlabel metal2 2123 16872 2135 16872 5 PcWe
rlabel metal2 2867 16872 2879 16872 5 PcEn
rlabel metal2 2939 16872 2951 16872 5 SysBus
<< end >>
