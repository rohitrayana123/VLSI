magic
tech c035u
timestamp 1394145165
<< metal1 >>
rect 805 970 935 980
rect 757 942 887 952
rect 0 57 599 67
rect 973 57 1008 67
<< m2contact >>
rect 791 968 805 982
rect 935 968 949 982
rect 743 940 757 954
rect 887 940 901 954
rect 599 55 613 69
rect 959 55 973 69
<< metal2 >>
rect 744 954 756 1023
rect 792 982 804 1023
rect 744 901 756 940
rect 792 901 804 968
rect 864 901 876 1023
rect 888 901 900 940
rect 936 901 948 968
rect 600 69 612 102
rect 744 0 756 102
rect 792 0 804 102
rect 960 69 972 102
use scanreg  scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 102
box 0 0 720 799
use rowcrosser  rowcrosser_0
timestamp 1386086759
transform 1 0 720 0 1 102
box 0 0 48 799
use rowcrosser  rowcrosser_1
timestamp 1386086759
transform 1 0 768 0 1 102
box 0 0 48 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 816 0 1 102
box 0 0 192 799
<< labels >>
rlabel metal1 0 57 0 67 3 Ir
rlabel metal1 1008 57 1008 67 7 Imm
rlabel metal2 744 1023 756 1023 5 Ext0
rlabel metal2 792 1023 804 1023 5 Ext1
rlabel metal2 864 1023 876 1023 5 ImmSel
rlabel metal2 744 0 756 0 1 Ext0
rlabel metal2 792 0 804 0 1 Ext1
<< end >>
