../../../Design/Implementation/verilog/behavioural/ram.sv