magic
tech c035u
timestamp 1395695751
<< checkpaint >>
rect -13483 -2099 14222 8465
<< metal1 >>
rect -12183 6766 -12133 7165
rect -419 7143 10115 7153
rect -3251 7117 -3233 7131
rect -2363 7117 -2345 7131
rect -1499 7119 9299 7129
rect -4595 7095 1955 7105
rect 6841 7095 6959 7105
rect 7657 7095 8159 7105
rect -10403 7069 -10385 7083
rect -8435 7071 -6289 7081
rect -4787 7071 -1321 7081
rect -803 7071 1139 7081
rect 3577 7071 3695 7081
rect 4309 7069 4327 7083
rect 6301 7071 12815 7081
rect -10811 7045 -10793 7059
rect -10427 7047 -9601 7057
rect -8579 7047 -7117 7057
rect -7043 7047 -2149 7057
rect -1643 7047 4403 7057
rect 6025 7047 9431 7057
rect -12099 7023 -6361 7033
rect -5051 7023 7667 7033
rect -12099 6999 1943 7009
rect 3565 6999 12743 7009
rect -11345 6975 -9265 6985
rect -9251 6975 -913 6985
rect -899 6975 5591 6985
rect 5605 6975 12047 6985
rect 12733 6975 12767 6985
rect -7967 6951 -7345 6961
rect -7139 6951 -4729 6961
rect -4655 6951 11879 6961
rect -6539 6927 455 6937
rect 469 6927 6863 6937
rect 6877 6927 10931 6937
rect 12757 6927 12838 6937
rect -3827 6903 7199 6913
rect 8029 6903 8483 6913
rect 8941 6903 11747 6913
rect 12805 6903 12838 6913
rect -587 6879 12743 6889
rect 12781 6879 12838 6889
rect 313 6855 11327 6865
rect 12757 6855 12838 6865
rect 1129 6831 8735 6841
rect 10285 6831 12791 6841
rect 12829 6831 12838 6841
rect -12183 6741 -12096 6766
rect -12183 989 -12133 6741
rect 12872 6121 12922 7165
rect 12744 6096 12922 6121
rect 7405 5998 8783 6008
rect -1667 5974 10967 5984
rect -1979 5950 -1033 5960
rect -1019 5950 5615 5960
rect 5629 5950 6455 5960
rect 6469 5950 7487 5960
rect 7501 5950 11687 5960
rect -2027 5926 11327 5936
rect -2075 5902 2327 5912
rect 2437 5902 7391 5912
rect 7405 5902 12263 5912
rect -2363 5878 -2353 5888
rect -2195 5878 2423 5888
rect -3419 5854 -1993 5864
rect -1811 5854 10151 5864
rect -3875 5830 -3817 5840
rect -3683 5830 10199 5840
rect -3947 5806 5255 5816
rect -4043 5782 1631 5792
rect -4403 5758 1871 5768
rect -4499 5734 -3409 5744
rect -2987 5734 -97 5744
rect -83 5734 1079 5744
rect 1093 5734 4271 5744
rect 4285 5734 4391 5744
rect 4405 5734 6695 5744
rect 6709 5734 8183 5744
rect 8197 5734 10103 5744
rect 10117 5734 10583 5744
rect -4619 5710 -3121 5720
rect -3107 5710 2687 5720
rect 2701 5710 11879 5720
rect -4715 5686 -3673 5696
rect -3659 5686 2351 5696
rect 2365 5686 2999 5696
rect 3013 5686 4343 5696
rect 4357 5686 5591 5696
rect 5605 5686 6791 5696
rect -4883 5662 -4801 5672
rect -4739 5662 -4729 5672
rect -4643 5662 -769 5672
rect 6229 5662 6335 5672
rect -4955 5638 1487 5648
rect 5149 5638 8975 5648
rect -4979 5614 9887 5624
rect -5219 5590 12455 5600
rect -5219 5566 10871 5576
rect -5315 5542 -49 5552
rect 4741 5542 11999 5552
rect -5435 5518 -1273 5528
rect -1211 5518 12838 5528
rect -5579 5494 -5329 5504
rect -5267 5494 10751 5504
rect 10765 5494 11231 5504
rect -5603 5470 -409 5480
rect 4477 5470 8231 5480
rect 8245 5470 9479 5480
rect -5651 5446 6671 5456
rect 11437 5446 11903 5456
rect -5747 5422 6527 5432
rect 10933 5422 11807 5432
rect -5987 5398 -5761 5408
rect -5699 5398 -2689 5408
rect -2675 5398 935 5408
rect 949 5398 2063 5408
rect 2077 5398 6671 5408
rect 6685 5398 8519 5408
rect 8533 5398 10919 5408
rect 10933 5398 11423 5408
rect -6059 5374 11279 5384
rect -6107 5350 -193 5360
rect 4261 5350 9239 5360
rect -6179 5326 -5977 5336
rect -5891 5326 6215 5336
rect -6203 5302 1847 5312
rect 1861 5302 6743 5312
rect 7165 5302 7367 5312
rect 7381 5302 7511 5312
rect 9781 5302 9791 5312
rect -6395 5278 1439 5288
rect 2317 5278 2399 5288
rect 4141 5278 9935 5288
rect -6467 5254 -5893 5264
rect -5879 5254 -5785 5264
rect -5771 5254 -5473 5264
rect -5459 5254 -5017 5264
rect -5003 5254 -4057 5264
rect -4043 5254 -2737 5264
rect -2723 5254 -2665 5264
rect -2651 5254 -2545 5264
rect -2531 5254 2951 5264
rect 2965 5254 4199 5264
rect 4213 5254 7151 5264
rect 7165 5254 9287 5264
rect 9301 5254 9767 5264
rect 9781 5254 11951 5264
rect -6467 5230 8159 5240
rect -6515 5206 9575 5216
rect -6515 5182 -1369 5192
rect -1283 5182 1079 5192
rect 2197 5182 6455 5192
rect 9373 5182 9455 5192
rect -6611 5158 12767 5168
rect -6635 5134 -2617 5144
rect -2603 5134 -2377 5144
rect -2363 5134 191 5144
rect 2101 5134 9359 5144
rect -6659 5110 8471 5120
rect -6683 5086 3767 5096
rect 3781 5086 8111 5096
rect -6731 5062 -1 5072
rect 2053 5062 10847 5072
rect -6827 5038 1559 5048
rect 2029 5038 3935 5048
rect 3997 5038 4967 5048
rect 4981 5038 6623 5048
rect 11485 5038 12119 5048
rect -6899 5014 -4273 5024
rect -4139 5014 -3433 5024
rect -3251 5014 -25 5024
rect 1933 5014 12239 5024
rect -7115 4990 -1249 5000
rect -1235 4990 8039 5000
rect 8053 4990 11471 5000
rect -7139 4966 -4513 4976
rect -4499 4966 12479 4976
rect -7211 4942 7295 4952
rect -7331 4918 -7321 4928
rect -7235 4918 8279 4928
rect -7451 4894 -4321 4904
rect -4307 4894 -2785 4904
rect -2771 4894 10655 4904
rect 10669 4894 11663 4904
rect 11677 4894 11735 4904
rect -7451 4870 12383 4880
rect -7619 4846 3239 4856
rect 3253 4846 5135 4856
rect 5149 4846 12047 4856
rect -7739 4822 -3793 4832
rect -3731 4822 -1201 4832
rect 1909 4822 4799 4832
rect 4861 4822 7031 4832
rect 7045 4822 7319 4832
rect 8725 4822 8735 4832
rect -7883 4798 -4705 4808
rect -4691 4798 12239 4808
rect -7907 4774 4031 4784
rect 4093 4774 6119 4784
rect 6133 4774 6983 4784
rect 6997 4774 12695 4784
rect -8075 4750 -5569 4760
rect -5435 4750 9527 4760
rect -8195 4726 -6817 4736
rect -6803 4726 -2185 4736
rect -2171 4726 -1129 4736
rect -1115 4726 2207 4736
rect 2221 4726 2255 4736
rect 2269 4726 3191 4736
rect 3205 4726 6287 4736
rect 6301 4726 8711 4736
rect -8219 4702 -6889 4712
rect -6875 4702 -4825 4712
rect -4811 4702 -4609 4712
rect -4595 4702 8231 4712
rect -8219 4678 -5545 4688
rect -5483 4678 2663 4688
rect 3757 4678 9335 4688
rect -8243 4654 -7705 4664
rect -7691 4654 -5401 4664
rect -5387 4654 -5161 4664
rect -5147 4654 -3145 4664
rect -3131 4654 -2761 4664
rect -2747 4654 -241 4664
rect -227 4654 2735 4664
rect 2941 4654 3887 4664
rect 3901 4654 12431 4664
rect -8315 4630 5903 4640
rect 5917 4630 6599 4640
rect -8771 4606 -5353 4616
rect -5339 4606 -4537 4616
rect -4523 4606 -2305 4616
rect -2291 4606 647 4616
rect 661 4606 2711 4616
rect 2725 4606 5975 4616
rect 5989 4606 10079 4616
rect -8795 4582 -8785 4592
rect -8651 4582 -625 4592
rect -611 4582 -397 4592
rect -383 4582 6383 4592
rect 6397 4582 7223 4592
rect 7237 4582 7367 4592
rect 7381 4582 9431 4592
rect 11869 4582 12599 4592
rect -8867 4558 -2641 4568
rect -2627 4558 11855 4568
rect -8891 4534 -505 4544
rect 1813 4534 7679 4544
rect -8915 4510 4223 4520
rect 4237 4510 10175 4520
rect -8939 4486 -8185 4496
rect -8123 4486 -6793 4496
rect -6779 4486 11519 4496
rect 11533 4486 11543 4496
rect 11557 4486 12527 4496
rect -8963 4462 6815 4472
rect 6925 4462 7079 4472
rect 7621 4462 7631 4472
rect -8987 4438 -6409 4448
rect -6395 4438 -6289 4448
rect -6275 4438 -337 4448
rect -323 4438 4655 4448
rect 4669 4438 8327 4448
rect -9059 4414 -3649 4424
rect -3467 4414 1199 4424
rect 1765 4414 11351 4424
rect -9083 4390 -3961 4400
rect -3947 4390 -3601 4400
rect -3539 4390 12095 4400
rect -9131 4366 8375 4376
rect -9155 4342 12191 4352
rect -9227 4318 -6433 4328
rect -6419 4318 10679 4328
rect -9299 4294 -8593 4304
rect -8579 4294 2975 4304
rect 2989 4294 3743 4304
rect 3757 4294 6143 4304
rect 6157 4294 7127 4304
rect 7141 4294 7607 4304
rect 7621 4294 8255 4304
rect 8269 4294 9503 4304
rect 9517 4294 11135 4304
rect -9419 4270 -1441 4280
rect -1307 4270 -1153 4280
rect -875 4270 -265 4280
rect 1597 4270 11087 4280
rect -9443 4246 -673 4256
rect 1525 4246 8423 4256
rect -9467 4222 -3241 4232
rect -3035 4222 -3025 4232
rect -2699 4222 -2593 4232
rect -2459 4222 -97 4232
rect 1477 4222 9311 4232
rect -9539 4198 -7873 4208
rect -7763 4198 -4177 4208
rect -4163 4198 -2905 4208
rect -2891 4198 2111 4208
rect 2125 4198 5639 4208
rect 5653 4198 6935 4208
rect 6949 4198 11399 4208
rect -9611 4174 -2857 4184
rect -2843 4174 8303 4184
rect -9659 4150 -3745 4160
rect -3731 4150 -2113 4160
rect -2099 4150 2135 4160
rect 2149 4150 5879 4160
rect 5893 4150 6911 4160
rect 6925 4150 7487 4160
rect -9683 4126 -7249 4136
rect -7235 4126 -2953 4136
rect -2939 4126 -145 4136
rect -131 4126 1127 4136
rect 1141 4126 2087 4136
rect 2101 4126 4895 4136
rect 5821 4126 12071 4136
rect -9923 4102 -3385 4112
rect -3371 4102 -73 4112
rect 685 4102 695 4112
rect 1285 4102 1295 4112
rect 1429 4102 10127 4112
rect -9971 4078 -9817 4088
rect -9803 4078 6479 4088
rect 10909 4078 11447 4088
rect -10019 4054 -9793 4064
rect -9779 4054 -6865 4064
rect -6851 4054 -6745 4064
rect -6731 4054 -6025 4064
rect -6011 4054 -4585 4064
rect -4571 4054 -4009 4064
rect -3995 4054 -2041 4064
rect -2027 4054 7463 4064
rect 7477 4054 11015 4064
rect 11029 4054 12143 4064
rect -10067 4030 11831 4040
rect -10091 4006 -6433 4016
rect -6419 4006 -4105 4016
rect -4091 4006 -1249 4016
rect -1235 4006 10895 4016
rect -10115 3982 -1009 3992
rect -923 3982 3647 3992
rect 3661 3982 8015 3992
rect -10283 3958 -3169 3968
rect -3059 3958 5783 3968
rect -10307 3934 -8497 3944
rect -8483 3934 -3673 3944
rect -3659 3934 -2137 3944
rect -2123 3934 1175 3944
rect 1261 3934 10703 3944
rect -10331 3910 -3649 3920
rect -3635 3910 -3313 3920
rect -3299 3910 9143 3920
rect 9157 3910 12311 3920
rect -10403 3886 -5665 3896
rect -5651 3886 -1177 3896
rect -1163 3886 5831 3896
rect 5845 3886 6239 3896
rect 6253 3886 7943 3896
rect 7957 3886 11495 3896
rect -10475 3862 1607 3872
rect 1717 3862 5039 3872
rect 5125 3862 5447 3872
rect 5509 3862 6023 3872
rect -10499 3838 -7801 3848
rect -7787 3838 -6457 3848
rect -6443 3838 -2617 3848
rect -2603 3838 -1321 3848
rect -1307 3838 -313 3848
rect -299 3838 1031 3848
rect 1045 3838 2855 3848
rect 2869 3838 3215 3848
rect 3229 3838 5111 3848
rect 5125 3838 6695 3848
rect 6709 3838 7175 3848
rect 7189 3838 7343 3848
rect 7357 3838 8975 3848
rect 8989 3838 10343 3848
rect 10357 3838 11591 3848
rect 11605 3838 12071 3848
rect -10523 3814 6503 3824
rect 9637 3814 12575 3824
rect -10571 3790 12359 3800
rect -10595 3766 -7585 3776
rect -7571 3766 4679 3776
rect 4693 3766 9047 3776
rect 9061 3766 12647 3776
rect -10619 3742 -2833 3752
rect -2819 3742 12623 3752
rect -10643 3718 -4801 3728
rect -4787 3718 2567 3728
rect 2629 3718 6407 3728
rect 7285 3718 7535 3728
rect 9205 3718 9383 3728
rect 9613 3718 10295 3728
rect -10643 3694 6959 3704
rect 7117 3694 7415 3704
rect 9085 3694 12838 3704
rect -10691 3670 -4753 3680
rect -4739 3670 -721 3680
rect 61 3670 9647 3680
rect 9997 3670 10775 3680
rect -10739 3646 -5473 3656
rect -5459 3646 4991 3656
rect 5005 3646 6095 3656
rect 6109 3646 8399 3656
rect 8629 3646 12743 3656
rect -10787 3622 -6841 3632
rect -6827 3622 -4921 3632
rect -4907 3622 2447 3632
rect 2605 3622 12491 3632
rect -10811 3598 -961 3608
rect -947 3598 5567 3608
rect 5581 3598 7823 3608
rect 7837 3598 12023 3608
rect -10883 3574 1727 3584
rect 1789 3574 11255 3584
rect -10883 3550 3695 3560
rect 3925 3550 10823 3560
rect 11317 3550 11555 3560
rect -10931 3526 -9889 3536
rect -9875 3526 -9577 3536
rect -9563 3526 -4561 3536
rect -4547 3526 -2881 3536
rect -2867 3526 1151 3536
rect 1165 3526 3431 3536
rect 3445 3526 5651 3536
rect 5665 3526 6767 3536
rect 6781 3526 9095 3536
rect 9109 3526 10463 3536
rect 10477 3526 11831 3536
rect 12421 3526 12671 3536
rect -10955 3502 -7297 3512
rect -7283 3502 3455 3512
rect 4213 3502 12599 3512
rect -11003 3478 -5809 3488
rect -5795 3478 -1057 3488
rect -923 3478 2975 3488
rect 2989 3478 7079 3488
rect 8173 3478 8183 3488
rect 8461 3478 9407 3488
rect 9925 3478 12551 3488
rect -11051 3454 -9769 3464
rect -9755 3454 -4345 3464
rect -4163 3454 1991 3464
rect 2533 3454 6419 3464
rect 6433 3454 12119 3464
rect -11099 3430 -5257 3440
rect -5171 3430 -2929 3440
rect -2915 3430 -2521 3440
rect -2507 3430 -2257 3440
rect -2243 3430 1247 3440
rect 1261 3430 4631 3440
rect 4645 3430 8495 3440
rect 8509 3430 11039 3440
rect 11053 3430 12143 3440
rect -11123 3406 -6145 3416
rect -6131 3406 -4225 3416
rect -4211 3406 -3769 3416
rect -3755 3406 -2281 3416
rect -2267 3406 -2161 3416
rect -2147 3406 7031 3416
rect 7045 3406 7271 3416
rect 7285 3406 9959 3416
rect 10093 3406 10103 3416
rect 11413 3406 11687 3416
rect -11123 3382 6359 3392
rect 6517 3382 12335 3392
rect -11195 3358 -10729 3368
rect -10715 3358 -3361 3368
rect -3347 3358 -1777 3368
rect -1763 3358 -769 3368
rect -707 3358 7295 3368
rect 7309 3358 11159 3368
rect -11315 3334 -10849 3344
rect -10835 3334 -8473 3344
rect -8459 3334 7799 3344
rect 9253 3334 9455 3344
rect -11411 3310 -2521 3320
rect -2507 3310 -817 3320
rect -467 3310 4559 3320
rect 4573 3310 8855 3320
rect 8869 3310 10031 3320
rect 10045 3310 10799 3320
rect -11459 3286 -9049 3296
rect -9035 3286 1367 3296
rect 1429 3286 4475 3296
rect 4489 3286 5447 3296
rect 5461 3286 10391 3296
rect -11483 3262 -3889 3272
rect -3875 3262 10607 3272
rect -11555 3238 -6097 3248
rect -6083 3238 6167 3248
rect 6181 3238 7463 3248
rect -11603 3214 -8521 3224
rect -8507 3214 5231 3224
rect 5893 3214 8543 3224
rect -11675 3190 -3577 3200
rect -3299 3190 -3169 3200
rect -3059 3190 10415 3200
rect -11819 3166 2807 3176
rect 2917 3166 5519 3176
rect 6181 3166 6239 3176
rect 6373 3166 6527 3176
rect 6853 3166 7199 3176
rect -11843 3142 -8761 3152
rect -8531 3142 -1873 3152
rect -1859 3142 671 3152
rect 685 3142 4055 3152
rect 4069 3142 7535 3152
rect 7549 3142 9167 3152
rect 9181 3142 11675 3152
rect -11891 3118 -7489 3128
rect -7403 3118 5351 3128
rect -11939 3094 -11233 3104
rect -11219 3094 -10489 3104
rect -10475 3094 -10441 3104
rect -10427 3094 -6121 3104
rect -6107 3094 -4105 3104
rect -4091 3094 -1849 3104
rect -1835 3094 2375 3104
rect 2389 3094 2495 3104
rect 2509 3094 2783 3104
rect 2797 3094 3263 3104
rect 3277 3094 4103 3104
rect 4117 3094 4367 3104
rect 4381 3094 5495 3104
rect 5509 3094 7559 3104
rect 7573 3094 9863 3104
rect 9877 3094 10991 3104
rect -11963 3070 -8041 3080
rect -8027 3070 5759 3080
rect -11963 3046 1655 3056
rect 2389 3046 2447 3056
rect 2677 3046 2687 3056
rect 2749 3046 2951 3056
rect 4117 3046 4223 3056
rect 4453 3046 11927 3056
rect -12011 3022 -8641 3032
rect -8627 3022 -4225 3032
rect -4211 3022 -361 3032
rect -347 3022 4247 3032
rect 5245 3022 5615 3032
rect -12011 2998 -11809 3008
rect -11723 2998 -4273 3008
rect -4115 2998 6095 3008
rect 6109 2998 9839 3008
rect -12035 2974 -11377 2984
rect -11363 2974 -5929 2984
rect -5915 2974 1271 2984
rect 1285 2974 3815 2984
rect 3829 2974 11735 2984
rect -12035 2950 7055 2960
rect -12059 2926 -8353 2936
rect -8339 2926 -8281 2936
rect -8267 2926 -4657 2936
rect -4643 2926 -2977 2936
rect -2963 2926 -2809 2936
rect -2795 2926 5471 2936
rect 5485 2926 9719 2936
rect 9733 2926 10655 2936
rect 10669 2926 11615 2936
rect 11629 2926 11927 2936
rect 11941 2926 12167 2936
rect -12099 2902 -5833 2912
rect -5819 2902 8783 2912
rect 11629 2902 11675 2912
rect -12099 2878 -3529 2888
rect -2987 2878 2591 2888
rect 2605 2878 8591 2888
rect -12059 2854 -7273 2864
rect -7259 2854 -5281 2864
rect -5267 2854 -5113 2864
rect -5099 2854 2279 2864
rect 2293 2854 5951 2864
rect 7069 2854 7223 2864
rect -11915 2830 -11041 2840
rect -11027 2830 -2233 2840
rect -2219 2830 -2065 2840
rect -2051 2830 4007 2840
rect 4021 2830 5015 2840
rect 5029 2830 5303 2840
rect 5317 2830 11039 2840
rect -11891 2806 -11257 2816
rect -11243 2806 -10921 2816
rect -10907 2806 -9337 2816
rect -9323 2806 -8713 2816
rect -8699 2806 -8449 2816
rect -8435 2806 4079 2816
rect 4093 2806 6071 2816
rect 6085 2806 6575 2816
rect 6589 2806 7919 2816
rect 7933 2806 11135 2816
rect 11149 2806 11639 2816
rect -11843 2782 -11161 2792
rect -11147 2782 5207 2792
rect 5485 2782 5651 2792
rect -11771 2758 -6049 2768
rect -5987 2758 9023 2768
rect -11315 2734 -9481 2744
rect -9467 2734 -8377 2744
rect -8363 2734 -4633 2744
rect -4619 2734 -4297 2744
rect -4283 2734 -1297 2744
rect -1283 2734 -529 2744
rect -515 2734 95 2744
rect 109 2734 3119 2744
rect 3133 2734 5687 2744
rect 5701 2734 5927 2744
rect 5941 2734 7583 2744
rect 7597 2734 11759 2744
rect 11773 2734 12215 2744
rect -11147 2710 -10297 2720
rect -10283 2710 -8809 2720
rect -8795 2710 -7345 2720
rect -7331 2710 3359 2720
rect 3373 2710 4415 2720
rect 4429 2710 5639 2720
rect 5653 2710 6479 2720
rect 6493 2710 6551 2720
rect 6565 2710 9119 2720
rect 9133 2710 9743 2720
rect 9757 2710 11183 2720
rect 11773 2710 12263 2720
rect -11075 2686 6047 2696
rect 6061 2686 10511 2696
rect -11051 2662 -7369 2672
rect -7355 2662 2639 2672
rect 2653 2662 3023 2672
rect 6061 2662 6119 2672
rect 6565 2662 6599 2672
rect 9037 2662 9335 2672
rect -11003 2638 5183 2648
rect 5197 2638 11303 2648
rect -10955 2614 -7993 2624
rect -7979 2614 3527 2624
rect 5197 2614 11447 2624
rect -10931 2590 -10393 2600
rect -10379 2590 -3865 2600
rect -3851 2590 5159 2600
rect 5173 2590 5927 2600
rect 9133 2590 9431 2600
rect -10715 2566 2471 2576
rect 2485 2566 5999 2576
rect -10667 2542 -289 2552
rect -275 2542 10943 2552
rect -10595 2518 -1945 2528
rect -1931 2518 10823 2528
rect 10837 2518 11711 2528
rect 11725 2518 12167 2528
rect -10571 2494 -8593 2504
rect -8579 2494 -5689 2504
rect -5675 2494 -2641 2504
rect -2627 2494 -217 2504
rect -203 2494 527 2504
rect 541 2494 8351 2504
rect 8365 2494 10559 2504
rect -10499 2470 -10009 2480
rect -9995 2470 719 2480
rect 733 2470 5399 2480
rect 5413 2470 5735 2480
rect 8365 2470 8927 2480
rect -10451 2446 1367 2456
rect 1381 2446 7007 2456
rect 7021 2446 8591 2456
rect -10379 2422 -7441 2432
rect -7427 2422 -4081 2432
rect -4067 2422 -3193 2432
rect -3179 2422 -649 2432
rect -635 2422 1343 2432
rect 1357 2422 2879 2432
rect 2893 2422 6023 2432
rect 6037 2422 7439 2432
rect 7453 2422 9719 2432
rect -10235 2398 4319 2408
rect 5413 2398 5903 2408
rect -10211 2374 6623 2384
rect -10163 2350 2879 2360
rect -9731 2326 -3865 2336
rect -3851 2326 -3217 2336
rect -3203 2326 -2713 2336
rect -2699 2326 1319 2336
rect 2485 2326 2567 2336
rect 2845 2326 9791 2336
rect -9587 2302 -6577 2312
rect -6563 2302 -457 2312
rect -443 2302 3623 2312
rect 3637 2302 8879 2312
rect -9563 2278 -1561 2288
rect -1547 2278 3551 2288
rect -9515 2254 10007 2264
rect -9395 2230 -8929 2240
rect -8867 2230 -841 2240
rect -515 2230 -397 2240
rect -347 2230 -265 2240
rect -203 2230 -25 2240
rect 37 2230 3143 2240
rect -9371 2206 -7681 2216
rect -7667 2206 -3913 2216
rect -3899 2206 2303 2216
rect 2317 2206 5855 2216
rect 5869 2206 7103 2216
rect -9347 2182 -9169 2192
rect -9155 2182 -3817 2192
rect -3803 2182 -3769 2192
rect -3755 2182 -2593 2192
rect -2579 2182 -553 2192
rect -539 2182 4151 2192
rect 4165 2182 5711 2192
rect 5725 2182 8279 2192
rect 8293 2182 8759 2192
rect -9323 2158 -7825 2168
rect -7811 2158 3551 2168
rect 3565 2158 5975 2168
rect -9251 2134 -8785 2144
rect -8771 2134 -4201 2144
rect -4187 2134 -2137 2144
rect -2123 2134 5375 2144
rect 5389 2134 5543 2144
rect 5557 2134 5831 2144
rect -8819 2110 -5545 2120
rect -5531 2110 -4729 2120
rect -4715 2110 2159 2120
rect -8435 2086 -1657 2096
rect -1403 2086 2543 2096
rect -8411 2062 3719 2072
rect -8387 2038 -577 2048
rect -563 2038 5279 2048
rect 5293 2038 11951 2048
rect -8363 2014 -7321 2024
rect -7307 2014 -5593 2024
rect -5579 2014 -3289 2024
rect -3275 2014 -1753 2024
rect -1739 2014 8207 2024
rect 8221 2014 10487 2024
rect 10501 2014 11207 2024
rect -8339 1990 -1153 2000
rect -899 1990 11375 2000
rect -8099 1966 -7681 1976
rect -7619 1966 -3841 1976
rect -3611 1966 -505 1976
rect -491 1966 3863 1976
rect 3877 1966 7415 1976
rect 7429 1966 9215 1976
rect 9229 1966 9815 1976
rect -7859 1942 6887 1952
rect -7811 1918 -6241 1928
rect -6227 1918 -433 1928
rect -323 1918 -193 1928
rect 181 1918 5327 1928
rect -7571 1894 5423 1904
rect -7523 1870 3095 1880
rect 5293 1870 5783 1880
rect -7355 1846 -4465 1856
rect -4451 1846 215 1856
rect 445 1846 7247 1856
rect 7261 1846 12287 1856
rect -7307 1822 1223 1832
rect -7187 1798 11111 1808
rect -7091 1774 -2833 1784
rect -2459 1774 8735 1784
rect 8749 1774 11555 1784
rect -7043 1750 -7033 1760
rect -6971 1750 6791 1760
rect 6805 1750 11783 1760
rect -6995 1726 10031 1736
rect 11797 1726 12491 1736
rect -6947 1702 2639 1712
rect -6755 1678 -6625 1688
rect -6563 1678 -5137 1688
rect -5123 1678 -2089 1688
rect -2075 1678 8567 1688
rect 8581 1678 8999 1688
rect -6707 1654 -6313 1664
rect -6299 1654 -5377 1664
rect -5363 1654 -3097 1664
rect -3083 1654 1319 1664
rect 1333 1654 2759 1664
rect 2773 1654 4175 1664
rect 9013 1654 9287 1664
rect -6683 1630 -5257 1640
rect -5243 1630 -3985 1640
rect -3971 1630 4583 1640
rect 4597 1630 11063 1640
rect -6491 1606 -6265 1616
rect -6251 1606 -3457 1616
rect -3443 1606 -3049 1616
rect -2435 1606 3791 1616
rect 4189 1606 4475 1616
rect -6347 1582 -6289 1592
rect -6203 1582 407 1592
rect 469 1582 11807 1592
rect -6299 1558 -3025 1568
rect -2387 1558 11975 1568
rect -6155 1534 71 1544
rect 805 1534 6311 1544
rect 11989 1534 12695 1544
rect -6083 1510 3935 1520
rect 3949 1510 4535 1520
rect 6325 1510 8663 1520
rect -5915 1486 -5893 1496
rect -5843 1486 9263 1496
rect -5867 1462 4751 1472
rect -5771 1438 -5761 1448
rect -5699 1438 -4873 1448
rect -4859 1438 2231 1448
rect -5675 1414 7967 1424
rect -5363 1390 -865 1400
rect -851 1390 359 1400
rect 373 1390 5711 1400
rect 5725 1390 6263 1400
rect 6277 1390 10247 1400
rect -5339 1366 12719 1376
rect -5147 1342 -1609 1352
rect -1115 1342 8831 1352
rect -5099 1318 -5065 1328
rect -5003 1318 -2353 1328
rect -2267 1318 -2041 1328
rect -1715 1318 4367 1328
rect 6277 1318 6419 1328
rect -4931 1294 6335 1304
rect 6349 1294 8687 1304
rect -4835 1270 -2929 1280
rect -2915 1270 -169 1280
rect -155 1270 -121 1280
rect -107 1270 5087 1280
rect 5101 1270 8807 1280
rect 8821 1270 10367 1280
rect 10381 1270 11207 1280
rect -4451 1246 6719 1256
rect -4403 1222 695 1232
rect 853 1222 7631 1232
rect -4187 1198 -4057 1208
rect -3923 1198 4295 1208
rect -4067 1174 9695 1184
rect -3539 1150 11903 1160
rect -3179 1126 -3121 1136
rect -2315 1126 7511 1136
rect -2027 1102 3839 1112
rect -827 1078 -601 1088
rect -227 1078 -49 1088
rect 1045 1078 1295 1088
rect 2245 1078 2327 1088
rect 12781 1078 12838 1088
rect -155 1054 2399 1064
rect 2413 1054 6191 1064
rect 12757 1054 12838 1064
rect -12183 964 -12096 989
rect -12183 -799 -12133 964
rect 12872 344 12922 6096
rect 12432 319 12922 344
rect -419 221 3047 231
rect -803 197 -25 207
rect 829 197 11567 207
rect -1019 173 2399 183
rect 2869 173 7223 183
rect -1067 149 2183 159
rect 2197 149 3023 159
rect 3037 149 7871 159
rect -3779 125 3983 135
rect -5891 101 -5881 111
rect -5627 101 -409 111
rect 781 101 3671 111
rect -5891 77 11543 87
rect -6179 53 -961 63
rect -947 53 2999 63
rect -6323 29 3143 39
rect -6371 5 -4297 15
rect -3995 5 -3601 15
rect -1451 5 503 15
rect 589 5 1943 15
rect 2797 5 8063 15
rect -6539 -19 -5185 -9
rect -5171 -19 -3361 -9
rect -3347 -19 -289 -9
rect 349 -19 3479 -9
rect -6659 -43 -4345 -33
rect -4019 -43 6407 -33
rect 6589 -43 7991 -33
rect -6779 -67 -3529 -57
rect -2339 -67 551 -57
rect 613 -67 911 -57
rect 1021 -67 2927 -57
rect 5341 -67 10943 -57
rect -6947 -91 -4561 -81
rect -4355 -91 -3721 -81
rect -3467 -91 -385 -81
rect -251 -91 7727 -81
rect -7043 -115 3575 -105
rect 3781 -115 10103 -105
rect -7139 -139 8543 -129
rect 8821 -139 9959 -129
rect -7403 -163 2615 -153
rect 2773 -163 10607 -153
rect -7523 -187 8855 -177
rect -7547 -211 -2881 -201
rect -2771 -211 5375 -201
rect 5437 -211 10247 -201
rect -7595 -235 -7225 -225
rect -7163 -235 119 -225
rect 325 -235 9143 -225
rect 9925 -237 9943 -223
rect 12421 -235 12455 -225
rect -8699 -259 2327 -249
rect 2701 -259 12838 -249
rect -8723 -283 3287 -273
rect 3397 -283 9983 -273
rect 12373 -283 12431 -273
rect -8771 -307 -5881 -297
rect -5867 -307 3815 -297
rect 3829 -307 7199 -297
rect 7213 -307 9071 -297
rect -9011 -331 8423 -321
rect -9035 -355 7415 -345
rect -9107 -379 -6937 -369
rect -6875 -379 12407 -369
rect -9131 -403 8639 -393
rect 8653 -403 8735 -393
rect 8749 -403 11231 -393
rect -9203 -427 -4729 -417
rect -4307 -427 -2209 -417
rect -1163 -427 11159 -417
rect -9227 -451 11687 -441
rect -9299 -475 -4921 -465
rect -4691 -475 3335 -465
rect -9491 -499 -8689 -489
rect -7667 -499 335 -489
rect 1405 -499 2135 -489
rect 2149 -499 8183 -489
rect -9539 -523 -49 -513
rect 1549 -523 4967 -513
rect -10139 -547 959 -537
rect -10259 -571 287 -561
rect -10307 -595 -3145 -585
rect -3131 -595 407 -585
rect 421 -595 9191 -585
rect -10355 -619 -4489 -609
rect -3971 -619 5759 -609
rect -10403 -643 -2569 -633
rect -2555 -643 6383 -633
rect 6397 -643 10799 -633
rect -10547 -667 -4441 -657
rect -3827 -667 887 -657
rect -10691 -691 8903 -681
rect -11171 -715 7631 -705
rect -12099 -739 -11977 -729
rect -11723 -739 -7129 -729
rect -7067 -739 -5065 -729
rect -5051 -739 7511 -729
rect 12469 -739 12838 -729
rect -12099 -763 -10849 -753
rect -10787 -763 4559 -753
rect 12445 -763 12838 -753
rect -6611 -787 -5869 -777
rect -5411 -787 263 -777
rect 12421 -787 12838 -777
rect 12872 -799 12922 319
<< m2contact >>
rect -433 7141 -419 7155
rect 10115 7141 10129 7155
rect -3265 7117 -3251 7131
rect -2377 7117 -2363 7131
rect -1513 7117 -1499 7131
rect 9299 7117 9313 7131
rect -4609 7093 -4595 7107
rect 1955 7093 1969 7107
rect 6827 7093 6841 7107
rect 6959 7093 6973 7107
rect 7643 7093 7657 7107
rect 8159 7093 8173 7107
rect -10417 7069 -10403 7083
rect -8449 7069 -8435 7083
rect -6289 7069 -6275 7083
rect -4801 7069 -4787 7083
rect -1321 7069 -1307 7083
rect -817 7069 -803 7083
rect 1139 7069 1153 7083
rect 3563 7069 3577 7083
rect 3695 7069 3709 7083
rect 4295 7069 4309 7083
rect 6287 7069 6301 7083
rect 12815 7069 12829 7083
rect -10825 7045 -10811 7059
rect -10441 7045 -10427 7059
rect -9601 7045 -9587 7059
rect -8593 7045 -8579 7059
rect -7117 7045 -7103 7059
rect -7057 7045 -7043 7059
rect -2149 7045 -2135 7059
rect -1657 7045 -1643 7059
rect 4403 7045 4417 7059
rect 6011 7045 6025 7059
rect 9431 7045 9445 7059
rect -12113 7021 -12099 7035
rect -6361 7021 -6347 7035
rect -5065 7021 -5051 7035
rect 7667 7021 7681 7035
rect -12113 6997 -12099 7011
rect 1943 6997 1957 7011
rect 3551 6997 3565 7011
rect 12743 6997 12757 7011
rect -11377 6973 -11345 6987
rect -9265 6973 -9251 6987
rect -913 6973 -899 6987
rect 5591 6973 5605 6987
rect 12047 6973 12061 6987
rect 12719 6973 12733 6987
rect 12767 6973 12781 6987
rect -7981 6949 -7967 6963
rect -7345 6949 -7331 6963
rect -7153 6949 -7139 6963
rect -4729 6949 -4715 6963
rect -4669 6949 -4655 6963
rect 11879 6949 11893 6963
rect -6553 6925 -6539 6939
rect 455 6925 469 6939
rect 6863 6925 6877 6939
rect 10931 6925 10945 6939
rect 12743 6925 12757 6939
rect 12838 6925 12852 6939
rect -3841 6901 -3827 6915
rect 7199 6901 7213 6915
rect 8015 6901 8029 6915
rect 8483 6901 8497 6915
rect 8927 6901 8941 6915
rect 11747 6901 11761 6915
rect 12791 6901 12805 6915
rect 12838 6901 12852 6915
rect -601 6877 -587 6891
rect 12743 6877 12757 6891
rect 12767 6877 12781 6891
rect 12838 6877 12852 6891
rect 299 6853 313 6867
rect 11327 6853 11341 6867
rect 12743 6853 12757 6867
rect 12838 6853 12852 6867
rect 1115 6829 1129 6843
rect 8735 6829 8749 6843
rect 10271 6829 10285 6843
rect 12791 6829 12805 6843
rect 12815 6829 12829 6843
rect 12838 6829 12852 6843
rect 7391 5996 7405 6010
rect 8783 5996 8797 6010
rect -1681 5972 -1667 5986
rect 10967 5972 10981 5986
rect -1993 5948 -1979 5962
rect -1033 5948 -1019 5962
rect 5615 5948 5629 5962
rect 6455 5948 6469 5962
rect 7487 5948 7501 5962
rect 11687 5948 11701 5962
rect -2041 5924 -2027 5938
rect 11327 5924 11341 5938
rect -2089 5900 -2075 5914
rect 2327 5900 2341 5914
rect 2423 5900 2437 5914
rect 7391 5900 7405 5914
rect 12263 5900 12277 5914
rect -2377 5876 -2363 5890
rect -2353 5876 -2339 5890
rect -2209 5876 -2195 5890
rect 2423 5876 2437 5890
rect -3433 5852 -3419 5866
rect -1993 5852 -1979 5866
rect -1825 5852 -1811 5866
rect 10151 5852 10165 5866
rect -3889 5828 -3875 5842
rect -3817 5828 -3803 5842
rect -3697 5828 -3683 5842
rect 10199 5828 10213 5842
rect -3961 5804 -3947 5818
rect 5255 5804 5269 5818
rect -4057 5780 -4043 5794
rect 1631 5780 1645 5794
rect -4417 5756 -4403 5770
rect 1871 5756 1885 5770
rect -4513 5732 -4499 5746
rect -3409 5732 -3395 5746
rect -3001 5732 -2987 5746
rect -97 5732 -83 5746
rect 1079 5732 1093 5746
rect 4271 5732 4285 5746
rect 4391 5732 4405 5746
rect 6695 5732 6709 5746
rect 8183 5732 8197 5746
rect 10103 5732 10117 5746
rect 10583 5732 10597 5746
rect -4633 5708 -4619 5722
rect -3121 5708 -3107 5722
rect 2687 5708 2701 5722
rect 11879 5708 11893 5722
rect -4729 5684 -4715 5698
rect -3673 5684 -3659 5698
rect 2351 5684 2365 5698
rect 2999 5684 3013 5698
rect 4343 5684 4357 5698
rect 5591 5684 5605 5698
rect 6791 5684 6805 5698
rect -4897 5660 -4883 5674
rect -4801 5660 -4787 5674
rect -4753 5660 -4739 5674
rect -4729 5660 -4715 5674
rect -4657 5660 -4643 5674
rect -769 5660 -755 5674
rect 6215 5660 6229 5674
rect 6335 5660 6349 5674
rect -4969 5636 -4955 5650
rect 1487 5636 1501 5650
rect 5135 5636 5149 5650
rect 8975 5636 8989 5650
rect -4993 5612 -4979 5626
rect 9887 5612 9901 5626
rect -5233 5588 -5219 5602
rect 12455 5588 12469 5602
rect -5233 5564 -5219 5578
rect 10871 5564 10885 5578
rect -5329 5540 -5315 5554
rect -49 5540 -35 5554
rect 4727 5540 4741 5554
rect 11999 5540 12013 5554
rect -5449 5516 -5435 5530
rect -1273 5516 -1259 5530
rect -1225 5516 -1211 5530
rect 12838 5516 12852 5530
rect -5593 5492 -5579 5506
rect -5329 5492 -5315 5506
rect -5281 5492 -5267 5506
rect 10751 5492 10765 5506
rect 11231 5492 11245 5506
rect -5617 5468 -5603 5482
rect -409 5468 -395 5482
rect 4463 5468 4477 5482
rect 8231 5468 8245 5482
rect 9479 5468 9493 5482
rect -5665 5444 -5651 5458
rect 6671 5444 6685 5458
rect 11423 5444 11437 5458
rect 11903 5444 11917 5458
rect -5761 5420 -5747 5434
rect 6527 5420 6541 5434
rect 10919 5420 10933 5434
rect 11807 5420 11821 5434
rect -6001 5396 -5987 5410
rect -5761 5396 -5747 5410
rect -5713 5396 -5699 5410
rect -2689 5396 -2675 5410
rect 935 5396 949 5410
rect 2063 5396 2077 5410
rect 6671 5396 6685 5410
rect 8519 5396 8533 5410
rect 10919 5396 10933 5410
rect 11423 5396 11437 5410
rect -6073 5372 -6059 5386
rect 11279 5372 11293 5386
rect -6121 5348 -6107 5362
rect -193 5348 -179 5362
rect 4247 5348 4261 5362
rect 9239 5348 9253 5362
rect -6193 5324 -6179 5338
rect -5977 5324 -5963 5338
rect -5905 5324 -5891 5338
rect 6215 5324 6229 5338
rect -6217 5300 -6203 5314
rect 1847 5300 1861 5314
rect 6743 5300 6757 5314
rect 7151 5300 7165 5314
rect 7367 5300 7381 5314
rect 7511 5300 7525 5314
rect 9767 5300 9781 5314
rect 9791 5300 9805 5314
rect -6409 5276 -6395 5290
rect 1439 5276 1453 5290
rect 2303 5276 2317 5290
rect 2399 5276 2413 5290
rect 4127 5276 4141 5290
rect 9935 5276 9949 5290
rect -6481 5252 -6467 5266
rect -5893 5252 -5879 5266
rect -5785 5252 -5771 5266
rect -5473 5252 -5459 5266
rect -5017 5252 -5003 5266
rect -4057 5252 -4043 5266
rect -2737 5252 -2723 5266
rect -2665 5252 -2651 5266
rect -2545 5252 -2531 5266
rect 2951 5252 2965 5266
rect 4199 5252 4213 5266
rect 7151 5252 7165 5266
rect 9287 5252 9301 5266
rect 9767 5252 9781 5266
rect 11951 5252 11965 5266
rect -6481 5228 -6467 5242
rect 8159 5228 8173 5242
rect -6529 5204 -6515 5218
rect 9575 5204 9589 5218
rect -6529 5180 -6515 5194
rect -1369 5180 -1355 5194
rect -1297 5180 -1283 5194
rect 1079 5180 1093 5194
rect 2183 5180 2197 5194
rect 6455 5180 6469 5194
rect 9359 5180 9373 5194
rect 9455 5180 9469 5194
rect -6625 5156 -6611 5170
rect 12767 5156 12781 5170
rect -6649 5132 -6635 5146
rect -2617 5132 -2603 5146
rect -2377 5132 -2363 5146
rect 191 5132 205 5146
rect 2087 5132 2101 5146
rect 9359 5132 9373 5146
rect -6673 5108 -6659 5122
rect 8471 5108 8485 5122
rect -6697 5084 -6683 5098
rect 3767 5084 3781 5098
rect 8111 5084 8125 5098
rect -6745 5060 -6731 5074
rect -1 5060 13 5074
rect 2039 5060 2053 5074
rect 10847 5060 10861 5074
rect -6841 5036 -6827 5050
rect 1559 5036 1573 5050
rect 2015 5036 2029 5050
rect 3935 5036 3949 5050
rect 3983 5036 3997 5050
rect 4967 5036 4981 5050
rect 6623 5036 6637 5050
rect 11471 5036 11485 5050
rect 12119 5036 12133 5050
rect -6913 5012 -6899 5026
rect -4273 5012 -4259 5026
rect -4153 5012 -4139 5026
rect -3433 5012 -3419 5026
rect -3265 5012 -3251 5026
rect -25 5012 -11 5026
rect 1919 5012 1933 5026
rect 12239 5012 12253 5026
rect -7129 4988 -7115 5002
rect -1249 4988 -1235 5002
rect 8039 4988 8053 5002
rect 11471 4988 11485 5002
rect -7153 4964 -7139 4978
rect -4513 4964 -4499 4978
rect 12479 4964 12493 4978
rect -7225 4940 -7211 4954
rect 7295 4940 7309 4954
rect -7345 4916 -7331 4930
rect -7321 4916 -7307 4930
rect -7249 4916 -7235 4930
rect 8279 4916 8293 4930
rect -7465 4892 -7451 4906
rect -4321 4892 -4307 4906
rect -2785 4892 -2771 4906
rect 10655 4892 10669 4906
rect 11663 4892 11677 4906
rect 11735 4892 11749 4906
rect -7465 4868 -7451 4882
rect 12383 4868 12397 4882
rect -7633 4844 -7619 4858
rect 3239 4844 3253 4858
rect 5135 4844 5149 4858
rect 12047 4844 12061 4858
rect -7753 4820 -7739 4834
rect -3793 4820 -3779 4834
rect -3745 4820 -3731 4834
rect -1201 4820 -1187 4834
rect 1895 4820 1909 4834
rect 4799 4820 4813 4834
rect 4847 4820 4861 4834
rect 7031 4820 7045 4834
rect 7319 4820 7333 4834
rect 8711 4820 8725 4834
rect 8735 4820 8749 4834
rect -7897 4796 -7883 4810
rect -4705 4796 -4691 4810
rect 12239 4796 12253 4810
rect -7921 4772 -7907 4786
rect 4031 4772 4045 4786
rect 4079 4772 4093 4786
rect 6119 4772 6133 4786
rect 6983 4772 6997 4786
rect 12695 4772 12709 4786
rect -8089 4748 -8075 4762
rect -5569 4748 -5555 4762
rect -5449 4748 -5435 4762
rect 9527 4748 9541 4762
rect -8209 4724 -8195 4738
rect -6817 4724 -6803 4738
rect -2185 4724 -2171 4738
rect -1129 4724 -1115 4738
rect 2207 4724 2221 4738
rect 2255 4724 2269 4738
rect 3191 4724 3205 4738
rect 6287 4724 6301 4738
rect 8711 4724 8725 4738
rect -8233 4700 -8219 4714
rect -6889 4700 -6875 4714
rect -4825 4700 -4811 4714
rect -4609 4700 -4595 4714
rect 8231 4700 8245 4714
rect -8233 4676 -8219 4690
rect -5545 4676 -5531 4690
rect -5497 4676 -5483 4690
rect 2663 4676 2677 4690
rect 3743 4676 3757 4690
rect 9335 4676 9349 4690
rect -8257 4652 -8243 4666
rect -7705 4652 -7691 4666
rect -5401 4652 -5387 4666
rect -5161 4652 -5147 4666
rect -3145 4652 -3131 4666
rect -2761 4652 -2747 4666
rect -241 4652 -227 4666
rect 2735 4652 2749 4666
rect 2927 4652 2941 4666
rect 3887 4652 3901 4666
rect 12431 4652 12445 4666
rect -8329 4628 -8315 4642
rect 5903 4628 5917 4642
rect 6599 4628 6613 4642
rect -8785 4604 -8771 4618
rect -5353 4604 -5339 4618
rect -4537 4604 -4523 4618
rect -2305 4604 -2291 4618
rect 647 4604 661 4618
rect 2711 4604 2725 4618
rect 5975 4604 5989 4618
rect 10079 4604 10093 4618
rect -8809 4580 -8795 4594
rect -8785 4580 -8771 4594
rect -8665 4580 -8651 4594
rect -625 4580 -611 4594
rect -397 4580 -383 4594
rect 6383 4580 6397 4594
rect 7223 4580 7237 4594
rect 7367 4580 7381 4594
rect 9431 4580 9445 4594
rect 11855 4580 11869 4594
rect 12599 4580 12613 4594
rect -8881 4556 -8867 4570
rect -2641 4556 -2627 4570
rect 11855 4556 11869 4570
rect -8905 4532 -8891 4546
rect -505 4532 -491 4546
rect 1799 4532 1813 4546
rect 7679 4532 7693 4546
rect -8929 4508 -8915 4522
rect 4223 4508 4237 4522
rect 10175 4508 10189 4522
rect -8953 4484 -8939 4498
rect -8185 4484 -8171 4498
rect -8137 4484 -8123 4498
rect -6793 4484 -6779 4498
rect 11519 4484 11533 4498
rect 11543 4484 11557 4498
rect 12527 4484 12541 4498
rect -8977 4460 -8963 4474
rect 6815 4460 6829 4474
rect 6911 4460 6925 4474
rect 7079 4460 7093 4474
rect 7607 4460 7621 4474
rect 7631 4460 7645 4474
rect -9001 4436 -8987 4450
rect -6409 4436 -6395 4450
rect -6289 4436 -6275 4450
rect -337 4436 -323 4450
rect 4655 4436 4669 4450
rect 8327 4436 8341 4450
rect -9073 4412 -9059 4426
rect -3649 4412 -3635 4426
rect -3481 4412 -3467 4426
rect 1199 4412 1213 4426
rect 1751 4412 1765 4426
rect 11351 4412 11365 4426
rect -9097 4388 -9083 4402
rect -3961 4388 -3947 4402
rect -3601 4388 -3587 4402
rect -3553 4388 -3539 4402
rect 12095 4388 12109 4402
rect -9145 4364 -9131 4378
rect 8375 4364 8389 4378
rect -9169 4340 -9155 4354
rect 12191 4340 12205 4354
rect -9241 4316 -9227 4330
rect -6433 4316 -6419 4330
rect 10679 4316 10693 4330
rect -9313 4292 -9299 4306
rect -8593 4292 -8579 4306
rect 2975 4292 2989 4306
rect 3743 4292 3757 4306
rect 6143 4292 6157 4306
rect 7127 4292 7141 4306
rect 7607 4292 7621 4306
rect 8255 4292 8269 4306
rect 9503 4292 9517 4306
rect 11135 4292 11149 4306
rect -9433 4268 -9419 4282
rect -1441 4268 -1427 4282
rect -1321 4268 -1307 4282
rect -1153 4268 -1139 4282
rect -889 4268 -875 4282
rect -265 4268 -251 4282
rect 1583 4268 1597 4282
rect 11087 4268 11101 4282
rect -9457 4244 -9443 4258
rect -673 4244 -659 4258
rect 1511 4244 1525 4258
rect 8423 4244 8437 4258
rect -9481 4220 -9467 4234
rect -3241 4220 -3227 4234
rect -3049 4220 -3035 4234
rect -3025 4220 -3011 4234
rect -2713 4220 -2699 4234
rect -2593 4220 -2579 4234
rect -2473 4220 -2459 4234
rect -97 4220 -83 4234
rect 1463 4220 1477 4234
rect 9311 4220 9325 4234
rect -9553 4196 -9539 4210
rect -7873 4196 -7859 4210
rect -7777 4196 -7763 4210
rect -4177 4196 -4163 4210
rect -2905 4196 -2891 4210
rect 2111 4196 2125 4210
rect 5639 4196 5653 4210
rect 6935 4196 6949 4210
rect 11399 4196 11413 4210
rect -9625 4172 -9611 4186
rect -2857 4172 -2843 4186
rect 8303 4172 8317 4186
rect -9673 4148 -9659 4162
rect -3745 4148 -3731 4162
rect -2113 4148 -2099 4162
rect 2135 4148 2149 4162
rect 5879 4148 5893 4162
rect 6911 4148 6925 4162
rect 7487 4148 7501 4162
rect -9697 4124 -9683 4138
rect -7249 4124 -7235 4138
rect -2953 4124 -2939 4138
rect -145 4124 -131 4138
rect 1127 4124 1141 4138
rect 2087 4124 2101 4138
rect 4895 4124 4909 4138
rect 5807 4124 5821 4138
rect 12071 4124 12085 4138
rect -9937 4100 -9923 4114
rect -3385 4100 -3371 4114
rect -73 4100 -59 4114
rect 671 4100 685 4114
rect 695 4100 709 4114
rect 1271 4100 1285 4114
rect 1295 4100 1309 4114
rect 1415 4100 1429 4114
rect 10127 4100 10141 4114
rect -9985 4076 -9971 4090
rect -9817 4076 -9803 4090
rect 6479 4076 6493 4090
rect 10895 4076 10909 4090
rect 11447 4076 11461 4090
rect -10033 4052 -10019 4066
rect -9793 4052 -9779 4066
rect -6865 4052 -6851 4066
rect -6745 4052 -6731 4066
rect -6025 4052 -6011 4066
rect -4585 4052 -4571 4066
rect -4009 4052 -3995 4066
rect -2041 4052 -2027 4066
rect 7463 4052 7477 4066
rect 11015 4052 11029 4066
rect 12143 4052 12157 4066
rect -10081 4028 -10067 4042
rect 11831 4028 11845 4042
rect -10105 4004 -10091 4018
rect -6433 4004 -6419 4018
rect -4105 4004 -4091 4018
rect -1249 4004 -1235 4018
rect 10895 4004 10909 4018
rect -10129 3980 -10115 3994
rect -1009 3980 -995 3994
rect -937 3980 -923 3994
rect 3647 3980 3661 3994
rect 8015 3980 8029 3994
rect -10297 3956 -10283 3970
rect -3169 3956 -3155 3970
rect -3073 3956 -3059 3970
rect 5783 3956 5797 3970
rect -10321 3932 -10307 3946
rect -8497 3932 -8483 3946
rect -3673 3932 -3659 3946
rect -2137 3932 -2123 3946
rect 1175 3932 1189 3946
rect 1247 3932 1261 3946
rect 10703 3932 10717 3946
rect -10345 3908 -10331 3922
rect -3649 3908 -3635 3922
rect -3313 3908 -3299 3922
rect 9143 3908 9157 3922
rect 12311 3908 12325 3922
rect -10417 3884 -10403 3898
rect -5665 3884 -5651 3898
rect -1177 3884 -1163 3898
rect 5831 3884 5845 3898
rect 6239 3884 6253 3898
rect 7943 3884 7957 3898
rect 11495 3884 11509 3898
rect -10489 3860 -10475 3874
rect 1607 3860 1621 3874
rect 1703 3860 1717 3874
rect 5039 3860 5053 3874
rect 5111 3860 5125 3874
rect 5447 3860 5461 3874
rect 5495 3860 5509 3874
rect 6023 3860 6037 3874
rect -10513 3836 -10499 3850
rect -7801 3836 -7787 3850
rect -6457 3836 -6443 3850
rect -2617 3836 -2603 3850
rect -1321 3836 -1307 3850
rect -313 3836 -299 3850
rect 1031 3836 1045 3850
rect 2855 3836 2869 3850
rect 3215 3836 3229 3850
rect 5111 3836 5125 3850
rect 6695 3836 6709 3850
rect 7175 3836 7189 3850
rect 7343 3836 7357 3850
rect 8975 3836 8989 3850
rect 10343 3836 10357 3850
rect 11591 3836 11605 3850
rect 12071 3836 12085 3850
rect -10537 3812 -10523 3826
rect 6503 3812 6517 3826
rect 9623 3812 9637 3826
rect 12575 3812 12589 3826
rect -10585 3788 -10571 3802
rect 12359 3788 12373 3802
rect -10609 3764 -10595 3778
rect -7585 3764 -7571 3778
rect 4679 3764 4693 3778
rect 9047 3764 9061 3778
rect 12647 3764 12661 3778
rect -10633 3740 -10619 3754
rect -2833 3740 -2819 3754
rect 12623 3740 12637 3754
rect -10657 3716 -10643 3730
rect -4801 3716 -4787 3730
rect 2567 3716 2581 3730
rect 2615 3716 2629 3730
rect 6407 3716 6421 3730
rect 7271 3716 7285 3730
rect 7535 3716 7549 3730
rect 9191 3716 9205 3730
rect 9383 3716 9397 3730
rect 9599 3716 9613 3730
rect 10295 3716 10309 3730
rect -10657 3692 -10643 3706
rect 6959 3692 6973 3706
rect 7103 3692 7117 3706
rect 7415 3692 7429 3706
rect 9071 3692 9085 3706
rect 12838 3692 12852 3706
rect -10705 3668 -10691 3682
rect -4753 3668 -4739 3682
rect -721 3668 -707 3682
rect 47 3668 61 3682
rect 9647 3668 9661 3682
rect 9983 3668 9997 3682
rect 10775 3668 10789 3682
rect -10753 3644 -10739 3658
rect -5473 3644 -5459 3658
rect 4991 3644 5005 3658
rect 6095 3644 6109 3658
rect 8399 3644 8413 3658
rect 8615 3644 8629 3658
rect 12743 3644 12757 3658
rect -10801 3620 -10787 3634
rect -6841 3620 -6827 3634
rect -4921 3620 -4907 3634
rect 2447 3620 2461 3634
rect 2591 3620 2605 3634
rect 12491 3620 12505 3634
rect -10825 3596 -10811 3610
rect -961 3596 -947 3610
rect 5567 3596 5581 3610
rect 7823 3596 7837 3610
rect 12023 3596 12037 3610
rect -10897 3572 -10883 3586
rect 1727 3572 1741 3586
rect 1775 3572 1789 3586
rect 11255 3572 11269 3586
rect -10897 3548 -10883 3562
rect 3695 3548 3709 3562
rect 3911 3548 3925 3562
rect 10823 3548 10837 3562
rect 11303 3548 11317 3562
rect 11555 3548 11569 3562
rect -10945 3524 -10931 3538
rect -9889 3524 -9875 3538
rect -9577 3524 -9563 3538
rect -4561 3524 -4547 3538
rect -2881 3524 -2867 3538
rect 1151 3524 1165 3538
rect 3431 3524 3445 3538
rect 5651 3524 5665 3538
rect 6767 3524 6781 3538
rect 9095 3524 9109 3538
rect 10463 3524 10477 3538
rect 11831 3524 11845 3538
rect 12407 3524 12421 3538
rect 12671 3524 12685 3538
rect -10969 3500 -10955 3514
rect -7297 3500 -7283 3514
rect 3455 3500 3469 3514
rect 4199 3500 4213 3514
rect 12599 3500 12613 3514
rect -11017 3476 -11003 3490
rect -5809 3476 -5795 3490
rect -1057 3476 -1043 3490
rect -937 3476 -923 3490
rect 2975 3476 2989 3490
rect 7079 3476 7093 3490
rect 8159 3476 8173 3490
rect 8183 3476 8197 3490
rect 8447 3476 8461 3490
rect 9407 3476 9421 3490
rect 9911 3476 9925 3490
rect 12551 3476 12565 3490
rect -11065 3452 -11051 3466
rect -9769 3452 -9755 3466
rect -4345 3452 -4331 3466
rect -4177 3452 -4163 3466
rect 1991 3452 2005 3466
rect 2519 3452 2533 3466
rect 6419 3452 6433 3466
rect 12119 3452 12133 3466
rect -11113 3428 -11099 3442
rect -5257 3428 -5243 3442
rect -5185 3428 -5171 3442
rect -2929 3428 -2915 3442
rect -2521 3428 -2507 3442
rect -2257 3428 -2243 3442
rect 1247 3428 1261 3442
rect 4631 3428 4645 3442
rect 8495 3428 8509 3442
rect 11039 3428 11053 3442
rect 12143 3428 12157 3442
rect -11137 3404 -11123 3418
rect -6145 3404 -6131 3418
rect -4225 3404 -4211 3418
rect -3769 3404 -3755 3418
rect -2281 3404 -2267 3418
rect -2161 3404 -2147 3418
rect 7031 3404 7045 3418
rect 7271 3404 7285 3418
rect 9959 3404 9973 3418
rect 10079 3404 10093 3418
rect 10103 3404 10117 3418
rect 11399 3404 11413 3418
rect 11687 3404 11701 3418
rect -11137 3380 -11123 3394
rect 6359 3380 6373 3394
rect 6503 3380 6517 3394
rect 12335 3380 12349 3394
rect -11209 3356 -11195 3370
rect -10729 3356 -10715 3370
rect -3361 3356 -3347 3370
rect -1777 3356 -1763 3370
rect -769 3356 -755 3370
rect -721 3356 -707 3370
rect 7295 3356 7309 3370
rect 11159 3356 11173 3370
rect -11329 3332 -11315 3346
rect -10849 3332 -10835 3346
rect -8473 3332 -8459 3346
rect 7799 3332 7813 3346
rect 9239 3332 9253 3346
rect 9455 3332 9469 3346
rect -11425 3308 -11411 3322
rect -2521 3308 -2507 3322
rect -817 3308 -803 3322
rect -481 3308 -467 3322
rect 4559 3308 4573 3322
rect 8855 3308 8869 3322
rect 10031 3308 10045 3322
rect 10799 3308 10813 3322
rect -11473 3284 -11459 3298
rect -9049 3284 -9035 3298
rect 1367 3284 1381 3298
rect 1415 3284 1429 3298
rect 4475 3284 4489 3298
rect 5447 3284 5461 3298
rect 10391 3284 10405 3298
rect -11497 3260 -11483 3274
rect -3889 3260 -3875 3274
rect 10607 3260 10621 3274
rect -11569 3236 -11555 3250
rect -6097 3236 -6083 3250
rect 6167 3236 6181 3250
rect 7463 3236 7477 3250
rect -11617 3212 -11603 3226
rect -8521 3212 -8507 3226
rect 5231 3212 5245 3226
rect 5879 3212 5893 3226
rect 8543 3212 8557 3226
rect -11689 3188 -11675 3202
rect -3577 3188 -3563 3202
rect -3313 3188 -3299 3202
rect -3169 3188 -3155 3202
rect -3073 3188 -3059 3202
rect 10415 3188 10429 3202
rect -11833 3164 -11819 3178
rect 2807 3164 2821 3178
rect 2903 3164 2917 3178
rect 5519 3164 5533 3178
rect 6167 3164 6181 3178
rect 6239 3164 6253 3178
rect 6359 3164 6373 3178
rect 6527 3164 6541 3178
rect 6839 3164 6853 3178
rect 7199 3164 7213 3178
rect -11857 3140 -11843 3154
rect -8761 3140 -8747 3154
rect -8545 3140 -8531 3154
rect -1873 3140 -1859 3154
rect 671 3140 685 3154
rect 4055 3140 4069 3154
rect 7535 3140 7549 3154
rect 9167 3140 9181 3154
rect 11675 3140 11689 3154
rect -11905 3116 -11891 3130
rect -7489 3116 -7475 3130
rect -7417 3116 -7403 3130
rect 5351 3116 5365 3130
rect -11953 3092 -11939 3106
rect -11233 3092 -11219 3106
rect -10489 3092 -10475 3106
rect -10441 3092 -10427 3106
rect -6121 3092 -6107 3106
rect -4105 3092 -4091 3106
rect -1849 3092 -1835 3106
rect 2375 3092 2389 3106
rect 2495 3092 2509 3106
rect 2783 3092 2797 3106
rect 3263 3092 3277 3106
rect 4103 3092 4117 3106
rect 4367 3092 4381 3106
rect 5495 3092 5509 3106
rect 7559 3092 7573 3106
rect 9863 3092 9877 3106
rect 10991 3092 11005 3106
rect -11977 3068 -11963 3082
rect -8041 3068 -8027 3082
rect 5759 3068 5773 3082
rect -11977 3044 -11963 3058
rect 1655 3044 1669 3058
rect 2375 3044 2389 3058
rect 2447 3044 2461 3058
rect 2663 3044 2677 3058
rect 2687 3044 2701 3058
rect 2735 3044 2749 3058
rect 2951 3044 2965 3058
rect 4103 3044 4117 3058
rect 4223 3044 4237 3058
rect 4439 3044 4453 3058
rect 11927 3044 11941 3058
rect -12025 3020 -12011 3034
rect -8641 3020 -8627 3034
rect -4225 3020 -4211 3034
rect -361 3020 -347 3034
rect 4247 3020 4261 3034
rect 5231 3020 5245 3034
rect 5615 3020 5629 3034
rect -12025 2996 -12011 3010
rect -11809 2996 -11795 3010
rect -11737 2996 -11723 3010
rect -4273 2996 -4259 3010
rect -4129 2996 -4115 3010
rect 6095 2996 6109 3010
rect 9839 2996 9853 3010
rect -12049 2972 -12035 2986
rect -11377 2972 -11363 2986
rect -5929 2972 -5915 2986
rect 1271 2972 1285 2986
rect 3815 2972 3829 2986
rect 11735 2972 11749 2986
rect -12049 2948 -12035 2962
rect 7055 2948 7069 2962
rect -12073 2924 -12059 2938
rect -8353 2924 -8339 2938
rect -8281 2924 -8267 2938
rect -4657 2924 -4643 2938
rect -2977 2924 -2963 2938
rect -2809 2924 -2795 2938
rect 5471 2924 5485 2938
rect 9719 2924 9733 2938
rect 10655 2924 10669 2938
rect 11615 2924 11629 2938
rect 11927 2924 11941 2938
rect 12167 2924 12181 2938
rect -12113 2900 -12099 2914
rect -5833 2900 -5819 2914
rect 8783 2900 8797 2914
rect 11615 2900 11629 2914
rect 11675 2900 11689 2914
rect -12113 2876 -12099 2890
rect -3529 2876 -3515 2890
rect -3001 2876 -2987 2890
rect 2591 2876 2605 2890
rect 8591 2876 8605 2890
rect -12073 2852 -12059 2866
rect -7273 2852 -7259 2866
rect -5281 2852 -5267 2866
rect -5113 2852 -5099 2866
rect 2279 2852 2293 2866
rect 5951 2852 5965 2866
rect 7055 2852 7069 2866
rect 7223 2852 7237 2866
rect -11929 2828 -11915 2842
rect -11041 2828 -11027 2842
rect -2233 2828 -2219 2842
rect -2065 2828 -2051 2842
rect 4007 2828 4021 2842
rect 5015 2828 5029 2842
rect 5303 2828 5317 2842
rect 11039 2828 11053 2842
rect -11905 2804 -11891 2818
rect -11257 2804 -11243 2818
rect -10921 2804 -10907 2818
rect -9337 2804 -9323 2818
rect -8713 2804 -8699 2818
rect -8449 2804 -8435 2818
rect 4079 2804 4093 2818
rect 6071 2804 6085 2818
rect 6575 2804 6589 2818
rect 7919 2804 7933 2818
rect 11135 2804 11149 2818
rect 11639 2804 11653 2818
rect -11857 2780 -11843 2794
rect -11161 2780 -11147 2794
rect 5207 2780 5221 2794
rect 5471 2780 5485 2794
rect 5651 2780 5665 2794
rect -11785 2756 -11771 2770
rect -6049 2756 -6035 2770
rect -6001 2756 -5987 2770
rect 9023 2756 9037 2770
rect -11329 2732 -11315 2746
rect -9481 2732 -9467 2746
rect -8377 2732 -8363 2746
rect -4633 2732 -4619 2746
rect -4297 2732 -4283 2746
rect -1297 2732 -1283 2746
rect -529 2732 -515 2746
rect 95 2732 109 2746
rect 3119 2732 3133 2746
rect 5687 2732 5701 2746
rect 5927 2732 5941 2746
rect 7583 2732 7597 2746
rect 11759 2732 11773 2746
rect 12215 2732 12229 2746
rect -11161 2708 -11147 2722
rect -10297 2708 -10283 2722
rect -8809 2708 -8795 2722
rect -7345 2708 -7331 2722
rect 3359 2708 3373 2722
rect 4415 2708 4429 2722
rect 5639 2708 5653 2722
rect 6479 2708 6493 2722
rect 6551 2708 6565 2722
rect 9119 2708 9133 2722
rect 9743 2708 9757 2722
rect 11183 2708 11197 2722
rect 11759 2708 11773 2722
rect 12263 2708 12277 2722
rect -11089 2684 -11075 2698
rect 6047 2684 6061 2698
rect 10511 2684 10525 2698
rect -11065 2660 -11051 2674
rect -7369 2660 -7355 2674
rect 2639 2660 2653 2674
rect 3023 2660 3037 2674
rect 6047 2660 6061 2674
rect 6119 2660 6133 2674
rect 6551 2660 6565 2674
rect 6599 2660 6613 2674
rect 9023 2660 9037 2674
rect 9335 2660 9349 2674
rect -11017 2636 -11003 2650
rect 5183 2636 5197 2650
rect 11303 2636 11317 2650
rect -10969 2612 -10955 2626
rect -7993 2612 -7979 2626
rect 3527 2612 3541 2626
rect 5183 2612 5197 2626
rect 11447 2612 11461 2626
rect -10945 2588 -10931 2602
rect -10393 2588 -10379 2602
rect -3865 2588 -3851 2602
rect 5159 2588 5173 2602
rect 5927 2588 5941 2602
rect 9119 2588 9133 2602
rect 9431 2588 9445 2602
rect -10729 2564 -10715 2578
rect 2471 2564 2485 2578
rect 5999 2564 6013 2578
rect -10681 2540 -10667 2554
rect -289 2540 -275 2554
rect 10943 2540 10957 2554
rect -10609 2516 -10595 2530
rect -1945 2516 -1931 2530
rect 10823 2516 10837 2530
rect 11711 2516 11725 2530
rect 12167 2516 12181 2530
rect -10585 2492 -10571 2506
rect -8593 2492 -8579 2506
rect -5689 2492 -5675 2506
rect -2641 2492 -2627 2506
rect -217 2492 -203 2506
rect 527 2492 541 2506
rect 8351 2492 8365 2506
rect 10559 2492 10573 2506
rect -10513 2468 -10499 2482
rect -10009 2468 -9995 2482
rect 719 2468 733 2482
rect 5399 2468 5413 2482
rect 5735 2468 5749 2482
rect 8351 2468 8365 2482
rect 8927 2468 8941 2482
rect -10465 2444 -10451 2458
rect 1367 2444 1381 2458
rect 7007 2444 7021 2458
rect 8591 2444 8605 2458
rect -10393 2420 -10379 2434
rect -7441 2420 -7427 2434
rect -4081 2420 -4067 2434
rect -3193 2420 -3179 2434
rect -649 2420 -635 2434
rect 1343 2420 1357 2434
rect 2879 2420 2893 2434
rect 6023 2420 6037 2434
rect 7439 2420 7453 2434
rect 9719 2420 9733 2434
rect -10249 2396 -10235 2410
rect 4319 2396 4333 2410
rect 5399 2396 5413 2410
rect 5903 2396 5917 2410
rect -10225 2372 -10211 2386
rect 6623 2372 6637 2386
rect -10177 2348 -10163 2362
rect 2879 2348 2893 2362
rect -9745 2324 -9731 2338
rect -3865 2324 -3851 2338
rect -3217 2324 -3203 2338
rect -2713 2324 -2699 2338
rect 1319 2324 1333 2338
rect 2471 2324 2485 2338
rect 2567 2324 2581 2338
rect 2831 2324 2845 2338
rect 9791 2324 9805 2338
rect -9601 2300 -9587 2314
rect -6577 2300 -6563 2314
rect -457 2300 -443 2314
rect 3623 2300 3637 2314
rect 8879 2300 8893 2314
rect -9577 2276 -9563 2290
rect -1561 2276 -1547 2290
rect 3551 2276 3565 2290
rect -9529 2252 -9515 2266
rect 10007 2252 10021 2266
rect -9409 2228 -9395 2242
rect -8929 2228 -8915 2242
rect -8881 2228 -8867 2242
rect -841 2228 -827 2242
rect -529 2228 -515 2242
rect -397 2228 -383 2242
rect -361 2228 -347 2242
rect -265 2228 -251 2242
rect -217 2228 -203 2242
rect -25 2228 -11 2242
rect 23 2228 37 2242
rect 3143 2228 3157 2242
rect -9385 2204 -9371 2218
rect -7681 2204 -7667 2218
rect -3913 2204 -3899 2218
rect 2303 2204 2317 2218
rect 5855 2204 5869 2218
rect 7103 2204 7117 2218
rect -9361 2180 -9347 2194
rect -9169 2180 -9155 2194
rect -3817 2180 -3803 2194
rect -3769 2180 -3755 2194
rect -2593 2180 -2579 2194
rect -553 2180 -539 2194
rect 4151 2180 4165 2194
rect 5711 2180 5725 2194
rect 8279 2180 8293 2194
rect 8759 2180 8773 2194
rect -9337 2156 -9323 2170
rect -7825 2156 -7811 2170
rect 3551 2156 3565 2170
rect 5975 2156 5989 2170
rect -9265 2132 -9251 2146
rect -8785 2132 -8771 2146
rect -4201 2132 -4187 2146
rect -2137 2132 -2123 2146
rect 5375 2132 5389 2146
rect 5543 2132 5557 2146
rect 5831 2132 5845 2146
rect -8833 2108 -8819 2122
rect -5545 2108 -5531 2122
rect -4729 2108 -4715 2122
rect 2159 2108 2173 2122
rect -8449 2084 -8435 2098
rect -1657 2084 -1643 2098
rect -1417 2084 -1403 2098
rect 2543 2084 2557 2098
rect -8425 2060 -8411 2074
rect 3719 2060 3733 2074
rect -8401 2036 -8387 2050
rect -577 2036 -563 2050
rect 5279 2036 5293 2050
rect 11951 2036 11965 2050
rect -8377 2012 -8363 2026
rect -7321 2012 -7307 2026
rect -5593 2012 -5579 2026
rect -3289 2012 -3275 2026
rect -1753 2012 -1739 2026
rect 8207 2012 8221 2026
rect 10487 2012 10501 2026
rect 11207 2012 11221 2026
rect -8353 1988 -8339 2002
rect -1153 1988 -1139 2002
rect -913 1988 -899 2002
rect 11375 1988 11389 2002
rect -8113 1964 -8099 1978
rect -7681 1964 -7667 1978
rect -7633 1964 -7619 1978
rect -3841 1964 -3827 1978
rect -3625 1964 -3611 1978
rect -505 1964 -491 1978
rect 3863 1964 3877 1978
rect 7415 1964 7429 1978
rect 9215 1964 9229 1978
rect 9815 1964 9829 1978
rect -7873 1940 -7859 1954
rect 6887 1940 6901 1954
rect -7825 1916 -7811 1930
rect -6241 1916 -6227 1930
rect -433 1916 -419 1930
rect -337 1916 -323 1930
rect -193 1916 -179 1930
rect 167 1916 181 1930
rect 5327 1916 5341 1930
rect -7585 1892 -7571 1906
rect 5423 1892 5437 1906
rect -7537 1868 -7523 1882
rect 3095 1868 3109 1882
rect 5279 1868 5293 1882
rect 5783 1868 5797 1882
rect -7369 1844 -7355 1858
rect -4465 1844 -4451 1858
rect 215 1844 229 1858
rect 431 1844 445 1858
rect 7247 1844 7261 1858
rect 12287 1844 12301 1858
rect -7321 1820 -7307 1834
rect 1223 1820 1237 1834
rect -7201 1796 -7187 1810
rect 11111 1796 11125 1810
rect -7105 1772 -7091 1786
rect -2833 1772 -2819 1786
rect -2473 1772 -2459 1786
rect 8735 1772 8749 1786
rect 11555 1772 11569 1786
rect -7057 1748 -7043 1762
rect -7033 1748 -7019 1762
rect -6985 1748 -6971 1762
rect 6791 1748 6805 1762
rect 11783 1748 11797 1762
rect -7009 1724 -6995 1738
rect 10031 1724 10045 1738
rect 11783 1724 11797 1738
rect 12491 1724 12505 1738
rect -6961 1700 -6947 1714
rect 2639 1700 2653 1714
rect -6769 1676 -6755 1690
rect -6625 1676 -6611 1690
rect -6577 1676 -6563 1690
rect -5137 1676 -5123 1690
rect -2089 1676 -2075 1690
rect 8567 1676 8581 1690
rect 8999 1676 9013 1690
rect -6721 1652 -6707 1666
rect -6313 1652 -6299 1666
rect -5377 1652 -5363 1666
rect -3097 1652 -3083 1666
rect 1319 1652 1333 1666
rect 2759 1652 2773 1666
rect 4175 1652 4189 1666
rect 8999 1652 9013 1666
rect 9287 1652 9301 1666
rect -6697 1628 -6683 1642
rect -5257 1628 -5243 1642
rect -3985 1628 -3971 1642
rect 4583 1628 4597 1642
rect 11063 1628 11077 1642
rect -6505 1604 -6491 1618
rect -6265 1604 -6251 1618
rect -3457 1604 -3443 1618
rect -3049 1604 -3035 1618
rect -2449 1604 -2435 1618
rect 3791 1604 3805 1618
rect 4175 1604 4189 1618
rect 4475 1604 4489 1618
rect -6361 1580 -6347 1594
rect -6289 1580 -6275 1594
rect -6217 1580 -6203 1594
rect 407 1580 421 1594
rect 455 1580 469 1594
rect 11807 1580 11821 1594
rect -6313 1556 -6299 1570
rect -3025 1556 -3011 1570
rect -2401 1556 -2387 1570
rect 11975 1556 11989 1570
rect -6169 1532 -6155 1546
rect 71 1532 85 1546
rect 791 1532 805 1546
rect 6311 1532 6325 1546
rect 11975 1532 11989 1546
rect 12695 1532 12709 1546
rect -6097 1508 -6083 1522
rect 3935 1508 3949 1522
rect 4535 1508 4549 1522
rect 6311 1508 6325 1522
rect 8663 1508 8677 1522
rect -5929 1484 -5915 1498
rect -5893 1484 -5879 1498
rect -5857 1484 -5843 1498
rect 9263 1484 9277 1498
rect -5881 1460 -5867 1474
rect 4751 1460 4765 1474
rect -5785 1436 -5771 1450
rect -5761 1436 -5747 1450
rect -5713 1436 -5699 1450
rect -4873 1436 -4859 1450
rect 2231 1436 2245 1450
rect -5689 1412 -5675 1426
rect 7967 1412 7981 1426
rect -5377 1388 -5363 1402
rect -865 1388 -851 1402
rect 359 1388 373 1402
rect 5711 1388 5725 1402
rect 6263 1388 6277 1402
rect 10247 1388 10261 1402
rect -5353 1364 -5339 1378
rect 12719 1364 12733 1378
rect -5161 1340 -5147 1354
rect -1609 1340 -1595 1354
rect -1129 1340 -1115 1354
rect 8831 1340 8845 1354
rect -5113 1316 -5099 1330
rect -5065 1316 -5051 1330
rect -5017 1316 -5003 1330
rect -2353 1316 -2339 1330
rect -2281 1316 -2267 1330
rect -2041 1316 -2027 1330
rect -1729 1316 -1715 1330
rect 4367 1316 4381 1330
rect 6263 1316 6277 1330
rect 6419 1316 6433 1330
rect -4945 1292 -4931 1306
rect 6335 1292 6349 1306
rect 8687 1292 8701 1306
rect -4849 1268 -4835 1282
rect -2929 1268 -2915 1282
rect -169 1268 -155 1282
rect -121 1268 -107 1282
rect 5087 1268 5101 1282
rect 8807 1268 8821 1282
rect 10367 1268 10381 1282
rect 11207 1268 11221 1282
rect -4465 1244 -4451 1258
rect 6719 1244 6733 1258
rect -4417 1220 -4403 1234
rect 695 1220 709 1234
rect 839 1220 853 1234
rect 7631 1220 7645 1234
rect -4201 1196 -4187 1210
rect -4057 1196 -4043 1210
rect -3937 1196 -3923 1210
rect 4295 1196 4309 1210
rect -4081 1172 -4067 1186
rect 9695 1172 9709 1186
rect -3553 1148 -3539 1162
rect 11903 1148 11917 1162
rect -3193 1124 -3179 1138
rect -3121 1124 -3107 1138
rect -2329 1124 -2315 1138
rect 7511 1124 7525 1138
rect -2041 1100 -2027 1114
rect 3839 1100 3853 1114
rect -841 1076 -827 1090
rect -601 1076 -587 1090
rect -241 1076 -227 1090
rect -49 1076 -35 1090
rect 1031 1076 1045 1090
rect 1295 1076 1309 1090
rect 2231 1076 2245 1090
rect 2327 1076 2341 1090
rect 12767 1076 12781 1090
rect 12838 1076 12852 1090
rect -169 1052 -155 1066
rect 2399 1052 2413 1066
rect 6191 1052 6205 1066
rect 12743 1052 12757 1066
rect 12838 1052 12852 1066
rect -433 219 -419 233
rect 3047 219 3061 233
rect -817 195 -803 209
rect -25 195 -11 209
rect 815 195 829 209
rect 11567 195 11581 209
rect -1033 171 -1019 185
rect 2399 171 2413 185
rect 2855 171 2869 185
rect 7223 171 7237 185
rect -1081 147 -1067 161
rect 2183 147 2197 161
rect 3023 147 3037 161
rect 7871 147 7885 161
rect -3793 123 -3779 137
rect 3983 123 3997 137
rect -5905 99 -5891 113
rect -5881 99 -5867 113
rect -5641 99 -5627 113
rect -409 99 -395 113
rect 767 99 781 113
rect 3671 99 3685 113
rect -5905 75 -5891 89
rect 11543 75 11557 89
rect -6193 51 -6179 65
rect -961 51 -947 65
rect 2999 51 3013 65
rect -6337 27 -6323 41
rect 3143 27 3157 41
rect -6385 3 -6371 17
rect -4297 3 -4283 17
rect -4009 3 -3995 17
rect -3601 3 -3587 17
rect -1465 3 -1451 17
rect 503 3 517 17
rect 575 3 589 17
rect 1943 3 1957 17
rect 2783 3 2797 17
rect 8063 3 8077 17
rect -6553 -21 -6539 -7
rect -5185 -21 -5171 -7
rect -3361 -21 -3347 -7
rect -289 -21 -275 -7
rect 335 -21 349 -7
rect 3479 -21 3493 -7
rect -6673 -45 -6659 -31
rect -4345 -45 -4331 -31
rect -4033 -45 -4019 -31
rect 6407 -45 6421 -31
rect 6575 -45 6589 -31
rect 7991 -45 8005 -31
rect -6793 -69 -6779 -55
rect -3529 -69 -3515 -55
rect -2353 -69 -2339 -55
rect 551 -69 565 -55
rect 599 -69 613 -55
rect 911 -69 925 -55
rect 1007 -69 1021 -55
rect 2927 -69 2941 -55
rect 5327 -69 5341 -55
rect 10943 -69 10957 -55
rect -6961 -93 -6947 -79
rect -4561 -93 -4547 -79
rect -4369 -93 -4355 -79
rect -3721 -93 -3707 -79
rect -3481 -93 -3467 -79
rect -385 -93 -371 -79
rect -265 -93 -251 -79
rect 7727 -93 7741 -79
rect -7057 -117 -7043 -103
rect 3575 -117 3589 -103
rect 3767 -117 3781 -103
rect 10103 -117 10117 -103
rect -7153 -141 -7139 -127
rect 8543 -141 8557 -127
rect 8807 -141 8821 -127
rect 9959 -141 9973 -127
rect -7417 -165 -7403 -151
rect 2615 -165 2629 -151
rect 2759 -165 2773 -151
rect 10607 -165 10621 -151
rect -7537 -189 -7523 -175
rect 8855 -189 8869 -175
rect -7561 -213 -7547 -199
rect -2881 -213 -2867 -199
rect -2785 -213 -2771 -199
rect 5375 -213 5389 -199
rect 5423 -213 5437 -199
rect 10247 -213 10261 -199
rect -7609 -237 -7595 -223
rect -7225 -237 -7211 -223
rect -7177 -237 -7163 -223
rect 119 -237 133 -223
rect 311 -237 325 -223
rect 9143 -237 9157 -223
rect 9911 -237 9925 -223
rect 12407 -237 12421 -223
rect 12455 -237 12469 -223
rect -8713 -261 -8699 -247
rect 2327 -261 2341 -247
rect 2687 -261 2701 -247
rect 12838 -261 12852 -247
rect -8737 -285 -8723 -271
rect 3287 -285 3301 -271
rect 3383 -285 3397 -271
rect 9983 -285 9997 -271
rect 12359 -285 12373 -271
rect 12431 -285 12445 -271
rect -8785 -309 -8771 -295
rect -5881 -309 -5867 -295
rect 3815 -309 3829 -295
rect 7199 -309 7213 -295
rect 9071 -309 9085 -295
rect -9025 -333 -9011 -319
rect 8423 -333 8437 -319
rect -9049 -357 -9035 -343
rect 7415 -357 7429 -343
rect -9121 -381 -9107 -367
rect -6937 -381 -6923 -367
rect -6889 -381 -6875 -367
rect 12407 -381 12421 -367
rect -9145 -405 -9131 -391
rect 8639 -405 8653 -391
rect 8735 -405 8749 -391
rect 11231 -405 11245 -391
rect -9217 -429 -9203 -415
rect -4729 -429 -4715 -415
rect -4321 -429 -4307 -415
rect -2209 -429 -2195 -415
rect -1177 -429 -1163 -415
rect 11159 -429 11173 -415
rect -9241 -453 -9227 -439
rect 11687 -453 11701 -439
rect -9313 -477 -9299 -463
rect -4921 -477 -4907 -463
rect -4705 -477 -4691 -463
rect 3335 -477 3349 -463
rect -9505 -501 -9491 -487
rect -8689 -501 -8675 -487
rect -7681 -501 -7667 -487
rect 335 -501 349 -487
rect 1391 -501 1405 -487
rect 2135 -501 2149 -487
rect 8183 -501 8197 -487
rect -9553 -525 -9539 -511
rect -49 -525 -35 -511
rect 1535 -525 1549 -511
rect 4967 -525 4981 -511
rect -10153 -549 -10139 -535
rect 959 -549 973 -535
rect -10273 -573 -10259 -559
rect 287 -573 301 -559
rect -10321 -597 -10307 -583
rect -3145 -597 -3131 -583
rect 407 -597 421 -583
rect 9191 -597 9205 -583
rect -10369 -621 -10355 -607
rect -4489 -621 -4475 -607
rect -3985 -621 -3971 -607
rect 5759 -621 5773 -607
rect -10417 -645 -10403 -631
rect -2569 -645 -2555 -631
rect 6383 -645 6397 -631
rect 10799 -645 10813 -631
rect -10561 -669 -10547 -655
rect -4441 -669 -4427 -655
rect -3841 -669 -3827 -655
rect 887 -669 901 -655
rect -10705 -693 -10691 -679
rect 8903 -693 8917 -679
rect -11185 -717 -11171 -703
rect 7631 -717 7645 -703
rect -12113 -741 -12099 -727
rect -11977 -741 -11963 -727
rect -11737 -741 -11723 -727
rect -7129 -741 -7115 -727
rect -7081 -741 -7067 -727
rect -5065 -741 -5051 -727
rect 7511 -741 7525 -727
rect 12455 -741 12469 -727
rect 12838 -741 12852 -727
rect -12113 -765 -12099 -751
rect -10849 -765 -10835 -751
rect -10801 -765 -10787 -751
rect 4559 -765 4573 -751
rect 12431 -765 12445 -751
rect 12838 -765 12852 -751
rect -6625 -789 -6611 -775
rect -5869 -789 -5855 -775
rect -5425 -789 -5411 -775
rect 263 -789 277 -775
rect 12407 -789 12421 -775
rect 12838 -789 12852 -775
<< metal2 >>
rect -12183 7022 -12113 7034
rect -12183 6998 -12113 7010
rect -11364 6987 -11352 7165
rect -10812 7059 -10800 7165
rect -10404 7083 -10392 7165
rect -10403 7069 -10385 7083
rect -10811 7045 -10793 7059
rect -11376 6819 -11364 6973
rect -10824 6819 -10812 7045
rect -10440 6819 -10428 7045
rect -10416 6819 -10404 7069
rect -9600 7059 -9588 7165
rect -9264 6819 -9252 6973
rect -8592 6819 -8580 7045
rect -8448 6819 -8436 7069
rect -7980 6963 -7968 7165
rect -7152 6963 -7140 7165
rect -7116 7059 -7104 7165
rect -6288 7083 -6276 7165
rect -7344 6819 -7332 6949
rect -7056 6819 -7044 7045
rect -6552 6819 -6540 6925
rect -6360 6819 -6348 7021
rect -5064 6819 -5052 7021
rect -4800 6819 -4788 7069
rect -4668 6963 -4656 7165
rect -4728 6819 -4716 6949
rect -4608 6819 -4596 7093
rect -3840 6915 -3828 7165
rect -3252 7131 -3240 7165
rect -2364 7131 -2352 7165
rect -3251 7117 -3233 7131
rect -2363 7117 -2345 7131
rect -3264 6819 -3252 7117
rect -2376 6819 -2364 7117
rect -2148 7059 -2136 7165
rect -1656 6819 -1644 7045
rect -1512 6819 -1500 7117
rect -1320 7083 -1308 7165
rect -912 6819 -900 6973
rect -816 6819 -804 7069
rect -600 6819 -588 6877
rect -432 6819 -420 7141
rect 300 6867 312 7165
rect 456 6819 468 6925
rect 1116 6843 1128 7165
rect 1140 7083 1152 7165
rect 1956 7107 1968 7165
rect 3564 7083 3576 7165
rect 4308 7083 4320 7165
rect 4309 7069 4327 7083
rect 1944 6819 1956 6997
rect 3552 6819 3564 6997
rect 3696 6819 3708 7069
rect 4296 6819 4308 7069
rect 4404 7059 4416 7165
rect 6012 7059 6024 7165
rect 6828 7107 6840 7165
rect 7644 7107 7656 7165
rect 5592 6819 5604 6973
rect 6288 6819 6300 7069
rect 6864 6819 6876 6925
rect 6960 6819 6972 7093
rect 7668 7035 7680 7165
rect 7200 6819 7212 6901
rect 8016 6819 8028 6901
rect 8160 6819 8172 7093
rect 8484 6915 8496 7165
rect 9300 7131 9312 7165
rect 10116 7155 10128 7165
rect 8736 6819 8748 6829
rect 8928 6819 8940 6901
rect 9432 6819 9444 7045
rect 10932 6939 10944 7165
rect 11748 6915 11760 7165
rect 10272 6819 10284 6829
rect 11328 6819 11340 6853
rect 11880 6819 11892 6949
rect 12048 6819 12060 6973
rect 12720 6819 12732 6973
rect 12744 6939 12756 6997
rect 12768 6891 12780 6973
rect 12744 6867 12756 6877
rect 12792 6843 12804 6901
rect 12816 6843 12828 7069
rect 12852 6926 12922 6938
rect 12852 6902 12922 6914
rect 12852 6878 12922 6890
rect 12852 6854 12922 6866
rect 12852 6830 12922 6842
rect -12072 2938 -12060 6020
rect -12048 2986 -12036 6020
rect -12024 3034 -12012 6020
rect -11976 3082 -11964 6020
rect -11952 3106 -11940 6020
rect -11904 3130 -11892 6020
rect -11856 3154 -11844 6020
rect -11832 3178 -11820 6020
rect -12183 2901 -12113 2913
rect -12183 2877 -12113 2889
rect -12072 1042 -12060 2852
rect -12048 1042 -12036 2948
rect -12024 1042 -12012 2996
rect -11976 1042 -11964 3044
rect -11808 3010 -11796 6020
rect -11928 1042 -11916 2828
rect -11904 1042 -11892 2804
rect -11856 1042 -11844 2780
rect -11784 2770 -11772 6020
rect -11736 3010 -11724 6020
rect -11688 3202 -11676 6020
rect -11616 3226 -11604 6020
rect -11568 3250 -11556 6020
rect -11496 3274 -11484 6020
rect -11472 3298 -11460 6020
rect -11424 3322 -11412 6020
rect -11328 3346 -11316 6020
rect -11376 1042 -11364 2972
rect -11256 2818 -11244 6020
rect -11232 3106 -11220 6020
rect -11208 3370 -11196 6020
rect -11160 2794 -11148 6020
rect -11136 3418 -11124 6020
rect -11112 3442 -11100 6020
rect -11064 3466 -11052 6020
rect -11328 1042 -11316 2732
rect -11160 1042 -11148 2708
rect -11136 1042 -11124 3380
rect -11040 2842 -11028 6020
rect -11016 3490 -11004 6020
rect -10968 3514 -10956 6020
rect -10944 3538 -10932 6020
rect -10920 2818 -10908 6020
rect -10896 3586 -10884 6020
rect -11088 1042 -11076 2684
rect -11064 1042 -11052 2660
rect -11016 1042 -11004 2636
rect -10968 1042 -10956 2612
rect -10944 1042 -10932 2588
rect -10896 1042 -10884 3548
rect -10848 3346 -10836 6020
rect -10824 3610 -10812 6020
rect -10800 3634 -10788 6020
rect -10752 3658 -10740 6020
rect -10728 3370 -10716 6020
rect -10704 3682 -10692 6020
rect -10656 3730 -10644 6020
rect -10632 3754 -10620 6020
rect -10608 3778 -10596 6020
rect -10584 3802 -10572 6020
rect -10536 3826 -10524 6020
rect -10512 3850 -10500 6020
rect -10488 3874 -10476 6020
rect -10728 1042 -10716 2564
rect -10680 1042 -10668 2540
rect -10656 1042 -10644 3692
rect -10440 3106 -10428 6020
rect -10416 3898 -10404 6020
rect -10608 1042 -10596 2516
rect -10584 1042 -10572 2492
rect -10512 1042 -10500 2468
rect -10488 1042 -10476 3092
rect -10392 2602 -10380 6020
rect -10344 3922 -10332 6020
rect -10320 3946 -10308 6020
rect -10296 3970 -10284 6020
rect -10464 1042 -10452 2444
rect -10392 1042 -10380 2420
rect -10296 1042 -10284 2708
rect -10248 2410 -10236 6020
rect -10224 2386 -10212 6020
rect -10176 2362 -10164 6020
rect -10128 3994 -10116 6020
rect -10104 4018 -10092 6020
rect -10080 4042 -10068 6020
rect -10032 4066 -10020 6020
rect -10008 2482 -9996 6020
rect -9984 4090 -9972 6020
rect -9936 4114 -9924 6020
rect -9888 3538 -9876 6020
rect -9816 4090 -9804 6020
rect -9792 1042 -9780 4052
rect -9768 3466 -9756 6020
rect -9696 4138 -9684 6020
rect -9672 4162 -9660 6020
rect -9624 4186 -9612 6020
rect -9576 3538 -9564 6020
rect -9552 4210 -9540 6020
rect -9744 1042 -9732 2324
rect -9600 1042 -9588 2300
rect -9576 1042 -9564 2276
rect -9528 2266 -9516 6020
rect -9480 4234 -9468 6020
rect -9456 4258 -9444 6020
rect -9480 1042 -9468 2732
rect -9432 1042 -9420 4268
rect -9408 2242 -9396 6020
rect -9336 2818 -9324 6020
rect -9312 4306 -9300 6020
rect -9240 4330 -9228 6020
rect -9168 4354 -9156 6020
rect -9144 4378 -9132 6020
rect -9096 4402 -9084 6020
rect -9384 1042 -9372 2204
rect -9360 1042 -9348 2180
rect -9336 1042 -9324 2156
rect -9264 1042 -9252 2132
rect -9168 1042 -9156 2180
rect -9072 1042 -9060 4412
rect -9048 3298 -9036 6020
rect -9000 4450 -8988 6020
rect -8928 4522 -8916 6020
rect -8880 4570 -8868 6020
rect -8808 4594 -8796 6020
rect -8784 4618 -8772 6020
rect -8976 1042 -8964 4460
rect -8952 1042 -8940 4484
rect -8928 1042 -8916 2228
rect -8904 1042 -8892 4532
rect -8880 1042 -8868 2228
rect -8832 1042 -8820 2108
rect -8808 1042 -8796 2708
rect -8784 2146 -8772 4580
rect -8760 3154 -8748 6020
rect -8712 2818 -8700 6020
rect -8664 4594 -8652 6020
rect -8592 4306 -8580 6020
rect -8544 3154 -8532 6020
rect -8640 1042 -8628 3020
rect -8592 1042 -8580 2492
rect -8520 1042 -8508 3212
rect -8496 1042 -8484 3932
rect -8472 3346 -8460 6020
rect -8448 2818 -8436 6020
rect -8448 1042 -8436 2084
rect -8424 2074 -8412 6020
rect -8376 2746 -8364 6020
rect -8352 2938 -8340 6020
rect -8328 4642 -8316 6020
rect -8280 2938 -8268 6020
rect -8256 4666 -8244 6020
rect -8232 4714 -8220 6020
rect -8208 4738 -8196 6020
rect -8400 1042 -8388 2036
rect -8376 1042 -8364 2012
rect -8352 1042 -8340 1988
rect -8232 1042 -8220 4676
rect -8184 4498 -8172 6020
rect -8136 4498 -8124 6020
rect -8112 1978 -8100 6020
rect -8088 4762 -8076 6020
rect -8040 3082 -8028 6020
rect -7992 2626 -7980 6020
rect -7920 4786 -7908 6020
rect -7896 4810 -7884 6020
rect -7872 4210 -7860 6020
rect -7824 2170 -7812 6020
rect -7800 3850 -7788 6020
rect -7776 4210 -7764 6020
rect -7752 4834 -7740 6020
rect -7704 4666 -7692 6020
rect -7680 2218 -7668 6020
rect -7632 4858 -7620 6020
rect -7584 3778 -7572 6020
rect -7872 1042 -7860 1940
rect -7824 1042 -7812 1916
rect -7680 1042 -7668 1964
rect -7632 1042 -7620 1964
rect -7584 1042 -7572 1892
rect -7536 1882 -7524 6020
rect -7464 4906 -7452 6020
rect -7488 1042 -7476 3116
rect -7464 1042 -7452 4868
rect -7440 2434 -7428 6020
rect -7416 3130 -7404 6020
rect -7368 2674 -7356 6020
rect -7344 4930 -7332 6020
rect -7368 1042 -7356 1844
rect -7344 1042 -7332 2708
rect -7320 2026 -7308 4916
rect -7296 3514 -7284 6020
rect -7248 4930 -7236 6020
rect -7224 4954 -7212 6020
rect -7320 1042 -7308 1820
rect -7272 1042 -7260 2852
rect -7248 1042 -7236 4124
rect -7200 1810 -7188 6020
rect -7152 4978 -7140 6020
rect -7128 5002 -7116 6020
rect -7104 1786 -7092 6020
rect -7056 1762 -7044 6020
rect -7032 1042 -7020 1748
rect -7008 1738 -6996 6020
rect -6984 1042 -6972 1748
rect -6960 1714 -6948 6020
rect -6912 1042 -6900 5012
rect -6888 4714 -6876 6020
rect -6864 4066 -6852 6020
rect -6840 5050 -6828 6020
rect -6840 1042 -6828 3620
rect -6816 1042 -6804 4724
rect -6792 4498 -6780 6020
rect -6768 1690 -6756 6020
rect -6744 5074 -6732 6020
rect -6696 5098 -6684 6020
rect -6672 5122 -6660 6020
rect -6648 5146 -6636 6020
rect -6624 5170 -6612 6020
rect -6744 1042 -6732 4052
rect -6576 2314 -6564 6020
rect -6528 5218 -6516 6020
rect -6480 5266 -6468 6020
rect -6720 1042 -6708 1652
rect -6696 1042 -6684 1628
rect -6624 1042 -6612 1676
rect -6576 1042 -6564 1676
rect -6528 1042 -6516 5180
rect -6504 1042 -6492 1604
rect -6480 1042 -6468 5228
rect -6456 3850 -6444 6020
rect -6432 4330 -6420 6020
rect -6408 5290 -6396 6020
rect -6432 1042 -6420 4004
rect -6408 1042 -6396 4436
rect -6360 1594 -6348 6020
rect -6312 1666 -6300 6020
rect -6288 4450 -6276 6020
rect -6264 1618 -6252 6020
rect -6216 5314 -6204 6020
rect -6192 5338 -6180 6020
rect -6312 1042 -6300 1556
rect -6288 1042 -6276 1580
rect -6240 1042 -6228 1916
rect -6216 1042 -6204 1580
rect -6168 1546 -6156 6020
rect -6120 5362 -6108 6020
rect -6144 1042 -6132 3404
rect -6096 3250 -6084 6020
rect -6072 5386 -6060 6020
rect -6024 4066 -6012 6020
rect -6000 5410 -5988 6020
rect -5976 5338 -5964 6020
rect -6120 1042 -6108 3092
rect -5928 2986 -5916 6020
rect -5904 5338 -5892 6020
rect -6096 1042 -6084 1508
rect -6048 1042 -6036 2756
rect -6000 1042 -5988 2756
rect -5892 1498 -5880 5252
rect -5856 1498 -5844 6020
rect -5808 3490 -5796 6020
rect -5784 5266 -5772 6020
rect -5760 5434 -5748 6020
rect -5712 5410 -5700 6020
rect -5928 1042 -5916 1484
rect -5880 1042 -5868 1460
rect -5832 1042 -5820 2900
rect -5760 1450 -5748 5396
rect -5688 2506 -5676 6020
rect -5664 5458 -5652 6020
rect -5616 5482 -5604 6020
rect -5592 5506 -5580 6020
rect -5568 4762 -5556 6020
rect -5544 4690 -5532 6020
rect -5496 4690 -5484 6020
rect -5472 5266 -5460 6020
rect -5448 5530 -5436 6020
rect -5784 1042 -5772 1436
rect -5712 1042 -5700 1436
rect -5688 1042 -5676 1412
rect -5664 1042 -5652 3884
rect -5592 1042 -5580 2012
rect -5544 1042 -5532 2108
rect -5472 1042 -5460 3644
rect -5448 1042 -5436 4748
rect -5400 4666 -5388 6020
rect -5376 1666 -5364 6020
rect -5352 4618 -5340 6020
rect -5328 5554 -5316 6020
rect -5280 5506 -5268 6020
rect -5376 1042 -5364 1388
rect -5352 1042 -5340 1364
rect -5328 1042 -5316 5492
rect -5256 3442 -5244 6020
rect -5232 5602 -5220 6020
rect -5280 1042 -5268 2852
rect -5256 1042 -5244 1628
rect -5232 1042 -5220 5564
rect -5184 3442 -5172 6020
rect -5160 4666 -5148 6020
rect -5112 2866 -5100 6020
rect -5160 1042 -5148 1340
rect -5136 1042 -5124 1676
rect -5064 1330 -5052 6020
rect -5016 5266 -5004 6020
rect -4992 5626 -4980 6020
rect -4968 5650 -4956 6020
rect -4920 3634 -4908 6020
rect -5112 1042 -5100 1316
rect -5016 1042 -5004 1316
rect -4944 1042 -4932 1292
rect -4896 1042 -4884 5660
rect -4872 1450 -4860 6020
rect -4800 5674 -4788 6020
rect -4752 5674 -4740 6020
rect -4728 5698 -4716 6020
rect -4848 1042 -4836 1268
rect -4824 1042 -4812 4700
rect -4800 1042 -4788 3716
rect -4752 1042 -4740 3668
rect -4728 2122 -4716 5660
rect -4704 4810 -4692 6020
rect -4656 5674 -4644 6020
rect -4632 5722 -4620 6020
rect -4656 1042 -4644 2924
rect -4632 1042 -4620 2732
rect -4608 1042 -4596 4700
rect -4584 1042 -4572 4052
rect -4560 3538 -4548 6020
rect -4536 4618 -4524 6020
rect -4512 5746 -4500 6020
rect -4512 1042 -4500 4964
rect -4464 1858 -4452 6020
rect -4416 5770 -4404 6020
rect -4344 3466 -4332 6020
rect -4320 4906 -4308 6020
rect -4296 2746 -4284 6020
rect -4272 5026 -4260 6020
rect -4224 3418 -4212 6020
rect -4464 1042 -4452 1244
rect -4416 1042 -4404 1220
rect -4272 1042 -4260 2996
rect -4224 1042 -4212 3020
rect -4200 2146 -4188 6020
rect -4176 4210 -4164 6020
rect -4152 5026 -4140 6020
rect -4104 4018 -4092 6020
rect -4200 1042 -4188 1196
rect -4176 1042 -4164 3452
rect -4128 1042 -4116 2996
rect -4104 1042 -4092 3092
rect -4080 2434 -4068 6020
rect -4056 5794 -4044 6020
rect -4056 1210 -4044 5252
rect -4008 4066 -3996 6020
rect -3984 1642 -3972 6020
rect -3960 5818 -3948 6020
rect -4080 1042 -4068 1172
rect -3960 1042 -3948 4388
rect -3912 2218 -3900 6020
rect -3888 5842 -3876 6020
rect -3936 1042 -3924 1196
rect -3888 1042 -3876 3260
rect -3864 2602 -3852 6020
rect -3864 1042 -3852 2324
rect -3840 1978 -3828 6020
rect -3816 2194 -3804 5828
rect -3792 4834 -3780 6020
rect -3768 3418 -3756 6020
rect -3744 4834 -3732 6020
rect -3696 5842 -3684 6020
rect -3672 5698 -3660 6020
rect -3648 4426 -3636 6020
rect -3600 4402 -3588 6020
rect -3768 1042 -3756 2180
rect -3744 1042 -3732 4148
rect -3672 1042 -3660 3932
rect -3648 1042 -3636 3908
rect -3576 3202 -3564 6020
rect -3552 4402 -3540 6020
rect -3528 2890 -3516 6020
rect -3480 4426 -3468 6020
rect -3624 1042 -3612 1964
rect -3456 1618 -3444 6020
rect -3432 5866 -3420 6020
rect -3552 1042 -3540 1148
rect -3432 1042 -3420 5012
rect -3408 1042 -3396 5732
rect -3384 4114 -3372 6020
rect -3360 3370 -3348 6020
rect -3312 3922 -3300 6020
rect -3264 5026 -3252 6020
rect -3312 1042 -3300 3188
rect -3288 1042 -3276 2012
rect -3240 1042 -3228 4220
rect -3216 2338 -3204 6020
rect -3192 2434 -3180 6020
rect -3144 4666 -3132 6020
rect -3168 3202 -3156 3956
rect -3120 1138 -3108 5708
rect -3096 1666 -3084 6020
rect -3072 3970 -3060 6020
rect -3048 4234 -3036 6020
rect -3000 5746 -2988 6020
rect -3192 1042 -3180 1124
rect -3072 1042 -3060 3188
rect -3048 1042 -3036 1604
rect -3024 1570 -3012 4220
rect -2976 2938 -2964 6020
rect -3000 1042 -2988 2876
rect -2952 1042 -2940 4124
rect -2928 3442 -2916 6020
rect -2928 1042 -2916 1268
rect -2904 1042 -2892 4196
rect -2880 3538 -2868 6020
rect -2856 4186 -2844 6020
rect -2832 3754 -2820 6020
rect -2784 4906 -2772 6020
rect -2760 4666 -2748 6020
rect -2832 1042 -2820 1772
rect -2808 1042 -2796 2924
rect -2736 1042 -2724 5252
rect -2712 4234 -2700 6020
rect -2712 1042 -2700 2324
rect -2688 1042 -2676 5396
rect -2664 5266 -2652 6020
rect -2640 4570 -2628 6020
rect -2616 5146 -2604 6020
rect -2544 5266 -2532 6020
rect -2640 1042 -2628 2492
rect -2616 1042 -2604 3836
rect -2592 2194 -2580 4220
rect -2520 3442 -2508 6020
rect -2472 4234 -2460 6020
rect -2520 1042 -2508 3308
rect -2472 1042 -2460 1772
rect -2448 1618 -2436 6020
rect -2376 5890 -2364 6020
rect -2400 1042 -2388 1556
rect -2376 1042 -2364 5132
rect -2352 1330 -2340 5876
rect -2328 1138 -2316 6020
rect -2304 1042 -2292 4604
rect -2280 3418 -2268 6020
rect -2208 5890 -2196 6020
rect -2184 4738 -2172 6020
rect -2136 3946 -2124 6020
rect -2088 5914 -2076 6020
rect -2280 1042 -2268 1316
rect -2256 1042 -2244 3428
rect -2232 1042 -2220 2828
rect -2160 1042 -2148 3404
rect -2136 1042 -2124 2132
rect -2112 1042 -2100 4148
rect -2064 2842 -2052 6020
rect -2040 5938 -2028 6020
rect -1992 5962 -1980 6020
rect -2088 1042 -2076 1676
rect -2040 1330 -2028 4052
rect -2040 1042 -2028 1100
rect -1992 1042 -1980 5852
rect -1944 2530 -1932 6020
rect -1872 3154 -1860 6020
rect -1848 3106 -1836 6020
rect -1824 5866 -1812 6020
rect -1776 3370 -1764 6020
rect -1752 2026 -1740 6020
rect -1728 1330 -1716 6020
rect -1680 5986 -1668 6020
rect -1656 2098 -1644 6020
rect -1608 1354 -1596 6020
rect -1560 2290 -1548 6020
rect -1440 4282 -1428 6020
rect -1416 2098 -1404 6020
rect -1368 5194 -1356 6020
rect -1320 4282 -1308 6020
rect -1296 5194 -1284 6020
rect -1272 5530 -1260 6020
rect -1248 5002 -1236 6020
rect -1224 5530 -1212 6020
rect -1320 1042 -1308 3836
rect -1296 1042 -1284 2732
rect -1248 1042 -1236 4004
rect -1200 1042 -1188 4820
rect -1176 3898 -1164 6020
rect -1128 4738 -1116 6020
rect -1152 2002 -1140 4268
rect -1056 3490 -1044 6020
rect -1032 5962 -1020 6020
rect -1008 3994 -996 6020
rect -960 3610 -948 6020
rect -936 3994 -924 6020
rect -888 4282 -876 6020
rect -1128 1042 -1116 1340
rect -936 1042 -924 3476
rect -840 2242 -828 6020
rect -816 3322 -804 6020
rect -768 5674 -756 6020
rect -720 3682 -708 6020
rect -672 4258 -660 6020
rect -912 1042 -900 1988
rect -864 1042 -852 1388
rect -840 1042 -828 1076
rect -768 1042 -756 3356
rect -720 1042 -708 3356
rect -648 1042 -636 2420
rect -624 1042 -612 4580
rect -600 1090 -588 6020
rect -552 2194 -540 6020
rect -528 2746 -516 6020
rect -504 4546 -492 6020
rect -576 1042 -564 2036
rect -528 1042 -516 2228
rect -504 1042 -492 1964
rect -480 1042 -468 3308
rect -456 2314 -444 6020
rect -432 1930 -420 6020
rect -408 5482 -396 6020
rect -396 2242 -384 4580
rect -360 3034 -348 6020
rect -336 4450 -324 6020
rect -312 3850 -300 6020
rect -288 2554 -276 6020
rect -240 4666 -228 6020
rect -264 2242 -252 4268
rect -216 2506 -204 6020
rect -360 1042 -348 2228
rect -336 1042 -324 1916
rect -240 1042 -228 1076
rect -216 1042 -204 2228
rect -192 1930 -180 5348
rect -168 1282 -156 6020
rect -168 1042 -156 1052
rect -144 1042 -132 4124
rect -120 1282 -108 6020
rect -96 5746 -84 6020
rect -96 1042 -84 4220
rect -72 4114 -60 6020
rect -48 1090 -36 5540
rect -24 2242 -12 5012
rect 0 1042 12 5060
rect 48 3682 60 6020
rect 24 1042 36 2228
rect 72 1042 84 1532
rect 96 1042 108 2732
rect 168 1042 180 1916
rect 192 1042 204 5132
rect 216 1042 228 1844
rect 408 1594 420 6020
rect 360 1042 372 1388
rect 432 1042 444 1844
rect 456 1042 468 1580
rect 528 1042 540 2492
rect 648 1042 660 4604
rect 672 4114 684 6020
rect 672 1042 684 3140
rect 696 1234 708 4100
rect 720 1042 732 2468
rect 792 1042 804 1532
rect 840 1042 852 1220
rect 936 1042 948 5396
rect 1032 3850 1044 6020
rect 1080 5746 1092 6020
rect 1032 1042 1044 1076
rect 1080 1042 1092 5180
rect 1128 1042 1140 4124
rect 1152 1042 1164 3524
rect 1176 1042 1188 3932
rect 1200 1042 1212 4412
rect 1224 1834 1236 6020
rect 1248 3946 1260 6020
rect 1272 4114 1284 6020
rect 1248 1042 1260 3428
rect 1272 1042 1284 2972
rect 1296 1090 1308 4100
rect 1320 2338 1332 6020
rect 1344 2434 1356 6020
rect 1368 3298 1380 6020
rect 1416 4114 1428 6020
rect 1440 5290 1452 6020
rect 1464 4234 1476 6020
rect 1488 5650 1500 6020
rect 1512 4258 1524 6020
rect 1560 5050 1572 6020
rect 1584 4282 1596 6020
rect 1608 3874 1620 6020
rect 1632 5794 1644 6020
rect 1320 1042 1332 1652
rect 1368 1042 1380 2444
rect 1416 1042 1428 3284
rect 1656 3058 1668 6020
rect 1704 3874 1716 6020
rect 1728 3586 1740 6020
rect 1752 4426 1764 6020
rect 1776 3586 1788 6020
rect 1800 4546 1812 6020
rect 1848 5314 1860 6020
rect 1872 5770 1884 6020
rect 1896 4834 1908 6020
rect 1920 5026 1932 6020
rect 1992 3466 2004 6020
rect 2016 5050 2028 6020
rect 2040 5074 2052 6020
rect 2064 5410 2076 6020
rect 2088 5146 2100 6020
rect 2088 1042 2100 4124
rect 2112 1042 2124 4196
rect 2136 4162 2148 6020
rect 2160 2122 2172 6020
rect 2184 5194 2196 6020
rect 2208 1042 2220 4724
rect 2232 1450 2244 6020
rect 2256 4738 2268 6020
rect 2304 5290 2316 6020
rect 2232 1042 2244 1076
rect 2280 1042 2292 2852
rect 2304 1042 2316 2204
rect 2328 1090 2340 5900
rect 2352 5698 2364 6020
rect 2376 3106 2388 6020
rect 2424 5914 2436 6020
rect 2376 1042 2388 3044
rect 2400 1066 2412 5276
rect 2424 1042 2436 5876
rect 2448 3058 2460 3620
rect 2472 2578 2484 6020
rect 2496 3106 2508 6020
rect 2472 1042 2484 2324
rect 2520 1042 2532 3452
rect 2544 2098 2556 6020
rect 2568 2338 2580 3716
rect 2592 3634 2604 6020
rect 2616 3730 2628 6020
rect 2592 1042 2604 2876
rect 2640 2674 2652 6020
rect 2664 4690 2676 6020
rect 2688 3058 2700 5708
rect 2712 4618 2724 6020
rect 2736 4666 2748 6020
rect 2640 1042 2652 1700
rect 2664 1042 2676 3044
rect 2736 1042 2748 3044
rect 2760 1666 2772 6020
rect 2784 3106 2796 6020
rect 2808 3178 2820 6020
rect 2856 3850 2868 6020
rect 2880 2434 2892 6020
rect 2928 4666 2940 6020
rect 2832 1042 2844 2324
rect 2880 1042 2892 2348
rect 2904 1042 2916 3164
rect 2952 3058 2964 5252
rect 2976 4306 2988 6020
rect 3000 5698 3012 6020
rect 2976 1042 2988 3476
rect 3024 2674 3036 6020
rect 3096 1042 3108 1868
rect 3120 1042 3132 2732
rect 3144 2242 3156 6020
rect 3192 1042 3204 4724
rect 3216 1042 3228 3836
rect 3240 1042 3252 4844
rect 3264 1042 3276 3092
rect 3360 1042 3372 2708
rect 3432 1042 3444 3524
rect 3456 1042 3468 3500
rect 3528 1042 3540 2612
rect 3552 2290 3564 6020
rect 3552 1042 3564 2156
rect 3624 1042 3636 2300
rect 3648 1042 3660 3980
rect 3696 3562 3708 6020
rect 3744 4690 3756 6020
rect 3768 5098 3780 6020
rect 3720 1042 3732 2060
rect 3744 1042 3756 4292
rect 3792 1618 3804 6020
rect 3816 2986 3828 6020
rect 3840 1114 3852 6020
rect 3888 4666 3900 6020
rect 3912 3562 3924 6020
rect 3936 5050 3948 6020
rect 3984 5050 3996 6020
rect 4008 2842 4020 6020
rect 4032 4786 4044 6020
rect 4080 4786 4092 6020
rect 3864 1042 3876 1964
rect 3936 1042 3948 1508
rect 4056 1042 4068 3140
rect 4104 3106 4116 6020
rect 4128 5290 4140 6020
rect 4080 1042 4092 2804
rect 4104 1042 4116 3044
rect 4152 1042 4164 2180
rect 4176 1666 4188 6020
rect 4200 5266 4212 6020
rect 4248 5362 4260 6020
rect 4176 1042 4188 1604
rect 4200 1042 4212 3500
rect 4224 3058 4236 4508
rect 4248 1042 4260 3020
rect 4272 1042 4284 5732
rect 4296 1210 4308 6020
rect 4344 5698 4356 6020
rect 4368 3106 4380 6020
rect 4320 1042 4332 2396
rect 4368 1042 4380 1316
rect 4392 1042 4404 5732
rect 4464 5482 4476 6020
rect 4416 1042 4428 2708
rect 4440 1042 4452 3044
rect 4476 1618 4488 3284
rect 4536 1522 4548 6020
rect 4560 3322 4572 6020
rect 4584 1642 4596 6020
rect 4632 3442 4644 6020
rect 4656 4450 4668 6020
rect 4680 3778 4692 6020
rect 4728 5554 4740 6020
rect 4752 1474 4764 6020
rect 4800 4834 4812 6020
rect 4848 4834 4860 6020
rect 4896 4138 4908 6020
rect 4968 5050 4980 6020
rect 4992 3658 5004 6020
rect 5016 2842 5028 6020
rect 5040 3874 5052 6020
rect 5088 1282 5100 6020
rect 5112 3874 5124 6020
rect 5136 5650 5148 6020
rect 5112 1042 5124 3836
rect 5136 1042 5148 4844
rect 5184 2650 5196 6020
rect 5208 2794 5220 6020
rect 5232 3226 5244 6020
rect 5160 1042 5172 2588
rect 5184 1042 5196 2612
rect 5232 1042 5244 3020
rect 5256 1042 5268 5804
rect 5280 2050 5292 6020
rect 5304 2842 5316 6020
rect 5328 1930 5340 6020
rect 5280 1042 5292 1868
rect 5352 1042 5364 3116
rect 5376 2146 5388 6020
rect 5400 2482 5412 6020
rect 5400 1042 5412 2396
rect 5424 1906 5436 6020
rect 5448 3298 5460 3860
rect 5472 2938 5484 6020
rect 5496 3874 5508 6020
rect 5520 3178 5532 6020
rect 5568 3610 5580 6020
rect 5472 1042 5484 2780
rect 5496 1042 5508 3092
rect 5544 1042 5556 2132
rect 5592 1042 5604 5684
rect 5616 3034 5628 5948
rect 5640 4210 5652 6020
rect 5652 2794 5664 3524
rect 5688 2746 5700 6020
rect 5640 1042 5652 2708
rect 5712 2194 5724 6020
rect 5736 2482 5748 6020
rect 5760 3082 5772 6020
rect 5808 4138 5820 6020
rect 5784 1882 5796 3956
rect 5832 3898 5844 6020
rect 5880 4162 5892 6020
rect 5712 1042 5724 1388
rect 5832 1042 5844 2132
rect 5856 1042 5868 2204
rect 5880 1042 5892 3212
rect 5904 2410 5916 4628
rect 5928 2746 5940 6020
rect 5952 2866 5964 6020
rect 5976 4618 5988 6020
rect 5928 1042 5940 2588
rect 6000 2578 6012 6020
rect 6024 2434 6036 3860
rect 6048 2698 6060 6020
rect 6096 3658 6108 6020
rect 5976 1042 5988 2156
rect 6048 1042 6060 2660
rect 6072 1042 6084 2804
rect 6096 1042 6108 2996
rect 6120 2674 6132 4772
rect 6144 1042 6156 4292
rect 6168 3250 6180 6020
rect 6168 1042 6180 3164
rect 6192 1066 6204 6020
rect 6216 5674 6228 6020
rect 6216 1042 6228 5324
rect 6240 3178 6252 3884
rect 6264 1402 6276 6020
rect 6264 1042 6276 1316
rect 6288 1042 6300 4724
rect 6312 1546 6324 6020
rect 6312 1042 6324 1508
rect 6336 1306 6348 5660
rect 6360 3394 6372 6020
rect 6384 4594 6396 6020
rect 6408 3730 6420 6020
rect 6456 5962 6468 6020
rect 6360 1042 6372 3164
rect 6420 1330 6432 3452
rect 6456 1042 6468 5180
rect 6480 4090 6492 6020
rect 6504 3826 6516 6020
rect 6480 1042 6492 2708
rect 6504 1042 6516 3380
rect 6528 3178 6540 5420
rect 6552 2722 6564 6020
rect 6576 2818 6588 6020
rect 6624 5050 6636 6020
rect 6672 5458 6684 6020
rect 6696 5746 6708 6020
rect 6600 2674 6612 4628
rect 6552 1042 6564 2660
rect 6624 1042 6636 2372
rect 6672 1042 6684 5396
rect 6696 1042 6708 3836
rect 6720 1258 6732 6020
rect 6744 1042 6756 5300
rect 6768 3538 6780 6020
rect 6792 5698 6804 6020
rect 6816 4474 6828 6020
rect 6792 1042 6804 1748
rect 6840 1042 6852 3164
rect 6888 1954 6900 6020
rect 6912 4474 6924 6020
rect 6912 1042 6924 4148
rect 6936 1042 6948 4196
rect 6960 3706 6972 6020
rect 6984 1042 6996 4772
rect 7008 2458 7020 6020
rect 7032 4834 7044 6020
rect 7032 1042 7044 3404
rect 7056 2962 7068 6020
rect 7080 3490 7092 4460
rect 7104 3706 7116 6020
rect 7128 4306 7140 6020
rect 7152 5314 7164 6020
rect 7056 1042 7068 2852
rect 7104 1042 7116 2204
rect 7152 1042 7164 5252
rect 7176 1042 7188 3836
rect 7200 3178 7212 6020
rect 7224 2866 7236 4580
rect 7248 1858 7260 6020
rect 7272 3730 7284 6020
rect 7296 4954 7308 6020
rect 7272 1042 7284 3404
rect 7296 1042 7308 3356
rect 7320 1042 7332 4820
rect 7344 3850 7356 6020
rect 7368 5314 7380 6020
rect 7392 6010 7404 6020
rect 7368 1042 7380 4580
rect 7392 1042 7404 5900
rect 7416 1978 7428 3692
rect 7440 2434 7452 6020
rect 7464 4066 7476 6020
rect 7488 5962 7500 6020
rect 7464 1042 7476 3236
rect 7488 1042 7500 4148
rect 7512 1138 7524 5300
rect 7608 4474 7620 6020
rect 7536 3154 7548 3716
rect 7560 1042 7572 3092
rect 7584 1042 7596 2732
rect 7608 1042 7620 4292
rect 7632 1234 7644 4460
rect 7680 1042 7692 4532
rect 7800 1042 7812 3332
rect 7824 1042 7836 3596
rect 7920 1042 7932 2804
rect 7944 1042 7956 3884
rect 7968 1426 7980 6020
rect 8016 3994 8028 6020
rect 8160 5242 8172 6020
rect 8040 1042 8052 4988
rect 8112 1042 8124 5084
rect 8184 3490 8196 5732
rect 8160 1042 8172 3476
rect 8208 2026 8220 6020
rect 8232 5482 8244 6020
rect 8232 1042 8244 4700
rect 8256 4306 8268 6020
rect 8280 4930 8292 6020
rect 8328 4450 8340 6020
rect 8280 1042 8292 2180
rect 8304 1042 8316 4172
rect 8352 2506 8364 6020
rect 8376 4378 8388 6020
rect 8424 4258 8436 6020
rect 8472 5122 8484 6020
rect 8352 1042 8364 2468
rect 8400 1042 8412 3644
rect 8448 1042 8460 3476
rect 8496 1042 8508 3428
rect 8520 1042 8532 5396
rect 8544 3226 8556 6020
rect 8568 1690 8580 6020
rect 8592 2890 8604 6020
rect 8616 3658 8628 6020
rect 8592 1042 8604 2444
rect 8664 1522 8676 6020
rect 8688 1306 8700 6020
rect 8712 4834 8724 6020
rect 8784 6010 8796 6020
rect 8712 1042 8724 4724
rect 8736 1786 8748 4820
rect 8760 1042 8772 2180
rect 8784 1042 8796 2900
rect 8808 1282 8820 6020
rect 8832 1354 8844 6020
rect 8856 3322 8868 6020
rect 8880 2314 8892 6020
rect 8928 2482 8940 6020
rect 8976 5650 8988 6020
rect 8976 1042 8988 3836
rect 9000 1690 9012 6020
rect 9024 2770 9036 6020
rect 9048 3778 9060 6020
rect 9072 3706 9084 6020
rect 9000 1042 9012 1652
rect 9024 1042 9036 2660
rect 9096 1042 9108 3524
rect 9120 2722 9132 6020
rect 9144 3922 9156 6020
rect 9168 3154 9180 6020
rect 9192 3730 9204 6020
rect 9240 5362 9252 6020
rect 9120 1042 9132 2588
rect 9216 1042 9228 1964
rect 9240 1042 9252 3332
rect 9264 1498 9276 6020
rect 9288 1666 9300 5252
rect 9312 4234 9324 6020
rect 9360 5194 9372 6020
rect 9336 2674 9348 4676
rect 9360 1042 9372 5132
rect 9384 3730 9396 6020
rect 9408 3490 9420 6020
rect 9480 5482 9492 6020
rect 9432 2602 9444 4580
rect 9456 3346 9468 5180
rect 9504 4306 9516 6020
rect 9528 4762 9540 6020
rect 9576 5218 9588 6020
rect 9600 3730 9612 6020
rect 9624 3826 9636 6020
rect 9648 3682 9660 6020
rect 9696 1186 9708 6020
rect 9720 2938 9732 6020
rect 9744 2722 9756 6020
rect 9768 5314 9780 6020
rect 9720 1042 9732 2420
rect 9768 1042 9780 5252
rect 9792 2338 9804 5300
rect 9816 1978 9828 6020
rect 9840 3010 9852 6020
rect 9864 3106 9876 6020
rect 9888 5626 9900 6020
rect 9936 5290 9948 6020
rect 9912 1042 9924 3476
rect 9960 3418 9972 6020
rect 9984 3682 9996 6020
rect 10032 3322 10044 6020
rect 10080 4618 10092 6020
rect 10152 5866 10164 6020
rect 10104 3418 10116 5732
rect 10176 4522 10188 6020
rect 10200 5842 10212 6020
rect 10008 1042 10020 2252
rect 10032 1042 10044 1724
rect 10080 1042 10092 3404
rect 10128 1042 10140 4100
rect 10248 1402 10260 6020
rect 10296 3730 10308 6020
rect 10344 3850 10356 6020
rect 10368 1282 10380 6020
rect 10392 3298 10404 6020
rect 10416 3202 10428 6020
rect 10464 3538 10476 6020
rect 10488 2026 10500 6020
rect 10512 2698 10524 6020
rect 10560 2506 10572 6020
rect 10584 5746 10596 6020
rect 10608 3274 10620 6020
rect 10656 4906 10668 6020
rect 10680 4330 10692 6020
rect 10704 3946 10716 6020
rect 10752 5506 10764 6020
rect 10776 3682 10788 6020
rect 10800 3322 10812 6020
rect 10824 3562 10836 6020
rect 10872 5578 10884 6020
rect 10656 1042 10668 2924
rect 10824 1042 10836 2516
rect 10848 1042 10860 5060
rect 10896 4090 10908 6020
rect 10920 5434 10932 6020
rect 10896 1042 10908 4004
rect 10920 1042 10932 5396
rect 10944 2554 10956 6020
rect 10968 5986 10980 6020
rect 11016 4066 11028 6020
rect 11040 3442 11052 6020
rect 10992 1042 11004 3092
rect 11040 1042 11052 2828
rect 11064 1642 11076 6020
rect 11088 4282 11100 6020
rect 11136 4306 11148 6020
rect 11160 3370 11172 6020
rect 11112 1042 11124 1796
rect 11136 1042 11148 2804
rect 11184 2722 11196 6020
rect 11208 2026 11220 6020
rect 11232 5506 11244 6020
rect 11280 5386 11292 6020
rect 11208 1042 11220 1268
rect 11256 1042 11268 3572
rect 11304 3562 11316 6020
rect 11304 1042 11316 2636
rect 11328 1042 11340 5924
rect 11352 1042 11364 4412
rect 11376 2002 11388 6020
rect 11400 4210 11412 6020
rect 11424 5458 11436 6020
rect 11400 1042 11412 3404
rect 11424 1042 11436 5396
rect 11472 5050 11484 6020
rect 11448 2626 11460 4076
rect 11472 1042 11484 4988
rect 11496 3898 11508 6020
rect 11544 4498 11556 6020
rect 11520 1042 11532 4484
rect 11592 3850 11604 6020
rect 11556 1786 11568 3548
rect 11616 2938 11628 6020
rect 11664 4906 11676 6020
rect 11688 3418 11700 5948
rect 11676 2914 11688 3140
rect 11616 1042 11628 2900
rect 11640 1042 11652 2804
rect 11712 2530 11724 6020
rect 11736 4906 11748 6020
rect 11736 1042 11748 2972
rect 11760 2746 11772 6020
rect 11760 1042 11772 2708
rect 11784 1762 11796 6020
rect 11784 1042 11796 1724
rect 11808 1594 11820 5420
rect 11832 4042 11844 6020
rect 11856 4594 11868 6020
rect 11832 1042 11844 3524
rect 11856 1042 11868 4556
rect 11880 1042 11892 5708
rect 11904 1162 11916 5444
rect 11928 3058 11940 6020
rect 11952 5266 11964 6020
rect 11928 1042 11940 2924
rect 11952 1042 11964 2036
rect 11976 1570 11988 6020
rect 11976 1042 11988 1532
rect 12000 1042 12012 5540
rect 12024 3610 12036 6020
rect 12048 1042 12060 4844
rect 12072 4138 12084 6020
rect 12072 1042 12084 3836
rect 12096 1042 12108 4388
rect 12120 3466 12132 5036
rect 12144 4066 12156 6020
rect 12144 1042 12156 3428
rect 12168 2938 12180 6020
rect 12168 1042 12180 2516
rect 12192 1042 12204 4340
rect 12216 2746 12228 6020
rect 12240 5026 12252 6020
rect 12240 1042 12252 4796
rect 12264 2722 12276 5900
rect 12312 3922 12324 6020
rect 12336 3394 12348 6020
rect 12384 4882 12396 6020
rect 12432 4666 12444 6020
rect 12456 5602 12468 6020
rect 12480 4978 12492 6020
rect 12528 4498 12540 6020
rect 12288 1042 12300 1844
rect 12360 1042 12372 3788
rect 12408 1042 12420 3524
rect 12492 1738 12504 3620
rect 12552 3490 12564 6020
rect 12576 3826 12588 6020
rect 12600 3514 12612 4580
rect 12624 3754 12636 6020
rect 12648 3778 12660 6020
rect 12672 3538 12684 6020
rect 12696 1546 12708 4772
rect 12720 1378 12732 6020
rect 12852 5517 12922 5529
rect 12744 1066 12756 3644
rect 12768 1090 12780 5156
rect 12852 3693 12922 3705
rect 12852 1077 12922 1089
rect 12852 1053 12922 1065
rect -11976 -727 -11964 243
rect -11736 -727 -11724 243
rect -11184 -703 -11172 243
rect -12183 -740 -12113 -728
rect -10848 -751 -10836 243
rect -10800 -751 -10788 243
rect -10704 -679 -10692 243
rect -10560 -655 -10548 243
rect -10416 -631 -10404 243
rect -10368 -607 -10356 243
rect -10320 -583 -10308 243
rect -10272 -559 -10260 243
rect -10152 -535 -10140 243
rect -9552 -511 -9540 243
rect -9504 -487 -9492 243
rect -9312 -463 -9300 243
rect -9240 -439 -9228 243
rect -9216 -415 -9204 243
rect -9144 -391 -9132 243
rect -9120 -367 -9108 243
rect -9048 -343 -9036 243
rect -9024 -319 -9012 243
rect -8784 -295 -8772 243
rect -8736 -271 -8724 243
rect -8712 -247 -8700 243
rect -8688 -487 -8676 243
rect -7680 -487 -7668 243
rect -7608 -223 -7596 243
rect -7560 -199 -7548 243
rect -7536 -175 -7524 243
rect -7416 -151 -7404 243
rect -7224 -223 -7212 243
rect -7176 -223 -7164 243
rect -7152 -127 -7140 243
rect -7128 -727 -7116 243
rect -7080 -727 -7068 243
rect -7056 -103 -7044 243
rect -6960 -79 -6948 243
rect -6936 -367 -6924 243
rect -6888 -367 -6876 243
rect -6792 -55 -6780 243
rect -6672 -31 -6660 243
rect -12183 -764 -12113 -752
rect -6624 -775 -6612 243
rect -6552 -7 -6540 243
rect -6384 17 -6372 243
rect -6336 41 -6324 243
rect -6192 65 -6180 243
rect -5904 113 -5892 243
rect -5640 113 -5628 243
rect -5904 -799 -5892 75
rect -5880 -295 -5868 99
rect -5424 -775 -5412 243
rect -5184 -7 -5172 243
rect -5064 -727 -5052 243
rect -4920 -463 -4908 243
rect -4728 -415 -4716 243
rect -4704 -463 -4692 243
rect -4560 -79 -4548 243
rect -4488 -607 -4476 243
rect -4440 -655 -4428 243
rect -4368 -79 -4356 243
rect -4344 -31 -4332 243
rect -4320 -415 -4308 243
rect -4296 17 -4284 243
rect -4032 -31 -4020 243
rect -4008 17 -3996 243
rect -3984 -607 -3972 243
rect -3840 -655 -3828 243
rect -3792 137 -3780 243
rect -3720 -79 -3708 243
rect -3600 17 -3588 243
rect -3528 -55 -3516 243
rect -3480 -79 -3468 243
rect -3360 -7 -3348 243
rect -3144 -583 -3132 243
rect -2880 -199 -2868 243
rect -2784 -199 -2772 243
rect -2568 -631 -2556 243
rect -2352 -55 -2340 243
rect -2208 -415 -2196 243
rect -1464 17 -1452 243
rect -1176 -415 -1164 243
rect -1080 161 -1068 243
rect -1032 185 -1020 243
rect -960 65 -948 243
rect -816 209 -804 243
rect -432 233 -420 243
rect -408 113 -396 243
rect -384 -79 -372 243
rect -288 -7 -276 243
rect -264 -79 -252 243
rect -48 -511 -36 243
rect -24 209 -12 243
rect 120 -223 132 243
rect 264 -775 276 243
rect 288 -559 300 243
rect 312 -223 324 243
rect 336 -7 348 243
rect -5868 -799 -5856 -789
rect 336 -799 348 -501
rect 408 -583 420 243
rect 504 17 516 243
rect 552 -55 564 243
rect 576 17 588 243
rect 600 -55 612 243
rect 768 113 780 243
rect 816 209 828 243
rect 888 -655 900 243
rect 912 -55 924 243
rect 960 -535 972 243
rect 1008 -55 1020 243
rect 1392 -487 1404 243
rect 1536 -511 1548 243
rect 1944 17 1956 243
rect 2136 -487 2148 243
rect 2184 161 2196 243
rect 2328 -247 2340 243
rect 2400 185 2412 243
rect 2616 -151 2628 243
rect 2688 -247 2700 243
rect 2760 -151 2772 243
rect 2784 17 2796 243
rect 2856 185 2868 243
rect 2928 -55 2940 243
rect 3000 65 3012 243
rect 3024 161 3036 243
rect 3048 233 3060 243
rect 3144 41 3156 243
rect 3288 -271 3300 243
rect 3336 -463 3348 243
rect 3384 -271 3396 243
rect 3480 -7 3492 243
rect 3576 -103 3588 243
rect 3672 113 3684 243
rect 3768 -103 3780 243
rect 3816 -295 3828 243
rect 3984 137 3996 243
rect 4560 -751 4572 243
rect 4968 -511 4980 243
rect 5328 -55 5340 243
rect 5376 -199 5388 243
rect 5424 -199 5436 243
rect 5760 -607 5772 243
rect 6384 -631 6396 243
rect 6408 -31 6420 243
rect 6576 -31 6588 243
rect 7200 -295 7212 243
rect 7224 185 7236 243
rect 7416 -343 7428 243
rect 7512 -727 7524 243
rect 7632 -703 7644 243
rect 7728 -79 7740 243
rect 7872 161 7884 243
rect 7992 -31 8004 243
rect 8064 17 8076 243
rect 8184 -487 8196 243
rect 8424 -319 8436 243
rect 8544 -127 8556 243
rect 8640 -391 8652 243
rect 8736 -391 8748 243
rect 8808 -127 8820 243
rect 8856 -175 8868 243
rect 8904 -679 8916 243
rect 9072 -295 9084 243
rect 9144 -223 9156 243
rect 9192 -583 9204 243
rect 9912 -223 9924 243
rect 9960 -127 9972 243
rect 9925 -237 9943 -223
rect 9924 -799 9936 -237
rect 9984 -271 9996 243
rect 10104 -103 10116 243
rect 10248 -199 10260 243
rect 10608 -151 10620 243
rect 10800 -631 10812 243
rect 10944 -55 10956 243
rect 11160 -415 11172 243
rect 11232 -391 11244 243
rect 11544 89 11556 243
rect 11568 209 11580 243
rect 11688 -439 11700 243
rect 12360 -271 12372 243
rect 12408 -223 12420 243
rect 12408 -775 12420 -381
rect 12432 -751 12444 -285
rect 12456 -727 12468 -237
rect 12852 -260 12922 -248
rect 12852 -740 12922 -728
rect 12852 -764 12922 -752
rect 12852 -788 12922 -776
use nand2  g8541
timestamp 1395695751
transform 1 0 -12096 0 1 6020
box -10 0 100 799
use nor2  g8462
timestamp 1395695751
transform 1 0 -12000 0 1 6020
box -3 0 125 799
use nand3  g8469
timestamp 1395695751
transform 1 0 -11880 0 1 6020
box -10 0 127 799
use inv  g8513
timestamp 1395695751
transform 1 0 -11760 0 1 6020
box 0 0 120 799
use inv  g8639
timestamp 1395695751
transform 1 0 -11640 0 1 6020
box 0 0 120 799
use nor2  g8774
timestamp 1395695751
transform 1 0 -11520 0 1 6020
box -3 0 125 799
use inv  g8756
timestamp 1395695751
transform 1 0 -11400 0 1 6020
box 0 0 120 799
use nand2  g8642
timestamp 1395695751
transform 1 0 -11280 0 1 6020
box -10 0 100 799
use nand2  g8545
timestamp 1395695751
transform 1 0 -11184 0 1 6020
box -10 0 100 799
use nand2  g8536
timestamp 1395695751
transform 1 0 -11088 0 1 6020
box -10 0 100 799
use nand3  g8724
timestamp 1395695751
transform 1 0 -10992 0 1 6020
box -10 0 127 799
use nand2  g8554
timestamp 1395695751
transform 1 0 -10872 0 1 6020
box -10 0 100 799
use nand2  g8477
timestamp 1395695751
transform 1 0 -10776 0 1 6020
box -10 0 100 799
use nand3  g8506
timestamp 1395695751
transform 1 0 -10680 0 1 6020
box -10 0 127 799
use nand2  g8758
timestamp 1395695751
transform 1 0 -10560 0 1 6020
box -10 0 100 799
use nand2  g8567
timestamp 1395695751
transform 1 0 -10464 0 1 6020
box -10 0 100 799
use nand2  g8623
timestamp 1395695751
transform 1 0 -10368 0 1 6020
box -10 0 100 799
use nor2  g8474
timestamp 1395695751
transform 1 0 -10272 0 1 6020
box -3 0 125 799
use nand2  g8585
timestamp 1395695751
transform 1 0 -10152 0 1 6020
box -10 0 100 799
use nand2  g8640
timestamp 1395695751
transform 1 0 -10056 0 1 6020
box -10 0 100 799
use inv  g8584
timestamp 1395695751
transform 1 0 -9960 0 1 6020
box 0 0 120 799
use inv  g8603
timestamp 1395695751
transform 1 0 -9840 0 1 6020
box 0 0 120 799
use and2  g8597
timestamp 1395695751
transform 1 0 -9720 0 1 6020
box -10 0 127 799
use nand2  g8472
timestamp 1395695751
transform 1 0 -9600 0 1 6020
box -10 0 100 799
use nor2  g8712
timestamp 1395695751
transform 1 0 -9504 0 1 6020
box -3 0 125 799
use mux2  g8655
timestamp 1395695751
transform 1 0 -9384 0 1 6020
box -4 0 195 799
use and2  g8749
timestamp 1395695751
transform 1 0 -9192 0 1 6020
box -10 0 127 799
use inv  g8741
timestamp 1395695751
transform 1 0 -9072 0 1 6020
box 0 0 120 799
use inv  g8572
timestamp 1395695751
transform 1 0 -8952 0 1 6020
box 0 0 120 799
use nand2  g8772
timestamp 1395695751
transform 1 0 -8832 0 1 6020
box -10 0 100 799
use inv  g8763
timestamp 1395695751
transform 1 0 -8736 0 1 6020
box 0 0 120 799
use inv  g8729
timestamp 1395695751
transform 1 0 -8616 0 1 6020
box 0 0 120 799
use nand2  g8761
timestamp 1395695751
transform 1 0 -8496 0 1 6020
box -10 0 100 799
use nand2  g8456
timestamp 1395695751
transform 1 0 -8400 0 1 6020
box -10 0 100 799
use nand4  g8450
timestamp 1395695751
transform 1 0 -8304 0 1 6020
box -10 0 154 799
use nand2  g8589
timestamp 1395695751
transform 1 0 -8160 0 1 6020
box -10 0 100 799
use inv  g8645
timestamp 1395695751
transform 1 0 -8064 0 1 6020
box 0 0 120 799
use nand2  g8649
timestamp 1395695751
transform 1 0 -7944 0 1 6020
box -10 0 100 799
use nand3  g8616
timestamp 1395695751
transform 1 0 -7848 0 1 6020
box -10 0 127 799
use and2  g8690
timestamp 1395695751
transform 1 0 -7728 0 1 6020
box -10 0 127 799
use inv  g8683
timestamp 1395695751
transform 1 0 -7608 0 1 6020
box 0 0 120 799
use nand2  g8667
timestamp 1395695751
transform 1 0 -7488 0 1 6020
box -10 0 100 799
use nor2  g8547
timestamp 1395695751
transform 1 0 -7392 0 1 6020
box -3 0 125 799
use nand2  g8493
timestamp 1395695751
transform 1 0 -7272 0 1 6020
box -10 0 100 799
use nand2  g8440
timestamp 1395695751
transform 1 0 -7176 0 1 6020
box -10 0 100 799
use rowcrosser  AluWe
timestamp 1395695751
transform 1 0 -7080 0 1 6020
box 0 0 48 799
use inv  g8504
timestamp 1395695751
transform 1 0 -7032 0 1 6020
box 0 0 120 799
use nand2  g8449
timestamp 1395695751
transform 1 0 -6912 0 1 6020
box -10 0 100 799
use nand2  g8414
timestamp 1395695751
transform 1 0 -6816 0 1 6020
box -10 0 100 799
use nand3  g8418
timestamp 1395695751
transform 1 0 -6720 0 1 6020
box -10 0 127 799
use nand2  g8636
timestamp 1395695751
transform 1 0 -6600 0 1 6020
box -10 0 100 799
use nand3  g8651
timestamp 1395695751
transform 1 0 -6504 0 1 6020
box -10 0 127 799
use rowcrosser  StatusRegEn
timestamp 1395695751
transform 1 0 -6384 0 1 6020
box 0 0 48 799
use nand2  g8620
timestamp 1395695751
transform 1 0 -6336 0 1 6020
box -10 0 100 799
use nand2  g8483
timestamp 1395695751
transform 1 0 -6240 0 1 6020
box -10 0 100 799
use nand2  g8717
timestamp 1395695751
transform 1 0 -6144 0 1 6020
box -10 0 100 799
use nand2  g8666
timestamp 1395695751
transform 1 0 -6048 0 1 6020
box -10 0 100 799
use nor2  g8511
timestamp 1395695751
transform 1 0 -5952 0 1 6020
box -3 0 125 799
use nand2  g8696
timestamp 1395695751
transform 1 0 -5832 0 1 6020
box -10 0 100 799
use nand2  g8407
timestamp 1395695751
transform 1 0 -5736 0 1 6020
box -10 0 100 799
use nand3  g8486
timestamp 1395695751
transform 1 0 -5640 0 1 6020
box -10 0 127 799
use nand2  g8618
timestamp 1395695751
transform 1 0 -5520 0 1 6020
box -10 0 100 799
use nand3  g8562
timestamp 1395695751
transform 1 0 -5424 0 1 6020
box -10 0 127 799
use nand2  g8703
timestamp 1395695751
transform 1 0 -5304 0 1 6020
box -10 0 100 799
use and2  g8489
timestamp 1395695751
transform 1 0 -5208 0 1 6020
box -10 0 127 799
use rowcrosser  IrWe
timestamp 1395695751
transform 1 0 -5088 0 1 6020
box 0 0 48 799
use nand2  g8723
timestamp 1395695751
transform 1 0 -5040 0 1 6020
box -10 0 100 799
use inv  g8735
timestamp 1395695751
transform 1 0 -4944 0 1 6020
box 0 0 120 799
use rowcrosser  ALE
timestamp 1395695751
transform 1 0 -4824 0 1 6020
box 0 0 48 799
use nand2  g8403
timestamp 1395695751
transform 1 0 -4776 0 1 6020
box -10 0 100 799
use nand2  g8612
timestamp 1395695751
transform 1 0 -4680 0 1 6020
box -10 0 100 799
use nand2  g8631
timestamp 1395695751
transform 1 0 -4584 0 1 6020
box -10 0 100 799
use inv  g8532
timestamp 1395695751
transform 1 0 -4488 0 1 6020
box 0 0 120 799
use nand3  g8529
timestamp 1395695751
transform 1 0 -4368 0 1 6020
box -10 0 127 799
use nand3  g8676
timestamp 1395695751
transform 1 0 -4248 0 1 6020
box -10 0 127 799
use nand2  g8538
timestamp 1395695751
transform 1 0 -4128 0 1 6020
box -10 0 100 799
use nand2  g8580
timestamp 1395695751
transform 1 0 -4032 0 1 6020
box -10 0 100 799
use nand3  g8594
timestamp 1395695751
transform 1 0 -3936 0 1 6020
box -10 0 127 799
use nand2  g8648
timestamp 1395695751
transform 1 0 -3816 0 1 6020
box -10 0 100 799
use nand2  g8425
timestamp 1395695751
transform 1 0 -3720 0 1 6020
box -10 0 100 799
use nand3  g8524
timestamp 1395695751
transform 1 0 -3624 0 1 6020
box -10 0 127 799
use nand2  g8609
timestamp 1395695751
transform 1 0 -3504 0 1 6020
box -10 0 100 799
use nor2  g8743
timestamp 1395695751
transform 1 0 -3408 0 1 6020
box -3 0 125 799
use rowcrosser  Flags_91_2_93_
timestamp 1395695751
transform 1 0 -3288 0 1 6020
box 0 0 48 799
use nor2  g8479
timestamp 1395695751
transform 1 0 -3240 0 1 6020
box -3 0 125 799
use nand2  g8728
timestamp 1395695751
transform 1 0 -3120 0 1 6020
box -10 0 100 799
use nor2  g8564
timestamp 1395695751
transform 1 0 -3024 0 1 6020
box -3 0 125 799
use nand2  g8699
timestamp 1395695751
transform 1 0 -2904 0 1 6020
box -10 0 100 799
use and2  g8694
timestamp 1395695751
transform 1 0 -2808 0 1 6020
box -10 0 127 799
use nand2  g8533
timestamp 1395695751
transform 1 0 -2688 0 1 6020
box -10 0 100 799
use mux2  g8700
timestamp 1395695751
transform 1 0 -2592 0 1 6020
box -4 0 195 799
use rowcrosser  WdSel
timestamp 1395695751
transform 1 0 -2400 0 1 6020
box 0 0 48 799
use inv  g8627
timestamp 1395695751
transform 1 0 -2352 0 1 6020
box 0 0 120 799
use and2  g8634
timestamp 1395695751
transform 1 0 -2232 0 1 6020
box -10 0 127 799
use nand2  g8731
timestamp 1395695751
transform 1 0 -2112 0 1 6020
box -10 0 100 799
use inv  g8746
timestamp 1395695751
transform 1 0 -2016 0 1 6020
box 0 0 120 799
use nand2  g8705
timestamp 1395695751
transform 1 0 -1896 0 1 6020
box -10 0 100 799
use nand2  g8431
timestamp 1395695751
transform 1 0 -1800 0 1 6020
box -10 0 100 799
use nor2  rm_assigns_buf_StatusReg_1
timestamp 1395695751
transform 1 0 -1704 0 1 6020
box -3 0 125 799
use buffer  g8421
timestamp 1395695751
transform 1 0 -1584 0 1 6020
box -5 0 120 799
use nor2  g8399
timestamp 1395695751
transform 1 0 -1464 0 1 6020
box -3 0 125 799
use nand4  g8778
timestamp 1395695751
transform 1 0 -1344 0 1 6020
box -10 0 154 799
use inv  g8507
timestamp 1395695751
transform 1 0 -1200 0 1 6020
box 0 0 120 799
use nand2  g8688
timestamp 1395695751
transform 1 0 -1080 0 1 6020
box -10 0 100 799
use nand3  g8411
timestamp 1395695751
transform 1 0 -984 0 1 6020
box -10 0 127 799
use nor2  g8553
timestamp 1395695751
transform 1 0 -864 0 1 6020
box -3 0 125 799
use inv  g8646
timestamp 1395695751
transform 1 0 -744 0 1 6020
box 0 0 120 799
use rowcrosser  PcEn
timestamp 1395695751
transform 1 0 -624 0 1 6020
box 0 0 48 799
use nand2  g8417
timestamp 1395695751
transform 1 0 -576 0 1 6020
box -10 0 100 799
use nand2  g8658
timestamp 1395695751
transform 1 0 -480 0 1 6020
box -10 0 100 799
use nand3  g8698
timestamp 1395695751
transform 1 0 -384 0 1 6020
box -10 0 127 799
use and2  g8641
timestamp 1395695751
transform 1 0 -264 0 1 6020
box -10 0 127 799
use nand2  StatusReg_reg_91_3_93_
timestamp 1395695751
transform 1 0 -144 0 1 6020
box -10 0 100 799
use scandtype  stateSub_reg_91_2_93_
timestamp 1395695751
transform 1 0 -48 0 1 6020
box -9 0 624 799
use scandtype  g8546
timestamp 1395695751
transform 1 0 576 0 1 6020
box -9 0 624 799
use nand2  g8750
timestamp 1395695751
transform 1 0 1200 0 1 6020
box -10 0 100 799
use nand2  g8444
timestamp 1395695751
transform 1 0 1296 0 1 6020
box -10 0 100 799
use nand4  g8466
timestamp 1395695751
transform 1 0 1392 0 1 6020
box -10 0 154 799
use nand4  g8468
timestamp 1395695751
transform 1 0 1536 0 1 6020
box -10 0 154 799
use nand4  g8433
timestamp 1395695751
transform 1 0 1680 0 1 6020
box -10 0 154 799
use nand4  g8420
timestamp 1395695751
transform 1 0 1824 0 1 6020
box -10 0 154 799
use nand4  g8624
timestamp 1395695751
transform 1 0 1968 0 1 6020
box -10 0 154 799
use nand2  g8668
timestamp 1395695751
transform 1 0 2112 0 1 6020
box -10 0 100 799
use and2  g8733
timestamp 1395695751
transform 1 0 2208 0 1 6020
box -10 0 127 799
use nor2  g8537
timestamp 1395695751
transform 1 0 2328 0 1 6020
box -3 0 125 799
use nor2  g8531
timestamp 1395695751
transform 1 0 2448 0 1 6020
box -3 0 125 799
use nand3  g8542
timestamp 1395695751
transform 1 0 2568 0 1 6020
box -10 0 127 799
use nand4  g8754
timestamp 1395695751
transform 1 0 2688 0 1 6020
box -10 0 154 799
use nor2  g8760
timestamp 1395695751
transform 1 0 2832 0 1 6020
box -3 0 125 799
use nand2  StatusReg_reg_91_1_93_
timestamp 1395695751
transform 1 0 2952 0 1 6020
box -10 0 100 799
use scandtype  g8435
timestamp 1395695751
transform 1 0 3048 0 1 6020
box -9 0 624 799
use rowcrosser  LrWe
timestamp 1395695751
transform 1 0 3672 0 1 6020
box 0 0 48 799
use nand4  g8452
timestamp 1395695751
transform 1 0 3720 0 1 6020
box -10 0 154 799
use nand2  g8710
timestamp 1395695751
transform 1 0 3864 0 1 6020
box -10 0 100 799
use nand2  g8610
timestamp 1395695751
transform 1 0 3960 0 1 6020
box -10 0 100 799
use nand2  g8635
timestamp 1395695751
transform 1 0 4056 0 1 6020
box -10 0 100 799
use nor2  g8713
timestamp 1395695751
transform 1 0 4152 0 1 6020
box -3 0 125 799
use rowcrosser  ImmSel
timestamp 1395695751
transform 1 0 4272 0 1 6020
box 0 0 48 799
use xor2  g8604
timestamp 1395695751
transform 1 0 4320 0 1 6020
box -3 0 202 799
use nand2  g8691
timestamp 1395695751
transform 1 0 4512 0 1 6020
box -10 0 100 799
use nand2  g8522
timestamp 1395695751
transform 1 0 4608 0 1 6020
box -10 0 100 799
use and2  g8656
timestamp 1395695751
transform 1 0 4704 0 1 6020
box -10 0 127 799
use inv  g8535
timestamp 1395695751
transform 1 0 4824 0 1 6020
box 0 0 120 799
use nand3  g8516
timestamp 1395695751
transform 1 0 4944 0 1 6020
box -10 0 127 799
use nand2  g8514
timestamp 1395695751
transform 1 0 5064 0 1 6020
box -10 0 100 799
use nand2  g8673
timestamp 1395695751
transform 1 0 5160 0 1 6020
box -10 0 100 799
use nand2  g8559
timestamp 1395695751
transform 1 0 5256 0 1 6020
box -10 0 100 799
use nand2  g8748
timestamp 1395695751
transform 1 0 5352 0 1 6020
box -10 0 100 799
use nand2  g8718
timestamp 1395695751
transform 1 0 5448 0 1 6020
box -10 0 100 799
use nor2  g8590
timestamp 1395695751
transform 1 0 5544 0 1 6020
box -3 0 125 799
use nand3  g8670
timestamp 1395695751
transform 1 0 5664 0 1 6020
box -10 0 127 799
use nor2  g8619
timestamp 1395695751
transform 1 0 5784 0 1 6020
box -3 0 125 799
use nand3  g8599
timestamp 1395695751
transform 1 0 5904 0 1 6020
box -10 0 127 799
use inv  g8480
timestamp 1395695751
transform 1 0 6024 0 1 6020
box 0 0 120 799
use nand2  g8436
timestamp 1395695751
transform 1 0 6144 0 1 6020
box -10 0 100 799
use nand2  g8586
timestamp 1395695751
transform 1 0 6240 0 1 6020
box -10 0 100 799
use nand2  g8548
timestamp 1395695751
transform 1 0 6336 0 1 6020
box -10 0 100 799
use nand2  g8740
timestamp 1395695751
transform 1 0 6432 0 1 6020
box -10 0 100 799
use nor2  g8653
timestamp 1395695751
transform 1 0 6528 0 1 6020
box -3 0 125 799
use nand2  g8595
timestamp 1395695751
transform 1 0 6648 0 1 6020
box -10 0 100 799
use nand2  g8720
timestamp 1395695751
transform 1 0 6744 0 1 6020
box -10 0 100 799
use nand2  g8573
timestamp 1395695751
transform 1 0 6840 0 1 6020
box -10 0 100 799
use rowcrosser  rowcrosser_0
timestamp 1395695751
transform 1 0 6936 0 1 6020
box 0 0 48 799
use nand2  g8701
timestamp 1395695751
transform 1 0 6984 0 1 6020
box -10 0 100 799
use nand2  g8674
timestamp 1395695751
transform 1 0 7080 0 1 6020
box -10 0 100 799
use rowcrosser  Flags_91_1_93_
timestamp 1395695751
transform 1 0 7176 0 1 6020
box 0 0 48 799
use nand2  g8630
timestamp 1395695751
transform 1 0 7224 0 1 6020
box -10 0 100 799
use nand2  g8732
timestamp 1395695751
transform 1 0 7320 0 1 6020
box -10 0 100 799
use nand2  StatusReg_reg_91_0_93_
timestamp 1395695751
transform 1 0 7416 0 1 6020
box -10 0 100 799
use scandtype  g8591
timestamp 1395695751
transform 1 0 7512 0 1 6020
box -9 0 624 799
use rowcrosser  AluEn
timestamp 1395695751
transform 1 0 8136 0 1 6020
box 0 0 48 799
use nand3  g8702
timestamp 1395695751
transform 1 0 8184 0 1 6020
box -10 0 127 799
use nand2  g8443
timestamp 1395695751
transform 1 0 8304 0 1 6020
box -10 0 100 799
use inv  g8427
timestamp 1395695751
transform 1 0 8400 0 1 6020
box 0 0 120 799
use nand3  g8432
timestamp 1395695751
transform 1 0 8520 0 1 6020
box -10 0 127 799
use nand3  g8424
timestamp 1395695751
transform 1 0 8640 0 1 6020
box -10 0 127 799
use nand4  g8410
timestamp 1395695751
transform 1 0 8760 0 1 6020
box -10 0 154 799
use rowcrosser  Op2Sel_91_1_93_
timestamp 1395695751
transform 1 0 8904 0 1 6020
box 0 0 48 799
use nand4  g8503
timestamp 1395695751
transform 1 0 8952 0 1 6020
box -10 0 154 799
use nand3  g8588
timestamp 1395695751
transform 1 0 9096 0 1 6020
box -10 0 127 799
use nor2  g8495
timestamp 1395695751
transform 1 0 9216 0 1 6020
box -3 0 125 799
use nand3  g8659
timestamp 1395695751
transform 1 0 9336 0 1 6020
box -10 0 127 799
use nand2  g8406
timestamp 1395695751
transform 1 0 9456 0 1 6020
box -10 0 100 799
use nand3  g8487
timestamp 1395695751
transform 1 0 9552 0 1 6020
box -10 0 127 799
use nand3  g8508
timestamp 1395695751
transform 1 0 9672 0 1 6020
box -10 0 127 799
use nand3  g8563
timestamp 1395695751
transform 1 0 9792 0 1 6020
box -10 0 127 799
use nand2  g8677
timestamp 1395695751
transform 1 0 9912 0 1 6020
box -10 0 100 799
use inv  g8706
timestamp 1395695751
transform 1 0 10008 0 1 6020
box 0 0 120 799
use nand2  g8439
timestamp 1395695751
transform 1 0 10128 0 1 6020
box -10 0 100 799
use nand2  g8473
timestamp 1395695751
transform 1 0 10224 0 1 6020
box -10 0 100 799
use nand3  g8600
timestamp 1395695751
transform 1 0 10320 0 1 6020
box -10 0 127 799
use nand2  g8695
timestamp 1395695751
transform 1 0 10440 0 1 6020
box -10 0 100 799
use nand2  g8637
timestamp 1395695751
transform 1 0 10536 0 1 6020
box -10 0 100 799
use nand2  g8494
timestamp 1395695751
transform 1 0 10632 0 1 6020
box -10 0 100 799
use nand3  g8465
timestamp 1395695751
transform 1 0 10728 0 1 6020
box -10 0 127 799
use nand4  g8523
timestamp 1395695751
transform 1 0 10848 0 1 6020
box -10 0 154 799
use nand3  g8615
timestamp 1395695751
transform 1 0 10992 0 1 6020
box -10 0 127 799
use nand4  g8455
timestamp 1395695751
transform 1 0 11112 0 1 6020
box -10 0 154 799
use nand2  g8650
timestamp 1395695751
transform 1 0 11256 0 1 6020
box -10 0 100 799
use nand2  g8478
timestamp 1395695751
transform 1 0 11352 0 1 6020
box -10 0 100 799
use and2  g8744
timestamp 1395695751
transform 1 0 11448 0 1 6020
box -10 0 127 799
use and2  g8663
timestamp 1395695751
transform 1 0 11568 0 1 6020
box -10 0 127 799
use nand3  g8447
timestamp 1395695751
transform 1 0 11688 0 1 6020
box -10 0 127 799
use nand2  g8575
timestamp 1395695751
transform 1 0 11808 0 1 6020
box -10 0 100 799
use nand2  g8759
timestamp 1395695751
transform 1 0 11904 0 1 6020
box -10 0 100 799
use nand2  g8714
timestamp 1395695751
transform 1 0 12000 0 1 6020
box -10 0 100 799
use mux2  g8540
timestamp 1395695751
transform 1 0 12096 0 1 6020
box -4 0 195 799
use and2  g8510
timestamp 1395695751
transform 1 0 12288 0 1 6020
box -10 0 127 799
use nand2  g8451
timestamp 1395695751
transform 1 0 12408 0 1 6020
box -10 0 100 799
use nand2  g8519
timestamp 1395695751
transform 1 0 12504 0 1 6020
box -10 0 100 799
use nand2  LrSel
timestamp 1395695751
transform 1 0 12600 0 1 6020
box -10 0 100 799
use rowcrosser  LrEn
timestamp 1395695751
transform 1 0 12696 0 1 6020
box 0 0 48 799
use nand2  g8747
timestamp 1395695751
transform 1 0 -12096 0 1 243
box -10 0 100 799
use rowcrosser  g8737
timestamp 1395695751
transform 1 0 -12000 0 1 243
box 0 0 48 799
use and2  stateSub_reg_91_0_93_
timestamp 1395695751
transform 1 0 -11952 0 1 243
box -10 0 127 799
use scandtype  g8625
timestamp 1395695751
transform 1 0 -11832 0 1 243
box -9 0 624 799
use nand2  g8552
timestamp 1395695751
transform 1 0 -11208 0 1 243
box -10 0 100 799
use nor2  g8558
timestamp 1395695751
transform 1 0 -11112 0 1 243
box -3 0 125 799
use and2  g8777
timestamp 1395695751
transform 1 0 -10992 0 1 243
box -10 0 127 799
use inv  g8430
timestamp 1395695751
transform 1 0 -10872 0 1 243
box 0 0 120 799
use nand3  g8697
timestamp 1395695751
transform 1 0 -10752 0 1 243
box -10 0 127 799
use nand2  g8614
timestamp 1395695751
transform 1 0 -10632 0 1 243
box -10 0 100 799
use nand2  g8629
timestamp 1395695751
transform 1 0 -10536 0 1 243
box -10 0 100 799
use nand2  g8543
timestamp 1395695751
transform 1 0 -10440 0 1 243
box -10 0 100 799
use nand2  state_reg_91_1_93_
timestamp 1395695751
transform 1 0 -10344 0 1 243
box -10 0 100 799
use scandtype  g8416
timestamp 1395695751
transform 1 0 -10248 0 1 243
box -9 0 624 799
use nand2  g8434
timestamp 1395695751
transform 1 0 -9624 0 1 243
box -10 0 100 799
use and2  g8578
timestamp 1395695751
transform 1 0 -9528 0 1 243
box -10 0 127 799
use nand3  g8556
timestamp 1395695751
transform 1 0 -9408 0 1 243
box -10 0 127 799
use nand2  g8566
timestamp 1395695751
transform 1 0 -9288 0 1 243
box -10 0 100 799
use nand2  g8611
timestamp 1395695751
transform 1 0 -9192 0 1 243
box -10 0 100 799
use nand2  g8429
timestamp 1395695751
transform 1 0 -9096 0 1 243
box -10 0 100 799
use nand4  g8726
timestamp 1395695751
transform 1 0 -9000 0 1 243
box -10 0 154 799
use nand2  g8458
timestamp 1395695751
transform 1 0 -8856 0 1 243
box -10 0 100 799
use nand2  g8736
timestamp 1395695751
transform 1 0 -8760 0 1 243
box -10 0 100 799
use inv  g8476
timestamp 1395695751
transform 1 0 -8664 0 1 243
box 0 0 120 799
use nor2  g8687
timestamp 1395695751
transform 1 0 -8544 0 1 243
box -3 0 125 799
use nand2  StatusReg_reg_91_2_93_
timestamp 1395695751
transform 1 0 -8424 0 1 243
box -10 0 100 799
use scandtype  g8498
timestamp 1395695751
transform 1 0 -8328 0 1 243
box -9 0 624 799
use rowcrosser  SysBus_91_3_93_
timestamp 1395695751
transform 1 0 -7704 0 1 243
box 0 0 48 799
use nand4  g8501
timestamp 1395695751
transform 1 0 -7656 0 1 243
box -10 0 154 799
use nor2  g8587
timestamp 1395695751
transform 1 0 -7512 0 1 243
box -3 0 125 799
use nand2  g8608
timestamp 1395695751
transform 1 0 -7392 0 1 243
box -10 0 100 799
use nand2  g8534
timestamp 1395695751
transform 1 0 -7296 0 1 243
box -10 0 100 799
use nand2  g8454
timestamp 1395695751
transform 1 0 -7200 0 1 243
box -10 0 100 799
use nand2  g8442
timestamp 1395695751
transform 1 0 -7104 0 1 243
box -10 0 100 799
use nand4  g8680
timestamp 1395695751
transform 1 0 -7008 0 1 243
box -10 0 154 799
use nand2  g8521
timestamp 1395695751
transform 1 0 -6864 0 1 243
box -10 0 100 799
use nand3  g8394
timestamp 1395695751
transform 1 0 -6768 0 1 243
box -10 0 127 799
use rowcrosser  AluOR_91_1_93_
timestamp 1395695751
transform 1 0 -6648 0 1 243
box 0 0 48 799
use nand4  g8692
timestamp 1395695751
transform 1 0 -6600 0 1 243
box -10 0 154 799
use nand2  g8453
timestamp 1395695751
transform 1 0 -6456 0 1 243
box -10 0 100 799
use nand2  g8719
timestamp 1395695751
transform 1 0 -6360 0 1 243
box -10 0 100 799
use nand2  g8644
timestamp 1395695751
transform 1 0 -6264 0 1 243
box -10 0 100 799
use nand2  g8461
timestamp 1395695751
transform 1 0 -6168 0 1 243
box -10 0 100 799
use inv  g8679
timestamp 1395695751
transform 1 0 -6072 0 1 243
box 0 0 120 799
use nand2  g8770
timestamp 1395695751
transform 1 0 -5952 0 1 243
box -10 0 100 799
use inv  g8661
timestamp 1395695751
transform 1 0 -5856 0 1 243
box 0 0 120 799
use nand3  g8776
timestamp 1395695751
transform 1 0 -5736 0 1 243
box -10 0 127 799
use inv  g8550
timestamp 1395695751
transform 1 0 -5616 0 1 243
box 0 0 120 799
use nand2  g8438
timestamp 1395695751
transform 1 0 -5496 0 1 243
box -10 0 100 799
use nand2  g8549
timestamp 1395695751
transform 1 0 -5400 0 1 243
box -10 0 100 799
use nand2  g8412
timestamp 1395695751
transform 1 0 -5304 0 1 243
box -10 0 100 799
use nand3  g8481
timestamp 1395695751
transform 1 0 -5208 0 1 243
box -10 0 127 799
use inv  g8457
timestamp 1395695751
transform 1 0 -5088 0 1 243
box 0 0 120 799
use nand2  g8518
timestamp 1395695751
transform 1 0 -4968 0 1 243
box -10 0 100 799
use nand2  g8515
timestamp 1395695751
transform 1 0 -4872 0 1 243
box -10 0 100 799
use nand2  g8484
timestamp 1395695751
transform 1 0 -4776 0 1 243
box -10 0 100 799
use nand4  g8496
timestamp 1395695751
transform 1 0 -4680 0 1 243
box -10 0 154 799
use nand4  g8470
timestamp 1395695751
transform 1 0 -4536 0 1 243
box -10 0 154 799
use nand4  g8707
timestamp 1395695751
transform 1 0 -4392 0 1 243
box -10 0 154 799
use nand2  g8574
timestamp 1395695751
transform 1 0 -4248 0 1 243
box -10 0 100 799
use nand2  g8426
timestamp 1395695751
transform 1 0 -4152 0 1 243
box -10 0 100 799
use nand4  g8660
timestamp 1395695751
transform 1 0 -4056 0 1 243
box -10 0 154 799
use nand2  g8579
timestamp 1395695751
transform 1 0 -3912 0 1 243
box -10 0 100 799
use nand3  g8509
timestamp 1395695751
transform 1 0 -3816 0 1 243
box -10 0 127 799
use nand3  g8592
timestamp 1395695751
transform 1 0 -3696 0 1 243
box -10 0 127 799
use and2  g8490
timestamp 1395695751
transform 1 0 -3576 0 1 243
box -10 0 127 799
use and2  g8500
timestamp 1395695751
transform 1 0 -3456 0 1 243
box -10 0 127 799
use nor2  g8605
timestamp 1395695751
transform 1 0 -3336 0 1 243
box -3 0 125 799
use inv  g8446
timestamp 1395695751
transform 1 0 -3216 0 1 243
box 0 0 120 799
use and2  g8560
timestamp 1395695751
transform 1 0 -3096 0 1 243
box -10 0 127 799
use nand3  g8459
timestamp 1395695751
transform 1 0 -2976 0 1 243
box -10 0 127 799
use nand2  g8753
timestamp 1395695751
transform 1 0 -2856 0 1 243
box -10 0 100 799
use nand2  g8684
timestamp 1395695751
transform 1 0 -2760 0 1 243
box -10 0 100 799
use and2  g8638
timestamp 1395695751
transform 1 0 -2664 0 1 243
box -10 0 127 799
use inv  g8527
timestamp 1395695751
transform 1 0 -2544 0 1 243
box 0 0 120 799
use nand2  g8570
timestamp 1395695751
transform 1 0 -2424 0 1 243
box -10 0 100 799
use nand4  g8530
timestamp 1395695751
transform 1 0 -2328 0 1 243
box -10 0 154 799
use nand3  IntStatus_reg
timestamp 1395695751
transform 1 0 -2184 0 1 243
box -10 0 127 799
use scanreg  g8745
timestamp 1395695751
transform 1 0 -2064 0 1 243
box -11 0 720 799
use and2  g8491
timestamp 1395695751
transform 1 0 -1344 0 1 243
box -10 0 127 799
use and2  g8721
timestamp 1395695751
transform 1 0 -1224 0 1 243
box -10 0 127 799
use inv  g8715
timestamp 1395695751
transform 1 0 -1104 0 1 243
box 0 0 120 799
use nand2  g8437
timestamp 1395695751
transform 1 0 -984 0 1 243
box -10 0 100 799
use nand2  g8755
timestamp 1395695751
transform 1 0 -888 0 1 243
box -10 0 100 799
use inv  g8752
timestamp 1395695751
transform 1 0 -792 0 1 243
box 0 0 120 799
use nor2  g8678
timestamp 1395695751
transform 1 0 -672 0 1 243
box -3 0 125 799
use nand2  g8526
timestamp 1395695751
transform 1 0 -552 0 1 243
box -10 0 100 799
use nand4  g8423
timestamp 1395695751
transform 1 0 -456 0 1 243
box -10 0 154 799
use nand3  g8601
timestamp 1395695751
transform 1 0 -312 0 1 243
box -10 0 127 799
use and2  g8405
timestamp 1395695751
transform 1 0 -192 0 1 243
box -10 0 127 799
use nand3  g8582
timestamp 1395695751
transform 1 0 -72 0 1 243
box -10 0 127 799
use nand2  g8632
timestamp 1395695751
transform 1 0 48 0 1 243
box -10 0 100 799
use nand2  g8464
timestamp 1395695751
transform 1 0 144 0 1 243
box -10 0 100 799
use nand4  g8568
timestamp 1395695751
transform 1 0 240 0 1 243
box -10 0 154 799
use nand2  g8460
timestamp 1395695751
transform 1 0 384 0 1 243
box -10 0 100 799
use nand4  g8626
timestamp 1395695751
transform 1 0 480 0 1 243
box -10 0 154 799
use and2  g8404
timestamp 1395695751
transform 1 0 624 0 1 243
box -10 0 127 799
use nand3  g8428
timestamp 1395695751
transform 1 0 744 0 1 243
box -10 0 127 799
use nand3  g8413
timestamp 1395695751
transform 1 0 864 0 1 243
box -10 0 127 799
use nor2  g8577
timestamp 1395695751
transform 1 0 984 0 1 243
box -3 0 125 799
use nand3  g8682
timestamp 1395695751
transform 1 0 1104 0 1 243
box -10 0 127 799
use and2  g8571
timestamp 1395695751
transform 1 0 1224 0 1 243
box -10 0 127 799
use nand2  IRQ2_reg
timestamp 1395695751
transform 1 0 1344 0 1 243
box -10 0 100 799
use scandtype  g8602
timestamp 1395695751
transform 1 0 1440 0 1 243
box -9 0 624 799
use nand2  g8669
timestamp 1395695751
transform 1 0 2064 0 1 243
box -10 0 100 799
use nand2  g8593
timestamp 1395695751
transform 1 0 2160 0 1 243
box -10 0 100 799
use nand2  g8686
timestamp 1395695751
transform 1 0 2256 0 1 243
box -10 0 100 799
use nand2  g8517
timestamp 1395695751
transform 1 0 2352 0 1 243
box -10 0 100 799
use inv  g8402
timestamp 1395695751
transform 1 0 2448 0 1 243
box 0 0 120 799
use nand4  g8738
timestamp 1395695751
transform 1 0 2568 0 1 243
box -10 0 154 799
use nand2  g8422
timestamp 1395695751
transform 1 0 2712 0 1 243
box -10 0 100 799
use nand4  g8622
timestamp 1395695751
transform 1 0 2808 0 1 243
box -10 0 154 799
use nand3  g8633
timestamp 1395695751
transform 1 0 2952 0 1 243
box -10 0 127 799
use nand2  g8488
timestamp 1395695751
transform 1 0 3072 0 1 243
box -10 0 100 799
use nand4  g8475
timestamp 1395695751
transform 1 0 3168 0 1 243
box -10 0 154 799
use nand2  g8598
timestamp 1395695751
transform 1 0 3312 0 1 243
box -10 0 100 799
use nand2  g8555
timestamp 1395695751
transform 1 0 3408 0 1 243
box -10 0 100 799
use nand2  g8415
timestamp 1395695751
transform 1 0 3504 0 1 243
box -10 0 100 799
use nand2  g8675
timestamp 1395695751
transform 1 0 3600 0 1 243
box -10 0 100 799
use nand2  g8725
timestamp 1395695751
transform 1 0 3696 0 1 243
box -10 0 100 799
use inv  g8643
timestamp 1395695751
transform 1 0 3792 0 1 243
box 0 0 120 799
use inv  g8742
timestamp 1395695751
transform 1 0 3912 0 1 243
box 0 0 120 799
use nand2  g8520
timestamp 1395695751
transform 1 0 4032 0 1 243
box -10 0 100 799
use nand2  g8708
timestamp 1395695751
transform 1 0 4128 0 1 243
box -10 0 100 799
use and2  g8617
timestamp 1395695751
transform 1 0 4224 0 1 243
box -10 0 127 799
use nand3  IRQ1_reg
timestamp 1395695751
transform 1 0 4344 0 1 243
box -10 0 127 799
use scandtype  g8502
timestamp 1395695751
transform 1 0 4464 0 1 243
box -9 0 624 799
use nand3  g8505
timestamp 1395695751
transform 1 0 5088 0 1 243
box -10 0 127 799
use nand2  g8419
timestamp 1395695751
transform 1 0 5208 0 1 243
box -10 0 100 799
use nand4  g8596
timestamp 1395695751
transform 1 0 5304 0 1 243
box -10 0 154 799
use and2  g8773
timestamp 1395695751
transform 1 0 5448 0 1 243
box -10 0 127 799
use inv  g8463
timestamp 1395695751
transform 1 0 5568 0 1 243
box 0 0 120 799
use inv  g8557
timestamp 1395695751
transform 1 0 5688 0 1 243
box 0 0 120 799
use nand2  g8757
timestamp 1395695751
transform 1 0 5808 0 1 243
box -10 0 100 799
use inv  g8607
timestamp 1395695751
transform 1 0 5904 0 1 243
box 0 0 120 799
use nand2  g8727
timestamp 1395695751
transform 1 0 6024 0 1 243
box -10 0 100 799
use nor2  g8471
timestamp 1395695751
transform 1 0 6120 0 1 243
box -3 0 125 799
use nand2  g8492
timestamp 1395695751
transform 1 0 6240 0 1 243
box -10 0 100 799
use nand2  g8583
timestamp 1395695751
transform 1 0 6336 0 1 243
box -10 0 100 799
use nand2  g8665
timestamp 1395695751
transform 1 0 6432 0 1 243
box -10 0 100 799
use nor2  g8685
timestamp 1395695751
transform 1 0 6528 0 1 243
box -3 0 125 799
use and2  g8662
timestamp 1395695751
transform 1 0 6648 0 1 243
box -10 0 127 799
use inv  g8621
timestamp 1395695751
transform 1 0 6768 0 1 243
box 0 0 120 799
use nor2  g8628
timestamp 1395695751
transform 1 0 6888 0 1 243
box -3 0 125 799
use and2  g8681
timestamp 1395695751
transform 1 0 7008 0 1 243
box -10 0 127 799
use nand3  g8657
timestamp 1395695751
transform 1 0 7128 0 1 243
box -10 0 127 799
use nand2  g8672
timestamp 1395695751
transform 1 0 7248 0 1 243
box -10 0 100 799
use nand2  g8482
timestamp 1395695751
transform 1 0 7344 0 1 243
box -10 0 100 799
use nand2  g8711
timestamp 1395695751
transform 1 0 7440 0 1 243
box -10 0 100 799
use nand3  g8467
timestamp 1395695751
transform 1 0 7536 0 1 243
box -10 0 127 799
use inv  g8722
timestamp 1395695751
transform 1 0 7656 0 1 243
box 0 0 120 799
use nor2  g8730
timestamp 1395695751
transform 1 0 7776 0 1 243
box -3 0 125 799
use nor2  g8647
timestamp 1395695751
transform 1 0 7896 0 1 243
box -3 0 125 799
use and2  g8539
timestamp 1395695751
transform 1 0 8016 0 1 243
box -10 0 127 799
use nor2  g8565
timestamp 1395695751
transform 1 0 8136 0 1 243
box -3 0 125 799
use and2  g8551
timestamp 1395695751
transform 1 0 8256 0 1 243
box -10 0 127 799
use nand2  g8704
timestamp 1395695751
transform 1 0 8376 0 1 243
box -10 0 100 799
use nand2  g8613
timestamp 1395695751
transform 1 0 8472 0 1 243
box -10 0 100 799
use inv  g8485
timestamp 1395695751
transform 1 0 8568 0 1 243
box 0 0 120 799
use nand4  g8497
timestamp 1395695751
transform 1 0 8688 0 1 243
box -10 0 154 799
use inv  g8751
timestamp 1395695751
transform 1 0 8832 0 1 243
box 0 0 120 799
use nand2  g8544
timestamp 1395695751
transform 1 0 8952 0 1 243
box -10 0 100 799
use nand3  g8569
timestamp 1395695751
transform 1 0 9048 0 1 243
box -10 0 127 799
use nand2  state_reg_91_0_93_
timestamp 1395695751
transform 1 0 9168 0 1 243
box -10 0 100 799
use scandtype  g8441
timestamp 1395695751
transform 1 0 9264 0 1 243
box -9 0 624 799
use rowcrosser  AluOR_91_0_93_
timestamp 1395695751
transform 1 0 9888 0 1 243
box 0 0 48 799
use nand3  g8654
timestamp 1395695751
transform 1 0 9936 0 1 243
box -10 0 127 799
use nand2  stateSub_reg_91_1_93_
timestamp 1395695751
transform 1 0 10056 0 1 243
box -10 0 100 799
use scandtype  g8652
timestamp 1395695751
transform 1 0 10152 0 1 243
box -9 0 624 799
use nand2  g8693
timestamp 1395695751
transform 1 0 10776 0 1 243
box -10 0 100 799
use nand2  g8767
timestamp 1395695751
transform 1 0 10872 0 1 243
box -10 0 100 799
use inv  g8525
timestamp 1395695751
transform 1 0 10968 0 1 243
box 0 0 120 799
use nand2  g8561
timestamp 1395695751
transform 1 0 11088 0 1 243
box -10 0 100 799
use nand2  g8528
timestamp 1395695751
transform 1 0 11184 0 1 243
box -10 0 100 799
use nand2  g8689
timestamp 1395695751
transform 1 0 11280 0 1 243
box -10 0 100 799
use and2  g8448
timestamp 1395695751
transform 1 0 11376 0 1 243
box -10 0 127 799
use nand2  g8739
timestamp 1395695751
transform 1 0 11496 0 1 243
box -10 0 100 799
use nor2  g8671
timestamp 1395695751
transform 1 0 11592 0 1 243
box -3 0 125 799
use nand2  g8606
timestamp 1395695751
transform 1 0 11712 0 1 243
box -10 0 100 799
use nand2  g8581
timestamp 1395695751
transform 1 0 11808 0 1 243
box -10 0 100 799
use nand3  g8576
timestamp 1395695751
transform 1 0 11904 0 1 243
box -10 0 127 799
use nand2  g8709
timestamp 1395695751
transform 1 0 12024 0 1 243
box -10 0 100 799
use nand2  g8734
timestamp 1395695751
transform 1 0 12120 0 1 243
box -10 0 100 799
use inv  SysBus_91_1_93_
timestamp 1395695751
transform 1 0 12216 0 1 243
box 0 0 120 799
use rowcrosser  SysBus_91_2_93_
timestamp 1395695751
transform 1 0 12336 0 1 243
box 0 0 48 799
use rowcrosser  nWE
timestamp 1395695751
transform 1 0 12384 0 1 243
box 0 0 48 799
<< labels >>
rlabel m2contact 12462 -230 12462 -230 8 AluOR[0]
rlabel m2contact 12462 -734 12462 -734 8 AluOR[0]
rlabel m2contact 12438 -278 12438 -278 8 AluOR[1]
rlabel m2contact 12438 -758 12438 -758 8 AluOR[1]
rlabel m2contact 12414 -374 12414 -374 8 ENB
rlabel m2contact 12414 -782 12414 -782 8 ENB
rlabel m2contact 12414 -230 12414 -230 8 AluOR[0]
rlabel m2contact 12366 -278 12366 -278 8 AluOR[1]
rlabel m2contact 11694 -446 11694 -446 8 n_11
rlabel m2contact 11574 202 11574 202 6 n_353
rlabel m2contact 11550 82 11550 82 6 SysBus[0]
rlabel m2contact 11238 -398 11238 -398 8 n_232
rlabel m2contact 11166 -422 11166 -422 8 n_129
rlabel m2contact 10950 -62 10950 -62 8 n_61
rlabel m2contact 10806 -638 10806 -638 8 n_106
rlabel m2contact 10614 -158 10614 -158 8 n_486
rlabel m2contact 10254 -206 10254 -206 8 n_337
rlabel m2contact 10110 -110 10110 -110 8 n_37
rlabel m2contact 9990 -278 9990 -278 8 n_316
rlabel m2contact 9966 -134 9966 -134 8 n_258
rlabel metal2 9936 -230 9936 -230 8 SysBus[3]
rlabel m2contact 9918 -230 9918 -230 8 SysBus[3]
rlabel m2contact 9198 -590 9198 -590 8 n_230
rlabel m2contact 9150 -230 9150 -230 8 n_181
rlabel m2contact 9078 -302 9078 -302 8 n_63
rlabel m2contact 8910 -686 8910 -686 8 n_291
rlabel m2contact 8862 -182 8862 -182 8 n_279
rlabel m2contact 8814 -134 8814 -134 8 n_258
rlabel m2contact 8742 -398 8742 -398 8 n_232
rlabel m2contact 8646 -398 8646 -398 8 n_232
rlabel m2contact 8550 -134 8550 -134 8 n_24
rlabel m2contact 8430 -326 8430 -326 8 n_123
rlabel m2contact 8190 -494 8190 -494 8 n_228
rlabel m2contact 8070 10 8070 10 6 n_16
rlabel m2contact 7998 -38 7998 -38 8 n_7
rlabel m2contact 7878 154 7878 154 6 n_46
rlabel m2contact 7734 -86 7734 -86 8 n_320
rlabel m2contact 7638 -710 7638 -710 8 n_18
rlabel m2contact 7518 -734 7518 -734 8 n_330
rlabel m2contact 7422 -350 7422 -350 8 n_21
rlabel m2contact 7230 178 7230 178 6 n_64
rlabel m2contact 7206 -302 7206 -302 8 n_63
rlabel m2contact 6582 -38 6582 -38 8 n_7
rlabel m2contact 6414 -38 6414 -38 8 n_309
rlabel m2contact 6390 -638 6390 -638 8 n_106
rlabel m2contact 5766 -614 5766 -614 8 n_306
rlabel m2contact 5430 -206 5430 -206 8 n_337
rlabel m2contact 5382 -206 5382 -206 8 n_287
rlabel m2contact 5334 -62 5334 -62 8 n_61
rlabel m2contact 4974 -518 4974 -518 8 IRQ1
rlabel m2contact 4566 -758 4566 -758 8 n_4
rlabel m2contact 3990 130 3990 130 6 n_132
rlabel m2contact 3822 -302 3822 -302 8 n_63
rlabel m2contact 3774 -110 3774 -110 8 n_37
rlabel m2contact 3678 106 3678 106 6 n_297
rlabel m2contact 3582 -110 3582 -110 8 n_259
rlabel m2contact 3486 -14 3486 -14 8 n_154
rlabel m2contact 3390 -278 3390 -278 8 n_316
rlabel m2contact 3342 -470 3342 -470 8 n_270
rlabel m2contact 3294 -278 3294 -278 8 n_225
rlabel m2contact 3150 34 3150 34 6 n_118
rlabel m2contact 3054 226 3054 226 6 n_71
rlabel m2contact 3030 154 3030 154 6 n_46
rlabel m2contact 3006 58 3006 58 6 n_56
rlabel m2contact 2934 -62 2934 -62 8 n_245
rlabel m2contact 2862 178 2862 178 6 n_64
rlabel m2contact 2790 10 2790 10 6 n_16
rlabel m2contact 2766 -158 2766 -158 8 n_486
rlabel m2contact 2694 -254 2694 -254 8 RegWe
rlabel m2contact 2622 -158 2622 -158 8 n_278
rlabel m2contact 2406 178 2406 178 6 n_29
rlabel m2contact 2334 -254 2334 -254 8 n_157
rlabel m2contact 2190 154 2190 154 6 n_46
rlabel m2contact 2142 -494 2142 -494 8 n_228
rlabel m2contact 1950 10 1950 10 6 IRQ2
rlabel m2contact 1542 -518 1542 -518 8 IRQ1
rlabel m2contact 1398 -494 1398 -494 8 n_228
rlabel m2contact 1014 -62 1014 -62 8 n_245
rlabel m2contact 966 -542 966 -542 8 n_265
rlabel m2contact 918 -62 918 -62 8 n_187
rlabel m2contact 894 -662 894 -662 8 n_102
rlabel m2contact 822 202 822 202 6 n_353
rlabel m2contact 774 106 774 106 6 n_297
rlabel m2contact 606 -62 606 -62 8 n_187
rlabel m2contact 582 10 582 10 6 IRQ2
rlabel m2contact 558 -62 558 -62 8 n_128
rlabel m2contact 510 10 510 10 6 IntStatus
rlabel m2contact 414 -590 414 -590 8 n_230
rlabel m2contact 342 -14 342 -14 8 n_154
rlabel m2contact 342 -494 342 -494 8 SysBus[2]
rlabel m2contact 318 -230 318 -230 8 n_181
rlabel m2contact 294 -566 294 -566 8 n_240
rlabel m2contact 270 -782 270 -782 8 n_236
rlabel m2contact 126 -230 126 -230 8 n_112
rlabel m2contact -18 202 -18 202 4 n_328
rlabel m2contact -42 -518 -42 -518 2 n_295
rlabel m2contact -258 -86 -258 -86 2 n_320
rlabel m2contact -282 -14 -282 -14 2 n_365
rlabel m2contact -378 -86 -378 -86 2 n_125
rlabel m2contact -402 106 -402 106 4 n_67
rlabel m2contact -426 226 -426 226 4 n_71
rlabel m2contact -810 202 -810 202 4 n_328
rlabel m2contact -954 58 -954 58 4 n_56
rlabel m2contact -1026 178 -1026 178 4 n_29
rlabel m2contact -1074 154 -1074 154 4 n_46
rlabel m2contact -1170 -422 -1170 -422 2 n_129
rlabel m2contact -1458 10 -1458 10 4 IntStatus
rlabel m2contact -2202 -422 -2202 -422 2 n_138
rlabel m2contact -2346 -62 -2346 -62 2 n_128
rlabel m2contact -2562 -638 -2562 -638 2 n_106
rlabel m2contact -2778 -206 -2778 -206 2 n_287
rlabel m2contact -2874 -206 -2874 -206 2 n_179
rlabel m2contact -3138 -590 -3138 -590 2 n_230
rlabel m2contact -3354 -14 -3354 -14 2 n_365
rlabel m2contact -3474 -86 -3474 -86 2 n_125
rlabel m2contact -3522 -62 -3522 -62 2 n_36
rlabel m2contact -3594 10 -3594 10 4 n_192
rlabel m2contact -3714 -86 -3714 -86 2 n_173
rlabel m2contact -3786 130 -3786 130 4 n_132
rlabel m2contact -3834 -662 -3834 -662 2 n_102
rlabel m2contact -3978 -614 -3978 -614 2 n_306
rlabel m2contact -4002 10 -4002 10 4 n_192
rlabel m2contact -4026 -38 -4026 -38 2 n_309
rlabel m2contact -4290 10 -4290 10 4 n_87
rlabel m2contact -4314 -422 -4314 -422 2 n_138
rlabel m2contact -4338 -38 -4338 -38 2 n_218
rlabel m2contact -4362 -86 -4362 -86 2 n_173
rlabel m2contact -4434 -662 -4434 -662 2 n_82
rlabel m2contact -4482 -614 -4482 -614 2 n_107
rlabel m2contact -4554 -86 -4554 -86 2 n_300
rlabel m2contact -4698 -470 -4698 -470 2 n_270
rlabel m2contact -4722 -422 -4722 -422 2 n_204
rlabel m2contact -4914 -470 -4914 -470 2 n_161
rlabel m2contact -5058 -734 -5058 -734 2 n_330
rlabel m2contact -5178 -14 -5178 -14 2 n_365
rlabel m2contact -5418 -782 -5418 -782 2 n_236
rlabel m2contact -5634 106 -5634 106 4 n_67
rlabel m2contact -5862 -782 -5862 -782 2 SysBus[1]
rlabel m2contact -5874 106 -5874 106 4 n_63
rlabel m2contact -5874 -302 -5874 -302 2 n_63
rlabel m2contact -5898 106 -5898 106 4 n_63
rlabel m2contact -5898 82 -5898 82 4 SysBus[0]
rlabel m2contact -6186 58 -6186 58 4 n_56
rlabel m2contact -6330 34 -6330 34 4 n_118
rlabel m2contact -6378 10 -6378 10 4 n_87
rlabel m2contact -6546 -14 -6546 -14 2 n_365
rlabel m2contact -6618 -782 -6618 -782 2 SysBus[1]
rlabel m2contact -6666 -38 -6666 -38 2 n_218
rlabel m2contact -6786 -62 -6786 -62 2 n_36
rlabel m2contact -6882 -374 -6882 -374 2 ENB
rlabel m2contact -6930 -374 -6930 -374 2 n_219
rlabel m2contact -6954 -86 -6954 -86 2 n_300
rlabel m2contact -7050 -110 -7050 -110 2 n_259
rlabel m2contact -7074 -734 -7074 -734 2 n_330
rlabel m2contact -7122 -734 -7122 -734 2 n_144
rlabel m2contact -7146 -134 -7146 -134 2 n_24
rlabel m2contact -7170 -230 -7170 -230 2 n_112
rlabel m2contact -7218 -230 -7218 -230 2 n_166
rlabel m2contact -7410 -158 -7410 -158 2 n_278
rlabel m2contact -7530 -182 -7530 -182 2 n_279
rlabel m2contact -7554 -206 -7554 -206 2 n_179
rlabel m2contact -7602 -230 -7602 -230 2 n_166
rlabel m2contact -7674 -494 -7674 -494 2 SysBus[2]
rlabel m2contact -8682 -494 -8682 -494 2 n_274
rlabel m2contact -8706 -254 -8706 -254 2 n_157
rlabel m2contact -8730 -278 -8730 -278 2 n_225
rlabel m2contact -8778 -302 -8778 -302 2 n_63
rlabel m2contact -9018 -326 -9018 -326 2 n_123
rlabel m2contact -9042 -350 -9042 -350 2 n_21
rlabel m2contact -9114 -374 -9114 -374 2 n_219
rlabel m2contact -9138 -398 -9138 -398 2 n_232
rlabel m2contact -9210 -422 -9210 -422 2 n_204
rlabel m2contact -9234 -446 -9234 -446 2 n_11
rlabel m2contact -9306 -470 -9306 -470 2 n_161
rlabel m2contact -9498 -494 -9498 -494 2 n_274
rlabel m2contact -9546 -518 -9546 -518 2 n_295
rlabel m2contact -10146 -542 -10146 -542 2 n_265
rlabel m2contact -10266 -566 -10266 -566 2 n_240
rlabel m2contact -10314 -590 -10314 -590 2 n_230
rlabel m2contact -10362 -614 -10362 -614 2 n_107
rlabel m2contact -10410 -638 -10410 -638 2 n_106
rlabel m2contact -10554 -662 -10554 -662 2 n_82
rlabel m2contact -10698 -686 -10698 -686 2 n_291
rlabel m2contact -10794 -758 -10794 -758 2 n_4
rlabel m2contact -10842 -758 -10842 -758 2 nIRQ
rlabel m2contact -11178 -710 -11178 -710 2 n_18
rlabel m2contact -11730 -734 -11730 -734 2 n_144
rlabel m2contact -11970 -734 -11970 -734 2 nWE
rlabel m2contact 12822 7076 12822 7076 6 Flags[0]
rlabel m2contact 12822 6836 12822 6836 6 Flags[0]
rlabel m2contact 12798 6908 12798 6908 6 Flags[3]
rlabel m2contact 12798 6836 12798 6836 6 Flags[3]
rlabel m2contact 12774 6980 12774 6980 6 Flags[2]
rlabel m2contact 12774 6884 12774 6884 6 Flags[2]
rlabel m2contact 12750 7004 12750 7004 6 CFlag
rlabel m2contact 12750 6932 12750 6932 6 CFlag
rlabel m2contact 12750 6884 12750 6884 6 Flags[1]
rlabel m2contact 12750 6860 12750 6860 6 Flags[1]
rlabel m2contact 12726 6980 12726 6980 6 Flags[2]
rlabel m2contact 12054 6980 12054 6980 6 OpcodeCondIn[0]
rlabel m2contact 11886 6956 11886 6956 6 MemEn
rlabel m2contact 11754 6908 11754 6908 6 StatusRegEn
rlabel m2contact 11334 6860 11334 6860 6 PcSel[0]
rlabel m2contact 10938 6932 10938 6932 6 StatusReg[3]
rlabel m2contact 10278 6836 10278 6836 6 Flags[3]
rlabel m2contact 10122 7148 10122 7148 6 StatusReg[2]
rlabel m2contact 9438 7052 9438 7052 6 Op2Sel[0]
rlabel m2contact 9306 7124 9306 7124 6 StatusReg[1]
rlabel m2contact 8934 6908 8934 6908 6 StatusRegEn
rlabel m2contact 8742 6836 8742 6836 6 PcSel[1]
rlabel m2contact 8490 6908 8490 6908 6 StatusReg[0]
rlabel m2contact 8166 7100 8166 7100 6 AluWe
rlabel m2contact 8022 6908 8022 6908 6 StatusReg[0]
rlabel m2contact 7674 7028 7674 7028 6 AluEn
rlabel m2contact 7650 7100 7650 7100 6 AluWe
rlabel m2contact 7206 6908 7206 6908 6 IrWe
rlabel m2contact 6966 7100 6966 7100 6 Op2Sel[1]
rlabel m2contact 6870 6932 6870 6932 6 StatusReg[3]
rlabel m2contact 6834 7100 6834 7100 6 Op2Sel[1]
rlabel m2contact 6294 7076 6294 7076 6 Flags[0]
rlabel m2contact 6018 7052 6018 7052 6 Op2Sel[0]
rlabel m2contact 5598 6980 5598 6980 6 OpcodeCondIn[0]
rlabel m2contact 4410 7052 4410 7052 6 Op1Sel
rlabel metal2 4320 7076 4320 7076 6 PcEn
rlabel m2contact 4302 7076 4302 7076 6 PcEn
rlabel m2contact 3702 7076 3702 7076 6 WdSel
rlabel m2contact 3570 7076 3570 7076 6 WdSel
rlabel m2contact 3558 7004 3558 7004 6 CFlag
rlabel m2contact 1962 7100 1962 7100 6 PcWe
rlabel m2contact 1950 7004 1950 7004 6 nME
rlabel m2contact 1146 7076 1146 7076 6 PcSel[2]
rlabel m2contact 1122 6836 1122 6836 6 PcSel[1]
rlabel m2contact 462 6932 462 6932 6 StatusReg[3]
rlabel m2contact 306 6860 306 6860 6 PcSel[0]
rlabel m2contact -426 7148 -426 7148 4 StatusReg[2]
rlabel m2contact -594 6884 -594 6884 4 Flags[1]
rlabel m2contact -810 7076 -810 7076 4 PcSel[2]
rlabel m2contact -906 6980 -906 6980 4 OpcodeCondIn[0]
rlabel m2contact -1314 7076 -1314 7076 4 LrEn
rlabel m2contact -1506 7124 -1506 7124 4 StatusReg[1]
rlabel m2contact -1650 7052 -1650 7052 4 Op1Sel
rlabel m2contact -2142 7052 -2142 7052 4 LrWe
rlabel metal2 -2352 7124 -2352 7124 4 LrSel
rlabel m2contact -2370 7124 -2370 7124 4 LrSel
rlabel metal2 -3240 7124 -3240 7124 4 ImmSel
rlabel m2contact -3258 7124 -3258 7124 4 ImmSel
rlabel m2contact -3834 6908 -3834 6908 4 IrWe
rlabel m2contact -4602 7100 -4602 7100 4 PcWe
rlabel m2contact -4662 6956 -4662 6956 4 MemEn
rlabel m2contact -4722 6956 -4722 6956 4 OpcodeCondIn[5]
rlabel m2contact -4794 7076 -4794 7076 4 LrEn
rlabel m2contact -5058 7028 -5058 7028 4 AluEn
rlabel m2contact -6282 7076 -6282 7076 4 OpcodeCondIn[7]
rlabel m2contact -6354 7028 -6354 7028 4 ALE
rlabel m2contact -6546 6932 -6546 6932 4 StatusReg[3]
rlabel m2contact -7050 7052 -7050 7052 4 LrWe
rlabel m2contact -7110 7052 -7110 7052 4 OpcodeCondIn[6]
rlabel m2contact -7146 6956 -7146 6956 4 OpcodeCondIn[5]
rlabel m2contact -7338 6956 -7338 6956 4 OpcodeCondIn[4]
rlabel m2contact -7974 6956 -7974 6956 4 OpcodeCondIn[4]
rlabel m2contact -8442 7076 -8442 7076 4 OpcodeCondIn[7]
rlabel m2contact -8586 7052 -8586 7052 4 OpcodeCondIn[6]
rlabel m2contact -9258 6980 -9258 6980 4 OpcodeCondIn[0]
rlabel m2contact -9594 7052 -9594 7052 4 OpcodeCondIn[3]
rlabel metal2 -10392 7076 -10392 7076 4 OpcodeCondIn[2]
rlabel m2contact -10410 7076 -10410 7076 4 OpcodeCondIn[2]
rlabel m2contact -10434 7052 -10434 7052 4 OpcodeCondIn[3]
rlabel metal2 -10800 7052 -10800 7052 4 OpcodeCondIn[1]
rlabel m2contact -10818 7052 -10818 7052 4 OpcodeCondIn[1]
rlabel m2contact -11352 6980 -11352 6980 4 OpcodeCondIn[0]
rlabel m2contact -11370 6980 -11370 6980 4 OpcodeCondIn[0]
rlabel m2contact 12774 5163 12774 5163 6 RwSel[0]
rlabel m2contact 12774 1083 12774 1083 6 RwSel[0]
rlabel m2contact 12750 3651 12750 3651 6 RwSel[1]
rlabel m2contact 12750 1059 12750 1059 6 RwSel[1]
rlabel m2contact 12726 1371 12726 1371 6 Flags[2]
rlabel m2contact 12702 4779 12702 4779 6 n_109
rlabel m2contact 12702 1539 12702 1539 6 n_109
rlabel m2contact 12678 3531 12678 3531 6 AluOR[0]
rlabel m2contact 12654 3771 12654 3771 6 n_310
rlabel m2contact 12630 3747 12630 3747 6 n_282
rlabel m2contact 12606 4587 12606 4587 6 n_266
rlabel m2contact 12606 3507 12606 3507 6 n_266
rlabel m2contact 12582 3819 12582 3819 6 n_349
rlabel m2contact 12558 3483 12558 3483 6 SysBus[3]
rlabel m2contact 12534 4491 12534 4491 6 n_351
rlabel m2contact 12498 3627 12498 3627 6 n_25
rlabel m2contact 12498 1731 12498 1731 6 n_25
rlabel m2contact 12486 4971 12486 4971 6 n_253
rlabel m2contact 12462 5595 12462 5595 6 n_163
rlabel m2contact 12438 4659 12438 4659 6 n_188
rlabel m2contact 12414 3531 12414 3531 6 AluOR[0]
rlabel m2contact 12390 4875 12390 4875 6 n_182
rlabel m2contact 12366 3795 12366 3795 6 AluOR[1]
rlabel m2contact 12342 3387 12342 3387 6 n_111
rlabel m2contact 12318 3915 12318 3915 6 n_190
rlabel m2contact 12294 1851 12294 1851 6 n_77
rlabel m2contact 12270 5907 12270 5907 6 n_20
rlabel m2contact 12270 2715 12270 2715 6 n_20
rlabel m2contact 12246 5019 12246 5019 6 n_32
rlabel m2contact 12246 4803 12246 4803 6 n_28
rlabel m2contact 12222 2739 12222 2739 6 stateSub[0]
rlabel m2contact 12198 4347 12198 4347 6 n_79
rlabel m2contact 12174 2523 12174 2523 6 n_81
rlabel m2contact 12174 2931 12174 2931 6 stateSub[1]
rlabel m2contact 12150 3435 12150 3435 6 n_215
rlabel m2contact 12150 4059 12150 4059 6 n_276
rlabel m2contact 12126 5043 12126 5043 6 n_332
rlabel m2contact 12126 3459 12126 3459 6 n_332
rlabel m2contact 12102 4395 12102 4395 6 n_198
rlabel m2contact 12078 4131 12078 4131 6 n_8
rlabel m2contact 12078 3843 12078 3843 6 n_248
rlabel m2contact 12054 4851 12054 4851 6 n_221
rlabel m2contact 12030 3603 12030 3603 6 OpcodeCondIn[1]
rlabel m2contact 12006 5547 12006 5547 6 n_126
rlabel m2contact 11982 1539 11982 1539 6 n_109
rlabel m2contact 11982 1563 11982 1563 6 n_113
rlabel m2contact 11958 5259 11958 5259 6 state[0]
rlabel m2contact 11958 2043 11958 2043 6 n_39
rlabel m2contact 11934 3051 11934 3051 6 n_74
rlabel m2contact 11934 2931 11934 2931 6 stateSub[1]
rlabel m2contact 11910 5451 11910 5451 6 n_91
rlabel m2contact 11910 1155 11910 1155 6 n_91
rlabel m2contact 11886 5715 11886 5715 6 n_374
rlabel m2contact 11862 4587 11862 4587 6 n_266
rlabel m2contact 11862 4563 11862 4563 6 n_85
rlabel m2contact 11838 4035 11838 4035 6 n_318
rlabel m2contact 11838 3531 11838 3531 6 n_185
rlabel m2contact 11814 5427 11814 5427 6 n_224
rlabel m2contact 11814 1587 11814 1587 6 n_224
rlabel m2contact 11790 1731 11790 1731 6 n_25
rlabel m2contact 11790 1755 11790 1755 6 n_89
rlabel m2contact 11766 2715 11766 2715 6 n_20
rlabel m2contact 11766 2739 11766 2739 6 stateSub[0]
rlabel m2contact 11742 4899 11742 4899 6 n_66
rlabel m2contact 11742 2979 11742 2979 6 n_30
rlabel m2contact 11718 2523 11718 2523 6 n_81
rlabel m2contact 11694 5955 11694 5955 6 n_250
rlabel m2contact 11694 3411 11694 3411 6 n_250
rlabel m2contact 11682 3147 11682 3147 6 n_122
rlabel m2contact 11682 2907 11682 2907 6 n_122
rlabel m2contact 11670 4899 11670 4899 6 n_66
rlabel m2contact 11646 2811 11646 2811 6 OpcodeCondIn[7]
rlabel m2contact 11622 2907 11622 2907 6 n_122
rlabel m2contact 11622 2931 11622 2931 6 stateSub[1]
rlabel m2contact 11598 3843 11598 3843 6 n_248
rlabel m2contact 11562 3555 11562 3555 6 n_340
rlabel m2contact 11562 1779 11562 1779 6 n_340
rlabel m2contact 11550 4491 11550 4491 6 n_351
rlabel m2contact 11526 4491 11526 4491 6 n_351
rlabel m2contact 11502 3891 11502 3891 6 OpcodeCondIn[2]
rlabel m2contact 11478 5043 11478 5043 6 n_332
rlabel m2contact 11478 4995 11478 4995 6 n_252
rlabel m2contact 11454 4083 11454 4083 6 n_222
rlabel m2contact 11454 2619 11454 2619 6 n_222
rlabel m2contact 11430 5451 11430 5451 6 n_91
rlabel m2contact 11430 5403 11430 5403 6 n_264
rlabel m2contact 11406 3411 11406 3411 6 n_250
rlabel m2contact 11406 4203 11406 4203 6 n_178
rlabel m2contact 11382 1995 11382 1995 6 n_57
rlabel m2contact 11358 4419 11358 4419 6 n_244
rlabel m2contact 11334 5931 11334 5931 6 n_95
rlabel m2contact 11310 3555 11310 3555 6 n_340
rlabel m2contact 11310 2643 11310 2643 6 n_243
rlabel m2contact 11286 5379 11286 5379 6 n_312
rlabel m2contact 11262 3579 11262 3579 6 n_233
rlabel m2contact 11238 5499 11238 5499 6 n_162
rlabel m2contact 11214 1275 11214 1275 6 n_268
rlabel m2contact 11214 2019 11214 2019 6 OpcodeCondIn[4]
rlabel m2contact 11190 2715 11190 2715 6 n_239
rlabel m2contact 11166 3363 11166 3363 6 n_75
rlabel m2contact 11142 4299 11142 4299 6 OpcodeCondIn[6]
rlabel m2contact 11142 2811 11142 2811 6 OpcodeCondIn[7]
rlabel m2contact 11118 1803 11118 1803 6 n_114
rlabel m2contact 11094 4275 11094 4275 6 n_216
rlabel m2contact 11070 1635 11070 1635 6 n_214
rlabel m2contact 11046 3435 11046 3435 6 n_215
rlabel m2contact 11046 2835 11046 2835 6 n_237
rlabel m2contact 11022 4059 11022 4059 6 n_276
rlabel m2contact 10998 3099 10998 3099 6 OpcodeCondIn[3]
rlabel m2contact 10974 5979 10974 5979 6 n_285
rlabel m2contact 10950 2547 10950 2547 6 n_284
rlabel m2contact 10926 5427 10926 5427 6 n_224
rlabel m2contact 10926 5403 10926 5403 6 n_264
rlabel m2contact 10902 4083 10902 4083 6 n_222
rlabel m2contact 10902 4011 10902 4011 6 n_86
rlabel m2contact 10878 5571 10878 5571 6 n_206
rlabel m2contact 10854 5067 10854 5067 6 n_104
rlabel m2contact 10830 3555 10830 3555 6 n_196
rlabel m2contact 10830 2523 10830 2523 6 n_81
rlabel m2contact 10806 3315 10806 3315 6 n_195
rlabel m2contact 10782 3675 10782 3675 6 n_140
rlabel m2contact 10758 5499 10758 5499 6 n_162
rlabel m2contact 10710 3939 10710 3939 6 n_43
rlabel m2contact 10686 4323 10686 4323 6 n_42
rlabel m2contact 10662 4899 10662 4899 6 n_66
rlabel m2contact 10662 2931 10662 2931 6 stateSub[1]
rlabel m2contact 10614 3267 10614 3267 6 n_101
rlabel m2contact 10590 5739 10590 5739 6 stateSub[2]
rlabel m2contact 10566 2499 10566 2499 6 n_84
rlabel m2contact 10518 2691 10518 2691 6 n_169
rlabel m2contact 10494 2019 10494 2019 6 OpcodeCondIn[4]
rlabel m2contact 10470 3531 10470 3531 6 n_185
rlabel m2contact 10422 3195 10422 3195 6 n_302
rlabel m2contact 10398 3291 10398 3291 6 n_267
rlabel m2contact 10374 1275 10374 1275 6 n_268
rlabel m2contact 10350 3843 10350 3843 6 n_248
rlabel m2contact 10302 3723 10302 3723 6 n_323
rlabel m2contact 10254 1395 10254 1395 6 n_327
rlabel m2contact 10206 5835 10206 5835 6 n_60
rlabel m2contact 10182 4515 10182 4515 6 n_26
rlabel m2contact 10158 5859 10158 5859 6 n_12
rlabel m2contact 10134 4107 10134 4107 6 n_97
rlabel m2contact 10110 5739 10110 5739 6 stateSub[2]
rlabel m2contact 10110 3411 10110 3411 6 stateSub[2]
rlabel m2contact 10086 3411 10086 3411 6 stateSub[2]
rlabel m2contact 10086 4611 10086 4611 6 n_151
rlabel m2contact 10038 3315 10038 3315 6 n_195
rlabel m2contact 10038 1731 10038 1731 6 n_354
rlabel m2contact 10014 2259 10014 2259 6 n_155
rlabel m2contact 9990 3675 9990 3675 6 n_140
rlabel m2contact 9966 3411 9966 3411 6 n_211
rlabel m2contact 9942 5283 9942 5283 6 n_108
rlabel m2contact 9918 3483 9918 3483 6 SysBus[3]
rlabel m2contact 9894 5619 9894 5619 6 n_149
rlabel m2contact 9870 3099 9870 3099 6 OpcodeCondIn[3]
rlabel m2contact 9846 3003 9846 3003 6 n_136
rlabel m2contact 9822 1971 9822 1971 6 n_189
rlabel m2contact 9798 5307 9798 5307 6 n_165
rlabel m2contact 9798 2331 9798 2331 6 n_165
rlabel m2contact 9774 5307 9774 5307 6 n_165
rlabel m2contact 9774 5259 9774 5259 6 state[0]
rlabel m2contact 9750 2715 9750 2715 6 n_239
rlabel m2contact 9726 2427 9726 2427 6 n_53
rlabel m2contact 9726 2931 9726 2931 6 stateSub[1]
rlabel m2contact 9702 1179 9702 1179 6 n_137
rlabel m2contact 9654 3675 9654 3675 6 n_371
rlabel m2contact 9630 3819 9630 3819 6 n_349
rlabel m2contact 9606 3723 9606 3723 6 n_323
rlabel m2contact 9582 5211 9582 5211 6 n_292
rlabel m2contact 9534 4755 9534 4755 6 n_51
rlabel m2contact 9510 4299 9510 4299 6 OpcodeCondIn[6]
rlabel m2contact 9486 5475 9486 5475 6 n_50
rlabel m2contact 9462 5187 9462 5187 6 n_231
rlabel m2contact 9462 3339 9462 3339 6 n_231
rlabel m2contact 9438 4587 9438 4587 6 n_121
rlabel m2contact 9438 2595 9438 2595 6 n_121
rlabel m2contact 9414 3483 9414 3483 6 n_234
rlabel m2contact 9390 3723 9390 3723 6 n_193
rlabel m2contact 9366 5187 9366 5187 6 n_231
rlabel m2contact 9366 5139 9366 5139 6 n_308
rlabel m2contact 9342 4683 9342 4683 6 n_17
rlabel m2contact 9342 2667 9342 2667 6 n_17
rlabel m2contact 9318 4227 9318 4227 6 n_110
rlabel m2contact 9294 5259 9294 5259 6 state[0]
rlabel m2contact 9294 1659 9294 1659 6 state[0]
rlabel m2contact 9270 1491 9270 1491 6 n_31
rlabel m2contact 9246 3339 9246 3339 6 n_231
rlabel m2contact 9246 5355 9246 5355 6 n_69
rlabel m2contact 9222 1971 9222 1971 6 n_189
rlabel m2contact 9198 3723 9198 3723 6 n_193
rlabel m2contact 9174 3147 9174 3147 6 n_122
rlabel m2contact 9150 3915 9150 3915 6 n_190
rlabel m2contact 9126 2595 9126 2595 6 n_121
rlabel m2contact 9126 2715 9126 2715 6 n_239
rlabel m2contact 9102 3531 9102 3531 6 n_185
rlabel m2contact 9078 3699 9078 3699 6 Rs1Sel[1]
rlabel m2contact 9054 3771 9054 3771 6 n_310
rlabel m2contact 9030 2667 9030 2667 6 n_17
rlabel m2contact 9030 2763 9030 2763 6 n_321
rlabel m2contact 9006 1659 9006 1659 6 state[0]
rlabel m2contact 9006 1683 9006 1683 6 n_364
rlabel m2contact 8982 5643 8982 5643 6 n_269
rlabel m2contact 8982 3843 8982 3843 6 n_248
rlabel m2contact 8934 2475 8934 2475 6 StatusRegEn
rlabel m2contact 8886 2307 8886 2307 6 n_294
rlabel m2contact 8862 3315 8862 3315 6 n_195
rlabel m2contact 8838 1347 8838 1347 6 n_172
rlabel m2contact 8814 1275 8814 1275 6 n_268
rlabel m2contact 8790 6003 8790 6003 6 n_105
rlabel m2contact 8790 2907 8790 2907 6 nWait
rlabel m2contact 8766 2187 8766 2187 6 n_257
rlabel m2contact 8742 4827 8742 4827 6 n_340
rlabel m2contact 8742 1779 8742 1779 6 n_340
rlabel m2contact 8718 4827 8718 4827 6 n_340
rlabel m2contact 8718 4731 8718 4731 6 n_288
rlabel m2contact 8694 1299 8694 1299 6 n_345
rlabel m2contact 8670 1515 8670 1515 6 n_335
rlabel m2contact 8622 3651 8622 3651 6 RwSel[1]
rlabel m2contact 8598 2883 8598 2883 6 n_359
rlabel m2contact 8598 2451 8598 2451 6 n_199
rlabel m2contact 8574 1683 8574 1683 6 n_364
rlabel m2contact 8550 3219 8550 3219 6 n_203
rlabel m2contact 8526 5403 8526 5403 6 n_264
rlabel m2contact 8502 3435 8502 3435 6 n_215
rlabel m2contact 8478 5115 8478 5115 6 n_296
rlabel m2contact 8454 3483 8454 3483 6 n_234
rlabel m2contact 8430 4251 8430 4251 6 n_281
rlabel m2contact 8406 3651 8406 3651 6 n_235
rlabel m2contact 8382 4371 8382 4371 6 n_80
rlabel m2contact 8358 2475 8358 2475 6 StatusRegEn
rlabel m2contact 8358 2499 8358 2499 6 n_84
rlabel m2contact 8334 4443 8334 4443 6 n_88
rlabel m2contact 8310 4179 8310 4179 6 n_226
rlabel m2contact 8286 4923 8286 4923 6 n_76
rlabel m2contact 8286 2187 8286 2187 6 n_257
rlabel m2contact 8262 4299 8262 4299 6 OpcodeCondIn[6]
rlabel m2contact 8238 5475 8238 5475 6 n_50
rlabel m2contact 8238 4707 8238 4707 6 n_289
rlabel m2contact 8214 2019 8214 2019 6 OpcodeCondIn[4]
rlabel m2contact 8190 5739 8190 5739 6 stateSub[2]
rlabel m2contact 8190 3483 8190 3483 6 stateSub[2]
rlabel m2contact 8166 3483 8166 3483 6 stateSub[2]
rlabel m2contact 8166 5235 8166 5235 6 AluWe
rlabel m2contact 8118 5091 8118 5091 6 n_314
rlabel m2contact 8046 4995 8046 4995 6 n_252
rlabel m2contact 8022 3987 8022 3987 6 StatusReg[0]
rlabel m2contact 7974 1419 7974 1419 6 n_484
rlabel m2contact 7950 3891 7950 3891 6 OpcodeCondIn[2]
rlabel m2contact 7926 2811 7926 2811 6 OpcodeCondIn[7]
rlabel m2contact 7830 3603 7830 3603 6 OpcodeCondIn[1]
rlabel m2contact 7806 3339 7806 3339 6 n_13
rlabel m2contact 7686 4539 7686 4539 6 n_305
rlabel m2contact 7638 4467 7638 4467 6 n_373
rlabel m2contact 7638 1227 7638 1227 6 n_373
rlabel m2contact 7614 4467 7614 4467 6 n_373
rlabel m2contact 7614 4299 7614 4299 6 OpcodeCondIn[6]
rlabel m2contact 7590 2739 7590 2739 6 stateSub[0]
rlabel m2contact 7566 3099 7566 3099 6 OpcodeCondIn[3]
rlabel m2contact 7542 3723 7542 3723 6 n_122
rlabel m2contact 7542 3147 7542 3147 6 n_122
rlabel m2contact 7518 5307 7518 5307 6 n_99
rlabel m2contact 7518 1131 7518 1131 6 n_99
rlabel m2contact 7494 5955 7494 5955 6 n_250
rlabel m2contact 7494 4155 7494 4155 6 n_209
rlabel m2contact 7470 4059 7470 4059 6 n_276
rlabel m2contact 7470 3243 7470 3243 6 n_313
rlabel m2contact 7446 2427 7446 2427 6 n_53
rlabel m2contact 7422 3699 7422 3699 6 n_189
rlabel m2contact 7422 1971 7422 1971 6 n_189
rlabel m2contact 7398 6003 7398 6003 6 n_105
rlabel m2contact 7398 5907 7398 5907 6 n_20
rlabel m2contact 7374 5307 7374 5307 6 n_99
rlabel m2contact 7374 4587 7374 4587 6 n_121
rlabel m2contact 7350 3843 7350 3843 6 n_248
rlabel m2contact 7326 4827 7326 4827 6 n_130
rlabel m2contact 7302 3363 7302 3363 6 n_75
rlabel m2contact 7302 4947 7302 4947 6 n_78
rlabel m2contact 7278 3723 7278 3723 6 n_122
rlabel m2contact 7278 3411 7278 3411 6 n_211
rlabel m2contact 7254 1851 7254 1851 6 n_77
rlabel m2contact 7230 4587 7230 4587 6 n_121
rlabel m2contact 7230 2859 7230 2859 6 n_121
rlabel m2contact 7206 3171 7206 3171 6 IrWe
rlabel m2contact 7182 3843 7182 3843 6 n_248
rlabel m2contact 7158 5307 7158 5307 6 n_99
rlabel m2contact 7158 5259 7158 5259 6 state[0]
rlabel m2contact 7134 4299 7134 4299 6 OpcodeCondIn[6]
rlabel m2contact 7110 3699 7110 3699 6 n_189
rlabel m2contact 7110 2211 7110 2211 6 n_160
rlabel m2contact 7086 4467 7086 4467 6 n_55
rlabel m2contact 7086 3483 7086 3483 6 n_55
rlabel m2contact 7062 2859 7062 2859 6 n_121
rlabel m2contact 7062 2955 7062 2955 6 n_200
rlabel m2contact 7038 4827 7038 4827 6 n_130
rlabel m2contact 7038 3411 7038 3411 6 n_211
rlabel m2contact 7014 2451 7014 2451 6 n_199
rlabel m2contact 6990 4779 6990 4779 6 n_109
rlabel m2contact 6966 3699 6966 3699 6 Op2Sel[1]
rlabel m2contact 6942 4203 6942 4203 6 n_178
rlabel m2contact 6918 4467 6918 4467 6 n_55
rlabel m2contact 6918 4155 6918 4155 6 n_209
rlabel m2contact 6894 1947 6894 1947 6 n_485
rlabel m2contact 6846 3171 6846 3171 6 IrWe
rlabel m2contact 6822 4467 6822 4467 6 n_156
rlabel m2contact 6798 5691 6798 5691 6 OpcodeCondIn[5]
rlabel m2contact 6798 1755 6798 1755 6 n_89
rlabel m2contact 6774 3531 6774 3531 6 n_185
rlabel m2contact 6750 5307 6750 5307 6 n_72
rlabel m2contact 6726 1251 6726 1251 6 n_103
rlabel m2contact 6702 5739 6702 5739 6 stateSub[2]
rlabel m2contact 6702 3843 6702 3843 6 n_248
rlabel m2contact 6678 5451 6678 5451 6 n_83
rlabel m2contact 6678 5403 6678 5403 6 n_264
rlabel m2contact 6630 5043 6630 5043 6 n_48
rlabel m2contact 6630 2379 6630 2379 6 n_23
rlabel m2contact 6606 4635 6606 4635 6 n_22
rlabel m2contact 6606 2667 6606 2667 6 n_22
rlabel m2contact 6582 2811 6582 2811 6 OpcodeCondIn[7]
rlabel m2contact 6558 2667 6558 2667 6 n_22
rlabel m2contact 6558 2715 6558 2715 6 n_239
rlabel m2contact 6534 5427 6534 5427 6 n_273
rlabel m2contact 6534 3171 6534 3171 6 n_273
rlabel m2contact 6510 3387 6510 3387 6 n_111
rlabel m2contact 6510 3819 6510 3819 6 n_207
rlabel m2contact 6486 4083 6486 4083 6 n_171
rlabel m2contact 6486 2715 6486 2715 6 n_239
rlabel m2contact 6462 5187 6462 5187 6 n_70
rlabel m2contact 6462 5955 6462 5955 6 n_250
rlabel m2contact 6426 3459 6426 3459 6 n_332
rlabel m2contact 6426 1323 6426 1323 6 n_332
rlabel m2contact 6414 3723 6414 3723 6 n_98
rlabel m2contact 6390 4587 6390 4587 6 n_121
rlabel m2contact 6366 3171 6366 3171 6 n_273
rlabel m2contact 6366 3387 6366 3387 6 n_44
rlabel m2contact 6342 5667 6342 5667 6 n_345
rlabel m2contact 6342 1299 6342 1299 6 n_345
rlabel m2contact 6318 1515 6318 1515 6 n_335
rlabel m2contact 6318 1539 6318 1539 6 n_329
rlabel m2contact 6294 4731 6294 4731 6 n_288
rlabel m2contact 6270 1323 6270 1323 6 n_332
rlabel m2contact 6270 1395 6270 1395 6 n_327
rlabel m2contact 6246 3891 6246 3891 6 OpcodeCondIn[2]
rlabel m2contact 6246 3171 6246 3171 6 OpcodeCondIn[2]
rlabel m2contact 6222 5667 6222 5667 6 n_345
rlabel m2contact 6222 5331 6222 5331 6 n_6
rlabel m2contact 6198 1059 6198 1059 6 n_167
rlabel m2contact 6174 3171 6174 3171 6 OpcodeCondIn[2]
rlabel m2contact 6174 3243 6174 3243 6 n_313
rlabel m2contact 6150 4299 6150 4299 6 OpcodeCondIn[6]
rlabel m2contact 6126 4779 6126 4779 6 n_109
rlabel m2contact 6126 2667 6126 2667 6 n_109
rlabel m2contact 6102 3003 6102 3003 6 n_136
rlabel m2contact 6102 3651 6102 3651 6 n_235
rlabel m2contact 6078 2811 6078 2811 6 OpcodeCondIn[7]
rlabel m2contact 6054 2667 6054 2667 6 n_109
rlabel m2contact 6054 2691 6054 2691 6 n_169
rlabel m2contact 6030 3867 6030 3867 6 n_53
rlabel m2contact 6030 2427 6030 2427 6 n_53
rlabel m2contact 6006 2571 6006 2571 6 n_183
rlabel m2contact 5982 4611 5982 4611 6 n_151
rlabel m2contact 5982 2163 5982 2163 6 n_159
rlabel m2contact 5958 2859 5958 2859 6 n_205
rlabel m2contact 5934 2595 5934 2595 6 n_220
rlabel m2contact 5934 2739 5934 2739 6 stateSub[0]
rlabel m2contact 5910 4635 5910 4635 6 n_22
rlabel m2contact 5910 2403 5910 2403 6 n_22
rlabel m2contact 5886 3219 5886 3219 6 n_203
rlabel m2contact 5886 4155 5886 4155 6 n_209
rlabel m2contact 5862 2211 5862 2211 6 n_160
rlabel m2contact 5838 2139 5838 2139 6 n_210
rlabel m2contact 5838 3891 5838 3891 6 OpcodeCondIn[2]
rlabel m2contact 5814 4131 5814 4131 6 n_8
rlabel m2contact 5790 3963 5790 3963 6 n_251
rlabel m2contact 5790 1875 5790 1875 6 n_251
rlabel m2contact 5766 3075 5766 3075 6 n_194
rlabel m2contact 5742 2475 5742 2475 6 n_170
rlabel m2contact 5718 1395 5718 1395 6 n_327
rlabel m2contact 5718 2187 5718 2187 6 n_257
rlabel m2contact 5694 2739 5694 2739 6 stateSub[0]
rlabel m2contact 5658 3531 5658 3531 6 n_185
rlabel m2contact 5658 2787 5658 2787 6 n_185
rlabel m2contact 5646 4203 5646 4203 6 n_178
rlabel m2contact 5646 2715 5646 2715 6 n_239
rlabel m2contact 5622 5955 5622 5955 6 n_250
rlabel m2contact 5622 3027 5622 3027 6 n_250
rlabel m2contact 5598 5691 5598 5691 6 OpcodeCondIn[5]
rlabel m2contact 5574 3603 5574 3603 6 OpcodeCondIn[1]
rlabel m2contact 5550 2139 5550 2139 6 n_210
rlabel m2contact 5526 3171 5526 3171 6 n_15
rlabel m2contact 5502 3867 5502 3867 6 n_53
rlabel m2contact 5502 3099 5502 3099 6 OpcodeCondIn[3]
rlabel m2contact 5478 2787 5478 2787 6 n_185
rlabel m2contact 5478 2931 5478 2931 6 stateSub[1]
rlabel m2contact 5454 3867 5454 3867 6 n_267
rlabel m2contact 5454 3291 5454 3291 6 n_267
rlabel m2contact 5430 1899 5430 1899 6 n_202
rlabel m2contact 5406 2403 5406 2403 6 n_22
rlabel m2contact 5406 2475 5406 2475 6 n_170
rlabel m2contact 5382 2139 5382 2139 6 n_210
rlabel m2contact 5358 3123 5358 3123 6 n_34
rlabel m2contact 5334 1923 5334 1923 6 n_38
rlabel m2contact 5310 2835 5310 2835 6 n_237
rlabel m2contact 5286 1875 5286 1875 6 n_251
rlabel m2contact 5286 2043 5286 2043 6 n_39
rlabel m2contact 5262 5811 5262 5811 6 n_208
rlabel m2contact 5238 3027 5238 3027 6 n_250
rlabel m2contact 5238 3219 5238 3219 6 n_271
rlabel m2contact 5214 2787 5214 2787 6 n_115
rlabel m2contact 5190 2619 5190 2619 6 n_222
rlabel m2contact 5190 2643 5190 2643 6 n_243
rlabel m2contact 5166 2595 5166 2595 6 n_220
rlabel m2contact 5142 5643 5142 5643 6 n_269
rlabel m2contact 5142 4851 5142 4851 6 n_221
rlabel m2contact 5118 3867 5118 3867 6 n_267
rlabel m2contact 5118 3843 5118 3843 6 n_248
rlabel m2contact 5094 1275 5094 1275 6 n_268
rlabel m2contact 5046 3867 5046 3867 6 n_262
rlabel m2contact 5022 2835 5022 2835 6 n_237
rlabel m2contact 4998 3651 4998 3651 6 n_235
rlabel m2contact 4974 5043 4974 5043 6 n_48
rlabel m2contact 4902 4131 4902 4131 6 n_174
rlabel m2contact 4854 4827 4854 4827 6 n_130
rlabel m2contact 4806 4827 4806 4827 6 n_148
rlabel m2contact 4758 1467 4758 1467 6 n_52
rlabel m2contact 4734 5547 4734 5547 6 n_126
rlabel m2contact 4686 3771 4686 3771 6 n_310
rlabel m2contact 4662 4443 4662 4443 6 n_88
rlabel m2contact 4638 3435 4638 3435 6 n_215
rlabel m2contact 4590 1635 4590 1635 6 n_214
rlabel m2contact 4566 3315 4566 3315 6 n_195
rlabel m2contact 4542 1515 4542 1515 6 n_131
rlabel m2contact 4482 3291 4482 3291 6 n_267
rlabel m2contact 4482 1611 4482 1611 6 n_267
rlabel m2contact 4470 5475 4470 5475 6 n_50
rlabel m2contact 4446 3051 4446 3051 6 n_74
rlabel m2contact 4422 2715 4422 2715 6 n_239
rlabel m2contact 4398 5739 4398 5739 6 stateSub[2]
rlabel m2contact 4374 1323 4374 1323 6 n_33
rlabel m2contact 4374 3099 4374 3099 6 OpcodeCondIn[3]
rlabel m2contact 4350 5691 4350 5691 6 OpcodeCondIn[5]
rlabel m2contact 4326 2403 4326 2403 6 n_45
rlabel m2contact 4302 1203 4302 1203 6 PcEn
rlabel m2contact 4278 5739 4278 5739 6 stateSub[2]
rlabel m2contact 4254 5355 4254 5355 6 n_69
rlabel m2contact 4254 3027 4254 3027 6 n_58
rlabel m2contact 4230 4515 4230 4515 6 n_26
rlabel m2contact 4230 3051 4230 3051 6 n_26
rlabel m2contact 4206 3507 4206 3507 6 n_266
rlabel m2contact 4206 5259 4206 5259 6 state[0]
rlabel m2contact 4182 1611 4182 1611 6 n_267
rlabel m2contact 4182 1659 4182 1659 6 n_217
rlabel m2contact 4158 2187 4158 2187 6 n_257
rlabel m2contact 4134 5283 4134 5283 6 n_108
rlabel m2contact 4110 3051 4110 3051 6 n_26
rlabel m2contact 4110 3099 4110 3099 6 OpcodeCondIn[3]
rlabel m2contact 4086 4779 4086 4779 6 n_109
rlabel m2contact 4086 2811 4086 2811 6 OpcodeCondIn[7]
rlabel m2contact 4062 3147 4062 3147 6 n_122
rlabel m2contact 4038 4779 4038 4779 6 n_49
rlabel m2contact 4014 2835 4014 2835 6 n_237
rlabel m2contact 3990 5043 3990 5043 6 n_48
rlabel m2contact 3942 5043 3942 5043 6 n_247
rlabel m2contact 3942 1515 3942 1515 6 n_131
rlabel m2contact 3918 3555 3918 3555 6 n_196
rlabel m2contact 3894 4659 3894 4659 6 n_188
rlabel m2contact 3870 1971 3870 1971 6 n_189
rlabel m2contact 3846 1107 3846 1107 6 n_315
rlabel m2contact 3822 2979 3822 2979 6 n_30
rlabel m2contact 3798 1611 3798 1611 6 n_263
rlabel m2contact 3774 5091 3774 5091 6 n_314
rlabel m2contact 3750 4683 3750 4683 6 n_17
rlabel m2contact 3750 4299 3750 4299 6 OpcodeCondIn[6]
rlabel m2contact 3726 2067 3726 2067 6 n_14
rlabel m2contact 3702 3555 3702 3555 6 WdSel
rlabel m2contact 3654 3987 3654 3987 6 StatusReg[0]
rlabel m2contact 3630 2307 3630 2307 6 n_294
rlabel m2contact 3558 2163 3558 2163 6 n_159
rlabel m2contact 3558 2283 3558 2283 6 CFlag
rlabel m2contact 3534 2619 3534 2619 6 n_255
rlabel m2contact 3462 3507 3462 3507 6 n_153
rlabel m2contact 3438 3531 3438 3531 6 n_185
rlabel m2contact 3366 2715 3366 2715 6 n_239
rlabel m2contact 3270 3099 3270 3099 6 OpcodeCondIn[3]
rlabel m2contact 3246 4851 3246 4851 6 n_221
rlabel m2contact 3222 3843 3222 3843 6 n_248
rlabel m2contact 3198 4731 3198 4731 6 n_288
rlabel m2contact 3150 2235 3150 2235 6 n_372
rlabel m2contact 3126 2739 3126 2739 6 stateSub[0]
rlabel m2contact 3102 1875 3102 1875 6 n_100
rlabel m2contact 3030 2667 3030 2667 6 n_146
rlabel m2contact 3006 5691 3006 5691 6 OpcodeCondIn[5]
rlabel m2contact 2982 3483 2982 3483 6 n_55
rlabel m2contact 2982 4299 2982 4299 6 OpcodeCondIn[6]
rlabel m2contact 2958 5259 2958 5259 6 state[0]
rlabel m2contact 2958 3051 2958 3051 6 state[0]
rlabel m2contact 2934 4659 2934 4659 6 n_188
rlabel m2contact 2910 3171 2910 3171 6 n_15
rlabel m2contact 2886 2355 2886 2355 6 n_96
rlabel m2contact 2886 2427 2886 2427 6 n_53
rlabel m2contact 2862 3843 2862 3843 6 n_248
rlabel m2contact 2838 2331 2838 2331 6 n_165
rlabel m2contact 2814 3171 2814 3171 6 n_142
rlabel m2contact 2790 3099 2790 3099 6 OpcodeCondIn[3]
rlabel m2contact 2766 1659 2766 1659 6 n_217
rlabel m2contact 2742 3051 2742 3051 6 state[0]
rlabel m2contact 2742 4659 2742 4659 6 n_150
rlabel m2contact 2718 4611 2718 4611 6 n_151
rlabel m2contact 2694 5715 2694 5715 6 n_374
rlabel m2contact 2694 3051 2694 3051 6 n_374
rlabel m2contact 2670 3051 2670 3051 6 n_374
rlabel m2contact 2670 4683 2670 4683 6 n_147
rlabel m2contact 2646 1707 2646 1707 6 n_362
rlabel m2contact 2646 2667 2646 2667 6 n_146
rlabel m2contact 2622 3723 2622 3723 6 n_98
rlabel m2contact 2598 3627 2598 3627 6 n_25
rlabel m2contact 2598 2883 2598 2883 6 n_359
rlabel m2contact 2574 3723 2574 3723 6 n_286
rlabel m2contact 2574 2331 2574 2331 6 n_286
rlabel m2contact 2550 2091 2550 2091 6 n_184
rlabel m2contact 2526 3459 2526 3459 6 n_332
rlabel m2contact 2502 3099 2502 3099 6 OpcodeCondIn[3]
rlabel m2contact 2478 2331 2478 2331 6 n_286
rlabel m2contact 2478 2571 2478 2571 6 n_183
rlabel m2contact 2454 3627 2454 3627 6 n_35
rlabel m2contact 2454 3051 2454 3051 6 n_35
rlabel m2contact 2430 5907 2430 5907 6 n_20
rlabel m2contact 2430 5883 2430 5883 6 n_62
rlabel m2contact 2406 5283 2406 5283 6 n_167
rlabel m2contact 2406 1059 2406 1059 6 n_167
rlabel m2contact 2382 3051 2382 3051 6 n_35
rlabel m2contact 2382 3099 2382 3099 6 OpcodeCondIn[3]
rlabel m2contact 2358 5691 2358 5691 6 OpcodeCondIn[5]
rlabel m2contact 2334 5907 2334 5907 6 n_47
rlabel m2contact 2334 1083 2334 1083 6 n_47
rlabel m2contact 2310 5283 2310 5283 6 n_167
rlabel m2contact 2310 2211 2310 2211 6 n_160
rlabel m2contact 2286 2859 2286 2859 6 n_205
rlabel m2contact 2262 4731 2262 4731 6 n_288
rlabel m2contact 2238 1083 2238 1083 6 n_47
rlabel m2contact 2238 1443 2238 1443 6 n_65
rlabel m2contact 2214 4731 2214 4731 6 n_288
rlabel m2contact 2190 5187 2190 5187 6 n_70
rlabel m2contact 2166 2115 2166 2115 6 n_19
rlabel m2contact 2142 4155 2142 4155 6 n_209
rlabel m2contact 2118 4203 2118 4203 6 n_178
rlabel m2contact 2094 5139 2094 5139 6 n_308
rlabel m2contact 2094 4131 2094 4131 6 n_174
rlabel m2contact 2070 5403 2070 5403 6 n_264
rlabel m2contact 2046 5067 2046 5067 6 n_104
rlabel m2contact 2022 5043 2022 5043 6 n_247
rlabel m2contact 1998 3459 1998 3459 6 n_59
rlabel m2contact 1926 5019 1926 5019 6 n_32
rlabel m2contact 1902 4827 1902 4827 6 n_148
rlabel m2contact 1878 5763 1878 5763 6 n_120
rlabel m2contact 1854 5307 1854 5307 6 n_72
rlabel m2contact 1806 4539 1806 4539 6 n_305
rlabel m2contact 1782 3579 1782 3579 6 n_233
rlabel m2contact 1758 4419 1758 4419 6 n_244
rlabel m2contact 1734 3579 1734 3579 6 n_186
rlabel m2contact 1710 3867 1710 3867 6 n_262
rlabel m2contact 1662 3051 1662 3051 6 nWE
rlabel m2contact 1638 5787 1638 5787 6 n_54
rlabel m2contact 1614 3867 1614 3867 6 n_249
rlabel m2contact 1590 4275 1590 4275 6 n_216
rlabel m2contact 1566 5043 1566 5043 6 n_277
rlabel m2contact 1518 4251 1518 4251 6 n_281
rlabel m2contact 1494 5643 1494 5643 6 n_197
rlabel m2contact 1470 4227 1470 4227 6 n_110
rlabel m2contact 1446 5283 1446 5283 6 n_68
rlabel m2contact 1422 3291 1422 3291 6 n_267
rlabel m2contact 1422 4107 1422 4107 6 n_97
rlabel m2contact 1374 2451 1374 2451 6 n_199
rlabel m2contact 1374 3291 1374 3291 6 n_27
rlabel m2contact 1350 2427 1350 2427 6 n_53
rlabel m2contact 1326 1659 1326 1659 6 n_217
rlabel m2contact 1326 2331 1326 2331 6 state[1]
rlabel m2contact 1302 4107 1302 4107 6 n_180
rlabel m2contact 1302 1083 1302 1083 6 n_180
rlabel m2contact 1278 4107 1278 4107 6 n_180
rlabel m2contact 1278 2979 1278 2979 6 n_30
rlabel m2contact 1254 3939 1254 3939 6 n_43
rlabel m2contact 1254 3435 1254 3435 6 n_215
rlabel m2contact 1230 1827 1230 1827 6 n_135
rlabel m2contact 1206 4419 1206 4419 6 n_175
rlabel m2contact 1182 3939 1182 3939 6 n_191
rlabel m2contact 1158 3531 1158 3531 6 n_185
rlabel m2contact 1134 4131 1134 4131 6 n_174
rlabel m2contact 1086 5187 1086 5187 6 n_299
rlabel m2contact 1086 5739 1086 5739 6 stateSub[2]
rlabel m2contact 1038 1083 1038 1083 6 n_180
rlabel m2contact 1038 3843 1038 3843 6 n_248
rlabel m2contact 942 5403 942 5403 6 n_264
rlabel m2contact 846 1227 846 1227 6 n_373
rlabel m2contact 798 1539 798 1539 6 n_329
rlabel m2contact 726 2475 726 2475 6 n_170
rlabel m2contact 702 4107 702 4107 6 n_280
rlabel m2contact 702 1227 702 1227 6 n_280
rlabel m2contact 678 4107 678 4107 6 n_280
rlabel m2contact 678 3147 678 3147 6 n_122
rlabel m2contact 654 4611 654 4611 6 n_151
rlabel m2contact 534 2499 534 2499 6 n_84
rlabel m2contact 462 1587 462 1587 6 n_224
rlabel m2contact 438 1851 438 1851 6 n_77
rlabel m2contact 414 1587 414 1587 6 n_487
rlabel m2contact 366 1395 366 1395 6 n_327
rlabel m2contact 222 1851 222 1851 6 n_119
rlabel m2contact 198 5139 198 5139 6 n_127
rlabel m2contact 174 1923 174 1923 6 n_38
rlabel m2contact 102 2739 102 2739 6 stateSub[0]
rlabel m2contact 78 1539 78 1539 6 n_73
rlabel m2contact 54 3675 54 3675 6 n_371
rlabel m2contact 30 2235 30 2235 6 n_372
rlabel m2contact 6 5067 6 5067 6 n_352
rlabel m2contact -18 5019 -18 5019 4 ImmSel
rlabel m2contact -18 2235 -18 2235 4 ImmSel
rlabel m2contact -42 5547 -42 5547 4 n_133
rlabel m2contact -42 1083 -42 1083 4 n_133
rlabel m2contact -66 4107 -66 4107 4 n_117
rlabel m2contact -90 4227 -90 4227 4 n_168
rlabel m2contact -90 5739 -90 5739 4 stateSub[2]
rlabel m2contact -114 1275 -114 1275 4 n_268
rlabel m2contact -138 4131 -138 4131 4 n_174
rlabel m2contact -162 1059 -162 1059 4 n_167
rlabel m2contact -162 1275 -162 1275 4 n_268
rlabel m2contact -186 5355 -186 5355 4 n_164
rlabel m2contact -186 1923 -186 1923 4 n_164
rlabel m2contact -210 2235 -210 2235 4 ImmSel
rlabel m2contact -210 2499 -210 2499 4 n_84
rlabel m2contact -234 1083 -234 1083 4 n_133
rlabel m2contact -234 4659 -234 4659 4 n_150
rlabel m2contact -258 4275 -258 4275 4 n_9
rlabel m2contact -258 2235 -258 2235 4 n_9
rlabel m2contact -282 2547 -282 2547 4 n_284
rlabel m2contact -306 3843 -306 3843 4 n_248
rlabel m2contact -330 1923 -330 1923 4 n_164
rlabel m2contact -330 4443 -330 4443 4 n_88
rlabel m2contact -354 2235 -354 2235 4 n_9
rlabel m2contact -354 3027 -354 3027 4 n_58
rlabel m2contact -390 4587 -390 4587 4 n_121
rlabel m2contact -390 2235 -390 2235 4 n_121
rlabel m2contact -402 5475 -402 5475 4 n_293
rlabel m2contact -426 1923 -426 1923 4 StatusReg[2]
rlabel m2contact -450 2307 -450 2307 4 n_294
rlabel m2contact -474 3315 -474 3315 4 n_195
rlabel m2contact -498 1971 -498 1971 4 n_189
rlabel m2contact -498 4539 -498 4539 4 n_93
rlabel m2contact -522 2235 -522 2235 4 n_121
rlabel m2contact -522 2739 -522 2739 4 stateSub[0]
rlabel m2contact -546 2187 -546 2187 4 n_257
rlabel m2contact -570 2043 -570 2043 4 n_39
rlabel m2contact -594 1083 -594 1083 4 Flags[1]
rlabel m2contact -618 4587 -618 4587 4 n_121
rlabel m2contact -642 2427 -642 2427 4 n_53
rlabel m2contact -666 4251 -666 4251 4 n_261
rlabel m2contact -714 3363 -714 3363 4 n_75
rlabel m2contact -714 3675 -714 3675 4 n_260
rlabel m2contact -762 5667 -762 5667 4 n_368
rlabel m2contact -762 3363 -762 3363 4 n_134
rlabel m2contact -810 3315 -810 3315 4 PcSel[2]
rlabel m2contact -834 1083 -834 1083 4 Flags[1]
rlabel m2contact -834 2235 -834 2235 4 n_348
rlabel m2contact -858 1395 -858 1395 4 n_327
rlabel m2contact -882 4275 -882 4275 4 n_9
rlabel m2contact -906 1995 -906 1995 4 n_57
rlabel m2contact -930 3483 -930 3483 4 n_55
rlabel m2contact -930 3987 -930 3987 4 StatusReg[0]
rlabel m2contact -954 3603 -954 3603 4 OpcodeCondIn[1]
rlabel m2contact -1002 3987 -1002 3987 4 n_275
rlabel m2contact -1026 5955 -1026 5955 4 n_250
rlabel m2contact -1050 3483 -1050 3483 4 n_272
rlabel m2contact -1122 1347 -1122 1347 4 n_172
rlabel m2contact -1122 4731 -1122 4731 4 n_288
rlabel m2contact -1146 4275 -1146 4275 4 n_40
rlabel m2contact -1146 1995 -1146 1995 4 n_40
rlabel m2contact -1170 3891 -1170 3891 4 OpcodeCondIn[2]
rlabel m2contact -1194 4827 -1194 4827 4 n_124
rlabel m2contact -1218 5523 -1218 5523 4 Rs1Sel[0]
rlabel m2contact -1242 4995 -1242 4995 4 n_252
rlabel m2contact -1242 4011 -1242 4011 4 n_86
rlabel m2contact -1266 5523 -1266 5523 4 n_176
rlabel m2contact -1290 5187 -1290 5187 4 n_299
rlabel m2contact -1290 2739 -1290 2739 4 stateSub[0]
rlabel m2contact -1314 4275 -1314 4275 4 n_40
rlabel m2contact -1314 3843 -1314 3843 4 n_248
rlabel m2contact -1362 5187 -1362 5187 4 n_336
rlabel m2contact -1410 2091 -1410 2091 4 n_184
rlabel m2contact -1434 4275 -1434 4275 4 n_317
rlabel m2contact -1554 2283 -1554 2283 4 CFlag
rlabel m2contact -1602 1347 -1602 1347 4 n_334
rlabel m2contact -1650 2091 -1650 2091 4 Op1Sel
rlabel m2contact -1674 5979 -1674 5979 4 n_285
rlabel m2contact -1722 1323 -1722 1323 4 n_33
rlabel m2contact -1746 2019 -1746 2019 4 OpcodeCondIn[4]
rlabel m2contact -1770 3363 -1770 3363 4 n_134
rlabel m2contact -1818 5859 -1818 5859 4 n_12
rlabel m2contact -1842 3099 -1842 3099 4 OpcodeCondIn[3]
rlabel m2contact -1866 3147 -1866 3147 4 n_122
rlabel m2contact -1938 2523 -1938 2523 4 n_81
rlabel m2contact -1986 5955 -1986 5955 4 n_250
rlabel m2contact -1986 5859 -1986 5859 4 n_213
rlabel m2contact -2034 1107 -2034 1107 4 n_315
rlabel m2contact -2034 5931 -2034 5931 4 n_95
rlabel m2contact -2034 4059 -2034 4059 4 n_276
rlabel m2contact -2034 1323 -2034 1323 4 n_276
rlabel m2contact -2058 2835 -2058 2835 4 n_237
rlabel m2contact -2082 5907 -2082 5907 4 n_47
rlabel m2contact -2082 1683 -2082 1683 4 n_364
rlabel m2contact -2106 4155 -2106 4155 4 n_209
rlabel m2contact -2130 2139 -2130 2139 4 n_210
rlabel m2contact -2130 3939 -2130 3939 4 n_191
rlabel m2contact -2154 3411 -2154 3411 4 n_211
rlabel m2contact -2178 4731 -2178 4731 4 n_288
rlabel m2contact -2202 5883 -2202 5883 4 n_62
rlabel m2contact -2226 2835 -2226 2835 4 n_237
rlabel m2contact -2250 3435 -2250 3435 4 n_215
rlabel m2contact -2274 1323 -2274 1323 4 n_276
rlabel m2contact -2274 3411 -2274 3411 4 n_211
rlabel m2contact -2298 4611 -2298 4611 4 n_151
rlabel m2contact -2322 1131 -2322 1131 4 n_99
rlabel m2contact -2346 5883 -2346 5883 4 LrSel
rlabel m2contact -2346 1323 -2346 1323 4 LrSel
rlabel m2contact -2370 5883 -2370 5883 4 LrSel
rlabel m2contact -2370 5139 -2370 5139 4 n_127
rlabel m2contact -2394 1563 -2394 1563 4 n_113
rlabel m2contact -2442 1611 -2442 1611 4 n_263
rlabel m2contact -2466 1779 -2466 1779 4 n_340
rlabel m2contact -2466 4227 -2466 4227 4 n_168
rlabel m2contact -2514 3435 -2514 3435 4 n_215
rlabel m2contact -2514 3315 -2514 3315 4 PcSel[2]
rlabel m2contact -2538 5259 -2538 5259 4 state[0]
rlabel m2contact -2586 4227 -2586 4227 4 n_257
rlabel m2contact -2586 2187 -2586 2187 4 n_257
rlabel m2contact -2610 5139 -2610 5139 4 n_127
rlabel m2contact -2610 3843 -2610 3843 4 n_248
rlabel m2contact -2634 4563 -2634 4563 4 n_85
rlabel m2contact -2634 2499 -2634 2499 4 n_84
rlabel m2contact -2658 5259 -2658 5259 4 state[0]
rlabel m2contact -2682 5403 -2682 5403 4 n_264
rlabel m2contact -2706 4227 -2706 4227 4 n_257
rlabel m2contact -2706 2331 -2706 2331 4 state[1]
rlabel m2contact -2730 5259 -2730 5259 4 state[0]
rlabel m2contact -2754 4659 -2754 4659 4 n_150
rlabel m2contact -2778 4899 -2778 4899 4 n_66
rlabel m2contact -2802 2931 -2802 2931 4 stateSub[1]
rlabel m2contact -2826 1779 -2826 1779 4 n_254
rlabel m2contact -2826 3747 -2826 3747 4 n_282
rlabel m2contact -2850 4179 -2850 4179 4 n_226
rlabel m2contact -2874 3531 -2874 3531 4 n_185
rlabel m2contact -2898 4203 -2898 4203 4 n_178
rlabel m2contact -2922 1275 -2922 1275 4 n_268
rlabel m2contact -2922 3435 -2922 3435 4 n_215
rlabel m2contact -2946 4131 -2946 4131 4 n_174
rlabel m2contact -2970 2931 -2970 2931 4 stateSub[1]
rlabel m2contact -2994 2883 -2994 2883 4 n_359
rlabel m2contact -2994 5739 -2994 5739 4 stateSub[2]
rlabel m2contact -3018 4227 -3018 4227 4 n_301
rlabel m2contact -3018 1563 -3018 1563 4 n_301
rlabel m2contact -3042 4227 -3042 4227 4 n_301
rlabel m2contact -3042 1611 -3042 1611 4 n_322
rlabel m2contact -3066 3195 -3066 3195 4 n_302
rlabel m2contact -3066 3963 -3066 3963 4 n_251
rlabel m2contact -3090 1659 -3090 1659 4 n_217
rlabel m2contact -3114 5715 -3114 5715 4 n_374
rlabel m2contact -3114 1131 -3114 1131 4 n_374
rlabel m2contact -3138 4659 -3138 4659 4 n_150
rlabel m2contact -3162 3963 -3162 3963 4 n_177
rlabel m2contact -3162 3195 -3162 3195 4 n_177
rlabel m2contact -3186 1131 -3186 1131 4 n_374
rlabel m2contact -3186 2427 -3186 2427 4 n_53
rlabel m2contact -3210 2331 -3210 2331 4 state[1]
rlabel m2contact -3234 4227 -3234 4227 4 n_223
rlabel m2contact -3258 5019 -3258 5019 4 ImmSel
rlabel m2contact -3282 2019 -3282 2019 4 OpcodeCondIn[4]
rlabel m2contact -3306 3195 -3306 3195 4 n_177
rlabel m2contact -3306 3915 -3306 3915 4 n_190
rlabel m2contact -3354 3363 -3354 3363 4 n_134
rlabel m2contact -3378 4107 -3378 4107 4 n_117
rlabel m2contact -3402 5739 -3402 5739 4 n_152
rlabel m2contact -3426 5859 -3426 5859 4 n_213
rlabel m2contact -3426 5019 -3426 5019 4 n_212
rlabel m2contact -3450 1611 -3450 1611 4 n_322
rlabel m2contact -3474 4419 -3474 4419 4 n_175
rlabel m2contact -3522 2883 -3522 2883 4 nOE
rlabel m2contact -3546 1155 -3546 1155 4 n_91
rlabel m2contact -3546 4395 -3546 4395 4 n_198
rlabel m2contact -3570 3195 -3570 3195 4 n_319
rlabel m2contact -3594 4395 -3594 4395 4 n_356
rlabel m2contact -3618 1971 -3618 1971 4 n_189
rlabel m2contact -3642 4419 -3642 4419 4 n_92
rlabel m2contact -3642 3915 -3642 3915 4 n_190
rlabel m2contact -3666 5691 -3666 5691 4 OpcodeCondIn[5]
rlabel m2contact -3666 3939 -3666 3939 4 n_191
rlabel m2contact -3690 5835 -3690 5835 4 n_60
rlabel m2contact -3738 4827 -3738 4827 4 n_124
rlabel m2contact -3738 4155 -3738 4155 4 n_209
rlabel m2contact -3762 2187 -3762 2187 4 n_257
rlabel m2contact -3762 3411 -3762 3411 4 n_211
rlabel m2contact -3786 4827 -3786 4827 4 n_41
rlabel m2contact -3810 5835 -3810 5835 4 n_257
rlabel m2contact -3810 2187 -3810 2187 4 n_257
rlabel m2contact -3834 1971 -3834 1971 4 n_158
rlabel m2contact -3858 2331 -3858 2331 4 state[1]
rlabel m2contact -3858 2595 -3858 2595 4 n_220
rlabel m2contact -3882 5835 -3882 5835 4 n_257
rlabel m2contact -3882 3267 -3882 3267 4 n_101
rlabel m2contact -3906 2211 -3906 2211 4 n_160
rlabel m2contact -3930 1203 -3930 1203 4 PcEn
rlabel m2contact -3954 5811 -3954 5811 4 n_208
rlabel m2contact -3954 4395 -3954 4395 4 n_356
rlabel m2contact -3978 1635 -3978 1635 4 n_214
rlabel m2contact -4002 4059 -4002 4059 4 n_276
rlabel m2contact -4050 5787 -4050 5787 4 n_54
rlabel m2contact -4050 5259 -4050 5259 4 state[0]
rlabel m2contact -4050 1203 -4050 1203 4 state[0]
rlabel m2contact -4074 1179 -4074 1179 4 n_137
rlabel m2contact -4074 2427 -4074 2427 4 n_53
rlabel m2contact -4098 4011 -4098 4011 4 n_86
rlabel m2contact -4098 3099 -4098 3099 4 OpcodeCondIn[3]
rlabel m2contact -4122 3003 -4122 3003 4 n_136
rlabel m2contact -4146 5019 -4146 5019 4 n_212
rlabel m2contact -4170 3459 -4170 3459 4 n_59
rlabel m2contact -4170 4203 -4170 4203 4 n_178
rlabel m2contact -4194 1203 -4194 1203 4 state[0]
rlabel m2contact -4194 2139 -4194 2139 4 n_210
rlabel m2contact -4218 3411 -4218 3411 4 n_211
rlabel m2contact -4218 3027 -4218 3027 4 n_58
rlabel m2contact -4266 5019 -4266 5019 4 n_242
rlabel m2contact -4266 3003 -4266 3003 4 n_304
rlabel m2contact -4290 2739 -4290 2739 4 stateSub[0]
rlabel m2contact -4314 4899 -4314 4899 4 n_66
rlabel m2contact -4338 3459 -4338 3459 4 n_238
rlabel m2contact -4410 1227 -4410 1227 4 n_280
rlabel m2contact -4410 5763 -4410 5763 4 n_120
rlabel m2contact -4458 1251 -4458 1251 4 n_103
rlabel m2contact -4458 1851 -4458 1851 4 n_119
rlabel m2contact -4506 5739 -4506 5739 4 n_152
rlabel m2contact -4506 4971 -4506 4971 4 n_253
rlabel m2contact -4530 4611 -4530 4611 4 n_151
rlabel m2contact -4554 3531 -4554 3531 4 n_185
rlabel m2contact -4578 4059 -4578 4059 4 n_276
rlabel m2contact -4602 4707 -4602 4707 4 n_289
rlabel m2contact -4626 5715 -4626 5715 4 n_374
rlabel m2contact -4626 2739 -4626 2739 4 stateSub[0]
rlabel m2contact -4650 5667 -4650 5667 4 n_368
rlabel m2contact -4650 2931 -4650 2931 4 stateSub[1]
rlabel m2contact -4698 4803 -4698 4803 4 n_28
rlabel m2contact -4722 5691 -4722 5691 4 OpcodeCondIn[5]
rlabel m2contact -4722 5667 -4722 5667 4 n_19
rlabel m2contact -4722 2115 -4722 2115 4 n_19
rlabel m2contact -4746 5667 -4746 5667 4 n_19
rlabel m2contact -4746 3675 -4746 3675 4 n_260
rlabel m2contact -4794 5667 -4794 5667 4 LrEn
rlabel m2contact -4794 3723 -4794 3723 4 n_286
rlabel m2contact -4818 4707 -4818 4707 4 n_289
rlabel m2contact -4842 1275 -4842 1275 4 n_268
rlabel m2contact -4866 1443 -4866 1443 4 n_65
rlabel m2contact -4890 5667 -4890 5667 4 LrEn
rlabel m2contact -4914 3627 -4914 3627 4 n_35
rlabel m2contact -4938 1299 -4938 1299 4 n_345
rlabel m2contact -4962 5643 -4962 5643 4 n_197
rlabel m2contact -4986 5619 -4986 5619 4 n_149
rlabel m2contact -5010 1323 -5010 1323 4 LrSel
rlabel m2contact -5010 5259 -5010 5259 4 state[0]
rlabel m2contact -5058 1323 -5058 1323 4 AluEn
rlabel m2contact -5106 1323 -5106 1323 4 AluEn
rlabel m2contact -5106 2859 -5106 2859 4 n_205
rlabel m2contact -5130 1683 -5130 1683 4 n_364
rlabel m2contact -5154 1347 -5154 1347 4 n_334
rlabel m2contact -5154 4659 -5154 4659 4 n_150
rlabel m2contact -5178 3435 -5178 3435 4 n_215
rlabel m2contact -5226 5595 -5226 5595 4 n_163
rlabel m2contact -5226 5571 -5226 5571 4 n_206
rlabel m2contact -5250 1635 -5250 1635 4 n_214
rlabel m2contact -5250 3435 -5250 3435 4 n_116
rlabel m2contact -5274 5499 -5274 5499 4 n_162
rlabel m2contact -5274 2859 -5274 2859 4 n_205
rlabel m2contact -5322 5547 -5322 5547 4 n_133
rlabel m2contact -5322 5499 -5322 5499 4 n_324
rlabel m2contact -5346 1371 -5346 1371 4 Flags[2]
rlabel m2contact -5346 4611 -5346 4611 4 n_151
rlabel m2contact -5370 1395 -5370 1395 4 n_327
rlabel m2contact -5370 1659 -5370 1659 4 n_217
rlabel m2contact -5394 4659 -5394 4659 4 n_150
rlabel m2contact -5442 5523 -5442 5523 4 n_176
rlabel m2contact -5442 4755 -5442 4755 4 n_51
rlabel m2contact -5466 5259 -5466 5259 4 state[0]
rlabel m2contact -5466 3651 -5466 3651 4 n_235
rlabel m2contact -5490 4683 -5490 4683 4 n_147
rlabel m2contact -5538 4683 -5538 4683 4 n_370
rlabel m2contact -5538 2115 -5538 2115 4 n_19
rlabel m2contact -5562 4755 -5562 4755 4 n_350
rlabel m2contact -5586 5499 -5586 5499 4 n_324
rlabel m2contact -5586 2019 -5586 2019 4 OpcodeCondIn[4]
rlabel m2contact -5610 5475 -5610 5475 4 n_293
rlabel m2contact -5658 5451 -5658 5451 4 n_83
rlabel m2contact -5658 3891 -5658 3891 4 OpcodeCondIn[2]
rlabel m2contact -5682 1419 -5682 1419 4 n_484
rlabel m2contact -5682 2499 -5682 2499 4 n_84
rlabel m2contact -5706 5403 -5706 5403 4 n_264
rlabel m2contact -5706 1443 -5706 1443 4 n_65
rlabel m2contact -5754 5427 -5754 5427 4 n_273
rlabel m2contact -5754 5403 -5754 5403 4 n_3
rlabel m2contact -5754 1443 -5754 1443 4 n_3
rlabel m2contact -5778 1443 -5778 1443 4 n_3
rlabel m2contact -5778 5259 -5778 5259 4 state[0]
rlabel m2contact -5802 3483 -5802 3483 4 n_272
rlabel m2contact -5826 2907 -5826 2907 4 nWait
rlabel m2contact -5850 1491 -5850 1491 4 n_31
rlabel m2contact -5874 1467 -5874 1467 4 n_52
rlabel m2contact -5886 5259 -5886 5259 4 state[0]
rlabel m2contact -5886 1491 -5886 1491 4 state[0]
rlabel m2contact -5898 5331 -5898 5331 4 n_6
rlabel m2contact -5922 1491 -5922 1491 4 state[0]
rlabel m2contact -5922 2979 -5922 2979 4 n_30
rlabel m2contact -5970 5331 -5970 5331 4 n_10
rlabel m2contact -5994 5403 -5994 5403 4 n_3
rlabel m2contact -5994 2763 -5994 2763 4 n_321
rlabel m2contact -6018 4059 -6018 4059 4 n_276
rlabel m2contact -6042 2763 -6042 2763 4 n_307
rlabel m2contact -6066 5379 -6066 5379 4 n_312
rlabel m2contact -6090 1515 -6090 1515 4 n_131
rlabel m2contact -6090 3243 -6090 3243 4 n_313
rlabel m2contact -6114 5355 -6114 5355 4 n_164
rlabel m2contact -6114 3099 -6114 3099 4 OpcodeCondIn[3]
rlabel m2contact -6138 3411 -6138 3411 4 n_211
rlabel m2contact -6162 1539 -6162 1539 4 n_73
rlabel m2contact -6186 5331 -6186 5331 4 n_10
rlabel m2contact -6210 5307 -6210 5307 4 n_72
rlabel m2contact -6210 1587 -6210 1587 4 n_487
rlabel m2contact -6234 1923 -6234 1923 4 StatusReg[2]
rlabel m2contact -6258 1611 -6258 1611 4 n_322
rlabel m2contact -6282 1587 -6282 1587 4 ALE
rlabel m2contact -6282 4443 -6282 4443 4 n_88
rlabel m2contact -6306 1563 -6306 1563 4 n_301
rlabel m2contact -6306 1659 -6306 1659 4 n_217
rlabel m2contact -6354 1587 -6354 1587 4 ALE
rlabel m2contact -6402 5283 -6402 5283 4 n_68
rlabel m2contact -6402 4443 -6402 4443 4 n_88
rlabel m2contact -6426 4323 -6426 4323 4 n_42
rlabel m2contact -6426 4011 -6426 4011 4 n_86
rlabel m2contact -6450 3843 -6450 3843 4 n_248
rlabel m2contact -6474 5259 -6474 5259 4 state[0]
rlabel m2contact -6474 5235 -6474 5235 4 AluWe
rlabel m2contact -6498 1611 -6498 1611 4 n_322
rlabel m2contact -6522 5211 -6522 5211 4 n_292
rlabel m2contact -6522 5187 -6522 5187 4 n_336
rlabel m2contact -6570 1683 -6570 1683 4 n_364
rlabel m2contact -6570 2307 -6570 2307 4 n_294
rlabel m2contact -6618 5163 -6618 5163 4 RwSel[0]
rlabel m2contact -6618 1683 -6618 1683 4 SysBus[1]
rlabel m2contact -6642 5139 -6642 5139 4 n_127
rlabel m2contact -6666 5115 -6666 5115 4 n_296
rlabel m2contact -6690 5091 -6690 5091 4 n_314
rlabel m2contact -6690 1635 -6690 1635 4 n_214
rlabel m2contact -6714 1659 -6714 1659 4 n_217
rlabel m2contact -6738 5067 -6738 5067 4 n_352
rlabel m2contact -6738 4059 -6738 4059 4 n_276
rlabel m2contact -6762 1683 -6762 1683 4 SysBus[1]
rlabel m2contact -6786 4491 -6786 4491 4 n_351
rlabel m2contact -6810 4731 -6810 4731 4 n_288
rlabel m2contact -6834 5043 -6834 5043 4 n_277
rlabel m2contact -6834 3627 -6834 3627 4 n_35
rlabel m2contact -6858 4059 -6858 4059 4 n_276
rlabel m2contact -6882 4707 -6882 4707 4 n_289
rlabel m2contact -6906 5019 -6906 5019 4 n_242
rlabel m2contact -6954 1707 -6954 1707 4 n_362
rlabel m2contact -6978 1755 -6978 1755 4 n_89
rlabel m2contact -7002 1731 -7002 1731 4 n_354
rlabel m2contact -7026 1755 -7026 1755 4 LrWe
rlabel m2contact -7050 1755 -7050 1755 4 LrWe
rlabel m2contact -7098 1779 -7098 1779 4 n_254
rlabel m2contact -7122 4995 -7122 4995 4 n_252
rlabel m2contact -7146 4971 -7146 4971 4 n_253
rlabel m2contact -7194 1803 -7194 1803 4 n_114
rlabel m2contact -7218 4947 -7218 4947 4 n_78
rlabel m2contact -7242 4923 -7242 4923 4 n_76
rlabel m2contact -7242 4131 -7242 4131 4 n_174
rlabel m2contact -7266 2859 -7266 2859 4 n_205
rlabel m2contact -7290 3507 -7290 3507 4 n_153
rlabel m2contact -7314 1827 -7314 1827 4 n_135
rlabel m2contact -7314 4923 -7314 4923 4 OpcodeCondIn[4]
rlabel m2contact -7314 2019 -7314 2019 4 OpcodeCondIn[4]
rlabel m2contact -7338 4923 -7338 4923 4 OpcodeCondIn[4]
rlabel m2contact -7338 2715 -7338 2715 4 n_239
rlabel m2contact -7362 1851 -7362 1851 4 n_119
rlabel m2contact -7362 2667 -7362 2667 4 n_146
rlabel m2contact -7410 3123 -7410 3123 4 n_34
rlabel m2contact -7434 2427 -7434 2427 4 n_53
rlabel m2contact -7458 4899 -7458 4899 4 n_66
rlabel m2contact -7458 4875 -7458 4875 4 n_182
rlabel m2contact -7482 3123 -7482 3123 4 n_241
rlabel m2contact -7530 1875 -7530 1875 4 n_100
rlabel m2contact -7578 1899 -7578 1899 4 n_202
rlabel m2contact -7578 3771 -7578 3771 4 n_310
rlabel m2contact -7626 4851 -7626 4851 4 n_221
rlabel m2contact -7626 1971 -7626 1971 4 n_158
rlabel m2contact -7674 1971 -7674 1971 4 SysBus[2]
rlabel m2contact -7674 2211 -7674 2211 4 n_160
rlabel m2contact -7698 4659 -7698 4659 4 n_150
rlabel m2contact -7746 4827 -7746 4827 4 n_41
rlabel m2contact -7770 4203 -7770 4203 4 n_178
rlabel m2contact -7794 3843 -7794 3843 4 n_248
rlabel m2contact -7818 1923 -7818 1923 4 StatusReg[2]
rlabel m2contact -7818 2163 -7818 2163 4 n_159
rlabel m2contact -7866 1947 -7866 1947 4 n_485
rlabel m2contact -7866 4203 -7866 4203 4 n_94
rlabel m2contact -7890 4803 -7890 4803 4 n_28
rlabel m2contact -7914 4779 -7914 4779 4 n_49
rlabel m2contact -7986 2619 -7986 2619 4 n_255
rlabel m2contact -8034 3075 -8034 3075 4 n_194
rlabel m2contact -8082 4755 -8082 4755 4 n_350
rlabel m2contact -8106 1971 -8106 1971 4 SysBus[2]
rlabel m2contact -8130 4491 -8130 4491 4 n_351
rlabel m2contact -8178 4491 -8178 4491 4 n_290
rlabel m2contact -8202 4731 -8202 4731 4 n_288
rlabel m2contact -8226 4707 -8226 4707 4 n_289
rlabel m2contact -8226 4683 -8226 4683 4 n_370
rlabel m2contact -8250 4659 -8250 4659 4 n_150
rlabel m2contact -8274 2931 -8274 2931 4 stateSub[1]
rlabel m2contact -8322 4635 -8322 4635 4 n_22
rlabel m2contact -8346 1995 -8346 1995 4 n_40
rlabel m2contact -8346 2931 -8346 2931 4 stateSub[1]
rlabel m2contact -8370 2019 -8370 2019 4 OpcodeCondIn[4]
rlabel m2contact -8370 2739 -8370 2739 4 stateSub[0]
rlabel m2contact -8394 2043 -8394 2043 4 n_39
rlabel m2contact -8418 2067 -8418 2067 4 n_14
rlabel m2contact -8442 2091 -8442 2091 4 Op1Sel
rlabel m2contact -8442 2811 -8442 2811 4 OpcodeCondIn[7]
rlabel m2contact -8466 3339 -8466 3339 4 n_13
rlabel m2contact -8490 3939 -8490 3939 4 n_191
rlabel m2contact -8514 3219 -8514 3219 4 n_271
rlabel m2contact -8538 3147 -8538 3147 4 n_122
rlabel m2contact -8586 4299 -8586 4299 4 OpcodeCondIn[6]
rlabel m2contact -8586 2499 -8586 2499 4 n_84
rlabel m2contact -8634 3027 -8634 3027 4 n_58
rlabel m2contact -8658 4587 -8658 4587 4 n_121
rlabel m2contact -8706 2811 -8706 2811 4 OpcodeCondIn[7]
rlabel m2contact -8754 3147 -8754 3147 4 n_201
rlabel m2contact -8778 4611 -8778 4611 4 n_151
rlabel m2contact -8778 4587 -8778 4587 4 n_210
rlabel m2contact -8778 2139 -8778 2139 4 n_210
rlabel m2contact -8802 4587 -8802 4587 4 n_210
rlabel m2contact -8802 2715 -8802 2715 4 n_239
rlabel m2contact -8826 2115 -8826 2115 4 n_19
rlabel m2contact -8874 4563 -8874 4563 4 n_85
rlabel m2contact -8874 2235 -8874 2235 4 n_348
rlabel m2contact -8898 4539 -8898 4539 4 n_93
rlabel m2contact -8922 4515 -8922 4515 4 n_26
rlabel m2contact -8922 2235 -8922 2235 4 n_303
rlabel m2contact -8946 4491 -8946 4491 4 n_290
rlabel m2contact -8970 4467 -8970 4467 4 n_156
rlabel m2contact -8994 4443 -8994 4443 4 n_88
rlabel m2contact -9042 3291 -9042 3291 4 n_27
rlabel m2contact -9066 4419 -9066 4419 4 n_92
rlabel m2contact -9090 4395 -9090 4395 4 n_356
rlabel m2contact -9138 4371 -9138 4371 4 n_80
rlabel m2contact -9162 4347 -9162 4347 4 n_79
rlabel m2contact -9162 2187 -9162 2187 4 n_257
rlabel m2contact -9234 4323 -9234 4323 4 n_42
rlabel m2contact -9258 2139 -9258 2139 4 n_210
rlabel m2contact -9306 4299 -9306 4299 4 OpcodeCondIn[6]
rlabel m2contact -9330 2163 -9330 2163 4 n_159
rlabel m2contact -9330 2811 -9330 2811 4 OpcodeCondIn[7]
rlabel m2contact -9354 2187 -9354 2187 4 n_257
rlabel m2contact -9378 2211 -9378 2211 4 n_160
rlabel m2contact -9402 2235 -9402 2235 4 n_303
rlabel m2contact -9426 4275 -9426 4275 4 n_317
rlabel m2contact -9450 4251 -9450 4251 4 n_261
rlabel m2contact -9474 4227 -9474 4227 4 n_223
rlabel m2contact -9474 2739 -9474 2739 4 stateSub[0]
rlabel m2contact -9522 2259 -9522 2259 4 n_155
rlabel m2contact -9546 4203 -9546 4203 4 n_94
rlabel m2contact -9570 2283 -9570 2283 4 CFlag
rlabel m2contact -9570 3531 -9570 3531 4 n_185
rlabel m2contact -9594 2307 -9594 2307 4 n_294
rlabel m2contact -9618 4179 -9618 4179 4 n_226
rlabel m2contact -9666 4155 -9666 4155 4 n_209
rlabel m2contact -9690 4131 -9690 4131 4 n_174
rlabel m2contact -9738 2331 -9738 2331 4 state[1]
rlabel m2contact -9762 3459 -9762 3459 4 n_238
rlabel m2contact -9786 4059 -9786 4059 4 n_276
rlabel m2contact -9810 4083 -9810 4083 4 n_171
rlabel m2contact -9882 3531 -9882 3531 4 n_185
rlabel m2contact -9930 4107 -9930 4107 4 n_117
rlabel m2contact -9978 4083 -9978 4083 4 n_171
rlabel m2contact -10002 2475 -10002 2475 4 n_170
rlabel m2contact -10026 4059 -10026 4059 4 n_276
rlabel m2contact -10074 4035 -10074 4035 4 n_318
rlabel m2contact -10098 4011 -10098 4011 4 n_86
rlabel m2contact -10122 3987 -10122 3987 4 n_275
rlabel m2contact -10170 2355 -10170 2355 4 n_96
rlabel m2contact -10218 2379 -10218 2379 4 n_23
rlabel m2contact -10242 2403 -10242 2403 4 n_45
rlabel m2contact -10290 3963 -10290 3963 4 n_177
rlabel m2contact -10290 2715 -10290 2715 4 n_239
rlabel m2contact -10314 3939 -10314 3939 4 n_191
rlabel m2contact -10338 3915 -10338 3915 4 n_190
rlabel m2contact -10386 2427 -10386 2427 4 n_53
rlabel m2contact -10386 2595 -10386 2595 4 n_220
rlabel m2contact -10410 3891 -10410 3891 4 OpcodeCondIn[2]
rlabel m2contact -10434 3099 -10434 3099 4 OpcodeCondIn[3]
rlabel m2contact -10458 2451 -10458 2451 4 n_199
rlabel m2contact -10482 3867 -10482 3867 4 n_249
rlabel m2contact -10482 3099 -10482 3099 4 OpcodeCondIn[3]
rlabel m2contact -10506 3843 -10506 3843 4 n_248
rlabel m2contact -10506 2475 -10506 2475 4 n_170
rlabel m2contact -10530 3819 -10530 3819 4 n_207
rlabel m2contact -10578 3795 -10578 3795 4 AluOR[1]
rlabel m2contact -10578 2499 -10578 2499 4 n_84
rlabel m2contact -10602 3771 -10602 3771 4 n_310
rlabel m2contact -10602 2523 -10602 2523 4 n_81
rlabel m2contact -10626 3747 -10626 3747 4 n_282
rlabel m2contact -10650 3723 -10650 3723 4 n_286
rlabel m2contact -10650 3699 -10650 3699 4 Op2Sel[1]
rlabel m2contact -10674 2547 -10674 2547 4 n_284
rlabel m2contact -10698 3675 -10698 3675 4 n_260
rlabel m2contact -10722 2571 -10722 2571 4 n_183
rlabel m2contact -10722 3363 -10722 3363 4 n_134
rlabel m2contact -10746 3651 -10746 3651 4 n_235
rlabel m2contact -10794 3627 -10794 3627 4 n_35
rlabel m2contact -10818 3603 -10818 3603 4 OpcodeCondIn[1]
rlabel m2contact -10842 3339 -10842 3339 4 n_13
rlabel m2contact -10890 3579 -10890 3579 4 n_186
rlabel m2contact -10890 3555 -10890 3555 4 WdSel
rlabel m2contact -10914 2811 -10914 2811 4 OpcodeCondIn[7]
rlabel m2contact -10938 3531 -10938 3531 4 n_185
rlabel m2contact -10938 2595 -10938 2595 4 n_220
rlabel m2contact -10962 3507 -10962 3507 4 n_153
rlabel m2contact -10962 2619 -10962 2619 4 n_255
rlabel m2contact -11010 3483 -11010 3483 4 n_272
rlabel m2contact -11010 2643 -11010 2643 4 n_243
rlabel m2contact -11034 2835 -11034 2835 4 n_237
rlabel m2contact -11058 3459 -11058 3459 4 n_238
rlabel m2contact -11058 2667 -11058 2667 4 n_146
rlabel m2contact -11082 2691 -11082 2691 4 n_169
rlabel m2contact -11106 3435 -11106 3435 4 n_116
rlabel m2contact -11130 3411 -11130 3411 4 n_211
rlabel m2contact -11130 3387 -11130 3387 4 n_44
rlabel m2contact -11154 2715 -11154 2715 4 n_239
rlabel m2contact -11154 2787 -11154 2787 4 n_115
rlabel m2contact -11202 3363 -11202 3363 4 n_134
rlabel m2contact -11226 3099 -11226 3099 4 OpcodeCondIn[3]
rlabel m2contact -11250 2811 -11250 2811 4 OpcodeCondIn[7]
rlabel m2contact -11322 3339 -11322 3339 4 n_13
rlabel m2contact -11322 2739 -11322 2739 4 stateSub[0]
rlabel m2contact -11370 2979 -11370 2979 4 n_30
rlabel m2contact -11418 3315 -11418 3315 4 PcSel[2]
rlabel m2contact -11466 3291 -11466 3291 4 n_27
rlabel m2contact -11490 3267 -11490 3267 4 n_101
rlabel m2contact -11562 3243 -11562 3243 4 n_313
rlabel m2contact -11610 3219 -11610 3219 4 n_271
rlabel m2contact -11682 3195 -11682 3195 4 n_319
rlabel m2contact -11730 3003 -11730 3003 4 n_304
rlabel m2contact -11778 2763 -11778 2763 4 n_307
rlabel m2contact -11802 3003 -11802 3003 4 n_246
rlabel m2contact -11826 3171 -11826 3171 4 n_142
rlabel m2contact -11850 3147 -11850 3147 4 n_201
rlabel m2contact -11850 2787 -11850 2787 4 n_115
rlabel m2contact -11898 3123 -11898 3123 4 n_241
rlabel m2contact -11898 2811 -11898 2811 4 OpcodeCondIn[7]
rlabel m2contact -11922 2835 -11922 2835 4 n_237
rlabel m2contact -11946 3099 -11946 3099 4 OpcodeCondIn[3]
rlabel m2contact -11970 3075 -11970 3075 4 n_194
rlabel m2contact -11970 3051 -11970 3051 4 nWE
rlabel m2contact -12018 3027 -12018 3027 4 n_58
rlabel m2contact -12018 3003 -12018 3003 4 n_246
rlabel m2contact -12042 2979 -12042 2979 4 n_30
rlabel m2contact -12042 2955 -12042 2955 4 n_200
rlabel m2contact -12066 2859 -12066 2859 4 n_205
rlabel m2contact -12066 2931 -12066 2931 4 stateSub[1]
rlabel metal1 12897 3183 12897 3183 6 GND!
rlabel metal1 -12158 3183 -12158 3183 4 Vdd!
rlabel metal2 11748 7165 11760 7165 6 StatusRegEn
rlabel metal2 10932 7165 10944 7165 6 StatusReg[3]
rlabel metal2 10116 7165 10128 7165 6 StatusReg[2]
rlabel metal2 9300 7165 9312 7165 6 StatusReg[1]
rlabel metal2 8484 7165 8496 7165 6 StatusReg[0]
rlabel metal2 7668 7165 7680 7165 6 AluEn
rlabel metal2 7644 7165 7656 7165 6 AluWe
rlabel metal2 6828 7165 6840 7165 6 Op2Sel[1]
rlabel metal2 6012 7165 6024 7165 6 Op2Sel[0]
rlabel metal2 4404 7165 4416 7165 6 Op1Sel
rlabel metal2 4308 7165 4320 7165 6 PcEn
rlabel metal2 3564 7165 3576 7165 6 WdSel
rlabel metal2 1956 7165 1968 7165 6 PcWe
rlabel metal2 1140 7165 1152 7165 6 PcSel[2]
rlabel metal2 1116 7165 1128 7165 6 PcSel[1]
rlabel metal2 300 7165 312 7165 6 PcSel[0]
rlabel metal2 -1320 7165 -1308 7165 4 LrEn
rlabel metal2 -2148 7165 -2136 7165 4 LrWe
rlabel metal2 -2364 7165 -2352 7165 4 LrSel
rlabel metal2 -3252 7165 -3240 7165 4 ImmSel
rlabel metal2 -3840 7165 -3828 7165 4 IrWe
rlabel metal2 -4668 7165 -4656 7165 4 MemEn
rlabel metal2 -6288 7165 -6276 7165 4 OpcodeCondIn[7]
rlabel metal2 -7116 7165 -7104 7165 4 OpcodeCondIn[6]
rlabel metal2 -7152 7165 -7140 7165 4 OpcodeCondIn[5]
rlabel metal2 -7980 7165 -7968 7165 4 OpcodeCondIn[4]
rlabel metal2 -9600 7165 -9588 7165 4 OpcodeCondIn[3]
rlabel metal2 -10404 7165 -10392 7165 4 OpcodeCondIn[2]
rlabel metal2 -10812 7165 -10800 7165 4 OpcodeCondIn[1]
rlabel metal2 -11364 7165 -11352 7165 4 OpcodeCondIn[0]
rlabel metal2 9924 -799 9936 -799 8 SysBus[3]
rlabel metal2 336 -799 348 -799 8 SysBus[2]
rlabel metal2 -5868 -799 -5856 -799 2 SysBus[1]
rlabel metal2 -5904 -799 -5892 -799 2 SysBus[0]
rlabel metal2 -12183 -740 -12183 -728 2 nWE
rlabel metal2 -12183 -764 -12183 -752 2 nIRQ
rlabel metal2 12922 -260 12922 -248 8 RegWe
rlabel metal2 12922 -740 12922 -728 8 AluOR[0]
rlabel metal2 12922 -764 12922 -752 8 AluOR[1]
rlabel metal2 12922 -788 12922 -776 8 ENB
rlabel metal2 -12183 2901 -12183 2913 4 nWait
rlabel metal2 -12183 2877 -12183 2889 4 nOE
rlabel metal2 12922 5517 12922 5529 6 Rs1Sel[0]
rlabel metal2 12922 3693 12922 3705 6 Rs1Sel[1]
rlabel metal2 12922 1077 12922 1089 6 RwSel[0]
rlabel metal2 12922 1053 12922 1065 6 RwSel[1]
rlabel metal2 -12183 7022 -12183 7034 4 ALE
rlabel metal2 -12183 6998 -12183 7010 4 nME
rlabel metal2 12922 6926 12922 6938 6 CFlag
rlabel metal2 12922 6902 12922 6914 6 Flags[3]
rlabel metal2 12922 6878 12922 6890 6 Flags[2]
rlabel metal2 12922 6854 12922 6866 6 Flags[1]
rlabel metal2 12922 6830 12922 6842 6 Flags[0]
<< end >>
