magic
tech c035u
timestamp 1393809735
<< metal1 >>
rect 2391 1680 14375 1690
rect 2391 1495 2401 1680
rect 3066 1655 13223 1665
rect 2908 1635 12071 1645
rect 2800 1615 10919 1625
rect 2678 1590 9767 1600
rect 2521 1557 8614 1569
rect 2614 1533 7462 1543
rect 2458 1506 6310 1517
rect 2245 1485 2401 1495
rect 5965 1485 14159 1495
rect 2005 1455 3053 1465
rect 5725 1455 13006 1465
rect 1766 1430 2895 1440
rect 5486 1430 11855 1440
rect 1526 1407 2784 1417
rect 5246 1407 10703 1417
rect 38 1383 1341 1393
rect 1360 1383 1583 1393
rect 1597 1383 1823 1393
rect 1837 1383 2063 1393
rect 3759 1383 5061 1393
rect 5080 1383 5303 1393
rect 5317 1383 5543 1393
rect 5557 1383 5783 1393
rect 325 1358 430 1368
rect 445 1358 911 1368
rect 925 1358 1391 1368
rect 1405 1358 1871 1368
rect 4045 1358 4150 1368
rect 4165 1358 4631 1368
rect 4645 1358 5111 1368
rect 5125 1358 5591 1368
rect 159 1332 887 1342
rect 901 1332 1127 1342
rect 1141 1332 1847 1342
rect 1861 1332 2087 1342
rect 3879 1332 4607 1342
rect 4621 1332 4847 1342
rect 4861 1332 5567 1342
rect 5581 1332 5807 1342
rect 86 1297 383 1307
rect 397 1297 623 1307
rect 637 1297 863 1307
rect 877 1297 1099 1307
rect 1286 1295 2664 1305
rect 3806 1297 4103 1307
rect 4117 1297 4343 1307
rect 4357 1297 4583 1307
rect 4597 1297 4819 1307
rect 5006 1295 9549 1305
rect 278 1275 670 1285
rect 686 1275 723 1285
rect 205 1246 406 1257
rect 422 1246 647 1257
rect 713 1257 723 1275
rect 1047 1273 2506 1283
rect 3998 1275 4390 1285
rect 4406 1275 4443 1285
rect 661 1246 1367 1257
rect 713 1208 723 1246
rect 1381 1246 1607 1257
rect 3925 1246 4126 1257
rect 4142 1246 4367 1257
rect 4433 1257 4443 1275
rect 4767 1273 8399 1283
rect 4381 1246 5087 1257
rect 806 1221 2598 1231
rect 713 1198 1151 1208
rect 1166 1198 1631 1208
rect 1645 1198 2111 1208
rect 4433 1208 4443 1246
rect 5101 1246 5327 1257
rect 4526 1221 7247 1231
rect 4433 1198 4871 1208
rect 4886 1198 5351 1208
rect 5365 1198 5831 1208
rect 565 1176 2444 1187
rect 4285 1176 6095 1187
rect 2894 1144 3023 1154
rect 3037 1144 6455 1154
rect 6469 1144 7607 1154
rect 7622 1144 8759 1154
rect 8773 1144 9911 1154
rect 9925 1144 11063 1154
rect 11077 1144 12214 1154
rect 12229 1144 13367 1154
rect 3613 1107 6023 1117
rect 6037 1107 6239 1117
rect 469 1074 503 1084
rect 709 1075 743 1085
rect 949 1075 983 1085
rect 1190 1080 1223 1090
rect 1429 1080 1463 1090
rect 1669 1080 1703 1090
rect 1909 1080 1943 1090
rect 2150 1080 2182 1090
rect 4189 1074 4223 1084
rect 4429 1075 4463 1085
rect 4669 1075 4703 1085
rect 4910 1080 4943 1090
rect 5149 1080 5183 1090
rect 5389 1080 5423 1090
rect 7044 1094 7175 1104
rect 5629 1080 5663 1090
rect 5870 1080 5902 1090
rect 7189 1094 7391 1104
rect 8196 1094 8327 1104
rect 8341 1094 8543 1104
rect 9348 1094 9479 1104
rect 9493 1094 9695 1104
rect 10500 1094 10631 1104
rect 10645 1094 10847 1104
rect 11652 1094 11783 1104
rect 11797 1094 11999 1104
rect 12804 1094 12935 1104
rect 12949 1094 13151 1104
rect 13956 1094 14087 1104
rect 14101 1094 14303 1104
rect 0 75 2303 85
rect 2317 75 14500 85
rect 0 40 6166 50
rect 6181 40 7318 50
rect 7333 40 8470 50
rect 8485 40 9623 50
rect 9638 40 10773 50
rect 10791 40 11925 50
rect 11943 40 13077 50
rect 13095 40 14231 50
rect 14245 40 14500 50
rect 0 5 6383 15
rect 6397 5 7535 15
rect 7549 5 8687 15
rect 8701 5 9839 15
rect 9854 5 10990 15
rect 11008 5 12142 15
rect 12160 5 13294 15
rect 13312 5 14447 15
rect 14461 5 14500 15
<< m2contact >>
rect 2231 1484 2245 1498
rect 14375 1679 14389 1693
rect 3050 1655 3066 1669
rect 13223 1654 13237 1668
rect 2893 1635 2908 1649
rect 12071 1631 12085 1645
rect 2783 1613 2800 1627
rect 10919 1611 10933 1625
rect 2663 1587 2678 1602
rect 9767 1589 9781 1603
rect 2505 1554 2521 1570
rect 8614 1555 8632 1570
rect 2600 1532 2614 1546
rect 7462 1531 7477 1545
rect 2444 1505 2458 1519
rect 6310 1505 6325 1519
rect 5951 1482 5965 1496
rect 14159 1484 14173 1498
rect 1991 1453 2005 1467
rect 3053 1454 3067 1468
rect 5711 1453 5725 1467
rect 13006 1453 13022 1467
rect 1751 1428 1766 1442
rect 2895 1429 2909 1443
rect 5471 1428 5486 1442
rect 11855 1429 11869 1443
rect 1510 1404 1526 1419
rect 2784 1405 2798 1419
rect 5230 1404 5246 1419
rect 10703 1405 10717 1419
rect 24 1382 38 1396
rect 1341 1381 1360 1397
rect 1583 1380 1597 1394
rect 1823 1382 1837 1396
rect 2063 1382 2078 1396
rect 3744 1382 3759 1396
rect 5061 1381 5080 1397
rect 5303 1380 5317 1394
rect 5543 1382 5557 1396
rect 5783 1382 5798 1396
rect 311 1357 325 1371
rect 430 1357 445 1371
rect 911 1357 925 1371
rect 1391 1357 1405 1371
rect 1871 1356 1886 1370
rect 4031 1357 4045 1371
rect 4150 1357 4165 1371
rect 4631 1357 4645 1371
rect 5111 1357 5125 1371
rect 5591 1356 5606 1370
rect 142 1330 159 1344
rect 887 1332 901 1346
rect 1127 1331 1141 1345
rect 1847 1331 1861 1345
rect 2087 1330 2102 1344
rect 3862 1330 3879 1344
rect 4607 1332 4621 1346
rect 4847 1331 4861 1345
rect 5567 1331 5581 1345
rect 5807 1330 5822 1344
rect 71 1295 86 1309
rect 383 1295 397 1309
rect 623 1296 637 1310
rect 863 1296 877 1310
rect 1099 1295 1116 1312
rect 1269 1293 1286 1307
rect 2664 1294 2678 1308
rect 3791 1295 3806 1309
rect 4103 1295 4117 1309
rect 4343 1296 4357 1310
rect 4583 1296 4597 1310
rect 4819 1295 4836 1312
rect 4989 1293 5006 1307
rect 9549 1293 9568 1310
rect 263 1273 278 1287
rect 670 1269 686 1287
rect 191 1245 205 1259
rect 406 1244 422 1258
rect 647 1245 661 1259
rect 1030 1270 1047 1285
rect 2506 1271 2520 1285
rect 3983 1273 3998 1287
rect 4390 1269 4406 1287
rect 1367 1245 1381 1259
rect 1607 1245 1621 1259
rect 3911 1245 3925 1259
rect 4126 1244 4142 1258
rect 4367 1245 4381 1259
rect 4750 1270 4767 1285
rect 8399 1271 8413 1285
rect 790 1219 806 1233
rect 2598 1220 2612 1234
rect 1151 1197 1166 1211
rect 1631 1197 1645 1211
rect 2111 1197 2125 1211
rect 5087 1245 5101 1259
rect 5327 1245 5341 1259
rect 4510 1219 4526 1233
rect 7247 1220 7262 1234
rect 4871 1197 4886 1211
rect 5351 1197 5365 1211
rect 5831 1197 5845 1211
rect 551 1176 565 1190
rect 2444 1175 2458 1189
rect 4271 1176 4285 1190
rect 6095 1175 6109 1189
rect 2878 1139 2894 1155
rect 3023 1141 3037 1155
rect 6455 1143 6469 1157
rect 7607 1143 7622 1157
rect 8759 1143 8773 1157
rect 9911 1143 9925 1157
rect 11063 1143 11077 1157
rect 12214 1142 12229 1156
rect 13367 1143 13382 1158
rect 3599 1105 3613 1119
rect 6023 1105 6037 1119
rect 6239 1104 6253 1118
rect 455 1071 469 1085
rect 503 1071 517 1085
rect 695 1074 709 1088
rect 743 1073 757 1087
rect 935 1074 949 1088
rect 983 1074 997 1088
rect 1175 1078 1190 1092
rect 1223 1078 1238 1092
rect 1414 1078 1429 1092
rect 1463 1078 1478 1092
rect 1655 1079 1669 1093
rect 1703 1078 1717 1092
rect 1895 1079 1909 1093
rect 1943 1078 1957 1092
rect 2135 1078 2150 1092
rect 2182 1078 2197 1092
rect 4175 1071 4189 1085
rect 4223 1071 4237 1085
rect 4415 1074 4429 1088
rect 4463 1073 4477 1087
rect 4655 1074 4669 1088
rect 4703 1074 4717 1088
rect 4895 1078 4910 1092
rect 4943 1078 4958 1092
rect 5134 1078 5149 1092
rect 5183 1078 5198 1092
rect 5375 1079 5389 1093
rect 5423 1078 5437 1092
rect 5615 1079 5629 1093
rect 7030 1092 7044 1106
rect 5663 1078 5677 1092
rect 5855 1078 5870 1092
rect 5902 1078 5917 1092
rect 7175 1091 7189 1105
rect 7391 1092 7405 1106
rect 8182 1092 8196 1106
rect 8327 1091 8341 1105
rect 8543 1092 8557 1106
rect 9334 1092 9348 1106
rect 9479 1091 9493 1105
rect 9695 1092 9709 1106
rect 10486 1092 10500 1106
rect 10631 1091 10645 1105
rect 10847 1092 10861 1106
rect 11638 1092 11652 1106
rect 11783 1091 11797 1105
rect 11999 1092 12013 1106
rect 12790 1092 12804 1106
rect 12935 1091 12949 1105
rect 13151 1092 13165 1106
rect 13942 1092 13956 1106
rect 14087 1091 14101 1105
rect 14303 1092 14317 1106
rect 2303 74 2317 88
rect 6166 38 6181 52
rect 7318 38 7333 52
rect 8470 38 8485 52
rect 9623 38 9638 53
rect 10773 38 10791 53
rect 11925 38 11943 53
rect 13077 38 13095 53
rect 14231 37 14245 52
rect 6383 4 6397 18
rect 7535 4 7549 18
rect 8687 4 8701 18
rect 9839 3 9854 18
rect 10990 0 11008 15
rect 12142 0 12160 15
rect 13294 0 13312 15
rect 14447 3 14461 18
<< metal2 >>
rect 24 1396 36 1895
rect 24 1068 36 1382
rect 144 1344 156 1895
rect 72 1068 84 1295
rect 144 1068 156 1330
rect 264 1287 276 1895
rect 192 1068 204 1245
rect 264 1068 276 1273
rect 312 1068 324 1357
rect 384 1068 396 1295
rect 408 1068 420 1244
rect 432 1068 444 1357
rect 456 1068 468 1071
rect 504 1068 516 1071
rect 552 1068 564 1176
rect 624 1068 636 1296
rect 648 1068 660 1245
rect 672 1068 684 1269
rect 696 1068 708 1074
rect 744 1068 756 1073
rect 792 1068 804 1219
rect 864 1068 876 1296
rect 888 1068 900 1332
rect 912 1068 924 1357
rect 936 1068 948 1074
rect 984 1068 996 1074
rect 1032 1068 1044 1270
rect 1104 1068 1116 1295
rect 1128 1068 1140 1331
rect 1152 1068 1164 1197
rect 1176 1068 1188 1078
rect 1224 1068 1236 1078
rect 1272 1068 1284 1293
rect 1344 1068 1356 1381
rect 1368 1068 1380 1245
rect 1392 1068 1404 1357
rect 1416 1068 1428 1078
rect 1464 1068 1476 1078
rect 1512 1068 1524 1404
rect 1584 1068 1596 1380
rect 1608 1068 1620 1245
rect 1632 1068 1644 1197
rect 1656 1068 1668 1079
rect 1704 1068 1716 1078
rect 1752 1068 1764 1428
rect 1824 1068 1836 1382
rect 1848 1068 1860 1331
rect 1872 1068 1884 1356
rect 1896 1068 1908 1079
rect 1944 1068 1956 1078
rect 1992 1068 2004 1453
rect 2064 1068 2076 1382
rect 2088 1068 2100 1330
rect 2112 1068 2124 1197
rect 2136 1068 2148 1078
rect 2184 1068 2196 1078
rect 2232 1068 2244 1484
rect 2352 1068 2364 1895
rect 2445 1189 2457 1505
rect 2507 1285 2519 1554
rect 2600 1234 2612 1532
rect 2665 1308 2677 1587
rect 2785 1419 2797 1613
rect 2895 1443 2907 1635
rect 3054 1468 3066 1655
rect 3094 1223 3106 1895
rect 3072 1211 3106 1223
rect 3744 1396 3756 1895
rect 2880 1068 2892 1139
rect 3024 1068 3036 1141
rect 3072 1068 3084 1211
rect 3600 1068 3612 1105
rect 3744 1068 3756 1382
rect 3864 1344 3876 1895
rect 3792 1068 3804 1295
rect 3864 1068 3876 1330
rect 3984 1287 3996 1895
rect 3912 1068 3924 1245
rect 3984 1068 3996 1273
rect 4032 1068 4044 1357
rect 4104 1068 4116 1295
rect 4128 1068 4140 1244
rect 4152 1068 4164 1357
rect 4176 1068 4188 1071
rect 4224 1068 4236 1071
rect 4272 1068 4284 1176
rect 4344 1068 4356 1296
rect 4368 1068 4380 1245
rect 4392 1068 4404 1269
rect 4416 1068 4428 1074
rect 4464 1068 4476 1073
rect 4512 1068 4524 1219
rect 4584 1068 4596 1296
rect 4608 1068 4620 1332
rect 4632 1068 4644 1357
rect 4656 1068 4668 1074
rect 4704 1068 4716 1074
rect 4752 1068 4764 1270
rect 4824 1068 4836 1295
rect 4848 1068 4860 1331
rect 4872 1068 4884 1197
rect 4896 1068 4908 1078
rect 4944 1068 4956 1078
rect 4992 1068 5004 1293
rect 5064 1068 5076 1381
rect 5088 1068 5100 1245
rect 5112 1068 5124 1357
rect 5136 1068 5148 1078
rect 5184 1068 5196 1078
rect 5232 1068 5244 1404
rect 5304 1068 5316 1380
rect 5328 1068 5340 1245
rect 5352 1068 5364 1197
rect 5376 1068 5388 1079
rect 5424 1068 5436 1078
rect 5472 1068 5484 1428
rect 5544 1068 5556 1382
rect 5568 1068 5580 1331
rect 5592 1068 5604 1356
rect 5616 1068 5628 1079
rect 5664 1068 5676 1078
rect 5712 1068 5724 1453
rect 5784 1068 5796 1382
rect 5808 1068 5820 1330
rect 5832 1068 5844 1197
rect 5856 1068 5868 1078
rect 5904 1068 5916 1078
rect 5952 1068 5964 1482
rect 6024 1068 6036 1105
rect 6096 1068 6108 1175
rect 6168 1068 6180 1194
rect 6240 1068 6252 1104
rect 6312 1068 6324 1505
rect 6456 1068 6468 1143
rect 6504 1068 6516 1895
rect 7032 1068 7044 1092
rect 7176 1068 7188 1091
rect 7248 1068 7260 1220
rect 7392 1068 7404 1092
rect 7464 1068 7476 1531
rect 7608 1068 7620 1143
rect 7656 1068 7668 1895
rect 8184 1068 8196 1092
rect 8328 1068 8340 1091
rect 8400 1068 8412 1271
rect 8544 1068 8556 1092
rect 8616 1068 8628 1555
rect 8760 1068 8772 1143
rect 8808 1068 8820 1895
rect 9336 1068 9348 1092
rect 9480 1068 9492 1091
rect 9552 1068 9564 1293
rect 9696 1068 9708 1092
rect 9768 1068 9780 1589
rect 9912 1068 9924 1143
rect 9960 1068 9972 1895
rect 10488 1068 10500 1092
rect 10632 1068 10644 1091
rect 10704 1068 10716 1405
rect 10848 1068 10860 1092
rect 10920 1068 10932 1611
rect 11064 1068 11076 1143
rect 11112 1068 11124 1895
rect 11640 1068 11652 1092
rect 11784 1068 11796 1091
rect 11856 1068 11868 1429
rect 12000 1068 12012 1092
rect 12072 1068 12084 1631
rect 12216 1068 12228 1142
rect 12264 1068 12276 1895
rect 12792 1068 12804 1092
rect 12936 1068 12948 1091
rect 13008 1068 13020 1453
rect 13152 1068 13164 1092
rect 13224 1068 13236 1654
rect 13368 1068 13380 1143
rect 13416 1068 13428 1895
rect 13944 1068 13956 1092
rect 14088 1068 14100 1091
rect 14160 1068 14172 1484
rect 14304 1068 14316 1092
rect 14376 1068 14388 1679
rect 2304 88 2316 269
rect 6168 52 6180 269
rect 6384 18 6396 269
rect 7320 52 7332 269
rect 7536 18 7548 269
rect 8472 52 8484 269
rect 8688 18 8700 269
rect 9624 53 9636 269
rect 9840 18 9852 269
rect 10776 53 10788 269
rect 10992 15 11004 269
rect 11928 53 11940 269
rect 12144 15 12156 269
rect 13080 53 13092 269
rect 13296 15 13308 269
rect 14232 52 14244 269
rect 14448 18 14460 269
use inv inv_11
timestamp 1386238110
transform 1 0 0 0 1 269
box 0 0 120 799
use inv inv_12
timestamp 1386238110
transform 1 0 120 0 1 269
box 0 0 120 799
use inv inv_13
timestamp 1386238110
transform 1 0 240 0 1 269
box 0 0 120 799
use nand3 nand3_8
timestamp 1386234893
transform 1 0 360 0 1 269
box 0 0 120 799
use inv inv_14
timestamp 1386238110
transform 1 0 480 0 1 269
box 0 0 120 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 600 0 1 269
box 0 0 120 799
use inv inv_15
timestamp 1386238110
transform 1 0 720 0 1 269
box 0 0 120 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 840 0 1 269
box 0 0 120 799
use inv inv_16
timestamp 1386238110
transform 1 0 960 0 1 269
box 0 0 120 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 1080 0 1 269
box 0 0 120 799
use inv inv_17
timestamp 1386238110
transform 1 0 1200 0 1 269
box 0 0 120 799
use nand3 nand3_12
timestamp 1386234893
transform 1 0 1320 0 1 269
box 0 0 120 799
use inv inv_18
timestamp 1386238110
transform 1 0 1440 0 1 269
box 0 0 120 799
use nand3 nand3_13
timestamp 1386234893
transform 1 0 1560 0 1 269
box 0 0 120 799
use inv inv_19
timestamp 1386238110
transform 1 0 1680 0 1 269
box 0 0 120 799
use nand3 nand3_14
timestamp 1386234893
transform 1 0 1800 0 1 269
box 0 0 120 799
use inv inv_20
timestamp 1386238110
transform 1 0 1920 0 1 269
box 0 0 120 799
use nand3 nand3_15
timestamp 1386234893
transform 1 0 2040 0 1 269
box 0 0 120 799
use inv inv_21
timestamp 1386238110
transform 1 0 2160 0 1 269
box 0 0 120 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 2280 0 1 269
box 0 0 720 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 3000 0 1 269
box 0 0 720 799
use inv inv_0
timestamp 1386238110
transform 1 0 3720 0 1 269
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 3840 0 1 269
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 3960 0 1 269
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 4080 0 1 269
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 4200 0 1 269
box 0 0 120 799
use nand3 nand3_1
timestamp 1386234893
transform 1 0 4320 0 1 269
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 4440 0 1 269
box 0 0 120 799
use nand3 nand3_2
timestamp 1386234893
transform 1 0 4560 0 1 269
box 0 0 120 799
use inv inv_5
timestamp 1386238110
transform 1 0 4680 0 1 269
box 0 0 120 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 4800 0 1 269
box 0 0 120 799
use inv inv_6
timestamp 1386238110
transform 1 0 4920 0 1 269
box 0 0 120 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 5040 0 1 269
box 0 0 120 799
use inv inv_7
timestamp 1386238110
transform 1 0 5160 0 1 269
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 5280 0 1 269
box 0 0 120 799
use inv inv_8
timestamp 1386238110
transform 1 0 5400 0 1 269
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 5520 0 1 269
box 0 0 120 799
use inv inv_9
timestamp 1386238110
transform 1 0 5640 0 1 269
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 5760 0 1 269
box 0 0 120 799
use inv inv_10
timestamp 1386238110
transform 1 0 5880 0 1 269
box 0 0 120 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 6000 0 1 269
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 6216 0 1 269
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 6432 0 1 269
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 7152 0 1 269
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 7368 0 1 269
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 7584 0 1 269
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 8304 0 1 269
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 8520 0 1 269
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 8736 0 1 269
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 9456 0 1 269
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 9672 0 1 269
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 9888 0 1 269
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 10608 0 1 269
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 10824 0 1 269
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 11040 0 1 269
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 11760 0 1 269
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 11976 0 1 269
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 12192 0 1 269
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 12912 0 1 269
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 13128 0 1 269
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 13344 0 1 269
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 14064 0 1 269
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 14280 0 1 269
box 0 0 216 799
<< labels >>
rlabel metal2 24 1895 36 1895 5 Rs2[0]
rlabel metal2 144 1895 156 1895 5 Rs2[1]
rlabel metal2 264 1895 276 1895 5 Rs2[2]
rlabel metal2 3744 1895 3756 1895 5 Rs1[0]
rlabel metal2 3864 1895 3876 1895 5 Rs1[1]
rlabel metal2 3984 1895 3996 1895 5 Rs1[2]
rlabel metal2 2352 1895 2364 1895 5 IRWe
rlabel metal1 0 75 0 85 3 Databus
rlabel metal1 0 40 0 50 3 Rd1[0]
rlabel metal1 0 5 0 15 3 Rd2[0]
rlabel metal1 14500 75 14500 85 7 Databus
rlabel metal1 14500 40 14500 50 7 Rd1[0]
rlabel metal1 14500 5 14500 15 7 Rd2[0]
rlabel metal2 3094 1895 3106 1895 5 WData[0]
rlabel metal2 6504 1895 6516 1895 5 WData[1]
rlabel metal2 7656 1895 7668 1895 5 WData[2]
rlabel metal2 8808 1895 8820 1895 5 WData[3]
rlabel metal2 9960 1895 9972 1895 5 WData[4]
rlabel metal2 11112 1895 11124 1895 5 WData[5]
rlabel metal2 12264 1895 12276 1895 5 WData[6]
rlabel metal2 13416 1895 13428 1895 5 WData[7]
<< end >>
