magic
tech c035u
timestamp 1394548889
<< checkpaint >>
rect 0 17608 25377 22003
rect 2009 -1208 25377 17608
<< metal1 >>
rect 481 21074 16244 21084
rect 16258 21074 23668 21084
rect 504 21050 16364 21060
rect 16378 21050 23668 21060
rect 527 21026 16484 21036
rect 16498 21026 23668 21036
rect 550 21002 16604 21012
rect 16618 21002 23668 21012
rect 573 20978 16724 20988
rect 16738 20978 23668 20988
rect 596 20954 5228 20964
rect 5242 20954 23668 20964
rect 619 20930 5420 20940
rect 5434 20930 23668 20940
rect 642 20906 5612 20916
rect 5626 20906 23668 20916
rect 665 20882 5276 20892
rect 5290 20882 23668 20892
rect 688 20858 5468 20868
rect 5482 20858 23668 20868
rect 711 20834 5660 20844
rect 5674 20834 23668 20844
rect 734 20810 6932 20820
rect 6946 20810 23668 20820
rect 757 20786 6908 20796
rect 6922 20786 22364 20796
rect 22378 20786 23668 20796
rect 780 20762 6884 20772
rect 6898 20762 22580 20772
rect 22594 20762 23668 20772
rect 803 20738 22700 20748
rect 22714 20738 23668 20748
rect 826 20714 22820 20724
rect 22834 20714 23668 20724
rect 0 17893 467 17903
rect 481 17893 832 17903
rect 0 17827 832 17837
rect 0 16717 490 16727
rect 504 16717 832 16727
rect 0 16651 832 16661
rect 0 15541 513 15551
rect 527 15541 832 15551
rect 0 15475 832 15485
rect 0 14365 536 14375
rect 550 14365 832 14375
rect 0 14299 832 14309
rect 0 13189 559 13199
rect 573 13189 832 13199
rect 0 13123 832 13133
rect 0 12013 582 12023
rect 596 12013 832 12023
rect 0 11947 832 11957
rect 0 10837 605 10847
rect 619 10837 832 10847
rect 0 10771 832 10781
rect 0 9661 628 9671
rect 642 9661 832 9671
rect 0 9595 832 9605
rect 0 8485 651 8495
rect 665 8485 832 8495
rect 0 8419 832 8429
rect 0 7309 674 7319
rect 688 7309 832 7319
rect 0 7243 832 7253
rect 0 6133 697 6143
rect 711 6133 832 6143
rect 0 6067 832 6077
rect 0 4957 720 4967
rect 734 4957 832 4967
rect 0 4891 832 4901
rect 0 3781 743 3791
rect 757 3781 832 3791
rect 0 3715 832 3725
rect 0 2605 766 2615
rect 780 2605 832 2615
rect 0 2539 832 2549
rect 0 1429 789 1439
rect 803 1429 832 1439
rect 0 1363 832 1373
rect 0 253 812 263
rect 826 253 832 263
rect 0 187 832 197
rect 2306 72 3524 82
rect 3538 72 23877 82
<< m2contact >>
rect 467 21072 481 21086
rect 16244 21073 16258 21087
rect 490 21048 504 21062
rect 16364 21048 16378 21062
rect 513 21024 527 21038
rect 16484 21024 16498 21038
rect 536 21000 550 21014
rect 16604 21000 16618 21014
rect 559 20976 573 20990
rect 16724 20976 16738 20990
rect 582 20952 596 20966
rect 5228 20952 5242 20966
rect 605 20928 619 20942
rect 5420 20928 5434 20942
rect 628 20904 642 20918
rect 5612 20904 5626 20918
rect 651 20880 665 20894
rect 5276 20880 5290 20894
rect 674 20856 688 20870
rect 5468 20856 5482 20870
rect 697 20832 711 20846
rect 5660 20832 5674 20846
rect 720 20808 734 20822
rect 6932 20808 6946 20822
rect 743 20784 757 20798
rect 6908 20784 6922 20798
rect 22364 20784 22378 20798
rect 766 20760 780 20774
rect 6884 20760 6898 20774
rect 22580 20759 22594 20773
rect 789 20736 803 20750
rect 22700 20736 22714 20750
rect 812 20712 826 20726
rect 22820 20712 22834 20726
rect 467 17891 481 17905
rect 490 16715 504 16729
rect 513 15539 527 15553
rect 536 14363 550 14377
rect 559 13187 573 13201
rect 582 12011 596 12025
rect 605 10835 619 10849
rect 628 9659 642 9673
rect 651 8483 665 8497
rect 674 7307 688 7321
rect 697 6131 711 6145
rect 720 4955 734 4969
rect 743 3779 757 3793
rect 766 2603 780 2617
rect 789 1427 803 1441
rect 812 251 826 265
rect 3524 70 3538 84
rect 23877 70 23891 84
<< metal2 >>
rect 468 17905 480 21072
rect 491 16729 503 21048
rect 514 15553 526 21024
rect 537 14377 549 21000
rect 560 13201 572 20976
rect 583 12025 595 20952
rect 606 10849 618 20928
rect 629 9673 641 20904
rect 652 8497 664 20880
rect 675 7321 687 20856
rect 698 6145 710 20832
rect 721 4969 733 20808
rect 744 3793 756 20784
rect 767 2617 779 20760
rect 790 1441 802 20736
rect 813 265 825 20712
rect 837 20703 1037 21230
rect 1053 20703 1065 21230
rect 1077 20703 1089 21230
rect 1101 20703 1113 21230
rect 1125 20703 1137 21230
rect 5205 20703 5217 21230
rect 5229 20703 5241 20952
rect 5277 20703 5289 20880
rect 5421 20703 5433 20928
rect 5469 20703 5481 20856
rect 5613 20703 5625 20904
rect 5661 20703 5673 20832
rect 5829 20703 5841 21230
rect 6575 20703 6587 21230
rect 6885 20703 6897 20760
rect 6909 20703 6921 20784
rect 6933 20703 6945 20808
rect 16245 20703 16257 21073
rect 16365 20703 16377 21048
rect 16485 20703 16497 21024
rect 16605 20703 16617 21000
rect 16725 20703 16737 20976
rect 17901 20703 17913 21230
rect 18333 20703 18345 21230
rect 18525 20703 18537 21230
rect 18597 20703 18609 21230
rect 18693 20703 18705 21230
rect 22365 20703 22377 20784
rect 22581 20703 22593 20759
rect 22701 20703 22713 20736
rect 22821 20703 22833 20712
rect 23205 20703 23217 21230
rect 23877 20703 24077 21230
rect 837 0 1037 92
rect 1053 0 1065 92
rect 1077 0 1089 92
rect 1101 0 1113 92
rect 1125 0 1137 92
rect 2373 0 2385 92
rect 3165 0 3177 93
rect 3525 84 3537 92
rect 3669 0 3681 92
rect 3885 0 3897 92
rect 4629 0 4641 92
rect 4797 0 4809 92
rect 5181 0 5193 92
rect 5397 0 5409 92
rect 6141 0 6153 92
rect 6309 0 6321 92
rect 15717 0 15729 92
rect 15909 0 15921 92
rect 16749 0 16761 92
rect 17037 0 17049 92
rect 19701 0 19713 92
rect 19749 0 19761 92
rect 19797 0 19809 92
rect 19845 0 19857 92
rect 19893 0 19905 92
rect 19941 0 19953 92
rect 19989 0 20001 92
rect 20037 0 20049 92
rect 20349 0 20361 92
rect 20397 0 20409 92
rect 20445 0 20457 92
rect 20493 0 20505 92
rect 20805 0 20817 92
rect 20853 0 20865 92
rect 21237 0 21249 92
rect 21477 0 21489 92
rect 21525 0 21537 92
rect 21573 0 21585 92
rect 21621 0 21633 92
rect 21669 0 21681 92
rect 21717 0 21729 92
rect 21765 0 21777 92
rect 21813 0 21825 92
rect 22125 0 22137 92
rect 22173 0 22185 92
rect 22221 0 22233 92
rect 22269 0 22281 92
rect 22581 0 22593 92
rect 22629 0 22641 92
rect 22941 0 22953 92
rect 23229 0 23241 92
rect 23637 0 23649 92
rect 23877 84 24077 92
rect 23891 70 24077 84
rect 23877 0 24077 70
use slice17 slice17_0
timestamp 1394548889
transform 1 0 5166 0 1 18908
box -4329 0 18911 1795
use leftbuf_slice leftbuf_slice_0
array 0 0 1469 0 15 1176
timestamp 1394489502
transform 1 0 832 0 1 98
box 0 -6 1469 1170
use IrAA IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 2301 0 1 9611
box 0 -111 1008 1065
use LLIcell_U LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1393855556
transform 1 0 23349 0 1 9611
box 0 0 192 1042
use IrBA IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 2301 0 1 6083
box 0 -111 1008 1065
use IrBB IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 2301 0 1 204
box 0 -112 1008 1064
use LLIcell_L LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23349 0 1 203
box 0 0 192 1042
use Datapath_slice Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394548889
transform 1 0 3309 0 1 92
box 0 0 20768 1176
<< labels >>
rlabel metal1 0 187 0 197 3 SysBus[0]
rlabel metal1 0 1363 0 1373 3 SysBus[1]
rlabel metal1 0 2539 0 2549 3 SysBus[2]
rlabel metal1 0 3715 0 3725 3 SysBus[3]
rlabel metal1 0 4891 0 4901 3 SysBus[4]
rlabel metal1 0 6067 0 6077 3 SysBus[5]
rlabel metal1 0 7243 0 7253 3 SysBus[6]
rlabel metal1 0 8419 0 8429 3 SysBus[7]
rlabel metal1 0 9595 0 9605 3 SysBus[8]
rlabel metal1 0 10771 0 10781 3 SysBus[9]
rlabel metal1 0 11947 0 11957 3 SysBus[10]
rlabel metal1 0 13123 0 13133 3 SysBus[11]
rlabel metal1 0 14299 0 14309 3 SysBus[12]
rlabel metal1 0 15475 0 15485 3 SysBus[13]
rlabel metal1 0 16651 0 16661 3 SysBus[14]
rlabel metal1 0 17827 0 17837 3 SysBus[15]
rlabel metal1 0 253 0 263 3 Ir[0]
rlabel metal1 0 1429 0 1439 3 Ir[1]
rlabel metal1 0 2605 0 2615 3 Ir[2]
rlabel metal1 0 3781 0 3791 3 Ir[3]
rlabel metal1 0 4957 0 4967 3 Ir[4]
rlabel metal1 0 6133 0 6143 3 Ir[5]
rlabel metal1 0 7309 0 7319 3 Ir[6]
rlabel metal1 0 8485 0 8495 3 Ir[7]
rlabel metal1 0 9661 0 9671 3 Ir[8]
rlabel metal1 0 10837 0 10847 3 Ir[9]
rlabel metal1 0 12013 0 12023 3 Ir[10]
rlabel metal1 0 13189 0 13199 3 Ir[11]
rlabel metal1 0 14365 0 14375 3 Ir[12]
rlabel metal1 0 15541 0 15551 3 Ir[13]
rlabel metal1 0 16717 0 16727 3 Ir[14]
rlabel metal1 0 17893 0 17903 3 Ir[15]
rlabel metal2 3669 0 3681 0 1 LrSel
rlabel metal2 3885 0 3897 0 1 LrWe
rlabel metal2 4629 0 4641 0 1 LrEn
rlabel metal2 4797 0 4809 0 1 PcSel[0]
rlabel metal2 5181 0 5193 0 1 PcSel[1]
rlabel metal2 5397 0 5409 0 1 PcWe
rlabel metal2 6141 0 6153 0 1 PcEn
rlabel metal2 6309 0 6321 0 1 WdSel
rlabel metal2 15909 0 15921 0 1 Op2Sel
rlabel metal2 15717 0 15729 0 1 Op1Sel
rlabel metal2 16749 0 16761 0 1 CIn_Slice
rlabel metal2 19749 0 19761 0 1 Sh8B_L
rlabel metal2 19797 0 19809 0 1 Sh8C_L
rlabel metal2 19701 0 19713 0 1 Sh8A_L
rlabel metal2 21813 0 21825 0 1 Sh8G_R
rlabel metal2 21765 0 21777 0 1 Sh8F_R
rlabel metal2 21717 0 21729 0 1 Sh8E_R
rlabel metal2 21669 0 21681 0 1 Sh8D_R
rlabel metal2 21621 0 21633 0 1 Sh8C_R
rlabel metal2 23229 0 23241 0 1 ShOut
rlabel metal2 22269 0 22281 0 1 Sh4B_R
rlabel metal2 22221 0 22233 0 1 Sh4A_R
rlabel metal2 22173 0 22185 0 1 Sh4Z_R
rlabel metal2 22581 0 22593 0 1 Sh2Z_R
rlabel metal2 22629 0 22641 0 1 Sh2A_R
rlabel metal2 22941 0 22953 0 1 Sh1_R_Out
rlabel metal2 22125 0 22137 0 1 Sh4Y_L
rlabel metal2 20037 0 20049 0 1 Sh8H_L
rlabel metal2 20349 0 20361 0 1 Sh4A_L
rlabel metal2 20805 0 20817 0 1 Sh2B_L
rlabel metal2 20853 0 20865 0 1 Sh2C_L
rlabel metal2 20397 0 20409 0 1 Sh4B_L
rlabel metal2 20445 0 20457 0 1 Sh4C_L
rlabel metal2 20493 0 20505 0 1 Sh4D_L
rlabel metal2 21573 0 21585 0 1 Sh8B_R
rlabel metal2 21525 0 21537 0 1 Sh8A_R
rlabel metal2 21477 0 21489 0 1 Sh8Z_R
rlabel metal2 21237 0 21249 0 1 Sh1_L_In
rlabel metal2 19845 0 19857 0 1 Sh8D_L
rlabel metal2 19893 0 19905 0 1 Sh8E_L
rlabel metal2 19941 0 19953 0 1 Sh8F_L
rlabel metal2 19989 0 20001 0 1 Sh8G_L
rlabel metal2 23877 0 24077 0 1 GND!
rlabel metal2 17037 0 17049 0 1 nZ_prev
rlabel metal2 23637 0 23649 0 1 AluEn
rlabel metal2 837 0 1037 0 1 Vdd!
rlabel metal2 1053 0 1065 0 1 SDI
rlabel metal2 1077 0 1089 0 1 Test
rlabel metal2 1101 0 1113 0 1 Clock
rlabel metal2 1125 0 1137 0 1 nReset
rlabel metal2 3165 0 3177 0 1 ImmSel
rlabel metal2 2373 0 2385 0 1 IrWe
rlabel m2contact 750 20781 750 20781 1 Ir[3]
rlabel metal2 727 20782 727 20782 1 Ir[4]
rlabel metal2 704 20781 704 20781 1 Ir[5]
rlabel metal2 681 20780 681 20780 1 Ir[6]
rlabel metal2 658 20779 658 20779 1 Ir[7]
rlabel metal2 635 20777 635 20777 1 Ir[8]
rlabel metal2 612 20777 612 20777 1 Ir[9]
rlabel metal2 589 20776 589 20776 1 Ir[10]
rlabel metal2 566 20777 566 20777 1 Ir[11]
rlabel metal2 543 20777 543 20777 1 Ir[12]
rlabel metal2 520 20776 520 20776 1 Ir[13]
rlabel metal2 497 20776 497 20776 1 Ir[14]
rlabel metal2 473 20777 473 20777 1 Ir[15]
rlabel metal2 1053 21230 1065 21230 1 SDI
rlabel metal2 1077 21230 1089 21230 1 Test
rlabel metal2 1101 21230 1113 21230 1 Clock
rlabel metal2 1125 21230 1137 21230 1 nReset
rlabel metal2 837 21230 1037 21230 5 Vdd!
rlabel metal2 5829 21230 5841 21230 5 RwSel
rlabel metal2 5205 21230 5217 21230 5 Rs1Sel
rlabel metal2 6575 21230 6587 21230 5 RegWe
rlabel metal2 17901 21230 17913 21230 5 CFlag
rlabel metal2 18333 21230 18345 21230 5 Flags[2]
rlabel metal2 18525 21230 18537 21230 5 Flags[1]
rlabel metal2 18597 21230 18609 21230 5 Flags[3]
rlabel metal2 23205 21230 23217 21230 5 AluEn
rlabel metal2 23877 21230 24077 21230 1 GND!
rlabel metal2 18693 21230 18705 21230 5 Flags[0]
rlabel metal1 5249 20959 5249 20959 1 Ir[10]
rlabel metal2 5234 20945 5234 20945 1 Ir[10]
rlabel metal2 5283 20872 5283 20872 1 Ir[7]
rlabel metal2 5426 20920 5426 20920 1 Ir[9]
rlabel metal2 5475 20849 5475 20849 1 Ir[6]
rlabel metal2 5618 20897 5618 20897 1 Ir[8]
rlabel metal2 5668 20826 5668 20826 1 Ir[5]
rlabel metal2 6889 20752 6889 20752 1 Ir[2]
rlabel metal2 6915 20776 6915 20776 1 Ir[3]
rlabel metal2 6938 20800 6938 20800 1 Ir[4]
rlabel metal2 16250 21066 16250 21066 1 Ir[15]
rlabel metal2 16369 21041 16369 21041 1 Ir[14]
rlabel metal2 16490 21018 16490 21018 1 Ir[13]
rlabel metal2 16611 20994 16611 20994 1 Ir[12]
rlabel metal2 16731 20969 16731 20969 1 Ir[11]
rlabel metal2 22371 20779 22371 20779 1 Ir[3]
rlabel metal2 22586 20754 22586 20754 1 Ir[2]
rlabel metal2 22706 20729 22706 20729 1 Ir[1]
rlabel metal2 22827 20707 22827 20707 1 Ir[0]
<< end >>
