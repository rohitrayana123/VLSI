../behavioural/opcodes.svh