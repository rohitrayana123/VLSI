magic
tech c035u
timestamp 1394633578
<< metal1 >>
rect 3085 1355 3263 1365
rect 3277 1355 3407 1365
rect 3421 1355 3551 1365
rect 3565 1355 3695 1365
rect 1093 1333 1247 1343
rect 2965 1333 3839 1343
rect 3853 1333 3983 1343
rect 3997 1333 4127 1343
rect 4141 1333 4535 1343
rect 6181 1334 6335 1344
rect 6877 1333 7223 1343
rect 997 1311 1151 1321
rect 1285 1311 1463 1321
rect 1501 1311 1559 1321
rect 2845 1311 3119 1321
rect 5005 1311 5207 1321
rect 5677 1311 5879 1321
rect 5917 1311 6215 1321
rect 6229 1311 6407 1321
rect 6421 1311 6527 1321
rect 6541 1311 6647 1321
rect 6997 1311 7199 1321
rect 877 1289 1127 1299
rect 1189 1289 1319 1299
rect 1381 1289 1535 1299
rect 1861 1289 1895 1299
rect 2125 1289 2399 1299
rect 2725 1289 4271 1299
rect 4285 1289 4391 1299
rect 4765 1289 4799 1299
rect 5149 1289 5183 1299
rect 5269 1289 5303 1299
rect 5821 1289 5855 1299
rect 6061 1289 6095 1299
rect 6277 1290 6311 1300
rect 7141 1289 7175 1299
rect 685 1267 959 1277
rect 973 1267 1055 1277
rect 1069 1267 3167 1277
rect 3181 1267 3311 1277
rect 3325 1267 3743 1277
rect 3757 1267 3887 1277
rect 3901 1267 4175 1277
rect 4189 1267 4439 1277
rect 4453 1267 4943 1277
rect 4957 1267 5639 1277
rect 5653 1267 7103 1277
rect 565 1245 1343 1255
rect 1357 1245 1656 1255
rect 1670 1245 3287 1255
rect 3301 1245 3431 1255
rect 3445 1245 4151 1255
rect 4165 1245 4295 1255
rect 4309 1245 4415 1255
rect 4429 1245 4559 1255
rect 4573 1245 4703 1255
rect 4717 1245 4919 1255
rect 445 1223 935 1233
rect 949 1223 2687 1233
rect 2701 1223 2927 1233
rect 2941 1223 5615 1233
rect 5629 1223 5759 1233
rect 5773 1223 6935 1233
rect 6949 1223 7079 1233
rect 325 1201 791 1211
rect 805 1201 1439 1211
rect 1453 1201 2663 1211
rect 2677 1201 2783 1211
rect 2797 1201 4679 1211
rect 4693 1201 4895 1211
rect 4909 1201 5591 1211
rect 5605 1201 5735 1211
rect 5749 1201 5975 1211
rect 5989 1201 6791 1211
rect 6805 1201 7055 1211
rect 205 1179 1631 1189
rect 1645 1179 2639 1189
rect 2653 1179 2759 1189
rect 2773 1179 2879 1189
rect 2893 1179 2999 1189
rect 3013 1179 4823 1189
rect 4837 1179 5567 1189
rect 5581 1179 5711 1189
rect 5725 1179 6767 1189
rect 6781 1179 6911 1189
rect 6925 1179 7031 1189
rect 0 1157 172 1167
rect 7320 1157 7822 1167
rect 0 1134 168 1144
rect 7320 1134 7822 1144
rect 0 1096 168 1121
rect 7320 1096 7822 1121
rect 0 451 168 476
rect 7320 451 7822 476
rect 0 428 168 438
rect 7317 428 7822 438
rect 0 405 169 415
rect 7320 405 7822 415
rect 0 382 168 392
rect 7320 382 7822 392
rect 253 360 911 370
rect 925 360 1415 370
rect 1429 360 5327 370
rect 5341 360 5951 370
rect 373 338 2903 348
rect 2917 338 3023 348
rect 3037 338 5039 348
rect 493 316 815 326
rect 829 316 1031 326
rect 1045 316 1223 326
rect 1237 316 1679 326
rect 1693 316 2807 326
rect 2821 316 3047 326
rect 3061 316 5351 326
rect 5365 316 5999 326
rect 613 294 3143 304
rect 3157 294 3575 304
rect 3589 294 3719 304
rect 3733 294 3863 304
rect 3877 294 4007 304
rect 4021 294 5063 304
rect 5077 294 5783 304
rect 5797 294 6119 304
rect 6133 294 6815 304
rect 6829 294 6959 304
rect 733 272 839 282
rect 853 272 3455 282
rect 3469 272 3599 282
rect 3613 272 4031 282
rect 4045 272 4583 282
rect 4597 272 4727 282
rect 4741 272 5087 282
rect 5101 272 6143 282
rect 6157 272 6839 282
rect 7309 272 7727 282
rect 349 250 1583 260
rect 1597 250 1919 260
rect 1933 250 2279 260
rect 4501 250 5471 260
rect 5533 250 5879 260
rect 7261 250 7319 260
rect 1741 228 1799 238
rect 3349 228 5447 238
rect 5509 228 6359 238
rect 517 206 2015 216
rect 4645 206 7487 216
rect 685 184 2087 194
rect 4357 177 5520 187
rect 6157 184 6479 194
rect 6733 184 6959 194
rect 709 162 2303 172
rect 781 140 2471 150
rect 997 118 2519 128
rect 85 96 3215 106
rect 1477 70 3359 80
rect 1837 48 3503 58
rect 2245 21 3647 31
rect 2581 -4 3791 6
rect 2893 -26 3935 -16
rect 3229 -48 4079 -38
rect 3397 -70 4223 -60
rect 3565 -92 5399 -82
rect 1141 -114 4847 -104
<< m2contact >>
rect 3071 1353 3085 1367
rect 3263 1353 3277 1367
rect 3407 1353 3421 1367
rect 3551 1353 3565 1367
rect 3695 1353 3709 1367
rect 1079 1331 1093 1345
rect 1247 1331 1261 1345
rect 2951 1331 2965 1345
rect 3839 1331 3853 1345
rect 3983 1331 3997 1345
rect 4127 1331 4141 1345
rect 4535 1331 4549 1345
rect 6167 1332 6181 1346
rect 6335 1332 6349 1346
rect 6863 1331 6877 1345
rect 7223 1331 7237 1345
rect 983 1309 997 1323
rect 1151 1309 1165 1323
rect 1271 1309 1285 1323
rect 1463 1309 1477 1323
rect 1487 1309 1501 1323
rect 1559 1309 1573 1323
rect 2831 1309 2845 1323
rect 3119 1309 3133 1323
rect 4991 1309 5005 1323
rect 5207 1309 5221 1323
rect 5663 1309 5677 1323
rect 5879 1309 5893 1323
rect 5903 1309 5917 1323
rect 6215 1309 6229 1323
rect 6407 1309 6421 1323
rect 6527 1309 6541 1323
rect 6647 1309 6661 1323
rect 6983 1309 6997 1323
rect 7199 1309 7213 1323
rect 863 1287 877 1301
rect 1127 1287 1141 1301
rect 1175 1288 1189 1302
rect 1319 1287 1333 1301
rect 1367 1287 1381 1301
rect 1535 1287 1549 1301
rect 1847 1287 1861 1301
rect 1895 1287 1909 1301
rect 2111 1287 2125 1301
rect 2399 1287 2413 1301
rect 2711 1287 2725 1301
rect 4271 1287 4285 1301
rect 4391 1287 4405 1301
rect 4751 1287 4765 1301
rect 4799 1287 4813 1301
rect 5135 1287 5149 1301
rect 5183 1287 5197 1301
rect 5255 1287 5269 1301
rect 5303 1287 5317 1301
rect 5807 1287 5821 1301
rect 5855 1287 5869 1301
rect 6047 1287 6061 1301
rect 6095 1287 6109 1301
rect 6263 1287 6277 1301
rect 6311 1287 6325 1301
rect 7127 1287 7141 1301
rect 7175 1287 7189 1301
rect 671 1265 685 1279
rect 959 1265 973 1279
rect 1055 1265 1069 1279
rect 3167 1265 3181 1279
rect 3311 1265 3325 1279
rect 3743 1265 3757 1279
rect 3887 1265 3901 1279
rect 4175 1265 4189 1279
rect 4439 1266 4453 1280
rect 4943 1264 4957 1278
rect 5639 1265 5653 1279
rect 7103 1265 7117 1279
rect 551 1243 565 1257
rect 1343 1243 1357 1257
rect 1656 1243 1670 1257
rect 3287 1243 3301 1257
rect 3431 1243 3445 1257
rect 4151 1243 4165 1257
rect 4295 1243 4309 1257
rect 4415 1243 4429 1257
rect 4559 1243 4573 1257
rect 4703 1243 4717 1257
rect 4919 1243 4933 1257
rect 431 1221 445 1235
rect 935 1221 949 1235
rect 2687 1221 2701 1235
rect 2927 1221 2941 1235
rect 5615 1221 5629 1235
rect 5759 1221 5773 1235
rect 6935 1221 6949 1235
rect 7079 1221 7093 1235
rect 311 1199 325 1213
rect 791 1199 805 1213
rect 1439 1199 1453 1213
rect 2663 1199 2677 1213
rect 2783 1199 2797 1213
rect 4679 1199 4693 1213
rect 4895 1199 4909 1213
rect 5591 1199 5605 1213
rect 5735 1199 5749 1213
rect 5975 1199 5989 1213
rect 6791 1199 6805 1213
rect 7055 1199 7069 1213
rect 191 1177 205 1191
rect 1631 1177 1645 1191
rect 2639 1177 2653 1191
rect 2759 1177 2773 1191
rect 2879 1177 2893 1191
rect 2999 1177 3013 1191
rect 4823 1177 4837 1191
rect 5567 1177 5581 1191
rect 5711 1177 5725 1191
rect 6767 1177 6781 1191
rect 6911 1177 6925 1191
rect 7031 1177 7045 1191
rect 239 358 253 372
rect 911 358 925 372
rect 1415 358 1429 372
rect 5327 358 5341 372
rect 5951 358 5965 372
rect 359 336 373 350
rect 2903 336 2917 350
rect 3023 336 3037 350
rect 5039 336 5053 350
rect 479 314 493 328
rect 815 314 829 328
rect 1031 314 1045 328
rect 1223 314 1237 328
rect 1679 314 1693 328
rect 2807 314 2821 328
rect 3047 314 3061 328
rect 5351 315 5365 329
rect 5999 314 6013 328
rect 599 292 613 306
rect 3143 292 3157 306
rect 3575 292 3589 306
rect 3719 292 3733 306
rect 3863 292 3877 306
rect 4007 292 4021 306
rect 5063 292 5077 306
rect 5783 292 5797 306
rect 6119 292 6133 306
rect 6815 292 6829 306
rect 6959 292 6973 306
rect 719 270 733 284
rect 839 270 853 284
rect 3455 269 3469 283
rect 3599 270 3613 284
rect 4031 270 4045 284
rect 4583 270 4597 284
rect 4727 270 4741 284
rect 5087 270 5101 284
rect 6143 270 6157 284
rect 6839 270 6853 284
rect 7295 270 7309 284
rect 7727 270 7741 284
rect 335 248 349 262
rect 1583 248 1597 262
rect 1919 248 1933 262
rect 2279 248 2293 262
rect 4487 248 4501 262
rect 5471 248 5485 262
rect 5519 248 5533 262
rect 5879 248 5893 262
rect 7247 248 7261 262
rect 7319 248 7333 262
rect 1727 226 1741 240
rect 1799 226 1813 240
rect 3335 226 3349 240
rect 5447 226 5461 240
rect 5495 226 5509 240
rect 6359 226 6373 240
rect 503 204 517 218
rect 2015 204 2029 218
rect 4631 204 4645 218
rect 7487 204 7501 218
rect 671 182 685 196
rect 2087 182 2101 196
rect 4343 175 4357 189
rect 5520 175 5534 189
rect 6143 182 6157 196
rect 6479 182 6493 196
rect 6719 182 6733 196
rect 6959 182 6973 196
rect 695 160 709 174
rect 2303 160 2317 174
rect 767 138 781 152
rect 2471 138 2485 152
rect 983 116 997 130
rect 2519 116 2533 130
rect 71 94 85 108
rect 3215 94 3229 108
rect 1463 68 1477 82
rect 3359 68 3373 82
rect 1823 46 1837 60
rect 3503 47 3517 61
rect 2231 19 2245 33
rect 3647 19 3661 33
rect 2567 -6 2581 8
rect 3791 -5 3805 9
rect 2879 -28 2893 -14
rect 3935 -28 3949 -14
rect 3215 -50 3229 -36
rect 4079 -50 4093 -36
rect 3383 -72 3397 -58
rect 4223 -71 4237 -57
rect 3551 -94 3565 -80
rect 5399 -94 5413 -80
rect 1127 -116 1141 -102
rect 4847 -116 4861 -102
<< metal2 >>
rect 192 1191 204 1659
rect 312 1213 324 1659
rect 432 1235 444 1659
rect 552 1257 564 1659
rect 672 1279 684 1659
rect 192 1174 204 1177
rect 312 1174 324 1199
rect 432 1174 444 1221
rect 552 1174 564 1243
rect 672 1174 684 1265
rect 792 1174 804 1199
rect 864 1174 876 1287
rect 936 1174 948 1221
rect 960 1174 972 1265
rect 984 1174 996 1309
rect 1056 1174 1068 1265
rect 1080 1174 1092 1331
rect 1128 1174 1140 1287
rect 1152 1174 1164 1309
rect 1176 1174 1188 1288
rect 1248 1174 1260 1331
rect 1272 1174 1284 1309
rect 1320 1174 1332 1287
rect 1344 1174 1356 1243
rect 1368 1174 1380 1287
rect 1440 1174 1452 1199
rect 1464 1174 1476 1309
rect 1488 1174 1500 1309
rect 1536 1174 1548 1287
rect 1560 1174 1572 1309
rect 1632 1174 1644 1177
rect 1656 1174 1668 1243
rect 1776 1174 1788 1659
rect 1848 1174 1860 1287
rect 1896 1174 1908 1287
rect 2112 1174 2124 1287
rect 2208 1174 2220 1659
rect 2400 1301 2412 1659
rect 2400 1174 2412 1287
rect 2472 1174 2484 1659
rect 2568 1174 2580 1659
rect 2640 1174 2652 1177
rect 2664 1174 2676 1199
rect 2688 1174 2700 1221
rect 2712 1174 2724 1287
rect 2760 1174 2772 1177
rect 2784 1174 2796 1199
rect 2832 1174 2844 1309
rect 2880 1174 2892 1177
rect 2928 1174 2940 1221
rect 2952 1174 2964 1331
rect 3000 1174 3012 1177
rect 3072 1174 3084 1353
rect 3120 1174 3132 1309
rect 3168 1174 3180 1265
rect 3264 1174 3276 1353
rect 3288 1174 3300 1243
rect 3312 1174 3324 1265
rect 3408 1174 3420 1353
rect 3432 1174 3444 1243
rect 3552 1174 3564 1353
rect 3696 1174 3708 1353
rect 3744 1174 3756 1265
rect 3840 1174 3852 1331
rect 3888 1174 3900 1265
rect 3984 1174 3996 1331
rect 4128 1174 4140 1331
rect 4152 1174 4164 1243
rect 4176 1174 4188 1265
rect 4272 1173 4284 1287
rect 4296 1174 4308 1243
rect 4392 1174 4404 1287
rect 4416 1174 4428 1243
rect 4440 1174 4452 1266
rect 4536 1174 4548 1331
rect 4560 1174 4572 1243
rect 4680 1174 4692 1199
rect 4704 1174 4716 1243
rect 4752 1174 4764 1287
rect 4800 1174 4812 1287
rect 4824 1174 4836 1177
rect 4896 1174 4908 1199
rect 4920 1174 4932 1243
rect 4944 1174 4956 1264
rect 4992 1174 5004 1309
rect 5136 1174 5148 1287
rect 5184 1174 5196 1287
rect 5208 1174 5220 1309
rect 5256 1174 5268 1287
rect 5304 1174 5316 1287
rect 5568 1174 5580 1177
rect 5592 1174 5604 1199
rect 5616 1174 5628 1221
rect 5640 1174 5652 1265
rect 5664 1174 5676 1309
rect 5712 1174 5724 1177
rect 5736 1174 5748 1199
rect 5760 1174 5772 1221
rect 5808 1174 5820 1287
rect 5856 1174 5868 1287
rect 5880 1174 5892 1309
rect 5904 1174 5916 1309
rect 5976 1174 5988 1199
rect 6048 1174 6060 1287
rect 6096 1174 6108 1287
rect 6168 1174 6180 1332
rect 6216 1174 6228 1309
rect 6240 1174 6252 1659
rect 6264 1174 6276 1287
rect 6312 1174 6324 1287
rect 6336 1174 6348 1332
rect 6408 1174 6420 1309
rect 6432 1174 6444 1659
rect 6528 1174 6540 1309
rect 6552 1174 6564 1659
rect 6648 1174 6660 1309
rect 6672 1174 6684 1659
rect 6768 1174 6780 1177
rect 6792 1174 6804 1199
rect 6864 1174 6876 1331
rect 6912 1174 6924 1177
rect 6936 1174 6948 1221
rect 6984 1174 6996 1309
rect 7032 1174 7044 1177
rect 7056 1174 7068 1199
rect 7080 1174 7092 1221
rect 7104 1174 7116 1265
rect 7128 1174 7140 1287
rect 7176 1174 7188 1287
rect 7200 1174 7212 1309
rect 7224 1174 7236 1331
rect 7296 1174 7308 1659
rect 240 372 252 375
rect 360 350 372 375
rect 480 328 492 375
rect 600 306 612 375
rect 720 284 732 375
rect 816 328 828 375
rect 840 284 852 375
rect 912 372 924 375
rect 1032 328 1044 375
rect 1224 328 1236 375
rect 1416 372 1428 375
rect 1584 262 1596 375
rect 1680 328 1692 375
rect 72 -200 84 94
rect 336 -200 348 248
rect 1728 240 1740 375
rect 1800 240 1812 375
rect 1920 262 1932 375
rect 2016 218 2028 375
rect 504 -200 516 204
rect 2088 196 2100 375
rect 2280 262 2292 375
rect 672 -200 684 182
rect 2304 174 2316 375
rect 696 -200 708 160
rect 2472 152 2484 375
rect 768 -200 780 138
rect 2520 130 2532 375
rect 2808 328 2820 375
rect 2904 350 2916 375
rect 3024 350 3036 375
rect 3048 328 3060 375
rect 3144 306 3156 375
rect 984 -200 996 116
rect 3216 108 3228 375
rect 1128 -200 1140 -116
rect 1464 -200 1476 68
rect 1824 -200 1836 46
rect 2232 -200 2244 19
rect 2568 -200 2580 -6
rect 2880 -200 2892 -28
rect 3216 -200 3228 -50
rect 3336 -200 3348 226
rect 3360 82 3372 375
rect 3456 283 3468 375
rect 3504 61 3516 375
rect 3576 306 3588 375
rect 3600 284 3612 375
rect 3648 33 3660 375
rect 3720 306 3732 375
rect 3792 9 3804 375
rect 3864 306 3876 375
rect 3936 -14 3948 375
rect 4008 306 4020 375
rect 4032 284 4044 375
rect 4080 -36 4092 375
rect 4224 -57 4236 375
rect 4344 189 4356 375
rect 4488 262 4500 375
rect 4584 284 4596 375
rect 4632 218 4644 375
rect 4728 284 4740 375
rect 3384 -200 3396 -72
rect 3552 -200 3564 -94
rect 4848 -102 4860 375
rect 5040 350 5052 375
rect 5064 306 5076 375
rect 5088 284 5100 375
rect 5328 372 5340 375
rect 5352 329 5364 375
rect 5400 -80 5412 375
rect 5448 240 5460 375
rect 5472 262 5484 375
rect 5520 262 5532 375
rect 5784 306 5796 375
rect 5952 372 5964 375
rect 6000 328 6012 375
rect 6120 306 6132 375
rect 6144 284 6156 375
rect 5496 -200 5508 226
rect 5521 -200 5533 175
rect 5880 -200 5892 248
rect 6360 240 6372 375
rect 6480 196 6492 375
rect 6144 -200 6156 182
rect 6600 -200 6612 375
rect 6720 196 6732 375
rect 6816 306 6828 375
rect 6840 284 6852 375
rect 6960 306 6972 375
rect 7248 262 7260 375
rect 7296 284 7308 375
rect 6960 -200 6972 182
rect 7320 -200 7332 248
rect 7488 -200 7500 204
rect 7728 -200 7740 270
use inv inv_0
timestamp 1386238110
transform 1 0 168 0 1 375
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 288 0 1 375
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 408 0 1 375
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 528 0 1 375
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 648 0 1 375
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 768 0 1 375
box 0 0 120 799
use nand3 nand3_1
timestamp 1386234893
transform 1 0 888 0 1 375
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 1008 0 1 375
box 0 0 96 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1104 0 1 375
box 0 0 96 799
use nand2 nand2_16
timestamp 1386234792
transform 1 0 1200 0 1 375
box 0 0 96 799
use nand2 nand2_17
timestamp 1386234792
transform 1 0 1296 0 1 375
box 0 0 96 799
use nand3 nand3_2
timestamp 1386234893
transform 1 0 1392 0 1 375
box 0 0 120 799
use nand2 nand2_18
timestamp 1386234792
transform 1 0 1512 0 1 375
box 0 0 96 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 1608 0 1 375
box 0 0 144 799
use and2 and2_4
timestamp 1386234845
transform 1 0 1752 0 1 375
box 0 0 120 799
use xor2 xor2_3
timestamp 1386237344
transform 1 0 1872 0 1 375
box 0 0 192 799
use xor2 xor2_4
timestamp 1386237344
transform 1 0 2064 0 1 375
box 0 0 192 799
use xor2 xor2_5
timestamp 1386237344
transform 1 0 2256 0 1 375
box 0 0 192 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 2448 0 1 375
box 0 0 48 799
use inv inv_6
timestamp 1386238110
transform 1 0 2496 0 1 375
box 0 0 120 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 2616 0 1 375
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 2736 0 1 375
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 2856 0 1 375
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 2976 0 1 375
box 0 0 120 799
use nor3 nor3_6
timestamp 1386235396
transform 1 0 3096 0 1 375
box 0 0 144 799
use nor3 nor3_7
timestamp 1386235396
transform 1 0 3240 0 1 375
box 0 0 144 799
use nor3 nor3_8
timestamp 1386235396
transform 1 0 3384 0 1 375
box 0 0 144 799
use nor3 nor3_9
timestamp 1386235396
transform 1 0 3528 0 1 375
box 0 0 144 799
use nor3 nor3_10
timestamp 1386235396
transform 1 0 3672 0 1 375
box 0 0 144 799
use nor3 nor3_11
timestamp 1386235396
transform 1 0 3816 0 1 375
box 0 0 144 799
use nor3 nor3_12
timestamp 1386235396
transform 1 0 3960 0 1 375
box 0 0 144 799
use nor3 nor3_13
timestamp 1386235396
transform 1 0 4104 0 1 375
box 0 0 144 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 4248 0 1 375
box 0 0 120 799
use nor3 nor3_15
timestamp 1386235396
transform 1 0 4368 0 1 375
box 0 0 144 799
use nor3 nor3_16
timestamp 1386235396
transform 1 0 4512 0 1 375
box 0 0 144 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 4656 0 1 375
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 4776 0 1 375
box 0 0 96 799
use nor3 nor3_2
timestamp 1386235396
transform 1 0 4872 0 1 375
box 0 0 144 799
use nor3 nor3_3
timestamp 1386235396
transform 1 0 5016 0 1 375
box 0 0 144 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 5160 0 1 375
box 0 0 120 799
use nor3 nor3_4
timestamp 1386235396
transform 1 0 5280 0 1 375
box 0 0 144 799
use and2 and2_3
timestamp 1386234845
transform 1 0 5424 0 1 375
box 0 0 120 799
use nand4 nand4_2
timestamp 1386234936
transform 1 0 5544 0 1 375
box 0 0 144 799
use nand4 nand4_3
timestamp 1386234936
transform 1 0 5688 0 1 375
box 0 0 144 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 5832 0 1 375
box 0 0 96 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 5928 0 1 375
box 0 0 144 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 6072 0 1 375
box 0 0 120 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 6192 0 1 375
box 0 0 96 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 6288 0 1 375
box 0 0 96 799
use and2 and2_0
timestamp 1386234845
transform 1 0 6384 0 1 375
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 6504 0 1 375
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 6624 0 1 375
box 0 0 120 799
use nand4 nand4_4
timestamp 1386234936
transform 1 0 6744 0 1 375
box 0 0 144 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 6888 0 1 375
box 0 0 120 799
use nand4 nand4_5
timestamp 1386234936
transform 1 0 7008 0 1 375
box 0 0 144 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 7152 0 1 375
box 0 0 120 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 7272 0 1 375
box 0 0 48 799
<< labels >>
rlabel metal1 504 322 504 322 1 nC
rlabel metal1 272 364 272 364 1 nA
rlabel metal1 378 342 378 342 1 nB
rlabel metal1 627 297 627 297 1 nD
rlabel metal1 0 1096 0 1121 3 Vdd!
rlabel metal1 0 451 0 476 3 GND!
rlabel metal2 2880 -200 2892 -200 1 NAND
rlabel metal2 336 -200 348 -200 1 SUB
rlabel metal2 504 -200 516 -200 1 CIn_slice
rlabel metal2 672 -200 684 -200 1 LastCIn
rlabel metal2 696 -200 708 -200 1 COut
rlabel metal2 984 -200 996 -200 1 nZ
rlabel metal2 1128 -200 1140 -200 1 FAOut
rlabel metal2 1464 -200 1476 -200 1 AND
rlabel metal2 1824 -200 1836 -200 1 OR
rlabel metal2 2232 -200 2244 -200 1 XOR
rlabel metal2 2568 -200 2580 -200 1 NOT
rlabel metal2 3552 -200 3564 -200 1 ShL
rlabel metal2 3336 -200 3348 -200 1 ASign
rlabel metal2 3384 -200 3396 -200 1 ShB
rlabel metal2 3216 -200 3228 -200 1 NOR
rlabel metal2 768 -200 780 -200 1 N
rlabel metal2 72 -200 84 -200 1 ZeroA
rlabel metal2 192 1659 204 1659 5 OpCode[4]
rlabel metal2 312 1659 324 1659 5 OpCode[3]
rlabel metal2 432 1659 444 1659 5 OpCode[2]
rlabel metal2 552 1659 564 1659 5 OpCode[1]
rlabel metal2 672 1659 684 1659 5 OpCode[0]
rlabel metal1 747 275 747 275 1 nE
rlabel metal1 1765 232 1765 232 1 UseC
rlabel metal2 2568 1659 2580 1659 5 Z
rlabel metal2 2472 1659 2484 1659 5 N
rlabel metal2 2208 1659 2220 1659 5 V
rlabel metal2 1776 1659 1788 1659 5 Cin
rlabel metal2 2400 1659 2412 1659 5 C
rlabel metal1 3101 1291 3101 1291 1 ABC
rlabel metal1 3096 1314 3096 1314 1 ABnC
rlabel metal1 3095 1337 3095 1337 1 AnBC
rlabel metal1 3096 1359 3096 1359 1 AnBnC
rlabel metal1 0 428 0 438 1 Clock
rlabel metal1 0 405 0 415 1 Test
rlabel metal1 0 382 0 392 1 nReset
rlabel metal1 0 1134 0 1144 3 Scan
rlabel metal1 0 1157 0 1167 3 ScanReturn
rlabel metal2 5880 -200 5892 -200 1 ShInBit
rlabel metal2 5496 -200 5508 -200 1 Sh8
rlabel metal2 6144 -200 6156 -200 1 Sh4
rlabel metal2 6960 -200 6972 -200 1 Sh1
rlabel metal2 5521 -200 5533 -200 1 ShR
rlabel metal2 6600 -200 6612 -200 1 Sh2
rlabel metal2 7320 -200 7332 -200 1 ShOut
rlabel metal2 7488 -200 7500 -200 1 LLI
rlabel metal2 7728 -200 7740 -200 1 OutEn
rlabel metal2 5911 1194 5911 1194 1 N
rlabel metal1 7822 1096 7822 1121 7 Vdd!
rlabel metal1 7822 451 7822 476 7 GND!
rlabel metal1 5418 254 5418 254 1 ShSign
rlabel metal2 6240 1659 6252 1659 5 imm4[3]
rlabel metal2 6672 1659 6684 1659 5 imm4[0]
rlabel metal2 6552 1659 6564 1659 5 imm4[1]
rlabel metal2 6432 1659 6444 1659 5 imm4[2]
rlabel metal2 7296 1659 7308 1659 5 OutEn
rlabel metal1 7822 1134 7822 1144 1 Scan
rlabel metal1 7822 1157 7822 1167 1 ScanReturn
rlabel metal1 7822 428 7822 438 7 Clock
rlabel metal1 7822 382 7822 392 7 nReset
rlabel metal1 7822 405 7822 415 7 Test
<< end >>
