magic
tech c035u
timestamp 1394829379
<< metal1 >>
rect 0 15600 58 15610
rect 48 15397 58 15600
rect 0 15360 82 15370
rect 48 15157 58 15335
rect 72 15157 82 15360
rect 0 15120 106 15130
rect 48 14917 58 15095
rect 72 14917 82 15095
rect 96 14917 106 15120
rect 0 14880 130 14890
rect 48 14677 58 14855
rect 72 14677 82 14855
rect 96 14677 106 14855
rect 120 14677 130 14880
rect 0 14640 154 14650
rect 48 14437 58 14615
rect 72 14437 82 14615
rect 96 14437 106 14615
rect 120 14437 130 14615
rect 144 14437 154 14640
rect 0 14400 178 14410
rect 48 14197 58 14375
rect 72 14197 82 14375
rect 96 14197 106 14375
rect 120 14197 130 14375
rect 144 14197 154 14375
rect 168 14197 178 14400
rect 0 14160 202 14170
rect 48 13957 58 14135
rect 72 13957 82 14135
rect 96 13957 106 14135
rect 120 13957 130 14135
rect 144 13957 154 14135
rect 168 13957 178 14135
rect 192 13957 202 14160
rect 0 13920 226 13930
rect 48 13717 58 13895
rect 72 13717 82 13895
rect 96 13717 106 13895
rect 120 13717 130 13895
rect 144 13717 154 13895
rect 168 13717 178 13895
rect 192 13717 202 13895
rect 216 13717 226 13920
rect 0 13680 250 13690
rect 48 13477 58 13655
rect 72 13477 82 13655
rect 96 13477 106 13655
rect 120 13477 130 13655
rect 144 13477 154 13655
rect 168 13477 178 13655
rect 192 13477 202 13655
rect 216 13477 226 13655
rect 240 13477 250 13680
rect 0 13440 274 13450
rect 48 13237 58 13415
rect 72 13237 82 13415
rect 96 13237 106 13415
rect 120 13237 130 13415
rect 144 13237 154 13415
rect 168 13237 178 13415
rect 192 13237 202 13415
rect 216 13237 226 13415
rect 240 13237 250 13415
rect 264 13237 274 13440
rect 0 13200 298 13210
rect 48 12997 58 13175
rect 72 12997 82 13175
rect 96 12997 106 13175
rect 120 12997 130 13175
rect 144 12997 154 13175
rect 168 12997 178 13175
rect 192 12997 202 13175
rect 216 12997 226 13175
rect 240 12997 250 13175
rect 264 12997 274 13175
rect 288 12997 298 13200
rect 0 12960 322 12970
rect 48 12757 58 12935
rect 72 12757 82 12935
rect 96 12757 106 12935
rect 120 12757 130 12935
rect 144 12757 154 12935
rect 168 12757 178 12935
rect 192 12757 202 12935
rect 216 12757 226 12935
rect 240 12757 250 12935
rect 264 12757 274 12935
rect 288 12757 298 12935
rect 312 12757 322 12960
rect 0 12720 346 12730
rect 48 12517 58 12695
rect 72 12517 82 12695
rect 96 12517 106 12695
rect 120 12517 130 12695
rect 144 12517 154 12695
rect 168 12517 178 12695
rect 192 12517 202 12695
rect 216 12517 226 12695
rect 240 12517 250 12695
rect 264 12517 274 12695
rect 288 12517 298 12695
rect 312 12517 322 12695
rect 336 12517 346 12720
rect 0 12480 370 12490
rect 48 12277 58 12455
rect 72 12277 82 12455
rect 96 12277 106 12455
rect 120 12277 130 12455
rect 144 12277 154 12455
rect 168 12277 178 12455
rect 192 12277 202 12455
rect 216 12277 226 12455
rect 240 12277 250 12455
rect 264 12277 274 12455
rect 288 12277 298 12455
rect 312 12277 322 12455
rect 336 12277 346 12455
rect 360 12277 370 12480
rect 0 12240 394 12250
rect 48 12037 58 12215
rect 72 12037 82 12215
rect 96 12037 106 12215
rect 120 12037 130 12215
rect 144 12037 154 12215
rect 168 12037 178 12215
rect 192 12037 202 12215
rect 216 12037 226 12215
rect 240 12037 250 12215
rect 264 12037 274 12215
rect 288 12037 298 12215
rect 312 12037 322 12215
rect 336 12037 346 12215
rect 360 12037 370 12215
rect 384 12037 394 12240
rect 0 12000 418 12010
rect 48 11797 58 11975
rect 72 11797 82 11975
rect 96 11797 106 11975
rect 120 11797 130 11975
rect 144 11797 154 11975
rect 168 11797 178 11975
rect 192 11797 202 11975
rect 216 11797 226 11975
rect 240 11797 250 11975
rect 264 11797 274 11975
rect 288 11797 298 11975
rect 312 11797 322 11975
rect 336 11797 346 11975
rect 360 11797 370 11975
rect 384 11797 394 11975
rect 408 11797 418 12000
rect 0 11760 442 11770
rect 48 11557 58 11735
rect 72 11557 82 11735
rect 96 11557 106 11735
rect 120 11557 130 11735
rect 144 11557 154 11735
rect 168 11557 178 11735
rect 192 11557 202 11735
rect 216 11557 226 11735
rect 240 11557 250 11735
rect 264 11557 274 11735
rect 288 11557 298 11735
rect 312 11557 322 11735
rect 336 11557 346 11735
rect 360 11557 370 11735
rect 384 11557 394 11735
rect 408 11557 418 11735
rect 432 11557 442 11760
rect 0 11520 466 11530
rect 48 11317 58 11495
rect 72 11317 82 11495
rect 96 11317 106 11495
rect 120 11317 130 11495
rect 144 11317 154 11495
rect 168 11317 178 11495
rect 192 11317 202 11495
rect 216 11317 226 11495
rect 240 11317 250 11495
rect 264 11317 274 11495
rect 288 11317 298 11495
rect 312 11317 322 11495
rect 336 11317 346 11495
rect 360 11317 370 11495
rect 384 11317 394 11495
rect 408 11317 418 11495
rect 432 11317 442 11495
rect 456 11317 466 11520
rect 0 11280 490 11290
rect 48 11077 58 11255
rect 72 11077 82 11255
rect 96 11077 106 11255
rect 120 11077 130 11255
rect 144 11077 154 11255
rect 168 11077 178 11255
rect 192 11077 202 11255
rect 216 11077 226 11255
rect 240 11077 250 11255
rect 264 11077 274 11255
rect 288 11077 298 11255
rect 312 11077 322 11255
rect 336 11077 346 11255
rect 360 11077 370 11255
rect 384 11077 394 11255
rect 408 11077 418 11255
rect 432 11077 442 11255
rect 456 11077 466 11255
rect 480 11077 490 11280
rect 0 11040 514 11050
rect 48 10837 58 11015
rect 72 10837 82 11015
rect 96 10837 106 11015
rect 120 10837 130 11015
rect 144 10837 154 11015
rect 168 10837 178 11015
rect 192 10837 202 11015
rect 216 10837 226 11015
rect 240 10837 250 11015
rect 264 10837 274 11015
rect 288 10837 298 11015
rect 312 10837 322 11015
rect 336 10837 346 11015
rect 360 10837 370 11015
rect 384 10837 394 11015
rect 408 10837 418 11015
rect 432 10837 442 11015
rect 456 10837 466 11015
rect 480 10837 490 11015
rect 504 10837 514 11040
rect 0 10800 538 10810
rect 48 10597 58 10775
rect 72 10597 82 10775
rect 96 10597 106 10775
rect 120 10597 130 10775
rect 144 10597 154 10775
rect 168 10597 178 10775
rect 192 10597 202 10775
rect 216 10597 226 10775
rect 240 10597 250 10775
rect 264 10597 274 10775
rect 288 10597 298 10775
rect 312 10597 322 10775
rect 336 10597 346 10775
rect 360 10597 370 10775
rect 384 10597 394 10775
rect 408 10597 418 10775
rect 432 10597 442 10775
rect 456 10597 466 10775
rect 480 10597 490 10775
rect 504 10597 514 10775
rect 528 10597 538 10800
rect 0 10560 562 10570
rect 48 10357 58 10535
rect 72 10357 82 10535
rect 96 10357 106 10535
rect 120 10357 130 10535
rect 144 10357 154 10535
rect 168 10357 178 10535
rect 192 10357 202 10535
rect 216 10357 226 10535
rect 240 10357 250 10535
rect 264 10357 274 10535
rect 288 10357 298 10535
rect 312 10357 322 10535
rect 336 10357 346 10535
rect 360 10357 370 10535
rect 384 10357 394 10535
rect 408 10357 418 10535
rect 432 10357 442 10535
rect 456 10357 466 10535
rect 480 10357 490 10535
rect 504 10357 514 10535
rect 528 10357 538 10535
rect 552 10357 562 10560
rect 0 10320 586 10330
rect 48 10117 58 10295
rect 72 10117 82 10295
rect 96 10117 106 10295
rect 120 10117 130 10295
rect 144 10117 154 10295
rect 168 10117 178 10295
rect 192 10117 202 10295
rect 216 10117 226 10295
rect 240 10117 250 10295
rect 264 10117 274 10295
rect 288 10117 298 10295
rect 312 10117 322 10295
rect 336 10117 346 10295
rect 360 10117 370 10295
rect 384 10117 394 10295
rect 408 10117 418 10295
rect 432 10117 442 10295
rect 456 10117 466 10295
rect 480 10117 490 10295
rect 504 10117 514 10295
rect 528 10117 538 10295
rect 552 10117 562 10295
rect 576 10117 586 10320
rect 0 10080 610 10090
rect 48 9877 58 10055
rect 72 9877 82 10055
rect 96 9877 106 10055
rect 120 9877 130 10055
rect 144 9877 154 10055
rect 168 9877 178 10055
rect 192 9877 202 10055
rect 216 9877 226 10055
rect 240 9877 250 10055
rect 264 9877 274 10055
rect 288 9877 298 10055
rect 312 9877 322 10055
rect 336 9877 346 10055
rect 360 9877 370 10055
rect 384 9877 394 10055
rect 408 9877 418 10055
rect 432 9877 442 10055
rect 456 9877 466 10055
rect 480 9877 490 10055
rect 504 9877 514 10055
rect 528 9877 538 10055
rect 552 9877 562 10055
rect 576 9877 586 10055
rect 600 9877 610 10080
rect 0 9840 634 9850
rect 48 9637 58 9815
rect 72 9637 82 9815
rect 96 9637 106 9815
rect 120 9637 130 9815
rect 144 9637 154 9815
rect 168 9637 178 9815
rect 192 9637 202 9815
rect 216 9637 226 9815
rect 240 9637 250 9815
rect 264 9637 274 9815
rect 288 9637 298 9815
rect 312 9637 322 9815
rect 336 9637 346 9815
rect 360 9637 370 9815
rect 384 9637 394 9815
rect 408 9637 418 9815
rect 432 9637 442 9815
rect 456 9637 466 9815
rect 480 9637 490 9815
rect 504 9637 514 9815
rect 528 9637 538 9815
rect 552 9637 562 9815
rect 576 9637 586 9815
rect 600 9637 610 9815
rect 624 9637 634 9840
rect 0 9600 658 9610
rect 48 9397 58 9575
rect 72 9397 82 9575
rect 96 9397 106 9575
rect 120 9397 130 9575
rect 144 9397 154 9575
rect 168 9397 178 9575
rect 192 9397 202 9575
rect 216 9397 226 9575
rect 240 9397 250 9575
rect 264 9397 274 9575
rect 288 9397 298 9575
rect 312 9397 322 9575
rect 336 9397 346 9575
rect 360 9397 370 9575
rect 384 9397 394 9575
rect 408 9397 418 9575
rect 432 9397 442 9575
rect 456 9397 466 9575
rect 480 9397 490 9575
rect 504 9397 514 9575
rect 528 9397 538 9575
rect 552 9397 562 9575
rect 576 9397 586 9575
rect 600 9397 610 9575
rect 624 9397 634 9575
rect 648 9397 658 9600
rect 0 9360 682 9370
rect 48 9157 58 9335
rect 72 9157 82 9335
rect 96 9157 106 9335
rect 120 9157 130 9335
rect 144 9157 154 9335
rect 168 9157 178 9335
rect 192 9157 202 9335
rect 216 9157 226 9335
rect 240 9157 250 9335
rect 264 9157 274 9335
rect 288 9157 298 9335
rect 312 9157 322 9335
rect 336 9157 346 9335
rect 360 9157 370 9335
rect 384 9157 394 9335
rect 408 9157 418 9335
rect 432 9157 442 9335
rect 456 9157 466 9335
rect 480 9157 490 9335
rect 504 9157 514 9335
rect 528 9157 538 9335
rect 552 9157 562 9335
rect 576 9157 586 9335
rect 600 9157 610 9335
rect 624 9157 634 9335
rect 648 9157 658 9335
rect 672 9157 682 9360
rect 0 9120 706 9130
rect 48 8917 58 9095
rect 72 8917 82 9095
rect 96 8917 106 9095
rect 120 8917 130 9095
rect 144 8917 154 9095
rect 168 8917 178 9095
rect 192 8917 202 9095
rect 216 8917 226 9095
rect 240 8917 250 9095
rect 264 8917 274 9095
rect 288 8917 298 9095
rect 312 8917 322 9095
rect 336 8917 346 9095
rect 360 8917 370 9095
rect 384 8917 394 9095
rect 408 8917 418 9095
rect 432 8917 442 9095
rect 456 8917 466 9095
rect 480 8917 490 9095
rect 504 8917 514 9095
rect 528 8917 538 9095
rect 552 8917 562 9095
rect 576 8917 586 9095
rect 600 8917 610 9095
rect 624 8917 634 9095
rect 648 8917 658 9095
rect 672 8917 682 9095
rect 696 8917 706 9120
rect 0 8880 730 8890
rect 48 8677 58 8855
rect 72 8677 82 8855
rect 96 8677 106 8855
rect 120 8677 130 8855
rect 144 8677 154 8855
rect 168 8677 178 8855
rect 192 8677 202 8855
rect 216 8677 226 8855
rect 240 8677 250 8855
rect 264 8677 274 8855
rect 288 8677 298 8855
rect 312 8677 322 8855
rect 336 8677 346 8855
rect 360 8677 370 8855
rect 384 8677 394 8855
rect 408 8677 418 8855
rect 432 8677 442 8855
rect 456 8677 466 8855
rect 480 8677 490 8855
rect 504 8677 514 8855
rect 528 8677 538 8855
rect 552 8677 562 8855
rect 576 8677 586 8855
rect 600 8677 610 8855
rect 624 8677 634 8855
rect 648 8677 658 8855
rect 672 8677 682 8855
rect 696 8677 706 8855
rect 720 8677 730 8880
rect 0 8640 754 8650
rect 48 8437 58 8615
rect 72 8437 82 8615
rect 96 8437 106 8615
rect 120 8437 130 8615
rect 144 8437 154 8615
rect 168 8437 178 8615
rect 192 8437 202 8615
rect 216 8437 226 8615
rect 240 8437 250 8615
rect 264 8437 274 8615
rect 288 8437 298 8615
rect 312 8437 322 8615
rect 336 8437 346 8615
rect 360 8437 370 8615
rect 384 8437 394 8615
rect 408 8437 418 8615
rect 432 8437 442 8615
rect 456 8437 466 8615
rect 480 8437 490 8615
rect 504 8437 514 8615
rect 528 8437 538 8615
rect 552 8437 562 8615
rect 576 8437 586 8615
rect 600 8437 610 8615
rect 624 8437 634 8615
rect 648 8437 658 8615
rect 672 8437 682 8615
rect 696 8437 706 8615
rect 720 8437 730 8615
rect 744 8437 754 8640
rect 0 8400 778 8410
rect 48 8197 58 8375
rect 72 8197 82 8375
rect 96 8197 106 8375
rect 120 8197 130 8375
rect 144 8197 154 8375
rect 168 8197 178 8375
rect 192 8197 202 8375
rect 216 8197 226 8375
rect 240 8197 250 8375
rect 264 8197 274 8375
rect 288 8197 298 8375
rect 312 8197 322 8375
rect 336 8197 346 8375
rect 360 8197 370 8375
rect 384 8197 394 8375
rect 408 8197 418 8375
rect 432 8197 442 8375
rect 456 8197 466 8375
rect 480 8197 490 8375
rect 504 8197 514 8375
rect 528 8197 538 8375
rect 552 8197 562 8375
rect 576 8197 586 8375
rect 600 8197 610 8375
rect 624 8197 634 8375
rect 648 8197 658 8375
rect 672 8197 682 8375
rect 696 8197 706 8375
rect 720 8197 730 8375
rect 744 8197 754 8375
rect 768 8197 778 8400
rect 0 8160 802 8170
rect 48 7957 58 8135
rect 72 7957 82 8135
rect 96 7957 106 8135
rect 120 7957 130 8135
rect 144 7957 154 8135
rect 168 7957 178 8135
rect 192 7957 202 8135
rect 216 7957 226 8135
rect 240 7957 250 8135
rect 264 7957 274 8135
rect 288 7957 298 8135
rect 312 7957 322 8135
rect 336 7957 346 8135
rect 360 7957 370 8135
rect 384 7957 394 8135
rect 408 7957 418 8135
rect 432 7957 442 8135
rect 456 7957 466 8135
rect 480 7957 490 8135
rect 504 7957 514 8135
rect 528 7957 538 8135
rect 552 7957 562 8135
rect 576 7957 586 8135
rect 600 7957 610 8135
rect 624 7957 634 8135
rect 648 7957 658 8135
rect 672 7957 682 8135
rect 696 7957 706 8135
rect 720 7957 730 8135
rect 744 7957 754 8135
rect 768 7957 778 8135
rect 792 7957 802 8160
rect 0 7920 826 7930
rect 48 7717 58 7895
rect 72 7717 82 7895
rect 96 7717 106 7895
rect 120 7717 130 7895
rect 144 7717 154 7895
rect 168 7717 178 7895
rect 192 7717 202 7895
rect 216 7717 226 7895
rect 240 7717 250 7895
rect 264 7717 274 7895
rect 288 7717 298 7895
rect 312 7717 322 7895
rect 336 7717 346 7895
rect 360 7717 370 7895
rect 384 7717 394 7895
rect 408 7717 418 7895
rect 432 7717 442 7895
rect 456 7717 466 7895
rect 480 7717 490 7895
rect 504 7717 514 7895
rect 528 7717 538 7895
rect 552 7717 562 7895
rect 576 7717 586 7895
rect 600 7717 610 7895
rect 624 7717 634 7895
rect 648 7717 658 7895
rect 672 7717 682 7895
rect 696 7717 706 7895
rect 720 7717 730 7895
rect 744 7717 754 7895
rect 768 7717 778 7895
rect 792 7717 802 7895
rect 816 7717 826 7920
rect 0 7680 850 7690
rect 48 7477 58 7655
rect 72 7477 82 7655
rect 96 7477 106 7655
rect 120 7477 130 7655
rect 144 7477 154 7655
rect 168 7477 178 7655
rect 192 7477 202 7655
rect 216 7477 226 7655
rect 240 7477 250 7655
rect 264 7477 274 7655
rect 288 7477 298 7655
rect 312 7477 322 7655
rect 336 7477 346 7655
rect 360 7477 370 7655
rect 384 7477 394 7655
rect 408 7477 418 7655
rect 432 7477 442 7655
rect 456 7477 466 7655
rect 480 7477 490 7655
rect 504 7477 514 7655
rect 528 7477 538 7655
rect 552 7477 562 7655
rect 576 7477 586 7655
rect 600 7477 610 7655
rect 624 7477 634 7655
rect 648 7477 658 7655
rect 672 7477 682 7655
rect 696 7477 706 7655
rect 720 7477 730 7655
rect 744 7477 754 7655
rect 768 7477 778 7655
rect 792 7477 802 7655
rect 816 7477 826 7655
rect 840 7477 850 7680
rect 0 7440 874 7450
rect 48 7237 58 7415
rect 72 7237 82 7415
rect 96 7237 106 7415
rect 120 7237 130 7415
rect 144 7237 154 7415
rect 168 7237 178 7415
rect 192 7237 202 7415
rect 216 7237 226 7415
rect 240 7237 250 7415
rect 264 7237 274 7415
rect 288 7237 298 7415
rect 312 7237 322 7415
rect 336 7237 346 7415
rect 360 7237 370 7415
rect 384 7237 394 7415
rect 408 7237 418 7415
rect 432 7237 442 7415
rect 456 7237 466 7415
rect 480 7237 490 7415
rect 504 7237 514 7415
rect 528 7237 538 7415
rect 552 7237 562 7415
rect 576 7237 586 7415
rect 600 7237 610 7415
rect 624 7237 634 7415
rect 648 7237 658 7415
rect 672 7237 682 7415
rect 696 7237 706 7415
rect 720 7237 730 7415
rect 744 7237 754 7415
rect 768 7237 778 7415
rect 792 7237 802 7415
rect 816 7237 826 7415
rect 840 7237 850 7415
rect 864 7237 874 7440
rect 0 7200 898 7210
rect 48 6997 58 7175
rect 72 6997 82 7175
rect 96 6997 106 7175
rect 120 6997 130 7175
rect 144 6997 154 7175
rect 168 6997 178 7175
rect 192 6997 202 7175
rect 216 6997 226 7175
rect 240 6997 250 7175
rect 264 6997 274 7175
rect 288 6997 298 7175
rect 312 6997 322 7175
rect 336 6997 346 7175
rect 360 6997 370 7175
rect 384 6997 394 7175
rect 408 6997 418 7175
rect 432 6997 442 7175
rect 456 6997 466 7175
rect 480 6997 490 7175
rect 504 6997 514 7175
rect 528 6997 538 7175
rect 552 6997 562 7175
rect 576 6997 586 7175
rect 600 6997 610 7175
rect 624 6997 634 7175
rect 648 6997 658 7175
rect 672 6997 682 7175
rect 696 6997 706 7175
rect 720 6997 730 7175
rect 744 6997 754 7175
rect 768 6997 778 7175
rect 792 6997 802 7175
rect 816 6997 826 7175
rect 840 6997 850 7175
rect 864 6997 874 7175
rect 888 6997 898 7200
rect 0 6960 922 6970
rect 48 6757 58 6935
rect 72 6757 82 6935
rect 96 6757 106 6935
rect 120 6757 130 6935
rect 144 6757 154 6935
rect 168 6757 178 6935
rect 192 6757 202 6935
rect 216 6757 226 6935
rect 240 6757 250 6935
rect 264 6757 274 6935
rect 288 6757 298 6935
rect 312 6757 322 6935
rect 336 6757 346 6935
rect 360 6757 370 6935
rect 384 6757 394 6935
rect 408 6757 418 6935
rect 432 6757 442 6935
rect 456 6757 466 6935
rect 480 6757 490 6935
rect 504 6757 514 6935
rect 528 6757 538 6935
rect 552 6757 562 6935
rect 576 6757 586 6935
rect 600 6757 610 6935
rect 624 6757 634 6935
rect 648 6757 658 6935
rect 672 6757 682 6935
rect 696 6757 706 6935
rect 720 6757 730 6935
rect 744 6757 754 6935
rect 768 6757 778 6935
rect 792 6757 802 6935
rect 816 6757 826 6935
rect 840 6757 850 6935
rect 864 6757 874 6935
rect 888 6757 898 6935
rect 912 6757 922 6960
rect 0 6720 946 6730
rect 48 6517 58 6695
rect 72 6517 82 6695
rect 96 6517 106 6695
rect 120 6517 130 6695
rect 144 6517 154 6695
rect 168 6517 178 6695
rect 192 6517 202 6695
rect 216 6517 226 6695
rect 240 6517 250 6695
rect 264 6517 274 6695
rect 288 6517 298 6695
rect 312 6517 322 6695
rect 336 6517 346 6695
rect 360 6517 370 6695
rect 384 6517 394 6695
rect 408 6517 418 6695
rect 432 6517 442 6695
rect 456 6517 466 6695
rect 480 6517 490 6695
rect 504 6517 514 6695
rect 528 6517 538 6695
rect 552 6517 562 6695
rect 576 6517 586 6695
rect 600 6517 610 6695
rect 624 6517 634 6695
rect 648 6517 658 6695
rect 672 6517 682 6695
rect 696 6517 706 6695
rect 720 6517 730 6695
rect 744 6517 754 6695
rect 768 6517 778 6695
rect 792 6517 802 6695
rect 816 6517 826 6695
rect 840 6517 850 6695
rect 864 6517 874 6695
rect 888 6517 898 6695
rect 912 6517 922 6695
rect 936 6517 946 6720
rect 0 6480 970 6490
rect 48 6277 58 6455
rect 72 6277 82 6455
rect 96 6277 106 6455
rect 120 6277 130 6455
rect 144 6277 154 6455
rect 168 6277 178 6455
rect 192 6277 202 6455
rect 216 6277 226 6455
rect 240 6277 250 6455
rect 264 6277 274 6455
rect 288 6277 298 6455
rect 312 6277 322 6455
rect 336 6277 346 6455
rect 360 6277 370 6455
rect 384 6277 394 6455
rect 408 6277 418 6455
rect 432 6277 442 6455
rect 456 6277 466 6455
rect 480 6277 490 6455
rect 504 6277 514 6455
rect 528 6277 538 6455
rect 552 6277 562 6455
rect 576 6277 586 6455
rect 600 6277 610 6455
rect 624 6277 634 6455
rect 648 6277 658 6455
rect 672 6277 682 6455
rect 696 6277 706 6455
rect 720 6277 730 6455
rect 744 6277 754 6455
rect 768 6277 778 6455
rect 792 6277 802 6455
rect 816 6277 826 6455
rect 840 6277 850 6455
rect 864 6277 874 6455
rect 888 6277 898 6455
rect 912 6277 922 6455
rect 936 6277 946 6455
rect 960 6277 970 6480
rect 0 6240 994 6250
rect 48 6037 58 6215
rect 72 6037 82 6215
rect 96 6037 106 6215
rect 120 6037 130 6215
rect 144 6037 154 6215
rect 168 6037 178 6215
rect 192 6037 202 6215
rect 216 6037 226 6215
rect 240 6037 250 6215
rect 264 6037 274 6215
rect 288 6037 298 6215
rect 312 6037 322 6215
rect 336 6037 346 6215
rect 360 6037 370 6215
rect 384 6037 394 6215
rect 408 6037 418 6215
rect 432 6037 442 6215
rect 456 6037 466 6215
rect 480 6037 490 6215
rect 504 6037 514 6215
rect 528 6037 538 6215
rect 552 6037 562 6215
rect 576 6037 586 6215
rect 600 6037 610 6215
rect 624 6037 634 6215
rect 648 6037 658 6215
rect 672 6037 682 6215
rect 696 6037 706 6215
rect 720 6037 730 6215
rect 744 6037 754 6215
rect 768 6037 778 6215
rect 792 6037 802 6215
rect 816 6037 826 6215
rect 840 6037 850 6215
rect 864 6037 874 6215
rect 888 6037 898 6215
rect 912 6037 922 6215
rect 936 6037 946 6215
rect 960 6037 970 6215
rect 984 6037 994 6240
rect 0 6000 1018 6010
rect 48 5797 58 5975
rect 72 5797 82 5975
rect 96 5797 106 5975
rect 120 5797 130 5975
rect 144 5797 154 5975
rect 168 5797 178 5975
rect 192 5797 202 5975
rect 216 5797 226 5975
rect 240 5797 250 5975
rect 264 5797 274 5975
rect 288 5797 298 5975
rect 312 5797 322 5975
rect 336 5797 346 5975
rect 360 5797 370 5975
rect 384 5797 394 5975
rect 408 5797 418 5975
rect 432 5797 442 5975
rect 456 5797 466 5975
rect 480 5797 490 5975
rect 504 5797 514 5975
rect 528 5797 538 5975
rect 552 5797 562 5975
rect 576 5797 586 5975
rect 600 5797 610 5975
rect 624 5797 634 5975
rect 648 5797 658 5975
rect 672 5797 682 5975
rect 696 5797 706 5975
rect 720 5797 730 5975
rect 744 5797 754 5975
rect 768 5797 778 5975
rect 792 5797 802 5975
rect 816 5797 826 5975
rect 840 5797 850 5975
rect 864 5797 874 5975
rect 888 5797 898 5975
rect 912 5797 922 5975
rect 936 5797 946 5975
rect 960 5797 970 5975
rect 984 5797 994 5975
rect 1008 5797 1018 6000
rect 0 5760 1042 5770
rect 48 5557 58 5735
rect 72 5557 82 5735
rect 96 5557 106 5735
rect 120 5557 130 5735
rect 144 5557 154 5735
rect 168 5557 178 5735
rect 192 5557 202 5735
rect 216 5557 226 5735
rect 240 5557 250 5735
rect 264 5557 274 5735
rect 288 5557 298 5735
rect 312 5557 322 5735
rect 336 5557 346 5735
rect 360 5557 370 5735
rect 384 5557 394 5735
rect 408 5557 418 5735
rect 432 5557 442 5735
rect 456 5557 466 5735
rect 480 5557 490 5735
rect 504 5557 514 5735
rect 528 5557 538 5735
rect 552 5557 562 5735
rect 576 5557 586 5735
rect 600 5557 610 5735
rect 624 5557 634 5735
rect 648 5557 658 5735
rect 672 5557 682 5735
rect 696 5557 706 5735
rect 720 5557 730 5735
rect 744 5557 754 5735
rect 768 5557 778 5735
rect 792 5557 802 5735
rect 816 5557 826 5735
rect 840 5557 850 5735
rect 864 5557 874 5735
rect 888 5557 898 5735
rect 912 5557 922 5735
rect 936 5557 946 5735
rect 960 5557 970 5735
rect 984 5557 994 5735
rect 1008 5557 1018 5735
rect 1032 5557 1042 5760
rect 0 5520 1066 5530
rect 48 5317 58 5495
rect 72 5317 82 5495
rect 96 5317 106 5495
rect 120 5317 130 5495
rect 144 5317 154 5495
rect 168 5317 178 5495
rect 192 5317 202 5495
rect 216 5317 226 5495
rect 240 5317 250 5495
rect 264 5317 274 5495
rect 288 5317 298 5495
rect 312 5317 322 5495
rect 336 5317 346 5495
rect 360 5317 370 5495
rect 384 5317 394 5495
rect 408 5317 418 5495
rect 432 5317 442 5495
rect 456 5317 466 5495
rect 480 5317 490 5495
rect 504 5317 514 5495
rect 528 5317 538 5495
rect 552 5317 562 5495
rect 576 5317 586 5495
rect 600 5317 610 5495
rect 624 5317 634 5495
rect 648 5317 658 5495
rect 672 5317 682 5495
rect 696 5317 706 5495
rect 720 5317 730 5495
rect 744 5317 754 5495
rect 768 5317 778 5495
rect 792 5317 802 5495
rect 816 5317 826 5495
rect 840 5317 850 5495
rect 864 5317 874 5495
rect 888 5317 898 5495
rect 912 5317 922 5495
rect 936 5317 946 5495
rect 960 5317 970 5495
rect 984 5317 994 5495
rect 1008 5317 1018 5495
rect 1032 5317 1042 5495
rect 1056 5317 1066 5520
rect 0 5280 1090 5290
rect 48 5077 58 5255
rect 72 5077 82 5255
rect 96 5077 106 5255
rect 120 5077 130 5255
rect 144 5077 154 5255
rect 168 5077 178 5255
rect 192 5077 202 5255
rect 216 5077 226 5255
rect 240 5077 250 5255
rect 264 5077 274 5255
rect 288 5077 298 5255
rect 312 5077 322 5255
rect 336 5077 346 5255
rect 360 5077 370 5255
rect 384 5077 394 5255
rect 408 5077 418 5255
rect 432 5077 442 5255
rect 456 5077 466 5255
rect 480 5077 490 5255
rect 504 5077 514 5255
rect 528 5077 538 5255
rect 552 5077 562 5255
rect 576 5077 586 5255
rect 600 5077 610 5255
rect 624 5077 634 5255
rect 648 5077 658 5255
rect 672 5077 682 5255
rect 696 5077 706 5255
rect 720 5077 730 5255
rect 744 5077 754 5255
rect 768 5077 778 5255
rect 792 5077 802 5255
rect 816 5077 826 5255
rect 840 5077 850 5255
rect 864 5077 874 5255
rect 888 5077 898 5255
rect 912 5077 922 5255
rect 936 5077 946 5255
rect 960 5077 970 5255
rect 984 5077 994 5255
rect 1008 5077 1018 5255
rect 1032 5077 1042 5255
rect 1056 5077 1066 5255
rect 1080 5077 1090 5280
rect 0 5040 1114 5050
rect 48 4837 58 5015
rect 72 4837 82 5015
rect 96 4837 106 5015
rect 120 4837 130 5015
rect 144 4837 154 5015
rect 168 4837 178 5015
rect 192 4837 202 5015
rect 216 4837 226 5015
rect 240 4837 250 5015
rect 264 4837 274 5015
rect 288 4837 298 5015
rect 312 4837 322 5015
rect 336 4837 346 5015
rect 360 4837 370 5015
rect 384 4837 394 5015
rect 408 4837 418 5015
rect 432 4837 442 5015
rect 456 4837 466 5015
rect 480 4837 490 5015
rect 504 4837 514 5015
rect 528 4837 538 5015
rect 552 4837 562 5015
rect 576 4837 586 5015
rect 600 4837 610 5015
rect 624 4837 634 5015
rect 648 4837 658 5015
rect 672 4837 682 5015
rect 696 4837 706 5015
rect 720 4837 730 5015
rect 744 4837 754 5015
rect 768 4837 778 5015
rect 792 4837 802 5015
rect 816 4837 826 5015
rect 840 4837 850 5015
rect 864 4837 874 5015
rect 888 4837 898 5015
rect 912 4837 922 5015
rect 936 4837 946 5015
rect 960 4837 970 5015
rect 984 4837 994 5015
rect 1008 4837 1018 5015
rect 1032 4837 1042 5015
rect 1056 4837 1066 5015
rect 1080 4837 1090 5015
rect 1104 4837 1114 5040
rect 0 4800 1138 4810
rect 48 4597 58 4775
rect 72 4597 82 4775
rect 96 4597 106 4775
rect 120 4597 130 4775
rect 144 4597 154 4775
rect 168 4597 178 4775
rect 192 4597 202 4775
rect 216 4597 226 4775
rect 240 4597 250 4775
rect 264 4597 274 4775
rect 288 4597 298 4775
rect 312 4597 322 4775
rect 336 4597 346 4775
rect 360 4597 370 4775
rect 384 4597 394 4775
rect 408 4597 418 4775
rect 432 4597 442 4775
rect 456 4597 466 4775
rect 480 4597 490 4775
rect 504 4597 514 4775
rect 528 4597 538 4775
rect 552 4597 562 4775
rect 576 4597 586 4775
rect 600 4597 610 4775
rect 624 4597 634 4775
rect 648 4597 658 4775
rect 672 4597 682 4775
rect 696 4597 706 4775
rect 720 4597 730 4775
rect 744 4597 754 4775
rect 768 4597 778 4775
rect 792 4597 802 4775
rect 816 4597 826 4775
rect 840 4597 850 4775
rect 864 4597 874 4775
rect 888 4597 898 4775
rect 912 4597 922 4775
rect 936 4597 946 4775
rect 960 4597 970 4775
rect 984 4597 994 4775
rect 1008 4597 1018 4775
rect 1032 4597 1042 4775
rect 1056 4597 1066 4775
rect 1080 4597 1090 4775
rect 1104 4597 1114 4775
rect 1128 4597 1138 4800
rect 0 4560 1162 4570
rect 48 4357 58 4535
rect 72 4357 82 4535
rect 96 4357 106 4535
rect 120 4357 130 4535
rect 144 4357 154 4535
rect 168 4357 178 4535
rect 192 4357 202 4535
rect 216 4357 226 4535
rect 240 4357 250 4535
rect 264 4357 274 4535
rect 288 4357 298 4535
rect 312 4357 322 4535
rect 336 4357 346 4535
rect 360 4357 370 4535
rect 384 4357 394 4535
rect 408 4357 418 4535
rect 432 4357 442 4535
rect 456 4357 466 4535
rect 480 4357 490 4535
rect 504 4357 514 4535
rect 528 4357 538 4535
rect 552 4357 562 4535
rect 576 4357 586 4535
rect 600 4357 610 4535
rect 624 4357 634 4535
rect 648 4357 658 4535
rect 672 4357 682 4535
rect 696 4357 706 4535
rect 720 4357 730 4535
rect 744 4357 754 4535
rect 768 4357 778 4535
rect 792 4357 802 4535
rect 816 4357 826 4535
rect 840 4357 850 4535
rect 864 4357 874 4535
rect 888 4357 898 4535
rect 912 4357 922 4535
rect 936 4357 946 4535
rect 960 4357 970 4535
rect 984 4357 994 4535
rect 1008 4357 1018 4535
rect 1032 4357 1042 4535
rect 1056 4357 1066 4535
rect 1080 4357 1090 4535
rect 1104 4357 1114 4535
rect 1128 4357 1138 4535
rect 1152 4357 1162 4560
rect 0 4320 1186 4330
rect 48 4117 58 4295
rect 72 4117 82 4295
rect 96 4117 106 4295
rect 120 4117 130 4295
rect 144 4117 154 4295
rect 168 4117 178 4295
rect 192 4117 202 4295
rect 216 4117 226 4295
rect 240 4117 250 4295
rect 264 4117 274 4295
rect 288 4117 298 4295
rect 312 4117 322 4295
rect 336 4117 346 4295
rect 360 4117 370 4295
rect 384 4117 394 4295
rect 408 4117 418 4295
rect 432 4117 442 4295
rect 456 4117 466 4295
rect 480 4117 490 4295
rect 504 4117 514 4295
rect 528 4117 538 4295
rect 552 4117 562 4295
rect 576 4117 586 4295
rect 600 4117 610 4295
rect 624 4117 634 4295
rect 648 4117 658 4295
rect 672 4117 682 4295
rect 696 4117 706 4295
rect 720 4117 730 4295
rect 744 4117 754 4295
rect 768 4117 778 4295
rect 792 4117 802 4295
rect 816 4117 826 4295
rect 840 4117 850 4295
rect 864 4117 874 4295
rect 888 4117 898 4295
rect 912 4117 922 4295
rect 936 4117 946 4295
rect 960 4117 970 4295
rect 984 4117 994 4295
rect 1008 4117 1018 4295
rect 1032 4117 1042 4295
rect 1056 4117 1066 4295
rect 1080 4117 1090 4295
rect 1104 4117 1114 4295
rect 1128 4117 1138 4295
rect 1152 4117 1162 4295
rect 1176 4117 1186 4320
rect 32461 4296 32519 4306
rect 32773 4296 32807 4306
rect 32869 4296 32927 4306
rect 32989 4296 33047 4306
rect 33085 4296 33143 4306
rect 27637 4272 27671 4282
rect 27925 4272 27959 4282
rect 28021 4272 28055 4282
rect 28117 4272 28151 4282
rect 32365 4272 32399 4282
rect 32437 4272 32615 4282
rect 32677 4272 32711 4282
rect 32749 4272 33287 4282
rect 27613 4248 27767 4258
rect 27829 4248 27863 4258
rect 27901 4248 28271 4258
rect 32341 4248 33407 4258
rect 27589 4224 28367 4234
rect 28429 4224 28463 4234
rect 32317 4224 33503 4234
rect 33565 4224 33599 4234
rect 35413 4224 35447 4234
rect 27061 4200 27095 4210
rect 27277 4200 27311 4210
rect 27349 4200 27431 4210
rect 27493 4200 27527 4210
rect 27565 4200 28559 4210
rect 28621 4200 28655 4210
rect 28717 4200 28751 4210
rect 28789 4200 28847 4210
rect 30493 4200 30551 4210
rect 32005 4200 32039 4210
rect 32101 4200 32135 4210
rect 32173 4200 32231 4210
rect 32293 4200 33695 4210
rect 35389 4200 35567 4210
rect 26917 4176 26975 4186
rect 27037 4176 27215 4186
rect 27253 4176 28943 4186
rect 30277 4176 30311 4186
rect 30349 4176 30407 4186
rect 30469 4176 30671 4186
rect 30709 4176 30791 4186
rect 31981 4176 33815 4186
rect 35269 4176 35327 4186
rect 35365 4176 35663 4186
rect 24589 4152 24623 4162
rect 26485 4152 26519 4162
rect 26821 4152 26855 4162
rect 26893 4152 29039 4162
rect 30037 4152 30095 4162
rect 30157 4152 30191 4162
rect 30253 4152 30911 4162
rect 31885 4152 31919 4162
rect 31957 4152 33935 4162
rect 33973 4152 34031 4162
rect 34069 4152 34127 4162
rect 34165 4152 34223 4162
rect 35149 4152 35207 4162
rect 35245 4152 35759 4162
rect 24565 4128 24719 4138
rect 26461 4128 26615 4138
rect 26677 4128 26735 4138
rect 26773 4128 29135 4138
rect 30013 4128 31031 4138
rect 31477 4128 31511 4138
rect 31573 4128 31607 4138
rect 31789 4128 31823 4138
rect 31861 4128 34343 4138
rect 34861 4128 34895 4138
rect 34933 4128 34991 4138
rect 35029 4128 35087 4138
rect 35125 4128 35855 4138
rect 24541 4104 24839 4114
rect 24877 4104 24959 4114
rect 25021 4104 25055 4114
rect 26437 4104 29255 4114
rect 29317 4104 29351 4114
rect 29461 4104 31151 4114
rect 31213 4104 31271 4114
rect 31453 4104 31727 4114
rect 31765 4104 34439 4114
rect 34477 4104 34535 4114
rect 34741 4104 34799 4114
rect 34837 4104 35951 4114
rect 35989 4104 36047 4114
rect 0 4080 1210 4090
rect 48 3877 58 4055
rect 72 3877 82 4055
rect 96 3877 106 4055
rect 120 3877 130 4055
rect 144 3877 154 4055
rect 168 3877 178 4055
rect 192 3877 202 4055
rect 216 3877 226 4055
rect 240 3877 250 4055
rect 264 3877 274 4055
rect 288 3877 298 4055
rect 312 3877 322 4055
rect 336 3877 346 4055
rect 360 3877 370 4055
rect 384 3877 394 4055
rect 408 3877 418 4055
rect 432 3877 442 4055
rect 456 3877 466 4055
rect 480 3877 490 4055
rect 504 3877 514 4055
rect 528 3877 538 4055
rect 552 3877 562 4055
rect 576 3877 586 4055
rect 600 3877 610 4055
rect 624 3877 634 4055
rect 648 3877 658 4055
rect 672 3877 682 4055
rect 696 3877 706 4055
rect 720 3877 730 4055
rect 744 3877 754 4055
rect 768 3877 778 4055
rect 792 3877 802 4055
rect 816 3877 826 4055
rect 840 3877 850 4055
rect 864 3877 874 4055
rect 888 3877 898 4055
rect 912 3877 922 4055
rect 936 3877 946 4055
rect 960 3877 970 4055
rect 984 3877 994 4055
rect 1008 3877 1018 4055
rect 1032 3877 1042 4055
rect 1056 3877 1066 4055
rect 1080 3877 1090 4055
rect 1104 3877 1114 4055
rect 1128 3877 1138 4055
rect 1152 3877 1162 4055
rect 1176 3877 1186 4055
rect 1200 3877 1210 4080
rect 24445 4080 24479 4090
rect 24517 4080 25151 4090
rect 25213 4080 25247 4090
rect 25285 4080 25367 4090
rect 25405 4080 25463 4090
rect 25501 4080 25559 4090
rect 25669 4080 26279 4090
rect 26341 4080 26375 4090
rect 26413 4080 31391 4090
rect 31429 4080 34631 4090
rect 34693 4080 34943 4090
rect 34957 4080 36143 4090
rect 24325 4056 24359 4066
rect 24397 4056 25103 4066
rect 25117 4056 26543 4066
rect 26557 4056 36263 4066
rect 36301 4056 36359 4066
rect 24301 4032 33479 4042
rect 33517 4032 36455 4042
rect 24085 4008 24119 4018
rect 24181 4008 24239 4018
rect 24277 4008 36023 4018
rect 36061 4008 36551 4018
rect 23725 3984 23759 3994
rect 23941 3984 23999 3994
rect 24037 3984 26999 3994
rect 27013 3984 27719 3994
rect 27733 3984 32951 3994
rect 32965 3984 34391 3994
rect 34405 3984 36682 3994
rect 23581 3960 23639 3970
rect 23701 3960 23807 3970
rect 23821 3960 23879 3970
rect 23917 3960 24887 3970
rect 24901 3960 24983 3970
rect 24997 3960 25295 3970
rect 25309 3960 26567 3970
rect 26581 3960 27119 3970
rect 27133 3960 31007 3970
rect 31045 3960 34007 3970
rect 34045 3960 36647 3970
rect 36672 3970 36682 3984
rect 36672 3960 36791 3970
rect 23365 3936 23399 3946
rect 23437 3936 23495 3946
rect 23557 3936 24143 3946
rect 24157 3936 35903 3946
rect 35917 3936 36887 3946
rect 36925 3936 37031 3946
rect 37069 3936 37127 3946
rect 37165 3936 37223 3946
rect 23341 3912 32495 3922
rect 32533 3912 37343 3922
rect 37405 3912 37463 3922
rect 37501 3912 37583 3922
rect 23197 3888 23255 3898
rect 23317 3888 35183 3898
rect 35221 3888 37679 3898
rect 37741 3888 37775 3898
rect 23173 3864 37823 3874
rect 0 3840 1234 3850
rect 48 3637 58 3815
rect 72 3637 82 3815
rect 96 3637 106 3815
rect 120 3637 130 3815
rect 144 3637 154 3815
rect 168 3637 178 3815
rect 192 3637 202 3815
rect 216 3637 226 3815
rect 240 3637 250 3815
rect 264 3637 274 3815
rect 288 3637 298 3815
rect 312 3637 322 3815
rect 336 3637 346 3815
rect 360 3637 370 3815
rect 384 3637 394 3815
rect 408 3637 418 3815
rect 432 3637 442 3815
rect 456 3637 466 3815
rect 480 3637 490 3815
rect 504 3637 514 3815
rect 528 3637 538 3815
rect 552 3637 562 3815
rect 576 3637 586 3815
rect 600 3637 610 3815
rect 624 3637 634 3815
rect 648 3637 658 3815
rect 672 3637 682 3815
rect 696 3637 706 3815
rect 720 3637 730 3815
rect 744 3637 754 3815
rect 768 3637 778 3815
rect 792 3637 802 3815
rect 816 3637 826 3815
rect 840 3637 850 3815
rect 864 3637 874 3815
rect 888 3637 898 3815
rect 912 3637 922 3815
rect 936 3637 946 3815
rect 960 3637 970 3815
rect 984 3637 994 3815
rect 1008 3637 1018 3815
rect 1032 3637 1042 3815
rect 1056 3637 1066 3815
rect 1080 3637 1090 3815
rect 1104 3637 1114 3815
rect 1128 3637 1138 3815
rect 1152 3637 1162 3815
rect 1176 3637 1186 3815
rect 1200 3637 1210 3815
rect 1224 3637 1234 3840
rect 23077 3840 23111 3850
rect 23149 3840 37871 3850
rect 37909 3840 37967 3850
rect 22861 3816 22919 3826
rect 22981 3816 23015 3826
rect 23053 3816 29111 3826
rect 29149 3816 38087 3826
rect 38125 3816 38183 3826
rect 22837 3792 38303 3802
rect 22477 3768 22559 3778
rect 22597 3768 22655 3778
rect 22717 3768 22775 3778
rect 22813 3768 38423 3778
rect 22381 3744 22415 3754
rect 22453 3744 33335 3754
rect 33349 3744 38351 3754
rect 38365 3744 38519 3754
rect 22285 3720 22319 3730
rect 22357 3720 27287 3730
rect 27325 3720 30719 3730
rect 30733 3720 36311 3730
rect 36325 3720 36935 3730
rect 36949 3720 38663 3730
rect 22261 3696 35303 3706
rect 35341 3696 38759 3706
rect 38917 3696 38951 3706
rect 39709 3696 39767 3706
rect 39805 3696 39863 3706
rect 39901 3696 39959 3706
rect 40501 3696 40559 3706
rect 40597 3696 40655 3706
rect 15109 3672 15143 3682
rect 15421 3672 15479 3682
rect 21661 3672 21695 3682
rect 21757 3672 21815 3682
rect 21877 3672 21935 3682
rect 21973 3672 22055 3682
rect 22093 3672 22151 3682
rect 22237 3672 30383 3682
rect 30421 3672 32375 3682
rect 32413 3672 38855 3682
rect 38893 3672 39047 3682
rect 39229 3672 39263 3682
rect 39301 3672 39359 3682
rect 39517 3672 39551 3682
rect 39613 3672 39647 3682
rect 39685 3672 40055 3682
rect 40405 3672 40439 3682
rect 40477 3672 40775 3682
rect 40813 3672 40871 3682
rect 41053 3672 41087 3682
rect 15085 3648 15335 3658
rect 15397 3648 15671 3658
rect 21637 3648 31703 3658
rect 31741 3648 37199 3658
rect 37237 3648 39167 3658
rect 39205 3648 39455 3658
rect 39493 3648 40151 3658
rect 40189 3648 40247 3658
rect 40285 3648 40343 3658
rect 40381 3648 40991 3658
rect 41029 3648 41183 3658
rect 41245 3648 41303 3658
rect 41341 3648 41399 3658
rect 14701 3624 14735 3634
rect 14773 3624 14831 3634
rect 14893 3624 14927 3634
rect 14989 3624 15023 3634
rect 15061 3624 15887 3634
rect 21133 3624 21167 3634
rect 21613 3624 32543 3634
rect 32557 3624 37439 3634
rect 37477 3624 41495 3634
rect 41869 3624 41903 3634
rect 0 3600 1258 3610
rect 48 3397 58 3575
rect 72 3397 82 3575
rect 96 3397 106 3575
rect 120 3397 130 3575
rect 144 3397 154 3575
rect 168 3397 178 3575
rect 192 3397 202 3575
rect 216 3397 226 3575
rect 240 3397 250 3575
rect 264 3397 274 3575
rect 288 3397 298 3575
rect 312 3397 322 3575
rect 336 3397 346 3575
rect 360 3397 370 3575
rect 384 3397 394 3575
rect 408 3397 418 3575
rect 432 3397 442 3575
rect 456 3397 466 3575
rect 480 3397 490 3575
rect 504 3397 514 3575
rect 528 3397 538 3575
rect 552 3397 562 3575
rect 576 3397 586 3575
rect 600 3397 610 3575
rect 624 3397 634 3575
rect 648 3397 658 3575
rect 672 3397 682 3575
rect 696 3397 706 3575
rect 720 3397 730 3575
rect 744 3397 754 3575
rect 768 3397 778 3575
rect 792 3397 802 3575
rect 816 3397 826 3575
rect 840 3397 850 3575
rect 864 3397 874 3575
rect 888 3397 898 3575
rect 912 3397 922 3575
rect 936 3397 946 3575
rect 960 3397 970 3575
rect 984 3397 994 3575
rect 1008 3397 1018 3575
rect 1032 3397 1042 3575
rect 1056 3397 1066 3575
rect 1080 3397 1090 3575
rect 1104 3397 1114 3575
rect 1128 3397 1138 3575
rect 1152 3397 1162 3575
rect 1176 3397 1186 3575
rect 1200 3397 1210 3575
rect 1224 3397 1234 3575
rect 1248 3397 1258 3600
rect 14605 3600 14639 3610
rect 14677 3600 16103 3610
rect 20245 3600 20447 3610
rect 20509 3600 20567 3610
rect 20605 3600 20663 3610
rect 20749 3600 20783 3610
rect 20845 3600 20879 3610
rect 21037 3600 21071 3610
rect 21109 3600 21215 3610
rect 21229 3600 21263 3610
rect 21325 3600 21359 3610
rect 21517 3600 21551 3610
rect 21589 3600 30215 3610
rect 30229 3600 32567 3610
rect 32581 3600 41615 3610
rect 41677 3600 41711 3610
rect 41749 3600 41807 3610
rect 41845 3600 41999 3610
rect 42037 3600 42119 3610
rect 14293 3576 14351 3586
rect 14413 3576 14447 3586
rect 14485 3576 14543 3586
rect 14581 3576 16319 3586
rect 19429 3576 19487 3586
rect 19525 3576 19583 3586
rect 19669 3576 19727 3586
rect 19837 3576 20975 3586
rect 21013 3576 21455 3586
rect 21493 3576 29015 3586
rect 29053 3576 30767 3586
rect 30805 3576 34967 3586
rect 35005 3576 40127 3586
rect 40165 3576 42215 3586
rect 13621 3552 13679 3562
rect 13717 3552 13775 3562
rect 13909 3552 13991 3562
rect 14053 3552 14207 3562
rect 14269 3552 14375 3562
rect 14389 3552 14783 3562
rect 14797 3552 14855 3562
rect 14869 3552 16535 3562
rect 19309 3552 19367 3562
rect 19405 3552 30071 3562
rect 30109 3552 36407 3562
rect 36421 3552 42335 3562
rect 13525 3528 13559 3538
rect 13597 3528 16751 3538
rect 19213 3528 19247 3538
rect 19285 3528 26951 3538
rect 26989 3528 42455 3538
rect 12853 3504 12887 3514
rect 13069 3504 13127 3514
rect 13165 3504 13223 3514
rect 13501 3504 16967 3514
rect 18997 3504 19055 3514
rect 19117 3504 19151 3514
rect 19189 3504 26591 3514
rect 26629 3504 37943 3514
rect 37981 3504 42599 3514
rect 12757 3480 12791 3490
rect 12829 3480 12983 3490
rect 13045 3480 13319 3490
rect 13405 3480 13439 3490
rect 13477 3480 14951 3490
rect 14965 3480 17183 3490
rect 18805 3480 18839 3490
rect 18901 3480 18935 3490
rect 18973 3480 28031 3490
rect 28069 3480 42047 3490
rect 42061 3480 42695 3490
rect 12661 3456 12695 3466
rect 12733 3456 17399 3466
rect 18685 3456 18743 3466
rect 18781 3456 25175 3466
rect 25189 3456 26303 3466
rect 26317 3456 27455 3466
rect 27469 3456 30839 3466
rect 30853 3456 32063 3466
rect 32077 3456 33311 3466
rect 33325 3456 33743 3466
rect 33757 3456 33839 3466
rect 33853 3456 34247 3466
rect 34261 3456 38639 3466
rect 38677 3456 41567 3466
rect 41581 3456 42815 3466
rect 12637 3432 17471 3442
rect 18589 3432 18623 3442
rect 18661 3432 24599 3442
rect 24637 3432 41687 3442
rect 41725 3432 42935 3442
rect 12397 3408 12455 3418
rect 12613 3408 17615 3418
rect 18493 3408 18527 3418
rect 18565 3408 29855 3418
rect 29869 3408 37799 3418
rect 37837 3408 41927 3418
rect 41941 3408 43055 3418
rect 43429 3408 43463 3418
rect 12301 3384 12335 3394
rect 12373 3384 12551 3394
rect 12589 3384 17831 3394
rect 18469 3384 26831 3394
rect 26869 3384 28199 3394
rect 28213 3384 43151 3394
rect 43213 3384 43271 3394
rect 43333 3384 43367 3394
rect 43405 3384 43559 3394
rect 43621 3384 43655 3394
rect 0 3360 1282 3370
rect 48 3157 58 3335
rect 72 3157 82 3335
rect 96 3157 106 3335
rect 120 3157 130 3335
rect 144 3157 154 3335
rect 168 3157 178 3335
rect 192 3157 202 3335
rect 216 3157 226 3335
rect 240 3157 250 3335
rect 264 3157 274 3335
rect 288 3157 298 3335
rect 312 3157 322 3335
rect 336 3157 346 3335
rect 360 3157 370 3335
rect 384 3157 394 3335
rect 408 3157 418 3335
rect 432 3157 442 3335
rect 456 3157 466 3335
rect 480 3157 490 3335
rect 504 3157 514 3335
rect 528 3157 538 3335
rect 552 3157 562 3335
rect 576 3157 586 3335
rect 600 3157 610 3335
rect 624 3157 634 3335
rect 648 3157 658 3335
rect 672 3157 682 3335
rect 696 3157 706 3335
rect 720 3157 730 3335
rect 744 3157 754 3335
rect 768 3157 778 3335
rect 792 3157 802 3335
rect 816 3157 826 3335
rect 840 3157 850 3335
rect 864 3157 874 3335
rect 888 3157 898 3335
rect 912 3157 922 3335
rect 936 3157 946 3335
rect 960 3157 970 3335
rect 984 3157 994 3335
rect 1008 3157 1018 3335
rect 1032 3157 1042 3335
rect 1056 3157 1066 3335
rect 1080 3157 1090 3335
rect 1104 3157 1114 3335
rect 1128 3157 1138 3335
rect 1152 3157 1162 3335
rect 1176 3157 1186 3335
rect 1200 3157 1210 3335
rect 1224 3157 1234 3335
rect 1248 3157 1258 3335
rect 1272 3157 1282 3360
rect 12205 3360 12239 3370
rect 12277 3360 17903 3370
rect 18373 3360 18407 3370
rect 18445 3360 28823 3370
rect 28861 3360 30119 3370
rect 30133 3360 33671 3370
rect 33709 3360 43751 3370
rect 12181 3336 18047 3346
rect 18349 3336 24815 3346
rect 24853 3336 37007 3346
rect 37045 3336 40007 3346
rect 40021 3336 40079 3346
rect 40093 3336 43079 3346
rect 43093 3336 43871 3346
rect 44029 3336 44063 3346
rect 12157 3312 18263 3322
rect 18325 3312 35831 3322
rect 35869 3312 43943 3322
rect 44005 3312 44183 3322
rect 12037 3288 12095 3298
rect 12133 3288 28535 3298
rect 28573 3288 41783 3298
rect 41821 3288 44351 3298
rect 44413 3288 44471 3298
rect 12013 3264 22535 3274
rect 22573 3264 26063 3274
rect 26077 3264 37079 3274
rect 37093 3264 37175 3274
rect 37189 3264 39407 3274
rect 39421 3264 40199 3274
rect 40213 3264 44567 3274
rect 11893 3240 11951 3250
rect 11989 3240 18815 3250
rect 18853 3240 20927 3250
rect 20941 3240 25439 3250
rect 25477 3240 31583 3250
rect 31621 3240 37631 3250
rect 37645 3240 43127 3250
rect 43165 3240 44711 3250
rect 11725 3216 11807 3226
rect 11845 3216 32639 3226
rect 32653 3216 44807 3226
rect 11629 3192 11663 3202
rect 11701 3192 25223 3202
rect 25261 3192 25511 3202
rect 25525 3192 26231 3202
rect 26245 3192 31367 3202
rect 31405 3192 33263 3202
rect 33301 3192 44903 3202
rect 11605 3168 20639 3178
rect 20677 3168 22895 3178
rect 22933 3168 31799 3178
rect 31837 3168 36959 3178
rect 36973 3168 39911 3178
rect 39925 3168 44999 3178
rect 11485 3144 11519 3154
rect 11581 3144 38711 3154
rect 38725 3144 41351 3154
rect 41365 3144 45119 3154
rect 0 3120 1306 3130
rect 48 2917 58 3095
rect 72 2917 82 3095
rect 96 2917 106 3095
rect 120 2917 130 3095
rect 144 2917 154 3095
rect 168 2917 178 3095
rect 192 2917 202 3095
rect 216 2917 226 3095
rect 240 2917 250 3095
rect 264 2917 274 3095
rect 288 2917 298 3095
rect 312 2917 322 3095
rect 336 2917 346 3095
rect 360 2917 370 3095
rect 384 2917 394 3095
rect 408 2917 418 3095
rect 432 2917 442 3095
rect 456 2917 466 3095
rect 480 2917 490 3095
rect 504 2917 514 3095
rect 528 2917 538 3095
rect 552 2917 562 3095
rect 576 2917 586 3095
rect 600 2917 610 3095
rect 624 2917 634 3095
rect 648 2917 658 3095
rect 672 2917 682 3095
rect 696 2917 706 3095
rect 720 2917 730 3095
rect 744 2917 754 3095
rect 768 2917 778 3095
rect 792 2917 802 3095
rect 816 2917 826 3095
rect 840 2917 850 3095
rect 864 2917 874 3095
rect 888 2917 898 3095
rect 912 2917 922 3095
rect 936 2917 946 3095
rect 960 2917 970 3095
rect 984 2917 994 3095
rect 1008 2917 1018 3095
rect 1032 2917 1042 3095
rect 1056 2917 1066 3095
rect 1080 2917 1090 3095
rect 1104 2917 1114 3095
rect 1128 2917 1138 3095
rect 1152 2917 1162 3095
rect 1176 2917 1186 3095
rect 1200 2917 1210 3095
rect 1224 2917 1234 3095
rect 1248 2917 1258 3095
rect 1272 2917 1282 3095
rect 1296 2917 1306 3120
rect 11389 3120 11423 3130
rect 11461 3120 13247 3130
rect 13261 3120 14903 3130
rect 14941 3120 21767 3130
rect 21781 3120 23951 3130
rect 23965 3120 24791 3130
rect 24805 3120 31295 3130
rect 31309 3120 38015 3130
rect 38029 3120 45215 3130
rect 11365 3096 19079 3106
rect 19093 3096 23615 3106
rect 23653 3096 26207 3106
rect 26221 3096 27791 3106
rect 27805 3096 28175 3106
rect 28189 3096 28295 3106
rect 28309 3096 28391 3106
rect 28405 3096 33911 3106
rect 33949 3096 37847 3106
rect 37885 3096 45335 3106
rect 11341 3072 20759 3082
rect 20797 3072 45455 3082
rect 11245 3048 11279 3058
rect 11317 3048 24215 3058
rect 24253 3048 26783 3058
rect 26797 3048 27983 3058
rect 27997 3048 28079 3058
rect 28093 3048 34319 3058
rect 34357 3048 37103 3058
rect 37141 3048 43343 3058
rect 43381 3048 45551 3058
rect 11149 3024 11183 3034
rect 11221 3024 18599 3034
rect 18637 3024 22391 3034
rect 22429 3024 45647 3034
rect 11101 3000 19031 3010
rect 19069 3000 26351 3010
rect 26389 3000 30287 3010
rect 30325 3000 45767 3010
rect 45829 3000 45863 3010
rect 45901 3000 45959 3010
rect 10981 2976 11039 2986
rect 11077 2976 23855 2986
rect 23893 2976 28487 2986
rect 28501 2976 28583 2986
rect 28597 2976 28679 2986
rect 28693 2976 28967 2986
rect 28981 2976 29279 2986
rect 29293 2976 33383 2986
rect 33421 2976 46055 2986
rect 46093 2976 46151 2986
rect 10885 2952 10919 2962
rect 10957 2952 20399 2962
rect 20413 2952 38279 2962
rect 38317 2952 46247 2962
rect 8629 2928 8663 2938
rect 8701 2928 8735 2938
rect 10861 2928 18719 2938
rect 18757 2928 31895 2938
rect 31933 2928 46367 2938
rect 8605 2904 8759 2914
rect 8797 2904 8855 2914
rect 10837 2904 46463 2914
rect 46501 2904 46559 2914
rect 46885 2904 46943 2914
rect 0 2880 1330 2890
rect 48 2677 58 2855
rect 72 2677 82 2855
rect 96 2677 106 2855
rect 120 2677 130 2855
rect 144 2677 154 2855
rect 168 2677 178 2855
rect 192 2677 202 2855
rect 216 2677 226 2855
rect 240 2677 250 2855
rect 264 2677 274 2855
rect 288 2677 298 2855
rect 312 2677 322 2855
rect 336 2677 346 2855
rect 360 2677 370 2855
rect 384 2677 394 2855
rect 408 2677 418 2855
rect 432 2677 442 2855
rect 456 2677 466 2855
rect 480 2677 490 2855
rect 504 2677 514 2855
rect 528 2677 538 2855
rect 552 2677 562 2855
rect 576 2677 586 2855
rect 600 2677 610 2855
rect 624 2677 634 2855
rect 648 2677 658 2855
rect 672 2677 682 2855
rect 696 2677 706 2855
rect 720 2677 730 2855
rect 744 2677 754 2855
rect 768 2677 778 2855
rect 792 2677 802 2855
rect 816 2677 826 2855
rect 840 2677 850 2855
rect 864 2677 874 2855
rect 888 2677 898 2855
rect 912 2677 922 2855
rect 936 2677 946 2855
rect 960 2677 970 2855
rect 984 2677 994 2855
rect 1008 2677 1018 2855
rect 1032 2677 1042 2855
rect 1056 2677 1066 2855
rect 1080 2677 1090 2855
rect 1104 2677 1114 2855
rect 1128 2677 1138 2855
rect 1152 2677 1162 2855
rect 1176 2677 1186 2855
rect 1200 2677 1210 2855
rect 1224 2677 1234 2855
rect 1248 2677 1258 2855
rect 1272 2677 1282 2855
rect 1296 2677 1306 2855
rect 1320 2677 1330 2880
rect 8365 2880 8423 2890
rect 8581 2880 8951 2890
rect 10741 2880 10775 2890
rect 10813 2880 46679 2890
rect 46717 2880 46823 2890
rect 46861 2880 47063 2890
rect 47101 2880 47159 2890
rect 8269 2856 8303 2866
rect 8341 2856 8519 2866
rect 8557 2856 9023 2866
rect 10717 2856 19343 2866
rect 19381 2856 47255 2866
rect 47557 2856 47591 2866
rect 8173 2832 8207 2842
rect 8245 2832 9047 2842
rect 10357 2832 10415 2842
rect 10693 2832 46799 2842
rect 46837 2832 47375 2842
rect 47533 2832 47711 2842
rect 47749 2832 47831 2842
rect 47965 2832 47999 2842
rect 8053 2808 8087 2818
rect 8125 2808 9143 2818
rect 10141 2808 10175 2818
rect 10213 2808 10271 2818
rect 10333 2808 10511 2818
rect 10549 2808 10607 2818
rect 10669 2808 45743 2818
rect 45781 2808 47471 2818
rect 47509 2808 48119 2818
rect 8029 2784 8135 2794
rect 8149 2784 9215 2794
rect 10045 2784 10079 2794
rect 10117 2784 12767 2794
rect 12805 2784 13175 2794
rect 13189 2784 21047 2794
rect 21085 2784 38495 2794
rect 38533 2784 44927 2794
rect 44941 2784 47207 2794
rect 47221 2784 47879 2794
rect 47893 2784 48263 2794
rect 7933 2760 7967 2770
rect 8005 2760 9239 2770
rect 9997 2760 36767 2770
rect 36805 2760 38399 2770
rect 38437 2760 45935 2770
rect 45973 2760 48383 2770
rect 48421 2760 48479 2770
rect 7909 2736 9335 2746
rect 9901 2736 9935 2746
rect 9973 2736 14615 2746
rect 14653 2736 21671 2746
rect 21709 2736 48575 2746
rect 7621 2712 7823 2722
rect 7861 2712 9431 2722
rect 9781 2712 9815 2722
rect 9853 2712 33527 2722
rect 33541 2712 34175 2722
rect 34189 2712 34487 2722
rect 34501 2712 34559 2722
rect 34573 2712 36239 2722
rect 36277 2712 36839 2722
rect 36853 2712 40823 2722
rect 40837 2712 48671 2722
rect 48733 2712 48767 2722
rect 7213 2688 9551 2698
rect 9757 2688 12911 2698
rect 12925 2688 14423 2698
rect 14461 2688 37247 2698
rect 37261 2688 43631 2698
rect 43669 2688 48863 2698
rect 6997 2664 9647 2674
rect 9709 2664 19463 2674
rect 19501 2664 26711 2674
rect 26749 2664 32687 2674
rect 32725 2664 37655 2674
rect 37693 2664 39839 2674
rect 39877 2664 44039 2674
rect 44077 2664 48959 2674
rect 0 2640 1354 2650
rect 48 2437 58 2615
rect 72 2437 82 2615
rect 96 2437 106 2615
rect 120 2437 130 2615
rect 144 2437 154 2615
rect 168 2437 178 2615
rect 192 2437 202 2615
rect 216 2437 226 2615
rect 240 2437 250 2615
rect 264 2437 274 2615
rect 288 2437 298 2615
rect 312 2437 322 2615
rect 336 2437 346 2615
rect 360 2437 370 2615
rect 384 2437 394 2615
rect 408 2437 418 2615
rect 432 2437 442 2615
rect 456 2437 466 2615
rect 480 2437 490 2615
rect 504 2437 514 2615
rect 528 2437 538 2615
rect 552 2437 562 2615
rect 576 2437 586 2615
rect 600 2437 610 2615
rect 624 2437 634 2615
rect 648 2437 658 2615
rect 672 2437 682 2615
rect 696 2437 706 2615
rect 720 2437 730 2615
rect 744 2437 754 2615
rect 768 2437 778 2615
rect 792 2437 802 2615
rect 816 2437 826 2615
rect 840 2437 850 2615
rect 864 2437 874 2615
rect 888 2437 898 2615
rect 912 2437 922 2615
rect 936 2437 946 2615
rect 960 2437 970 2615
rect 984 2437 994 2615
rect 1008 2437 1018 2615
rect 1032 2437 1042 2615
rect 1056 2437 1066 2615
rect 1080 2437 1090 2615
rect 1104 2437 1114 2615
rect 1128 2437 1138 2615
rect 1152 2437 1162 2615
rect 1176 2437 1186 2615
rect 1200 2437 1210 2615
rect 1224 2437 1234 2615
rect 1248 2437 1258 2615
rect 1272 2437 1282 2615
rect 1296 2437 1306 2615
rect 1320 2437 1330 2615
rect 1344 2437 1354 2640
rect 5773 2640 5831 2650
rect 5869 2640 5951 2650
rect 5989 2640 6071 2650
rect 6133 2640 6167 2650
rect 6325 2640 6383 2650
rect 6949 2640 44759 2650
rect 44773 2640 45023 2650
rect 45037 2640 49055 2650
rect 49093 2640 49151 2650
rect 5749 2616 6263 2626
rect 6301 2616 6479 2626
rect 6589 2616 10751 2626
rect 10789 2616 11543 2626
rect 11557 2616 40511 2626
rect 40525 2616 49247 2626
rect 5653 2592 5687 2602
rect 5725 2592 13367 2602
rect 13381 2592 19703 2602
rect 19741 2592 24455 2602
rect 24493 2592 28895 2602
rect 28909 2592 29087 2602
rect 29101 2592 34103 2602
rect 34141 2592 36071 2602
rect 36085 2592 38831 2602
rect 38869 2592 49343 2602
rect 5557 2568 5591 2578
rect 5629 2568 9527 2578
rect 9565 2568 11255 2578
rect 11293 2568 39335 2578
rect 39373 2568 45623 2578
rect 45661 2568 49439 2578
rect 5533 2544 12431 2554
rect 12469 2544 28127 2554
rect 28165 2544 28319 2554
rect 28333 2544 49535 2554
rect 5413 2520 5447 2530
rect 5485 2520 7871 2530
rect 7885 2520 22991 2530
rect 23029 2520 37991 2530
rect 38005 2520 46991 2530
rect 47005 2520 47279 2530
rect 47293 2520 49631 2530
rect 5317 2496 5351 2506
rect 5389 2496 9623 2506
rect 9661 2496 37703 2506
rect 37717 2496 41639 2506
rect 41653 2496 43295 2506
rect 43309 2496 49727 2506
rect 5293 2472 9119 2482
rect 9157 2472 14711 2482
rect 14749 2472 48095 2482
rect 48133 2472 49391 2482
rect 49405 2472 49847 2482
rect 50029 2472 50063 2482
rect 5197 2448 5231 2458
rect 5269 2448 6455 2458
rect 6493 2448 12311 2458
rect 12349 2448 26015 2458
rect 26029 2448 35615 2458
rect 35629 2448 37607 2458
rect 37621 2448 38255 2458
rect 38269 2448 47111 2458
rect 47125 2448 49967 2458
rect 50005 2448 50159 2458
rect 5173 2424 8831 2434
rect 8869 2424 8879 2434
rect 8893 2424 9071 2434
rect 9085 2424 9263 2434
rect 9277 2424 13535 2434
rect 13573 2424 25415 2434
rect 25429 2424 30743 2434
rect 30757 2424 34079 2434
rect 34093 2424 39095 2434
rect 39109 2424 40895 2434
rect 40909 2424 44975 2434
rect 45013 2424 46751 2434
rect 46765 2424 48599 2434
rect 48613 2424 49559 2434
rect 49573 2424 49655 2434
rect 49669 2424 50255 2434
rect 0 2400 1378 2410
rect 48 2197 58 2375
rect 72 2197 82 2375
rect 96 2197 106 2375
rect 120 2197 130 2375
rect 144 2197 154 2375
rect 168 2197 178 2375
rect 192 2197 202 2375
rect 216 2197 226 2375
rect 240 2197 250 2375
rect 264 2197 274 2375
rect 288 2197 298 2375
rect 312 2197 322 2375
rect 336 2197 346 2375
rect 360 2197 370 2375
rect 384 2197 394 2375
rect 408 2197 418 2375
rect 432 2197 442 2375
rect 456 2197 466 2375
rect 480 2197 490 2375
rect 504 2197 514 2375
rect 528 2197 538 2375
rect 552 2197 562 2375
rect 576 2197 586 2375
rect 600 2197 610 2375
rect 624 2197 634 2375
rect 648 2197 658 2375
rect 672 2197 682 2375
rect 696 2197 706 2375
rect 720 2197 730 2375
rect 744 2197 754 2375
rect 768 2197 778 2375
rect 792 2197 802 2375
rect 816 2197 826 2375
rect 840 2197 850 2375
rect 864 2197 874 2375
rect 888 2197 898 2375
rect 912 2197 922 2375
rect 936 2197 946 2375
rect 960 2197 970 2375
rect 984 2197 994 2375
rect 1008 2197 1018 2375
rect 1032 2197 1042 2375
rect 1056 2197 1066 2375
rect 1080 2197 1090 2375
rect 1104 2197 1114 2375
rect 1128 2197 1138 2375
rect 1152 2197 1162 2375
rect 1176 2197 1186 2375
rect 1200 2197 1210 2375
rect 1224 2197 1234 2375
rect 1248 2197 1258 2375
rect 1272 2197 1282 2375
rect 1296 2197 1306 2375
rect 1320 2197 1330 2375
rect 1344 2197 1354 2375
rect 1368 2197 1378 2400
rect 5077 2400 5111 2410
rect 5149 2400 7799 2410
rect 7837 2400 35999 2410
rect 36013 2400 39311 2410
rect 39325 2400 43223 2410
rect 43237 2400 46199 2410
rect 46213 2400 47615 2410
rect 47629 2400 48191 2410
rect 48205 2400 48311 2410
rect 48325 2400 48527 2410
rect 48541 2400 50351 2410
rect 5053 2376 8927 2386
rect 8965 2376 13655 2386
rect 13693 2376 46127 2386
rect 46165 2376 46175 2386
rect 46189 2376 50831 2386
rect 4933 2352 4991 2362
rect 5029 2352 6143 2362
rect 6181 2352 6215 2362
rect 6229 2352 6431 2362
rect 6445 2352 7775 2362
rect 7789 2352 32207 2362
rect 32245 2352 34775 2362
rect 34813 2352 43727 2362
rect 43765 2352 50879 2362
rect 51037 2352 51071 2362
rect 4909 2328 27071 2338
rect 27109 2328 29207 2338
rect 29221 2328 32999 2338
rect 33013 2328 51167 2338
rect 51229 2328 51263 2338
rect 4789 2304 4847 2314
rect 4885 2304 36431 2314
rect 36469 2304 39935 2314
rect 39973 2304 44327 2314
rect 44365 2304 50135 2314
rect 50173 2304 51383 2314
rect 4765 2280 5495 2290
rect 5509 2280 15119 2290
rect 15157 2280 44615 2290
rect 44629 2280 44951 2290
rect 44965 2280 45047 2290
rect 45061 2280 47399 2290
rect 47413 2280 51503 2290
rect 4621 2256 10439 2266
rect 10477 2256 15455 2266
rect 15493 2256 21383 2266
rect 21397 2256 24935 2266
rect 24973 2256 43799 2266
rect 43813 2256 46967 2266
rect 46981 2256 51599 2266
rect 51685 2256 51719 2266
rect 4573 2232 43487 2242
rect 43525 2232 50855 2242
rect 50893 2232 51359 2242
rect 51397 2232 51863 2242
rect 4213 2208 8279 2218
rect 8317 2208 12047 2218
rect 12061 2208 21983 2218
rect 21997 2208 36335 2218
rect 36373 2208 36383 2218
rect 36397 2208 36719 2218
rect 36733 2208 36815 2218
rect 36829 2208 38231 2218
rect 38245 2208 38687 2218
rect 38701 2208 42671 2218
rect 42709 2208 49679 2218
rect 49693 2208 51983 2218
rect 3997 2184 21719 2194
rect 21733 2184 28799 2194
rect 28813 2184 30599 2194
rect 30613 2184 39983 2194
rect 39997 2184 40703 2194
rect 40717 2184 41255 2194
rect 41269 2184 47663 2194
rect 47677 2184 52103 2194
rect 0 2160 1402 2170
rect 48 1957 58 2135
rect 72 1957 82 2135
rect 96 1957 106 2135
rect 120 1957 130 2135
rect 144 1957 154 2135
rect 168 1957 178 2135
rect 192 1957 202 2135
rect 216 1957 226 2135
rect 240 1957 250 2135
rect 264 1957 274 2135
rect 288 1957 298 2135
rect 312 1957 322 2135
rect 336 1957 346 2135
rect 360 1957 370 2135
rect 384 1957 394 2135
rect 408 1957 418 2135
rect 432 1957 442 2135
rect 456 1957 466 2135
rect 480 1957 490 2135
rect 504 1957 514 2135
rect 528 1957 538 2135
rect 552 1957 562 2135
rect 576 1957 586 2135
rect 600 1957 610 2135
rect 624 1957 634 2135
rect 648 1957 658 2135
rect 672 1957 682 2135
rect 696 1957 706 2135
rect 720 1957 730 2135
rect 744 1957 754 2135
rect 768 1957 778 2135
rect 792 1957 802 2135
rect 816 1957 826 2135
rect 840 1957 850 2135
rect 864 1957 874 2135
rect 888 1957 898 2135
rect 912 1957 922 2135
rect 936 1957 946 2135
rect 960 1957 970 2135
rect 984 1957 994 2135
rect 1008 1957 1018 2135
rect 1032 1957 1042 2135
rect 1056 1957 1066 2135
rect 1080 1957 1090 2135
rect 1104 1957 1114 2135
rect 1128 1957 1138 2135
rect 1152 1957 1162 2135
rect 1176 1957 1186 2135
rect 1200 1957 1210 2135
rect 1224 1957 1234 2135
rect 1248 1957 1258 2135
rect 1272 1957 1282 2135
rect 1296 1957 1306 2135
rect 1320 1957 1330 2135
rect 1344 1957 1354 2135
rect 1368 1957 1378 2135
rect 1392 1957 1402 2160
rect 3949 2160 22727 2170
rect 22741 2160 52199 2170
rect 3445 2136 3479 2146
rect 3589 2136 8639 2146
rect 8677 2136 47687 2146
rect 47725 2136 49367 2146
rect 49381 2136 52319 2146
rect 3421 2112 9311 2122
rect 9349 2112 13751 2122
rect 13789 2112 18503 2122
rect 18541 2112 28727 2122
rect 28765 2112 42431 2122
rect 42469 2112 51191 2122
rect 51205 2112 51407 2122
rect 51421 2112 52439 2122
rect 3229 2088 3263 2098
rect 3301 2088 3359 2098
rect 3397 2088 6239 2098
rect 6277 2088 27743 2098
rect 27781 2088 34871 2098
rect 34909 2088 44231 2098
rect 44245 2088 44423 2098
rect 44437 2088 52559 2098
rect 3133 2064 3167 2074
rect 3205 2064 8495 2074
rect 8533 2064 10895 2074
rect 10933 2064 45839 2074
rect 45877 2064 52487 2074
rect 52501 2064 52679 2074
rect 3109 2040 8399 2050
rect 8437 2040 45311 2050
rect 45349 2040 52799 2050
rect 3085 2016 22199 2026
rect 22213 2016 38159 2026
rect 38197 2016 40535 2026
rect 40573 2016 48455 2026
rect 48493 2016 49175 2026
rect 49189 2016 50183 2026
rect 50197 2016 52895 2026
rect 2989 1992 3023 2002
rect 3061 1992 11855 2002
rect 11869 1992 48167 2002
rect 48181 1992 49751 2002
rect 49765 1992 53015 2002
rect 2965 1968 6359 1978
rect 6397 1968 25127 1978
rect 25165 1968 51839 1978
rect 51877 1968 53135 1978
rect 2941 1944 30575 1954
rect 30589 1944 33623 1954
rect 33637 1944 35927 1954
rect 35965 1944 40319 1954
rect 40357 1944 46919 1954
rect 46957 1944 50087 1954
rect 50101 1944 53231 1954
rect 0 1920 1426 1930
rect 48 1717 58 1895
rect 72 1717 82 1895
rect 96 1717 106 1895
rect 120 1717 130 1895
rect 144 1717 154 1895
rect 168 1717 178 1895
rect 192 1717 202 1895
rect 216 1717 226 1895
rect 240 1717 250 1895
rect 264 1717 274 1895
rect 288 1717 298 1895
rect 312 1717 322 1895
rect 336 1717 346 1895
rect 360 1717 370 1895
rect 384 1717 394 1895
rect 408 1717 418 1895
rect 432 1717 442 1895
rect 456 1717 466 1895
rect 480 1717 490 1895
rect 504 1717 514 1895
rect 528 1717 538 1895
rect 552 1717 562 1895
rect 576 1717 586 1895
rect 600 1717 610 1895
rect 624 1717 634 1895
rect 648 1717 658 1895
rect 672 1717 682 1895
rect 696 1717 706 1895
rect 720 1717 730 1895
rect 744 1717 754 1895
rect 768 1717 778 1895
rect 792 1717 802 1895
rect 816 1717 826 1895
rect 840 1717 850 1895
rect 864 1717 874 1895
rect 888 1717 898 1895
rect 912 1717 922 1895
rect 936 1717 946 1895
rect 960 1717 970 1895
rect 984 1717 994 1895
rect 1008 1717 1018 1895
rect 1032 1717 1042 1895
rect 1056 1717 1066 1895
rect 1080 1717 1090 1895
rect 1104 1717 1114 1895
rect 1128 1717 1138 1895
rect 1152 1717 1162 1895
rect 1176 1717 1186 1895
rect 1200 1717 1210 1895
rect 1224 1717 1234 1895
rect 1248 1717 1258 1895
rect 1272 1717 1282 1895
rect 1296 1717 1306 1895
rect 1320 1717 1330 1895
rect 1344 1717 1354 1895
rect 1368 1717 1378 1895
rect 1392 1717 1402 1895
rect 1416 1717 1426 1920
rect 2845 1920 2879 1930
rect 2917 1920 21239 1930
rect 21277 1920 25343 1930
rect 25381 1920 28871 1930
rect 28885 1920 32831 1930
rect 32845 1920 42887 1930
rect 42901 1920 44087 1930
rect 44101 1920 52607 1930
rect 52621 1920 52727 1930
rect 52741 1920 53375 1930
rect 2821 1896 5927 1906
rect 5965 1896 11159 1906
rect 11197 1896 28343 1906
rect 28381 1896 53471 1906
rect 2797 1872 11735 1882
rect 11749 1872 22031 1882
rect 22069 1872 30167 1882
rect 30205 1872 36743 1882
rect 36757 1872 38999 1882
rect 39013 1872 42983 1882
rect 42997 1872 44735 1882
rect 44749 1872 45719 1882
rect 45733 1872 45791 1882
rect 45805 1872 45911 1882
rect 45925 1872 52871 1882
rect 52909 1872 53543 1882
rect 2677 1848 2735 1858
rect 2773 1848 24647 1858
rect 24661 1848 27839 1858
rect 27877 1848 39815 1858
rect 39829 1848 42503 1858
rect 42517 1848 48623 1858
rect 48637 1848 51287 1858
rect 51301 1848 51431 1858
rect 51445 1848 52007 1858
rect 52021 1848 53591 1858
rect 2581 1824 2615 1834
rect 2653 1824 3335 1834
rect 3373 1824 6047 1834
rect 6085 1824 8447 1834
rect 8461 1824 12527 1834
rect 12565 1824 14519 1834
rect 14557 1824 21527 1834
rect 21565 1824 33791 1834
rect 33829 1824 43535 1834
rect 43573 1824 48551 1834
rect 48589 1824 53111 1834
rect 53149 1824 53639 1834
rect 2557 1800 3239 1810
rect 3277 1800 9455 1810
rect 9493 1800 12479 1810
rect 12493 1800 14327 1810
rect 14365 1800 53663 1810
rect 2413 1776 9287 1786
rect 9301 1776 17663 1786
rect 17677 1776 53615 1786
rect 53653 1776 53687 1786
rect 2365 1752 53783 1762
rect 2005 1728 3455 1738
rect 3493 1728 9407 1738
rect 9469 1728 15431 1738
rect 15445 1728 22511 1738
rect 22525 1728 43583 1738
rect 43597 1728 53903 1738
rect 1789 1704 9095 1714
rect 9109 1704 13823 1714
rect 13837 1704 53999 1714
rect 0 1680 1450 1690
rect 1440 1666 1450 1680
rect 1741 1680 53639 1690
rect 53677 1680 54071 1690
rect 1440 1656 9503 1666
rect 9517 1656 12503 1666
rect 12517 1656 46607 1666
rect 46621 1656 50207 1666
rect 50221 1656 54119 1666
rect 48 1477 58 1655
rect 72 1477 82 1655
rect 96 1477 106 1655
rect 120 1477 130 1655
rect 144 1477 154 1655
rect 168 1477 178 1655
rect 192 1477 202 1655
rect 216 1477 226 1655
rect 240 1477 250 1655
rect 264 1477 274 1655
rect 288 1477 298 1655
rect 312 1477 322 1655
rect 336 1477 346 1655
rect 360 1477 370 1655
rect 384 1477 394 1655
rect 408 1477 418 1655
rect 432 1477 442 1655
rect 456 1477 466 1655
rect 480 1477 490 1655
rect 504 1477 514 1655
rect 528 1477 538 1655
rect 552 1477 562 1655
rect 576 1477 586 1655
rect 600 1477 610 1655
rect 624 1477 634 1655
rect 648 1477 658 1655
rect 672 1477 682 1655
rect 696 1477 706 1655
rect 720 1477 730 1655
rect 744 1477 754 1655
rect 768 1477 778 1655
rect 792 1477 802 1655
rect 816 1477 826 1655
rect 840 1477 850 1655
rect 864 1477 874 1655
rect 888 1477 898 1655
rect 912 1477 922 1655
rect 936 1477 946 1655
rect 960 1477 970 1655
rect 984 1477 994 1655
rect 1008 1477 1018 1655
rect 1032 1477 1042 1655
rect 1056 1477 1066 1655
rect 1080 1477 1090 1655
rect 1104 1477 1114 1655
rect 1128 1477 1138 1655
rect 1152 1477 1162 1655
rect 1176 1477 1186 1655
rect 1200 1477 1210 1655
rect 1224 1477 1234 1655
rect 1248 1477 1258 1655
rect 1272 1474 1282 1655
rect 1296 1498 1306 1655
rect 1320 1522 1330 1655
rect 1344 1546 1354 1655
rect 1368 1594 1378 1655
rect 1392 1618 1402 1655
rect 1416 1642 1426 1655
rect 1416 1632 46895 1642
rect 46909 1632 49199 1642
rect 49213 1632 54215 1642
rect 1392 1608 9383 1618
rect 9445 1608 35639 1618
rect 35677 1608 41279 1618
rect 41317 1608 42263 1618
rect 42277 1608 45095 1618
rect 45133 1608 48983 1618
rect 48997 1608 49775 1618
rect 49789 1608 51527 1618
rect 51541 1608 54095 1618
rect 54133 1608 54167 1618
rect 54181 1608 54311 1618
rect 1368 1584 9191 1594
rect 9229 1584 13199 1594
rect 13237 1584 33575 1594
rect 33613 1584 51143 1594
rect 51181 1584 54370 1594
rect 54360 1573 54370 1584
rect 1381 1560 5327 1570
rect 5365 1560 9215 1570
rect 9253 1560 41375 1570
rect 41413 1560 41543 1570
rect 41557 1560 42863 1570
rect 42877 1560 42959 1570
rect 42973 1560 44495 1570
rect 44509 1560 48359 1570
rect 48397 1560 54335 1570
rect 1344 1536 8999 1546
rect 9037 1536 44159 1546
rect 44197 1536 51695 1546
rect 51733 1536 54407 1546
rect 1320 1512 8711 1522
rect 8749 1512 8975 1522
rect 8989 1512 9167 1522
rect 9181 1512 9359 1522
rect 9373 1512 12863 1522
rect 12901 1512 27503 1522
rect 27541 1512 32591 1522
rect 32629 1512 39743 1522
rect 39781 1512 43919 1522
rect 43933 1512 53351 1522
rect 53389 1512 54551 1522
rect 1296 1488 33455 1498
rect 33469 1488 35495 1498
rect 35509 1488 44135 1498
rect 44149 1488 54671 1498
rect 1272 1464 54791 1474
rect 0 1440 3311 1450
rect 3325 1440 40295 1450
rect 40309 1440 52055 1450
rect 52069 1440 54887 1450
rect 1261 1416 5423 1426
rect 5461 1416 9719 1426
rect 9733 1416 21335 1426
rect 21373 1416 28511 1426
rect 28525 1416 42527 1426
rect 42541 1416 45479 1426
rect 45493 1416 46415 1426
rect 46429 1416 53207 1426
rect 53245 1416 54287 1426
rect 54373 1416 54983 1426
rect 48 1237 58 1415
rect 72 1237 82 1415
rect 96 1237 106 1415
rect 120 1237 130 1415
rect 144 1237 154 1415
rect 168 1237 178 1415
rect 192 1237 202 1415
rect 216 1237 226 1415
rect 240 1237 250 1415
rect 264 1237 274 1415
rect 288 1237 298 1415
rect 312 1237 322 1415
rect 336 1237 346 1415
rect 360 1237 370 1415
rect 384 1237 394 1415
rect 408 1237 418 1415
rect 432 1237 442 1415
rect 456 1237 466 1415
rect 480 1237 490 1415
rect 504 1237 514 1415
rect 528 1237 538 1415
rect 552 1237 562 1415
rect 576 1237 586 1415
rect 600 1237 610 1415
rect 624 1237 634 1415
rect 648 1237 658 1415
rect 672 1237 682 1415
rect 696 1237 706 1415
rect 720 1237 730 1415
rect 744 1237 754 1415
rect 768 1237 778 1415
rect 792 1237 802 1415
rect 816 1237 826 1415
rect 840 1237 850 1415
rect 864 1237 874 1415
rect 888 1237 898 1415
rect 912 1237 922 1415
rect 936 1237 946 1415
rect 960 1237 970 1415
rect 984 1237 994 1415
rect 1008 1237 1018 1415
rect 1032 1237 1042 1415
rect 1056 1234 1066 1415
rect 1080 1258 1090 1415
rect 1104 1282 1114 1415
rect 1128 1306 1138 1415
rect 1152 1330 1162 1415
rect 1176 1354 1186 1415
rect 1200 1378 1210 1415
rect 1224 1402 1234 1415
rect 1224 1392 19127 1402
rect 19165 1392 28439 1402
rect 28477 1392 37367 1402
rect 37381 1392 41879 1402
rect 41917 1392 55079 1402
rect 1200 1368 5567 1378
rect 5605 1368 11111 1378
rect 11125 1368 23735 1378
rect 23773 1368 31631 1378
rect 31645 1368 35039 1378
rect 35053 1368 38039 1378
rect 38053 1368 46775 1378
rect 46789 1368 53759 1378
rect 53797 1368 54263 1378
rect 54349 1368 55175 1378
rect 1176 1344 23375 1354
rect 23413 1344 45527 1354
rect 45565 1344 47975 1354
rect 48013 1344 53711 1354
rect 53725 1344 55295 1354
rect 1152 1320 4823 1330
rect 4861 1320 10247 1330
rect 10285 1320 12215 1330
rect 12253 1320 32111 1330
rect 32149 1320 40415 1330
rect 40453 1320 47351 1330
rect 47389 1320 49271 1330
rect 49285 1320 54767 1330
rect 54805 1320 55415 1330
rect 1128 1296 12959 1306
rect 12997 1296 20855 1306
rect 20893 1296 23207 1306
rect 23221 1296 23591 1306
rect 23605 1296 23663 1306
rect 23677 1296 41951 1306
rect 41965 1296 44855 1306
rect 44869 1296 51815 1306
rect 51829 1296 53303 1306
rect 53317 1296 53855 1306
rect 53869 1296 54695 1306
rect 54709 1296 55535 1306
rect 1104 1272 9791 1282
rect 9829 1272 33023 1282
rect 33061 1272 38927 1282
rect 38965 1272 41423 1282
rect 41437 1272 46031 1282
rect 46069 1272 47135 1282
rect 47173 1272 47183 1282
rect 47197 1272 51479 1282
rect 51517 1272 52175 1282
rect 52213 1272 54047 1282
rect 54085 1272 54143 1282
rect 54157 1272 55631 1282
rect 1080 1248 5663 1258
rect 5701 1248 24095 1258
rect 24133 1248 27383 1258
rect 27397 1248 43823 1258
rect 43837 1248 55151 1258
rect 55189 1248 55751 1258
rect 1056 1224 11495 1234
rect 11533 1224 27407 1234
rect 27445 1224 29159 1234
rect 29173 1224 38447 1234
rect 38461 1224 40967 1234
rect 41005 1224 46439 1234
rect 46477 1224 49607 1234
rect 49645 1224 53831 1234
rect 53845 1224 55679 1234
rect 55693 1224 55847 1234
rect 0 1200 20471 1210
rect 20485 1200 31175 1210
rect 31189 1200 35807 1210
rect 35821 1200 37511 1210
rect 37525 1200 38807 1210
rect 38821 1200 40103 1210
rect 40117 1200 45503 1210
rect 45517 1200 47903 1210
rect 47917 1200 49295 1210
rect 49309 1200 54839 1210
rect 54853 1200 55954 1210
rect 1045 1176 9911 1186
rect 9949 1176 14999 1186
rect 15037 1176 23231 1186
rect 23269 1176 31247 1186
rect 31285 1176 31655 1186
rect 31669 1176 37319 1186
rect 37357 1176 37559 1186
rect 37597 1176 42095 1186
rect 42133 1176 47807 1186
rect 47845 1176 49871 1186
rect 49885 1176 55055 1186
rect 55093 1176 55919 1186
rect 55944 1186 55954 1200
rect 56053 1200 56471 1210
rect 55944 1176 56639 1186
rect 48 997 58 1175
rect 72 997 82 1175
rect 96 997 106 1175
rect 120 997 130 1175
rect 144 997 154 1175
rect 168 997 178 1175
rect 192 997 202 1175
rect 216 997 226 1175
rect 240 997 250 1175
rect 264 997 274 1175
rect 288 997 298 1175
rect 312 997 322 1175
rect 336 997 346 1175
rect 360 997 370 1175
rect 384 997 394 1175
rect 408 997 418 1175
rect 432 997 442 1175
rect 456 997 466 1175
rect 480 997 490 1175
rect 504 997 514 1175
rect 528 997 538 1175
rect 552 997 562 1175
rect 576 997 586 1175
rect 600 997 610 1175
rect 624 997 634 1175
rect 648 997 658 1175
rect 672 997 682 1175
rect 696 997 706 1175
rect 720 997 730 1175
rect 744 997 754 1175
rect 768 997 778 1175
rect 792 997 802 1175
rect 816 997 826 1175
rect 840 994 850 1175
rect 864 1018 874 1175
rect 888 1042 898 1175
rect 912 1066 922 1175
rect 936 1090 946 1175
rect 960 1114 970 1175
rect 984 1138 994 1175
rect 1008 1162 1018 1175
rect 1008 1152 10055 1162
rect 10093 1152 19631 1162
rect 19645 1152 41591 1162
rect 41629 1152 42143 1162
rect 42157 1152 44879 1162
rect 44917 1152 48647 1162
rect 48685 1152 52703 1162
rect 52717 1152 56687 1162
rect 984 1128 43031 1138
rect 43069 1128 49943 1138
rect 49981 1128 50303 1138
rect 50317 1128 51767 1138
rect 51781 1128 54071 1138
rect 54085 1128 56783 1138
rect 960 1104 5879 1114
rect 5893 1104 23471 1114
rect 23509 1104 29231 1114
rect 29269 1104 39623 1114
rect 39661 1104 42743 1114
rect 42757 1104 47447 1114
rect 47485 1104 53159 1114
rect 53173 1104 55727 1114
rect 55765 1104 56879 1114
rect 936 1080 7943 1090
rect 7981 1080 30887 1090
rect 30925 1080 38063 1090
rect 38101 1080 40631 1090
rect 40669 1080 44447 1090
rect 44485 1080 46583 1090
rect 46597 1080 52415 1090
rect 52453 1080 56975 1090
rect 912 1056 2855 1066
rect 2893 1056 4799 1066
rect 4813 1056 8471 1066
rect 8485 1056 10991 1066
rect 11005 1056 11759 1066
rect 11773 1056 21431 1066
rect 21469 1056 25031 1066
rect 25069 1056 27167 1066
rect 27181 1056 30863 1066
rect 30877 1056 41759 1066
rect 41773 1056 51911 1066
rect 51925 1056 57095 1066
rect 888 1032 8063 1042
rect 8101 1032 21143 1042
rect 21181 1032 29063 1042
rect 29077 1032 44111 1042
rect 44125 1032 45695 1042
rect 45709 1032 46271 1042
rect 46285 1032 51095 1042
rect 51109 1032 53399 1042
rect 53413 1032 54527 1042
rect 54565 1032 57167 1042
rect 864 1008 8183 1018
rect 8221 1008 44543 1018
rect 44581 1008 48695 1018
rect 48709 1008 51119 1018
rect 51133 1008 53519 1018
rect 53557 1008 55511 1018
rect 55549 1008 57191 1018
rect 840 984 5807 994
rect 5845 984 10583 994
rect 10621 984 12671 994
rect 12709 984 38735 994
rect 38773 984 49223 994
rect 49261 984 53927 994
rect 53941 984 57287 994
rect 0 960 20519 970
rect 20533 960 28991 970
rect 29005 960 34271 970
rect 34285 960 37271 970
rect 37285 960 49583 970
rect 49597 960 54719 970
rect 54733 960 55031 970
rect 55045 960 55799 970
rect 55813 960 55895 970
rect 55909 960 57359 970
rect 829 936 11639 946
rect 11677 936 20183 946
rect 20197 936 38591 946
rect 38605 936 44303 946
rect 44317 936 46727 946
rect 46741 936 48911 946
rect 48925 936 52631 946
rect 52645 936 55439 946
rect 55453 936 57119 946
rect 57133 936 57383 946
rect 48 757 58 935
rect 72 757 82 935
rect 96 757 106 935
rect 120 757 130 935
rect 144 757 154 935
rect 168 757 178 935
rect 192 757 202 935
rect 216 757 226 935
rect 240 757 250 935
rect 264 757 274 935
rect 288 757 298 935
rect 312 757 322 935
rect 336 757 346 935
rect 360 757 370 935
rect 384 757 394 935
rect 408 757 418 935
rect 432 757 442 935
rect 456 757 466 935
rect 480 757 490 935
rect 504 757 514 935
rect 528 757 538 935
rect 552 757 562 935
rect 576 757 586 935
rect 600 757 610 935
rect 624 757 634 935
rect 648 754 658 935
rect 672 778 682 935
rect 696 802 706 935
rect 720 826 730 935
rect 744 874 754 935
rect 768 898 778 935
rect 792 922 802 935
rect 792 912 10151 922
rect 10189 912 42911 922
rect 42949 912 50039 922
rect 50077 912 56903 922
rect 56917 912 57479 922
rect 768 888 13415 898
rect 13453 888 36863 898
rect 36901 888 46391 898
rect 46405 888 52535 898
rect 52573 888 56711 898
rect 56725 888 57599 898
rect 744 864 1151 874
rect 1165 864 8903 874
rect 8917 864 17879 874
rect 17917 864 18383 874
rect 18421 864 33983 874
rect 33997 864 40679 874
rect 40693 864 42623 874
rect 42637 864 46223 874
rect 46261 864 50327 874
rect 50365 864 54479 874
rect 54493 864 54575 874
rect 54589 864 57647 874
rect 57661 864 57695 874
rect 757 840 5087 850
rect 5125 840 9023 850
rect 9061 840 10487 850
rect 10525 840 30647 850
rect 30685 840 35543 850
rect 35581 840 50231 850
rect 50269 840 55391 850
rect 55429 840 57815 850
rect 720 816 13295 826
rect 13333 816 19223 826
rect 19261 816 28919 826
rect 28957 816 32783 826
rect 32821 816 37751 826
rect 37789 816 41975 826
rect 42013 816 49511 826
rect 49549 816 55607 826
rect 55645 816 57887 826
rect 696 792 12071 802
rect 12109 792 22751 802
rect 22789 792 27935 802
rect 27973 792 34415 802
rect 34453 792 35063 802
rect 35101 792 40031 802
rect 40069 792 47039 802
rect 47077 792 50111 802
rect 50125 792 53663 802
rect 53701 792 57071 802
rect 57109 792 57791 802
rect 57829 792 57911 802
rect 672 768 4967 778
rect 5005 768 10391 778
rect 10429 768 13103 778
rect 13141 768 21191 778
rect 21205 768 24407 778
rect 24421 768 31055 778
rect 31069 768 34367 778
rect 34381 768 38975 778
rect 38989 768 39383 778
rect 39397 768 45191 778
rect 45229 768 46655 778
rect 46693 768 49703 778
rect 49741 768 51791 778
rect 51805 768 57215 778
rect 57229 768 57335 778
rect 57373 768 57935 778
rect 648 744 11399 754
rect 11437 744 29327 754
rect 29365 744 33767 754
rect 33781 744 42191 754
rect 42229 744 49319 754
rect 49357 744 57263 754
rect 57301 744 57671 754
rect 57709 744 58031 754
rect 0 720 23831 730
rect 23845 720 24191 730
rect 24205 720 45407 730
rect 45421 720 55703 730
rect 55717 720 57047 730
rect 57061 720 57407 730
rect 57421 720 57959 730
rect 57973 720 58127 730
rect 637 696 2999 706
rect 3037 696 4943 706
rect 4957 696 27191 706
rect 27229 696 27695 706
rect 27709 696 34511 706
rect 34549 696 35471 706
rect 35485 696 39431 706
rect 39469 696 50447 706
rect 50461 696 56447 706
rect 56485 696 58234 706
rect 48 517 58 695
rect 72 517 82 695
rect 96 517 106 695
rect 120 517 130 695
rect 144 517 154 695
rect 168 517 178 695
rect 192 517 202 695
rect 216 517 226 695
rect 240 517 250 695
rect 264 517 274 695
rect 288 517 298 695
rect 312 517 322 695
rect 336 517 346 695
rect 360 517 370 695
rect 384 517 394 695
rect 408 517 418 695
rect 432 517 442 695
rect 456 514 466 695
rect 480 538 490 695
rect 504 562 514 695
rect 528 610 538 695
rect 552 634 562 695
rect 576 658 586 695
rect 600 682 610 695
rect 600 672 3143 682
rect 3181 672 11903 682
rect 11917 672 50279 682
rect 50293 672 54383 682
rect 54421 672 55559 682
rect 55573 672 57455 682
rect 57493 672 58199 682
rect 58224 682 58234 696
rect 58224 672 58319 682
rect 576 648 11783 658
rect 11821 648 28631 658
rect 28669 648 30815 658
rect 30829 648 30935 658
rect 30949 648 31079 658
rect 31093 648 31319 658
rect 31333 648 31535 658
rect 31549 648 36119 658
rect 36157 648 37919 658
rect 37933 648 38327 658
rect 38341 648 38783 658
rect 38797 648 42791 658
rect 42829 648 46007 658
rect 46021 648 46103 658
rect 46117 648 46295 658
rect 46309 648 51575 658
rect 51613 648 51959 658
rect 51997 648 53063 658
rect 53077 648 58391 658
rect 552 624 11927 634
rect 11965 624 19559 634
rect 19597 624 22295 634
rect 22333 624 22871 634
rect 22885 624 42311 634
rect 42349 624 52823 634
rect 52837 624 53567 634
rect 53605 624 54815 634
rect 54829 624 54911 634
rect 54925 624 55463 634
rect 55477 624 55871 634
rect 55885 624 58439 634
rect 528 600 9575 610
rect 9589 600 11015 610
rect 11053 600 20375 610
rect 20389 600 26255 610
rect 26293 600 31487 610
rect 31525 600 52655 610
rect 52693 600 54863 610
rect 54901 600 58079 610
rect 58093 600 58247 610
rect 58261 600 58559 610
rect 541 576 5999 586
rect 6013 576 8807 586
rect 8821 576 18095 586
rect 18109 576 56615 586
rect 56653 576 57431 586
rect 57445 576 58055 586
rect 58069 576 58607 586
rect 58621 576 58655 586
rect 504 552 20423 562
rect 20461 552 36215 562
rect 36229 552 39575 562
rect 39589 552 43895 562
rect 43909 552 48791 562
rect 48805 552 49007 562
rect 49021 552 49103 562
rect 49117 552 51311 562
rect 51325 552 51887 562
rect 51901 552 52031 562
rect 52045 552 54455 562
rect 54469 552 55223 562
rect 55237 552 57311 562
rect 57349 552 57623 562
rect 57637 552 58343 562
rect 58357 552 58703 562
rect 480 528 41159 538
rect 41197 528 45263 538
rect 45277 528 49031 538
rect 49069 528 54599 538
rect 54613 528 55247 538
rect 55261 528 55319 538
rect 55333 528 57143 538
rect 57181 528 57575 538
rect 57613 528 58727 538
rect 456 504 2591 514
rect 2629 504 2687 514
rect 2701 504 5783 514
rect 5797 504 9863 514
rect 9877 504 10007 514
rect 10021 504 37823 514
rect 37837 504 41111 514
rect 41125 504 43247 514
rect 43285 504 45575 514
rect 45589 504 49823 514
rect 49861 504 56759 514
rect 56797 504 57527 514
rect 57541 504 57863 514
rect 57925 504 58775 514
rect 0 480 14495 490
rect 14509 480 33239 490
rect 33253 480 36983 490
rect 36997 480 40919 490
rect 40933 480 47423 490
rect 47437 480 47759 490
rect 47773 480 53327 490
rect 53341 480 58175 490
rect 58189 480 58463 490
rect 58477 480 58583 490
rect 58597 480 58823 490
rect 445 456 2711 466
rect 2749 456 14807 466
rect 14845 456 27647 466
rect 27685 456 44255 466
rect 44269 456 52367 466
rect 52381 456 56855 466
rect 56893 456 58415 466
rect 58453 456 58871 466
rect 48 277 58 455
rect 72 277 82 455
rect 96 277 106 455
rect 120 277 130 455
rect 144 277 154 455
rect 168 277 178 455
rect 192 277 202 455
rect 216 277 226 455
rect 240 274 250 455
rect 264 298 274 455
rect 288 322 298 455
rect 312 346 322 455
rect 336 370 346 455
rect 360 394 370 455
rect 384 418 394 455
rect 408 442 418 455
rect 408 432 15647 442
rect 15685 432 45983 442
rect 45997 432 48887 442
rect 48901 432 54647 442
rect 54685 432 58943 442
rect 384 408 15863 418
rect 15901 408 23783 418
rect 23797 408 32879 418
rect 32893 408 35711 418
rect 35725 408 40607 418
rect 40621 408 47303 418
rect 47317 408 51743 418
rect 51757 408 55775 418
rect 55789 408 57239 418
rect 57253 408 58991 418
rect 360 384 16079 394
rect 16117 384 23087 394
rect 23125 384 46511 394
rect 46525 384 47639 394
rect 47653 384 48287 394
rect 48301 384 48503 394
rect 48517 384 52247 394
rect 52261 384 57167 394
rect 57205 384 59063 394
rect 336 360 16295 370
rect 16333 360 20903 370
rect 20917 360 46343 370
rect 46381 360 48839 370
rect 48877 360 49415 370
rect 49453 360 57359 370
rect 57397 360 58679 370
rect 58741 360 58967 370
rect 59005 360 59111 370
rect 312 336 16511 346
rect 16549 336 21911 346
rect 21949 336 44831 346
rect 44845 336 45383 346
rect 45397 336 52991 346
rect 53029 336 55271 346
rect 55309 336 58631 346
rect 58669 336 59159 346
rect 288 312 14183 322
rect 14221 312 15167 322
rect 15181 312 15503 322
rect 15517 312 15719 322
rect 15733 312 15935 322
rect 15949 312 16151 322
rect 16165 312 16367 322
rect 16381 312 16583 322
rect 16597 312 16799 322
rect 16813 312 17015 322
rect 17029 312 17231 322
rect 17245 312 17447 322
rect 17485 312 32903 322
rect 32941 312 35591 322
rect 35605 312 35687 322
rect 35701 312 35783 322
rect 35797 312 35879 322
rect 35893 312 36599 322
rect 36613 312 39143 322
rect 39181 312 43439 322
rect 43477 312 51239 322
rect 51277 312 59087 322
rect 59125 312 59207 322
rect 264 288 16727 298
rect 16765 288 20951 298
rect 20989 288 24335 298
rect 24373 288 49127 298
rect 49165 288 53975 298
rect 54013 288 54239 298
rect 54325 288 56591 298
rect 56605 288 57743 298
rect 57757 288 58271 298
rect 58285 288 58919 298
rect 58957 288 59039 298
rect 59077 288 59303 298
rect 240 264 16943 274
rect 16981 264 22631 274
rect 22669 264 26495 274
rect 26533 264 42575 274
rect 42613 264 43679 274
rect 43693 264 43847 274
rect 43885 264 47567 274
rect 47605 264 58295 274
rect 58333 264 59351 274
rect 0 240 30959 250
rect 30973 240 31223 250
rect 31237 240 31679 250
rect 31693 240 33191 250
rect 33205 240 33863 250
rect 33877 240 34751 250
rect 34765 240 42551 250
rect 42565 240 44639 250
rect 44653 240 51335 250
rect 51349 240 53087 250
rect 53101 240 53279 250
rect 53293 240 54935 250
rect 54949 240 59279 250
rect 59317 240 59423 250
rect 229 216 17159 226
rect 17197 216 21407 226
rect 21421 216 23279 226
rect 23293 216 27143 226
rect 27157 216 34703 226
rect 34717 216 36191 226
rect 36205 216 38567 226
rect 38581 216 41471 226
rect 41509 216 44687 226
rect 44725 216 47327 226
rect 47341 216 49487 226
rect 49501 216 56951 226
rect 56989 216 58751 226
rect 58789 216 59482 226
rect 48 34 58 215
rect 72 58 82 215
rect 96 82 106 215
rect 120 130 130 215
rect 144 154 154 215
rect 168 178 178 215
rect 192 202 202 215
rect 192 192 15311 202
rect 15349 192 18863 202
rect 18877 192 20711 202
rect 20725 192 20807 202
rect 20821 192 21287 202
rect 21301 192 24695 202
rect 24733 192 33119 202
rect 33157 192 35423 202
rect 35461 192 48743 202
rect 48781 192 48815 202
rect 48829 192 50999 202
rect 51013 192 52127 202
rect 52141 192 53879 202
rect 53917 192 56807 202
rect 56821 192 58847 202
rect 58885 192 59447 202
rect 59472 202 59482 216
rect 59472 192 59543 202
rect 168 168 17375 178
rect 17413 168 33431 178
rect 33445 168 36527 178
rect 36565 168 41063 178
rect 41101 168 44783 178
rect 44821 168 48047 178
rect 48061 168 52775 178
rect 52813 168 54959 178
rect 54997 168 55103 178
rect 55117 168 58103 178
rect 58141 168 58151 178
rect 58165 168 58487 178
rect 58501 168 59591 178
rect 144 144 17591 154
rect 17629 144 21791 154
rect 21829 144 22487 154
rect 22501 144 24767 154
rect 24781 144 25079 154
rect 25093 144 26639 154
rect 26653 144 31127 154
rect 31165 144 32015 154
rect 32053 144 39239 154
rect 39277 144 50807 154
rect 50845 144 52295 154
rect 52333 144 54191 154
rect 54229 144 56639 154
rect 56653 144 56735 154
rect 56749 144 56831 154
rect 56845 144 57719 154
rect 57733 144 59639 154
rect 120 120 6191 130
rect 6205 120 17807 130
rect 17845 120 25535 130
rect 25573 120 27359 130
rect 27373 120 29183 130
rect 29197 120 34607 130
rect 34645 120 40847 130
rect 40885 120 46535 130
rect 46573 120 53447 130
rect 53485 120 56663 130
rect 56701 120 57911 130
rect 57949 120 57983 130
rect 57997 120 59519 130
rect 59557 120 59722 130
rect 133 96 5207 106
rect 5245 96 8735 106
rect 8773 96 30527 106
rect 30565 96 40751 106
rect 40789 96 52079 106
rect 52117 96 53543 106
rect 53557 96 57503 106
rect 57517 96 57839 106
rect 57901 96 59687 106
rect 59712 106 59722 120
rect 59712 96 59759 106
rect 96 72 6407 82
rect 6421 72 13967 82
rect 14005 72 14111 82
rect 14125 72 15239 82
rect 15253 72 15575 82
rect 15589 72 15791 82
rect 15805 72 16007 82
rect 16021 72 16223 82
rect 16237 72 16439 82
rect 16453 72 16655 82
rect 16669 72 16871 82
rect 16885 72 17087 82
rect 17101 72 17303 82
rect 17317 72 17519 82
rect 17533 72 17735 82
rect 17749 72 17951 82
rect 17965 72 18167 82
rect 18181 72 22127 82
rect 22165 72 23975 82
rect 24013 72 24047 82
rect 24061 72 34199 82
rect 34237 72 36479 82
rect 36493 72 39023 82
rect 39061 72 39071 82
rect 39085 72 45143 82
rect 45157 72 48935 82
rect 48973 72 49463 82
rect 49477 72 49895 82
rect 49909 72 52943 82
rect 52957 72 55823 82
rect 55861 72 59567 82
rect 59605 72 59842 82
rect 72 48 6095 58
rect 6109 48 18023 58
rect 18061 48 20543 58
rect 20581 48 21839 58
rect 21853 48 22943 58
rect 22957 48 28247 58
rect 28285 48 35735 58
rect 35773 48 40223 58
rect 40261 48 47231 58
rect 47269 48 48239 58
rect 48277 48 48431 58
rect 48445 48 51647 58
rect 51661 48 55007 58
rect 55021 48 55343 58
rect 55357 48 57023 58
rect 57037 48 59327 58
rect 59365 48 59807 58
rect 59832 58 59842 72
rect 59832 48 59879 58
rect 48 24 18250 34
rect 7752 13 7762 24
rect 18240 13 18250 24
rect 18277 24 18922 34
rect 18912 13 18922 24
rect 18949 24 39538 34
rect 33216 13 33226 24
rect 39528 13 39538 24
rect 39565 24 45442 34
rect 42384 13 42394 24
rect 45432 13 45442 24
rect 45469 24 51058 34
rect 51048 13 51058 24
rect 51085 24 58018 34
rect 58008 13 58018 24
rect 58045 24 58378 34
rect 58368 13 58378 24
rect 58405 24 58546 34
rect 58536 13 58546 24
rect 58573 24 58810 34
rect 58800 13 58810 24
rect 58837 24 59410 34
rect 59400 13 59410 24
rect 59437 24 59938 34
rect 59928 13 59938 24
<< m2contact >>
rect 47 15383 61 15397
rect 47 15335 61 15349
rect 47 15143 61 15157
rect 71 15143 85 15157
rect 47 15095 61 15109
rect 71 15095 85 15109
rect 47 14903 61 14917
rect 71 14903 85 14917
rect 95 14903 109 14917
rect 47 14855 61 14869
rect 71 14855 85 14869
rect 95 14855 109 14869
rect 47 14663 61 14677
rect 71 14663 85 14677
rect 95 14663 109 14677
rect 119 14663 133 14677
rect 47 14615 61 14629
rect 71 14615 85 14629
rect 95 14615 109 14629
rect 119 14615 133 14629
rect 47 14423 61 14437
rect 71 14423 85 14437
rect 95 14423 109 14437
rect 119 14423 133 14437
rect 143 14423 157 14437
rect 47 14375 61 14389
rect 71 14375 85 14389
rect 95 14375 109 14389
rect 119 14375 133 14389
rect 143 14375 157 14389
rect 47 14183 61 14197
rect 71 14183 85 14197
rect 95 14183 109 14197
rect 119 14183 133 14197
rect 143 14183 157 14197
rect 167 14183 181 14197
rect 47 14135 61 14149
rect 71 14135 85 14149
rect 95 14135 109 14149
rect 119 14135 133 14149
rect 143 14135 157 14149
rect 167 14135 181 14149
rect 47 13943 61 13957
rect 71 13943 85 13957
rect 95 13943 109 13957
rect 119 13943 133 13957
rect 143 13943 157 13957
rect 167 13943 181 13957
rect 191 13943 205 13957
rect 47 13895 61 13909
rect 71 13895 85 13909
rect 95 13895 109 13909
rect 119 13895 133 13909
rect 143 13895 157 13909
rect 167 13895 181 13909
rect 191 13895 205 13909
rect 47 13703 61 13717
rect 71 13703 85 13717
rect 95 13703 109 13717
rect 119 13703 133 13717
rect 143 13703 157 13717
rect 167 13703 181 13717
rect 191 13703 205 13717
rect 215 13703 229 13717
rect 47 13655 61 13669
rect 71 13655 85 13669
rect 95 13655 109 13669
rect 119 13655 133 13669
rect 143 13655 157 13669
rect 167 13655 181 13669
rect 191 13655 205 13669
rect 215 13655 229 13669
rect 47 13463 61 13477
rect 71 13463 85 13477
rect 95 13463 109 13477
rect 119 13463 133 13477
rect 143 13463 157 13477
rect 167 13463 181 13477
rect 191 13463 205 13477
rect 215 13463 229 13477
rect 239 13463 253 13477
rect 47 13415 61 13429
rect 71 13415 85 13429
rect 95 13415 109 13429
rect 119 13415 133 13429
rect 143 13415 157 13429
rect 167 13415 181 13429
rect 191 13415 205 13429
rect 215 13415 229 13429
rect 239 13415 253 13429
rect 47 13223 61 13237
rect 71 13223 85 13237
rect 95 13223 109 13237
rect 119 13223 133 13237
rect 143 13223 157 13237
rect 167 13223 181 13237
rect 191 13223 205 13237
rect 215 13223 229 13237
rect 239 13223 253 13237
rect 263 13223 277 13237
rect 47 13175 61 13189
rect 71 13175 85 13189
rect 95 13175 109 13189
rect 119 13175 133 13189
rect 143 13175 157 13189
rect 167 13175 181 13189
rect 191 13175 205 13189
rect 215 13175 229 13189
rect 239 13175 253 13189
rect 263 13175 277 13189
rect 47 12983 61 12997
rect 71 12983 85 12997
rect 95 12983 109 12997
rect 119 12983 133 12997
rect 143 12983 157 12997
rect 167 12983 181 12997
rect 191 12983 205 12997
rect 215 12983 229 12997
rect 239 12983 253 12997
rect 263 12983 277 12997
rect 287 12983 301 12997
rect 47 12935 61 12949
rect 71 12935 85 12949
rect 95 12935 109 12949
rect 119 12935 133 12949
rect 143 12935 157 12949
rect 167 12935 181 12949
rect 191 12935 205 12949
rect 215 12935 229 12949
rect 239 12935 253 12949
rect 263 12935 277 12949
rect 287 12935 301 12949
rect 47 12743 61 12757
rect 71 12743 85 12757
rect 95 12743 109 12757
rect 119 12743 133 12757
rect 143 12743 157 12757
rect 167 12743 181 12757
rect 191 12743 205 12757
rect 215 12743 229 12757
rect 239 12743 253 12757
rect 263 12743 277 12757
rect 287 12743 301 12757
rect 311 12743 325 12757
rect 47 12695 61 12709
rect 71 12695 85 12709
rect 95 12695 109 12709
rect 119 12695 133 12709
rect 143 12695 157 12709
rect 167 12695 181 12709
rect 191 12695 205 12709
rect 215 12695 229 12709
rect 239 12695 253 12709
rect 263 12695 277 12709
rect 287 12695 301 12709
rect 311 12695 325 12709
rect 47 12503 61 12517
rect 71 12503 85 12517
rect 95 12503 109 12517
rect 119 12503 133 12517
rect 143 12503 157 12517
rect 167 12503 181 12517
rect 191 12503 205 12517
rect 215 12503 229 12517
rect 239 12503 253 12517
rect 263 12503 277 12517
rect 287 12503 301 12517
rect 311 12503 325 12517
rect 335 12503 349 12517
rect 47 12455 61 12469
rect 71 12455 85 12469
rect 95 12455 109 12469
rect 119 12455 133 12469
rect 143 12455 157 12469
rect 167 12455 181 12469
rect 191 12455 205 12469
rect 215 12455 229 12469
rect 239 12455 253 12469
rect 263 12455 277 12469
rect 287 12455 301 12469
rect 311 12455 325 12469
rect 335 12455 349 12469
rect 47 12263 61 12277
rect 71 12263 85 12277
rect 95 12263 109 12277
rect 119 12263 133 12277
rect 143 12263 157 12277
rect 167 12263 181 12277
rect 191 12263 205 12277
rect 215 12263 229 12277
rect 239 12263 253 12277
rect 263 12263 277 12277
rect 287 12263 301 12277
rect 311 12263 325 12277
rect 335 12263 349 12277
rect 359 12263 373 12277
rect 47 12215 61 12229
rect 71 12215 85 12229
rect 95 12215 109 12229
rect 119 12215 133 12229
rect 143 12215 157 12229
rect 167 12215 181 12229
rect 191 12215 205 12229
rect 215 12215 229 12229
rect 239 12215 253 12229
rect 263 12215 277 12229
rect 287 12215 301 12229
rect 311 12215 325 12229
rect 335 12215 349 12229
rect 359 12215 373 12229
rect 47 12023 61 12037
rect 71 12023 85 12037
rect 95 12023 109 12037
rect 119 12023 133 12037
rect 143 12023 157 12037
rect 167 12023 181 12037
rect 191 12023 205 12037
rect 215 12023 229 12037
rect 239 12023 253 12037
rect 263 12023 277 12037
rect 287 12023 301 12037
rect 311 12023 325 12037
rect 335 12023 349 12037
rect 359 12023 373 12037
rect 383 12023 397 12037
rect 47 11975 61 11989
rect 71 11975 85 11989
rect 95 11975 109 11989
rect 119 11975 133 11989
rect 143 11975 157 11989
rect 167 11975 181 11989
rect 191 11975 205 11989
rect 215 11975 229 11989
rect 239 11975 253 11989
rect 263 11975 277 11989
rect 287 11975 301 11989
rect 311 11975 325 11989
rect 335 11975 349 11989
rect 359 11975 373 11989
rect 383 11975 397 11989
rect 47 11783 61 11797
rect 71 11783 85 11797
rect 95 11783 109 11797
rect 119 11783 133 11797
rect 143 11783 157 11797
rect 167 11783 181 11797
rect 191 11783 205 11797
rect 215 11783 229 11797
rect 239 11783 253 11797
rect 263 11783 277 11797
rect 287 11783 301 11797
rect 311 11783 325 11797
rect 335 11783 349 11797
rect 359 11783 373 11797
rect 383 11783 397 11797
rect 407 11783 421 11797
rect 47 11735 61 11749
rect 71 11735 85 11749
rect 95 11735 109 11749
rect 119 11735 133 11749
rect 143 11735 157 11749
rect 167 11735 181 11749
rect 191 11735 205 11749
rect 215 11735 229 11749
rect 239 11735 253 11749
rect 263 11735 277 11749
rect 287 11735 301 11749
rect 311 11735 325 11749
rect 335 11735 349 11749
rect 359 11735 373 11749
rect 383 11735 397 11749
rect 407 11735 421 11749
rect 47 11543 61 11557
rect 71 11543 85 11557
rect 95 11543 109 11557
rect 119 11543 133 11557
rect 143 11543 157 11557
rect 167 11543 181 11557
rect 191 11543 205 11557
rect 215 11543 229 11557
rect 239 11543 253 11557
rect 263 11543 277 11557
rect 287 11543 301 11557
rect 311 11543 325 11557
rect 335 11543 349 11557
rect 359 11543 373 11557
rect 383 11543 397 11557
rect 407 11543 421 11557
rect 431 11543 445 11557
rect 47 11495 61 11509
rect 71 11495 85 11509
rect 95 11495 109 11509
rect 119 11495 133 11509
rect 143 11495 157 11509
rect 167 11495 181 11509
rect 191 11495 205 11509
rect 215 11495 229 11509
rect 239 11495 253 11509
rect 263 11495 277 11509
rect 287 11495 301 11509
rect 311 11495 325 11509
rect 335 11495 349 11509
rect 359 11495 373 11509
rect 383 11495 397 11509
rect 407 11495 421 11509
rect 431 11495 445 11509
rect 47 11303 61 11317
rect 71 11303 85 11317
rect 95 11303 109 11317
rect 119 11303 133 11317
rect 143 11303 157 11317
rect 167 11303 181 11317
rect 191 11303 205 11317
rect 215 11303 229 11317
rect 239 11303 253 11317
rect 263 11303 277 11317
rect 287 11303 301 11317
rect 311 11303 325 11317
rect 335 11303 349 11317
rect 359 11303 373 11317
rect 383 11303 397 11317
rect 407 11303 421 11317
rect 431 11303 445 11317
rect 455 11303 469 11317
rect 47 11255 61 11269
rect 71 11255 85 11269
rect 95 11255 109 11269
rect 119 11255 133 11269
rect 143 11255 157 11269
rect 167 11255 181 11269
rect 191 11255 205 11269
rect 215 11255 229 11269
rect 239 11255 253 11269
rect 263 11255 277 11269
rect 287 11255 301 11269
rect 311 11255 325 11269
rect 335 11255 349 11269
rect 359 11255 373 11269
rect 383 11255 397 11269
rect 407 11255 421 11269
rect 431 11255 445 11269
rect 455 11255 469 11269
rect 47 11063 61 11077
rect 71 11063 85 11077
rect 95 11063 109 11077
rect 119 11063 133 11077
rect 143 11063 157 11077
rect 167 11063 181 11077
rect 191 11063 205 11077
rect 215 11063 229 11077
rect 239 11063 253 11077
rect 263 11063 277 11077
rect 287 11063 301 11077
rect 311 11063 325 11077
rect 335 11063 349 11077
rect 359 11063 373 11077
rect 383 11063 397 11077
rect 407 11063 421 11077
rect 431 11063 445 11077
rect 455 11063 469 11077
rect 479 11063 493 11077
rect 47 11015 61 11029
rect 71 11015 85 11029
rect 95 11015 109 11029
rect 119 11015 133 11029
rect 143 11015 157 11029
rect 167 11015 181 11029
rect 191 11015 205 11029
rect 215 11015 229 11029
rect 239 11015 253 11029
rect 263 11015 277 11029
rect 287 11015 301 11029
rect 311 11015 325 11029
rect 335 11015 349 11029
rect 359 11015 373 11029
rect 383 11015 397 11029
rect 407 11015 421 11029
rect 431 11015 445 11029
rect 455 11015 469 11029
rect 479 11015 493 11029
rect 47 10823 61 10837
rect 71 10823 85 10837
rect 95 10823 109 10837
rect 119 10823 133 10837
rect 143 10823 157 10837
rect 167 10823 181 10837
rect 191 10823 205 10837
rect 215 10823 229 10837
rect 239 10823 253 10837
rect 263 10823 277 10837
rect 287 10823 301 10837
rect 311 10823 325 10837
rect 335 10823 349 10837
rect 359 10823 373 10837
rect 383 10823 397 10837
rect 407 10823 421 10837
rect 431 10823 445 10837
rect 455 10823 469 10837
rect 479 10823 493 10837
rect 503 10823 517 10837
rect 47 10775 61 10789
rect 71 10775 85 10789
rect 95 10775 109 10789
rect 119 10775 133 10789
rect 143 10775 157 10789
rect 167 10775 181 10789
rect 191 10775 205 10789
rect 215 10775 229 10789
rect 239 10775 253 10789
rect 263 10775 277 10789
rect 287 10775 301 10789
rect 311 10775 325 10789
rect 335 10775 349 10789
rect 359 10775 373 10789
rect 383 10775 397 10789
rect 407 10775 421 10789
rect 431 10775 445 10789
rect 455 10775 469 10789
rect 479 10775 493 10789
rect 503 10775 517 10789
rect 47 10583 61 10597
rect 71 10583 85 10597
rect 95 10583 109 10597
rect 119 10583 133 10597
rect 143 10583 157 10597
rect 167 10583 181 10597
rect 191 10583 205 10597
rect 215 10583 229 10597
rect 239 10583 253 10597
rect 263 10583 277 10597
rect 287 10583 301 10597
rect 311 10583 325 10597
rect 335 10583 349 10597
rect 359 10583 373 10597
rect 383 10583 397 10597
rect 407 10583 421 10597
rect 431 10583 445 10597
rect 455 10583 469 10597
rect 479 10583 493 10597
rect 503 10583 517 10597
rect 527 10583 541 10597
rect 47 10535 61 10549
rect 71 10535 85 10549
rect 95 10535 109 10549
rect 119 10535 133 10549
rect 143 10535 157 10549
rect 167 10535 181 10549
rect 191 10535 205 10549
rect 215 10535 229 10549
rect 239 10535 253 10549
rect 263 10535 277 10549
rect 287 10535 301 10549
rect 311 10535 325 10549
rect 335 10535 349 10549
rect 359 10535 373 10549
rect 383 10535 397 10549
rect 407 10535 421 10549
rect 431 10535 445 10549
rect 455 10535 469 10549
rect 479 10535 493 10549
rect 503 10535 517 10549
rect 527 10535 541 10549
rect 47 10343 61 10357
rect 71 10343 85 10357
rect 95 10343 109 10357
rect 119 10343 133 10357
rect 143 10343 157 10357
rect 167 10343 181 10357
rect 191 10343 205 10357
rect 215 10343 229 10357
rect 239 10343 253 10357
rect 263 10343 277 10357
rect 287 10343 301 10357
rect 311 10343 325 10357
rect 335 10343 349 10357
rect 359 10343 373 10357
rect 383 10343 397 10357
rect 407 10343 421 10357
rect 431 10343 445 10357
rect 455 10343 469 10357
rect 479 10343 493 10357
rect 503 10343 517 10357
rect 527 10343 541 10357
rect 551 10343 565 10357
rect 47 10295 61 10309
rect 71 10295 85 10309
rect 95 10295 109 10309
rect 119 10295 133 10309
rect 143 10295 157 10309
rect 167 10295 181 10309
rect 191 10295 205 10309
rect 215 10295 229 10309
rect 239 10295 253 10309
rect 263 10295 277 10309
rect 287 10295 301 10309
rect 311 10295 325 10309
rect 335 10295 349 10309
rect 359 10295 373 10309
rect 383 10295 397 10309
rect 407 10295 421 10309
rect 431 10295 445 10309
rect 455 10295 469 10309
rect 479 10295 493 10309
rect 503 10295 517 10309
rect 527 10295 541 10309
rect 551 10295 565 10309
rect 47 10103 61 10117
rect 71 10103 85 10117
rect 95 10103 109 10117
rect 119 10103 133 10117
rect 143 10103 157 10117
rect 167 10103 181 10117
rect 191 10103 205 10117
rect 215 10103 229 10117
rect 239 10103 253 10117
rect 263 10103 277 10117
rect 287 10103 301 10117
rect 311 10103 325 10117
rect 335 10103 349 10117
rect 359 10103 373 10117
rect 383 10103 397 10117
rect 407 10103 421 10117
rect 431 10103 445 10117
rect 455 10103 469 10117
rect 479 10103 493 10117
rect 503 10103 517 10117
rect 527 10103 541 10117
rect 551 10103 565 10117
rect 575 10103 589 10117
rect 47 10055 61 10069
rect 71 10055 85 10069
rect 95 10055 109 10069
rect 119 10055 133 10069
rect 143 10055 157 10069
rect 167 10055 181 10069
rect 191 10055 205 10069
rect 215 10055 229 10069
rect 239 10055 253 10069
rect 263 10055 277 10069
rect 287 10055 301 10069
rect 311 10055 325 10069
rect 335 10055 349 10069
rect 359 10055 373 10069
rect 383 10055 397 10069
rect 407 10055 421 10069
rect 431 10055 445 10069
rect 455 10055 469 10069
rect 479 10055 493 10069
rect 503 10055 517 10069
rect 527 10055 541 10069
rect 551 10055 565 10069
rect 575 10055 589 10069
rect 47 9863 61 9877
rect 71 9863 85 9877
rect 95 9863 109 9877
rect 119 9863 133 9877
rect 143 9863 157 9877
rect 167 9863 181 9877
rect 191 9863 205 9877
rect 215 9863 229 9877
rect 239 9863 253 9877
rect 263 9863 277 9877
rect 287 9863 301 9877
rect 311 9863 325 9877
rect 335 9863 349 9877
rect 359 9863 373 9877
rect 383 9863 397 9877
rect 407 9863 421 9877
rect 431 9863 445 9877
rect 455 9863 469 9877
rect 479 9863 493 9877
rect 503 9863 517 9877
rect 527 9863 541 9877
rect 551 9863 565 9877
rect 575 9863 589 9877
rect 599 9863 613 9877
rect 47 9815 61 9829
rect 71 9815 85 9829
rect 95 9815 109 9829
rect 119 9815 133 9829
rect 143 9815 157 9829
rect 167 9815 181 9829
rect 191 9815 205 9829
rect 215 9815 229 9829
rect 239 9815 253 9829
rect 263 9815 277 9829
rect 287 9815 301 9829
rect 311 9815 325 9829
rect 335 9815 349 9829
rect 359 9815 373 9829
rect 383 9815 397 9829
rect 407 9815 421 9829
rect 431 9815 445 9829
rect 455 9815 469 9829
rect 479 9815 493 9829
rect 503 9815 517 9829
rect 527 9815 541 9829
rect 551 9815 565 9829
rect 575 9815 589 9829
rect 599 9815 613 9829
rect 47 9623 61 9637
rect 71 9623 85 9637
rect 95 9623 109 9637
rect 119 9623 133 9637
rect 143 9623 157 9637
rect 167 9623 181 9637
rect 191 9623 205 9637
rect 215 9623 229 9637
rect 239 9623 253 9637
rect 263 9623 277 9637
rect 287 9623 301 9637
rect 311 9623 325 9637
rect 335 9623 349 9637
rect 359 9623 373 9637
rect 383 9623 397 9637
rect 407 9623 421 9637
rect 431 9623 445 9637
rect 455 9623 469 9637
rect 479 9623 493 9637
rect 503 9623 517 9637
rect 527 9623 541 9637
rect 551 9623 565 9637
rect 575 9623 589 9637
rect 599 9623 613 9637
rect 623 9623 637 9637
rect 47 9575 61 9589
rect 71 9575 85 9589
rect 95 9575 109 9589
rect 119 9575 133 9589
rect 143 9575 157 9589
rect 167 9575 181 9589
rect 191 9575 205 9589
rect 215 9575 229 9589
rect 239 9575 253 9589
rect 263 9575 277 9589
rect 287 9575 301 9589
rect 311 9575 325 9589
rect 335 9575 349 9589
rect 359 9575 373 9589
rect 383 9575 397 9589
rect 407 9575 421 9589
rect 431 9575 445 9589
rect 455 9575 469 9589
rect 479 9575 493 9589
rect 503 9575 517 9589
rect 527 9575 541 9589
rect 551 9575 565 9589
rect 575 9575 589 9589
rect 599 9575 613 9589
rect 623 9575 637 9589
rect 47 9383 61 9397
rect 71 9383 85 9397
rect 95 9383 109 9397
rect 119 9383 133 9397
rect 143 9383 157 9397
rect 167 9383 181 9397
rect 191 9383 205 9397
rect 215 9383 229 9397
rect 239 9383 253 9397
rect 263 9383 277 9397
rect 287 9383 301 9397
rect 311 9383 325 9397
rect 335 9383 349 9397
rect 359 9383 373 9397
rect 383 9383 397 9397
rect 407 9383 421 9397
rect 431 9383 445 9397
rect 455 9383 469 9397
rect 479 9383 493 9397
rect 503 9383 517 9397
rect 527 9383 541 9397
rect 551 9383 565 9397
rect 575 9383 589 9397
rect 599 9383 613 9397
rect 623 9383 637 9397
rect 647 9383 661 9397
rect 47 9335 61 9349
rect 71 9335 85 9349
rect 95 9335 109 9349
rect 119 9335 133 9349
rect 143 9335 157 9349
rect 167 9335 181 9349
rect 191 9335 205 9349
rect 215 9335 229 9349
rect 239 9335 253 9349
rect 263 9335 277 9349
rect 287 9335 301 9349
rect 311 9335 325 9349
rect 335 9335 349 9349
rect 359 9335 373 9349
rect 383 9335 397 9349
rect 407 9335 421 9349
rect 431 9335 445 9349
rect 455 9335 469 9349
rect 479 9335 493 9349
rect 503 9335 517 9349
rect 527 9335 541 9349
rect 551 9335 565 9349
rect 575 9335 589 9349
rect 599 9335 613 9349
rect 623 9335 637 9349
rect 647 9335 661 9349
rect 47 9143 61 9157
rect 71 9143 85 9157
rect 95 9143 109 9157
rect 119 9143 133 9157
rect 143 9143 157 9157
rect 167 9143 181 9157
rect 191 9143 205 9157
rect 215 9143 229 9157
rect 239 9143 253 9157
rect 263 9143 277 9157
rect 287 9143 301 9157
rect 311 9143 325 9157
rect 335 9143 349 9157
rect 359 9143 373 9157
rect 383 9143 397 9157
rect 407 9143 421 9157
rect 431 9143 445 9157
rect 455 9143 469 9157
rect 479 9143 493 9157
rect 503 9143 517 9157
rect 527 9143 541 9157
rect 551 9143 565 9157
rect 575 9143 589 9157
rect 599 9143 613 9157
rect 623 9143 637 9157
rect 647 9143 661 9157
rect 671 9143 685 9157
rect 47 9095 61 9109
rect 71 9095 85 9109
rect 95 9095 109 9109
rect 119 9095 133 9109
rect 143 9095 157 9109
rect 167 9095 181 9109
rect 191 9095 205 9109
rect 215 9095 229 9109
rect 239 9095 253 9109
rect 263 9095 277 9109
rect 287 9095 301 9109
rect 311 9095 325 9109
rect 335 9095 349 9109
rect 359 9095 373 9109
rect 383 9095 397 9109
rect 407 9095 421 9109
rect 431 9095 445 9109
rect 455 9095 469 9109
rect 479 9095 493 9109
rect 503 9095 517 9109
rect 527 9095 541 9109
rect 551 9095 565 9109
rect 575 9095 589 9109
rect 599 9095 613 9109
rect 623 9095 637 9109
rect 647 9095 661 9109
rect 671 9095 685 9109
rect 47 8903 61 8917
rect 71 8903 85 8917
rect 95 8903 109 8917
rect 119 8903 133 8917
rect 143 8903 157 8917
rect 167 8903 181 8917
rect 191 8903 205 8917
rect 215 8903 229 8917
rect 239 8903 253 8917
rect 263 8903 277 8917
rect 287 8903 301 8917
rect 311 8903 325 8917
rect 335 8903 349 8917
rect 359 8903 373 8917
rect 383 8903 397 8917
rect 407 8903 421 8917
rect 431 8903 445 8917
rect 455 8903 469 8917
rect 479 8903 493 8917
rect 503 8903 517 8917
rect 527 8903 541 8917
rect 551 8903 565 8917
rect 575 8903 589 8917
rect 599 8903 613 8917
rect 623 8903 637 8917
rect 647 8903 661 8917
rect 671 8903 685 8917
rect 695 8903 709 8917
rect 47 8855 61 8869
rect 71 8855 85 8869
rect 95 8855 109 8869
rect 119 8855 133 8869
rect 143 8855 157 8869
rect 167 8855 181 8869
rect 191 8855 205 8869
rect 215 8855 229 8869
rect 239 8855 253 8869
rect 263 8855 277 8869
rect 287 8855 301 8869
rect 311 8855 325 8869
rect 335 8855 349 8869
rect 359 8855 373 8869
rect 383 8855 397 8869
rect 407 8855 421 8869
rect 431 8855 445 8869
rect 455 8855 469 8869
rect 479 8855 493 8869
rect 503 8855 517 8869
rect 527 8855 541 8869
rect 551 8855 565 8869
rect 575 8855 589 8869
rect 599 8855 613 8869
rect 623 8855 637 8869
rect 647 8855 661 8869
rect 671 8855 685 8869
rect 695 8855 709 8869
rect 47 8663 61 8677
rect 71 8663 85 8677
rect 95 8663 109 8677
rect 119 8663 133 8677
rect 143 8663 157 8677
rect 167 8663 181 8677
rect 191 8663 205 8677
rect 215 8663 229 8677
rect 239 8663 253 8677
rect 263 8663 277 8677
rect 287 8663 301 8677
rect 311 8663 325 8677
rect 335 8663 349 8677
rect 359 8663 373 8677
rect 383 8663 397 8677
rect 407 8663 421 8677
rect 431 8663 445 8677
rect 455 8663 469 8677
rect 479 8663 493 8677
rect 503 8663 517 8677
rect 527 8663 541 8677
rect 551 8663 565 8677
rect 575 8663 589 8677
rect 599 8663 613 8677
rect 623 8663 637 8677
rect 647 8663 661 8677
rect 671 8663 685 8677
rect 695 8663 709 8677
rect 719 8663 733 8677
rect 47 8615 61 8629
rect 71 8615 85 8629
rect 95 8615 109 8629
rect 119 8615 133 8629
rect 143 8615 157 8629
rect 167 8615 181 8629
rect 191 8615 205 8629
rect 215 8615 229 8629
rect 239 8615 253 8629
rect 263 8615 277 8629
rect 287 8615 301 8629
rect 311 8615 325 8629
rect 335 8615 349 8629
rect 359 8615 373 8629
rect 383 8615 397 8629
rect 407 8615 421 8629
rect 431 8615 445 8629
rect 455 8615 469 8629
rect 479 8615 493 8629
rect 503 8615 517 8629
rect 527 8615 541 8629
rect 551 8615 565 8629
rect 575 8615 589 8629
rect 599 8615 613 8629
rect 623 8615 637 8629
rect 647 8615 661 8629
rect 671 8615 685 8629
rect 695 8615 709 8629
rect 719 8615 733 8629
rect 47 8423 61 8437
rect 71 8423 85 8437
rect 95 8423 109 8437
rect 119 8423 133 8437
rect 143 8423 157 8437
rect 167 8423 181 8437
rect 191 8423 205 8437
rect 215 8423 229 8437
rect 239 8423 253 8437
rect 263 8423 277 8437
rect 287 8423 301 8437
rect 311 8423 325 8437
rect 335 8423 349 8437
rect 359 8423 373 8437
rect 383 8423 397 8437
rect 407 8423 421 8437
rect 431 8423 445 8437
rect 455 8423 469 8437
rect 479 8423 493 8437
rect 503 8423 517 8437
rect 527 8423 541 8437
rect 551 8423 565 8437
rect 575 8423 589 8437
rect 599 8423 613 8437
rect 623 8423 637 8437
rect 647 8423 661 8437
rect 671 8423 685 8437
rect 695 8423 709 8437
rect 719 8423 733 8437
rect 743 8423 757 8437
rect 47 8375 61 8389
rect 71 8375 85 8389
rect 95 8375 109 8389
rect 119 8375 133 8389
rect 143 8375 157 8389
rect 167 8375 181 8389
rect 191 8375 205 8389
rect 215 8375 229 8389
rect 239 8375 253 8389
rect 263 8375 277 8389
rect 287 8375 301 8389
rect 311 8375 325 8389
rect 335 8375 349 8389
rect 359 8375 373 8389
rect 383 8375 397 8389
rect 407 8375 421 8389
rect 431 8375 445 8389
rect 455 8375 469 8389
rect 479 8375 493 8389
rect 503 8375 517 8389
rect 527 8375 541 8389
rect 551 8375 565 8389
rect 575 8375 589 8389
rect 599 8375 613 8389
rect 623 8375 637 8389
rect 647 8375 661 8389
rect 671 8375 685 8389
rect 695 8375 709 8389
rect 719 8375 733 8389
rect 743 8375 757 8389
rect 47 8183 61 8197
rect 71 8183 85 8197
rect 95 8183 109 8197
rect 119 8183 133 8197
rect 143 8183 157 8197
rect 167 8183 181 8197
rect 191 8183 205 8197
rect 215 8183 229 8197
rect 239 8183 253 8197
rect 263 8183 277 8197
rect 287 8183 301 8197
rect 311 8183 325 8197
rect 335 8183 349 8197
rect 359 8183 373 8197
rect 383 8183 397 8197
rect 407 8183 421 8197
rect 431 8183 445 8197
rect 455 8183 469 8197
rect 479 8183 493 8197
rect 503 8183 517 8197
rect 527 8183 541 8197
rect 551 8183 565 8197
rect 575 8183 589 8197
rect 599 8183 613 8197
rect 623 8183 637 8197
rect 647 8183 661 8197
rect 671 8183 685 8197
rect 695 8183 709 8197
rect 719 8183 733 8197
rect 743 8183 757 8197
rect 767 8183 781 8197
rect 47 8135 61 8149
rect 71 8135 85 8149
rect 95 8135 109 8149
rect 119 8135 133 8149
rect 143 8135 157 8149
rect 167 8135 181 8149
rect 191 8135 205 8149
rect 215 8135 229 8149
rect 239 8135 253 8149
rect 263 8135 277 8149
rect 287 8135 301 8149
rect 311 8135 325 8149
rect 335 8135 349 8149
rect 359 8135 373 8149
rect 383 8135 397 8149
rect 407 8135 421 8149
rect 431 8135 445 8149
rect 455 8135 469 8149
rect 479 8135 493 8149
rect 503 8135 517 8149
rect 527 8135 541 8149
rect 551 8135 565 8149
rect 575 8135 589 8149
rect 599 8135 613 8149
rect 623 8135 637 8149
rect 647 8135 661 8149
rect 671 8135 685 8149
rect 695 8135 709 8149
rect 719 8135 733 8149
rect 743 8135 757 8149
rect 767 8135 781 8149
rect 47 7943 61 7957
rect 71 7943 85 7957
rect 95 7943 109 7957
rect 119 7943 133 7957
rect 143 7943 157 7957
rect 167 7943 181 7957
rect 191 7943 205 7957
rect 215 7943 229 7957
rect 239 7943 253 7957
rect 263 7943 277 7957
rect 287 7943 301 7957
rect 311 7943 325 7957
rect 335 7943 349 7957
rect 359 7943 373 7957
rect 383 7943 397 7957
rect 407 7943 421 7957
rect 431 7943 445 7957
rect 455 7943 469 7957
rect 479 7943 493 7957
rect 503 7943 517 7957
rect 527 7943 541 7957
rect 551 7943 565 7957
rect 575 7943 589 7957
rect 599 7943 613 7957
rect 623 7943 637 7957
rect 647 7943 661 7957
rect 671 7943 685 7957
rect 695 7943 709 7957
rect 719 7943 733 7957
rect 743 7943 757 7957
rect 767 7943 781 7957
rect 791 7943 805 7957
rect 47 7895 61 7909
rect 71 7895 85 7909
rect 95 7895 109 7909
rect 119 7895 133 7909
rect 143 7895 157 7909
rect 167 7895 181 7909
rect 191 7895 205 7909
rect 215 7895 229 7909
rect 239 7895 253 7909
rect 263 7895 277 7909
rect 287 7895 301 7909
rect 311 7895 325 7909
rect 335 7895 349 7909
rect 359 7895 373 7909
rect 383 7895 397 7909
rect 407 7895 421 7909
rect 431 7895 445 7909
rect 455 7895 469 7909
rect 479 7895 493 7909
rect 503 7895 517 7909
rect 527 7895 541 7909
rect 551 7895 565 7909
rect 575 7895 589 7909
rect 599 7895 613 7909
rect 623 7895 637 7909
rect 647 7895 661 7909
rect 671 7895 685 7909
rect 695 7895 709 7909
rect 719 7895 733 7909
rect 743 7895 757 7909
rect 767 7895 781 7909
rect 791 7895 805 7909
rect 47 7703 61 7717
rect 71 7703 85 7717
rect 95 7703 109 7717
rect 119 7703 133 7717
rect 143 7703 157 7717
rect 167 7703 181 7717
rect 191 7703 205 7717
rect 215 7703 229 7717
rect 239 7703 253 7717
rect 263 7703 277 7717
rect 287 7703 301 7717
rect 311 7703 325 7717
rect 335 7703 349 7717
rect 359 7703 373 7717
rect 383 7703 397 7717
rect 407 7703 421 7717
rect 431 7703 445 7717
rect 455 7703 469 7717
rect 479 7703 493 7717
rect 503 7703 517 7717
rect 527 7703 541 7717
rect 551 7703 565 7717
rect 575 7703 589 7717
rect 599 7703 613 7717
rect 623 7703 637 7717
rect 647 7703 661 7717
rect 671 7703 685 7717
rect 695 7703 709 7717
rect 719 7703 733 7717
rect 743 7703 757 7717
rect 767 7703 781 7717
rect 791 7703 805 7717
rect 815 7703 829 7717
rect 47 7655 61 7669
rect 71 7655 85 7669
rect 95 7655 109 7669
rect 119 7655 133 7669
rect 143 7655 157 7669
rect 167 7655 181 7669
rect 191 7655 205 7669
rect 215 7655 229 7669
rect 239 7655 253 7669
rect 263 7655 277 7669
rect 287 7655 301 7669
rect 311 7655 325 7669
rect 335 7655 349 7669
rect 359 7655 373 7669
rect 383 7655 397 7669
rect 407 7655 421 7669
rect 431 7655 445 7669
rect 455 7655 469 7669
rect 479 7655 493 7669
rect 503 7655 517 7669
rect 527 7655 541 7669
rect 551 7655 565 7669
rect 575 7655 589 7669
rect 599 7655 613 7669
rect 623 7655 637 7669
rect 647 7655 661 7669
rect 671 7655 685 7669
rect 695 7655 709 7669
rect 719 7655 733 7669
rect 743 7655 757 7669
rect 767 7655 781 7669
rect 791 7655 805 7669
rect 815 7655 829 7669
rect 47 7463 61 7477
rect 71 7463 85 7477
rect 95 7463 109 7477
rect 119 7463 133 7477
rect 143 7463 157 7477
rect 167 7463 181 7477
rect 191 7463 205 7477
rect 215 7463 229 7477
rect 239 7463 253 7477
rect 263 7463 277 7477
rect 287 7463 301 7477
rect 311 7463 325 7477
rect 335 7463 349 7477
rect 359 7463 373 7477
rect 383 7463 397 7477
rect 407 7463 421 7477
rect 431 7463 445 7477
rect 455 7463 469 7477
rect 479 7463 493 7477
rect 503 7463 517 7477
rect 527 7463 541 7477
rect 551 7463 565 7477
rect 575 7463 589 7477
rect 599 7463 613 7477
rect 623 7463 637 7477
rect 647 7463 661 7477
rect 671 7463 685 7477
rect 695 7463 709 7477
rect 719 7463 733 7477
rect 743 7463 757 7477
rect 767 7463 781 7477
rect 791 7463 805 7477
rect 815 7463 829 7477
rect 839 7463 853 7477
rect 47 7415 61 7429
rect 71 7415 85 7429
rect 95 7415 109 7429
rect 119 7415 133 7429
rect 143 7415 157 7429
rect 167 7415 181 7429
rect 191 7415 205 7429
rect 215 7415 229 7429
rect 239 7415 253 7429
rect 263 7415 277 7429
rect 287 7415 301 7429
rect 311 7415 325 7429
rect 335 7415 349 7429
rect 359 7415 373 7429
rect 383 7415 397 7429
rect 407 7415 421 7429
rect 431 7415 445 7429
rect 455 7415 469 7429
rect 479 7415 493 7429
rect 503 7415 517 7429
rect 527 7415 541 7429
rect 551 7415 565 7429
rect 575 7415 589 7429
rect 599 7415 613 7429
rect 623 7415 637 7429
rect 647 7415 661 7429
rect 671 7415 685 7429
rect 695 7415 709 7429
rect 719 7415 733 7429
rect 743 7415 757 7429
rect 767 7415 781 7429
rect 791 7415 805 7429
rect 815 7415 829 7429
rect 839 7415 853 7429
rect 47 7223 61 7237
rect 71 7223 85 7237
rect 95 7223 109 7237
rect 119 7223 133 7237
rect 143 7223 157 7237
rect 167 7223 181 7237
rect 191 7223 205 7237
rect 215 7223 229 7237
rect 239 7223 253 7237
rect 263 7223 277 7237
rect 287 7223 301 7237
rect 311 7223 325 7237
rect 335 7223 349 7237
rect 359 7223 373 7237
rect 383 7223 397 7237
rect 407 7223 421 7237
rect 431 7223 445 7237
rect 455 7223 469 7237
rect 479 7223 493 7237
rect 503 7223 517 7237
rect 527 7223 541 7237
rect 551 7223 565 7237
rect 575 7223 589 7237
rect 599 7223 613 7237
rect 623 7223 637 7237
rect 647 7223 661 7237
rect 671 7223 685 7237
rect 695 7223 709 7237
rect 719 7223 733 7237
rect 743 7223 757 7237
rect 767 7223 781 7237
rect 791 7223 805 7237
rect 815 7223 829 7237
rect 839 7223 853 7237
rect 863 7223 877 7237
rect 47 7175 61 7189
rect 71 7175 85 7189
rect 95 7175 109 7189
rect 119 7175 133 7189
rect 143 7175 157 7189
rect 167 7175 181 7189
rect 191 7175 205 7189
rect 215 7175 229 7189
rect 239 7175 253 7189
rect 263 7175 277 7189
rect 287 7175 301 7189
rect 311 7175 325 7189
rect 335 7175 349 7189
rect 359 7175 373 7189
rect 383 7175 397 7189
rect 407 7175 421 7189
rect 431 7175 445 7189
rect 455 7175 469 7189
rect 479 7175 493 7189
rect 503 7175 517 7189
rect 527 7175 541 7189
rect 551 7175 565 7189
rect 575 7175 589 7189
rect 599 7175 613 7189
rect 623 7175 637 7189
rect 647 7175 661 7189
rect 671 7175 685 7189
rect 695 7175 709 7189
rect 719 7175 733 7189
rect 743 7175 757 7189
rect 767 7175 781 7189
rect 791 7175 805 7189
rect 815 7175 829 7189
rect 839 7175 853 7189
rect 863 7175 877 7189
rect 47 6983 61 6997
rect 71 6983 85 6997
rect 95 6983 109 6997
rect 119 6983 133 6997
rect 143 6983 157 6997
rect 167 6983 181 6997
rect 191 6983 205 6997
rect 215 6983 229 6997
rect 239 6983 253 6997
rect 263 6983 277 6997
rect 287 6983 301 6997
rect 311 6983 325 6997
rect 335 6983 349 6997
rect 359 6983 373 6997
rect 383 6983 397 6997
rect 407 6983 421 6997
rect 431 6983 445 6997
rect 455 6983 469 6997
rect 479 6983 493 6997
rect 503 6983 517 6997
rect 527 6983 541 6997
rect 551 6983 565 6997
rect 575 6983 589 6997
rect 599 6983 613 6997
rect 623 6983 637 6997
rect 647 6983 661 6997
rect 671 6983 685 6997
rect 695 6983 709 6997
rect 719 6983 733 6997
rect 743 6983 757 6997
rect 767 6983 781 6997
rect 791 6983 805 6997
rect 815 6983 829 6997
rect 839 6983 853 6997
rect 863 6983 877 6997
rect 887 6983 901 6997
rect 47 6935 61 6949
rect 71 6935 85 6949
rect 95 6935 109 6949
rect 119 6935 133 6949
rect 143 6935 157 6949
rect 167 6935 181 6949
rect 191 6935 205 6949
rect 215 6935 229 6949
rect 239 6935 253 6949
rect 263 6935 277 6949
rect 287 6935 301 6949
rect 311 6935 325 6949
rect 335 6935 349 6949
rect 359 6935 373 6949
rect 383 6935 397 6949
rect 407 6935 421 6949
rect 431 6935 445 6949
rect 455 6935 469 6949
rect 479 6935 493 6949
rect 503 6935 517 6949
rect 527 6935 541 6949
rect 551 6935 565 6949
rect 575 6935 589 6949
rect 599 6935 613 6949
rect 623 6935 637 6949
rect 647 6935 661 6949
rect 671 6935 685 6949
rect 695 6935 709 6949
rect 719 6935 733 6949
rect 743 6935 757 6949
rect 767 6935 781 6949
rect 791 6935 805 6949
rect 815 6935 829 6949
rect 839 6935 853 6949
rect 863 6935 877 6949
rect 887 6935 901 6949
rect 47 6743 61 6757
rect 71 6743 85 6757
rect 95 6743 109 6757
rect 119 6743 133 6757
rect 143 6743 157 6757
rect 167 6743 181 6757
rect 191 6743 205 6757
rect 215 6743 229 6757
rect 239 6743 253 6757
rect 263 6743 277 6757
rect 287 6743 301 6757
rect 311 6743 325 6757
rect 335 6743 349 6757
rect 359 6743 373 6757
rect 383 6743 397 6757
rect 407 6743 421 6757
rect 431 6743 445 6757
rect 455 6743 469 6757
rect 479 6743 493 6757
rect 503 6743 517 6757
rect 527 6743 541 6757
rect 551 6743 565 6757
rect 575 6743 589 6757
rect 599 6743 613 6757
rect 623 6743 637 6757
rect 647 6743 661 6757
rect 671 6743 685 6757
rect 695 6743 709 6757
rect 719 6743 733 6757
rect 743 6743 757 6757
rect 767 6743 781 6757
rect 791 6743 805 6757
rect 815 6743 829 6757
rect 839 6743 853 6757
rect 863 6743 877 6757
rect 887 6743 901 6757
rect 911 6743 925 6757
rect 47 6695 61 6709
rect 71 6695 85 6709
rect 95 6695 109 6709
rect 119 6695 133 6709
rect 143 6695 157 6709
rect 167 6695 181 6709
rect 191 6695 205 6709
rect 215 6695 229 6709
rect 239 6695 253 6709
rect 263 6695 277 6709
rect 287 6695 301 6709
rect 311 6695 325 6709
rect 335 6695 349 6709
rect 359 6695 373 6709
rect 383 6695 397 6709
rect 407 6695 421 6709
rect 431 6695 445 6709
rect 455 6695 469 6709
rect 479 6695 493 6709
rect 503 6695 517 6709
rect 527 6695 541 6709
rect 551 6695 565 6709
rect 575 6695 589 6709
rect 599 6695 613 6709
rect 623 6695 637 6709
rect 647 6695 661 6709
rect 671 6695 685 6709
rect 695 6695 709 6709
rect 719 6695 733 6709
rect 743 6695 757 6709
rect 767 6695 781 6709
rect 791 6695 805 6709
rect 815 6695 829 6709
rect 839 6695 853 6709
rect 863 6695 877 6709
rect 887 6695 901 6709
rect 911 6695 925 6709
rect 47 6503 61 6517
rect 71 6503 85 6517
rect 95 6503 109 6517
rect 119 6503 133 6517
rect 143 6503 157 6517
rect 167 6503 181 6517
rect 191 6503 205 6517
rect 215 6503 229 6517
rect 239 6503 253 6517
rect 263 6503 277 6517
rect 287 6503 301 6517
rect 311 6503 325 6517
rect 335 6503 349 6517
rect 359 6503 373 6517
rect 383 6503 397 6517
rect 407 6503 421 6517
rect 431 6503 445 6517
rect 455 6503 469 6517
rect 479 6503 493 6517
rect 503 6503 517 6517
rect 527 6503 541 6517
rect 551 6503 565 6517
rect 575 6503 589 6517
rect 599 6503 613 6517
rect 623 6503 637 6517
rect 647 6503 661 6517
rect 671 6503 685 6517
rect 695 6503 709 6517
rect 719 6503 733 6517
rect 743 6503 757 6517
rect 767 6503 781 6517
rect 791 6503 805 6517
rect 815 6503 829 6517
rect 839 6503 853 6517
rect 863 6503 877 6517
rect 887 6503 901 6517
rect 911 6503 925 6517
rect 935 6503 949 6517
rect 47 6455 61 6469
rect 71 6455 85 6469
rect 95 6455 109 6469
rect 119 6455 133 6469
rect 143 6455 157 6469
rect 167 6455 181 6469
rect 191 6455 205 6469
rect 215 6455 229 6469
rect 239 6455 253 6469
rect 263 6455 277 6469
rect 287 6455 301 6469
rect 311 6455 325 6469
rect 335 6455 349 6469
rect 359 6455 373 6469
rect 383 6455 397 6469
rect 407 6455 421 6469
rect 431 6455 445 6469
rect 455 6455 469 6469
rect 479 6455 493 6469
rect 503 6455 517 6469
rect 527 6455 541 6469
rect 551 6455 565 6469
rect 575 6455 589 6469
rect 599 6455 613 6469
rect 623 6455 637 6469
rect 647 6455 661 6469
rect 671 6455 685 6469
rect 695 6455 709 6469
rect 719 6455 733 6469
rect 743 6455 757 6469
rect 767 6455 781 6469
rect 791 6455 805 6469
rect 815 6455 829 6469
rect 839 6455 853 6469
rect 863 6455 877 6469
rect 887 6455 901 6469
rect 911 6455 925 6469
rect 935 6455 949 6469
rect 47 6263 61 6277
rect 71 6263 85 6277
rect 95 6263 109 6277
rect 119 6263 133 6277
rect 143 6263 157 6277
rect 167 6263 181 6277
rect 191 6263 205 6277
rect 215 6263 229 6277
rect 239 6263 253 6277
rect 263 6263 277 6277
rect 287 6263 301 6277
rect 311 6263 325 6277
rect 335 6263 349 6277
rect 359 6263 373 6277
rect 383 6263 397 6277
rect 407 6263 421 6277
rect 431 6263 445 6277
rect 455 6263 469 6277
rect 479 6263 493 6277
rect 503 6263 517 6277
rect 527 6263 541 6277
rect 551 6263 565 6277
rect 575 6263 589 6277
rect 599 6263 613 6277
rect 623 6263 637 6277
rect 647 6263 661 6277
rect 671 6263 685 6277
rect 695 6263 709 6277
rect 719 6263 733 6277
rect 743 6263 757 6277
rect 767 6263 781 6277
rect 791 6263 805 6277
rect 815 6263 829 6277
rect 839 6263 853 6277
rect 863 6263 877 6277
rect 887 6263 901 6277
rect 911 6263 925 6277
rect 935 6263 949 6277
rect 959 6263 973 6277
rect 47 6215 61 6229
rect 71 6215 85 6229
rect 95 6215 109 6229
rect 119 6215 133 6229
rect 143 6215 157 6229
rect 167 6215 181 6229
rect 191 6215 205 6229
rect 215 6215 229 6229
rect 239 6215 253 6229
rect 263 6215 277 6229
rect 287 6215 301 6229
rect 311 6215 325 6229
rect 335 6215 349 6229
rect 359 6215 373 6229
rect 383 6215 397 6229
rect 407 6215 421 6229
rect 431 6215 445 6229
rect 455 6215 469 6229
rect 479 6215 493 6229
rect 503 6215 517 6229
rect 527 6215 541 6229
rect 551 6215 565 6229
rect 575 6215 589 6229
rect 599 6215 613 6229
rect 623 6215 637 6229
rect 647 6215 661 6229
rect 671 6215 685 6229
rect 695 6215 709 6229
rect 719 6215 733 6229
rect 743 6215 757 6229
rect 767 6215 781 6229
rect 791 6215 805 6229
rect 815 6215 829 6229
rect 839 6215 853 6229
rect 863 6215 877 6229
rect 887 6215 901 6229
rect 911 6215 925 6229
rect 935 6215 949 6229
rect 959 6215 973 6229
rect 47 6023 61 6037
rect 71 6023 85 6037
rect 95 6023 109 6037
rect 119 6023 133 6037
rect 143 6023 157 6037
rect 167 6023 181 6037
rect 191 6023 205 6037
rect 215 6023 229 6037
rect 239 6023 253 6037
rect 263 6023 277 6037
rect 287 6023 301 6037
rect 311 6023 325 6037
rect 335 6023 349 6037
rect 359 6023 373 6037
rect 383 6023 397 6037
rect 407 6023 421 6037
rect 431 6023 445 6037
rect 455 6023 469 6037
rect 479 6023 493 6037
rect 503 6023 517 6037
rect 527 6023 541 6037
rect 551 6023 565 6037
rect 575 6023 589 6037
rect 599 6023 613 6037
rect 623 6023 637 6037
rect 647 6023 661 6037
rect 671 6023 685 6037
rect 695 6023 709 6037
rect 719 6023 733 6037
rect 743 6023 757 6037
rect 767 6023 781 6037
rect 791 6023 805 6037
rect 815 6023 829 6037
rect 839 6023 853 6037
rect 863 6023 877 6037
rect 887 6023 901 6037
rect 911 6023 925 6037
rect 935 6023 949 6037
rect 959 6023 973 6037
rect 983 6023 997 6037
rect 47 5975 61 5989
rect 71 5975 85 5989
rect 95 5975 109 5989
rect 119 5975 133 5989
rect 143 5975 157 5989
rect 167 5975 181 5989
rect 191 5975 205 5989
rect 215 5975 229 5989
rect 239 5975 253 5989
rect 263 5975 277 5989
rect 287 5975 301 5989
rect 311 5975 325 5989
rect 335 5975 349 5989
rect 359 5975 373 5989
rect 383 5975 397 5989
rect 407 5975 421 5989
rect 431 5975 445 5989
rect 455 5975 469 5989
rect 479 5975 493 5989
rect 503 5975 517 5989
rect 527 5975 541 5989
rect 551 5975 565 5989
rect 575 5975 589 5989
rect 599 5975 613 5989
rect 623 5975 637 5989
rect 647 5975 661 5989
rect 671 5975 685 5989
rect 695 5975 709 5989
rect 719 5975 733 5989
rect 743 5975 757 5989
rect 767 5975 781 5989
rect 791 5975 805 5989
rect 815 5975 829 5989
rect 839 5975 853 5989
rect 863 5975 877 5989
rect 887 5975 901 5989
rect 911 5975 925 5989
rect 935 5975 949 5989
rect 959 5975 973 5989
rect 983 5975 997 5989
rect 47 5783 61 5797
rect 71 5783 85 5797
rect 95 5783 109 5797
rect 119 5783 133 5797
rect 143 5783 157 5797
rect 167 5783 181 5797
rect 191 5783 205 5797
rect 215 5783 229 5797
rect 239 5783 253 5797
rect 263 5783 277 5797
rect 287 5783 301 5797
rect 311 5783 325 5797
rect 335 5783 349 5797
rect 359 5783 373 5797
rect 383 5783 397 5797
rect 407 5783 421 5797
rect 431 5783 445 5797
rect 455 5783 469 5797
rect 479 5783 493 5797
rect 503 5783 517 5797
rect 527 5783 541 5797
rect 551 5783 565 5797
rect 575 5783 589 5797
rect 599 5783 613 5797
rect 623 5783 637 5797
rect 647 5783 661 5797
rect 671 5783 685 5797
rect 695 5783 709 5797
rect 719 5783 733 5797
rect 743 5783 757 5797
rect 767 5783 781 5797
rect 791 5783 805 5797
rect 815 5783 829 5797
rect 839 5783 853 5797
rect 863 5783 877 5797
rect 887 5783 901 5797
rect 911 5783 925 5797
rect 935 5783 949 5797
rect 959 5783 973 5797
rect 983 5783 997 5797
rect 1007 5783 1021 5797
rect 47 5735 61 5749
rect 71 5735 85 5749
rect 95 5735 109 5749
rect 119 5735 133 5749
rect 143 5735 157 5749
rect 167 5735 181 5749
rect 191 5735 205 5749
rect 215 5735 229 5749
rect 239 5735 253 5749
rect 263 5735 277 5749
rect 287 5735 301 5749
rect 311 5735 325 5749
rect 335 5735 349 5749
rect 359 5735 373 5749
rect 383 5735 397 5749
rect 407 5735 421 5749
rect 431 5735 445 5749
rect 455 5735 469 5749
rect 479 5735 493 5749
rect 503 5735 517 5749
rect 527 5735 541 5749
rect 551 5735 565 5749
rect 575 5735 589 5749
rect 599 5735 613 5749
rect 623 5735 637 5749
rect 647 5735 661 5749
rect 671 5735 685 5749
rect 695 5735 709 5749
rect 719 5735 733 5749
rect 743 5735 757 5749
rect 767 5735 781 5749
rect 791 5735 805 5749
rect 815 5735 829 5749
rect 839 5735 853 5749
rect 863 5735 877 5749
rect 887 5735 901 5749
rect 911 5735 925 5749
rect 935 5735 949 5749
rect 959 5735 973 5749
rect 983 5735 997 5749
rect 1007 5735 1021 5749
rect 47 5543 61 5557
rect 71 5543 85 5557
rect 95 5543 109 5557
rect 119 5543 133 5557
rect 143 5543 157 5557
rect 167 5543 181 5557
rect 191 5543 205 5557
rect 215 5543 229 5557
rect 239 5543 253 5557
rect 263 5543 277 5557
rect 287 5543 301 5557
rect 311 5543 325 5557
rect 335 5543 349 5557
rect 359 5543 373 5557
rect 383 5543 397 5557
rect 407 5543 421 5557
rect 431 5543 445 5557
rect 455 5543 469 5557
rect 479 5543 493 5557
rect 503 5543 517 5557
rect 527 5543 541 5557
rect 551 5543 565 5557
rect 575 5543 589 5557
rect 599 5543 613 5557
rect 623 5543 637 5557
rect 647 5543 661 5557
rect 671 5543 685 5557
rect 695 5543 709 5557
rect 719 5543 733 5557
rect 743 5543 757 5557
rect 767 5543 781 5557
rect 791 5543 805 5557
rect 815 5543 829 5557
rect 839 5543 853 5557
rect 863 5543 877 5557
rect 887 5543 901 5557
rect 911 5543 925 5557
rect 935 5543 949 5557
rect 959 5543 973 5557
rect 983 5543 997 5557
rect 1007 5543 1021 5557
rect 1031 5543 1045 5557
rect 47 5495 61 5509
rect 71 5495 85 5509
rect 95 5495 109 5509
rect 119 5495 133 5509
rect 143 5495 157 5509
rect 167 5495 181 5509
rect 191 5495 205 5509
rect 215 5495 229 5509
rect 239 5495 253 5509
rect 263 5495 277 5509
rect 287 5495 301 5509
rect 311 5495 325 5509
rect 335 5495 349 5509
rect 359 5495 373 5509
rect 383 5495 397 5509
rect 407 5495 421 5509
rect 431 5495 445 5509
rect 455 5495 469 5509
rect 479 5495 493 5509
rect 503 5495 517 5509
rect 527 5495 541 5509
rect 551 5495 565 5509
rect 575 5495 589 5509
rect 599 5495 613 5509
rect 623 5495 637 5509
rect 647 5495 661 5509
rect 671 5495 685 5509
rect 695 5495 709 5509
rect 719 5495 733 5509
rect 743 5495 757 5509
rect 767 5495 781 5509
rect 791 5495 805 5509
rect 815 5495 829 5509
rect 839 5495 853 5509
rect 863 5495 877 5509
rect 887 5495 901 5509
rect 911 5495 925 5509
rect 935 5495 949 5509
rect 959 5495 973 5509
rect 983 5495 997 5509
rect 1007 5495 1021 5509
rect 1031 5495 1045 5509
rect 47 5303 61 5317
rect 71 5303 85 5317
rect 95 5303 109 5317
rect 119 5303 133 5317
rect 143 5303 157 5317
rect 167 5303 181 5317
rect 191 5303 205 5317
rect 215 5303 229 5317
rect 239 5303 253 5317
rect 263 5303 277 5317
rect 287 5303 301 5317
rect 311 5303 325 5317
rect 335 5303 349 5317
rect 359 5303 373 5317
rect 383 5303 397 5317
rect 407 5303 421 5317
rect 431 5303 445 5317
rect 455 5303 469 5317
rect 479 5303 493 5317
rect 503 5303 517 5317
rect 527 5303 541 5317
rect 551 5303 565 5317
rect 575 5303 589 5317
rect 599 5303 613 5317
rect 623 5303 637 5317
rect 647 5303 661 5317
rect 671 5303 685 5317
rect 695 5303 709 5317
rect 719 5303 733 5317
rect 743 5303 757 5317
rect 767 5303 781 5317
rect 791 5303 805 5317
rect 815 5303 829 5317
rect 839 5303 853 5317
rect 863 5303 877 5317
rect 887 5303 901 5317
rect 911 5303 925 5317
rect 935 5303 949 5317
rect 959 5303 973 5317
rect 983 5303 997 5317
rect 1007 5303 1021 5317
rect 1031 5303 1045 5317
rect 1055 5303 1069 5317
rect 47 5255 61 5269
rect 71 5255 85 5269
rect 95 5255 109 5269
rect 119 5255 133 5269
rect 143 5255 157 5269
rect 167 5255 181 5269
rect 191 5255 205 5269
rect 215 5255 229 5269
rect 239 5255 253 5269
rect 263 5255 277 5269
rect 287 5255 301 5269
rect 311 5255 325 5269
rect 335 5255 349 5269
rect 359 5255 373 5269
rect 383 5255 397 5269
rect 407 5255 421 5269
rect 431 5255 445 5269
rect 455 5255 469 5269
rect 479 5255 493 5269
rect 503 5255 517 5269
rect 527 5255 541 5269
rect 551 5255 565 5269
rect 575 5255 589 5269
rect 599 5255 613 5269
rect 623 5255 637 5269
rect 647 5255 661 5269
rect 671 5255 685 5269
rect 695 5255 709 5269
rect 719 5255 733 5269
rect 743 5255 757 5269
rect 767 5255 781 5269
rect 791 5255 805 5269
rect 815 5255 829 5269
rect 839 5255 853 5269
rect 863 5255 877 5269
rect 887 5255 901 5269
rect 911 5255 925 5269
rect 935 5255 949 5269
rect 959 5255 973 5269
rect 983 5255 997 5269
rect 1007 5255 1021 5269
rect 1031 5255 1045 5269
rect 1055 5255 1069 5269
rect 47 5063 61 5077
rect 71 5063 85 5077
rect 95 5063 109 5077
rect 119 5063 133 5077
rect 143 5063 157 5077
rect 167 5063 181 5077
rect 191 5063 205 5077
rect 215 5063 229 5077
rect 239 5063 253 5077
rect 263 5063 277 5077
rect 287 5063 301 5077
rect 311 5063 325 5077
rect 335 5063 349 5077
rect 359 5063 373 5077
rect 383 5063 397 5077
rect 407 5063 421 5077
rect 431 5063 445 5077
rect 455 5063 469 5077
rect 479 5063 493 5077
rect 503 5063 517 5077
rect 527 5063 541 5077
rect 551 5063 565 5077
rect 575 5063 589 5077
rect 599 5063 613 5077
rect 623 5063 637 5077
rect 647 5063 661 5077
rect 671 5063 685 5077
rect 695 5063 709 5077
rect 719 5063 733 5077
rect 743 5063 757 5077
rect 767 5063 781 5077
rect 791 5063 805 5077
rect 815 5063 829 5077
rect 839 5063 853 5077
rect 863 5063 877 5077
rect 887 5063 901 5077
rect 911 5063 925 5077
rect 935 5063 949 5077
rect 959 5063 973 5077
rect 983 5063 997 5077
rect 1007 5063 1021 5077
rect 1031 5063 1045 5077
rect 1055 5063 1069 5077
rect 1079 5063 1093 5077
rect 47 5015 61 5029
rect 71 5015 85 5029
rect 95 5015 109 5029
rect 119 5015 133 5029
rect 143 5015 157 5029
rect 167 5015 181 5029
rect 191 5015 205 5029
rect 215 5015 229 5029
rect 239 5015 253 5029
rect 263 5015 277 5029
rect 287 5015 301 5029
rect 311 5015 325 5029
rect 335 5015 349 5029
rect 359 5015 373 5029
rect 383 5015 397 5029
rect 407 5015 421 5029
rect 431 5015 445 5029
rect 455 5015 469 5029
rect 479 5015 493 5029
rect 503 5015 517 5029
rect 527 5015 541 5029
rect 551 5015 565 5029
rect 575 5015 589 5029
rect 599 5015 613 5029
rect 623 5015 637 5029
rect 647 5015 661 5029
rect 671 5015 685 5029
rect 695 5015 709 5029
rect 719 5015 733 5029
rect 743 5015 757 5029
rect 767 5015 781 5029
rect 791 5015 805 5029
rect 815 5015 829 5029
rect 839 5015 853 5029
rect 863 5015 877 5029
rect 887 5015 901 5029
rect 911 5015 925 5029
rect 935 5015 949 5029
rect 959 5015 973 5029
rect 983 5015 997 5029
rect 1007 5015 1021 5029
rect 1031 5015 1045 5029
rect 1055 5015 1069 5029
rect 1079 5015 1093 5029
rect 47 4823 61 4837
rect 71 4823 85 4837
rect 95 4823 109 4837
rect 119 4823 133 4837
rect 143 4823 157 4837
rect 167 4823 181 4837
rect 191 4823 205 4837
rect 215 4823 229 4837
rect 239 4823 253 4837
rect 263 4823 277 4837
rect 287 4823 301 4837
rect 311 4823 325 4837
rect 335 4823 349 4837
rect 359 4823 373 4837
rect 383 4823 397 4837
rect 407 4823 421 4837
rect 431 4823 445 4837
rect 455 4823 469 4837
rect 479 4823 493 4837
rect 503 4823 517 4837
rect 527 4823 541 4837
rect 551 4823 565 4837
rect 575 4823 589 4837
rect 599 4823 613 4837
rect 623 4823 637 4837
rect 647 4823 661 4837
rect 671 4823 685 4837
rect 695 4823 709 4837
rect 719 4823 733 4837
rect 743 4823 757 4837
rect 767 4823 781 4837
rect 791 4823 805 4837
rect 815 4823 829 4837
rect 839 4823 853 4837
rect 863 4823 877 4837
rect 887 4823 901 4837
rect 911 4823 925 4837
rect 935 4823 949 4837
rect 959 4823 973 4837
rect 983 4823 997 4837
rect 1007 4823 1021 4837
rect 1031 4823 1045 4837
rect 1055 4823 1069 4837
rect 1079 4823 1093 4837
rect 1103 4823 1117 4837
rect 47 4775 61 4789
rect 71 4775 85 4789
rect 95 4775 109 4789
rect 119 4775 133 4789
rect 143 4775 157 4789
rect 167 4775 181 4789
rect 191 4775 205 4789
rect 215 4775 229 4789
rect 239 4775 253 4789
rect 263 4775 277 4789
rect 287 4775 301 4789
rect 311 4775 325 4789
rect 335 4775 349 4789
rect 359 4775 373 4789
rect 383 4775 397 4789
rect 407 4775 421 4789
rect 431 4775 445 4789
rect 455 4775 469 4789
rect 479 4775 493 4789
rect 503 4775 517 4789
rect 527 4775 541 4789
rect 551 4775 565 4789
rect 575 4775 589 4789
rect 599 4775 613 4789
rect 623 4775 637 4789
rect 647 4775 661 4789
rect 671 4775 685 4789
rect 695 4775 709 4789
rect 719 4775 733 4789
rect 743 4775 757 4789
rect 767 4775 781 4789
rect 791 4775 805 4789
rect 815 4775 829 4789
rect 839 4775 853 4789
rect 863 4775 877 4789
rect 887 4775 901 4789
rect 911 4775 925 4789
rect 935 4775 949 4789
rect 959 4775 973 4789
rect 983 4775 997 4789
rect 1007 4775 1021 4789
rect 1031 4775 1045 4789
rect 1055 4775 1069 4789
rect 1079 4775 1093 4789
rect 1103 4775 1117 4789
rect 47 4583 61 4597
rect 71 4583 85 4597
rect 95 4583 109 4597
rect 119 4583 133 4597
rect 143 4583 157 4597
rect 167 4583 181 4597
rect 191 4583 205 4597
rect 215 4583 229 4597
rect 239 4583 253 4597
rect 263 4583 277 4597
rect 287 4583 301 4597
rect 311 4583 325 4597
rect 335 4583 349 4597
rect 359 4583 373 4597
rect 383 4583 397 4597
rect 407 4583 421 4597
rect 431 4583 445 4597
rect 455 4583 469 4597
rect 479 4583 493 4597
rect 503 4583 517 4597
rect 527 4583 541 4597
rect 551 4583 565 4597
rect 575 4583 589 4597
rect 599 4583 613 4597
rect 623 4583 637 4597
rect 647 4583 661 4597
rect 671 4583 685 4597
rect 695 4583 709 4597
rect 719 4583 733 4597
rect 743 4583 757 4597
rect 767 4583 781 4597
rect 791 4583 805 4597
rect 815 4583 829 4597
rect 839 4583 853 4597
rect 863 4583 877 4597
rect 887 4583 901 4597
rect 911 4583 925 4597
rect 935 4583 949 4597
rect 959 4583 973 4597
rect 983 4583 997 4597
rect 1007 4583 1021 4597
rect 1031 4583 1045 4597
rect 1055 4583 1069 4597
rect 1079 4583 1093 4597
rect 1103 4583 1117 4597
rect 1127 4583 1141 4597
rect 47 4535 61 4549
rect 71 4535 85 4549
rect 95 4535 109 4549
rect 119 4535 133 4549
rect 143 4535 157 4549
rect 167 4535 181 4549
rect 191 4535 205 4549
rect 215 4535 229 4549
rect 239 4535 253 4549
rect 263 4535 277 4549
rect 287 4535 301 4549
rect 311 4535 325 4549
rect 335 4535 349 4549
rect 359 4535 373 4549
rect 383 4535 397 4549
rect 407 4535 421 4549
rect 431 4535 445 4549
rect 455 4535 469 4549
rect 479 4535 493 4549
rect 503 4535 517 4549
rect 527 4535 541 4549
rect 551 4535 565 4549
rect 575 4535 589 4549
rect 599 4535 613 4549
rect 623 4535 637 4549
rect 647 4535 661 4549
rect 671 4535 685 4549
rect 695 4535 709 4549
rect 719 4535 733 4549
rect 743 4535 757 4549
rect 767 4535 781 4549
rect 791 4535 805 4549
rect 815 4535 829 4549
rect 839 4535 853 4549
rect 863 4535 877 4549
rect 887 4535 901 4549
rect 911 4535 925 4549
rect 935 4535 949 4549
rect 959 4535 973 4549
rect 983 4535 997 4549
rect 1007 4535 1021 4549
rect 1031 4535 1045 4549
rect 1055 4535 1069 4549
rect 1079 4535 1093 4549
rect 1103 4535 1117 4549
rect 1127 4535 1141 4549
rect 47 4343 61 4357
rect 71 4343 85 4357
rect 95 4343 109 4357
rect 119 4343 133 4357
rect 143 4343 157 4357
rect 167 4343 181 4357
rect 191 4343 205 4357
rect 215 4343 229 4357
rect 239 4343 253 4357
rect 263 4343 277 4357
rect 287 4343 301 4357
rect 311 4343 325 4357
rect 335 4343 349 4357
rect 359 4343 373 4357
rect 383 4343 397 4357
rect 407 4343 421 4357
rect 431 4343 445 4357
rect 455 4343 469 4357
rect 479 4343 493 4357
rect 503 4343 517 4357
rect 527 4343 541 4357
rect 551 4343 565 4357
rect 575 4343 589 4357
rect 599 4343 613 4357
rect 623 4343 637 4357
rect 647 4343 661 4357
rect 671 4343 685 4357
rect 695 4343 709 4357
rect 719 4343 733 4357
rect 743 4343 757 4357
rect 767 4343 781 4357
rect 791 4343 805 4357
rect 815 4343 829 4357
rect 839 4343 853 4357
rect 863 4343 877 4357
rect 887 4343 901 4357
rect 911 4343 925 4357
rect 935 4343 949 4357
rect 959 4343 973 4357
rect 983 4343 997 4357
rect 1007 4343 1021 4357
rect 1031 4343 1045 4357
rect 1055 4343 1069 4357
rect 1079 4343 1093 4357
rect 1103 4343 1117 4357
rect 1127 4343 1141 4357
rect 1151 4343 1165 4357
rect 47 4295 61 4309
rect 71 4295 85 4309
rect 95 4295 109 4309
rect 119 4295 133 4309
rect 143 4295 157 4309
rect 167 4295 181 4309
rect 191 4295 205 4309
rect 215 4295 229 4309
rect 239 4295 253 4309
rect 263 4295 277 4309
rect 287 4295 301 4309
rect 311 4295 325 4309
rect 335 4295 349 4309
rect 359 4295 373 4309
rect 383 4295 397 4309
rect 407 4295 421 4309
rect 431 4295 445 4309
rect 455 4295 469 4309
rect 479 4295 493 4309
rect 503 4295 517 4309
rect 527 4295 541 4309
rect 551 4295 565 4309
rect 575 4295 589 4309
rect 599 4295 613 4309
rect 623 4295 637 4309
rect 647 4295 661 4309
rect 671 4295 685 4309
rect 695 4295 709 4309
rect 719 4295 733 4309
rect 743 4295 757 4309
rect 767 4295 781 4309
rect 791 4295 805 4309
rect 815 4295 829 4309
rect 839 4295 853 4309
rect 863 4295 877 4309
rect 887 4295 901 4309
rect 911 4295 925 4309
rect 935 4295 949 4309
rect 959 4295 973 4309
rect 983 4295 997 4309
rect 1007 4295 1021 4309
rect 1031 4295 1045 4309
rect 1055 4295 1069 4309
rect 1079 4295 1093 4309
rect 1103 4295 1117 4309
rect 1127 4295 1141 4309
rect 1151 4295 1165 4309
rect 32447 4295 32461 4309
rect 32519 4295 32533 4309
rect 32759 4295 32773 4309
rect 32807 4295 32821 4309
rect 32855 4295 32869 4309
rect 32927 4295 32941 4309
rect 32975 4295 32989 4309
rect 33047 4295 33061 4309
rect 33071 4295 33085 4309
rect 33143 4295 33157 4309
rect 27623 4271 27637 4285
rect 27671 4271 27685 4285
rect 27911 4271 27925 4285
rect 27959 4271 27973 4285
rect 28007 4271 28021 4285
rect 28055 4271 28069 4285
rect 28103 4271 28117 4285
rect 28151 4271 28165 4285
rect 32351 4271 32365 4285
rect 32399 4271 32413 4285
rect 32423 4271 32437 4285
rect 32615 4271 32629 4285
rect 32663 4271 32677 4285
rect 32711 4271 32725 4285
rect 32735 4271 32749 4285
rect 33287 4271 33301 4285
rect 27599 4247 27613 4261
rect 27767 4247 27781 4261
rect 27815 4247 27829 4261
rect 27863 4247 27877 4261
rect 27887 4247 27901 4261
rect 28271 4247 28285 4261
rect 32327 4247 32341 4261
rect 33407 4247 33421 4261
rect 27575 4223 27589 4237
rect 28367 4223 28381 4237
rect 28415 4223 28429 4237
rect 28463 4223 28477 4237
rect 32303 4223 32317 4237
rect 33503 4223 33517 4237
rect 33551 4223 33565 4237
rect 33599 4223 33613 4237
rect 35399 4223 35413 4237
rect 35447 4223 35461 4237
rect 27047 4199 27061 4213
rect 27095 4199 27109 4213
rect 27263 4199 27277 4213
rect 27311 4199 27325 4213
rect 27335 4199 27349 4213
rect 27431 4199 27445 4213
rect 27479 4199 27493 4213
rect 27527 4199 27541 4213
rect 27551 4199 27565 4213
rect 28559 4199 28573 4213
rect 28607 4199 28621 4213
rect 28655 4199 28669 4213
rect 28703 4199 28717 4213
rect 28751 4199 28765 4213
rect 28775 4199 28789 4213
rect 28847 4199 28861 4213
rect 30479 4199 30493 4213
rect 30551 4199 30565 4213
rect 31991 4199 32005 4213
rect 32039 4199 32053 4213
rect 32087 4199 32101 4213
rect 32135 4199 32149 4213
rect 32159 4199 32173 4213
rect 32231 4199 32245 4213
rect 32279 4199 32293 4213
rect 33695 4199 33709 4213
rect 35375 4199 35389 4213
rect 35567 4199 35581 4213
rect 26903 4175 26917 4189
rect 26975 4175 26989 4189
rect 27023 4175 27037 4189
rect 27215 4175 27229 4189
rect 27239 4175 27253 4189
rect 28943 4175 28957 4189
rect 30263 4175 30277 4189
rect 30311 4175 30325 4189
rect 30335 4175 30349 4189
rect 30407 4175 30421 4189
rect 30455 4175 30469 4189
rect 30671 4175 30685 4189
rect 30695 4175 30709 4189
rect 30791 4175 30805 4189
rect 31967 4175 31981 4189
rect 33815 4175 33829 4189
rect 35255 4175 35269 4189
rect 35327 4175 35341 4189
rect 35351 4175 35365 4189
rect 35663 4175 35677 4189
rect 24575 4151 24589 4165
rect 24623 4151 24637 4165
rect 26471 4151 26485 4165
rect 26519 4151 26533 4165
rect 26807 4151 26821 4165
rect 26855 4151 26869 4165
rect 26879 4151 26893 4165
rect 29039 4151 29053 4165
rect 30023 4151 30037 4165
rect 30095 4151 30109 4165
rect 30143 4151 30157 4165
rect 30191 4151 30205 4165
rect 30239 4151 30253 4165
rect 30911 4151 30925 4165
rect 31871 4151 31885 4165
rect 31919 4151 31933 4165
rect 31943 4151 31957 4165
rect 33935 4151 33949 4165
rect 33959 4151 33973 4165
rect 34031 4151 34045 4165
rect 34055 4151 34069 4165
rect 34127 4151 34141 4165
rect 34151 4151 34165 4165
rect 34223 4151 34237 4165
rect 35135 4151 35149 4165
rect 35207 4151 35221 4165
rect 35231 4151 35245 4165
rect 35759 4151 35773 4165
rect 24551 4127 24565 4141
rect 24719 4127 24733 4141
rect 26447 4127 26461 4141
rect 26615 4127 26629 4141
rect 26663 4127 26677 4141
rect 26735 4127 26749 4141
rect 26759 4127 26773 4141
rect 29135 4127 29149 4141
rect 29999 4127 30013 4141
rect 31031 4127 31045 4141
rect 31463 4127 31477 4141
rect 31511 4127 31525 4141
rect 31559 4127 31573 4141
rect 31607 4127 31621 4141
rect 31775 4127 31789 4141
rect 31823 4127 31837 4141
rect 31847 4127 31861 4141
rect 34343 4127 34357 4141
rect 34847 4127 34861 4141
rect 34895 4127 34909 4141
rect 34919 4127 34933 4141
rect 34991 4127 35005 4141
rect 35015 4127 35029 4141
rect 35087 4127 35101 4141
rect 35111 4127 35125 4141
rect 35855 4127 35869 4141
rect 47 4103 61 4117
rect 71 4103 85 4117
rect 95 4103 109 4117
rect 119 4103 133 4117
rect 143 4103 157 4117
rect 167 4103 181 4117
rect 191 4103 205 4117
rect 215 4103 229 4117
rect 239 4103 253 4117
rect 263 4103 277 4117
rect 287 4103 301 4117
rect 311 4103 325 4117
rect 335 4103 349 4117
rect 359 4103 373 4117
rect 383 4103 397 4117
rect 407 4103 421 4117
rect 431 4103 445 4117
rect 455 4103 469 4117
rect 479 4103 493 4117
rect 503 4103 517 4117
rect 527 4103 541 4117
rect 551 4103 565 4117
rect 575 4103 589 4117
rect 599 4103 613 4117
rect 623 4103 637 4117
rect 647 4103 661 4117
rect 671 4103 685 4117
rect 695 4103 709 4117
rect 719 4103 733 4117
rect 743 4103 757 4117
rect 767 4103 781 4117
rect 791 4103 805 4117
rect 815 4103 829 4117
rect 839 4103 853 4117
rect 863 4103 877 4117
rect 887 4103 901 4117
rect 911 4103 925 4117
rect 935 4103 949 4117
rect 959 4103 973 4117
rect 983 4103 997 4117
rect 1007 4103 1021 4117
rect 1031 4103 1045 4117
rect 1055 4103 1069 4117
rect 1079 4103 1093 4117
rect 1103 4103 1117 4117
rect 1127 4103 1141 4117
rect 1151 4103 1165 4117
rect 1175 4103 1189 4117
rect 24527 4103 24541 4117
rect 24839 4103 24853 4117
rect 24863 4103 24877 4117
rect 24959 4103 24973 4117
rect 25007 4103 25021 4117
rect 25055 4103 25069 4117
rect 26423 4103 26437 4117
rect 29255 4103 29269 4117
rect 29303 4103 29317 4117
rect 29351 4103 29365 4117
rect 29447 4103 29461 4117
rect 31151 4103 31165 4117
rect 31199 4103 31213 4117
rect 31271 4103 31285 4117
rect 31439 4103 31453 4117
rect 31727 4103 31741 4117
rect 31751 4103 31765 4117
rect 34439 4103 34453 4117
rect 34463 4103 34477 4117
rect 34535 4103 34549 4117
rect 34727 4103 34741 4117
rect 34799 4103 34813 4117
rect 34823 4103 34837 4117
rect 35951 4103 35965 4117
rect 35975 4103 35989 4117
rect 36047 4103 36061 4117
rect 47 4055 61 4069
rect 71 4055 85 4069
rect 95 4055 109 4069
rect 119 4055 133 4069
rect 143 4055 157 4069
rect 167 4055 181 4069
rect 191 4055 205 4069
rect 215 4055 229 4069
rect 239 4055 253 4069
rect 263 4055 277 4069
rect 287 4055 301 4069
rect 311 4055 325 4069
rect 335 4055 349 4069
rect 359 4055 373 4069
rect 383 4055 397 4069
rect 407 4055 421 4069
rect 431 4055 445 4069
rect 455 4055 469 4069
rect 479 4055 493 4069
rect 503 4055 517 4069
rect 527 4055 541 4069
rect 551 4055 565 4069
rect 575 4055 589 4069
rect 599 4055 613 4069
rect 623 4055 637 4069
rect 647 4055 661 4069
rect 671 4055 685 4069
rect 695 4055 709 4069
rect 719 4055 733 4069
rect 743 4055 757 4069
rect 767 4055 781 4069
rect 791 4055 805 4069
rect 815 4055 829 4069
rect 839 4055 853 4069
rect 863 4055 877 4069
rect 887 4055 901 4069
rect 911 4055 925 4069
rect 935 4055 949 4069
rect 959 4055 973 4069
rect 983 4055 997 4069
rect 1007 4055 1021 4069
rect 1031 4055 1045 4069
rect 1055 4055 1069 4069
rect 1079 4055 1093 4069
rect 1103 4055 1117 4069
rect 1127 4055 1141 4069
rect 1151 4055 1165 4069
rect 1175 4055 1189 4069
rect 24431 4079 24445 4093
rect 24479 4079 24493 4093
rect 24503 4079 24517 4093
rect 25151 4079 25165 4093
rect 25199 4079 25213 4093
rect 25247 4079 25261 4093
rect 25271 4079 25285 4093
rect 25367 4079 25381 4093
rect 25391 4079 25405 4093
rect 25463 4079 25477 4093
rect 25487 4079 25501 4093
rect 25559 4079 25573 4093
rect 25655 4079 25669 4093
rect 26279 4079 26293 4093
rect 26327 4079 26341 4093
rect 26375 4079 26389 4093
rect 26399 4079 26413 4093
rect 31391 4079 31405 4093
rect 31415 4079 31429 4093
rect 34631 4079 34645 4093
rect 34679 4079 34693 4093
rect 34943 4079 34957 4093
rect 36143 4079 36157 4093
rect 24311 4055 24325 4069
rect 24359 4055 24373 4069
rect 24383 4055 24397 4069
rect 25103 4055 25117 4069
rect 26543 4055 26557 4069
rect 36263 4055 36277 4069
rect 36287 4055 36301 4069
rect 36359 4055 36373 4069
rect 24287 4031 24301 4045
rect 33479 4031 33493 4045
rect 33503 4031 33517 4045
rect 36455 4031 36469 4045
rect 24071 4007 24085 4021
rect 24119 4007 24133 4021
rect 24167 4007 24181 4021
rect 24239 4007 24253 4021
rect 24263 4007 24277 4021
rect 36023 4007 36037 4021
rect 36047 4007 36061 4021
rect 36551 4007 36565 4021
rect 23711 3983 23725 3997
rect 23759 3983 23773 3997
rect 23927 3983 23941 3997
rect 23999 3983 24013 3997
rect 24023 3983 24037 3997
rect 26999 3983 27013 3997
rect 27719 3983 27733 3997
rect 32951 3983 32965 3997
rect 34391 3983 34405 3997
rect 23567 3959 23581 3973
rect 23639 3959 23653 3973
rect 23687 3959 23701 3973
rect 23807 3959 23821 3973
rect 23879 3959 23893 3973
rect 23903 3959 23917 3973
rect 24887 3959 24901 3973
rect 24983 3959 24997 3973
rect 25295 3959 25309 3973
rect 26567 3959 26581 3973
rect 27119 3959 27133 3973
rect 31007 3959 31021 3973
rect 31031 3959 31045 3973
rect 34007 3959 34021 3973
rect 34031 3959 34045 3973
rect 36647 3959 36661 3973
rect 36791 3959 36805 3973
rect 23351 3935 23365 3949
rect 23399 3935 23413 3949
rect 23423 3935 23437 3949
rect 23495 3935 23509 3949
rect 23543 3935 23557 3949
rect 24143 3935 24157 3949
rect 35903 3935 35917 3949
rect 36887 3935 36901 3949
rect 36911 3935 36925 3949
rect 37031 3935 37045 3949
rect 37055 3935 37069 3949
rect 37127 3935 37141 3949
rect 37151 3935 37165 3949
rect 37223 3935 37237 3949
rect 23327 3911 23341 3925
rect 32495 3911 32509 3925
rect 32519 3911 32533 3925
rect 37343 3911 37357 3925
rect 37391 3911 37405 3925
rect 37463 3911 37477 3925
rect 37487 3911 37501 3925
rect 37583 3911 37597 3925
rect 23183 3887 23197 3901
rect 23255 3887 23269 3901
rect 23303 3887 23317 3901
rect 35183 3887 35197 3901
rect 35207 3887 35221 3901
rect 37679 3887 37693 3901
rect 37727 3887 37741 3901
rect 37775 3887 37789 3901
rect 47 3863 61 3877
rect 71 3863 85 3877
rect 95 3863 109 3877
rect 119 3863 133 3877
rect 143 3863 157 3877
rect 167 3863 181 3877
rect 191 3863 205 3877
rect 215 3863 229 3877
rect 239 3863 253 3877
rect 263 3863 277 3877
rect 287 3863 301 3877
rect 311 3863 325 3877
rect 335 3863 349 3877
rect 359 3863 373 3877
rect 383 3863 397 3877
rect 407 3863 421 3877
rect 431 3863 445 3877
rect 455 3863 469 3877
rect 479 3863 493 3877
rect 503 3863 517 3877
rect 527 3863 541 3877
rect 551 3863 565 3877
rect 575 3863 589 3877
rect 599 3863 613 3877
rect 623 3863 637 3877
rect 647 3863 661 3877
rect 671 3863 685 3877
rect 695 3863 709 3877
rect 719 3863 733 3877
rect 743 3863 757 3877
rect 767 3863 781 3877
rect 791 3863 805 3877
rect 815 3863 829 3877
rect 839 3863 853 3877
rect 863 3863 877 3877
rect 887 3863 901 3877
rect 911 3863 925 3877
rect 935 3863 949 3877
rect 959 3863 973 3877
rect 983 3863 997 3877
rect 1007 3863 1021 3877
rect 1031 3863 1045 3877
rect 1055 3863 1069 3877
rect 1079 3863 1093 3877
rect 1103 3863 1117 3877
rect 1127 3863 1141 3877
rect 1151 3863 1165 3877
rect 1175 3863 1189 3877
rect 1199 3863 1213 3877
rect 23159 3863 23173 3877
rect 37823 3863 37837 3877
rect 47 3815 61 3829
rect 71 3815 85 3829
rect 95 3815 109 3829
rect 119 3815 133 3829
rect 143 3815 157 3829
rect 167 3815 181 3829
rect 191 3815 205 3829
rect 215 3815 229 3829
rect 239 3815 253 3829
rect 263 3815 277 3829
rect 287 3815 301 3829
rect 311 3815 325 3829
rect 335 3815 349 3829
rect 359 3815 373 3829
rect 383 3815 397 3829
rect 407 3815 421 3829
rect 431 3815 445 3829
rect 455 3815 469 3829
rect 479 3815 493 3829
rect 503 3815 517 3829
rect 527 3815 541 3829
rect 551 3815 565 3829
rect 575 3815 589 3829
rect 599 3815 613 3829
rect 623 3815 637 3829
rect 647 3815 661 3829
rect 671 3815 685 3829
rect 695 3815 709 3829
rect 719 3815 733 3829
rect 743 3815 757 3829
rect 767 3815 781 3829
rect 791 3815 805 3829
rect 815 3815 829 3829
rect 839 3815 853 3829
rect 863 3815 877 3829
rect 887 3815 901 3829
rect 911 3815 925 3829
rect 935 3815 949 3829
rect 959 3815 973 3829
rect 983 3815 997 3829
rect 1007 3815 1021 3829
rect 1031 3815 1045 3829
rect 1055 3815 1069 3829
rect 1079 3815 1093 3829
rect 1103 3815 1117 3829
rect 1127 3815 1141 3829
rect 1151 3815 1165 3829
rect 1175 3815 1189 3829
rect 1199 3815 1213 3829
rect 23063 3839 23077 3853
rect 23111 3839 23125 3853
rect 23135 3839 23149 3853
rect 37871 3839 37885 3853
rect 37895 3839 37909 3853
rect 37967 3839 37981 3853
rect 22847 3815 22861 3829
rect 22919 3815 22933 3829
rect 22967 3815 22981 3829
rect 23015 3815 23029 3829
rect 23039 3815 23053 3829
rect 29111 3815 29125 3829
rect 29135 3815 29149 3829
rect 38087 3815 38101 3829
rect 38111 3815 38125 3829
rect 38183 3815 38197 3829
rect 22823 3791 22837 3805
rect 38303 3791 38317 3805
rect 22463 3767 22477 3781
rect 22559 3767 22573 3781
rect 22583 3767 22597 3781
rect 22655 3767 22669 3781
rect 22703 3767 22717 3781
rect 22775 3767 22789 3781
rect 22799 3767 22813 3781
rect 38423 3767 38437 3781
rect 22367 3743 22381 3757
rect 22415 3743 22429 3757
rect 22439 3743 22453 3757
rect 33335 3743 33349 3757
rect 38351 3743 38365 3757
rect 38519 3743 38533 3757
rect 22271 3719 22285 3733
rect 22319 3719 22333 3733
rect 22343 3719 22357 3733
rect 27287 3719 27301 3733
rect 27311 3719 27325 3733
rect 30719 3719 30733 3733
rect 36311 3719 36325 3733
rect 36935 3719 36949 3733
rect 38663 3719 38677 3733
rect 22247 3695 22261 3709
rect 35303 3695 35317 3709
rect 35327 3695 35341 3709
rect 38759 3695 38773 3709
rect 38903 3695 38917 3709
rect 38951 3695 38965 3709
rect 39695 3695 39709 3709
rect 39767 3695 39781 3709
rect 39791 3695 39805 3709
rect 39863 3695 39877 3709
rect 39887 3695 39901 3709
rect 39959 3695 39973 3709
rect 40487 3695 40501 3709
rect 40559 3695 40573 3709
rect 40583 3695 40597 3709
rect 40655 3695 40669 3709
rect 15095 3671 15109 3685
rect 15143 3671 15157 3685
rect 15407 3671 15421 3685
rect 15479 3671 15493 3685
rect 21647 3671 21661 3685
rect 21695 3671 21709 3685
rect 21743 3671 21757 3685
rect 21815 3671 21829 3685
rect 21863 3671 21877 3685
rect 21935 3671 21949 3685
rect 21959 3671 21973 3685
rect 22055 3671 22069 3685
rect 22079 3671 22093 3685
rect 22151 3671 22165 3685
rect 22223 3671 22237 3685
rect 30383 3671 30397 3685
rect 30407 3671 30421 3685
rect 32375 3671 32389 3685
rect 32399 3671 32413 3685
rect 38855 3671 38869 3685
rect 38879 3671 38893 3685
rect 39047 3671 39061 3685
rect 39215 3671 39229 3685
rect 39263 3671 39277 3685
rect 39287 3671 39301 3685
rect 39359 3671 39373 3685
rect 39503 3671 39517 3685
rect 39551 3671 39565 3685
rect 39599 3671 39613 3685
rect 39647 3671 39661 3685
rect 39671 3671 39685 3685
rect 40055 3671 40069 3685
rect 40391 3671 40405 3685
rect 40439 3671 40453 3685
rect 40463 3671 40477 3685
rect 40775 3671 40789 3685
rect 40799 3671 40813 3685
rect 40871 3671 40885 3685
rect 41039 3671 41053 3685
rect 41087 3671 41101 3685
rect 15071 3647 15085 3661
rect 15335 3647 15349 3661
rect 15383 3647 15397 3661
rect 15671 3647 15685 3661
rect 21623 3647 21637 3661
rect 31703 3647 31717 3661
rect 31727 3647 31741 3661
rect 37199 3647 37213 3661
rect 37223 3647 37237 3661
rect 39167 3647 39181 3661
rect 39191 3647 39205 3661
rect 39455 3647 39469 3661
rect 39479 3647 39493 3661
rect 40151 3647 40165 3661
rect 40175 3647 40189 3661
rect 40247 3647 40261 3661
rect 40271 3647 40285 3661
rect 40343 3647 40357 3661
rect 40367 3647 40381 3661
rect 40991 3647 41005 3661
rect 41015 3647 41029 3661
rect 41183 3647 41197 3661
rect 41231 3647 41245 3661
rect 41303 3647 41317 3661
rect 41327 3647 41341 3661
rect 41399 3647 41413 3661
rect 47 3623 61 3637
rect 71 3623 85 3637
rect 95 3623 109 3637
rect 119 3623 133 3637
rect 143 3623 157 3637
rect 167 3623 181 3637
rect 191 3623 205 3637
rect 215 3623 229 3637
rect 239 3623 253 3637
rect 263 3623 277 3637
rect 287 3623 301 3637
rect 311 3623 325 3637
rect 335 3623 349 3637
rect 359 3623 373 3637
rect 383 3623 397 3637
rect 407 3623 421 3637
rect 431 3623 445 3637
rect 455 3623 469 3637
rect 479 3623 493 3637
rect 503 3623 517 3637
rect 527 3623 541 3637
rect 551 3623 565 3637
rect 575 3623 589 3637
rect 599 3623 613 3637
rect 623 3623 637 3637
rect 647 3623 661 3637
rect 671 3623 685 3637
rect 695 3623 709 3637
rect 719 3623 733 3637
rect 743 3623 757 3637
rect 767 3623 781 3637
rect 791 3623 805 3637
rect 815 3623 829 3637
rect 839 3623 853 3637
rect 863 3623 877 3637
rect 887 3623 901 3637
rect 911 3623 925 3637
rect 935 3623 949 3637
rect 959 3623 973 3637
rect 983 3623 997 3637
rect 1007 3623 1021 3637
rect 1031 3623 1045 3637
rect 1055 3623 1069 3637
rect 1079 3623 1093 3637
rect 1103 3623 1117 3637
rect 1127 3623 1141 3637
rect 1151 3623 1165 3637
rect 1175 3623 1189 3637
rect 1199 3623 1213 3637
rect 1223 3623 1237 3637
rect 14687 3623 14701 3637
rect 14735 3623 14749 3637
rect 14759 3623 14773 3637
rect 14831 3623 14845 3637
rect 14879 3623 14893 3637
rect 14927 3623 14941 3637
rect 14975 3623 14989 3637
rect 15023 3623 15037 3637
rect 15047 3623 15061 3637
rect 15887 3623 15901 3637
rect 21119 3623 21133 3637
rect 21167 3623 21181 3637
rect 21599 3623 21613 3637
rect 32543 3623 32557 3637
rect 37439 3623 37453 3637
rect 37463 3623 37477 3637
rect 41495 3623 41509 3637
rect 41855 3623 41869 3637
rect 41903 3623 41917 3637
rect 47 3575 61 3589
rect 71 3575 85 3589
rect 95 3575 109 3589
rect 119 3575 133 3589
rect 143 3575 157 3589
rect 167 3575 181 3589
rect 191 3575 205 3589
rect 215 3575 229 3589
rect 239 3575 253 3589
rect 263 3575 277 3589
rect 287 3575 301 3589
rect 311 3575 325 3589
rect 335 3575 349 3589
rect 359 3575 373 3589
rect 383 3575 397 3589
rect 407 3575 421 3589
rect 431 3575 445 3589
rect 455 3575 469 3589
rect 479 3575 493 3589
rect 503 3575 517 3589
rect 527 3575 541 3589
rect 551 3575 565 3589
rect 575 3575 589 3589
rect 599 3575 613 3589
rect 623 3575 637 3589
rect 647 3575 661 3589
rect 671 3575 685 3589
rect 695 3575 709 3589
rect 719 3575 733 3589
rect 743 3575 757 3589
rect 767 3575 781 3589
rect 791 3575 805 3589
rect 815 3575 829 3589
rect 839 3575 853 3589
rect 863 3575 877 3589
rect 887 3575 901 3589
rect 911 3575 925 3589
rect 935 3575 949 3589
rect 959 3575 973 3589
rect 983 3575 997 3589
rect 1007 3575 1021 3589
rect 1031 3575 1045 3589
rect 1055 3575 1069 3589
rect 1079 3575 1093 3589
rect 1103 3575 1117 3589
rect 1127 3575 1141 3589
rect 1151 3575 1165 3589
rect 1175 3575 1189 3589
rect 1199 3575 1213 3589
rect 1223 3575 1237 3589
rect 14591 3599 14605 3613
rect 14639 3599 14653 3613
rect 14663 3599 14677 3613
rect 16103 3599 16117 3613
rect 20231 3599 20245 3613
rect 20447 3599 20461 3613
rect 20495 3599 20509 3613
rect 20567 3599 20581 3613
rect 20591 3599 20605 3613
rect 20663 3599 20677 3613
rect 20735 3599 20749 3613
rect 20783 3599 20797 3613
rect 20831 3599 20845 3613
rect 20879 3599 20893 3613
rect 21023 3599 21037 3613
rect 21071 3599 21085 3613
rect 21095 3599 21109 3613
rect 21215 3599 21229 3613
rect 21263 3599 21277 3613
rect 21311 3599 21325 3613
rect 21359 3599 21373 3613
rect 21503 3599 21517 3613
rect 21551 3599 21565 3613
rect 21575 3599 21589 3613
rect 30215 3599 30229 3613
rect 32567 3599 32581 3613
rect 41615 3599 41629 3613
rect 41663 3599 41677 3613
rect 41711 3599 41725 3613
rect 41735 3599 41749 3613
rect 41807 3599 41821 3613
rect 41831 3599 41845 3613
rect 41999 3599 42013 3613
rect 42023 3599 42037 3613
rect 42119 3599 42133 3613
rect 14279 3575 14293 3589
rect 14351 3575 14365 3589
rect 14399 3575 14413 3589
rect 14447 3575 14461 3589
rect 14471 3575 14485 3589
rect 14543 3575 14557 3589
rect 14567 3575 14581 3589
rect 16319 3575 16333 3589
rect 19415 3575 19429 3589
rect 19487 3575 19501 3589
rect 19511 3575 19525 3589
rect 19583 3575 19597 3589
rect 19655 3575 19669 3589
rect 19727 3575 19741 3589
rect 19823 3575 19837 3589
rect 20975 3575 20989 3589
rect 20999 3575 21013 3589
rect 21455 3575 21469 3589
rect 21479 3575 21493 3589
rect 29015 3575 29029 3589
rect 29039 3575 29053 3589
rect 30767 3575 30781 3589
rect 30791 3575 30805 3589
rect 34967 3575 34981 3589
rect 34991 3575 35005 3589
rect 40127 3575 40141 3589
rect 40151 3575 40165 3589
rect 42215 3575 42229 3589
rect 13607 3551 13621 3565
rect 13679 3551 13693 3565
rect 13703 3551 13717 3565
rect 13775 3551 13789 3565
rect 13895 3551 13909 3565
rect 13991 3551 14005 3565
rect 14039 3551 14053 3565
rect 14207 3551 14221 3565
rect 14255 3551 14269 3565
rect 14375 3551 14389 3565
rect 14783 3551 14797 3565
rect 14855 3551 14869 3565
rect 16535 3551 16549 3565
rect 19295 3551 19309 3565
rect 19367 3551 19381 3565
rect 19391 3551 19405 3565
rect 30071 3551 30085 3565
rect 30095 3551 30109 3565
rect 36407 3551 36421 3565
rect 42335 3551 42349 3565
rect 13511 3527 13525 3541
rect 13559 3527 13573 3541
rect 13583 3527 13597 3541
rect 16751 3527 16765 3541
rect 19199 3527 19213 3541
rect 19247 3527 19261 3541
rect 19271 3527 19285 3541
rect 26951 3527 26965 3541
rect 26975 3527 26989 3541
rect 42455 3527 42469 3541
rect 12839 3503 12853 3517
rect 12887 3503 12901 3517
rect 13055 3503 13069 3517
rect 13127 3503 13141 3517
rect 13151 3503 13165 3517
rect 13223 3503 13237 3517
rect 13487 3503 13501 3517
rect 16967 3503 16981 3517
rect 18983 3503 18997 3517
rect 19055 3503 19069 3517
rect 19103 3503 19117 3517
rect 19151 3503 19165 3517
rect 19175 3503 19189 3517
rect 26591 3503 26605 3517
rect 26615 3503 26629 3517
rect 37943 3503 37957 3517
rect 37967 3503 37981 3517
rect 42599 3503 42613 3517
rect 12743 3479 12757 3493
rect 12791 3479 12805 3493
rect 12815 3479 12829 3493
rect 12983 3479 12997 3493
rect 13031 3479 13045 3493
rect 13319 3479 13333 3493
rect 13391 3479 13405 3493
rect 13439 3479 13453 3493
rect 13463 3479 13477 3493
rect 14951 3479 14965 3493
rect 17183 3479 17197 3493
rect 18791 3479 18805 3493
rect 18839 3479 18853 3493
rect 18887 3479 18901 3493
rect 18935 3479 18949 3493
rect 18959 3479 18973 3493
rect 28031 3479 28045 3493
rect 28055 3479 28069 3493
rect 42047 3479 42061 3493
rect 42695 3479 42709 3493
rect 12647 3455 12661 3469
rect 12695 3455 12709 3469
rect 12719 3455 12733 3469
rect 17399 3455 17413 3469
rect 18671 3455 18685 3469
rect 18743 3455 18757 3469
rect 18767 3455 18781 3469
rect 25175 3455 25189 3469
rect 26303 3455 26317 3469
rect 27455 3455 27469 3469
rect 30839 3455 30853 3469
rect 32063 3455 32077 3469
rect 33311 3455 33325 3469
rect 33743 3455 33757 3469
rect 33839 3455 33853 3469
rect 34247 3455 34261 3469
rect 38639 3455 38653 3469
rect 38663 3455 38677 3469
rect 41567 3455 41581 3469
rect 42815 3455 42829 3469
rect 12623 3431 12637 3445
rect 17471 3431 17485 3445
rect 18575 3431 18589 3445
rect 18623 3431 18637 3445
rect 18647 3431 18661 3445
rect 24599 3431 24613 3445
rect 24623 3431 24637 3445
rect 41687 3431 41701 3445
rect 41711 3431 41725 3445
rect 42935 3431 42949 3445
rect 12383 3407 12397 3421
rect 12455 3407 12469 3421
rect 12599 3407 12613 3421
rect 17615 3407 17629 3421
rect 18479 3407 18493 3421
rect 18527 3407 18541 3421
rect 18551 3407 18565 3421
rect 29855 3407 29869 3421
rect 37799 3407 37813 3421
rect 37823 3407 37837 3421
rect 41927 3407 41941 3421
rect 43055 3407 43069 3421
rect 43415 3407 43429 3421
rect 43463 3407 43477 3421
rect 47 3383 61 3397
rect 71 3383 85 3397
rect 95 3383 109 3397
rect 119 3383 133 3397
rect 143 3383 157 3397
rect 167 3383 181 3397
rect 191 3383 205 3397
rect 215 3383 229 3397
rect 239 3383 253 3397
rect 263 3383 277 3397
rect 287 3383 301 3397
rect 311 3383 325 3397
rect 335 3383 349 3397
rect 359 3383 373 3397
rect 383 3383 397 3397
rect 407 3383 421 3397
rect 431 3383 445 3397
rect 455 3383 469 3397
rect 479 3383 493 3397
rect 503 3383 517 3397
rect 527 3383 541 3397
rect 551 3383 565 3397
rect 575 3383 589 3397
rect 599 3383 613 3397
rect 623 3383 637 3397
rect 647 3383 661 3397
rect 671 3383 685 3397
rect 695 3383 709 3397
rect 719 3383 733 3397
rect 743 3383 757 3397
rect 767 3383 781 3397
rect 791 3383 805 3397
rect 815 3383 829 3397
rect 839 3383 853 3397
rect 863 3383 877 3397
rect 887 3383 901 3397
rect 911 3383 925 3397
rect 935 3383 949 3397
rect 959 3383 973 3397
rect 983 3383 997 3397
rect 1007 3383 1021 3397
rect 1031 3383 1045 3397
rect 1055 3383 1069 3397
rect 1079 3383 1093 3397
rect 1103 3383 1117 3397
rect 1127 3383 1141 3397
rect 1151 3383 1165 3397
rect 1175 3383 1189 3397
rect 1199 3383 1213 3397
rect 1223 3383 1237 3397
rect 1247 3383 1261 3397
rect 12287 3383 12301 3397
rect 12335 3383 12349 3397
rect 12359 3383 12373 3397
rect 12551 3383 12565 3397
rect 12575 3383 12589 3397
rect 17831 3383 17845 3397
rect 18455 3383 18469 3397
rect 26831 3383 26845 3397
rect 26855 3383 26869 3397
rect 28199 3383 28213 3397
rect 43151 3383 43165 3397
rect 43199 3383 43213 3397
rect 43271 3383 43285 3397
rect 43319 3383 43333 3397
rect 43367 3383 43381 3397
rect 43391 3383 43405 3397
rect 43559 3383 43573 3397
rect 43607 3383 43621 3397
rect 43655 3383 43669 3397
rect 47 3335 61 3349
rect 71 3335 85 3349
rect 95 3335 109 3349
rect 119 3335 133 3349
rect 143 3335 157 3349
rect 167 3335 181 3349
rect 191 3335 205 3349
rect 215 3335 229 3349
rect 239 3335 253 3349
rect 263 3335 277 3349
rect 287 3335 301 3349
rect 311 3335 325 3349
rect 335 3335 349 3349
rect 359 3335 373 3349
rect 383 3335 397 3349
rect 407 3335 421 3349
rect 431 3335 445 3349
rect 455 3335 469 3349
rect 479 3335 493 3349
rect 503 3335 517 3349
rect 527 3335 541 3349
rect 551 3335 565 3349
rect 575 3335 589 3349
rect 599 3335 613 3349
rect 623 3335 637 3349
rect 647 3335 661 3349
rect 671 3335 685 3349
rect 695 3335 709 3349
rect 719 3335 733 3349
rect 743 3335 757 3349
rect 767 3335 781 3349
rect 791 3335 805 3349
rect 815 3335 829 3349
rect 839 3335 853 3349
rect 863 3335 877 3349
rect 887 3335 901 3349
rect 911 3335 925 3349
rect 935 3335 949 3349
rect 959 3335 973 3349
rect 983 3335 997 3349
rect 1007 3335 1021 3349
rect 1031 3335 1045 3349
rect 1055 3335 1069 3349
rect 1079 3335 1093 3349
rect 1103 3335 1117 3349
rect 1127 3335 1141 3349
rect 1151 3335 1165 3349
rect 1175 3335 1189 3349
rect 1199 3335 1213 3349
rect 1223 3335 1237 3349
rect 1247 3335 1261 3349
rect 12191 3359 12205 3373
rect 12239 3359 12253 3373
rect 12263 3359 12277 3373
rect 17903 3359 17917 3373
rect 18359 3359 18373 3373
rect 18407 3359 18421 3373
rect 18431 3359 18445 3373
rect 28823 3359 28837 3373
rect 28847 3359 28861 3373
rect 30119 3359 30133 3373
rect 33671 3359 33685 3373
rect 33695 3359 33709 3373
rect 43751 3359 43765 3373
rect 12167 3335 12181 3349
rect 18047 3335 18061 3349
rect 18335 3335 18349 3349
rect 24815 3335 24829 3349
rect 24839 3335 24853 3349
rect 37007 3335 37021 3349
rect 37031 3335 37045 3349
rect 40007 3335 40021 3349
rect 40079 3335 40093 3349
rect 43079 3335 43093 3349
rect 43871 3335 43885 3349
rect 44015 3335 44029 3349
rect 44063 3335 44077 3349
rect 12143 3311 12157 3325
rect 18263 3311 18277 3325
rect 18311 3311 18325 3325
rect 35831 3311 35845 3325
rect 35855 3311 35869 3325
rect 43943 3311 43957 3325
rect 43991 3311 44005 3325
rect 44183 3311 44197 3325
rect 12023 3287 12037 3301
rect 12095 3287 12109 3301
rect 12119 3287 12133 3301
rect 28535 3287 28549 3301
rect 28559 3287 28573 3301
rect 41783 3287 41797 3301
rect 41807 3287 41821 3301
rect 44351 3287 44365 3301
rect 44399 3287 44413 3301
rect 44471 3287 44485 3301
rect 11999 3263 12013 3277
rect 22535 3263 22549 3277
rect 22559 3263 22573 3277
rect 26063 3263 26077 3277
rect 37079 3263 37093 3277
rect 37175 3263 37189 3277
rect 39407 3263 39421 3277
rect 40199 3263 40213 3277
rect 44567 3263 44581 3277
rect 11879 3239 11893 3253
rect 11951 3239 11965 3253
rect 11975 3239 11989 3253
rect 18815 3239 18829 3253
rect 18839 3239 18853 3253
rect 20927 3239 20941 3253
rect 25439 3239 25453 3253
rect 25463 3239 25477 3253
rect 31583 3239 31597 3253
rect 31607 3239 31621 3253
rect 37631 3239 37645 3253
rect 43127 3239 43141 3253
rect 43151 3239 43165 3253
rect 44711 3239 44725 3253
rect 11711 3215 11725 3229
rect 11807 3215 11821 3229
rect 11831 3215 11845 3229
rect 32639 3215 32653 3229
rect 44807 3215 44821 3229
rect 11615 3191 11629 3205
rect 11663 3191 11677 3205
rect 11687 3191 11701 3205
rect 25223 3191 25237 3205
rect 25247 3191 25261 3205
rect 25511 3191 25525 3205
rect 26231 3191 26245 3205
rect 31367 3191 31381 3205
rect 31391 3191 31405 3205
rect 33263 3191 33277 3205
rect 33287 3191 33301 3205
rect 44903 3191 44917 3205
rect 11591 3167 11605 3181
rect 20639 3167 20653 3181
rect 20663 3167 20677 3181
rect 22895 3167 22909 3181
rect 22919 3167 22933 3181
rect 31799 3167 31813 3181
rect 31823 3167 31837 3181
rect 36959 3167 36973 3181
rect 39911 3167 39925 3181
rect 44999 3167 45013 3181
rect 47 3143 61 3157
rect 71 3143 85 3157
rect 95 3143 109 3157
rect 119 3143 133 3157
rect 143 3143 157 3157
rect 167 3143 181 3157
rect 191 3143 205 3157
rect 215 3143 229 3157
rect 239 3143 253 3157
rect 263 3143 277 3157
rect 287 3143 301 3157
rect 311 3143 325 3157
rect 335 3143 349 3157
rect 359 3143 373 3157
rect 383 3143 397 3157
rect 407 3143 421 3157
rect 431 3143 445 3157
rect 455 3143 469 3157
rect 479 3143 493 3157
rect 503 3143 517 3157
rect 527 3143 541 3157
rect 551 3143 565 3157
rect 575 3143 589 3157
rect 599 3143 613 3157
rect 623 3143 637 3157
rect 647 3143 661 3157
rect 671 3143 685 3157
rect 695 3143 709 3157
rect 719 3143 733 3157
rect 743 3143 757 3157
rect 767 3143 781 3157
rect 791 3143 805 3157
rect 815 3143 829 3157
rect 839 3143 853 3157
rect 863 3143 877 3157
rect 887 3143 901 3157
rect 911 3143 925 3157
rect 935 3143 949 3157
rect 959 3143 973 3157
rect 983 3143 997 3157
rect 1007 3143 1021 3157
rect 1031 3143 1045 3157
rect 1055 3143 1069 3157
rect 1079 3143 1093 3157
rect 1103 3143 1117 3157
rect 1127 3143 1141 3157
rect 1151 3143 1165 3157
rect 1175 3143 1189 3157
rect 1199 3143 1213 3157
rect 1223 3143 1237 3157
rect 1247 3143 1261 3157
rect 1271 3143 1285 3157
rect 11471 3143 11485 3157
rect 11519 3143 11533 3157
rect 11567 3143 11581 3157
rect 38711 3143 38725 3157
rect 41351 3143 41365 3157
rect 45119 3143 45133 3157
rect 47 3095 61 3109
rect 71 3095 85 3109
rect 95 3095 109 3109
rect 119 3095 133 3109
rect 143 3095 157 3109
rect 167 3095 181 3109
rect 191 3095 205 3109
rect 215 3095 229 3109
rect 239 3095 253 3109
rect 263 3095 277 3109
rect 287 3095 301 3109
rect 311 3095 325 3109
rect 335 3095 349 3109
rect 359 3095 373 3109
rect 383 3095 397 3109
rect 407 3095 421 3109
rect 431 3095 445 3109
rect 455 3095 469 3109
rect 479 3095 493 3109
rect 503 3095 517 3109
rect 527 3095 541 3109
rect 551 3095 565 3109
rect 575 3095 589 3109
rect 599 3095 613 3109
rect 623 3095 637 3109
rect 647 3095 661 3109
rect 671 3095 685 3109
rect 695 3095 709 3109
rect 719 3095 733 3109
rect 743 3095 757 3109
rect 767 3095 781 3109
rect 791 3095 805 3109
rect 815 3095 829 3109
rect 839 3095 853 3109
rect 863 3095 877 3109
rect 887 3095 901 3109
rect 911 3095 925 3109
rect 935 3095 949 3109
rect 959 3095 973 3109
rect 983 3095 997 3109
rect 1007 3095 1021 3109
rect 1031 3095 1045 3109
rect 1055 3095 1069 3109
rect 1079 3095 1093 3109
rect 1103 3095 1117 3109
rect 1127 3095 1141 3109
rect 1151 3095 1165 3109
rect 1175 3095 1189 3109
rect 1199 3095 1213 3109
rect 1223 3095 1237 3109
rect 1247 3095 1261 3109
rect 1271 3095 1285 3109
rect 11375 3119 11389 3133
rect 11423 3119 11437 3133
rect 11447 3119 11461 3133
rect 13247 3119 13261 3133
rect 14903 3119 14917 3133
rect 14927 3119 14941 3133
rect 21767 3119 21781 3133
rect 23951 3119 23965 3133
rect 24791 3119 24805 3133
rect 31295 3119 31309 3133
rect 38015 3119 38029 3133
rect 45215 3119 45229 3133
rect 11351 3095 11365 3109
rect 19079 3095 19093 3109
rect 23615 3095 23629 3109
rect 23639 3095 23653 3109
rect 26207 3095 26221 3109
rect 27791 3095 27805 3109
rect 28175 3095 28189 3109
rect 28295 3095 28309 3109
rect 28391 3095 28405 3109
rect 33911 3095 33925 3109
rect 33935 3095 33949 3109
rect 37847 3095 37861 3109
rect 37871 3095 37885 3109
rect 45335 3095 45349 3109
rect 11327 3071 11341 3085
rect 20759 3071 20773 3085
rect 20783 3071 20797 3085
rect 45455 3071 45469 3085
rect 11231 3047 11245 3061
rect 11279 3047 11293 3061
rect 11303 3047 11317 3061
rect 24215 3047 24229 3061
rect 24239 3047 24253 3061
rect 26783 3047 26797 3061
rect 27983 3047 27997 3061
rect 28079 3047 28093 3061
rect 34319 3047 34333 3061
rect 34343 3047 34357 3061
rect 37103 3047 37117 3061
rect 37127 3047 37141 3061
rect 43343 3047 43357 3061
rect 43367 3047 43381 3061
rect 45551 3047 45565 3061
rect 11135 3023 11149 3037
rect 11183 3023 11197 3037
rect 11207 3023 11221 3037
rect 18599 3023 18613 3037
rect 18623 3023 18637 3037
rect 22391 3023 22405 3037
rect 22415 3023 22429 3037
rect 45647 3023 45661 3037
rect 11087 2999 11101 3013
rect 19031 2999 19045 3013
rect 19055 2999 19069 3013
rect 26351 2999 26365 3013
rect 26375 2999 26389 3013
rect 30287 2999 30301 3013
rect 30311 2999 30325 3013
rect 45767 2999 45781 3013
rect 45815 2999 45829 3013
rect 45863 2999 45877 3013
rect 45887 2999 45901 3013
rect 45959 2999 45973 3013
rect 10967 2975 10981 2989
rect 11039 2975 11053 2989
rect 11063 2975 11077 2989
rect 23855 2975 23869 2989
rect 23879 2975 23893 2989
rect 28487 2975 28501 2989
rect 28583 2975 28597 2989
rect 28679 2975 28693 2989
rect 28967 2975 28981 2989
rect 29279 2975 29293 2989
rect 33383 2975 33397 2989
rect 33407 2975 33421 2989
rect 46055 2975 46069 2989
rect 46079 2975 46093 2989
rect 46151 2975 46165 2989
rect 10871 2951 10885 2965
rect 10919 2951 10933 2965
rect 10943 2951 10957 2965
rect 20399 2951 20413 2965
rect 38279 2951 38293 2965
rect 38303 2951 38317 2965
rect 46247 2951 46261 2965
rect 8615 2927 8629 2941
rect 8663 2927 8677 2941
rect 8687 2927 8701 2941
rect 8735 2927 8749 2941
rect 10847 2927 10861 2941
rect 18719 2927 18733 2941
rect 18743 2927 18757 2941
rect 31895 2927 31909 2941
rect 31919 2927 31933 2941
rect 46367 2927 46381 2941
rect 47 2903 61 2917
rect 71 2903 85 2917
rect 95 2903 109 2917
rect 119 2903 133 2917
rect 143 2903 157 2917
rect 167 2903 181 2917
rect 191 2903 205 2917
rect 215 2903 229 2917
rect 239 2903 253 2917
rect 263 2903 277 2917
rect 287 2903 301 2917
rect 311 2903 325 2917
rect 335 2903 349 2917
rect 359 2903 373 2917
rect 383 2903 397 2917
rect 407 2903 421 2917
rect 431 2903 445 2917
rect 455 2903 469 2917
rect 479 2903 493 2917
rect 503 2903 517 2917
rect 527 2903 541 2917
rect 551 2903 565 2917
rect 575 2903 589 2917
rect 599 2903 613 2917
rect 623 2903 637 2917
rect 647 2903 661 2917
rect 671 2903 685 2917
rect 695 2903 709 2917
rect 719 2903 733 2917
rect 743 2903 757 2917
rect 767 2903 781 2917
rect 791 2903 805 2917
rect 815 2903 829 2917
rect 839 2903 853 2917
rect 863 2903 877 2917
rect 887 2903 901 2917
rect 911 2903 925 2917
rect 935 2903 949 2917
rect 959 2903 973 2917
rect 983 2903 997 2917
rect 1007 2903 1021 2917
rect 1031 2903 1045 2917
rect 1055 2903 1069 2917
rect 1079 2903 1093 2917
rect 1103 2903 1117 2917
rect 1127 2903 1141 2917
rect 1151 2903 1165 2917
rect 1175 2903 1189 2917
rect 1199 2903 1213 2917
rect 1223 2903 1237 2917
rect 1247 2903 1261 2917
rect 1271 2903 1285 2917
rect 1295 2903 1309 2917
rect 8591 2903 8605 2917
rect 8759 2903 8773 2917
rect 8783 2903 8797 2917
rect 8855 2903 8869 2917
rect 10823 2903 10837 2917
rect 46463 2903 46477 2917
rect 46487 2903 46501 2917
rect 46559 2903 46573 2917
rect 46871 2903 46885 2917
rect 46943 2903 46957 2917
rect 47 2855 61 2869
rect 71 2855 85 2869
rect 95 2855 109 2869
rect 119 2855 133 2869
rect 143 2855 157 2869
rect 167 2855 181 2869
rect 191 2855 205 2869
rect 215 2855 229 2869
rect 239 2855 253 2869
rect 263 2855 277 2869
rect 287 2855 301 2869
rect 311 2855 325 2869
rect 335 2855 349 2869
rect 359 2855 373 2869
rect 383 2855 397 2869
rect 407 2855 421 2869
rect 431 2855 445 2869
rect 455 2855 469 2869
rect 479 2855 493 2869
rect 503 2855 517 2869
rect 527 2855 541 2869
rect 551 2855 565 2869
rect 575 2855 589 2869
rect 599 2855 613 2869
rect 623 2855 637 2869
rect 647 2855 661 2869
rect 671 2855 685 2869
rect 695 2855 709 2869
rect 719 2855 733 2869
rect 743 2855 757 2869
rect 767 2855 781 2869
rect 791 2855 805 2869
rect 815 2855 829 2869
rect 839 2855 853 2869
rect 863 2855 877 2869
rect 887 2855 901 2869
rect 911 2855 925 2869
rect 935 2855 949 2869
rect 959 2855 973 2869
rect 983 2855 997 2869
rect 1007 2855 1021 2869
rect 1031 2855 1045 2869
rect 1055 2855 1069 2869
rect 1079 2855 1093 2869
rect 1103 2855 1117 2869
rect 1127 2855 1141 2869
rect 1151 2855 1165 2869
rect 1175 2855 1189 2869
rect 1199 2855 1213 2869
rect 1223 2855 1237 2869
rect 1247 2855 1261 2869
rect 1271 2855 1285 2869
rect 1295 2855 1309 2869
rect 8351 2879 8365 2893
rect 8423 2879 8437 2893
rect 8567 2879 8581 2893
rect 8951 2879 8965 2893
rect 10727 2879 10741 2893
rect 10775 2879 10789 2893
rect 10799 2879 10813 2893
rect 46679 2879 46693 2893
rect 46703 2879 46717 2893
rect 46823 2879 46837 2893
rect 46847 2879 46861 2893
rect 47063 2879 47077 2893
rect 47087 2879 47101 2893
rect 47159 2879 47173 2893
rect 8255 2855 8269 2869
rect 8303 2855 8317 2869
rect 8327 2855 8341 2869
rect 8519 2855 8533 2869
rect 8543 2855 8557 2869
rect 9023 2855 9037 2869
rect 10703 2855 10717 2869
rect 19343 2855 19357 2869
rect 19367 2855 19381 2869
rect 47255 2855 47269 2869
rect 47543 2855 47557 2869
rect 47591 2855 47605 2869
rect 8159 2831 8173 2845
rect 8207 2831 8221 2845
rect 8231 2831 8245 2845
rect 9047 2831 9061 2845
rect 10343 2831 10357 2845
rect 10415 2831 10429 2845
rect 10679 2831 10693 2845
rect 46799 2831 46813 2845
rect 46823 2831 46837 2845
rect 47375 2831 47389 2845
rect 47519 2831 47533 2845
rect 47711 2831 47725 2845
rect 47735 2831 47749 2845
rect 47831 2831 47845 2845
rect 47951 2831 47965 2845
rect 47999 2831 48013 2845
rect 8039 2807 8053 2821
rect 8087 2807 8101 2821
rect 8111 2807 8125 2821
rect 9143 2807 9157 2821
rect 10127 2807 10141 2821
rect 10175 2807 10189 2821
rect 10199 2807 10213 2821
rect 10271 2807 10285 2821
rect 10319 2807 10333 2821
rect 10511 2807 10525 2821
rect 10535 2807 10549 2821
rect 10607 2807 10621 2821
rect 10655 2807 10669 2821
rect 45743 2807 45757 2821
rect 45767 2807 45781 2821
rect 47471 2807 47485 2821
rect 47495 2807 47509 2821
rect 48119 2807 48133 2821
rect 8015 2783 8029 2797
rect 8135 2783 8149 2797
rect 9215 2783 9229 2797
rect 10031 2783 10045 2797
rect 10079 2783 10093 2797
rect 10103 2783 10117 2797
rect 12767 2783 12781 2797
rect 12791 2783 12805 2797
rect 13175 2783 13189 2797
rect 21047 2783 21061 2797
rect 21071 2783 21085 2797
rect 38495 2783 38509 2797
rect 38519 2783 38533 2797
rect 44927 2783 44941 2797
rect 47207 2783 47221 2797
rect 47879 2783 47893 2797
rect 48263 2783 48277 2797
rect 7919 2759 7933 2773
rect 7967 2759 7981 2773
rect 7991 2759 8005 2773
rect 9239 2759 9253 2773
rect 9983 2759 9997 2773
rect 36767 2759 36781 2773
rect 36791 2759 36805 2773
rect 38399 2759 38413 2773
rect 38423 2759 38437 2773
rect 45935 2759 45949 2773
rect 45959 2759 45973 2773
rect 48383 2759 48397 2773
rect 48407 2759 48421 2773
rect 48479 2759 48493 2773
rect 7895 2735 7909 2749
rect 9335 2735 9349 2749
rect 9887 2735 9901 2749
rect 9935 2735 9949 2749
rect 9959 2735 9973 2749
rect 14615 2735 14629 2749
rect 14639 2735 14653 2749
rect 21671 2735 21685 2749
rect 21695 2735 21709 2749
rect 48575 2735 48589 2749
rect 7607 2711 7621 2725
rect 7823 2711 7837 2725
rect 7847 2711 7861 2725
rect 9431 2711 9445 2725
rect 9767 2711 9781 2725
rect 9815 2711 9829 2725
rect 9839 2711 9853 2725
rect 33527 2711 33541 2725
rect 34175 2711 34189 2725
rect 34487 2711 34501 2725
rect 34559 2711 34573 2725
rect 36239 2711 36253 2725
rect 36263 2711 36277 2725
rect 36839 2711 36853 2725
rect 40823 2711 40837 2725
rect 48671 2711 48685 2725
rect 48719 2711 48733 2725
rect 48767 2711 48781 2725
rect 7199 2687 7213 2701
rect 9551 2687 9565 2701
rect 9743 2687 9757 2701
rect 12911 2687 12925 2701
rect 14423 2687 14437 2701
rect 14447 2687 14461 2701
rect 37247 2687 37261 2701
rect 43631 2687 43645 2701
rect 43655 2687 43669 2701
rect 48863 2687 48877 2701
rect 47 2663 61 2677
rect 71 2663 85 2677
rect 95 2663 109 2677
rect 119 2663 133 2677
rect 143 2663 157 2677
rect 167 2663 181 2677
rect 191 2663 205 2677
rect 215 2663 229 2677
rect 239 2663 253 2677
rect 263 2663 277 2677
rect 287 2663 301 2677
rect 311 2663 325 2677
rect 335 2663 349 2677
rect 359 2663 373 2677
rect 383 2663 397 2677
rect 407 2663 421 2677
rect 431 2663 445 2677
rect 455 2663 469 2677
rect 479 2663 493 2677
rect 503 2663 517 2677
rect 527 2663 541 2677
rect 551 2663 565 2677
rect 575 2663 589 2677
rect 599 2663 613 2677
rect 623 2663 637 2677
rect 647 2663 661 2677
rect 671 2663 685 2677
rect 695 2663 709 2677
rect 719 2663 733 2677
rect 743 2663 757 2677
rect 767 2663 781 2677
rect 791 2663 805 2677
rect 815 2663 829 2677
rect 839 2663 853 2677
rect 863 2663 877 2677
rect 887 2663 901 2677
rect 911 2663 925 2677
rect 935 2663 949 2677
rect 959 2663 973 2677
rect 983 2663 997 2677
rect 1007 2663 1021 2677
rect 1031 2663 1045 2677
rect 1055 2663 1069 2677
rect 1079 2663 1093 2677
rect 1103 2663 1117 2677
rect 1127 2663 1141 2677
rect 1151 2663 1165 2677
rect 1175 2663 1189 2677
rect 1199 2663 1213 2677
rect 1223 2663 1237 2677
rect 1247 2663 1261 2677
rect 1271 2663 1285 2677
rect 1295 2663 1309 2677
rect 1319 2663 1333 2677
rect 6983 2663 6997 2677
rect 9647 2663 9661 2677
rect 9695 2663 9709 2677
rect 19463 2663 19477 2677
rect 19487 2663 19501 2677
rect 26711 2663 26725 2677
rect 26735 2663 26749 2677
rect 32687 2663 32701 2677
rect 32711 2663 32725 2677
rect 37655 2663 37669 2677
rect 37679 2663 37693 2677
rect 39839 2663 39853 2677
rect 39863 2663 39877 2677
rect 44039 2663 44053 2677
rect 44063 2663 44077 2677
rect 48959 2663 48973 2677
rect 47 2615 61 2629
rect 71 2615 85 2629
rect 95 2615 109 2629
rect 119 2615 133 2629
rect 143 2615 157 2629
rect 167 2615 181 2629
rect 191 2615 205 2629
rect 215 2615 229 2629
rect 239 2615 253 2629
rect 263 2615 277 2629
rect 287 2615 301 2629
rect 311 2615 325 2629
rect 335 2615 349 2629
rect 359 2615 373 2629
rect 383 2615 397 2629
rect 407 2615 421 2629
rect 431 2615 445 2629
rect 455 2615 469 2629
rect 479 2615 493 2629
rect 503 2615 517 2629
rect 527 2615 541 2629
rect 551 2615 565 2629
rect 575 2615 589 2629
rect 599 2615 613 2629
rect 623 2615 637 2629
rect 647 2615 661 2629
rect 671 2615 685 2629
rect 695 2615 709 2629
rect 719 2615 733 2629
rect 743 2615 757 2629
rect 767 2615 781 2629
rect 791 2615 805 2629
rect 815 2615 829 2629
rect 839 2615 853 2629
rect 863 2615 877 2629
rect 887 2615 901 2629
rect 911 2615 925 2629
rect 935 2615 949 2629
rect 959 2615 973 2629
rect 983 2615 997 2629
rect 1007 2615 1021 2629
rect 1031 2615 1045 2629
rect 1055 2615 1069 2629
rect 1079 2615 1093 2629
rect 1103 2615 1117 2629
rect 1127 2615 1141 2629
rect 1151 2615 1165 2629
rect 1175 2615 1189 2629
rect 1199 2615 1213 2629
rect 1223 2615 1237 2629
rect 1247 2615 1261 2629
rect 1271 2615 1285 2629
rect 1295 2615 1309 2629
rect 1319 2615 1333 2629
rect 5759 2639 5773 2653
rect 5831 2639 5845 2653
rect 5855 2639 5869 2653
rect 5951 2639 5965 2653
rect 5975 2639 5989 2653
rect 6071 2639 6085 2653
rect 6119 2639 6133 2653
rect 6167 2639 6181 2653
rect 6311 2639 6325 2653
rect 6383 2639 6397 2653
rect 6935 2639 6949 2653
rect 44759 2639 44773 2653
rect 45023 2639 45037 2653
rect 49055 2639 49069 2653
rect 49079 2639 49093 2653
rect 49151 2639 49165 2653
rect 5735 2615 5749 2629
rect 6263 2615 6277 2629
rect 6287 2615 6301 2629
rect 6479 2615 6493 2629
rect 6575 2615 6589 2629
rect 10751 2615 10765 2629
rect 10775 2615 10789 2629
rect 11543 2615 11557 2629
rect 40511 2615 40525 2629
rect 49247 2615 49261 2629
rect 5639 2591 5653 2605
rect 5687 2591 5701 2605
rect 5711 2591 5725 2605
rect 13367 2591 13381 2605
rect 19703 2591 19717 2605
rect 19727 2591 19741 2605
rect 24455 2591 24469 2605
rect 24479 2591 24493 2605
rect 28895 2591 28909 2605
rect 29087 2591 29101 2605
rect 34103 2591 34117 2605
rect 34127 2591 34141 2605
rect 36071 2591 36085 2605
rect 38831 2591 38845 2605
rect 38855 2591 38869 2605
rect 49343 2591 49357 2605
rect 5543 2567 5557 2581
rect 5591 2567 5605 2581
rect 5615 2567 5629 2581
rect 9527 2567 9541 2581
rect 9551 2567 9565 2581
rect 11255 2567 11269 2581
rect 11279 2567 11293 2581
rect 39335 2567 39349 2581
rect 39359 2567 39373 2581
rect 45623 2567 45637 2581
rect 45647 2567 45661 2581
rect 49439 2567 49453 2581
rect 5519 2543 5533 2557
rect 12431 2543 12445 2557
rect 12455 2543 12469 2557
rect 28127 2543 28141 2557
rect 28151 2543 28165 2557
rect 28319 2543 28333 2557
rect 49535 2543 49549 2557
rect 5399 2519 5413 2533
rect 5447 2519 5461 2533
rect 5471 2519 5485 2533
rect 7871 2519 7885 2533
rect 22991 2519 23005 2533
rect 23015 2519 23029 2533
rect 37991 2519 38005 2533
rect 46991 2519 47005 2533
rect 47279 2519 47293 2533
rect 49631 2519 49645 2533
rect 5303 2495 5317 2509
rect 5351 2495 5365 2509
rect 5375 2495 5389 2509
rect 9623 2495 9637 2509
rect 9647 2495 9661 2509
rect 37703 2495 37717 2509
rect 41639 2495 41653 2509
rect 43295 2495 43309 2509
rect 49727 2495 49741 2509
rect 5279 2471 5293 2485
rect 9119 2471 9133 2485
rect 9143 2471 9157 2485
rect 14711 2471 14725 2485
rect 14735 2471 14749 2485
rect 48095 2471 48109 2485
rect 48119 2471 48133 2485
rect 49391 2471 49405 2485
rect 49847 2471 49861 2485
rect 50015 2471 50029 2485
rect 50063 2471 50077 2485
rect 5183 2447 5197 2461
rect 5231 2447 5245 2461
rect 5255 2447 5269 2461
rect 6455 2447 6469 2461
rect 6479 2447 6493 2461
rect 12311 2447 12325 2461
rect 12335 2447 12349 2461
rect 26015 2447 26029 2461
rect 35615 2447 35629 2461
rect 37607 2447 37621 2461
rect 38255 2447 38269 2461
rect 47111 2447 47125 2461
rect 49967 2447 49981 2461
rect 49991 2447 50005 2461
rect 50159 2447 50173 2461
rect 47 2423 61 2437
rect 71 2423 85 2437
rect 95 2423 109 2437
rect 119 2423 133 2437
rect 143 2423 157 2437
rect 167 2423 181 2437
rect 191 2423 205 2437
rect 215 2423 229 2437
rect 239 2423 253 2437
rect 263 2423 277 2437
rect 287 2423 301 2437
rect 311 2423 325 2437
rect 335 2423 349 2437
rect 359 2423 373 2437
rect 383 2423 397 2437
rect 407 2423 421 2437
rect 431 2423 445 2437
rect 455 2423 469 2437
rect 479 2423 493 2437
rect 503 2423 517 2437
rect 527 2423 541 2437
rect 551 2423 565 2437
rect 575 2423 589 2437
rect 599 2423 613 2437
rect 623 2423 637 2437
rect 647 2423 661 2437
rect 671 2423 685 2437
rect 695 2423 709 2437
rect 719 2423 733 2437
rect 743 2423 757 2437
rect 767 2423 781 2437
rect 791 2423 805 2437
rect 815 2423 829 2437
rect 839 2423 853 2437
rect 863 2423 877 2437
rect 887 2423 901 2437
rect 911 2423 925 2437
rect 935 2423 949 2437
rect 959 2423 973 2437
rect 983 2423 997 2437
rect 1007 2423 1021 2437
rect 1031 2423 1045 2437
rect 1055 2423 1069 2437
rect 1079 2423 1093 2437
rect 1103 2423 1117 2437
rect 1127 2423 1141 2437
rect 1151 2423 1165 2437
rect 1175 2423 1189 2437
rect 1199 2423 1213 2437
rect 1223 2423 1237 2437
rect 1247 2423 1261 2437
rect 1271 2423 1285 2437
rect 1295 2423 1309 2437
rect 1319 2423 1333 2437
rect 1343 2423 1357 2437
rect 5159 2423 5173 2437
rect 8831 2423 8845 2437
rect 8855 2423 8869 2437
rect 8879 2423 8893 2437
rect 9071 2423 9085 2437
rect 9263 2423 9277 2437
rect 13535 2423 13549 2437
rect 13559 2423 13573 2437
rect 25415 2423 25429 2437
rect 30743 2423 30757 2437
rect 34079 2423 34093 2437
rect 39095 2423 39109 2437
rect 40895 2423 40909 2437
rect 44975 2423 44989 2437
rect 44999 2423 45013 2437
rect 46751 2423 46765 2437
rect 48599 2423 48613 2437
rect 49559 2423 49573 2437
rect 49655 2423 49669 2437
rect 50255 2423 50269 2437
rect 47 2375 61 2389
rect 71 2375 85 2389
rect 95 2375 109 2389
rect 119 2375 133 2389
rect 143 2375 157 2389
rect 167 2375 181 2389
rect 191 2375 205 2389
rect 215 2375 229 2389
rect 239 2375 253 2389
rect 263 2375 277 2389
rect 287 2375 301 2389
rect 311 2375 325 2389
rect 335 2375 349 2389
rect 359 2375 373 2389
rect 383 2375 397 2389
rect 407 2375 421 2389
rect 431 2375 445 2389
rect 455 2375 469 2389
rect 479 2375 493 2389
rect 503 2375 517 2389
rect 527 2375 541 2389
rect 551 2375 565 2389
rect 575 2375 589 2389
rect 599 2375 613 2389
rect 623 2375 637 2389
rect 647 2375 661 2389
rect 671 2375 685 2389
rect 695 2375 709 2389
rect 719 2375 733 2389
rect 743 2375 757 2389
rect 767 2375 781 2389
rect 791 2375 805 2389
rect 815 2375 829 2389
rect 839 2375 853 2389
rect 863 2375 877 2389
rect 887 2375 901 2389
rect 911 2375 925 2389
rect 935 2375 949 2389
rect 959 2375 973 2389
rect 983 2375 997 2389
rect 1007 2375 1021 2389
rect 1031 2375 1045 2389
rect 1055 2375 1069 2389
rect 1079 2375 1093 2389
rect 1103 2375 1117 2389
rect 1127 2375 1141 2389
rect 1151 2375 1165 2389
rect 1175 2375 1189 2389
rect 1199 2375 1213 2389
rect 1223 2375 1237 2389
rect 1247 2375 1261 2389
rect 1271 2375 1285 2389
rect 1295 2375 1309 2389
rect 1319 2375 1333 2389
rect 1343 2375 1357 2389
rect 5063 2399 5077 2413
rect 5111 2399 5125 2413
rect 5135 2399 5149 2413
rect 7799 2399 7813 2413
rect 7823 2399 7837 2413
rect 35999 2399 36013 2413
rect 39311 2399 39325 2413
rect 43223 2399 43237 2413
rect 46199 2399 46213 2413
rect 47615 2399 47629 2413
rect 48191 2399 48205 2413
rect 48311 2399 48325 2413
rect 48527 2399 48541 2413
rect 50351 2399 50365 2413
rect 5039 2375 5053 2389
rect 8927 2375 8941 2389
rect 8951 2375 8965 2389
rect 13655 2375 13669 2389
rect 13679 2375 13693 2389
rect 46127 2375 46141 2389
rect 46151 2375 46165 2389
rect 46175 2375 46189 2389
rect 50831 2375 50845 2389
rect 4919 2351 4933 2365
rect 4991 2351 5005 2365
rect 5015 2351 5029 2365
rect 6143 2351 6157 2365
rect 6167 2351 6181 2365
rect 6215 2351 6229 2365
rect 6431 2351 6445 2365
rect 7775 2351 7789 2365
rect 32207 2351 32221 2365
rect 32231 2351 32245 2365
rect 34775 2351 34789 2365
rect 34799 2351 34813 2365
rect 43727 2351 43741 2365
rect 43751 2351 43765 2365
rect 50879 2351 50893 2365
rect 51023 2351 51037 2365
rect 51071 2351 51085 2365
rect 4895 2327 4909 2341
rect 27071 2327 27085 2341
rect 27095 2327 27109 2341
rect 29207 2327 29221 2341
rect 32999 2327 33013 2341
rect 51167 2327 51181 2341
rect 51215 2327 51229 2341
rect 51263 2327 51277 2341
rect 4775 2303 4789 2317
rect 4847 2303 4861 2317
rect 4871 2303 4885 2317
rect 36431 2303 36445 2317
rect 36455 2303 36469 2317
rect 39935 2303 39949 2317
rect 39959 2303 39973 2317
rect 44327 2303 44341 2317
rect 44351 2303 44365 2317
rect 50135 2303 50149 2317
rect 50159 2303 50173 2317
rect 51383 2303 51397 2317
rect 4751 2279 4765 2293
rect 5495 2279 5509 2293
rect 15119 2279 15133 2293
rect 15143 2279 15157 2293
rect 44615 2279 44629 2293
rect 44951 2279 44965 2293
rect 45047 2279 45061 2293
rect 47399 2279 47413 2293
rect 51503 2279 51517 2293
rect 4607 2255 4621 2269
rect 10439 2255 10453 2269
rect 10463 2255 10477 2269
rect 15455 2255 15469 2269
rect 15479 2255 15493 2269
rect 21383 2255 21397 2269
rect 24935 2255 24949 2269
rect 24959 2255 24973 2269
rect 43799 2255 43813 2269
rect 46967 2255 46981 2269
rect 51599 2255 51613 2269
rect 51671 2255 51685 2269
rect 51719 2255 51733 2269
rect 4559 2231 4573 2245
rect 43487 2231 43501 2245
rect 43511 2231 43525 2245
rect 50855 2231 50869 2245
rect 50879 2231 50893 2245
rect 51359 2231 51373 2245
rect 51383 2231 51397 2245
rect 51863 2231 51877 2245
rect 4199 2207 4213 2221
rect 8279 2207 8293 2221
rect 8303 2207 8317 2221
rect 12047 2207 12061 2221
rect 21983 2207 21997 2221
rect 36335 2207 36349 2221
rect 36359 2207 36373 2221
rect 36383 2207 36397 2221
rect 36719 2207 36733 2221
rect 36815 2207 36829 2221
rect 38231 2207 38245 2221
rect 38687 2207 38701 2221
rect 42671 2207 42685 2221
rect 42695 2207 42709 2221
rect 49679 2207 49693 2221
rect 51983 2207 51997 2221
rect 47 2183 61 2197
rect 71 2183 85 2197
rect 95 2183 109 2197
rect 119 2183 133 2197
rect 143 2183 157 2197
rect 167 2183 181 2197
rect 191 2183 205 2197
rect 215 2183 229 2197
rect 239 2183 253 2197
rect 263 2183 277 2197
rect 287 2183 301 2197
rect 311 2183 325 2197
rect 335 2183 349 2197
rect 359 2183 373 2197
rect 383 2183 397 2197
rect 407 2183 421 2197
rect 431 2183 445 2197
rect 455 2183 469 2197
rect 479 2183 493 2197
rect 503 2183 517 2197
rect 527 2183 541 2197
rect 551 2183 565 2197
rect 575 2183 589 2197
rect 599 2183 613 2197
rect 623 2183 637 2197
rect 647 2183 661 2197
rect 671 2183 685 2197
rect 695 2183 709 2197
rect 719 2183 733 2197
rect 743 2183 757 2197
rect 767 2183 781 2197
rect 791 2183 805 2197
rect 815 2183 829 2197
rect 839 2183 853 2197
rect 863 2183 877 2197
rect 887 2183 901 2197
rect 911 2183 925 2197
rect 935 2183 949 2197
rect 959 2183 973 2197
rect 983 2183 997 2197
rect 1007 2183 1021 2197
rect 1031 2183 1045 2197
rect 1055 2183 1069 2197
rect 1079 2183 1093 2197
rect 1103 2183 1117 2197
rect 1127 2183 1141 2197
rect 1151 2183 1165 2197
rect 1175 2183 1189 2197
rect 1199 2183 1213 2197
rect 1223 2183 1237 2197
rect 1247 2183 1261 2197
rect 1271 2183 1285 2197
rect 1295 2183 1309 2197
rect 1319 2183 1333 2197
rect 1343 2183 1357 2197
rect 1367 2183 1381 2197
rect 3983 2183 3997 2197
rect 21719 2183 21733 2197
rect 28799 2183 28813 2197
rect 30599 2183 30613 2197
rect 39983 2183 39997 2197
rect 40703 2183 40717 2197
rect 41255 2183 41269 2197
rect 47663 2183 47677 2197
rect 52103 2183 52117 2197
rect 47 2135 61 2149
rect 71 2135 85 2149
rect 95 2135 109 2149
rect 119 2135 133 2149
rect 143 2135 157 2149
rect 167 2135 181 2149
rect 191 2135 205 2149
rect 215 2135 229 2149
rect 239 2135 253 2149
rect 263 2135 277 2149
rect 287 2135 301 2149
rect 311 2135 325 2149
rect 335 2135 349 2149
rect 359 2135 373 2149
rect 383 2135 397 2149
rect 407 2135 421 2149
rect 431 2135 445 2149
rect 455 2135 469 2149
rect 479 2135 493 2149
rect 503 2135 517 2149
rect 527 2135 541 2149
rect 551 2135 565 2149
rect 575 2135 589 2149
rect 599 2135 613 2149
rect 623 2135 637 2149
rect 647 2135 661 2149
rect 671 2135 685 2149
rect 695 2135 709 2149
rect 719 2135 733 2149
rect 743 2135 757 2149
rect 767 2135 781 2149
rect 791 2135 805 2149
rect 815 2135 829 2149
rect 839 2135 853 2149
rect 863 2135 877 2149
rect 887 2135 901 2149
rect 911 2135 925 2149
rect 935 2135 949 2149
rect 959 2135 973 2149
rect 983 2135 997 2149
rect 1007 2135 1021 2149
rect 1031 2135 1045 2149
rect 1055 2135 1069 2149
rect 1079 2135 1093 2149
rect 1103 2135 1117 2149
rect 1127 2135 1141 2149
rect 1151 2135 1165 2149
rect 1175 2135 1189 2149
rect 1199 2135 1213 2149
rect 1223 2135 1237 2149
rect 1247 2135 1261 2149
rect 1271 2135 1285 2149
rect 1295 2135 1309 2149
rect 1319 2135 1333 2149
rect 1343 2135 1357 2149
rect 1367 2135 1381 2149
rect 3935 2159 3949 2173
rect 22727 2159 22741 2173
rect 52199 2159 52213 2173
rect 3431 2135 3445 2149
rect 3479 2135 3493 2149
rect 3575 2135 3589 2149
rect 8639 2135 8653 2149
rect 8663 2135 8677 2149
rect 47687 2135 47701 2149
rect 47711 2135 47725 2149
rect 49367 2135 49381 2149
rect 52319 2135 52333 2149
rect 3407 2111 3421 2125
rect 9311 2111 9325 2125
rect 9335 2111 9349 2125
rect 13751 2111 13765 2125
rect 13775 2111 13789 2125
rect 18503 2111 18517 2125
rect 18527 2111 18541 2125
rect 28727 2111 28741 2125
rect 28751 2111 28765 2125
rect 42431 2111 42445 2125
rect 42455 2111 42469 2125
rect 51191 2111 51205 2125
rect 51407 2111 51421 2125
rect 52439 2111 52453 2125
rect 3215 2087 3229 2101
rect 3263 2087 3277 2101
rect 3287 2087 3301 2101
rect 3359 2087 3373 2101
rect 3383 2087 3397 2101
rect 6239 2087 6253 2101
rect 6263 2087 6277 2101
rect 27743 2087 27757 2101
rect 27767 2087 27781 2101
rect 34871 2087 34885 2101
rect 34895 2087 34909 2101
rect 44231 2087 44245 2101
rect 44423 2087 44437 2101
rect 52559 2087 52573 2101
rect 3119 2063 3133 2077
rect 3167 2063 3181 2077
rect 3191 2063 3205 2077
rect 8495 2063 8509 2077
rect 8519 2063 8533 2077
rect 10895 2063 10909 2077
rect 10919 2063 10933 2077
rect 45839 2063 45853 2077
rect 45863 2063 45877 2077
rect 52487 2063 52501 2077
rect 52679 2063 52693 2077
rect 3095 2039 3109 2053
rect 8399 2039 8413 2053
rect 8423 2039 8437 2053
rect 45311 2039 45325 2053
rect 45335 2039 45349 2053
rect 52799 2039 52813 2053
rect 3071 2015 3085 2029
rect 22199 2015 22213 2029
rect 38159 2015 38173 2029
rect 38183 2015 38197 2029
rect 40535 2015 40549 2029
rect 40559 2015 40573 2029
rect 48455 2015 48469 2029
rect 48479 2015 48493 2029
rect 49175 2015 49189 2029
rect 50183 2015 50197 2029
rect 52895 2015 52909 2029
rect 2975 1991 2989 2005
rect 3023 1991 3037 2005
rect 3047 1991 3061 2005
rect 11855 1991 11869 2005
rect 48167 1991 48181 2005
rect 49751 1991 49765 2005
rect 53015 1991 53029 2005
rect 2951 1967 2965 1981
rect 6359 1967 6373 1981
rect 6383 1967 6397 1981
rect 25127 1967 25141 1981
rect 25151 1967 25165 1981
rect 51839 1967 51853 1981
rect 51863 1967 51877 1981
rect 53135 1967 53149 1981
rect 47 1943 61 1957
rect 71 1943 85 1957
rect 95 1943 109 1957
rect 119 1943 133 1957
rect 143 1943 157 1957
rect 167 1943 181 1957
rect 191 1943 205 1957
rect 215 1943 229 1957
rect 239 1943 253 1957
rect 263 1943 277 1957
rect 287 1943 301 1957
rect 311 1943 325 1957
rect 335 1943 349 1957
rect 359 1943 373 1957
rect 383 1943 397 1957
rect 407 1943 421 1957
rect 431 1943 445 1957
rect 455 1943 469 1957
rect 479 1943 493 1957
rect 503 1943 517 1957
rect 527 1943 541 1957
rect 551 1943 565 1957
rect 575 1943 589 1957
rect 599 1943 613 1957
rect 623 1943 637 1957
rect 647 1943 661 1957
rect 671 1943 685 1957
rect 695 1943 709 1957
rect 719 1943 733 1957
rect 743 1943 757 1957
rect 767 1943 781 1957
rect 791 1943 805 1957
rect 815 1943 829 1957
rect 839 1943 853 1957
rect 863 1943 877 1957
rect 887 1943 901 1957
rect 911 1943 925 1957
rect 935 1943 949 1957
rect 959 1943 973 1957
rect 983 1943 997 1957
rect 1007 1943 1021 1957
rect 1031 1943 1045 1957
rect 1055 1943 1069 1957
rect 1079 1943 1093 1957
rect 1103 1943 1117 1957
rect 1127 1943 1141 1957
rect 1151 1943 1165 1957
rect 1175 1943 1189 1957
rect 1199 1943 1213 1957
rect 1223 1943 1237 1957
rect 1247 1943 1261 1957
rect 1271 1943 1285 1957
rect 1295 1943 1309 1957
rect 1319 1943 1333 1957
rect 1343 1943 1357 1957
rect 1367 1943 1381 1957
rect 1391 1943 1405 1957
rect 2927 1943 2941 1957
rect 30575 1943 30589 1957
rect 33623 1943 33637 1957
rect 35927 1943 35941 1957
rect 35951 1943 35965 1957
rect 40319 1943 40333 1957
rect 40343 1943 40357 1957
rect 46919 1943 46933 1957
rect 46943 1943 46957 1957
rect 50087 1943 50101 1957
rect 53231 1943 53245 1957
rect 47 1895 61 1909
rect 71 1895 85 1909
rect 95 1895 109 1909
rect 119 1895 133 1909
rect 143 1895 157 1909
rect 167 1895 181 1909
rect 191 1895 205 1909
rect 215 1895 229 1909
rect 239 1895 253 1909
rect 263 1895 277 1909
rect 287 1895 301 1909
rect 311 1895 325 1909
rect 335 1895 349 1909
rect 359 1895 373 1909
rect 383 1895 397 1909
rect 407 1895 421 1909
rect 431 1895 445 1909
rect 455 1895 469 1909
rect 479 1895 493 1909
rect 503 1895 517 1909
rect 527 1895 541 1909
rect 551 1895 565 1909
rect 575 1895 589 1909
rect 599 1895 613 1909
rect 623 1895 637 1909
rect 647 1895 661 1909
rect 671 1895 685 1909
rect 695 1895 709 1909
rect 719 1895 733 1909
rect 743 1895 757 1909
rect 767 1895 781 1909
rect 791 1895 805 1909
rect 815 1895 829 1909
rect 839 1895 853 1909
rect 863 1895 877 1909
rect 887 1895 901 1909
rect 911 1895 925 1909
rect 935 1895 949 1909
rect 959 1895 973 1909
rect 983 1895 997 1909
rect 1007 1895 1021 1909
rect 1031 1895 1045 1909
rect 1055 1895 1069 1909
rect 1079 1895 1093 1909
rect 1103 1895 1117 1909
rect 1127 1895 1141 1909
rect 1151 1895 1165 1909
rect 1175 1895 1189 1909
rect 1199 1895 1213 1909
rect 1223 1895 1237 1909
rect 1247 1895 1261 1909
rect 1271 1895 1285 1909
rect 1295 1895 1309 1909
rect 1319 1895 1333 1909
rect 1343 1895 1357 1909
rect 1367 1895 1381 1909
rect 1391 1895 1405 1909
rect 2831 1919 2845 1933
rect 2879 1919 2893 1933
rect 2903 1919 2917 1933
rect 21239 1919 21253 1933
rect 21263 1919 21277 1933
rect 25343 1919 25357 1933
rect 25367 1919 25381 1933
rect 28871 1919 28885 1933
rect 32831 1919 32845 1933
rect 42887 1919 42901 1933
rect 44087 1919 44101 1933
rect 52607 1919 52621 1933
rect 52727 1919 52741 1933
rect 53375 1919 53389 1933
rect 2807 1895 2821 1909
rect 5927 1895 5941 1909
rect 5951 1895 5965 1909
rect 11159 1895 11173 1909
rect 11183 1895 11197 1909
rect 28343 1895 28357 1909
rect 28367 1895 28381 1909
rect 53471 1895 53485 1909
rect 2783 1871 2797 1885
rect 11735 1871 11749 1885
rect 22031 1871 22045 1885
rect 22055 1871 22069 1885
rect 30167 1871 30181 1885
rect 30191 1871 30205 1885
rect 36743 1871 36757 1885
rect 38999 1871 39013 1885
rect 42983 1871 42997 1885
rect 44735 1871 44749 1885
rect 45719 1871 45733 1885
rect 45791 1871 45805 1885
rect 45911 1871 45925 1885
rect 52871 1871 52885 1885
rect 52895 1871 52909 1885
rect 53543 1871 53557 1885
rect 2663 1847 2677 1861
rect 2735 1847 2749 1861
rect 2759 1847 2773 1861
rect 24647 1847 24661 1861
rect 27839 1847 27853 1861
rect 27863 1847 27877 1861
rect 39815 1847 39829 1861
rect 42503 1847 42517 1861
rect 48623 1847 48637 1861
rect 51287 1847 51301 1861
rect 51431 1847 51445 1861
rect 52007 1847 52021 1861
rect 53591 1847 53605 1861
rect 2567 1823 2581 1837
rect 2615 1823 2629 1837
rect 2639 1823 2653 1837
rect 3335 1823 3349 1837
rect 3359 1823 3373 1837
rect 6047 1823 6061 1837
rect 6071 1823 6085 1837
rect 8447 1823 8461 1837
rect 12527 1823 12541 1837
rect 12551 1823 12565 1837
rect 14519 1823 14533 1837
rect 14543 1823 14557 1837
rect 21527 1823 21541 1837
rect 21551 1823 21565 1837
rect 33791 1823 33805 1837
rect 33815 1823 33829 1837
rect 43535 1823 43549 1837
rect 43559 1823 43573 1837
rect 48551 1823 48565 1837
rect 48575 1823 48589 1837
rect 53111 1823 53125 1837
rect 53135 1823 53149 1837
rect 53639 1823 53653 1837
rect 2543 1799 2557 1813
rect 3239 1799 3253 1813
rect 3263 1799 3277 1813
rect 9455 1799 9469 1813
rect 9479 1799 9493 1813
rect 12479 1799 12493 1813
rect 14327 1799 14341 1813
rect 14351 1799 14365 1813
rect 53663 1799 53677 1813
rect 2399 1775 2413 1789
rect 9287 1775 9301 1789
rect 17663 1775 17677 1789
rect 53615 1775 53629 1789
rect 53639 1775 53653 1789
rect 53687 1775 53701 1789
rect 2351 1751 2365 1765
rect 53783 1751 53797 1765
rect 1991 1727 2005 1741
rect 3455 1727 3469 1741
rect 3479 1727 3493 1741
rect 9407 1727 9421 1741
rect 9455 1727 9469 1741
rect 15431 1727 15445 1741
rect 22511 1727 22525 1741
rect 43583 1727 43597 1741
rect 53903 1727 53917 1741
rect 47 1703 61 1717
rect 71 1703 85 1717
rect 95 1703 109 1717
rect 119 1703 133 1717
rect 143 1703 157 1717
rect 167 1703 181 1717
rect 191 1703 205 1717
rect 215 1703 229 1717
rect 239 1703 253 1717
rect 263 1703 277 1717
rect 287 1703 301 1717
rect 311 1703 325 1717
rect 335 1703 349 1717
rect 359 1703 373 1717
rect 383 1703 397 1717
rect 407 1703 421 1717
rect 431 1703 445 1717
rect 455 1703 469 1717
rect 479 1703 493 1717
rect 503 1703 517 1717
rect 527 1703 541 1717
rect 551 1703 565 1717
rect 575 1703 589 1717
rect 599 1703 613 1717
rect 623 1703 637 1717
rect 647 1703 661 1717
rect 671 1703 685 1717
rect 695 1703 709 1717
rect 719 1703 733 1717
rect 743 1703 757 1717
rect 767 1703 781 1717
rect 791 1703 805 1717
rect 815 1703 829 1717
rect 839 1703 853 1717
rect 863 1703 877 1717
rect 887 1703 901 1717
rect 911 1703 925 1717
rect 935 1703 949 1717
rect 959 1703 973 1717
rect 983 1703 997 1717
rect 1007 1703 1021 1717
rect 1031 1703 1045 1717
rect 1055 1703 1069 1717
rect 1079 1703 1093 1717
rect 1103 1703 1117 1717
rect 1127 1703 1141 1717
rect 1151 1703 1165 1717
rect 1175 1703 1189 1717
rect 1199 1703 1213 1717
rect 1223 1703 1237 1717
rect 1247 1703 1261 1717
rect 1271 1703 1285 1717
rect 1295 1703 1309 1717
rect 1319 1703 1333 1717
rect 1343 1703 1357 1717
rect 1367 1703 1381 1717
rect 1391 1703 1405 1717
rect 1415 1703 1429 1717
rect 1775 1703 1789 1717
rect 9095 1703 9109 1717
rect 13823 1703 13837 1717
rect 53999 1703 54013 1717
rect 47 1655 61 1669
rect 71 1655 85 1669
rect 95 1655 109 1669
rect 119 1655 133 1669
rect 143 1655 157 1669
rect 167 1655 181 1669
rect 191 1655 205 1669
rect 215 1655 229 1669
rect 239 1655 253 1669
rect 263 1655 277 1669
rect 287 1655 301 1669
rect 311 1655 325 1669
rect 335 1655 349 1669
rect 359 1655 373 1669
rect 383 1655 397 1669
rect 407 1655 421 1669
rect 431 1655 445 1669
rect 455 1655 469 1669
rect 479 1655 493 1669
rect 503 1655 517 1669
rect 527 1655 541 1669
rect 551 1655 565 1669
rect 575 1655 589 1669
rect 599 1655 613 1669
rect 623 1655 637 1669
rect 647 1655 661 1669
rect 671 1655 685 1669
rect 695 1655 709 1669
rect 719 1655 733 1669
rect 743 1655 757 1669
rect 767 1655 781 1669
rect 791 1655 805 1669
rect 815 1655 829 1669
rect 839 1655 853 1669
rect 863 1655 877 1669
rect 887 1655 901 1669
rect 911 1655 925 1669
rect 935 1655 949 1669
rect 959 1655 973 1669
rect 983 1655 997 1669
rect 1007 1655 1021 1669
rect 1031 1655 1045 1669
rect 1055 1655 1069 1669
rect 1079 1655 1093 1669
rect 1103 1655 1117 1669
rect 1127 1655 1141 1669
rect 1151 1655 1165 1669
rect 1175 1655 1189 1669
rect 1199 1655 1213 1669
rect 1223 1655 1237 1669
rect 1247 1655 1261 1669
rect 1271 1655 1285 1669
rect 1295 1655 1309 1669
rect 1319 1655 1333 1669
rect 1343 1655 1357 1669
rect 1367 1655 1381 1669
rect 1391 1655 1405 1669
rect 1415 1655 1429 1669
rect 1727 1679 1741 1693
rect 53639 1679 53653 1693
rect 53663 1679 53677 1693
rect 54071 1679 54085 1693
rect 9503 1655 9517 1669
rect 12503 1655 12517 1669
rect 46607 1655 46621 1669
rect 50207 1655 50221 1669
rect 54119 1655 54133 1669
rect 47 1463 61 1477
rect 71 1463 85 1477
rect 95 1463 109 1477
rect 119 1463 133 1477
rect 143 1463 157 1477
rect 167 1463 181 1477
rect 191 1463 205 1477
rect 215 1463 229 1477
rect 239 1463 253 1477
rect 263 1463 277 1477
rect 287 1463 301 1477
rect 311 1463 325 1477
rect 335 1463 349 1477
rect 359 1463 373 1477
rect 383 1463 397 1477
rect 407 1463 421 1477
rect 431 1463 445 1477
rect 455 1463 469 1477
rect 479 1463 493 1477
rect 503 1463 517 1477
rect 527 1463 541 1477
rect 551 1463 565 1477
rect 575 1463 589 1477
rect 599 1463 613 1477
rect 623 1463 637 1477
rect 647 1463 661 1477
rect 671 1463 685 1477
rect 695 1463 709 1477
rect 719 1463 733 1477
rect 743 1463 757 1477
rect 767 1463 781 1477
rect 791 1463 805 1477
rect 815 1463 829 1477
rect 839 1463 853 1477
rect 863 1463 877 1477
rect 887 1463 901 1477
rect 911 1463 925 1477
rect 935 1463 949 1477
rect 959 1463 973 1477
rect 983 1463 997 1477
rect 1007 1463 1021 1477
rect 1031 1463 1045 1477
rect 1055 1463 1069 1477
rect 1079 1463 1093 1477
rect 1103 1463 1117 1477
rect 1127 1463 1141 1477
rect 1151 1463 1165 1477
rect 1175 1463 1189 1477
rect 1199 1463 1213 1477
rect 1223 1463 1237 1477
rect 1247 1463 1261 1477
rect 46895 1631 46909 1645
rect 49199 1631 49213 1645
rect 54215 1631 54229 1645
rect 9383 1607 9397 1621
rect 9431 1607 9445 1621
rect 35639 1607 35653 1621
rect 35663 1607 35677 1621
rect 41279 1607 41293 1621
rect 41303 1607 41317 1621
rect 42263 1607 42277 1621
rect 45095 1607 45109 1621
rect 45119 1607 45133 1621
rect 48983 1607 48997 1621
rect 49775 1607 49789 1621
rect 51527 1607 51541 1621
rect 54095 1607 54109 1621
rect 54119 1607 54133 1621
rect 54167 1607 54181 1621
rect 54311 1607 54325 1621
rect 9191 1583 9205 1597
rect 9215 1583 9229 1597
rect 13199 1583 13213 1597
rect 13223 1583 13237 1597
rect 33575 1583 33589 1597
rect 33599 1583 33613 1597
rect 51143 1583 51157 1597
rect 51167 1583 51181 1597
rect 1367 1559 1381 1573
rect 5327 1559 5341 1573
rect 5351 1559 5365 1573
rect 9215 1559 9229 1573
rect 9239 1559 9253 1573
rect 41375 1559 41389 1573
rect 41399 1559 41413 1573
rect 41543 1559 41557 1573
rect 42863 1559 42877 1573
rect 42959 1559 42973 1573
rect 44495 1559 44509 1573
rect 48359 1559 48373 1573
rect 48383 1559 48397 1573
rect 54335 1559 54349 1573
rect 54359 1559 54373 1573
rect 8999 1535 9013 1549
rect 9023 1535 9037 1549
rect 44159 1535 44173 1549
rect 44183 1535 44197 1549
rect 51695 1535 51709 1549
rect 51719 1535 51733 1549
rect 54407 1535 54421 1549
rect 8711 1511 8725 1525
rect 8735 1511 8749 1525
rect 8975 1511 8989 1525
rect 9167 1511 9181 1525
rect 9359 1511 9373 1525
rect 12863 1511 12877 1525
rect 12887 1511 12901 1525
rect 27503 1511 27517 1525
rect 27527 1511 27541 1525
rect 32591 1511 32605 1525
rect 32615 1511 32629 1525
rect 39743 1511 39757 1525
rect 39767 1511 39781 1525
rect 43919 1511 43933 1525
rect 53351 1511 53365 1525
rect 53375 1511 53389 1525
rect 54551 1511 54565 1525
rect 33455 1487 33469 1501
rect 35495 1487 35509 1501
rect 44135 1487 44149 1501
rect 54671 1487 54685 1501
rect 54791 1463 54805 1477
rect 3311 1439 3325 1453
rect 40295 1439 40309 1453
rect 52055 1439 52069 1453
rect 54887 1439 54901 1453
rect 47 1415 61 1429
rect 71 1415 85 1429
rect 95 1415 109 1429
rect 119 1415 133 1429
rect 143 1415 157 1429
rect 167 1415 181 1429
rect 191 1415 205 1429
rect 215 1415 229 1429
rect 239 1415 253 1429
rect 263 1415 277 1429
rect 287 1415 301 1429
rect 311 1415 325 1429
rect 335 1415 349 1429
rect 359 1415 373 1429
rect 383 1415 397 1429
rect 407 1415 421 1429
rect 431 1415 445 1429
rect 455 1415 469 1429
rect 479 1415 493 1429
rect 503 1415 517 1429
rect 527 1415 541 1429
rect 551 1415 565 1429
rect 575 1415 589 1429
rect 599 1415 613 1429
rect 623 1415 637 1429
rect 647 1415 661 1429
rect 671 1415 685 1429
rect 695 1415 709 1429
rect 719 1415 733 1429
rect 743 1415 757 1429
rect 767 1415 781 1429
rect 791 1415 805 1429
rect 815 1415 829 1429
rect 839 1415 853 1429
rect 863 1415 877 1429
rect 887 1415 901 1429
rect 911 1415 925 1429
rect 935 1415 949 1429
rect 959 1415 973 1429
rect 983 1415 997 1429
rect 1007 1415 1021 1429
rect 1031 1415 1045 1429
rect 1055 1415 1069 1429
rect 1079 1415 1093 1429
rect 1103 1415 1117 1429
rect 1127 1415 1141 1429
rect 1151 1415 1165 1429
rect 1175 1415 1189 1429
rect 1199 1415 1213 1429
rect 1223 1415 1237 1429
rect 1247 1415 1261 1429
rect 5423 1415 5437 1429
rect 5447 1415 5461 1429
rect 9719 1415 9733 1429
rect 21335 1415 21349 1429
rect 21359 1415 21373 1429
rect 28511 1415 28525 1429
rect 42527 1415 42541 1429
rect 45479 1415 45493 1429
rect 46415 1415 46429 1429
rect 53207 1415 53221 1429
rect 53231 1415 53245 1429
rect 54287 1415 54301 1429
rect 54359 1415 54373 1429
rect 54983 1415 54997 1429
rect 47 1223 61 1237
rect 71 1223 85 1237
rect 95 1223 109 1237
rect 119 1223 133 1237
rect 143 1223 157 1237
rect 167 1223 181 1237
rect 191 1223 205 1237
rect 215 1223 229 1237
rect 239 1223 253 1237
rect 263 1223 277 1237
rect 287 1223 301 1237
rect 311 1223 325 1237
rect 335 1223 349 1237
rect 359 1223 373 1237
rect 383 1223 397 1237
rect 407 1223 421 1237
rect 431 1223 445 1237
rect 455 1223 469 1237
rect 479 1223 493 1237
rect 503 1223 517 1237
rect 527 1223 541 1237
rect 551 1223 565 1237
rect 575 1223 589 1237
rect 599 1223 613 1237
rect 623 1223 637 1237
rect 647 1223 661 1237
rect 671 1223 685 1237
rect 695 1223 709 1237
rect 719 1223 733 1237
rect 743 1223 757 1237
rect 767 1223 781 1237
rect 791 1223 805 1237
rect 815 1223 829 1237
rect 839 1223 853 1237
rect 863 1223 877 1237
rect 887 1223 901 1237
rect 911 1223 925 1237
rect 935 1223 949 1237
rect 959 1223 973 1237
rect 983 1223 997 1237
rect 1007 1223 1021 1237
rect 1031 1223 1045 1237
rect 19127 1391 19141 1405
rect 19151 1391 19165 1405
rect 28439 1391 28453 1405
rect 28463 1391 28477 1405
rect 37367 1391 37381 1405
rect 41879 1391 41893 1405
rect 41903 1391 41917 1405
rect 55079 1391 55093 1405
rect 5567 1367 5581 1381
rect 5591 1367 5605 1381
rect 11111 1367 11125 1381
rect 23735 1367 23749 1381
rect 23759 1367 23773 1381
rect 31631 1367 31645 1381
rect 35039 1367 35053 1381
rect 38039 1367 38053 1381
rect 46775 1367 46789 1381
rect 53759 1367 53773 1381
rect 53783 1367 53797 1381
rect 54263 1367 54277 1381
rect 54335 1367 54349 1381
rect 55175 1367 55189 1381
rect 23375 1343 23389 1357
rect 23399 1343 23413 1357
rect 45527 1343 45541 1357
rect 45551 1343 45565 1357
rect 47975 1343 47989 1357
rect 47999 1343 48013 1357
rect 53711 1343 53725 1357
rect 55295 1343 55309 1357
rect 4823 1319 4837 1333
rect 4847 1319 4861 1333
rect 10247 1319 10261 1333
rect 10271 1319 10285 1333
rect 12215 1319 12229 1333
rect 12239 1319 12253 1333
rect 32111 1319 32125 1333
rect 32135 1319 32149 1333
rect 40415 1319 40429 1333
rect 40439 1319 40453 1333
rect 47351 1319 47365 1333
rect 47375 1319 47389 1333
rect 49271 1319 49285 1333
rect 54767 1319 54781 1333
rect 54791 1319 54805 1333
rect 55415 1319 55429 1333
rect 12959 1295 12973 1309
rect 12983 1295 12997 1309
rect 20855 1295 20869 1309
rect 20879 1295 20893 1309
rect 23207 1295 23221 1309
rect 23591 1295 23605 1309
rect 23663 1295 23677 1309
rect 41951 1295 41965 1309
rect 44855 1295 44869 1309
rect 51815 1295 51829 1309
rect 53303 1295 53317 1309
rect 53855 1295 53869 1309
rect 54695 1295 54709 1309
rect 55535 1295 55549 1309
rect 9791 1271 9805 1285
rect 9815 1271 9829 1285
rect 33023 1271 33037 1285
rect 33047 1271 33061 1285
rect 38927 1271 38941 1285
rect 38951 1271 38965 1285
rect 41423 1271 41437 1285
rect 46031 1271 46045 1285
rect 46055 1271 46069 1285
rect 47135 1271 47149 1285
rect 47159 1271 47173 1285
rect 47183 1271 47197 1285
rect 51479 1271 51493 1285
rect 51503 1271 51517 1285
rect 52175 1271 52189 1285
rect 52199 1271 52213 1285
rect 54047 1271 54061 1285
rect 54071 1271 54085 1285
rect 54143 1271 54157 1285
rect 55631 1271 55645 1285
rect 5663 1247 5677 1261
rect 5687 1247 5701 1261
rect 24095 1247 24109 1261
rect 24119 1247 24133 1261
rect 27383 1247 27397 1261
rect 43823 1247 43837 1261
rect 55151 1247 55165 1261
rect 55175 1247 55189 1261
rect 55751 1247 55765 1261
rect 11495 1223 11509 1237
rect 11519 1223 11533 1237
rect 27407 1223 27421 1237
rect 27431 1223 27445 1237
rect 29159 1223 29173 1237
rect 38447 1223 38461 1237
rect 40967 1223 40981 1237
rect 40991 1223 41005 1237
rect 46439 1223 46453 1237
rect 46463 1223 46477 1237
rect 49607 1223 49621 1237
rect 49631 1223 49645 1237
rect 53831 1223 53845 1237
rect 55679 1223 55693 1237
rect 55847 1223 55861 1237
rect 20471 1199 20485 1213
rect 31175 1199 31189 1213
rect 35807 1199 35821 1213
rect 37511 1199 37525 1213
rect 38807 1199 38821 1213
rect 40103 1199 40117 1213
rect 45503 1199 45517 1213
rect 47903 1199 47917 1213
rect 49295 1199 49309 1213
rect 54839 1199 54853 1213
rect 47 1175 61 1189
rect 71 1175 85 1189
rect 95 1175 109 1189
rect 119 1175 133 1189
rect 143 1175 157 1189
rect 167 1175 181 1189
rect 191 1175 205 1189
rect 215 1175 229 1189
rect 239 1175 253 1189
rect 263 1175 277 1189
rect 287 1175 301 1189
rect 311 1175 325 1189
rect 335 1175 349 1189
rect 359 1175 373 1189
rect 383 1175 397 1189
rect 407 1175 421 1189
rect 431 1175 445 1189
rect 455 1175 469 1189
rect 479 1175 493 1189
rect 503 1175 517 1189
rect 527 1175 541 1189
rect 551 1175 565 1189
rect 575 1175 589 1189
rect 599 1175 613 1189
rect 623 1175 637 1189
rect 647 1175 661 1189
rect 671 1175 685 1189
rect 695 1175 709 1189
rect 719 1175 733 1189
rect 743 1175 757 1189
rect 767 1175 781 1189
rect 791 1175 805 1189
rect 815 1175 829 1189
rect 839 1175 853 1189
rect 863 1175 877 1189
rect 887 1175 901 1189
rect 911 1175 925 1189
rect 935 1175 949 1189
rect 959 1175 973 1189
rect 983 1175 997 1189
rect 1007 1175 1021 1189
rect 1031 1175 1045 1189
rect 9911 1175 9925 1189
rect 9935 1175 9949 1189
rect 14999 1175 15013 1189
rect 15023 1175 15037 1189
rect 23231 1175 23245 1189
rect 23255 1175 23269 1189
rect 31247 1175 31261 1189
rect 31271 1175 31285 1189
rect 31655 1175 31669 1189
rect 37319 1175 37333 1189
rect 37343 1175 37357 1189
rect 37559 1175 37573 1189
rect 37583 1175 37597 1189
rect 42095 1175 42109 1189
rect 42119 1175 42133 1189
rect 47807 1175 47821 1189
rect 47831 1175 47845 1189
rect 49871 1175 49885 1189
rect 55055 1175 55069 1189
rect 55079 1175 55093 1189
rect 55919 1175 55933 1189
rect 56039 1199 56053 1213
rect 56471 1199 56485 1213
rect 56639 1175 56653 1189
rect 47 983 61 997
rect 71 983 85 997
rect 95 983 109 997
rect 119 983 133 997
rect 143 983 157 997
rect 167 983 181 997
rect 191 983 205 997
rect 215 983 229 997
rect 239 983 253 997
rect 263 983 277 997
rect 287 983 301 997
rect 311 983 325 997
rect 335 983 349 997
rect 359 983 373 997
rect 383 983 397 997
rect 407 983 421 997
rect 431 983 445 997
rect 455 983 469 997
rect 479 983 493 997
rect 503 983 517 997
rect 527 983 541 997
rect 551 983 565 997
rect 575 983 589 997
rect 599 983 613 997
rect 623 983 637 997
rect 647 983 661 997
rect 671 983 685 997
rect 695 983 709 997
rect 719 983 733 997
rect 743 983 757 997
rect 767 983 781 997
rect 791 983 805 997
rect 815 983 829 997
rect 10055 1151 10069 1165
rect 10079 1151 10093 1165
rect 19631 1151 19645 1165
rect 41591 1151 41605 1165
rect 41615 1151 41629 1165
rect 42143 1151 42157 1165
rect 44879 1151 44893 1165
rect 44903 1151 44917 1165
rect 48647 1151 48661 1165
rect 48671 1151 48685 1165
rect 52703 1151 52717 1165
rect 56687 1151 56701 1165
rect 43031 1127 43045 1141
rect 43055 1127 43069 1141
rect 49943 1127 49957 1141
rect 49967 1127 49981 1141
rect 50303 1127 50317 1141
rect 51767 1127 51781 1141
rect 54071 1127 54085 1141
rect 56783 1127 56797 1141
rect 5879 1103 5893 1117
rect 23471 1103 23485 1117
rect 23495 1103 23509 1117
rect 29231 1103 29245 1117
rect 29255 1103 29269 1117
rect 39623 1103 39637 1117
rect 39647 1103 39661 1117
rect 42743 1103 42757 1117
rect 47447 1103 47461 1117
rect 47471 1103 47485 1117
rect 53159 1103 53173 1117
rect 55727 1103 55741 1117
rect 55751 1103 55765 1117
rect 56879 1103 56893 1117
rect 7943 1079 7957 1093
rect 7967 1079 7981 1093
rect 30887 1079 30901 1093
rect 30911 1079 30925 1093
rect 38063 1079 38077 1093
rect 38087 1079 38101 1093
rect 40631 1079 40645 1093
rect 40655 1079 40669 1093
rect 44447 1079 44461 1093
rect 44471 1079 44485 1093
rect 46583 1079 46597 1093
rect 52415 1079 52429 1093
rect 52439 1079 52453 1093
rect 56975 1079 56989 1093
rect 2855 1055 2869 1069
rect 2879 1055 2893 1069
rect 4799 1055 4813 1069
rect 8471 1055 8485 1069
rect 10991 1055 11005 1069
rect 11759 1055 11773 1069
rect 21431 1055 21445 1069
rect 21455 1055 21469 1069
rect 25031 1055 25045 1069
rect 25055 1055 25069 1069
rect 27167 1055 27181 1069
rect 30863 1055 30877 1069
rect 41759 1055 41773 1069
rect 51911 1055 51925 1069
rect 57095 1055 57109 1069
rect 8063 1031 8077 1045
rect 8087 1031 8101 1045
rect 21143 1031 21157 1045
rect 21167 1031 21181 1045
rect 29063 1031 29077 1045
rect 44111 1031 44125 1045
rect 45695 1031 45709 1045
rect 46271 1031 46285 1045
rect 51095 1031 51109 1045
rect 53399 1031 53413 1045
rect 54527 1031 54541 1045
rect 54551 1031 54565 1045
rect 57167 1031 57181 1045
rect 8183 1007 8197 1021
rect 8207 1007 8221 1021
rect 44543 1007 44557 1021
rect 44567 1007 44581 1021
rect 48695 1007 48709 1021
rect 51119 1007 51133 1021
rect 53519 1007 53533 1021
rect 53543 1007 53557 1021
rect 55511 1007 55525 1021
rect 55535 1007 55549 1021
rect 57191 1007 57205 1021
rect 5807 983 5821 997
rect 5831 983 5845 997
rect 10583 983 10597 997
rect 10607 983 10621 997
rect 12671 983 12685 997
rect 12695 983 12709 997
rect 38735 983 38749 997
rect 38759 983 38773 997
rect 49223 983 49237 997
rect 49247 983 49261 997
rect 53927 983 53941 997
rect 57287 983 57301 997
rect 20519 959 20533 973
rect 28991 959 29005 973
rect 34271 959 34285 973
rect 37271 959 37285 973
rect 49583 959 49597 973
rect 54719 959 54733 973
rect 55031 959 55045 973
rect 55799 959 55813 973
rect 55895 959 55909 973
rect 57359 959 57373 973
rect 47 935 61 949
rect 71 935 85 949
rect 95 935 109 949
rect 119 935 133 949
rect 143 935 157 949
rect 167 935 181 949
rect 191 935 205 949
rect 215 935 229 949
rect 239 935 253 949
rect 263 935 277 949
rect 287 935 301 949
rect 311 935 325 949
rect 335 935 349 949
rect 359 935 373 949
rect 383 935 397 949
rect 407 935 421 949
rect 431 935 445 949
rect 455 935 469 949
rect 479 935 493 949
rect 503 935 517 949
rect 527 935 541 949
rect 551 935 565 949
rect 575 935 589 949
rect 599 935 613 949
rect 623 935 637 949
rect 647 935 661 949
rect 671 935 685 949
rect 695 935 709 949
rect 719 935 733 949
rect 743 935 757 949
rect 767 935 781 949
rect 791 935 805 949
rect 815 935 829 949
rect 11639 935 11653 949
rect 11663 935 11677 949
rect 20183 935 20197 949
rect 38591 935 38605 949
rect 44303 935 44317 949
rect 46727 935 46741 949
rect 48911 935 48925 949
rect 52631 935 52645 949
rect 55439 935 55453 949
rect 57119 935 57133 949
rect 57383 935 57397 949
rect 47 743 61 757
rect 71 743 85 757
rect 95 743 109 757
rect 119 743 133 757
rect 143 743 157 757
rect 167 743 181 757
rect 191 743 205 757
rect 215 743 229 757
rect 239 743 253 757
rect 263 743 277 757
rect 287 743 301 757
rect 311 743 325 757
rect 335 743 349 757
rect 359 743 373 757
rect 383 743 397 757
rect 407 743 421 757
rect 431 743 445 757
rect 455 743 469 757
rect 479 743 493 757
rect 503 743 517 757
rect 527 743 541 757
rect 551 743 565 757
rect 575 743 589 757
rect 599 743 613 757
rect 623 743 637 757
rect 10151 911 10165 925
rect 10175 911 10189 925
rect 42911 911 42925 925
rect 42935 911 42949 925
rect 50039 911 50053 925
rect 50063 911 50077 925
rect 56903 911 56917 925
rect 57479 911 57493 925
rect 13415 887 13429 901
rect 13439 887 13453 901
rect 36863 887 36877 901
rect 36887 887 36901 901
rect 46391 887 46405 901
rect 52535 887 52549 901
rect 52559 887 52573 901
rect 56711 887 56725 901
rect 57599 887 57613 901
rect 1151 863 1165 877
rect 8903 863 8917 877
rect 17879 863 17893 877
rect 17903 863 17917 877
rect 18383 863 18397 877
rect 18407 863 18421 877
rect 33983 863 33997 877
rect 40679 863 40693 877
rect 42623 863 42637 877
rect 46223 863 46237 877
rect 46247 863 46261 877
rect 50327 863 50341 877
rect 50351 863 50365 877
rect 54479 863 54493 877
rect 54575 863 54589 877
rect 57647 863 57661 877
rect 57695 863 57709 877
rect 743 839 757 853
rect 5087 839 5101 853
rect 5111 839 5125 853
rect 9023 839 9037 853
rect 9047 839 9061 853
rect 10487 839 10501 853
rect 10511 839 10525 853
rect 30647 839 30661 853
rect 30671 839 30685 853
rect 35543 839 35557 853
rect 35567 839 35581 853
rect 50231 839 50245 853
rect 50255 839 50269 853
rect 55391 839 55405 853
rect 55415 839 55429 853
rect 57815 839 57829 853
rect 13295 815 13309 829
rect 13319 815 13333 829
rect 19223 815 19237 829
rect 19247 815 19261 829
rect 28919 815 28933 829
rect 28943 815 28957 829
rect 32783 815 32797 829
rect 32807 815 32821 829
rect 37751 815 37765 829
rect 37775 815 37789 829
rect 41975 815 41989 829
rect 41999 815 42013 829
rect 49511 815 49525 829
rect 49535 815 49549 829
rect 55607 815 55621 829
rect 55631 815 55645 829
rect 57887 815 57901 829
rect 12071 791 12085 805
rect 12095 791 12109 805
rect 22751 791 22765 805
rect 22775 791 22789 805
rect 27935 791 27949 805
rect 27959 791 27973 805
rect 34415 791 34429 805
rect 34439 791 34453 805
rect 35063 791 35077 805
rect 35087 791 35101 805
rect 40031 791 40045 805
rect 40055 791 40069 805
rect 47039 791 47053 805
rect 47063 791 47077 805
rect 50111 791 50125 805
rect 53663 791 53677 805
rect 53687 791 53701 805
rect 57071 791 57085 805
rect 57095 791 57109 805
rect 57791 791 57805 805
rect 57815 791 57829 805
rect 57911 791 57925 805
rect 4967 767 4981 781
rect 4991 767 5005 781
rect 10391 767 10405 781
rect 10415 767 10429 781
rect 13103 767 13117 781
rect 13127 767 13141 781
rect 21191 767 21205 781
rect 24407 767 24421 781
rect 31055 767 31069 781
rect 34367 767 34381 781
rect 38975 767 38989 781
rect 39383 767 39397 781
rect 45191 767 45205 781
rect 45215 767 45229 781
rect 46655 767 46669 781
rect 46679 767 46693 781
rect 49703 767 49717 781
rect 49727 767 49741 781
rect 51791 767 51805 781
rect 57215 767 57229 781
rect 57335 767 57349 781
rect 57359 767 57373 781
rect 57935 767 57949 781
rect 11399 743 11413 757
rect 11423 743 11437 757
rect 29327 743 29341 757
rect 29351 743 29365 757
rect 33767 743 33781 757
rect 42191 743 42205 757
rect 42215 743 42229 757
rect 49319 743 49333 757
rect 49343 743 49357 757
rect 57263 743 57277 757
rect 57287 743 57301 757
rect 57671 743 57685 757
rect 57695 743 57709 757
rect 58031 743 58045 757
rect 23831 719 23845 733
rect 24191 719 24205 733
rect 45407 719 45421 733
rect 55703 719 55717 733
rect 57047 719 57061 733
rect 57407 719 57421 733
rect 57959 719 57973 733
rect 58127 719 58141 733
rect 47 695 61 709
rect 71 695 85 709
rect 95 695 109 709
rect 119 695 133 709
rect 143 695 157 709
rect 167 695 181 709
rect 191 695 205 709
rect 215 695 229 709
rect 239 695 253 709
rect 263 695 277 709
rect 287 695 301 709
rect 311 695 325 709
rect 335 695 349 709
rect 359 695 373 709
rect 383 695 397 709
rect 407 695 421 709
rect 431 695 445 709
rect 455 695 469 709
rect 479 695 493 709
rect 503 695 517 709
rect 527 695 541 709
rect 551 695 565 709
rect 575 695 589 709
rect 599 695 613 709
rect 623 695 637 709
rect 2999 695 3013 709
rect 3023 695 3037 709
rect 4943 695 4957 709
rect 27191 695 27205 709
rect 27215 695 27229 709
rect 27695 695 27709 709
rect 34511 695 34525 709
rect 34535 695 34549 709
rect 35471 695 35485 709
rect 39431 695 39445 709
rect 39455 695 39469 709
rect 50447 695 50461 709
rect 56447 695 56461 709
rect 56471 695 56485 709
rect 47 503 61 517
rect 71 503 85 517
rect 95 503 109 517
rect 119 503 133 517
rect 143 503 157 517
rect 167 503 181 517
rect 191 503 205 517
rect 215 503 229 517
rect 239 503 253 517
rect 263 503 277 517
rect 287 503 301 517
rect 311 503 325 517
rect 335 503 349 517
rect 359 503 373 517
rect 383 503 397 517
rect 407 503 421 517
rect 431 503 445 517
rect 3143 671 3157 685
rect 3167 671 3181 685
rect 11903 671 11917 685
rect 50279 671 50293 685
rect 54383 671 54397 685
rect 54407 671 54421 685
rect 55559 671 55573 685
rect 57455 671 57469 685
rect 57479 671 57493 685
rect 58199 671 58213 685
rect 58319 671 58333 685
rect 11783 647 11797 661
rect 11807 647 11821 661
rect 28631 647 28645 661
rect 28655 647 28669 661
rect 30815 647 30829 661
rect 30935 647 30949 661
rect 31079 647 31093 661
rect 31319 647 31333 661
rect 31535 647 31549 661
rect 36119 647 36133 661
rect 36143 647 36157 661
rect 37919 647 37933 661
rect 38327 647 38341 661
rect 38783 647 38797 661
rect 42791 647 42805 661
rect 42815 647 42829 661
rect 46007 647 46021 661
rect 46103 647 46117 661
rect 46295 647 46309 661
rect 51575 647 51589 661
rect 51599 647 51613 661
rect 51959 647 51973 661
rect 51983 647 51997 661
rect 53063 647 53077 661
rect 58391 647 58405 661
rect 11927 623 11941 637
rect 11951 623 11965 637
rect 19559 623 19573 637
rect 19583 623 19597 637
rect 22295 623 22309 637
rect 22319 623 22333 637
rect 22871 623 22885 637
rect 42311 623 42325 637
rect 42335 623 42349 637
rect 52823 623 52837 637
rect 53567 623 53581 637
rect 53591 623 53605 637
rect 54815 623 54829 637
rect 54911 623 54925 637
rect 55463 623 55477 637
rect 55871 623 55885 637
rect 58439 623 58453 637
rect 9575 599 9589 613
rect 11015 599 11029 613
rect 11039 599 11053 613
rect 20375 599 20389 613
rect 26255 599 26269 613
rect 26279 599 26293 613
rect 31487 599 31501 613
rect 31511 599 31525 613
rect 52655 599 52669 613
rect 52679 599 52693 613
rect 54863 599 54877 613
rect 54887 599 54901 613
rect 58079 599 58093 613
rect 58247 599 58261 613
rect 58559 599 58573 613
rect 527 575 541 589
rect 5999 575 6013 589
rect 8807 575 8821 589
rect 18095 575 18109 589
rect 56615 575 56629 589
rect 56639 575 56653 589
rect 57431 575 57445 589
rect 58055 575 58069 589
rect 58607 575 58621 589
rect 58655 575 58669 589
rect 20423 551 20437 565
rect 20447 551 20461 565
rect 36215 551 36229 565
rect 39575 551 39589 565
rect 43895 551 43909 565
rect 48791 551 48805 565
rect 49007 551 49021 565
rect 49103 551 49117 565
rect 51311 551 51325 565
rect 51887 551 51901 565
rect 52031 551 52045 565
rect 54455 551 54469 565
rect 55223 551 55237 565
rect 57311 551 57325 565
rect 57335 551 57349 565
rect 57623 551 57637 565
rect 58343 551 58357 565
rect 58703 551 58717 565
rect 41159 527 41173 541
rect 41183 527 41197 541
rect 45263 527 45277 541
rect 49031 527 49045 541
rect 49055 527 49069 541
rect 54599 527 54613 541
rect 55247 527 55261 541
rect 55319 527 55333 541
rect 57143 527 57157 541
rect 57167 527 57181 541
rect 57575 527 57589 541
rect 57599 527 57613 541
rect 58727 527 58741 541
rect 2591 503 2605 517
rect 2615 503 2629 517
rect 2687 503 2701 517
rect 5783 503 5797 517
rect 9863 503 9877 517
rect 10007 503 10021 517
rect 37823 503 37837 517
rect 41111 503 41125 517
rect 43247 503 43261 517
rect 43271 503 43285 517
rect 45575 503 45589 517
rect 49823 503 49837 517
rect 49847 503 49861 517
rect 56759 503 56773 517
rect 56783 503 56797 517
rect 57527 503 57541 517
rect 57863 503 57877 517
rect 57911 503 57925 517
rect 58775 503 58789 517
rect 14495 479 14509 493
rect 33239 479 33253 493
rect 36983 479 36997 493
rect 40919 479 40933 493
rect 47423 479 47437 493
rect 47759 479 47773 493
rect 53327 479 53341 493
rect 58175 479 58189 493
rect 58463 479 58477 493
rect 58583 479 58597 493
rect 58823 479 58837 493
rect 47 455 61 469
rect 71 455 85 469
rect 95 455 109 469
rect 119 455 133 469
rect 143 455 157 469
rect 167 455 181 469
rect 191 455 205 469
rect 215 455 229 469
rect 239 455 253 469
rect 263 455 277 469
rect 287 455 301 469
rect 311 455 325 469
rect 335 455 349 469
rect 359 455 373 469
rect 383 455 397 469
rect 407 455 421 469
rect 431 455 445 469
rect 2711 455 2725 469
rect 2735 455 2749 469
rect 14807 455 14821 469
rect 14831 455 14845 469
rect 27647 455 27661 469
rect 27671 455 27685 469
rect 44255 455 44269 469
rect 52367 455 52381 469
rect 56855 455 56869 469
rect 56879 455 56893 469
rect 58415 455 58429 469
rect 58439 455 58453 469
rect 58871 455 58885 469
rect 47 263 61 277
rect 71 263 85 277
rect 95 263 109 277
rect 119 263 133 277
rect 143 263 157 277
rect 167 263 181 277
rect 191 263 205 277
rect 215 263 229 277
rect 15647 431 15661 445
rect 15671 431 15685 445
rect 45983 431 45997 445
rect 48887 431 48901 445
rect 54647 431 54661 445
rect 54671 431 54685 445
rect 58943 431 58957 445
rect 15863 407 15877 421
rect 15887 407 15901 421
rect 23783 407 23797 421
rect 32879 407 32893 421
rect 35711 407 35725 421
rect 40607 407 40621 421
rect 47303 407 47317 421
rect 51743 407 51757 421
rect 55775 407 55789 421
rect 57239 407 57253 421
rect 58991 407 59005 421
rect 16079 383 16093 397
rect 16103 383 16117 397
rect 23087 383 23101 397
rect 23111 383 23125 397
rect 46511 383 46525 397
rect 47639 383 47653 397
rect 48287 383 48301 397
rect 48503 383 48517 397
rect 52247 383 52261 397
rect 57167 383 57181 397
rect 57191 383 57205 397
rect 59063 383 59077 397
rect 16295 359 16309 373
rect 16319 359 16333 373
rect 20903 359 20917 373
rect 46343 359 46357 373
rect 46367 359 46381 373
rect 48839 359 48853 373
rect 48863 359 48877 373
rect 49415 359 49429 373
rect 49439 359 49453 373
rect 57359 359 57373 373
rect 57383 359 57397 373
rect 58679 359 58693 373
rect 58727 359 58741 373
rect 58967 359 58981 373
rect 58991 359 59005 373
rect 59111 359 59125 373
rect 16511 335 16525 349
rect 16535 335 16549 349
rect 21911 335 21925 349
rect 21935 335 21949 349
rect 44831 335 44845 349
rect 45383 335 45397 349
rect 52991 335 53005 349
rect 53015 335 53029 349
rect 55271 335 55285 349
rect 55295 335 55309 349
rect 58631 335 58645 349
rect 58655 335 58669 349
rect 59159 335 59173 349
rect 14183 311 14197 325
rect 14207 311 14221 325
rect 15167 311 15181 325
rect 15503 311 15517 325
rect 15719 311 15733 325
rect 15935 311 15949 325
rect 16151 311 16165 325
rect 16367 311 16381 325
rect 16583 311 16597 325
rect 16799 311 16813 325
rect 17015 311 17029 325
rect 17231 311 17245 325
rect 17447 311 17461 325
rect 17471 311 17485 325
rect 32903 311 32917 325
rect 32927 311 32941 325
rect 35591 311 35605 325
rect 35687 311 35701 325
rect 35783 311 35797 325
rect 35879 311 35893 325
rect 36599 311 36613 325
rect 39143 311 39157 325
rect 39167 311 39181 325
rect 43439 311 43453 325
rect 43463 311 43477 325
rect 51239 311 51253 325
rect 51263 311 51277 325
rect 59087 311 59101 325
rect 59111 311 59125 325
rect 59207 311 59221 325
rect 16727 287 16741 301
rect 16751 287 16765 301
rect 20951 287 20965 301
rect 20975 287 20989 301
rect 24335 287 24349 301
rect 24359 287 24373 301
rect 49127 287 49141 301
rect 49151 287 49165 301
rect 53975 287 53989 301
rect 53999 287 54013 301
rect 54239 287 54253 301
rect 54311 287 54325 301
rect 56591 287 56605 301
rect 57743 287 57757 301
rect 58271 287 58285 301
rect 58919 287 58933 301
rect 58943 287 58957 301
rect 59039 287 59053 301
rect 59063 287 59077 301
rect 59303 287 59317 301
rect 16943 263 16957 277
rect 16967 263 16981 277
rect 22631 263 22645 277
rect 22655 263 22669 277
rect 26495 263 26509 277
rect 26519 263 26533 277
rect 42575 263 42589 277
rect 42599 263 42613 277
rect 43679 263 43693 277
rect 43847 263 43861 277
rect 43871 263 43885 277
rect 47567 263 47581 277
rect 47591 263 47605 277
rect 58295 263 58309 277
rect 58319 263 58333 277
rect 59351 263 59365 277
rect 30959 239 30973 253
rect 31223 239 31237 253
rect 31679 239 31693 253
rect 33191 239 33205 253
rect 33863 239 33877 253
rect 34751 239 34765 253
rect 42551 239 42565 253
rect 44639 239 44653 253
rect 51335 239 51349 253
rect 53087 239 53101 253
rect 53279 239 53293 253
rect 54935 239 54949 253
rect 59279 239 59293 253
rect 59303 239 59317 253
rect 59423 239 59437 253
rect 47 215 61 229
rect 71 215 85 229
rect 95 215 109 229
rect 119 215 133 229
rect 143 215 157 229
rect 167 215 181 229
rect 191 215 205 229
rect 215 215 229 229
rect 17159 215 17173 229
rect 17183 215 17197 229
rect 21407 215 21421 229
rect 23279 215 23293 229
rect 27143 215 27157 229
rect 34703 215 34717 229
rect 36191 215 36205 229
rect 38567 215 38581 229
rect 41471 215 41485 229
rect 41495 215 41509 229
rect 44687 215 44701 229
rect 44711 215 44725 229
rect 47327 215 47341 229
rect 49487 215 49501 229
rect 56951 215 56965 229
rect 56975 215 56989 229
rect 58751 215 58765 229
rect 58775 215 58789 229
rect 15311 191 15325 205
rect 15335 191 15349 205
rect 18863 191 18877 205
rect 20711 191 20725 205
rect 20807 191 20821 205
rect 21287 191 21301 205
rect 24695 191 24709 205
rect 24719 191 24733 205
rect 33119 191 33133 205
rect 33143 191 33157 205
rect 35423 191 35437 205
rect 35447 191 35461 205
rect 48743 191 48757 205
rect 48767 191 48781 205
rect 48815 191 48829 205
rect 50999 191 51013 205
rect 52127 191 52141 205
rect 53879 191 53893 205
rect 53903 191 53917 205
rect 56807 191 56821 205
rect 58847 191 58861 205
rect 58871 191 58885 205
rect 59447 191 59461 205
rect 59543 191 59557 205
rect 17375 167 17389 181
rect 17399 167 17413 181
rect 33431 167 33445 181
rect 36527 167 36541 181
rect 36551 167 36565 181
rect 41063 167 41077 181
rect 41087 167 41101 181
rect 44783 167 44797 181
rect 44807 167 44821 181
rect 48047 167 48061 181
rect 52775 167 52789 181
rect 52799 167 52813 181
rect 54959 167 54973 181
rect 54983 167 54997 181
rect 55103 167 55117 181
rect 58103 167 58117 181
rect 58127 167 58141 181
rect 58151 167 58165 181
rect 58487 167 58501 181
rect 59591 167 59605 181
rect 17591 143 17605 157
rect 17615 143 17629 157
rect 21791 143 21805 157
rect 21815 143 21829 157
rect 22487 143 22501 157
rect 24767 143 24781 157
rect 25079 143 25093 157
rect 26639 143 26653 157
rect 31127 143 31141 157
rect 31151 143 31165 157
rect 32015 143 32029 157
rect 32039 143 32053 157
rect 39239 143 39253 157
rect 39263 143 39277 157
rect 50807 143 50821 157
rect 50831 143 50845 157
rect 52295 143 52309 157
rect 52319 143 52333 157
rect 54191 143 54205 157
rect 54215 143 54229 157
rect 56639 143 56653 157
rect 56735 143 56749 157
rect 56831 143 56845 157
rect 57719 143 57733 157
rect 59639 143 59653 157
rect 6191 119 6205 133
rect 17807 119 17821 133
rect 17831 119 17845 133
rect 25535 119 25549 133
rect 25559 119 25573 133
rect 27359 119 27373 133
rect 29183 119 29197 133
rect 34607 119 34621 133
rect 34631 119 34645 133
rect 40847 119 40861 133
rect 40871 119 40885 133
rect 46535 119 46549 133
rect 46559 119 46573 133
rect 53447 119 53461 133
rect 53471 119 53485 133
rect 56663 119 56677 133
rect 56687 119 56701 133
rect 57911 119 57925 133
rect 57935 119 57949 133
rect 57983 119 57997 133
rect 59519 119 59533 133
rect 59543 119 59557 133
rect 119 95 133 109
rect 5207 95 5221 109
rect 5231 95 5245 109
rect 8735 95 8749 109
rect 8759 95 8773 109
rect 30527 95 30541 109
rect 30551 95 30565 109
rect 40751 95 40765 109
rect 40775 95 40789 109
rect 52079 95 52093 109
rect 52103 95 52117 109
rect 53543 95 53557 109
rect 57503 95 57517 109
rect 57839 95 57853 109
rect 57887 95 57901 109
rect 59687 95 59701 109
rect 59759 95 59773 109
rect 6407 71 6421 85
rect 13967 71 13981 85
rect 13991 71 14005 85
rect 14111 71 14125 85
rect 15239 71 15253 85
rect 15575 71 15589 85
rect 15791 71 15805 85
rect 16007 71 16021 85
rect 16223 71 16237 85
rect 16439 71 16453 85
rect 16655 71 16669 85
rect 16871 71 16885 85
rect 17087 71 17101 85
rect 17303 71 17317 85
rect 17519 71 17533 85
rect 17735 71 17749 85
rect 17951 71 17965 85
rect 18167 71 18181 85
rect 22127 71 22141 85
rect 22151 71 22165 85
rect 23975 71 23989 85
rect 23999 71 24013 85
rect 24047 71 24061 85
rect 34199 71 34213 85
rect 34223 71 34237 85
rect 36479 71 36493 85
rect 39023 71 39037 85
rect 39047 71 39061 85
rect 39071 71 39085 85
rect 45143 71 45157 85
rect 48935 71 48949 85
rect 48959 71 48973 85
rect 49463 71 49477 85
rect 49895 71 49909 85
rect 52943 71 52957 85
rect 55823 71 55837 85
rect 55847 71 55861 85
rect 59567 71 59581 85
rect 59591 71 59605 85
rect 6095 47 6109 61
rect 18023 47 18037 61
rect 18047 47 18061 61
rect 20543 47 20557 61
rect 20567 47 20581 61
rect 21839 47 21853 61
rect 22943 47 22957 61
rect 28247 47 28261 61
rect 28271 47 28285 61
rect 35735 47 35749 61
rect 35759 47 35773 61
rect 40223 47 40237 61
rect 40247 47 40261 61
rect 47231 47 47245 61
rect 47255 47 47269 61
rect 48239 47 48253 61
rect 48263 47 48277 61
rect 48431 47 48445 61
rect 51647 47 51661 61
rect 55007 47 55021 61
rect 55343 47 55357 61
rect 57023 47 57037 61
rect 59327 47 59341 61
rect 59351 47 59365 61
rect 59807 47 59821 61
rect 59879 47 59893 61
rect 18263 23 18277 37
rect 18935 23 18949 37
rect 39551 23 39565 37
rect 45455 23 45469 37
rect 51071 23 51085 37
rect 58031 23 58045 37
rect 58391 23 58405 37
rect 58559 23 58573 37
rect 58823 23 58837 37
rect 59423 23 59437 37
rect 7751 -1 7765 13
rect 18239 -1 18253 13
rect 18911 -1 18925 13
rect 33215 -1 33229 13
rect 39527 -1 39541 13
rect 42383 -1 42397 13
rect 45431 -1 45445 13
rect 51047 -1 51061 13
rect 58007 -1 58021 13
rect 58367 -1 58381 13
rect 58535 -1 58549 13
rect 58799 -1 58813 13
rect 59399 -1 59413 13
rect 59927 -1 59941 13
<< metal2 >>
rect 48 15349 60 15383
rect 48 15109 60 15143
rect 72 15109 84 15143
rect 48 14869 60 14903
rect 72 14869 84 14903
rect 96 14869 108 14903
rect 48 14629 60 14663
rect 72 14629 84 14663
rect 96 14629 108 14663
rect 120 14629 132 14663
rect 48 14389 60 14423
rect 72 14389 84 14423
rect 96 14389 108 14423
rect 120 14389 132 14423
rect 144 14389 156 14423
rect 48 14149 60 14183
rect 72 14149 84 14183
rect 96 14149 108 14183
rect 120 14149 132 14183
rect 144 14149 156 14183
rect 168 14149 180 14183
rect 48 13909 60 13943
rect 72 13909 84 13943
rect 96 13909 108 13943
rect 120 13909 132 13943
rect 144 13909 156 13943
rect 168 13909 180 13943
rect 192 13909 204 13943
rect 48 13669 60 13703
rect 72 13669 84 13703
rect 96 13669 108 13703
rect 120 13669 132 13703
rect 144 13669 156 13703
rect 168 13669 180 13703
rect 192 13669 204 13703
rect 216 13669 228 13703
rect 48 13429 60 13463
rect 72 13429 84 13463
rect 96 13429 108 13463
rect 120 13429 132 13463
rect 144 13429 156 13463
rect 168 13429 180 13463
rect 192 13429 204 13463
rect 216 13429 228 13463
rect 240 13429 252 13463
rect 48 13189 60 13223
rect 72 13189 84 13223
rect 96 13189 108 13223
rect 120 13189 132 13223
rect 144 13189 156 13223
rect 168 13189 180 13223
rect 192 13189 204 13223
rect 216 13189 228 13223
rect 240 13189 252 13223
rect 264 13189 276 13223
rect 48 12949 60 12983
rect 72 12949 84 12983
rect 96 12949 108 12983
rect 120 12949 132 12983
rect 144 12949 156 12983
rect 168 12949 180 12983
rect 192 12949 204 12983
rect 216 12949 228 12983
rect 240 12949 252 12983
rect 264 12949 276 12983
rect 288 12949 300 12983
rect 48 12709 60 12743
rect 72 12709 84 12743
rect 96 12709 108 12743
rect 120 12709 132 12743
rect 144 12709 156 12743
rect 168 12709 180 12743
rect 192 12709 204 12743
rect 216 12709 228 12743
rect 240 12709 252 12743
rect 264 12709 276 12743
rect 288 12709 300 12743
rect 312 12709 324 12743
rect 48 12469 60 12503
rect 72 12469 84 12503
rect 96 12469 108 12503
rect 120 12469 132 12503
rect 144 12469 156 12503
rect 168 12469 180 12503
rect 192 12469 204 12503
rect 216 12469 228 12503
rect 240 12469 252 12503
rect 264 12469 276 12503
rect 288 12469 300 12503
rect 312 12469 324 12503
rect 336 12469 348 12503
rect 48 12229 60 12263
rect 72 12229 84 12263
rect 96 12229 108 12263
rect 120 12229 132 12263
rect 144 12229 156 12263
rect 168 12229 180 12263
rect 192 12229 204 12263
rect 216 12229 228 12263
rect 240 12229 252 12263
rect 264 12229 276 12263
rect 288 12229 300 12263
rect 312 12229 324 12263
rect 336 12229 348 12263
rect 360 12229 372 12263
rect 48 11989 60 12023
rect 72 11989 84 12023
rect 96 11989 108 12023
rect 120 11989 132 12023
rect 144 11989 156 12023
rect 168 11989 180 12023
rect 192 11989 204 12023
rect 216 11989 228 12023
rect 240 11989 252 12023
rect 264 11989 276 12023
rect 288 11989 300 12023
rect 312 11989 324 12023
rect 336 11989 348 12023
rect 360 11989 372 12023
rect 384 11989 396 12023
rect 48 11749 60 11783
rect 72 11749 84 11783
rect 96 11749 108 11783
rect 120 11749 132 11783
rect 144 11749 156 11783
rect 168 11749 180 11783
rect 192 11749 204 11783
rect 216 11749 228 11783
rect 240 11749 252 11783
rect 264 11749 276 11783
rect 288 11749 300 11783
rect 312 11749 324 11783
rect 336 11749 348 11783
rect 360 11749 372 11783
rect 384 11749 396 11783
rect 408 11749 420 11783
rect 48 11509 60 11543
rect 72 11509 84 11543
rect 96 11509 108 11543
rect 120 11509 132 11543
rect 144 11509 156 11543
rect 168 11509 180 11543
rect 192 11509 204 11543
rect 216 11509 228 11543
rect 240 11509 252 11543
rect 264 11509 276 11543
rect 288 11509 300 11543
rect 312 11509 324 11543
rect 336 11509 348 11543
rect 360 11509 372 11543
rect 384 11509 396 11543
rect 408 11509 420 11543
rect 432 11509 444 11543
rect 48 11269 60 11303
rect 72 11269 84 11303
rect 96 11269 108 11303
rect 120 11269 132 11303
rect 144 11269 156 11303
rect 168 11269 180 11303
rect 192 11269 204 11303
rect 216 11269 228 11303
rect 240 11269 252 11303
rect 264 11269 276 11303
rect 288 11269 300 11303
rect 312 11269 324 11303
rect 336 11269 348 11303
rect 360 11269 372 11303
rect 384 11269 396 11303
rect 408 11269 420 11303
rect 432 11269 444 11303
rect 456 11269 468 11303
rect 48 11029 60 11063
rect 72 11029 84 11063
rect 96 11029 108 11063
rect 120 11029 132 11063
rect 144 11029 156 11063
rect 168 11029 180 11063
rect 192 11029 204 11063
rect 216 11029 228 11063
rect 240 11029 252 11063
rect 264 11029 276 11063
rect 288 11029 300 11063
rect 312 11029 324 11063
rect 336 11029 348 11063
rect 360 11029 372 11063
rect 384 11029 396 11063
rect 408 11029 420 11063
rect 432 11029 444 11063
rect 456 11029 468 11063
rect 480 11029 492 11063
rect 48 10789 60 10823
rect 72 10789 84 10823
rect 96 10789 108 10823
rect 120 10789 132 10823
rect 144 10789 156 10823
rect 168 10789 180 10823
rect 192 10789 204 10823
rect 216 10789 228 10823
rect 240 10789 252 10823
rect 264 10789 276 10823
rect 288 10789 300 10823
rect 312 10789 324 10823
rect 336 10789 348 10823
rect 360 10789 372 10823
rect 384 10789 396 10823
rect 408 10789 420 10823
rect 432 10789 444 10823
rect 456 10789 468 10823
rect 480 10789 492 10823
rect 504 10789 516 10823
rect 48 10549 60 10583
rect 72 10549 84 10583
rect 96 10549 108 10583
rect 120 10549 132 10583
rect 144 10549 156 10583
rect 168 10549 180 10583
rect 192 10549 204 10583
rect 216 10549 228 10583
rect 240 10549 252 10583
rect 264 10549 276 10583
rect 288 10549 300 10583
rect 312 10549 324 10583
rect 336 10549 348 10583
rect 360 10549 372 10583
rect 384 10549 396 10583
rect 408 10549 420 10583
rect 432 10549 444 10583
rect 456 10549 468 10583
rect 480 10549 492 10583
rect 504 10549 516 10583
rect 528 10549 540 10583
rect 48 10309 60 10343
rect 72 10309 84 10343
rect 96 10309 108 10343
rect 120 10309 132 10343
rect 144 10309 156 10343
rect 168 10309 180 10343
rect 192 10309 204 10343
rect 216 10309 228 10343
rect 240 10309 252 10343
rect 264 10309 276 10343
rect 288 10309 300 10343
rect 312 10309 324 10343
rect 336 10309 348 10343
rect 360 10309 372 10343
rect 384 10309 396 10343
rect 408 10309 420 10343
rect 432 10309 444 10343
rect 456 10309 468 10343
rect 480 10309 492 10343
rect 504 10309 516 10343
rect 528 10309 540 10343
rect 552 10309 564 10343
rect 48 10069 60 10103
rect 72 10069 84 10103
rect 96 10069 108 10103
rect 120 10069 132 10103
rect 144 10069 156 10103
rect 168 10069 180 10103
rect 192 10069 204 10103
rect 216 10069 228 10103
rect 240 10069 252 10103
rect 264 10069 276 10103
rect 288 10069 300 10103
rect 312 10069 324 10103
rect 336 10069 348 10103
rect 360 10069 372 10103
rect 384 10069 396 10103
rect 408 10069 420 10103
rect 432 10069 444 10103
rect 456 10069 468 10103
rect 480 10069 492 10103
rect 504 10069 516 10103
rect 528 10069 540 10103
rect 552 10069 564 10103
rect 576 10069 588 10103
rect 48 9829 60 9863
rect 72 9829 84 9863
rect 96 9829 108 9863
rect 120 9829 132 9863
rect 144 9829 156 9863
rect 168 9829 180 9863
rect 192 9829 204 9863
rect 216 9829 228 9863
rect 240 9829 252 9863
rect 264 9829 276 9863
rect 288 9829 300 9863
rect 312 9829 324 9863
rect 336 9829 348 9863
rect 360 9829 372 9863
rect 384 9829 396 9863
rect 408 9829 420 9863
rect 432 9829 444 9863
rect 456 9829 468 9863
rect 480 9829 492 9863
rect 504 9829 516 9863
rect 528 9829 540 9863
rect 552 9829 564 9863
rect 576 9829 588 9863
rect 600 9829 612 9863
rect 48 9589 60 9623
rect 72 9589 84 9623
rect 96 9589 108 9623
rect 120 9589 132 9623
rect 144 9589 156 9623
rect 168 9589 180 9623
rect 192 9589 204 9623
rect 216 9589 228 9623
rect 240 9589 252 9623
rect 264 9589 276 9623
rect 288 9589 300 9623
rect 312 9589 324 9623
rect 336 9589 348 9623
rect 360 9589 372 9623
rect 384 9589 396 9623
rect 408 9589 420 9623
rect 432 9589 444 9623
rect 456 9589 468 9623
rect 480 9589 492 9623
rect 504 9589 516 9623
rect 528 9589 540 9623
rect 552 9589 564 9623
rect 576 9589 588 9623
rect 600 9589 612 9623
rect 624 9589 636 9623
rect 48 9349 60 9383
rect 72 9349 84 9383
rect 96 9349 108 9383
rect 120 9349 132 9383
rect 144 9349 156 9383
rect 168 9349 180 9383
rect 192 9349 204 9383
rect 216 9349 228 9383
rect 240 9349 252 9383
rect 264 9349 276 9383
rect 288 9349 300 9383
rect 312 9349 324 9383
rect 336 9349 348 9383
rect 360 9349 372 9383
rect 384 9349 396 9383
rect 408 9349 420 9383
rect 432 9349 444 9383
rect 456 9349 468 9383
rect 480 9349 492 9383
rect 504 9349 516 9383
rect 528 9349 540 9383
rect 552 9349 564 9383
rect 576 9349 588 9383
rect 600 9349 612 9383
rect 624 9349 636 9383
rect 648 9349 660 9383
rect 48 9109 60 9143
rect 72 9109 84 9143
rect 96 9109 108 9143
rect 120 9109 132 9143
rect 144 9109 156 9143
rect 168 9109 180 9143
rect 192 9109 204 9143
rect 216 9109 228 9143
rect 240 9109 252 9143
rect 264 9109 276 9143
rect 288 9109 300 9143
rect 312 9109 324 9143
rect 336 9109 348 9143
rect 360 9109 372 9143
rect 384 9109 396 9143
rect 408 9109 420 9143
rect 432 9109 444 9143
rect 456 9109 468 9143
rect 480 9109 492 9143
rect 504 9109 516 9143
rect 528 9109 540 9143
rect 552 9109 564 9143
rect 576 9109 588 9143
rect 600 9109 612 9143
rect 624 9109 636 9143
rect 648 9109 660 9143
rect 672 9109 684 9143
rect 48 8869 60 8903
rect 72 8869 84 8903
rect 96 8869 108 8903
rect 120 8869 132 8903
rect 144 8869 156 8903
rect 168 8869 180 8903
rect 192 8869 204 8903
rect 216 8869 228 8903
rect 240 8869 252 8903
rect 264 8869 276 8903
rect 288 8869 300 8903
rect 312 8869 324 8903
rect 336 8869 348 8903
rect 360 8869 372 8903
rect 384 8869 396 8903
rect 408 8869 420 8903
rect 432 8869 444 8903
rect 456 8869 468 8903
rect 480 8869 492 8903
rect 504 8869 516 8903
rect 528 8869 540 8903
rect 552 8869 564 8903
rect 576 8869 588 8903
rect 600 8869 612 8903
rect 624 8869 636 8903
rect 648 8869 660 8903
rect 672 8869 684 8903
rect 696 8869 708 8903
rect 48 8629 60 8663
rect 72 8629 84 8663
rect 96 8629 108 8663
rect 120 8629 132 8663
rect 144 8629 156 8663
rect 168 8629 180 8663
rect 192 8629 204 8663
rect 216 8629 228 8663
rect 240 8629 252 8663
rect 264 8629 276 8663
rect 288 8629 300 8663
rect 312 8629 324 8663
rect 336 8629 348 8663
rect 360 8629 372 8663
rect 384 8629 396 8663
rect 408 8629 420 8663
rect 432 8629 444 8663
rect 456 8629 468 8663
rect 480 8629 492 8663
rect 504 8629 516 8663
rect 528 8629 540 8663
rect 552 8629 564 8663
rect 576 8629 588 8663
rect 600 8629 612 8663
rect 624 8629 636 8663
rect 648 8629 660 8663
rect 672 8629 684 8663
rect 696 8629 708 8663
rect 720 8629 732 8663
rect 48 8389 60 8423
rect 72 8389 84 8423
rect 96 8389 108 8423
rect 120 8389 132 8423
rect 144 8389 156 8423
rect 168 8389 180 8423
rect 192 8389 204 8423
rect 216 8389 228 8423
rect 240 8389 252 8423
rect 264 8389 276 8423
rect 288 8389 300 8423
rect 312 8389 324 8423
rect 336 8389 348 8423
rect 360 8389 372 8423
rect 384 8389 396 8423
rect 408 8389 420 8423
rect 432 8389 444 8423
rect 456 8389 468 8423
rect 480 8389 492 8423
rect 504 8389 516 8423
rect 528 8389 540 8423
rect 552 8389 564 8423
rect 576 8389 588 8423
rect 600 8389 612 8423
rect 624 8389 636 8423
rect 648 8389 660 8423
rect 672 8389 684 8423
rect 696 8389 708 8423
rect 720 8389 732 8423
rect 744 8389 756 8423
rect 48 8149 60 8183
rect 72 8149 84 8183
rect 96 8149 108 8183
rect 120 8149 132 8183
rect 144 8149 156 8183
rect 168 8149 180 8183
rect 192 8149 204 8183
rect 216 8149 228 8183
rect 240 8149 252 8183
rect 264 8149 276 8183
rect 288 8149 300 8183
rect 312 8149 324 8183
rect 336 8149 348 8183
rect 360 8149 372 8183
rect 384 8149 396 8183
rect 408 8149 420 8183
rect 432 8149 444 8183
rect 456 8149 468 8183
rect 480 8149 492 8183
rect 504 8149 516 8183
rect 528 8149 540 8183
rect 552 8149 564 8183
rect 576 8149 588 8183
rect 600 8149 612 8183
rect 624 8149 636 8183
rect 648 8149 660 8183
rect 672 8149 684 8183
rect 696 8149 708 8183
rect 720 8149 732 8183
rect 744 8149 756 8183
rect 768 8149 780 8183
rect 48 7909 60 7943
rect 72 7909 84 7943
rect 96 7909 108 7943
rect 120 7909 132 7943
rect 144 7909 156 7943
rect 168 7909 180 7943
rect 192 7909 204 7943
rect 216 7909 228 7943
rect 240 7909 252 7943
rect 264 7909 276 7943
rect 288 7909 300 7943
rect 312 7909 324 7943
rect 336 7909 348 7943
rect 360 7909 372 7943
rect 384 7909 396 7943
rect 408 7909 420 7943
rect 432 7909 444 7943
rect 456 7909 468 7943
rect 480 7909 492 7943
rect 504 7909 516 7943
rect 528 7909 540 7943
rect 552 7909 564 7943
rect 576 7909 588 7943
rect 600 7909 612 7943
rect 624 7909 636 7943
rect 648 7909 660 7943
rect 672 7909 684 7943
rect 696 7909 708 7943
rect 720 7909 732 7943
rect 744 7909 756 7943
rect 768 7909 780 7943
rect 792 7909 804 7943
rect 48 7669 60 7703
rect 72 7669 84 7703
rect 96 7669 108 7703
rect 120 7669 132 7703
rect 144 7669 156 7703
rect 168 7669 180 7703
rect 192 7669 204 7703
rect 216 7669 228 7703
rect 240 7669 252 7703
rect 264 7669 276 7703
rect 288 7669 300 7703
rect 312 7669 324 7703
rect 336 7669 348 7703
rect 360 7669 372 7703
rect 384 7669 396 7703
rect 408 7669 420 7703
rect 432 7669 444 7703
rect 456 7669 468 7703
rect 480 7669 492 7703
rect 504 7669 516 7703
rect 528 7669 540 7703
rect 552 7669 564 7703
rect 576 7669 588 7703
rect 600 7669 612 7703
rect 624 7669 636 7703
rect 648 7669 660 7703
rect 672 7669 684 7703
rect 696 7669 708 7703
rect 720 7669 732 7703
rect 744 7669 756 7703
rect 768 7669 780 7703
rect 792 7669 804 7703
rect 816 7669 828 7703
rect 48 7429 60 7463
rect 72 7429 84 7463
rect 96 7429 108 7463
rect 120 7429 132 7463
rect 144 7429 156 7463
rect 168 7429 180 7463
rect 192 7429 204 7463
rect 216 7429 228 7463
rect 240 7429 252 7463
rect 264 7429 276 7463
rect 288 7429 300 7463
rect 312 7429 324 7463
rect 336 7429 348 7463
rect 360 7429 372 7463
rect 384 7429 396 7463
rect 408 7429 420 7463
rect 432 7429 444 7463
rect 456 7429 468 7463
rect 480 7429 492 7463
rect 504 7429 516 7463
rect 528 7429 540 7463
rect 552 7429 564 7463
rect 576 7429 588 7463
rect 600 7429 612 7463
rect 624 7429 636 7463
rect 648 7429 660 7463
rect 672 7429 684 7463
rect 696 7429 708 7463
rect 720 7429 732 7463
rect 744 7429 756 7463
rect 768 7429 780 7463
rect 792 7429 804 7463
rect 816 7429 828 7463
rect 840 7429 852 7463
rect 48 7189 60 7223
rect 72 7189 84 7223
rect 96 7189 108 7223
rect 120 7189 132 7223
rect 144 7189 156 7223
rect 168 7189 180 7223
rect 192 7189 204 7223
rect 216 7189 228 7223
rect 240 7189 252 7223
rect 264 7189 276 7223
rect 288 7189 300 7223
rect 312 7189 324 7223
rect 336 7189 348 7223
rect 360 7189 372 7223
rect 384 7189 396 7223
rect 408 7189 420 7223
rect 432 7189 444 7223
rect 456 7189 468 7223
rect 480 7189 492 7223
rect 504 7189 516 7223
rect 528 7189 540 7223
rect 552 7189 564 7223
rect 576 7189 588 7223
rect 600 7189 612 7223
rect 624 7189 636 7223
rect 648 7189 660 7223
rect 672 7189 684 7223
rect 696 7189 708 7223
rect 720 7189 732 7223
rect 744 7189 756 7223
rect 768 7189 780 7223
rect 792 7189 804 7223
rect 816 7189 828 7223
rect 840 7189 852 7223
rect 864 7189 876 7223
rect 48 6949 60 6983
rect 72 6949 84 6983
rect 96 6949 108 6983
rect 120 6949 132 6983
rect 144 6949 156 6983
rect 168 6949 180 6983
rect 192 6949 204 6983
rect 216 6949 228 6983
rect 240 6949 252 6983
rect 264 6949 276 6983
rect 288 6949 300 6983
rect 312 6949 324 6983
rect 336 6949 348 6983
rect 360 6949 372 6983
rect 384 6949 396 6983
rect 408 6949 420 6983
rect 432 6949 444 6983
rect 456 6949 468 6983
rect 480 6949 492 6983
rect 504 6949 516 6983
rect 528 6949 540 6983
rect 552 6949 564 6983
rect 576 6949 588 6983
rect 600 6949 612 6983
rect 624 6949 636 6983
rect 648 6949 660 6983
rect 672 6949 684 6983
rect 696 6949 708 6983
rect 720 6949 732 6983
rect 744 6949 756 6983
rect 768 6949 780 6983
rect 792 6949 804 6983
rect 816 6949 828 6983
rect 840 6949 852 6983
rect 864 6949 876 6983
rect 888 6949 900 6983
rect 48 6709 60 6743
rect 72 6709 84 6743
rect 96 6709 108 6743
rect 120 6709 132 6743
rect 144 6709 156 6743
rect 168 6709 180 6743
rect 192 6709 204 6743
rect 216 6709 228 6743
rect 240 6709 252 6743
rect 264 6709 276 6743
rect 288 6709 300 6743
rect 312 6709 324 6743
rect 336 6709 348 6743
rect 360 6709 372 6743
rect 384 6709 396 6743
rect 408 6709 420 6743
rect 432 6709 444 6743
rect 456 6709 468 6743
rect 480 6709 492 6743
rect 504 6709 516 6743
rect 528 6709 540 6743
rect 552 6709 564 6743
rect 576 6709 588 6743
rect 600 6709 612 6743
rect 624 6709 636 6743
rect 648 6709 660 6743
rect 672 6709 684 6743
rect 696 6709 708 6743
rect 720 6709 732 6743
rect 744 6709 756 6743
rect 768 6709 780 6743
rect 792 6709 804 6743
rect 816 6709 828 6743
rect 840 6709 852 6743
rect 864 6709 876 6743
rect 888 6709 900 6743
rect 912 6709 924 6743
rect 48 6469 60 6503
rect 72 6469 84 6503
rect 96 6469 108 6503
rect 120 6469 132 6503
rect 144 6469 156 6503
rect 168 6469 180 6503
rect 192 6469 204 6503
rect 216 6469 228 6503
rect 240 6469 252 6503
rect 264 6469 276 6503
rect 288 6469 300 6503
rect 312 6469 324 6503
rect 336 6469 348 6503
rect 360 6469 372 6503
rect 384 6469 396 6503
rect 408 6469 420 6503
rect 432 6469 444 6503
rect 456 6469 468 6503
rect 480 6469 492 6503
rect 504 6469 516 6503
rect 528 6469 540 6503
rect 552 6469 564 6503
rect 576 6469 588 6503
rect 600 6469 612 6503
rect 624 6469 636 6503
rect 648 6469 660 6503
rect 672 6469 684 6503
rect 696 6469 708 6503
rect 720 6469 732 6503
rect 744 6469 756 6503
rect 768 6469 780 6503
rect 792 6469 804 6503
rect 816 6469 828 6503
rect 840 6469 852 6503
rect 864 6469 876 6503
rect 888 6469 900 6503
rect 912 6469 924 6503
rect 936 6469 948 6503
rect 48 6229 60 6263
rect 72 6229 84 6263
rect 96 6229 108 6263
rect 120 6229 132 6263
rect 144 6229 156 6263
rect 168 6229 180 6263
rect 192 6229 204 6263
rect 216 6229 228 6263
rect 240 6229 252 6263
rect 264 6229 276 6263
rect 288 6229 300 6263
rect 312 6229 324 6263
rect 336 6229 348 6263
rect 360 6229 372 6263
rect 384 6229 396 6263
rect 408 6229 420 6263
rect 432 6229 444 6263
rect 456 6229 468 6263
rect 480 6229 492 6263
rect 504 6229 516 6263
rect 528 6229 540 6263
rect 552 6229 564 6263
rect 576 6229 588 6263
rect 600 6229 612 6263
rect 624 6229 636 6263
rect 648 6229 660 6263
rect 672 6229 684 6263
rect 696 6229 708 6263
rect 720 6229 732 6263
rect 744 6229 756 6263
rect 768 6229 780 6263
rect 792 6229 804 6263
rect 816 6229 828 6263
rect 840 6229 852 6263
rect 864 6229 876 6263
rect 888 6229 900 6263
rect 912 6229 924 6263
rect 936 6229 948 6263
rect 960 6229 972 6263
rect 48 5989 60 6023
rect 72 5989 84 6023
rect 96 5989 108 6023
rect 120 5989 132 6023
rect 144 5989 156 6023
rect 168 5989 180 6023
rect 192 5989 204 6023
rect 216 5989 228 6023
rect 240 5989 252 6023
rect 264 5989 276 6023
rect 288 5989 300 6023
rect 312 5989 324 6023
rect 336 5989 348 6023
rect 360 5989 372 6023
rect 384 5989 396 6023
rect 408 5989 420 6023
rect 432 5989 444 6023
rect 456 5989 468 6023
rect 480 5989 492 6023
rect 504 5989 516 6023
rect 528 5989 540 6023
rect 552 5989 564 6023
rect 576 5989 588 6023
rect 600 5989 612 6023
rect 624 5989 636 6023
rect 648 5989 660 6023
rect 672 5989 684 6023
rect 696 5989 708 6023
rect 720 5989 732 6023
rect 744 5989 756 6023
rect 768 5989 780 6023
rect 792 5989 804 6023
rect 816 5989 828 6023
rect 840 5989 852 6023
rect 864 5989 876 6023
rect 888 5989 900 6023
rect 912 5989 924 6023
rect 936 5989 948 6023
rect 960 5989 972 6023
rect 984 5989 996 6023
rect 48 5749 60 5783
rect 72 5749 84 5783
rect 96 5749 108 5783
rect 120 5749 132 5783
rect 144 5749 156 5783
rect 168 5749 180 5783
rect 192 5749 204 5783
rect 216 5749 228 5783
rect 240 5749 252 5783
rect 264 5749 276 5783
rect 288 5749 300 5783
rect 312 5749 324 5783
rect 336 5749 348 5783
rect 360 5749 372 5783
rect 384 5749 396 5783
rect 408 5749 420 5783
rect 432 5749 444 5783
rect 456 5749 468 5783
rect 480 5749 492 5783
rect 504 5749 516 5783
rect 528 5749 540 5783
rect 552 5749 564 5783
rect 576 5749 588 5783
rect 600 5749 612 5783
rect 624 5749 636 5783
rect 648 5749 660 5783
rect 672 5749 684 5783
rect 696 5749 708 5783
rect 720 5749 732 5783
rect 744 5749 756 5783
rect 768 5749 780 5783
rect 792 5749 804 5783
rect 816 5749 828 5783
rect 840 5749 852 5783
rect 864 5749 876 5783
rect 888 5749 900 5783
rect 912 5749 924 5783
rect 936 5749 948 5783
rect 960 5749 972 5783
rect 984 5749 996 5783
rect 1008 5749 1020 5783
rect 48 5509 60 5543
rect 72 5509 84 5543
rect 96 5509 108 5543
rect 120 5509 132 5543
rect 144 5509 156 5543
rect 168 5509 180 5543
rect 192 5509 204 5543
rect 216 5509 228 5543
rect 240 5509 252 5543
rect 264 5509 276 5543
rect 288 5509 300 5543
rect 312 5509 324 5543
rect 336 5509 348 5543
rect 360 5509 372 5543
rect 384 5509 396 5543
rect 408 5509 420 5543
rect 432 5509 444 5543
rect 456 5509 468 5543
rect 480 5509 492 5543
rect 504 5509 516 5543
rect 528 5509 540 5543
rect 552 5509 564 5543
rect 576 5509 588 5543
rect 600 5509 612 5543
rect 624 5509 636 5543
rect 648 5509 660 5543
rect 672 5509 684 5543
rect 696 5509 708 5543
rect 720 5509 732 5543
rect 744 5509 756 5543
rect 768 5509 780 5543
rect 792 5509 804 5543
rect 816 5509 828 5543
rect 840 5509 852 5543
rect 864 5509 876 5543
rect 888 5509 900 5543
rect 912 5509 924 5543
rect 936 5509 948 5543
rect 960 5509 972 5543
rect 984 5509 996 5543
rect 1008 5509 1020 5543
rect 1032 5509 1044 5543
rect 48 5269 60 5303
rect 72 5269 84 5303
rect 96 5269 108 5303
rect 120 5269 132 5303
rect 144 5269 156 5303
rect 168 5269 180 5303
rect 192 5269 204 5303
rect 216 5269 228 5303
rect 240 5269 252 5303
rect 264 5269 276 5303
rect 288 5269 300 5303
rect 312 5269 324 5303
rect 336 5269 348 5303
rect 360 5269 372 5303
rect 384 5269 396 5303
rect 408 5269 420 5303
rect 432 5269 444 5303
rect 456 5269 468 5303
rect 480 5269 492 5303
rect 504 5269 516 5303
rect 528 5269 540 5303
rect 552 5269 564 5303
rect 576 5269 588 5303
rect 600 5269 612 5303
rect 624 5269 636 5303
rect 648 5269 660 5303
rect 672 5269 684 5303
rect 696 5269 708 5303
rect 720 5269 732 5303
rect 744 5269 756 5303
rect 768 5269 780 5303
rect 792 5269 804 5303
rect 816 5269 828 5303
rect 840 5269 852 5303
rect 864 5269 876 5303
rect 888 5269 900 5303
rect 912 5269 924 5303
rect 936 5269 948 5303
rect 960 5269 972 5303
rect 984 5269 996 5303
rect 1008 5269 1020 5303
rect 1032 5269 1044 5303
rect 1056 5269 1068 5303
rect 48 5029 60 5063
rect 72 5029 84 5063
rect 96 5029 108 5063
rect 120 5029 132 5063
rect 144 5029 156 5063
rect 168 5029 180 5063
rect 192 5029 204 5063
rect 216 5029 228 5063
rect 240 5029 252 5063
rect 264 5029 276 5063
rect 288 5029 300 5063
rect 312 5029 324 5063
rect 336 5029 348 5063
rect 360 5029 372 5063
rect 384 5029 396 5063
rect 408 5029 420 5063
rect 432 5029 444 5063
rect 456 5029 468 5063
rect 480 5029 492 5063
rect 504 5029 516 5063
rect 528 5029 540 5063
rect 552 5029 564 5063
rect 576 5029 588 5063
rect 600 5029 612 5063
rect 624 5029 636 5063
rect 648 5029 660 5063
rect 672 5029 684 5063
rect 696 5029 708 5063
rect 720 5029 732 5063
rect 744 5029 756 5063
rect 768 5029 780 5063
rect 792 5029 804 5063
rect 816 5029 828 5063
rect 840 5029 852 5063
rect 864 5029 876 5063
rect 888 5029 900 5063
rect 912 5029 924 5063
rect 936 5029 948 5063
rect 960 5029 972 5063
rect 984 5029 996 5063
rect 1008 5029 1020 5063
rect 1032 5029 1044 5063
rect 1056 5029 1068 5063
rect 1080 5029 1092 5063
rect 48 4789 60 4823
rect 72 4789 84 4823
rect 96 4789 108 4823
rect 120 4789 132 4823
rect 144 4789 156 4823
rect 168 4789 180 4823
rect 192 4789 204 4823
rect 216 4789 228 4823
rect 240 4789 252 4823
rect 264 4789 276 4823
rect 288 4789 300 4823
rect 312 4789 324 4823
rect 336 4789 348 4823
rect 360 4789 372 4823
rect 384 4789 396 4823
rect 408 4789 420 4823
rect 432 4789 444 4823
rect 456 4789 468 4823
rect 480 4789 492 4823
rect 504 4789 516 4823
rect 528 4789 540 4823
rect 552 4789 564 4823
rect 576 4789 588 4823
rect 600 4789 612 4823
rect 624 4789 636 4823
rect 648 4789 660 4823
rect 672 4789 684 4823
rect 696 4789 708 4823
rect 720 4789 732 4823
rect 744 4789 756 4823
rect 768 4789 780 4823
rect 792 4789 804 4823
rect 816 4789 828 4823
rect 840 4789 852 4823
rect 864 4789 876 4823
rect 888 4789 900 4823
rect 912 4789 924 4823
rect 936 4789 948 4823
rect 960 4789 972 4823
rect 984 4789 996 4823
rect 1008 4789 1020 4823
rect 1032 4789 1044 4823
rect 1056 4789 1068 4823
rect 1080 4789 1092 4823
rect 1104 4789 1116 4823
rect 48 4549 60 4583
rect 72 4549 84 4583
rect 96 4549 108 4583
rect 120 4549 132 4583
rect 144 4549 156 4583
rect 168 4549 180 4583
rect 192 4549 204 4583
rect 216 4549 228 4583
rect 240 4549 252 4583
rect 264 4549 276 4583
rect 288 4549 300 4583
rect 312 4549 324 4583
rect 336 4549 348 4583
rect 360 4549 372 4583
rect 384 4549 396 4583
rect 408 4549 420 4583
rect 432 4549 444 4583
rect 456 4549 468 4583
rect 480 4549 492 4583
rect 504 4549 516 4583
rect 528 4549 540 4583
rect 552 4549 564 4583
rect 576 4549 588 4583
rect 600 4549 612 4583
rect 624 4549 636 4583
rect 648 4549 660 4583
rect 672 4549 684 4583
rect 696 4549 708 4583
rect 720 4549 732 4583
rect 744 4549 756 4583
rect 768 4549 780 4583
rect 792 4549 804 4583
rect 816 4549 828 4583
rect 840 4549 852 4583
rect 864 4549 876 4583
rect 888 4549 900 4583
rect 912 4549 924 4583
rect 936 4549 948 4583
rect 960 4549 972 4583
rect 984 4549 996 4583
rect 1008 4549 1020 4583
rect 1032 4549 1044 4583
rect 1056 4549 1068 4583
rect 1080 4549 1092 4583
rect 1104 4549 1116 4583
rect 1128 4549 1140 4583
rect 48 4309 60 4343
rect 72 4309 84 4343
rect 96 4309 108 4343
rect 120 4309 132 4343
rect 144 4309 156 4343
rect 168 4309 180 4343
rect 192 4309 204 4343
rect 216 4309 228 4343
rect 240 4309 252 4343
rect 264 4309 276 4343
rect 288 4309 300 4343
rect 312 4309 324 4343
rect 336 4309 348 4343
rect 360 4309 372 4343
rect 384 4309 396 4343
rect 408 4309 420 4343
rect 432 4309 444 4343
rect 456 4309 468 4343
rect 480 4309 492 4343
rect 504 4309 516 4343
rect 528 4309 540 4343
rect 552 4309 564 4343
rect 576 4309 588 4343
rect 600 4309 612 4343
rect 624 4309 636 4343
rect 648 4309 660 4343
rect 672 4309 684 4343
rect 696 4309 708 4343
rect 720 4309 732 4343
rect 744 4309 756 4343
rect 768 4309 780 4343
rect 792 4309 804 4343
rect 816 4309 828 4343
rect 840 4309 852 4343
rect 864 4309 876 4343
rect 888 4309 900 4343
rect 912 4309 924 4343
rect 936 4309 948 4343
rect 960 4309 972 4343
rect 984 4309 996 4343
rect 1008 4309 1020 4343
rect 1032 4309 1044 4343
rect 1056 4309 1068 4343
rect 1080 4309 1092 4343
rect 1104 4309 1116 4343
rect 1128 4309 1140 4343
rect 1152 4309 1164 4343
rect 48 4069 60 4103
rect 72 4069 84 4103
rect 96 4069 108 4103
rect 120 4069 132 4103
rect 144 4069 156 4103
rect 168 4069 180 4103
rect 192 4069 204 4103
rect 216 4069 228 4103
rect 240 4069 252 4103
rect 264 4069 276 4103
rect 288 4069 300 4103
rect 312 4069 324 4103
rect 336 4069 348 4103
rect 360 4069 372 4103
rect 384 4069 396 4103
rect 408 4069 420 4103
rect 432 4069 444 4103
rect 456 4069 468 4103
rect 480 4069 492 4103
rect 504 4069 516 4103
rect 528 4069 540 4103
rect 552 4069 564 4103
rect 576 4069 588 4103
rect 600 4069 612 4103
rect 624 4069 636 4103
rect 648 4069 660 4103
rect 672 4069 684 4103
rect 696 4069 708 4103
rect 720 4069 732 4103
rect 744 4069 756 4103
rect 768 4069 780 4103
rect 792 4069 804 4103
rect 816 4069 828 4103
rect 840 4069 852 4103
rect 864 4069 876 4103
rect 888 4069 900 4103
rect 912 4069 924 4103
rect 936 4069 948 4103
rect 960 4069 972 4103
rect 984 4069 996 4103
rect 1008 4069 1020 4103
rect 1032 4069 1044 4103
rect 1056 4069 1068 4103
rect 1080 4069 1092 4103
rect 1104 4069 1116 4103
rect 1128 4069 1140 4103
rect 1152 4069 1164 4103
rect 1176 4069 1188 4103
rect 48 3829 60 3863
rect 72 3829 84 3863
rect 96 3829 108 3863
rect 120 3829 132 3863
rect 144 3829 156 3863
rect 168 3829 180 3863
rect 192 3829 204 3863
rect 216 3829 228 3863
rect 240 3829 252 3863
rect 264 3829 276 3863
rect 288 3829 300 3863
rect 312 3829 324 3863
rect 336 3829 348 3863
rect 360 3829 372 3863
rect 384 3829 396 3863
rect 408 3829 420 3863
rect 432 3829 444 3863
rect 456 3829 468 3863
rect 480 3829 492 3863
rect 504 3829 516 3863
rect 528 3829 540 3863
rect 552 3829 564 3863
rect 576 3829 588 3863
rect 600 3829 612 3863
rect 624 3829 636 3863
rect 648 3829 660 3863
rect 672 3829 684 3863
rect 696 3829 708 3863
rect 720 3829 732 3863
rect 744 3829 756 3863
rect 768 3829 780 3863
rect 792 3829 804 3863
rect 816 3829 828 3863
rect 840 3829 852 3863
rect 864 3829 876 3863
rect 888 3829 900 3863
rect 912 3829 924 3863
rect 936 3829 948 3863
rect 960 3829 972 3863
rect 984 3829 996 3863
rect 1008 3829 1020 3863
rect 1032 3829 1044 3863
rect 1056 3829 1068 3863
rect 1080 3829 1092 3863
rect 1104 3829 1116 3863
rect 1128 3829 1140 3863
rect 1152 3829 1164 3863
rect 1176 3829 1188 3863
rect 1200 3829 1212 3863
rect 48 3589 60 3623
rect 72 3589 84 3623
rect 96 3589 108 3623
rect 120 3589 132 3623
rect 144 3589 156 3623
rect 168 3589 180 3623
rect 192 3589 204 3623
rect 216 3589 228 3623
rect 240 3589 252 3623
rect 264 3589 276 3623
rect 288 3589 300 3623
rect 312 3589 324 3623
rect 336 3589 348 3623
rect 360 3589 372 3623
rect 384 3589 396 3623
rect 408 3589 420 3623
rect 432 3589 444 3623
rect 456 3589 468 3623
rect 480 3589 492 3623
rect 504 3589 516 3623
rect 528 3589 540 3623
rect 552 3589 564 3623
rect 576 3589 588 3623
rect 600 3589 612 3623
rect 624 3589 636 3623
rect 648 3589 660 3623
rect 672 3589 684 3623
rect 696 3589 708 3623
rect 720 3589 732 3623
rect 744 3589 756 3623
rect 768 3589 780 3623
rect 792 3589 804 3623
rect 816 3589 828 3623
rect 840 3589 852 3623
rect 864 3589 876 3623
rect 888 3589 900 3623
rect 912 3589 924 3623
rect 936 3589 948 3623
rect 960 3589 972 3623
rect 984 3589 996 3623
rect 1008 3589 1020 3623
rect 1032 3589 1044 3623
rect 1056 3589 1068 3623
rect 1080 3589 1092 3623
rect 1104 3589 1116 3623
rect 1128 3589 1140 3623
rect 1152 3589 1164 3623
rect 1176 3589 1188 3623
rect 1200 3589 1212 3623
rect 1224 3589 1236 3623
rect 48 3349 60 3383
rect 72 3349 84 3383
rect 96 3349 108 3383
rect 120 3349 132 3383
rect 144 3349 156 3383
rect 168 3349 180 3383
rect 192 3349 204 3383
rect 216 3349 228 3383
rect 240 3349 252 3383
rect 264 3349 276 3383
rect 288 3349 300 3383
rect 312 3349 324 3383
rect 336 3349 348 3383
rect 360 3349 372 3383
rect 384 3349 396 3383
rect 408 3349 420 3383
rect 432 3349 444 3383
rect 456 3349 468 3383
rect 480 3349 492 3383
rect 504 3349 516 3383
rect 528 3349 540 3383
rect 552 3349 564 3383
rect 576 3349 588 3383
rect 600 3349 612 3383
rect 624 3349 636 3383
rect 648 3349 660 3383
rect 672 3349 684 3383
rect 696 3349 708 3383
rect 720 3349 732 3383
rect 744 3349 756 3383
rect 768 3349 780 3383
rect 792 3349 804 3383
rect 816 3349 828 3383
rect 840 3349 852 3383
rect 864 3349 876 3383
rect 888 3349 900 3383
rect 912 3349 924 3383
rect 936 3349 948 3383
rect 960 3349 972 3383
rect 984 3349 996 3383
rect 1008 3349 1020 3383
rect 1032 3349 1044 3383
rect 1056 3349 1068 3383
rect 1080 3349 1092 3383
rect 1104 3349 1116 3383
rect 1128 3349 1140 3383
rect 1152 3349 1164 3383
rect 1176 3349 1188 3383
rect 1200 3349 1212 3383
rect 1224 3349 1236 3383
rect 1248 3349 1260 3383
rect 48 3109 60 3143
rect 72 3109 84 3143
rect 96 3109 108 3143
rect 120 3109 132 3143
rect 144 3109 156 3143
rect 168 3109 180 3143
rect 192 3109 204 3143
rect 216 3109 228 3143
rect 240 3109 252 3143
rect 264 3109 276 3143
rect 288 3109 300 3143
rect 312 3109 324 3143
rect 336 3109 348 3143
rect 360 3109 372 3143
rect 384 3109 396 3143
rect 408 3109 420 3143
rect 432 3109 444 3143
rect 456 3109 468 3143
rect 480 3109 492 3143
rect 504 3109 516 3143
rect 528 3109 540 3143
rect 552 3109 564 3143
rect 576 3109 588 3143
rect 600 3109 612 3143
rect 624 3109 636 3143
rect 648 3109 660 3143
rect 672 3109 684 3143
rect 696 3109 708 3143
rect 720 3109 732 3143
rect 744 3109 756 3143
rect 768 3109 780 3143
rect 792 3109 804 3143
rect 816 3109 828 3143
rect 840 3109 852 3143
rect 864 3109 876 3143
rect 888 3109 900 3143
rect 912 3109 924 3143
rect 936 3109 948 3143
rect 960 3109 972 3143
rect 984 3109 996 3143
rect 1008 3109 1020 3143
rect 1032 3109 1044 3143
rect 1056 3109 1068 3143
rect 1080 3109 1092 3143
rect 1104 3109 1116 3143
rect 1128 3109 1140 3143
rect 1152 3109 1164 3143
rect 1176 3109 1188 3143
rect 1200 3109 1212 3143
rect 1224 3109 1236 3143
rect 1248 3109 1260 3143
rect 1272 3109 1284 3143
rect 48 2869 60 2903
rect 72 2869 84 2903
rect 96 2869 108 2903
rect 120 2869 132 2903
rect 144 2869 156 2903
rect 168 2869 180 2903
rect 192 2869 204 2903
rect 216 2869 228 2903
rect 240 2869 252 2903
rect 264 2869 276 2903
rect 288 2869 300 2903
rect 312 2869 324 2903
rect 336 2869 348 2903
rect 360 2869 372 2903
rect 384 2869 396 2903
rect 408 2869 420 2903
rect 432 2869 444 2903
rect 456 2869 468 2903
rect 480 2869 492 2903
rect 504 2869 516 2903
rect 528 2869 540 2903
rect 552 2869 564 2903
rect 576 2869 588 2903
rect 600 2869 612 2903
rect 624 2869 636 2903
rect 648 2869 660 2903
rect 672 2869 684 2903
rect 696 2869 708 2903
rect 720 2869 732 2903
rect 744 2869 756 2903
rect 768 2869 780 2903
rect 792 2869 804 2903
rect 816 2869 828 2903
rect 840 2869 852 2903
rect 864 2869 876 2903
rect 888 2869 900 2903
rect 912 2869 924 2903
rect 936 2869 948 2903
rect 960 2869 972 2903
rect 984 2869 996 2903
rect 1008 2869 1020 2903
rect 1032 2869 1044 2903
rect 1056 2869 1068 2903
rect 1080 2869 1092 2903
rect 1104 2869 1116 2903
rect 1128 2869 1140 2903
rect 1152 2869 1164 2903
rect 1176 2869 1188 2903
rect 1200 2869 1212 2903
rect 1224 2869 1236 2903
rect 1248 2869 1260 2903
rect 1272 2869 1284 2903
rect 1296 2869 1308 2903
rect 48 2629 60 2663
rect 72 2629 84 2663
rect 96 2629 108 2663
rect 120 2629 132 2663
rect 144 2629 156 2663
rect 168 2629 180 2663
rect 192 2629 204 2663
rect 216 2629 228 2663
rect 240 2629 252 2663
rect 264 2629 276 2663
rect 288 2629 300 2663
rect 312 2629 324 2663
rect 336 2629 348 2663
rect 360 2629 372 2663
rect 384 2629 396 2663
rect 408 2629 420 2663
rect 432 2629 444 2663
rect 456 2629 468 2663
rect 480 2629 492 2663
rect 504 2629 516 2663
rect 528 2629 540 2663
rect 552 2629 564 2663
rect 576 2629 588 2663
rect 600 2629 612 2663
rect 624 2629 636 2663
rect 648 2629 660 2663
rect 672 2629 684 2663
rect 696 2629 708 2663
rect 720 2629 732 2663
rect 744 2629 756 2663
rect 768 2629 780 2663
rect 792 2629 804 2663
rect 816 2629 828 2663
rect 840 2629 852 2663
rect 864 2629 876 2663
rect 888 2629 900 2663
rect 912 2629 924 2663
rect 936 2629 948 2663
rect 960 2629 972 2663
rect 984 2629 996 2663
rect 1008 2629 1020 2663
rect 1032 2629 1044 2663
rect 1056 2629 1068 2663
rect 1080 2629 1092 2663
rect 1104 2629 1116 2663
rect 1128 2629 1140 2663
rect 1152 2629 1164 2663
rect 1176 2629 1188 2663
rect 1200 2629 1212 2663
rect 1224 2629 1236 2663
rect 1248 2629 1260 2663
rect 1272 2629 1284 2663
rect 1296 2629 1308 2663
rect 1320 2629 1332 2663
rect 48 2389 60 2423
rect 72 2389 84 2423
rect 96 2389 108 2423
rect 120 2389 132 2423
rect 144 2389 156 2423
rect 168 2389 180 2423
rect 192 2389 204 2423
rect 216 2389 228 2423
rect 240 2389 252 2423
rect 264 2389 276 2423
rect 288 2389 300 2423
rect 312 2389 324 2423
rect 336 2389 348 2423
rect 360 2389 372 2423
rect 384 2389 396 2423
rect 408 2389 420 2423
rect 432 2389 444 2423
rect 456 2389 468 2423
rect 480 2389 492 2423
rect 504 2389 516 2423
rect 528 2389 540 2423
rect 552 2389 564 2423
rect 576 2389 588 2423
rect 600 2389 612 2423
rect 624 2389 636 2423
rect 648 2389 660 2423
rect 672 2389 684 2423
rect 696 2389 708 2423
rect 720 2389 732 2423
rect 744 2389 756 2423
rect 768 2389 780 2423
rect 792 2389 804 2423
rect 816 2389 828 2423
rect 840 2389 852 2423
rect 864 2389 876 2423
rect 888 2389 900 2423
rect 912 2389 924 2423
rect 936 2389 948 2423
rect 960 2389 972 2423
rect 984 2389 996 2423
rect 1008 2389 1020 2423
rect 1032 2389 1044 2423
rect 1056 2389 1068 2423
rect 1080 2389 1092 2423
rect 1104 2389 1116 2423
rect 1128 2389 1140 2423
rect 1152 2389 1164 2423
rect 1176 2389 1188 2423
rect 1200 2389 1212 2423
rect 1224 2389 1236 2423
rect 1248 2389 1260 2423
rect 1272 2389 1284 2423
rect 1296 2389 1308 2423
rect 1320 2389 1332 2423
rect 1344 2389 1356 2423
rect 48 2149 60 2183
rect 72 2149 84 2183
rect 96 2149 108 2183
rect 120 2149 132 2183
rect 144 2149 156 2183
rect 168 2149 180 2183
rect 192 2149 204 2183
rect 216 2149 228 2183
rect 240 2149 252 2183
rect 264 2149 276 2183
rect 288 2149 300 2183
rect 312 2149 324 2183
rect 336 2149 348 2183
rect 360 2149 372 2183
rect 384 2149 396 2183
rect 408 2149 420 2183
rect 432 2149 444 2183
rect 456 2149 468 2183
rect 480 2149 492 2183
rect 504 2149 516 2183
rect 528 2149 540 2183
rect 552 2149 564 2183
rect 576 2149 588 2183
rect 600 2149 612 2183
rect 624 2149 636 2183
rect 648 2149 660 2183
rect 672 2149 684 2183
rect 696 2149 708 2183
rect 720 2149 732 2183
rect 744 2149 756 2183
rect 768 2149 780 2183
rect 792 2149 804 2183
rect 816 2149 828 2183
rect 840 2149 852 2183
rect 864 2149 876 2183
rect 888 2149 900 2183
rect 912 2149 924 2183
rect 936 2149 948 2183
rect 960 2149 972 2183
rect 984 2149 996 2183
rect 1008 2149 1020 2183
rect 1032 2149 1044 2183
rect 1056 2149 1068 2183
rect 1080 2149 1092 2183
rect 1104 2149 1116 2183
rect 1128 2149 1140 2183
rect 1152 2149 1164 2183
rect 1176 2149 1188 2183
rect 1200 2149 1212 2183
rect 1224 2149 1236 2183
rect 1248 2149 1260 2183
rect 1272 2149 1284 2183
rect 1296 2149 1308 2183
rect 1320 2149 1332 2183
rect 1344 2149 1356 2183
rect 1368 2149 1380 2183
rect 48 1909 60 1943
rect 72 1909 84 1943
rect 96 1909 108 1943
rect 120 1909 132 1943
rect 144 1909 156 1943
rect 168 1909 180 1943
rect 192 1909 204 1943
rect 216 1909 228 1943
rect 240 1909 252 1943
rect 264 1909 276 1943
rect 288 1909 300 1943
rect 312 1909 324 1943
rect 336 1909 348 1943
rect 360 1909 372 1943
rect 384 1909 396 1943
rect 408 1909 420 1943
rect 432 1909 444 1943
rect 456 1909 468 1943
rect 480 1909 492 1943
rect 504 1909 516 1943
rect 528 1909 540 1943
rect 552 1909 564 1943
rect 576 1909 588 1943
rect 600 1909 612 1943
rect 624 1909 636 1943
rect 648 1909 660 1943
rect 672 1909 684 1943
rect 696 1909 708 1943
rect 720 1909 732 1943
rect 744 1909 756 1943
rect 768 1909 780 1943
rect 792 1909 804 1943
rect 816 1909 828 1943
rect 840 1909 852 1943
rect 864 1909 876 1943
rect 888 1909 900 1943
rect 912 1909 924 1943
rect 936 1909 948 1943
rect 960 1909 972 1943
rect 984 1909 996 1943
rect 1008 1909 1020 1943
rect 1032 1909 1044 1943
rect 1056 1909 1068 1943
rect 1080 1909 1092 1943
rect 1104 1909 1116 1943
rect 1128 1909 1140 1943
rect 1152 1909 1164 1943
rect 1176 1909 1188 1943
rect 1200 1909 1212 1943
rect 1224 1909 1236 1943
rect 1248 1909 1260 1943
rect 1272 1909 1284 1943
rect 1296 1909 1308 1943
rect 1320 1909 1332 1943
rect 1344 1909 1356 1943
rect 1368 1909 1380 1943
rect 1392 1909 1404 1943
rect 48 1669 60 1703
rect 72 1669 84 1703
rect 96 1669 108 1703
rect 120 1669 132 1703
rect 144 1669 156 1703
rect 168 1669 180 1703
rect 192 1669 204 1703
rect 216 1669 228 1703
rect 240 1669 252 1703
rect 264 1669 276 1703
rect 288 1669 300 1703
rect 312 1669 324 1703
rect 336 1669 348 1703
rect 360 1669 372 1703
rect 384 1669 396 1703
rect 408 1669 420 1703
rect 432 1669 444 1703
rect 456 1669 468 1703
rect 480 1669 492 1703
rect 504 1669 516 1703
rect 528 1669 540 1703
rect 552 1669 564 1703
rect 576 1669 588 1703
rect 600 1669 612 1703
rect 624 1669 636 1703
rect 648 1669 660 1703
rect 672 1669 684 1703
rect 696 1669 708 1703
rect 720 1669 732 1703
rect 744 1669 756 1703
rect 768 1669 780 1703
rect 792 1669 804 1703
rect 816 1669 828 1703
rect 840 1669 852 1703
rect 864 1669 876 1703
rect 888 1669 900 1703
rect 912 1669 924 1703
rect 936 1669 948 1703
rect 960 1669 972 1703
rect 984 1669 996 1703
rect 1008 1669 1020 1703
rect 1032 1669 1044 1703
rect 1056 1669 1068 1703
rect 1080 1669 1092 1703
rect 1104 1669 1116 1703
rect 1128 1669 1140 1703
rect 1152 1669 1164 1703
rect 1176 1669 1188 1703
rect 1200 1669 1212 1703
rect 1224 1669 1236 1703
rect 1248 1669 1260 1703
rect 1272 1669 1284 1703
rect 1296 1669 1308 1703
rect 1320 1669 1332 1703
rect 1344 1669 1356 1703
rect 1368 1669 1380 1703
rect 1392 1669 1404 1703
rect 1416 1669 1428 1703
rect 48 1429 60 1463
rect 72 1429 84 1463
rect 96 1429 108 1463
rect 120 1429 132 1463
rect 144 1429 156 1463
rect 168 1429 180 1463
rect 192 1429 204 1463
rect 216 1429 228 1463
rect 240 1429 252 1463
rect 264 1429 276 1463
rect 288 1429 300 1463
rect 312 1429 324 1463
rect 336 1429 348 1463
rect 360 1429 372 1463
rect 384 1429 396 1463
rect 408 1429 420 1463
rect 432 1429 444 1463
rect 456 1429 468 1463
rect 480 1429 492 1463
rect 504 1429 516 1463
rect 528 1429 540 1463
rect 552 1429 564 1463
rect 576 1429 588 1463
rect 600 1429 612 1463
rect 624 1429 636 1463
rect 648 1429 660 1463
rect 672 1429 684 1463
rect 696 1429 708 1463
rect 720 1429 732 1463
rect 744 1429 756 1463
rect 768 1429 780 1463
rect 792 1429 804 1463
rect 816 1429 828 1463
rect 840 1429 852 1463
rect 864 1429 876 1463
rect 888 1429 900 1463
rect 912 1429 924 1463
rect 936 1429 948 1463
rect 960 1429 972 1463
rect 984 1429 996 1463
rect 1008 1429 1020 1463
rect 1032 1429 1044 1463
rect 1056 1429 1068 1463
rect 1080 1429 1092 1463
rect 1104 1429 1116 1463
rect 1128 1429 1140 1463
rect 1152 1429 1164 1463
rect 1176 1429 1188 1463
rect 1200 1429 1212 1463
rect 1224 1429 1236 1463
rect 1248 1429 1260 1463
rect 48 1189 60 1223
rect 72 1189 84 1223
rect 96 1189 108 1223
rect 120 1189 132 1223
rect 144 1189 156 1223
rect 168 1189 180 1223
rect 192 1189 204 1223
rect 216 1189 228 1223
rect 240 1189 252 1223
rect 264 1189 276 1223
rect 288 1189 300 1223
rect 312 1189 324 1223
rect 336 1189 348 1223
rect 360 1189 372 1223
rect 384 1189 396 1223
rect 408 1189 420 1223
rect 432 1189 444 1223
rect 456 1189 468 1223
rect 480 1189 492 1223
rect 504 1189 516 1223
rect 528 1189 540 1223
rect 552 1189 564 1223
rect 576 1189 588 1223
rect 600 1189 612 1223
rect 624 1189 636 1223
rect 648 1189 660 1223
rect 672 1189 684 1223
rect 696 1189 708 1223
rect 720 1189 732 1223
rect 744 1189 756 1223
rect 768 1189 780 1223
rect 792 1189 804 1223
rect 816 1189 828 1223
rect 840 1189 852 1223
rect 864 1189 876 1223
rect 888 1189 900 1223
rect 912 1189 924 1223
rect 936 1189 948 1223
rect 960 1189 972 1223
rect 984 1189 996 1223
rect 1008 1189 1020 1223
rect 1032 1189 1044 1223
rect 48 949 60 983
rect 72 949 84 983
rect 96 949 108 983
rect 120 949 132 983
rect 144 949 156 983
rect 168 949 180 983
rect 192 949 204 983
rect 216 949 228 983
rect 240 949 252 983
rect 264 949 276 983
rect 288 949 300 983
rect 312 949 324 983
rect 336 949 348 983
rect 360 949 372 983
rect 384 949 396 983
rect 408 949 420 983
rect 432 949 444 983
rect 456 949 468 983
rect 480 949 492 983
rect 504 949 516 983
rect 528 949 540 983
rect 552 949 564 983
rect 576 949 588 983
rect 600 949 612 983
rect 624 949 636 983
rect 648 949 660 983
rect 672 949 684 983
rect 696 949 708 983
rect 720 949 732 983
rect 744 949 756 983
rect 768 949 780 983
rect 792 949 804 983
rect 816 949 828 983
rect 48 709 60 743
rect 72 709 84 743
rect 96 709 108 743
rect 120 709 132 743
rect 144 709 156 743
rect 168 709 180 743
rect 192 709 204 743
rect 216 709 228 743
rect 240 709 252 743
rect 264 709 276 743
rect 288 709 300 743
rect 312 709 324 743
rect 336 709 348 743
rect 360 709 372 743
rect 384 709 396 743
rect 408 709 420 743
rect 432 709 444 743
rect 456 709 468 743
rect 480 709 492 743
rect 504 709 516 743
rect 528 709 540 743
rect 552 709 564 743
rect 576 709 588 743
rect 600 709 612 743
rect 624 709 636 743
rect 48 469 60 503
rect 72 469 84 503
rect 96 469 108 503
rect 120 469 132 503
rect 144 469 156 503
rect 168 469 180 503
rect 192 469 204 503
rect 216 469 228 503
rect 240 469 252 503
rect 264 469 276 503
rect 288 469 300 503
rect 312 469 324 503
rect 336 469 348 503
rect 360 469 372 503
rect 384 469 396 503
rect 408 469 420 503
rect 432 469 444 503
rect 48 229 60 263
rect 72 229 84 263
rect 96 229 108 263
rect 120 229 132 263
rect 144 229 156 263
rect 168 229 180 263
rect 192 229 204 263
rect 216 229 228 263
rect 120 -24 132 95
rect 528 -24 540 575
rect 744 -24 756 839
rect 1152 -24 1164 863
rect 1368 -24 1380 1559
rect 1728 -24 1740 1679
rect 1776 -24 1788 1703
rect 1992 -24 2004 1727
rect 2352 -24 2364 1751
rect 2400 -24 2412 1775
rect 2544 -24 2556 1799
rect 2568 -24 2580 1823
rect 2616 517 2628 1823
rect 2592 -24 2604 503
rect 2640 -24 2652 1823
rect 2664 -24 2676 1847
rect 2688 -24 2700 503
rect 2736 469 2748 1847
rect 2712 -24 2724 455
rect 2760 -24 2772 1847
rect 2784 -24 2796 1871
rect 2808 -24 2820 1895
rect 2832 -24 2844 1919
rect 2880 1069 2892 1919
rect 2856 -24 2868 1055
rect 2904 -24 2916 1919
rect 2928 -24 2940 1943
rect 2952 -24 2964 1967
rect 2976 -24 2988 1991
rect 3024 709 3036 1991
rect 3000 -24 3012 695
rect 3048 -24 3060 1991
rect 3072 -24 3084 2015
rect 3096 -24 3108 2039
rect 3120 -24 3132 2063
rect 3168 685 3180 2063
rect 3144 -24 3156 671
rect 3192 -24 3204 2063
rect 3216 -24 3228 2087
rect 3264 1813 3276 2087
rect 3240 -24 3252 1799
rect 3288 -24 3300 2087
rect 3360 1837 3372 2087
rect 3312 -24 3324 1439
rect 3336 -24 3348 1823
rect 3384 -24 3396 2087
rect 3408 -24 3420 2111
rect 3432 -24 3444 2135
rect 3480 1741 3492 2135
rect 3456 -24 3468 1727
rect 3576 -24 3588 2135
rect 3936 -24 3948 2159
rect 3984 -24 3996 2183
rect 4200 -24 4212 2207
rect 4560 -24 4572 2231
rect 4608 -24 4620 2255
rect 4752 -24 4764 2279
rect 4776 -24 4788 2303
rect 4848 1333 4860 2303
rect 4800 -24 4812 1055
rect 4824 -24 4836 1319
rect 4872 -24 4884 2303
rect 4896 -24 4908 2327
rect 4920 -24 4932 2351
rect 4992 781 5004 2351
rect 4944 -24 4956 695
rect 4968 -24 4980 767
rect 5016 -24 5028 2351
rect 5040 -24 5052 2375
rect 5064 -24 5076 2399
rect 5112 853 5124 2399
rect 5088 -24 5100 839
rect 5136 -24 5148 2399
rect 5160 -24 5172 2423
rect 5184 -24 5196 2447
rect 5232 109 5244 2447
rect 5208 -24 5220 95
rect 5256 -24 5268 2447
rect 5280 -24 5292 2471
rect 5304 -24 5316 2495
rect 5352 1573 5364 2495
rect 5328 -24 5340 1559
rect 5376 -24 5388 2495
rect 5400 -24 5412 2519
rect 5448 1429 5460 2519
rect 5424 -24 5436 1415
rect 5472 -24 5484 2519
rect 5496 -24 5508 2279
rect 5520 -24 5532 2543
rect 5544 -24 5556 2567
rect 5592 1381 5604 2567
rect 5568 -24 5580 1367
rect 5616 -24 5628 2567
rect 5640 -24 5652 2591
rect 5688 1261 5700 2591
rect 5664 -24 5676 1247
rect 5712 -24 5724 2591
rect 5736 -24 5748 2615
rect 5760 -24 5772 2639
rect 5832 997 5844 2639
rect 5784 -24 5796 503
rect 5808 -24 5820 983
rect 5856 -24 5868 2639
rect 5952 1909 5964 2639
rect 5880 -24 5892 1103
rect 5928 -24 5940 1895
rect 5976 -24 5988 2639
rect 6072 1837 6084 2639
rect 6000 -24 6012 575
rect 6048 -24 6060 1823
rect 6096 -24 6108 47
rect 6120 -24 6132 2639
rect 6168 2365 6180 2639
rect 6144 -24 6156 2351
rect 6192 -24 6204 119
rect 6216 -24 6228 2351
rect 6264 2101 6276 2615
rect 6240 -24 6252 2087
rect 6288 -24 6300 2615
rect 6312 -24 6324 2639
rect 6384 1981 6396 2639
rect 6480 2461 6492 2615
rect 6360 -24 6372 1967
rect 6408 -24 6420 71
rect 6432 -24 6444 2351
rect 6456 -24 6468 2447
rect 6576 -24 6588 2615
rect 6936 -24 6948 2639
rect 6984 -24 6996 2663
rect 7200 -24 7212 2687
rect 7608 -24 7620 2711
rect 7824 2413 7836 2711
rect 7752 -24 7764 -1
rect 7776 -24 7788 2351
rect 7800 -24 7812 2399
rect 7848 -24 7860 2711
rect 7872 -24 7884 2519
rect 7896 -24 7908 2735
rect 7920 -24 7932 2759
rect 7968 1093 7980 2759
rect 7944 -24 7956 1079
rect 7992 -24 8004 2759
rect 8016 -24 8028 2783
rect 8040 -24 8052 2807
rect 8088 1045 8100 2807
rect 8064 -24 8076 1031
rect 8112 -24 8124 2807
rect 8136 -24 8148 2783
rect 8160 -24 8172 2831
rect 8208 1021 8220 2831
rect 8184 -24 8196 1007
rect 8232 -24 8244 2831
rect 8256 -24 8268 2855
rect 8304 2221 8316 2855
rect 8280 -24 8292 2207
rect 8328 -24 8340 2855
rect 8352 -24 8364 2879
rect 8424 2053 8436 2879
rect 8520 2077 8532 2855
rect 8400 -24 8412 2039
rect 8448 -24 8460 1823
rect 8472 -24 8484 1055
rect 8496 -24 8508 2063
rect 8544 -24 8556 2855
rect 8568 -24 8580 2879
rect 8592 -24 8604 2903
rect 8616 -24 8628 2927
rect 8664 2149 8676 2927
rect 8640 -24 8652 2135
rect 8688 -24 8700 2927
rect 8736 1525 8748 2927
rect 8712 -24 8724 1511
rect 8760 109 8772 2903
rect 8736 -24 8748 95
rect 8784 -24 8796 2903
rect 8856 2437 8868 2903
rect 8808 -24 8820 575
rect 8832 -24 8844 2423
rect 8880 -24 8892 2423
rect 8952 2389 8964 2879
rect 8904 -24 8916 863
rect 8928 -24 8940 2375
rect 9024 1549 9036 2855
rect 8976 -24 8988 1511
rect 9000 -24 9012 1535
rect 9048 853 9060 2831
rect 9144 2485 9156 2807
rect 9024 -24 9036 839
rect 9072 -24 9084 2423
rect 9096 -24 9108 1703
rect 9120 -24 9132 2471
rect 9216 1597 9228 2783
rect 9168 -24 9180 1511
rect 9192 -24 9204 1583
rect 9240 1573 9252 2759
rect 9216 -24 9228 1559
rect 9264 -24 9276 2423
rect 9336 2125 9348 2735
rect 9288 -24 9300 1775
rect 9312 -24 9324 2111
rect 9360 -24 9372 1511
rect 9384 -24 9396 1607
rect 9408 -24 9420 1727
rect 9432 1621 9444 2711
rect 9552 2581 9564 2687
rect 9456 1741 9468 1799
rect 9456 -24 9468 1727
rect 9480 -24 9492 1799
rect 9504 -24 9516 1655
rect 9528 -24 9540 2567
rect 9648 2509 9660 2663
rect 9576 -24 9588 599
rect 9624 -24 9636 2495
rect 9696 -24 9708 2663
rect 9720 -24 9732 1415
rect 9744 -24 9756 2687
rect 9768 -24 9780 2711
rect 9816 1285 9828 2711
rect 9792 -24 9804 1271
rect 9840 -24 9852 2711
rect 9864 -24 9876 503
rect 9888 -24 9900 2735
rect 9936 1189 9948 2735
rect 9912 -24 9924 1175
rect 9960 -24 9972 2735
rect 9984 -24 9996 2759
rect 10008 -24 10020 503
rect 10032 -24 10044 2783
rect 10080 1165 10092 2783
rect 10056 -24 10068 1151
rect 10104 -24 10116 2783
rect 10128 -24 10140 2807
rect 10176 925 10188 2807
rect 10152 -24 10164 911
rect 10200 -24 10212 2807
rect 10272 1333 10284 2807
rect 10248 -24 10260 1319
rect 10320 -24 10332 2807
rect 10344 -24 10356 2831
rect 10416 781 10428 2831
rect 10392 -24 10404 767
rect 10440 -24 10452 2255
rect 10464 -24 10476 2255
rect 10512 853 10524 2807
rect 10488 -24 10500 839
rect 10536 -24 10548 2807
rect 10608 997 10620 2807
rect 10584 -24 10596 983
rect 10656 -24 10668 2807
rect 10680 -24 10692 2831
rect 10704 -24 10716 2855
rect 10728 -24 10740 2879
rect 10776 2629 10788 2879
rect 10752 -24 10764 2615
rect 10800 -24 10812 2879
rect 10824 -24 10836 2903
rect 10848 -24 10860 2927
rect 10872 -24 10884 2951
rect 10920 2077 10932 2951
rect 10896 -24 10908 2063
rect 10944 -24 10956 2951
rect 10968 -24 10980 2975
rect 10992 -24 11004 1055
rect 11040 613 11052 2975
rect 11016 -24 11028 599
rect 11064 -24 11076 2975
rect 11088 -24 11100 2999
rect 11112 -24 11124 1367
rect 11136 -24 11148 3023
rect 11184 1909 11196 3023
rect 11160 -24 11172 1895
rect 11208 -24 11220 3023
rect 11232 -24 11244 3047
rect 11280 2581 11292 3047
rect 11256 -24 11268 2567
rect 11304 -24 11316 3047
rect 11328 -24 11340 3071
rect 11352 -24 11364 3095
rect 11376 -24 11388 3119
rect 11424 757 11436 3119
rect 11400 -24 11412 743
rect 11448 -24 11460 3119
rect 11472 -24 11484 3143
rect 11520 1237 11532 3143
rect 11496 -24 11508 1223
rect 11544 -24 11556 2615
rect 11568 -24 11580 3143
rect 11592 -24 11604 3167
rect 11616 -24 11628 3191
rect 11664 949 11676 3191
rect 11640 -24 11652 935
rect 11688 -24 11700 3191
rect 11712 -24 11724 3215
rect 11736 -24 11748 1871
rect 11760 -24 11772 1055
rect 11808 661 11820 3215
rect 11784 -24 11796 647
rect 11832 -24 11844 3215
rect 11856 -24 11868 1991
rect 11880 -24 11892 3239
rect 11904 -24 11916 671
rect 11952 637 11964 3239
rect 11928 -24 11940 623
rect 11976 -24 11988 3239
rect 12000 -24 12012 3263
rect 12024 -24 12036 3287
rect 12048 -24 12060 2207
rect 12096 805 12108 3287
rect 12072 -24 12084 791
rect 12120 -24 12132 3287
rect 12144 -24 12156 3311
rect 12168 -24 12180 3335
rect 12192 -24 12204 3359
rect 12240 1333 12252 3359
rect 12216 -24 12228 1319
rect 12264 -24 12276 3359
rect 12288 -24 12300 3383
rect 12336 2461 12348 3383
rect 12312 -24 12324 2447
rect 12360 -24 12372 3383
rect 12384 -24 12396 3407
rect 12456 2557 12468 3407
rect 12432 -24 12444 2543
rect 12552 1837 12564 3383
rect 12480 -24 12492 1799
rect 12504 -24 12516 1655
rect 12528 -24 12540 1823
rect 12576 -24 12588 3383
rect 12600 -24 12612 3407
rect 12624 -24 12636 3431
rect 12648 -24 12660 3455
rect 12696 997 12708 3455
rect 12672 -24 12684 983
rect 12720 -24 12732 3455
rect 12744 -24 12756 3479
rect 12792 2797 12804 3479
rect 12768 -24 12780 2783
rect 12816 -24 12828 3479
rect 12840 -24 12852 3503
rect 12888 1525 12900 3503
rect 12864 -24 12876 1511
rect 12912 -24 12924 2687
rect 12984 1309 12996 3479
rect 12960 -24 12972 1295
rect 13032 -24 13044 3479
rect 13056 -24 13068 3503
rect 13128 781 13140 3503
rect 13104 -24 13116 767
rect 13152 -24 13164 3503
rect 13176 -24 13188 2783
rect 13224 1597 13236 3503
rect 13200 -24 13212 1583
rect 13248 -24 13260 3119
rect 13320 829 13332 3479
rect 13296 -24 13308 815
rect 13368 -24 13380 2591
rect 13392 -24 13404 3479
rect 13440 901 13452 3479
rect 13416 -24 13428 887
rect 13464 -24 13476 3479
rect 13488 -24 13500 3503
rect 13512 -24 13524 3527
rect 13560 2437 13572 3527
rect 13536 -24 13548 2423
rect 13584 -24 13596 3527
rect 13608 -24 13620 3551
rect 13680 2389 13692 3551
rect 13656 -24 13668 2375
rect 13704 -24 13716 3551
rect 13776 2125 13788 3551
rect 13752 -24 13764 2111
rect 13824 -24 13836 1703
rect 13896 -24 13908 3551
rect 13992 85 14004 3551
rect 13968 -24 13980 71
rect 14040 -24 14052 3551
rect 14208 325 14220 3551
rect 14112 -24 14124 71
rect 14184 -24 14196 311
rect 14256 -24 14268 3551
rect 14280 -24 14292 3575
rect 14352 1813 14364 3575
rect 14328 -24 14340 1799
rect 14376 -24 14388 3551
rect 14400 -24 14412 3575
rect 14448 2701 14460 3575
rect 14424 -24 14436 2687
rect 14472 -24 14484 3575
rect 14544 1837 14556 3575
rect 14496 -24 14508 479
rect 14520 -24 14532 1823
rect 14568 -24 14580 3575
rect 14592 -24 14604 3599
rect 14640 2749 14652 3599
rect 14616 -24 14628 2735
rect 14664 -24 14676 3599
rect 14688 -24 14700 3623
rect 14736 2485 14748 3623
rect 14712 -24 14724 2471
rect 14760 -24 14772 3623
rect 14784 -24 14796 3551
rect 14832 469 14844 3623
rect 14808 -24 14820 455
rect 14856 -24 14868 3551
rect 14880 -24 14892 3623
rect 14928 3133 14940 3623
rect 14904 -24 14916 3119
rect 14952 -24 14964 3479
rect 14976 -24 14988 3623
rect 15024 1189 15036 3623
rect 15000 -24 15012 1175
rect 15048 -24 15060 3623
rect 15072 -24 15084 3647
rect 15096 -24 15108 3671
rect 15144 2293 15156 3671
rect 15120 -24 15132 2279
rect 15168 -24 15180 311
rect 15336 205 15348 3647
rect 15240 -24 15252 71
rect 15312 -24 15324 191
rect 15384 -24 15396 3647
rect 15408 -24 15420 3671
rect 15480 2269 15492 3671
rect 15432 -24 15444 1727
rect 15456 -24 15468 2255
rect 15672 445 15684 3647
rect 15504 -24 15516 311
rect 15576 -24 15588 71
rect 15648 -24 15660 431
rect 15888 421 15900 3623
rect 15720 -24 15732 311
rect 15792 -24 15804 71
rect 15864 -24 15876 407
rect 16104 397 16116 3599
rect 15936 -24 15948 311
rect 16008 -24 16020 71
rect 16080 -24 16092 383
rect 16320 373 16332 3575
rect 16152 -24 16164 311
rect 16224 -24 16236 71
rect 16296 -24 16308 359
rect 16536 349 16548 3551
rect 16368 -24 16380 311
rect 16440 -24 16452 71
rect 16512 -24 16524 335
rect 16584 -24 16596 311
rect 16752 301 16764 3527
rect 16656 -24 16668 71
rect 16728 -24 16740 287
rect 16800 -24 16812 311
rect 16968 277 16980 3503
rect 16872 -24 16884 71
rect 16944 -24 16956 263
rect 17016 -24 17028 311
rect 17184 229 17196 3479
rect 17088 -24 17100 71
rect 17160 -24 17172 215
rect 17232 -24 17244 311
rect 17400 181 17412 3455
rect 17472 325 17484 3431
rect 17304 -24 17316 71
rect 17376 -24 17388 167
rect 17448 -24 17460 311
rect 17616 157 17628 3407
rect 17520 -24 17532 71
rect 17592 -24 17604 143
rect 17664 -24 17676 1775
rect 17832 133 17844 3383
rect 17904 877 17916 3359
rect 17736 -24 17748 71
rect 17808 -24 17820 119
rect 17880 -24 17892 863
rect 17952 -24 17964 71
rect 18048 61 18060 3335
rect 18024 -24 18036 47
rect 18096 -24 18108 575
rect 18168 -24 18180 71
rect 18264 37 18276 3311
rect 18240 -24 18252 -1
rect 18312 -24 18324 3311
rect 18336 -24 18348 3335
rect 18360 -24 18372 3359
rect 18408 877 18420 3359
rect 18384 -24 18396 863
rect 18432 -24 18444 3359
rect 18456 -24 18468 3383
rect 18480 -24 18492 3407
rect 18528 2125 18540 3407
rect 18504 -24 18516 2111
rect 18552 -24 18564 3407
rect 18576 -24 18588 3431
rect 18624 3037 18636 3431
rect 18600 -24 18612 3023
rect 18648 -24 18660 3431
rect 18672 -24 18684 3455
rect 18744 2941 18756 3455
rect 18720 -24 18732 2927
rect 18768 -24 18780 3455
rect 18792 -24 18804 3479
rect 18840 3253 18852 3479
rect 18816 -24 18828 3239
rect 18864 -24 18876 191
rect 18888 -24 18900 3479
rect 18936 37 18948 3479
rect 18912 -24 18924 -1
rect 18960 -24 18972 3479
rect 18984 -24 18996 3503
rect 19056 3013 19068 3503
rect 19032 -24 19044 2999
rect 19080 -24 19092 3095
rect 19104 -24 19116 3503
rect 19152 1405 19164 3503
rect 19128 -24 19140 1391
rect 19176 -24 19188 3503
rect 19200 -24 19212 3527
rect 19248 829 19260 3527
rect 19224 -24 19236 815
rect 19272 -24 19284 3527
rect 19296 -24 19308 3551
rect 19368 2869 19380 3551
rect 19344 -24 19356 2855
rect 19392 -24 19404 3551
rect 19416 -24 19428 3575
rect 19488 2677 19500 3575
rect 19464 -24 19476 2663
rect 19512 -24 19524 3575
rect 19584 637 19596 3575
rect 19560 -24 19572 623
rect 19632 -24 19644 1151
rect 19656 -24 19668 3575
rect 19728 2605 19740 3575
rect 19704 -24 19716 2591
rect 19824 -24 19836 3575
rect 20184 -24 20196 935
rect 20232 -24 20244 3599
rect 20376 -24 20388 599
rect 20400 -24 20412 2951
rect 20448 565 20460 3599
rect 20424 -24 20436 551
rect 20472 -24 20484 1199
rect 20496 -24 20508 3599
rect 20520 -24 20532 959
rect 20568 61 20580 3599
rect 20544 -24 20556 47
rect 20592 -24 20604 3599
rect 20664 3181 20676 3599
rect 20640 -24 20652 3167
rect 20712 -24 20724 191
rect 20736 -24 20748 3599
rect 20784 3085 20796 3599
rect 20760 -24 20772 3071
rect 20808 -24 20820 191
rect 20832 -24 20844 3599
rect 20880 1309 20892 3599
rect 20856 -24 20868 1295
rect 20904 -24 20916 359
rect 20928 -24 20940 3239
rect 20976 301 20988 3575
rect 20952 -24 20964 287
rect 21000 -24 21012 3575
rect 21024 -24 21036 3599
rect 21072 2797 21084 3599
rect 21048 -24 21060 2783
rect 21096 -24 21108 3599
rect 21120 -24 21132 3623
rect 21168 1045 21180 3623
rect 21144 -24 21156 1031
rect 21192 -24 21204 767
rect 21216 -24 21228 3599
rect 21264 1933 21276 3599
rect 21240 -24 21252 1919
rect 21288 -24 21300 191
rect 21312 -24 21324 3599
rect 21360 1429 21372 3599
rect 21336 -24 21348 1415
rect 21384 -24 21396 2255
rect 21456 1069 21468 3575
rect 21408 -24 21420 215
rect 21432 -24 21444 1055
rect 21480 -24 21492 3575
rect 21504 -24 21516 3599
rect 21552 1837 21564 3599
rect 21528 -24 21540 1823
rect 21576 -24 21588 3599
rect 21600 -24 21612 3623
rect 21624 -24 21636 3647
rect 21648 -24 21660 3671
rect 21696 2749 21708 3671
rect 21672 -24 21684 2735
rect 21720 -24 21732 2183
rect 21744 -24 21756 3671
rect 21768 -24 21780 3119
rect 21816 157 21828 3671
rect 21792 -24 21804 143
rect 21840 -24 21852 47
rect 21864 -24 21876 3671
rect 21936 349 21948 3671
rect 21912 -24 21924 335
rect 21960 -24 21972 3671
rect 21984 -24 21996 2207
rect 22056 1885 22068 3671
rect 22032 -24 22044 1871
rect 22080 -24 22092 3671
rect 22152 85 22164 3671
rect 22128 -24 22140 71
rect 22200 -24 22212 2015
rect 22224 -24 22236 3671
rect 22248 -24 22260 3695
rect 22272 -24 22284 3719
rect 22320 637 22332 3719
rect 22296 -24 22308 623
rect 22344 -24 22356 3719
rect 22368 -24 22380 3743
rect 22416 3037 22428 3743
rect 22392 -24 22404 3023
rect 22440 -24 22452 3743
rect 22464 -24 22476 3767
rect 22560 3277 22572 3767
rect 22488 -24 22500 143
rect 22512 -24 22524 1727
rect 22536 -24 22548 3263
rect 22584 -24 22596 3767
rect 22656 277 22668 3767
rect 22632 -24 22644 263
rect 22704 -24 22716 3767
rect 22728 -24 22740 2159
rect 22776 805 22788 3767
rect 22752 -24 22764 791
rect 22800 -24 22812 3767
rect 22824 -24 22836 3791
rect 22848 -24 22860 3815
rect 22920 3181 22932 3815
rect 22872 -24 22884 623
rect 22896 -24 22908 3167
rect 22944 -24 22956 47
rect 22968 -24 22980 3815
rect 23016 2533 23028 3815
rect 22992 -24 23004 2519
rect 23040 -24 23052 3815
rect 23064 -24 23076 3839
rect 23112 397 23124 3839
rect 23088 -24 23100 383
rect 23136 -24 23148 3839
rect 23160 -24 23172 3863
rect 23184 -24 23196 3887
rect 23208 -24 23220 1295
rect 23256 1189 23268 3887
rect 23232 -24 23244 1175
rect 23280 -24 23292 215
rect 23304 -24 23316 3887
rect 23328 -24 23340 3911
rect 23352 -24 23364 3935
rect 23400 1357 23412 3935
rect 23376 -24 23388 1343
rect 23424 -24 23436 3935
rect 23496 1117 23508 3935
rect 23472 -24 23484 1103
rect 23544 -24 23556 3935
rect 23568 -24 23580 3959
rect 23640 3109 23652 3959
rect 23592 -24 23604 1295
rect 23616 -24 23628 3095
rect 23664 -24 23676 1295
rect 23688 -24 23700 3959
rect 23712 -24 23724 3983
rect 23760 1381 23772 3983
rect 23736 -24 23748 1367
rect 23784 -24 23796 407
rect 23808 -24 23820 3959
rect 23880 2989 23892 3959
rect 23832 -24 23844 719
rect 23856 -24 23868 2975
rect 23904 -24 23916 3959
rect 23928 -24 23940 3983
rect 23952 -24 23964 3119
rect 24000 85 24012 3983
rect 23976 -24 23988 71
rect 24024 -24 24036 3983
rect 24048 -24 24060 71
rect 24072 -24 24084 4007
rect 24120 1261 24132 4007
rect 24096 -24 24108 1247
rect 24144 -24 24156 3935
rect 24168 -24 24180 4007
rect 24240 3061 24252 4007
rect 24192 -24 24204 719
rect 24216 -24 24228 3047
rect 24264 -24 24276 4007
rect 24288 -24 24300 4031
rect 24312 -24 24324 4055
rect 24360 301 24372 4055
rect 24336 -24 24348 287
rect 24384 -24 24396 4055
rect 24408 -24 24420 767
rect 24432 -24 24444 4079
rect 24480 2605 24492 4079
rect 24456 -24 24468 2591
rect 24504 -24 24516 4079
rect 24528 -24 24540 4103
rect 24552 -24 24564 4127
rect 24576 -24 24588 4151
rect 24624 3445 24636 4151
rect 24600 -24 24612 3431
rect 24648 -24 24660 1847
rect 24720 205 24732 4127
rect 24840 3349 24852 4103
rect 24696 -24 24708 191
rect 24768 -24 24780 143
rect 24792 -24 24804 3119
rect 24816 -24 24828 3335
rect 24864 -24 24876 4103
rect 24888 -24 24900 3959
rect 24960 2269 24972 4103
rect 24936 -24 24948 2255
rect 24984 -24 24996 3959
rect 25008 -24 25020 4103
rect 25056 1069 25068 4103
rect 25032 -24 25044 1055
rect 25080 -24 25092 143
rect 25104 -24 25116 4055
rect 25152 1981 25164 4079
rect 25128 -24 25140 1967
rect 25176 -24 25188 3455
rect 25200 -24 25212 4079
rect 25248 3205 25260 4079
rect 25224 -24 25236 3191
rect 25272 -24 25284 4079
rect 25296 -24 25308 3959
rect 25368 1933 25380 4079
rect 25344 -24 25356 1919
rect 25392 -24 25404 4079
rect 25464 3253 25476 4079
rect 25416 -24 25428 2423
rect 25440 -24 25452 3239
rect 25488 -24 25500 4079
rect 25512 -24 25524 3191
rect 25560 133 25572 4079
rect 25536 -24 25548 119
rect 25656 -24 25668 4079
rect 26016 -24 26028 2447
rect 26064 -24 26076 3263
rect 26208 -24 26220 3095
rect 26232 -24 26244 3191
rect 26280 613 26292 4079
rect 26256 -24 26268 599
rect 26304 -24 26316 3455
rect 26328 -24 26340 4079
rect 26376 3013 26388 4079
rect 26352 -24 26364 2999
rect 26400 -24 26412 4079
rect 26424 -24 26436 4103
rect 26448 -24 26460 4127
rect 26472 -24 26484 4151
rect 26520 277 26532 4151
rect 26496 -24 26508 263
rect 26544 -24 26556 4055
rect 26568 -24 26580 3959
rect 26616 3517 26628 4127
rect 26592 -24 26604 3503
rect 26640 -24 26652 143
rect 26664 -24 26676 4127
rect 26736 2677 26748 4127
rect 26712 -24 26724 2663
rect 26760 -24 26772 4127
rect 26784 -24 26796 3047
rect 26808 -24 26820 4151
rect 26856 3397 26868 4151
rect 26832 -24 26844 3383
rect 26880 -24 26892 4151
rect 26904 -24 26916 4175
rect 26976 3541 26988 4175
rect 26952 -24 26964 3527
rect 27000 -24 27012 3983
rect 27024 -24 27036 4175
rect 27048 -24 27060 4199
rect 27096 2341 27108 4199
rect 27072 -24 27084 2327
rect 27120 -24 27132 3959
rect 27144 -24 27156 215
rect 27168 -24 27180 1055
rect 27216 709 27228 4175
rect 27192 -24 27204 695
rect 27240 -24 27252 4175
rect 27264 -24 27276 4199
rect 27312 3733 27324 4199
rect 27288 -24 27300 3719
rect 27336 -24 27348 4199
rect 27360 -24 27372 119
rect 27384 -24 27396 1247
rect 27432 1237 27444 4199
rect 27408 -24 27420 1223
rect 27456 -24 27468 3455
rect 27480 -24 27492 4199
rect 27528 1525 27540 4199
rect 27504 -24 27516 1511
rect 27552 -24 27564 4199
rect 27576 -24 27588 4223
rect 27600 -24 27612 4247
rect 27624 -24 27636 4271
rect 27672 469 27684 4271
rect 27648 -24 27660 455
rect 27696 -24 27708 695
rect 27720 -24 27732 3983
rect 27768 2101 27780 4247
rect 27744 -24 27756 2087
rect 27792 -24 27804 3095
rect 27816 -24 27828 4247
rect 27864 1861 27876 4247
rect 27840 -24 27852 1847
rect 27888 -24 27900 4247
rect 27912 -24 27924 4271
rect 27960 805 27972 4271
rect 27936 -24 27948 791
rect 27984 -24 27996 3047
rect 28008 -24 28020 4271
rect 28056 3493 28068 4271
rect 28032 -24 28044 3479
rect 28080 -24 28092 3047
rect 28104 -24 28116 4271
rect 28152 2557 28164 4271
rect 28128 -24 28140 2543
rect 28176 -24 28188 3095
rect 28200 -24 28212 3383
rect 28272 61 28284 4247
rect 28248 -24 28260 47
rect 28296 -24 28308 3095
rect 28320 -24 28332 2543
rect 28368 1909 28380 4223
rect 28344 -24 28356 1895
rect 28392 -24 28404 3095
rect 28416 -24 28428 4223
rect 28464 1405 28476 4223
rect 28560 3301 28572 4199
rect 28440 -24 28452 1391
rect 28488 -24 28500 2975
rect 28512 -24 28524 1415
rect 28536 -24 28548 3287
rect 28584 -24 28596 2975
rect 28608 -24 28620 4199
rect 28656 661 28668 4199
rect 28632 -24 28644 647
rect 28680 -24 28692 2975
rect 28704 -24 28716 4199
rect 28752 2125 28764 4199
rect 28728 -24 28740 2111
rect 28776 -24 28788 4199
rect 28848 3373 28860 4199
rect 28800 -24 28812 2183
rect 28824 -24 28836 3359
rect 28872 -24 28884 1919
rect 28896 -24 28908 2591
rect 28944 829 28956 4175
rect 29040 3589 29052 4151
rect 29136 3829 29148 4127
rect 28920 -24 28932 815
rect 28968 -24 28980 2975
rect 28992 -24 29004 959
rect 29016 -24 29028 3575
rect 29064 -24 29076 1031
rect 29088 -24 29100 2591
rect 29112 -24 29124 3815
rect 29160 -24 29172 1223
rect 29184 -24 29196 119
rect 29208 -24 29220 2327
rect 29256 1117 29268 4103
rect 29232 -24 29244 1103
rect 29280 -24 29292 2975
rect 29304 -24 29316 4103
rect 29352 757 29364 4103
rect 29328 -24 29340 743
rect 29448 -24 29460 4103
rect 29856 -24 29868 3407
rect 30000 -24 30012 4127
rect 30024 -24 30036 4151
rect 30096 3565 30108 4151
rect 30072 -24 30084 3551
rect 30120 -24 30132 3359
rect 30144 -24 30156 4151
rect 30192 1885 30204 4151
rect 30168 -24 30180 1871
rect 30216 -24 30228 3599
rect 30240 -24 30252 4151
rect 30264 -24 30276 4175
rect 30312 3013 30324 4175
rect 30288 -24 30300 2999
rect 30336 -24 30348 4175
rect 30408 3685 30420 4175
rect 30384 -24 30396 3671
rect 30456 -24 30468 4175
rect 30480 -24 30492 4199
rect 30552 109 30564 4199
rect 30528 -24 30540 95
rect 30576 -24 30588 1943
rect 30600 -24 30612 2183
rect 30672 853 30684 4175
rect 30648 -24 30660 839
rect 30696 -24 30708 4175
rect 30720 -24 30732 3719
rect 30792 3589 30804 4175
rect 30744 -24 30756 2423
rect 30768 -24 30780 3575
rect 30816 -24 30828 647
rect 30840 -24 30852 3455
rect 30912 1093 30924 4151
rect 31032 3973 31044 4127
rect 30864 -24 30876 1055
rect 30888 -24 30900 1079
rect 30936 -24 30948 647
rect 30960 -24 30972 239
rect 31008 -24 31020 3959
rect 31056 -24 31068 767
rect 31080 -24 31092 647
rect 31152 157 31164 4103
rect 31128 -24 31140 143
rect 31176 -24 31188 1199
rect 31200 -24 31212 4103
rect 31272 1189 31284 4103
rect 31392 3205 31404 4079
rect 31224 -24 31236 239
rect 31248 -24 31260 1175
rect 31296 -24 31308 3119
rect 31320 -24 31332 647
rect 31368 -24 31380 3191
rect 31416 -24 31428 4079
rect 31440 -24 31452 4103
rect 31464 -24 31476 4127
rect 31512 613 31524 4127
rect 31488 -24 31500 599
rect 31536 -24 31548 647
rect 31560 -24 31572 4127
rect 31608 3253 31620 4127
rect 31728 3661 31740 4103
rect 31584 -24 31596 3239
rect 31632 -24 31644 1367
rect 31656 -24 31668 1175
rect 31680 -24 31692 239
rect 31704 -24 31716 3647
rect 31752 -24 31764 4103
rect 31776 -24 31788 4127
rect 31824 3181 31836 4127
rect 31800 -24 31812 3167
rect 31848 -24 31860 4127
rect 31872 -24 31884 4151
rect 31920 2941 31932 4151
rect 31896 -24 31908 2927
rect 31944 -24 31956 4151
rect 31968 -24 31980 4175
rect 31992 -24 32004 4199
rect 32040 157 32052 4199
rect 32016 -24 32028 143
rect 32064 -24 32076 3455
rect 32088 -24 32100 4199
rect 32136 1333 32148 4199
rect 32112 -24 32124 1319
rect 32160 -24 32172 4199
rect 32232 2365 32244 4199
rect 32208 -24 32220 2351
rect 32280 -24 32292 4199
rect 32304 -24 32316 4223
rect 32328 -24 32340 4247
rect 32352 -24 32364 4271
rect 32400 3685 32412 4271
rect 32376 -24 32388 3671
rect 32424 -24 32436 4271
rect 32448 -24 32460 4295
rect 32520 3925 32532 4295
rect 32496 -24 32508 3911
rect 32544 -24 32556 3623
rect 32568 -24 32580 3599
rect 32616 1525 32628 4271
rect 32592 -24 32604 1511
rect 32640 -24 32652 3215
rect 32664 -24 32676 4271
rect 32712 2677 32724 4271
rect 32688 -24 32700 2663
rect 32736 -24 32748 4271
rect 32760 -24 32772 4295
rect 32808 829 32820 4295
rect 32784 -24 32796 815
rect 32832 -24 32844 1919
rect 32856 -24 32868 4295
rect 32880 -24 32892 407
rect 32928 325 32940 4295
rect 32904 -24 32916 311
rect 32952 -24 32964 3983
rect 32976 -24 32988 4295
rect 33000 -24 33012 2327
rect 33048 1285 33060 4295
rect 33024 -24 33036 1271
rect 33072 -24 33084 4295
rect 33144 205 33156 4295
rect 33288 3205 33300 4271
rect 33120 -24 33132 191
rect 33192 -24 33204 239
rect 33216 -24 33228 -1
rect 33240 -24 33252 479
rect 33264 -24 33276 3191
rect 33312 -24 33324 3455
rect 33336 -24 33348 3743
rect 33408 2989 33420 4247
rect 33504 4045 33516 4223
rect 33384 -24 33396 2975
rect 33432 -24 33444 167
rect 33456 -24 33468 1487
rect 33480 -24 33492 4031
rect 33528 -24 33540 2711
rect 33552 -24 33564 4223
rect 33600 1597 33612 4223
rect 33696 3373 33708 4199
rect 33576 -24 33588 1583
rect 33624 -24 33636 1943
rect 33672 -24 33684 3359
rect 33744 -24 33756 3455
rect 33816 1837 33828 4175
rect 33768 -24 33780 743
rect 33792 -24 33804 1823
rect 33840 -24 33852 3455
rect 33936 3109 33948 4151
rect 33864 -24 33876 239
rect 33912 -24 33924 3095
rect 33960 -24 33972 4151
rect 34032 3973 34044 4151
rect 33984 -24 33996 863
rect 34008 -24 34020 3959
rect 34056 -24 34068 4151
rect 34128 2605 34140 4151
rect 34080 -24 34092 2423
rect 34104 -24 34116 2591
rect 34152 -24 34164 4151
rect 34176 -24 34188 2711
rect 34224 85 34236 4151
rect 34200 -24 34212 71
rect 34248 -24 34260 3455
rect 34344 3061 34356 4127
rect 34272 -24 34284 959
rect 34320 -24 34332 3047
rect 34368 -24 34380 767
rect 34392 -24 34404 3983
rect 34440 805 34452 4103
rect 34416 -24 34428 791
rect 34464 -24 34476 4103
rect 34488 -24 34500 2711
rect 34536 709 34548 4103
rect 34512 -24 34524 695
rect 34560 -24 34572 2711
rect 34632 133 34644 4079
rect 34608 -24 34620 119
rect 34680 -24 34692 4079
rect 34704 -24 34716 215
rect 34728 -24 34740 4103
rect 34800 2365 34812 4103
rect 34752 -24 34764 239
rect 34776 -24 34788 2351
rect 34824 -24 34836 4103
rect 34848 -24 34860 4127
rect 34896 2101 34908 4127
rect 34872 -24 34884 2087
rect 34920 -24 34932 4127
rect 34944 -24 34956 4079
rect 34992 3589 35004 4127
rect 34968 -24 34980 3575
rect 35016 -24 35028 4127
rect 35040 -24 35052 1367
rect 35088 805 35100 4127
rect 35064 -24 35076 791
rect 35112 -24 35124 4127
rect 35136 -24 35148 4151
rect 35208 3901 35220 4151
rect 35184 -24 35196 3887
rect 35232 -24 35244 4151
rect 35256 -24 35268 4175
rect 35328 3709 35340 4175
rect 35304 -24 35316 3695
rect 35352 -24 35364 4175
rect 35376 -24 35388 4199
rect 35400 -24 35412 4223
rect 35448 205 35460 4223
rect 35424 -24 35436 191
rect 35472 -24 35484 695
rect 35496 -24 35508 1487
rect 35568 853 35580 4199
rect 35544 -24 35556 839
rect 35592 -24 35604 311
rect 35616 -24 35628 2447
rect 35664 1621 35676 4175
rect 35640 -24 35652 1607
rect 35688 -24 35700 311
rect 35712 -24 35724 407
rect 35760 61 35772 4151
rect 35856 3325 35868 4127
rect 35736 -24 35748 47
rect 35784 -24 35796 311
rect 35808 -24 35820 1199
rect 35832 -24 35844 3311
rect 35880 -24 35892 311
rect 35904 -24 35916 3935
rect 35952 1957 35964 4103
rect 35928 -24 35940 1943
rect 35976 -24 35988 4103
rect 36048 4021 36060 4103
rect 36000 -24 36012 2399
rect 36024 -24 36036 4007
rect 36072 -24 36084 2591
rect 36144 661 36156 4079
rect 36264 2725 36276 4055
rect 36120 -24 36132 647
rect 36192 -24 36204 215
rect 36216 -24 36228 551
rect 36240 -24 36252 2711
rect 36288 -24 36300 4055
rect 36312 -24 36324 3719
rect 36360 2221 36372 4055
rect 36336 -24 36348 2207
rect 36384 -24 36396 2207
rect 36408 -24 36420 3551
rect 36456 2317 36468 4031
rect 36432 -24 36444 2303
rect 36552 181 36564 4007
rect 36480 -24 36492 71
rect 36528 -24 36540 167
rect 36600 -24 36612 311
rect 36648 -24 36660 3959
rect 36792 2773 36804 3959
rect 36720 -24 36732 2207
rect 36744 -24 36756 1871
rect 36768 -24 36780 2759
rect 36816 -24 36828 2207
rect 36840 -24 36852 2711
rect 36888 901 36900 3935
rect 36864 -24 36876 887
rect 36912 -24 36924 3935
rect 36936 -24 36948 3719
rect 37032 3349 37044 3935
rect 36960 -24 36972 3167
rect 36984 -24 36996 479
rect 37008 -24 37020 3335
rect 37056 -24 37068 3935
rect 37080 -24 37092 3263
rect 37128 3061 37140 3935
rect 37104 -24 37116 3047
rect 37152 -24 37164 3935
rect 37224 3661 37236 3935
rect 37176 -24 37188 3263
rect 37200 -24 37212 3647
rect 37248 -24 37260 2687
rect 37344 1189 37356 3911
rect 37272 -24 37284 959
rect 37320 -24 37332 1175
rect 37368 -24 37380 1391
rect 37392 -24 37404 3911
rect 37464 3637 37476 3911
rect 37440 -24 37452 3623
rect 37488 -24 37500 3911
rect 37512 -24 37524 1199
rect 37584 1189 37596 3911
rect 37560 -24 37572 1175
rect 37608 -24 37620 2447
rect 37632 -24 37644 3239
rect 37680 2677 37692 3887
rect 37656 -24 37668 2663
rect 37704 -24 37716 2495
rect 37728 -24 37740 3887
rect 37776 829 37788 3887
rect 37824 3421 37836 3863
rect 37752 -24 37764 815
rect 37800 -24 37812 3407
rect 37872 3109 37884 3839
rect 37824 -24 37836 503
rect 37848 -24 37860 3095
rect 37896 -24 37908 3839
rect 37968 3517 37980 3839
rect 37920 -24 37932 647
rect 37944 -24 37956 3503
rect 37992 -24 38004 2519
rect 38016 -24 38028 3119
rect 38040 -24 38052 1367
rect 38088 1093 38100 3815
rect 38064 -24 38076 1079
rect 38112 -24 38124 3815
rect 38184 2029 38196 3815
rect 38304 2965 38316 3791
rect 38160 -24 38172 2015
rect 38232 -24 38244 2207
rect 38256 -24 38268 2447
rect 38280 -24 38292 2951
rect 38328 -24 38340 647
rect 38352 -24 38364 3743
rect 38424 2773 38436 3767
rect 38520 2797 38532 3743
rect 38664 3469 38676 3719
rect 38400 -24 38412 2759
rect 38448 -24 38460 1223
rect 38496 -24 38508 2783
rect 38568 -24 38580 215
rect 38592 -24 38604 935
rect 38640 -24 38652 3455
rect 38688 -24 38700 2207
rect 38712 -24 38724 3143
rect 38760 997 38772 3695
rect 38856 2605 38868 3671
rect 38736 -24 38748 983
rect 38784 -24 38796 647
rect 38808 -24 38820 1199
rect 38832 -24 38844 2591
rect 38880 -24 38892 3671
rect 38904 -24 38916 3695
rect 38952 1285 38964 3695
rect 38928 -24 38940 1271
rect 38976 -24 38988 767
rect 39000 -24 39012 1871
rect 39048 85 39060 3671
rect 39024 -24 39036 71
rect 39072 -24 39084 71
rect 39096 -24 39108 2423
rect 39168 325 39180 3647
rect 39144 -24 39156 311
rect 39192 -24 39204 3647
rect 39216 -24 39228 3671
rect 39264 157 39276 3671
rect 39240 -24 39252 143
rect 39288 -24 39300 3671
rect 39360 2581 39372 3671
rect 39312 -24 39324 2399
rect 39336 -24 39348 2567
rect 39384 -24 39396 767
rect 39408 -24 39420 3263
rect 39456 709 39468 3647
rect 39432 -24 39444 695
rect 39480 -24 39492 3647
rect 39504 -24 39516 3671
rect 39552 37 39564 3671
rect 39528 -24 39540 -1
rect 39576 -24 39588 551
rect 39600 -24 39612 3671
rect 39648 1117 39660 3671
rect 39624 -24 39636 1103
rect 39672 -24 39684 3671
rect 39696 -24 39708 3695
rect 39768 1525 39780 3695
rect 39744 -24 39756 1511
rect 39792 -24 39804 3695
rect 39864 2677 39876 3695
rect 39816 -24 39828 1847
rect 39840 -24 39852 2663
rect 39888 -24 39900 3695
rect 39912 -24 39924 3167
rect 39960 2317 39972 3695
rect 39936 -24 39948 2303
rect 39984 -24 39996 2183
rect 40008 -24 40020 3335
rect 40056 805 40068 3671
rect 40152 3589 40164 3647
rect 40032 -24 40044 791
rect 40080 -24 40092 3335
rect 40104 -24 40116 1199
rect 40128 -24 40140 3575
rect 40176 -24 40188 3647
rect 40200 -24 40212 3263
rect 40248 61 40260 3647
rect 40224 -24 40236 47
rect 40272 -24 40284 3647
rect 40344 1957 40356 3647
rect 40296 -24 40308 1439
rect 40320 -24 40332 1943
rect 40368 -24 40380 3647
rect 40392 -24 40404 3671
rect 40440 1333 40452 3671
rect 40416 -24 40428 1319
rect 40464 -24 40476 3671
rect 40488 -24 40500 3695
rect 40512 -24 40524 2615
rect 40560 2029 40572 3695
rect 40536 -24 40548 2015
rect 40584 -24 40596 3695
rect 40656 1093 40668 3695
rect 40608 -24 40620 407
rect 40632 -24 40644 1079
rect 40680 -24 40692 863
rect 40704 -24 40716 2183
rect 40776 109 40788 3671
rect 40752 -24 40764 95
rect 40800 -24 40812 3671
rect 40824 -24 40836 2711
rect 40872 133 40884 3671
rect 40848 -24 40860 119
rect 40896 -24 40908 2423
rect 40992 1237 41004 3647
rect 40920 -24 40932 479
rect 40968 -24 40980 1223
rect 41016 -24 41028 3647
rect 41040 -24 41052 3671
rect 41088 181 41100 3671
rect 41184 541 41196 3647
rect 41064 -24 41076 167
rect 41112 -24 41124 503
rect 41160 -24 41172 527
rect 41232 -24 41244 3647
rect 41256 -24 41268 2183
rect 41304 1621 41316 3647
rect 41280 -24 41292 1607
rect 41328 -24 41340 3647
rect 41352 -24 41364 3143
rect 41400 1573 41412 3647
rect 41376 -24 41388 1559
rect 41424 -24 41436 1271
rect 41496 229 41508 3623
rect 41472 -24 41484 215
rect 41544 -24 41556 1559
rect 41568 -24 41580 3455
rect 41616 1165 41628 3599
rect 41592 -24 41604 1151
rect 41640 -24 41652 2495
rect 41664 -24 41676 3599
rect 41712 3445 41724 3599
rect 41688 -24 41700 3431
rect 41736 -24 41748 3599
rect 41808 3301 41820 3599
rect 41760 -24 41772 1055
rect 41784 -24 41796 3287
rect 41832 -24 41844 3599
rect 41856 -24 41868 3623
rect 41904 1405 41916 3623
rect 41880 -24 41892 1391
rect 41928 -24 41940 3407
rect 41952 -24 41964 1295
rect 42000 829 42012 3599
rect 41976 -24 41988 815
rect 42024 -24 42036 3599
rect 42048 -24 42060 3479
rect 42120 1189 42132 3599
rect 42096 -24 42108 1175
rect 42144 -24 42156 1151
rect 42216 757 42228 3575
rect 42192 -24 42204 743
rect 42264 -24 42276 1607
rect 42336 637 42348 3551
rect 42456 2125 42468 3527
rect 42312 -24 42324 623
rect 42384 -24 42396 -1
rect 42432 -24 42444 2111
rect 42504 -24 42516 1847
rect 42528 -24 42540 1415
rect 42600 277 42612 3503
rect 42696 2221 42708 3479
rect 42552 -24 42564 239
rect 42576 -24 42588 263
rect 42624 -24 42636 863
rect 42672 -24 42684 2207
rect 42744 -24 42756 1103
rect 42816 661 42828 3455
rect 42792 -24 42804 647
rect 42864 -24 42876 1559
rect 42888 -24 42900 1919
rect 42936 925 42948 3431
rect 42912 -24 42924 911
rect 42960 -24 42972 1559
rect 42984 -24 42996 1871
rect 43056 1141 43068 3407
rect 43032 -24 43044 1127
rect 43080 -24 43092 3335
rect 43152 3253 43164 3383
rect 43128 -24 43140 3239
rect 43200 -24 43212 3383
rect 43224 -24 43236 2399
rect 43272 517 43284 3383
rect 43248 -24 43260 503
rect 43296 -24 43308 2495
rect 43320 -24 43332 3383
rect 43368 3061 43380 3383
rect 43344 -24 43356 3047
rect 43392 -24 43404 3383
rect 43416 -24 43428 3407
rect 43464 325 43476 3407
rect 43440 -24 43452 311
rect 43488 -24 43500 2231
rect 43512 -24 43524 2231
rect 43560 1837 43572 3383
rect 43536 -24 43548 1823
rect 43584 -24 43596 1727
rect 43608 -24 43620 3383
rect 43656 2701 43668 3383
rect 43632 -24 43644 2687
rect 43752 2365 43764 3359
rect 43680 -24 43692 263
rect 43728 -24 43740 2351
rect 43800 -24 43812 2255
rect 43824 -24 43836 1247
rect 43872 277 43884 3335
rect 43848 -24 43860 263
rect 43896 -24 43908 551
rect 43920 -24 43932 1511
rect 43944 -24 43956 3311
rect 43992 -24 44004 3311
rect 44016 -24 44028 3335
rect 44064 2677 44076 3335
rect 44040 -24 44052 2663
rect 44088 -24 44100 1919
rect 44184 1549 44196 3311
rect 44352 2317 44364 3287
rect 44112 -24 44124 1031
rect 44136 -24 44148 1487
rect 44160 -24 44172 1535
rect 44232 -24 44244 2087
rect 44256 -24 44268 455
rect 44304 -24 44316 935
rect 44328 -24 44340 2303
rect 44400 -24 44412 3287
rect 44424 -24 44436 2087
rect 44472 1093 44484 3287
rect 44448 -24 44460 1079
rect 44496 -24 44508 1559
rect 44568 1021 44580 3263
rect 44544 -24 44556 1007
rect 44616 -24 44628 2279
rect 44640 -24 44652 239
rect 44712 229 44724 3239
rect 44688 -24 44700 215
rect 44736 -24 44748 1871
rect 44760 -24 44772 2639
rect 44808 181 44820 3215
rect 44784 -24 44796 167
rect 44832 -24 44844 335
rect 44856 -24 44868 1295
rect 44904 1165 44916 3191
rect 44880 -24 44892 1151
rect 44928 -24 44940 2783
rect 45000 2437 45012 3167
rect 44952 -24 44964 2279
rect 44976 -24 44988 2423
rect 45024 -24 45036 2639
rect 45048 -24 45060 2279
rect 45120 1621 45132 3143
rect 45096 -24 45108 1607
rect 45216 781 45228 3119
rect 45336 2053 45348 3095
rect 45144 -24 45156 71
rect 45192 -24 45204 767
rect 45264 -24 45276 527
rect 45312 -24 45324 2039
rect 45384 -24 45396 335
rect 45408 -24 45420 719
rect 45456 37 45468 3071
rect 45432 -24 45444 -1
rect 45480 -24 45492 1415
rect 45552 1357 45564 3047
rect 45648 2581 45660 3023
rect 45768 2821 45780 2999
rect 45504 -24 45516 1199
rect 45528 -24 45540 1343
rect 45576 -24 45588 503
rect 45624 -24 45636 2567
rect 45696 -24 45708 1031
rect 45720 -24 45732 1871
rect 45744 -24 45756 2807
rect 45792 -24 45804 1871
rect 45816 -24 45828 2999
rect 45864 2077 45876 2999
rect 45840 -24 45852 2063
rect 45888 -24 45900 2999
rect 45960 2773 45972 2999
rect 45912 -24 45924 1871
rect 45936 -24 45948 2759
rect 46056 1285 46068 2975
rect 45984 -24 45996 431
rect 46008 -24 46020 647
rect 46032 -24 46044 1271
rect 46080 -24 46092 2975
rect 46152 2389 46164 2975
rect 46104 -24 46116 647
rect 46128 -24 46140 2375
rect 46176 -24 46188 2375
rect 46200 -24 46212 2399
rect 46248 877 46260 2951
rect 46224 -24 46236 863
rect 46272 -24 46284 1031
rect 46296 -24 46308 647
rect 46368 373 46380 2927
rect 46344 -24 46356 359
rect 46392 -24 46404 887
rect 46416 -24 46428 1415
rect 46464 1237 46476 2903
rect 46440 -24 46452 1223
rect 46488 -24 46500 2903
rect 46512 -24 46524 383
rect 46560 133 46572 2903
rect 46536 -24 46548 119
rect 46584 -24 46596 1079
rect 46608 -24 46620 1655
rect 46680 781 46692 2879
rect 46656 -24 46668 767
rect 46704 -24 46716 2879
rect 46824 2845 46836 2879
rect 46728 -24 46740 935
rect 46752 -24 46764 2423
rect 46776 -24 46788 1367
rect 46800 -24 46812 2831
rect 46848 -24 46860 2879
rect 46872 -24 46884 2903
rect 46944 1957 46956 2903
rect 46896 -24 46908 1631
rect 46920 -24 46932 1943
rect 46968 -24 46980 2255
rect 46992 -24 47004 2519
rect 47064 805 47076 2879
rect 47040 -24 47052 791
rect 47088 -24 47100 2879
rect 47112 -24 47124 2447
rect 47160 1285 47172 2879
rect 47136 -24 47148 1271
rect 47184 -24 47196 1271
rect 47208 -24 47220 2783
rect 47256 61 47268 2855
rect 47232 -24 47244 47
rect 47280 -24 47292 2519
rect 47376 1333 47388 2831
rect 47304 -24 47316 407
rect 47328 -24 47340 215
rect 47352 -24 47364 1319
rect 47400 -24 47412 2279
rect 47472 1117 47484 2807
rect 47424 -24 47436 479
rect 47448 -24 47460 1103
rect 47496 -24 47508 2807
rect 47520 -24 47532 2831
rect 47544 -24 47556 2855
rect 47592 277 47604 2855
rect 47568 -24 47580 263
rect 47616 -24 47628 2399
rect 47640 -24 47652 383
rect 47664 -24 47676 2183
rect 47712 2149 47724 2831
rect 47688 -24 47700 2135
rect 47736 -24 47748 2831
rect 47832 1189 47844 2831
rect 47760 -24 47772 479
rect 47808 -24 47820 1175
rect 47880 -24 47892 2783
rect 47904 -24 47916 1199
rect 47952 -24 47964 2831
rect 48000 1357 48012 2831
rect 48120 2485 48132 2807
rect 47976 -24 47988 1343
rect 48048 -24 48060 167
rect 48096 -24 48108 2471
rect 48168 -24 48180 1991
rect 48192 -24 48204 2399
rect 48264 61 48276 2783
rect 48240 -24 48252 47
rect 48288 -24 48300 383
rect 48312 -24 48324 2399
rect 48384 1573 48396 2759
rect 48360 -24 48372 1559
rect 48408 -24 48420 2759
rect 48480 2029 48492 2759
rect 48432 -24 48444 47
rect 48456 -24 48468 2015
rect 48504 -24 48516 383
rect 48528 -24 48540 2399
rect 48576 1837 48588 2735
rect 48552 -24 48564 1823
rect 48600 -24 48612 2423
rect 48624 -24 48636 1847
rect 48672 1165 48684 2711
rect 48648 -24 48660 1151
rect 48696 -24 48708 1007
rect 48720 -24 48732 2711
rect 48768 205 48780 2711
rect 48744 -24 48756 191
rect 48792 -24 48804 551
rect 48864 373 48876 2687
rect 48816 -24 48828 191
rect 48840 -24 48852 359
rect 48888 -24 48900 431
rect 48912 -24 48924 935
rect 48960 85 48972 2663
rect 48936 -24 48948 71
rect 48984 -24 48996 1607
rect 49008 -24 49020 551
rect 49056 541 49068 2639
rect 49032 -24 49044 527
rect 49080 -24 49092 2639
rect 49104 -24 49116 551
rect 49152 301 49164 2639
rect 49128 -24 49140 287
rect 49176 -24 49188 2015
rect 49200 -24 49212 1631
rect 49248 997 49260 2615
rect 49224 -24 49236 983
rect 49272 -24 49284 1319
rect 49296 -24 49308 1199
rect 49344 757 49356 2591
rect 49320 -24 49332 743
rect 49368 -24 49380 2135
rect 49392 -24 49404 2471
rect 49440 373 49452 2567
rect 49536 829 49548 2543
rect 49416 -24 49428 359
rect 49464 -24 49476 71
rect 49488 -24 49500 215
rect 49512 -24 49524 815
rect 49560 -24 49572 2423
rect 49632 1237 49644 2519
rect 49584 -24 49596 959
rect 49608 -24 49620 1223
rect 49656 -24 49668 2423
rect 49680 -24 49692 2207
rect 49728 781 49740 2495
rect 49704 -24 49716 767
rect 49752 -24 49764 1991
rect 49776 -24 49788 1607
rect 49848 517 49860 2471
rect 49824 -24 49836 503
rect 49872 -24 49884 1175
rect 49968 1141 49980 2447
rect 49896 -24 49908 71
rect 49944 -24 49956 1127
rect 49992 -24 50004 2447
rect 50016 -24 50028 2471
rect 50064 925 50076 2471
rect 50160 2317 50172 2447
rect 50040 -24 50052 911
rect 50088 -24 50100 1943
rect 50112 -24 50124 791
rect 50136 -24 50148 2303
rect 50184 -24 50196 2015
rect 50208 -24 50220 1655
rect 50256 853 50268 2423
rect 50232 -24 50244 839
rect 50280 -24 50292 671
rect 50304 -24 50316 1127
rect 50352 877 50364 2399
rect 50328 -24 50340 863
rect 50448 -24 50460 695
rect 50832 157 50844 2375
rect 50880 2245 50892 2351
rect 50808 -24 50820 143
rect 50856 -24 50868 2231
rect 51000 -24 51012 191
rect 51024 -24 51036 2351
rect 51072 37 51084 2351
rect 51168 1597 51180 2327
rect 51048 -24 51060 -1
rect 51096 -24 51108 1031
rect 51120 -24 51132 1007
rect 51144 -24 51156 1583
rect 51192 -24 51204 2111
rect 51216 -24 51228 2327
rect 51264 325 51276 2327
rect 51384 2245 51396 2303
rect 51240 -24 51252 311
rect 51288 -24 51300 1847
rect 51312 -24 51324 551
rect 51336 -24 51348 239
rect 51360 -24 51372 2231
rect 51408 -24 51420 2111
rect 51432 -24 51444 1847
rect 51504 1285 51516 2279
rect 51480 -24 51492 1271
rect 51528 -24 51540 1607
rect 51600 661 51612 2255
rect 51576 -24 51588 647
rect 51648 -24 51660 47
rect 51672 -24 51684 2255
rect 51720 1549 51732 2255
rect 51864 1981 51876 2231
rect 51696 -24 51708 1535
rect 51744 -24 51756 407
rect 51768 -24 51780 1127
rect 51792 -24 51804 767
rect 51816 -24 51828 1295
rect 51840 -24 51852 1967
rect 51888 -24 51900 551
rect 51912 -24 51924 1055
rect 51984 661 51996 2207
rect 51960 -24 51972 647
rect 52008 -24 52020 1847
rect 52032 -24 52044 551
rect 52056 -24 52068 1439
rect 52104 109 52116 2183
rect 52200 1285 52212 2159
rect 52080 -24 52092 95
rect 52128 -24 52140 191
rect 52176 -24 52188 1271
rect 52248 -24 52260 383
rect 52320 157 52332 2135
rect 52440 1093 52452 2111
rect 52296 -24 52308 143
rect 52368 -24 52380 455
rect 52416 -24 52428 1079
rect 52488 -24 52500 2063
rect 52560 901 52572 2087
rect 52536 -24 52548 887
rect 52608 -24 52620 1919
rect 52632 -24 52644 935
rect 52680 613 52692 2063
rect 52656 -24 52668 599
rect 52704 -24 52716 1151
rect 52728 -24 52740 1919
rect 52800 181 52812 2039
rect 52896 1885 52908 2015
rect 52776 -24 52788 167
rect 52824 -24 52836 623
rect 52872 -24 52884 1871
rect 53016 349 53028 1991
rect 53136 1837 53148 1967
rect 52944 -24 52956 71
rect 52992 -24 53004 335
rect 53064 -24 53076 647
rect 53088 -24 53100 239
rect 53112 -24 53124 1823
rect 53232 1429 53244 1943
rect 53376 1525 53388 1919
rect 53160 -24 53172 1103
rect 53208 -24 53220 1415
rect 53280 -24 53292 239
rect 53304 -24 53316 1295
rect 53328 -24 53340 479
rect 53352 -24 53364 1511
rect 53400 -24 53412 1031
rect 53472 133 53484 1895
rect 53544 1021 53556 1871
rect 53448 -24 53460 119
rect 53520 -24 53532 1007
rect 53592 637 53604 1847
rect 53640 1789 53652 1823
rect 53544 -24 53556 95
rect 53568 -24 53580 623
rect 53616 -24 53628 1775
rect 53664 1693 53676 1799
rect 53640 -24 53652 1679
rect 53688 805 53700 1775
rect 53784 1381 53796 1751
rect 53664 -24 53676 791
rect 53712 -24 53724 1343
rect 53760 -24 53772 1367
rect 53832 -24 53844 1223
rect 53856 -24 53868 1295
rect 53904 205 53916 1727
rect 53880 -24 53892 191
rect 53928 -24 53940 983
rect 54000 301 54012 1703
rect 54072 1285 54084 1679
rect 54120 1621 54132 1655
rect 53976 -24 53988 287
rect 54048 -24 54060 1271
rect 54072 -24 54084 1127
rect 54096 -24 54108 1607
rect 54144 -24 54156 1271
rect 54168 -24 54180 1607
rect 54216 157 54228 1631
rect 54192 -24 54204 143
rect 54240 -24 54252 287
rect 54264 -24 54276 1367
rect 54288 -24 54300 1415
rect 54312 301 54324 1607
rect 54336 1381 54348 1559
rect 54360 1429 54372 1559
rect 54336 -24 54348 1367
rect 54408 685 54420 1535
rect 54552 1045 54564 1511
rect 54384 -24 54396 671
rect 54456 -24 54468 551
rect 54480 -24 54492 863
rect 54528 -24 54540 1031
rect 54576 -24 54588 863
rect 54600 -24 54612 527
rect 54672 445 54684 1487
rect 54792 1333 54804 1463
rect 54648 -24 54660 431
rect 54696 -24 54708 1295
rect 54720 -24 54732 959
rect 54768 -24 54780 1319
rect 54816 -24 54828 623
rect 54840 -24 54852 1199
rect 54888 613 54900 1439
rect 54864 -24 54876 599
rect 54912 -24 54924 623
rect 54936 -24 54948 239
rect 54984 181 54996 1415
rect 55080 1189 55092 1391
rect 55176 1261 55188 1367
rect 54960 -24 54972 167
rect 55008 -24 55020 47
rect 55032 -24 55044 959
rect 55056 -24 55068 1175
rect 55104 -24 55116 167
rect 55152 -24 55164 1247
rect 55224 -24 55236 551
rect 55248 -24 55260 527
rect 55296 349 55308 1343
rect 55416 853 55428 1319
rect 55536 1021 55548 1295
rect 55272 -24 55284 335
rect 55320 -24 55332 527
rect 55344 -24 55356 47
rect 55392 -24 55404 839
rect 55440 -24 55452 935
rect 55464 -24 55476 623
rect 55512 -24 55524 1007
rect 55632 829 55644 1271
rect 55560 -24 55572 671
rect 55608 -24 55620 815
rect 55680 -24 55692 1223
rect 55752 1117 55764 1247
rect 55704 -24 55716 719
rect 55728 -24 55740 1103
rect 55776 -24 55788 407
rect 55800 -24 55812 959
rect 55848 85 55860 1223
rect 55824 -24 55836 71
rect 55872 -24 55884 623
rect 55896 -24 55908 959
rect 55920 -24 55932 1175
rect 56040 -24 56052 1199
rect 56472 709 56484 1199
rect 56448 -24 56460 695
rect 56640 589 56652 1175
rect 56592 -24 56604 287
rect 56616 -24 56628 575
rect 56640 -24 56652 143
rect 56688 133 56700 1151
rect 56664 -24 56676 119
rect 56712 -24 56724 887
rect 56784 517 56796 1127
rect 56736 -24 56748 143
rect 56760 -24 56772 503
rect 56880 469 56892 1103
rect 56808 -24 56820 191
rect 56832 -24 56844 143
rect 56856 -24 56868 455
rect 56904 -24 56916 911
rect 56976 229 56988 1079
rect 57096 805 57108 1055
rect 56952 -24 56964 215
rect 57024 -24 57036 47
rect 57048 -24 57060 719
rect 57072 -24 57084 791
rect 57120 -24 57132 935
rect 57168 541 57180 1031
rect 57144 -24 57156 527
rect 57192 397 57204 1007
rect 57168 -24 57180 383
rect 57216 -24 57228 767
rect 57288 757 57300 983
rect 57360 781 57372 959
rect 57240 -24 57252 407
rect 57264 -24 57276 743
rect 57336 565 57348 767
rect 57312 -24 57324 551
rect 57336 -24 57348 551
rect 57384 373 57396 935
rect 57360 -24 57372 359
rect 57408 -24 57420 719
rect 57480 685 57492 911
rect 57432 -24 57444 575
rect 57456 -24 57468 671
rect 57600 541 57612 887
rect 57504 -24 57516 95
rect 57528 -24 57540 503
rect 57576 -24 57588 527
rect 57624 -24 57636 551
rect 57648 -24 57660 863
rect 57696 757 57708 863
rect 57816 805 57828 839
rect 57672 -24 57684 743
rect 57720 -24 57732 143
rect 57744 -24 57756 287
rect 57792 -24 57804 791
rect 57840 -24 57852 95
rect 57864 -24 57876 503
rect 57888 109 57900 815
rect 57912 517 57924 791
rect 57936 133 57948 767
rect 57912 -24 57924 119
rect 57960 -24 57972 719
rect 57984 -24 57996 119
rect 58032 37 58044 743
rect 58008 -24 58020 -1
rect 58056 -24 58068 575
rect 58080 -24 58092 599
rect 58128 181 58140 719
rect 58104 -24 58116 167
rect 58152 -24 58164 167
rect 58176 -24 58188 479
rect 58200 -24 58212 671
rect 58248 -24 58260 599
rect 58272 -24 58284 287
rect 58320 277 58332 671
rect 58296 -24 58308 263
rect 58344 -24 58356 551
rect 58392 37 58404 647
rect 58440 469 58452 623
rect 58368 -24 58380 -1
rect 58416 -24 58428 455
rect 58464 -24 58476 479
rect 58488 -24 58500 167
rect 58560 37 58572 599
rect 58536 -24 58548 -1
rect 58584 -24 58596 479
rect 58608 -24 58620 575
rect 58656 349 58668 575
rect 58632 -24 58644 335
rect 58680 -24 58692 359
rect 58704 -24 58716 551
rect 58728 373 58740 527
rect 58776 229 58788 503
rect 58752 -24 58764 215
rect 58824 37 58836 479
rect 58872 205 58884 455
rect 58944 301 58956 431
rect 58992 373 59004 407
rect 58800 -24 58812 -1
rect 58848 -24 58860 191
rect 58920 -24 58932 287
rect 58968 -24 58980 359
rect 59064 301 59076 383
rect 59112 325 59124 359
rect 59040 -24 59052 287
rect 59088 -24 59100 311
rect 59160 -24 59172 335
rect 59208 -24 59220 311
rect 59304 253 59316 287
rect 59280 -24 59292 239
rect 59352 61 59364 263
rect 59328 -24 59340 47
rect 59424 37 59436 239
rect 59400 -24 59412 -1
rect 59448 -24 59460 191
rect 59544 133 59556 191
rect 59520 -24 59532 119
rect 59592 85 59604 167
rect 59568 -24 59580 71
rect 59640 -24 59652 143
rect 59688 -24 59700 95
rect 59760 -24 59772 95
rect 59808 -24 59820 47
rect 59880 -24 59892 47
rect 59928 -24 59940 -1
use scandtype StatusReg_reg_0
timestamp 1386241841
transform 1 0 24 0 1 -823
box 0 0 624 799
use scandtype StatusReg_reg_1
timestamp 1386241841
transform 1 0 648 0 1 -823
box 0 0 624 799
use scandtype StatusReg_reg_2
timestamp 1386241841
transform 1 0 1272 0 1 -823
box 0 0 624 799
use scandtype StatusReg_reg_3
timestamp 1386241841
transform 1 0 1896 0 1 -823
box 0 0 624 799
use nand2 g11910
timestamp 1386234792
transform 1 0 2520 0 1 -823
box 0 0 96 799
use nand3 g11904
timestamp 1386234893
transform 1 0 2616 0 1 -823
box 0 0 120 799
use nand4 g11889
timestamp 1386234936
transform 1 0 2736 0 1 -823
box 0 0 144 799
use nand4 g11898
timestamp 1386234936
transform 1 0 2880 0 1 -823
box 0 0 144 799
use nand4 g11888
timestamp 1386234936
transform 1 0 3024 0 1 -823
box 0 0 144 799
use nand2 g11922
timestamp 1386234792
transform 1 0 3168 0 1 -823
box 0 0 96 799
use nand2 g11930
timestamp 1386234792
transform 1 0 3264 0 1 -823
box 0 0 96 799
use nand3 g11905
timestamp 1386234893
transform 1 0 3360 0 1 -823
box 0 0 120 799
use scandtype stateSub_reg_0
timestamp 1386241841
transform 1 0 3480 0 1 -823
box 0 0 624 799
use scandtype InISR_reg
timestamp 1386241841
transform 1 0 4104 0 1 -823
box 0 0 624 799
use nand3 g11909
timestamp 1386234893
transform 1 0 4728 0 1 -823
box 0 0 120 799
use nand4 g11925
timestamp 1386234936
transform 1 0 4848 0 1 -823
box 0 0 144 799
use nand3 g11902
timestamp 1386234893
transform 1 0 4992 0 1 -823
box 0 0 120 799
use nand3 g11900
timestamp 1386234893
transform 1 0 5112 0 1 -823
box 0 0 120 799
use nand3 g11903
timestamp 1386234893
transform 1 0 5232 0 1 -823
box 0 0 120 799
use nand2 g11957
timestamp 1386234792
transform 1 0 5352 0 1 -823
box 0 0 96 799
use nand4 g11906
timestamp 1386234936
transform 1 0 5448 0 1 -823
box 0 0 144 799
use nand2 g11921
timestamp 1386234792
transform 1 0 5592 0 1 -823
box 0 0 96 799
use nand4 g11911
timestamp 1386234936
transform 1 0 5688 0 1 -823
box 0 0 144 799
use nor2 g11907
timestamp 1386235306
transform 1 0 5832 0 1 -823
box 0 0 120 799
use nor2 g11931
timestamp 1386235306
transform 1 0 5952 0 1 -823
box 0 0 120 799
use nand2 g11914
timestamp 1386234792
transform 1 0 6072 0 1 -823
box 0 0 96 799
use nand2 g11916
timestamp 1386234792
transform 1 0 6168 0 1 -823
box 0 0 96 799
use and2 g11939
timestamp 1386234845
transform 1 0 6264 0 1 -823
box 0 0 120 799
use nand2 g11915
timestamp 1386234792
transform 1 0 6384 0 1 -823
box 0 0 96 799
use scandtype state_reg_0
timestamp 1386241841
transform 1 0 6480 0 1 -823
box 0 0 624 799
use scandtype state_reg_1
timestamp 1386241841
transform 1 0 7104 0 1 -823
box 0 0 624 799
use nand2 g11913
timestamp 1386234792
transform 1 0 7728 0 1 -823
box 0 0 96 799
use nand4 g11942
timestamp 1386234936
transform 1 0 7824 0 1 -823
box 0 0 144 799
use nand3 g11973
timestamp 1386234893
transform 1 0 7968 0 1 -823
box 0 0 120 799
use nand3 g11947
timestamp 1386234893
transform 1 0 8088 0 1 -823
box 0 0 120 799
use nand2 g11943
timestamp 1386234792
transform 1 0 8208 0 1 -823
box 0 0 96 799
use nor2 g11894
timestamp 1386235306
transform 1 0 8304 0 1 -823
box 0 0 120 799
use nand2 g11945
timestamp 1386234792
transform 1 0 8424 0 1 -823
box 0 0 96 799
use nand4 g11946
timestamp 1386234936
transform 1 0 8520 0 1 -823
box 0 0 144 799
use nand2 g11968
timestamp 1386234792
transform 1 0 8664 0 1 -823
box 0 0 96 799
use nand2 g11926
timestamp 1386234792
transform 1 0 8760 0 1 -823
box 0 0 96 799
use nand2 g11927
timestamp 1386234792
transform 1 0 8856 0 1 -823
box 0 0 96 799
use nand2 g11970
timestamp 1386234792
transform 1 0 8952 0 1 -823
box 0 0 96 799
use nand2 g11928
timestamp 1386234792
transform 1 0 9048 0 1 -823
box 0 0 96 799
use nand2 g11971
timestamp 1386234792
transform 1 0 9144 0 1 -823
box 0 0 96 799
use nand2 g11929
timestamp 1386234792
transform 1 0 9240 0 1 -823
box 0 0 96 799
use nand2 g11972
timestamp 1386234792
transform 1 0 9336 0 1 -823
box 0 0 96 799
use nand3 g11932
timestamp 1386234893
transform 1 0 9432 0 1 -823
box 0 0 120 799
use inv g11992
timestamp 1386238110
transform 1 0 9552 0 1 -823
box 0 0 120 799
use nand4 g11923
timestamp 1386234936
transform 1 0 9672 0 1 -823
box 0 0 144 799
use nand3 g11912
timestamp 1386234893
transform 1 0 9816 0 1 -823
box 0 0 120 799
use nand4 g11901
timestamp 1386234936
transform 1 0 9936 0 1 -823
box 0 0 144 799
use nand2 g11962
timestamp 1386234792
transform 1 0 10080 0 1 -823
box 0 0 96 799
use inv g11952
timestamp 1386238110
transform 1 0 10176 0 1 -823
box 0 0 120 799
use nor2 g11955
timestamp 1386235306
transform 1 0 10296 0 1 -823
box 0 0 120 799
use nand2 g11967
timestamp 1386234792
transform 1 0 10416 0 1 -823
box 0 0 96 799
use inv g11976
timestamp 1386238110
transform 1 0 10512 0 1 -823
box 0 0 120 799
use nand4 g11908
timestamp 1386234936
transform 1 0 10632 0 1 -823
box 0 0 144 799
use nand4 g11896
timestamp 1386234936
transform 1 0 10776 0 1 -823
box 0 0 144 799
use nand3 g11993
timestamp 1386234893
transform 1 0 10920 0 1 -823
box 0 0 120 799
use nand4 g11917
timestamp 1386234936
transform 1 0 11040 0 1 -823
box 0 0 144 799
use nand2 g11941
timestamp 1386234792
transform 1 0 11184 0 1 -823
box 0 0 96 799
use nand4 g11948
timestamp 1386234936
transform 1 0 11280 0 1 -823
box 0 0 144 799
use nand2 g11964
timestamp 1386234792
transform 1 0 11424 0 1 -823
box 0 0 96 799
use nand4 g11899
timestamp 1386234936
transform 1 0 11520 0 1 -823
box 0 0 144 799
use nand4 g11974
timestamp 1386234936
transform 1 0 11664 0 1 -823
box 0 0 144 799
use nand4 g11897
timestamp 1386234936
transform 1 0 11808 0 1 -823
box 0 0 144 799
use nand4 g11951
timestamp 1386234936
transform 1 0 11952 0 1 -823
box 0 0 144 799
use nand4 g11953
timestamp 1386234936
transform 1 0 12096 0 1 -823
box 0 0 144 799
use nand2 g11954
timestamp 1386234792
transform 1 0 12240 0 1 -823
box 0 0 96 799
use and2 g11958
timestamp 1386234845
transform 1 0 12336 0 1 -823
box 0 0 120 799
use nand2 g11963
timestamp 1386234792
transform 1 0 12456 0 1 -823
box 0 0 96 799
use nand4 g11977
timestamp 1386234936
transform 1 0 12552 0 1 -823
box 0 0 144 799
use nand2 g11983
timestamp 1386234792
transform 1 0 12696 0 1 -823
box 0 0 96 799
use nand2 g11984
timestamp 1386234792
transform 1 0 12792 0 1 -823
box 0 0 96 799
use inv g11985
timestamp 1386238110
transform 1 0 12888 0 1 -823
box 0 0 120 799
use and2 g11988
timestamp 1386234845
transform 1 0 13008 0 1 -823
box 0 0 120 799
use nand2 g11990
timestamp 1386234792
transform 1 0 13128 0 1 -823
box 0 0 96 799
use inv g11995
timestamp 1386238110
transform 1 0 13224 0 1 -823
box 0 0 120 799
use nand2 g11960
timestamp 1386234792
transform 1 0 13344 0 1 -823
box 0 0 96 799
use nand3 g11944
timestamp 1386234893
transform 1 0 13440 0 1 -823
box 0 0 120 799
use and2 g12002
timestamp 1386234845
transform 1 0 13560 0 1 -823
box 0 0 120 799
use inv g12006
timestamp 1386238110
transform 1 0 13680 0 1 -823
box 0 0 120 799
use trisbuf g746
timestamp 1386237216
transform 1 0 13800 0 1 -823
box 0 0 216 799
use trisbuf g738
timestamp 1386237216
transform 1 0 14016 0 1 -823
box 0 0 216 799
use and2 g11981
timestamp 1386234845
transform 1 0 14232 0 1 -823
box 0 0 120 799
use nand2 g11986
timestamp 1386234792
transform 1 0 14352 0 1 -823
box 0 0 96 799
use nand2 g11987
timestamp 1386234792
transform 1 0 14448 0 1 -823
box 0 0 96 799
use nand2 g11937
timestamp 1386234792
transform 1 0 14544 0 1 -823
box 0 0 96 799
use nand2 g11991
timestamp 1386234792
transform 1 0 14640 0 1 -823
box 0 0 96 799
use nand2 g11938
timestamp 1386234792
transform 1 0 14736 0 1 -823
box 0 0 96 799
use nand2 g11996
timestamp 1386234792
transform 1 0 14832 0 1 -823
box 0 0 96 799
use nand2 g11940
timestamp 1386234792
transform 1 0 14928 0 1 -823
box 0 0 96 799
use nand3 g11999
timestamp 1386234893
transform 1 0 15024 0 1 -823
box 0 0 120 799
use trisbuf g742
timestamp 1386237216
transform 1 0 15144 0 1 -823
box 0 0 216 799
use nand3 g12000
timestamp 1386234893
transform 1 0 15360 0 1 -823
box 0 0 120 799
use trisbuf g1
timestamp 1386237216
transform 1 0 15480 0 1 -823
box 0 0 216 799
use trisbuf g734
timestamp 1386237216
transform 1 0 15696 0 1 -823
box 0 0 216 799
use trisbuf g735
timestamp 1386237216
transform 1 0 15912 0 1 -823
box 0 0 216 799
use trisbuf g736
timestamp 1386237216
transform 1 0 16128 0 1 -823
box 0 0 216 799
use trisbuf g737
timestamp 1386237216
transform 1 0 16344 0 1 -823
box 0 0 216 799
use trisbuf g739
timestamp 1386237216
transform 1 0 16560 0 1 -823
box 0 0 216 799
use trisbuf g740
timestamp 1386237216
transform 1 0 16776 0 1 -823
box 0 0 216 799
use trisbuf g741
timestamp 1386237216
transform 1 0 16992 0 1 -823
box 0 0 216 799
use trisbuf g743
timestamp 1386237216
transform 1 0 17208 0 1 -823
box 0 0 216 799
use trisbuf g744
timestamp 1386237216
transform 1 0 17424 0 1 -823
box 0 0 216 799
use trisbuf g745
timestamp 1386237216
transform 1 0 17640 0 1 -823
box 0 0 216 799
use trisbuf g747
timestamp 1386237216
transform 1 0 17856 0 1 -823
box 0 0 216 799
use trisbuf g748
timestamp 1386237216
transform 1 0 18072 0 1 -823
box 0 0 216 799
use nand3 g12004
timestamp 1386234893
transform 1 0 18288 0 1 -823
box 0 0 120 799
use nand3 g12007
timestamp 1386234893
transform 1 0 18408 0 1 -823
box 0 0 120 799
use nand2 g11961
timestamp 1386234792
transform 1 0 18528 0 1 -823
box 0 0 96 799
use nor2 g11924
timestamp 1386235306
transform 1 0 18624 0 1 -823
box 0 0 120 799
use nand2 g12035
timestamp 1386234792
transform 1 0 18744 0 1 -823
box 0 0 96 799
use nand2 g12036
timestamp 1386234792
transform 1 0 18840 0 1 -823
box 0 0 96 799
use and2 g11969
timestamp 1386234845
transform 1 0 18936 0 1 -823
box 0 0 120 799
use nand2 g11997
timestamp 1386234792
transform 1 0 19056 0 1 -823
box 0 0 96 799
use nand2 g12043
timestamp 1386234792
transform 1 0 19152 0 1 -823
box 0 0 96 799
use nor2 g11933
timestamp 1386235306
transform 1 0 19248 0 1 -823
box 0 0 120 799
use nor2 g11982
timestamp 1386235306
transform 1 0 19368 0 1 -823
box 0 0 120 799
use inv g11935
timestamp 1386238110
transform 1 0 19488 0 1 -823
box 0 0 120 799
use and2 g11994
timestamp 1386234845
transform 1 0 19608 0 1 -823
box 0 0 120 799
use scandtype stateSub_reg_2
timestamp 1386241841
transform 1 0 19728 0 1 -823
box 0 0 624 799
use nand2 g12020
timestamp 1386234792
transform 1 0 20352 0 1 -823
box 0 0 96 799
use nand3 g12005
timestamp 1386234893
transform 1 0 20448 0 1 -823
box 0 0 120 799
use inv g11949
timestamp 1386238110
transform 1 0 20568 0 1 -823
box 0 0 120 799
use nand2 g12014
timestamp 1386234792
transform 1 0 20688 0 1 -823
box 0 0 96 799
use nand2 g12015
timestamp 1386234792
transform 1 0 20784 0 1 -823
box 0 0 96 799
use nand2 g12017
timestamp 1386234792
transform 1 0 20880 0 1 -823
box 0 0 96 799
use nand2 g12018
timestamp 1386234792
transform 1 0 20976 0 1 -823
box 0 0 96 799
use nand2 g12022
timestamp 1386234792
transform 1 0 21072 0 1 -823
box 0 0 96 799
use nand2 g12025
timestamp 1386234792
transform 1 0 21168 0 1 -823
box 0 0 96 799
use nand2 g12027
timestamp 1386234792
transform 1 0 21264 0 1 -823
box 0 0 96 799
use nand2 g12028
timestamp 1386234792
transform 1 0 21360 0 1 -823
box 0 0 96 799
use nand2 g12030
timestamp 1386234792
transform 1 0 21456 0 1 -823
box 0 0 96 799
use nand4 g11966
timestamp 1386234936
transform 1 0 21552 0 1 -823
box 0 0 144 799
use nand3 g12032
timestamp 1386234893
transform 1 0 21696 0 1 -823
box 0 0 120 799
use and2 g12038
timestamp 1386234845
transform 1 0 21816 0 1 -823
box 0 0 120 799
use and2 g12040
timestamp 1386234845
transform 1 0 21936 0 1 -823
box 0 0 120 799
use inv g12044
timestamp 1386238110
transform 1 0 22056 0 1 -823
box 0 0 120 799
use nand4 g11936
timestamp 1386234936
transform 1 0 22176 0 1 -823
box 0 0 144 799
use nand2 g11989
timestamp 1386234792
transform 1 0 22320 0 1 -823
box 0 0 96 799
use nand4 g11998
timestamp 1386234936
transform 1 0 22416 0 1 -823
box 0 0 144 799
use inv g12008
timestamp 1386238110
transform 1 0 22560 0 1 -823
box 0 0 120 799
use nand2 g12010
timestamp 1386234792
transform 1 0 22680 0 1 -823
box 0 0 96 799
use nand4 g11950
timestamp 1386234936
transform 1 0 22776 0 1 -823
box 0 0 144 799
use nand2 g12013
timestamp 1386234792
transform 1 0 22920 0 1 -823
box 0 0 96 799
use nand2 g12019
timestamp 1386234792
transform 1 0 23016 0 1 -823
box 0 0 96 799
use nand4 g11965
timestamp 1386234936
transform 1 0 23112 0 1 -823
box 0 0 144 799
use nand4 g11959
timestamp 1386234936
transform 1 0 23256 0 1 -823
box 0 0 144 799
use inv g12100
timestamp 1386238110
transform 1 0 23400 0 1 -823
box 0 0 120 799
use nand3 g12033
timestamp 1386234893
transform 1 0 23520 0 1 -823
box 0 0 120 799
use nand3 g12037
timestamp 1386234893
transform 1 0 23640 0 1 -823
box 0 0 120 799
use nand3 g12042
timestamp 1386234893
transform 1 0 23760 0 1 -823
box 0 0 120 799
use nand3 g12045
timestamp 1386234893
transform 1 0 23880 0 1 -823
box 0 0 120 799
use nand3 g12046
timestamp 1386234893
transform 1 0 24000 0 1 -823
box 0 0 120 799
use nand3 g12047
timestamp 1386234893
transform 1 0 24120 0 1 -823
box 0 0 120 799
use nand3 g12048
timestamp 1386234893
transform 1 0 24240 0 1 -823
box 0 0 120 799
use nand3 g12049
timestamp 1386234893
transform 1 0 24360 0 1 -823
box 0 0 120 799
use nand4 g11934
timestamp 1386234936
transform 1 0 24480 0 1 -823
box 0 0 144 799
use inv g12062
timestamp 1386238110
transform 1 0 24624 0 1 -823
box 0 0 120 799
use nand2 g12068
timestamp 1386234792
transform 1 0 24744 0 1 -823
box 0 0 96 799
use and2 g12069
timestamp 1386234845
transform 1 0 24840 0 1 -823
box 0 0 120 799
use nand2 g12070
timestamp 1386234792
transform 1 0 24960 0 1 -823
box 0 0 96 799
use nand2 g12073
timestamp 1386234792
transform 1 0 25056 0 1 -823
box 0 0 96 799
use nand2 g12080
timestamp 1386234792
transform 1 0 25152 0 1 -823
box 0 0 96 799
use and2 g12085
timestamp 1386234845
transform 1 0 25248 0 1 -823
box 0 0 120 799
use nand2 g12087
timestamp 1386234792
transform 1 0 25368 0 1 -823
box 0 0 96 799
use nand2 g12088
timestamp 1386234792
transform 1 0 25464 0 1 -823
box 0 0 96 799
use scandtype stateSub_reg_1
timestamp 1386241841
transform 1 0 25560 0 1 -823
box 0 0 624 799
use nand2 g12090
timestamp 1386234792
transform 1 0 26184 0 1 -823
box 0 0 96 799
use nand2 g12001
timestamp 1386234792
transform 1 0 26280 0 1 -823
box 0 0 96 799
use nand4 g12009
timestamp 1386234936
transform 1 0 26376 0 1 -823
box 0 0 144 799
use nand2 g12091
timestamp 1386234792
transform 1 0 26520 0 1 -823
box 0 0 96 799
use and2 g12012
timestamp 1386234845
transform 1 0 26616 0 1 -823
box 0 0 120 799
use nand3 g12021
timestamp 1386234893
transform 1 0 26736 0 1 -823
box 0 0 120 799
use and2 g11956
timestamp 1386234845
transform 1 0 26856 0 1 -823
box 0 0 120 799
use nand3 g12024
timestamp 1386234893
transform 1 0 26976 0 1 -823
box 0 0 120 799
use nand3 g12029
timestamp 1386234893
transform 1 0 27096 0 1 -823
box 0 0 120 799
use nand2 g12031
timestamp 1386234792
transform 1 0 27216 0 1 -823
box 0 0 96 799
use nand3 g12099
timestamp 1386234893
transform 1 0 27312 0 1 -823
box 0 0 120 799
use nand2 g12041
timestamp 1386234792
transform 1 0 27432 0 1 -823
box 0 0 96 799
use nand4 g11975
timestamp 1386234936
transform 1 0 27528 0 1 -823
box 0 0 144 799
use nand2 g12098
timestamp 1386234792
transform 1 0 27672 0 1 -823
box 0 0 96 799
use nand2 g12063
timestamp 1386234792
transform 1 0 27768 0 1 -823
box 0 0 96 799
use nand2 g12065
timestamp 1386234792
transform 1 0 27864 0 1 -823
box 0 0 96 799
use nand2 g12066
timestamp 1386234792
transform 1 0 27960 0 1 -823
box 0 0 96 799
use nand2 g12067
timestamp 1386234792
transform 1 0 28056 0 1 -823
box 0 0 96 799
use and2 g12097
timestamp 1386234845
transform 1 0 28152 0 1 -823
box 0 0 120 799
use nand2 g12074
timestamp 1386234792
transform 1 0 28272 0 1 -823
box 0 0 96 799
use nand2 g12075
timestamp 1386234792
transform 1 0 28368 0 1 -823
box 0 0 96 799
use nand2 g12076
timestamp 1386234792
transform 1 0 28464 0 1 -823
box 0 0 96 799
use nand2 g12077
timestamp 1386234792
transform 1 0 28560 0 1 -823
box 0 0 96 799
use nand2 g12078
timestamp 1386234792
transform 1 0 28656 0 1 -823
box 0 0 96 799
use nand2 g12081
timestamp 1386234792
transform 1 0 28752 0 1 -823
box 0 0 96 799
use nand2 g12082
timestamp 1386234792
transform 1 0 28848 0 1 -823
box 0 0 96 799
use nand2 g12084
timestamp 1386234792
transform 1 0 28944 0 1 -823
box 0 0 96 799
use nand2 g12086
timestamp 1386234792
transform 1 0 29040 0 1 -823
box 0 0 96 799
use nand3 g12101
timestamp 1386234893
transform 1 0 29136 0 1 -823
box 0 0 120 799
use nand2 g12089
timestamp 1386234792
transform 1 0 29256 0 1 -823
box 0 0 96 799
use scandtype IntReq_reg
timestamp 1386241841
transform 1 0 29352 0 1 -823
box 0 0 624 799
use and2 g12092
timestamp 1386234845
transform 1 0 29976 0 1 -823
box 0 0 120 799
use nand2 g12096
timestamp 1386234792
transform 1 0 30096 0 1 -823
box 0 0 96 799
use nand3 g12053
timestamp 1386234893
transform 1 0 30192 0 1 -823
box 0 0 120 799
use inv g12054
timestamp 1386238110
transform 1 0 30312 0 1 -823
box 0 0 120 799
use nor2 g12056
timestamp 1386235306
transform 1 0 30432 0 1 -823
box 0 0 120 799
use nor2 g12058
timestamp 1386235306
transform 1 0 30552 0 1 -823
box 0 0 120 799
use nand3 g12003
timestamp 1386234893
transform 1 0 30672 0 1 -823
box 0 0 120 799
use nand3 g12105
timestamp 1386234893
transform 1 0 30792 0 1 -823
box 0 0 120 799
use and2 g12120
timestamp 1386234845
transform 1 0 30912 0 1 -823
box 0 0 120 799
use and2 g12121
timestamp 1386234845
transform 1 0 31032 0 1 -823
box 0 0 120 799
use nand3 g12011
timestamp 1386234893
transform 1 0 31152 0 1 -823
box 0 0 120 799
use and2 g12130
timestamp 1386234845
transform 1 0 31272 0 1 -823
box 0 0 120 799
use nand3 g12016
timestamp 1386234893
transform 1 0 31392 0 1 -823
box 0 0 120 799
use nand2 g12139
timestamp 1386234792
transform 1 0 31512 0 1 -823
box 0 0 96 799
use nand3 g12023
timestamp 1386234893
transform 1 0 31608 0 1 -823
box 0 0 120 799
use nand2 g12026
timestamp 1386234792
transform 1 0 31728 0 1 -823
box 0 0 96 799
use nand2 g12034
timestamp 1386234792
transform 1 0 31824 0 1 -823
box 0 0 96 799
use nand3 g12039
timestamp 1386234893
transform 1 0 31920 0 1 -823
box 0 0 120 799
use nand2 g12094
timestamp 1386234792
transform 1 0 32040 0 1 -823
box 0 0 96 799
use inv g12051
timestamp 1386238110
transform 1 0 32136 0 1 -823
box 0 0 120 799
use nand4 g12055
timestamp 1386234936
transform 1 0 32256 0 1 -823
box 0 0 144 799
use nor2 g12057
timestamp 1386235306
transform 1 0 32400 0 1 -823
box 0 0 120 799
use nand2 g12060
timestamp 1386234792
transform 1 0 32520 0 1 -823
box 0 0 96 799
use nand2 g12061
timestamp 1386234792
transform 1 0 32616 0 1 -823
box 0 0 96 799
use nand2 g12064
timestamp 1386234792
transform 1 0 32712 0 1 -823
box 0 0 96 799
use nand3 g12083
timestamp 1386234893
transform 1 0 32808 0 1 -823
box 0 0 120 799
use nand3 g12102
timestamp 1386234893
transform 1 0 32928 0 1 -823
box 0 0 120 799
use inv g12103
timestamp 1386238110
transform 1 0 33048 0 1 -823
box 0 0 120 799
use nand3 g12106
timestamp 1386234893
transform 1 0 33168 0 1 -823
box 0 0 120 799
use and2 g12117
timestamp 1386234845
transform 1 0 33288 0 1 -823
box 0 0 120 799
use nand2 g12118
timestamp 1386234792
transform 1 0 33408 0 1 -823
box 0 0 96 799
use nand2 g12123
timestamp 1386234792
transform 1 0 33504 0 1 -823
box 0 0 96 799
use inv g12124
timestamp 1386238110
transform 1 0 33600 0 1 -823
box 0 0 120 799
use nand2 g12128
timestamp 1386234792
transform 1 0 33720 0 1 -823
box 0 0 96 799
use and2 g12129
timestamp 1386234845
transform 1 0 33816 0 1 -823
box 0 0 120 799
use nand2 g12132
timestamp 1386234792
transform 1 0 33936 0 1 -823
box 0 0 96 799
use nand2 g12135
timestamp 1386234792
transform 1 0 34032 0 1 -823
box 0 0 96 799
use nand2 g12136
timestamp 1386234792
transform 1 0 34128 0 1 -823
box 0 0 96 799
use and2 g12138
timestamp 1386234845
transform 1 0 34224 0 1 -823
box 0 0 120 799
use nand2 g12143
timestamp 1386234792
transform 1 0 34344 0 1 -823
box 0 0 96 799
use nand2 g12147
timestamp 1386234792
transform 1 0 34440 0 1 -823
box 0 0 96 799
use inv g12179
timestamp 1386238110
transform 1 0 34536 0 1 -823
box 0 0 120 799
use nand4 g12052
timestamp 1386234936
transform 1 0 34656 0 1 -823
box 0 0 144 799
use nand2 g12059
timestamp 1386234792
transform 1 0 34800 0 1 -823
box 0 0 96 799
use nand2 g12071
timestamp 1386234792
transform 1 0 34896 0 1 -823
box 0 0 96 799
use nand2 g12072
timestamp 1386234792
transform 1 0 34992 0 1 -823
box 0 0 96 799
use and2 g12079
timestamp 1386234845
transform 1 0 35088 0 1 -823
box 0 0 120 799
use and2 g12095
timestamp 1386234845
transform 1 0 35208 0 1 -823
box 0 0 120 799
use nand3 g12104
timestamp 1386234893
transform 1 0 35328 0 1 -823
box 0 0 120 799
use nor2 g12107
timestamp 1386235306
transform 1 0 35448 0 1 -823
box 0 0 120 799
use nand2 g12113
timestamp 1386234792
transform 1 0 35568 0 1 -823
box 0 0 96 799
use nand2 g12115
timestamp 1386234792
transform 1 0 35664 0 1 -823
box 0 0 96 799
use nand2 g12119
timestamp 1386234792
transform 1 0 35760 0 1 -823
box 0 0 96 799
use nand2 g12125
timestamp 1386234792
transform 1 0 35856 0 1 -823
box 0 0 96 799
use nand2 g12126
timestamp 1386234792
transform 1 0 35952 0 1 -823
box 0 0 96 799
use inv g12174
timestamp 1386238110
transform 1 0 36048 0 1 -823
box 0 0 120 799
use nand2 g12180
timestamp 1386234792
transform 1 0 36168 0 1 -823
box 0 0 96 799
use nand2 g12182
timestamp 1386234792
transform 1 0 36264 0 1 -823
box 0 0 96 799
use nand2 g12183
timestamp 1386234792
transform 1 0 36360 0 1 -823
box 0 0 96 799
use inv g12184
timestamp 1386238110
transform 1 0 36456 0 1 -823
box 0 0 120 799
use inv g12187
timestamp 1386238110
transform 1 0 36576 0 1 -823
box 0 0 120 799
use nand2 g12192
timestamp 1386234792
transform 1 0 36696 0 1 -823
box 0 0 96 799
use nand2 g12194
timestamp 1386234792
transform 1 0 36792 0 1 -823
box 0 0 96 799
use nand4 g12050
timestamp 1386234936
transform 1 0 36888 0 1 -823
box 0 0 144 799
use nand2 g12093
timestamp 1386234792
transform 1 0 37032 0 1 -823
box 0 0 96 799
use nand2 g12108
timestamp 1386234792
transform 1 0 37128 0 1 -823
box 0 0 96 799
use nor2 g12110
timestamp 1386235306
transform 1 0 37224 0 1 -823
box 0 0 120 799
use nor2 g12111
timestamp 1386235306
transform 1 0 37344 0 1 -823
box 0 0 120 799
use nor2 g12112
timestamp 1386235306
transform 1 0 37464 0 1 -823
box 0 0 120 799
use nand2 g12114
timestamp 1386234792
transform 1 0 37584 0 1 -823
box 0 0 96 799
use nand2 g12134
timestamp 1386234792
transform 1 0 37680 0 1 -823
box 0 0 96 799
use nand2 g12141
timestamp 1386234792
transform 1 0 37776 0 1 -823
box 0 0 96 799
use nand2 g12144
timestamp 1386234792
transform 1 0 37872 0 1 -823
box 0 0 96 799
use nand3 g12146
timestamp 1386234893
transform 1 0 37968 0 1 -823
box 0 0 120 799
use inv g12148
timestamp 1386238110
transform 1 0 38088 0 1 -823
box 0 0 120 799
use nand2 g12161
timestamp 1386234792
transform 1 0 38208 0 1 -823
box 0 0 96 799
use and2 g12162
timestamp 1386234845
transform 1 0 38304 0 1 -823
box 0 0 120 799
use inv g12163
timestamp 1386238110
transform 1 0 38424 0 1 -823
box 0 0 120 799
use and2 g12165
timestamp 1386234845
transform 1 0 38544 0 1 -823
box 0 0 120 799
use nand2 g12173
timestamp 1386234792
transform 1 0 38664 0 1 -823
box 0 0 96 799
use nand2 g12175
timestamp 1386234792
transform 1 0 38760 0 1 -823
box 0 0 96 799
use nand2 g12181
timestamp 1386234792
transform 1 0 38856 0 1 -823
box 0 0 96 799
use nand2 g12185
timestamp 1386234792
transform 1 0 38952 0 1 -823
box 0 0 96 799
use nor2 g12188
timestamp 1386235306
transform 1 0 39048 0 1 -823
box 0 0 120 799
use nand2 g12191
timestamp 1386234792
transform 1 0 39168 0 1 -823
box 0 0 96 799
use nand2 g12199
timestamp 1386234792
transform 1 0 39264 0 1 -823
box 0 0 96 799
use nand2 g12201
timestamp 1386234792
transform 1 0 39360 0 1 -823
box 0 0 96 799
use nand2 g12202
timestamp 1386234792
transform 1 0 39456 0 1 -823
box 0 0 96 799
use nand2 g12203
timestamp 1386234792
transform 1 0 39552 0 1 -823
box 0 0 96 799
use nor2 g12109
timestamp 1386235306
transform 1 0 39648 0 1 -823
box 0 0 120 799
use nand2 g12116
timestamp 1386234792
transform 1 0 39768 0 1 -823
box 0 0 96 799
use nand2 g12122
timestamp 1386234792
transform 1 0 39864 0 1 -823
box 0 0 96 799
use nand2 g12131
timestamp 1386234792
transform 1 0 39960 0 1 -823
box 0 0 96 799
use nand2 g12137
timestamp 1386234792
transform 1 0 40056 0 1 -823
box 0 0 96 799
use nand2 g12140
timestamp 1386234792
transform 1 0 40152 0 1 -823
box 0 0 96 799
use nand2 g12142
timestamp 1386234792
transform 1 0 40248 0 1 -823
box 0 0 96 799
use nand2 g12145
timestamp 1386234792
transform 1 0 40344 0 1 -823
box 0 0 96 799
use nand3 g12149
timestamp 1386234893
transform 1 0 40440 0 1 -823
box 0 0 120 799
use nand2 g12153
timestamp 1386234792
transform 1 0 40560 0 1 -823
box 0 0 96 799
use nor2 g12155
timestamp 1386235306
transform 1 0 40656 0 1 -823
box 0 0 120 799
use nand2 g12160
timestamp 1386234792
transform 1 0 40776 0 1 -823
box 0 0 96 799
use nor2 g12164
timestamp 1386235306
transform 1 0 40872 0 1 -823
box 0 0 120 799
use nand2 g12166
timestamp 1386234792
transform 1 0 40992 0 1 -823
box 0 0 96 799
use inv g12167
timestamp 1386238110
transform 1 0 41088 0 1 -823
box 0 0 120 799
use nand2 g12169
timestamp 1386234792
transform 1 0 41208 0 1 -823
box 0 0 96 799
use nand2 g12178
timestamp 1386234792
transform 1 0 41304 0 1 -823
box 0 0 96 799
use inv g12254
timestamp 1386238110
transform 1 0 41400 0 1 -823
box 0 0 120 799
use nand2 g12190
timestamp 1386234792
transform 1 0 41520 0 1 -823
box 0 0 96 799
use nand2 g12195
timestamp 1386234792
transform 1 0 41616 0 1 -823
box 0 0 96 799
use nand2 g12196
timestamp 1386234792
transform 1 0 41712 0 1 -823
box 0 0 96 799
use nand2 g12197
timestamp 1386234792
transform 1 0 41808 0 1 -823
box 0 0 96 799
use nand2 g12200
timestamp 1386234792
transform 1 0 41904 0 1 -823
box 0 0 96 799
use nor2 g12206
timestamp 1386235306
transform 1 0 42000 0 1 -823
box 0 0 120 799
use inv g12222
timestamp 1386238110
transform 1 0 42120 0 1 -823
box 0 0 120 799
use inv g12227
timestamp 1386238110
transform 1 0 42240 0 1 -823
box 0 0 120 799
use inv g12243
timestamp 1386238110
transform 1 0 42360 0 1 -823
box 0 0 120 799
use nand3 g12256
timestamp 1386234893
transform 1 0 42480 0 1 -823
box 0 0 120 799
use inv g12258
timestamp 1386238110
transform 1 0 42600 0 1 -823
box 0 0 120 799
use inv g12261
timestamp 1386238110
transform 1 0 42720 0 1 -823
box 0 0 120 799
use nand2 g12189
timestamp 1386234792
transform 1 0 42840 0 1 -823
box 0 0 96 799
use and2 g12186
timestamp 1386234845
transform 1 0 42936 0 1 -823
box 0 0 120 799
use inv g12170
timestamp 1386238110
transform 1 0 43056 0 1 -823
box 0 0 120 799
use nand2 g12168
timestamp 1386234792
transform 1 0 43176 0 1 -823
box 0 0 96 799
use nand2 g12133
timestamp 1386234792
transform 1 0 43272 0 1 -823
box 0 0 96 799
use nand2 g12150
timestamp 1386234792
transform 1 0 43368 0 1 -823
box 0 0 96 799
use nand2 g12151
timestamp 1386234792
transform 1 0 43464 0 1 -823
box 0 0 96 799
use nand2 g12154
timestamp 1386234792
transform 1 0 43560 0 1 -823
box 0 0 96 799
use inv g12176
timestamp 1386238110
transform 1 0 43656 0 1 -823
box 0 0 120 799
use nand2 g12177
timestamp 1386234792
transform 1 0 43776 0 1 -823
box 0 0 96 799
use nand2 g12193
timestamp 1386234792
transform 1 0 43872 0 1 -823
box 0 0 96 799
use nand2 g12204
timestamp 1386234792
transform 1 0 43968 0 1 -823
box 0 0 96 799
use nand3 g12205
timestamp 1386234893
transform 1 0 44064 0 1 -823
box 0 0 120 799
use mux2 g12207
timestamp 1386235218
transform 1 0 44184 0 1 -823
box 0 0 192 799
use nand2 g12213
timestamp 1386234792
transform 1 0 44376 0 1 -823
box 0 0 96 799
use inv g12215
timestamp 1386238110
transform 1 0 44472 0 1 -823
box 0 0 120 799
use nor2 g12218
timestamp 1386235306
transform 1 0 44592 0 1 -823
box 0 0 120 799
use nand2 g12221
timestamp 1386234792
transform 1 0 44712 0 1 -823
box 0 0 96 799
use nand2 g12223
timestamp 1386234792
transform 1 0 44808 0 1 -823
box 0 0 96 799
use nand2 g12226
timestamp 1386234792
transform 1 0 44904 0 1 -823
box 0 0 96 799
use nor2 g12228
timestamp 1386235306
transform 1 0 45000 0 1 -823
box 0 0 120 799
use inv g12231
timestamp 1386238110
transform 1 0 45120 0 1 -823
box 0 0 120 799
use inv g12233
timestamp 1386238110
transform 1 0 45240 0 1 -823
box 0 0 120 799
use nand2 g12244
timestamp 1386234792
transform 1 0 45360 0 1 -823
box 0 0 96 799
use nand2 g12248
timestamp 1386234792
transform 1 0 45456 0 1 -823
box 0 0 96 799
use inv g12249
timestamp 1386238110
transform 1 0 45552 0 1 -823
box 0 0 120 799
use nand2 g12251
timestamp 1386234792
transform 1 0 45672 0 1 -823
box 0 0 96 799
use nand2 g12252
timestamp 1386234792
transform 1 0 45768 0 1 -823
box 0 0 96 799
use nand2 g12253
timestamp 1386234792
transform 1 0 45864 0 1 -823
box 0 0 96 799
use nand2 g12255
timestamp 1386234792
transform 1 0 45960 0 1 -823
box 0 0 96 799
use nand2 g12257
timestamp 1386234792
transform 1 0 46056 0 1 -823
box 0 0 96 799
use nand2 g12259
timestamp 1386234792
transform 1 0 46152 0 1 -823
box 0 0 96 799
use and2 g12263
timestamp 1386234845
transform 1 0 46248 0 1 -823
box 0 0 120 799
use nand2 g12269
timestamp 1386234792
transform 1 0 46368 0 1 -823
box 0 0 96 799
use nand2 g12217
timestamp 1386234792
transform 1 0 46464 0 1 -823
box 0 0 96 799
use and2 g12237
timestamp 1386234845
transform 1 0 46560 0 1 -823
box 0 0 120 799
use nand4 g12127
timestamp 1386234936
transform 1 0 46680 0 1 -823
box 0 0 144 799
use nand3 g12152
timestamp 1386234893
transform 1 0 46824 0 1 -823
box 0 0 120 799
use and2 g12156
timestamp 1386234845
transform 1 0 46944 0 1 -823
box 0 0 120 799
use nand2 g12157
timestamp 1386234792
transform 1 0 47064 0 1 -823
box 0 0 96 799
use nand2 g12158
timestamp 1386234792
transform 1 0 47160 0 1 -823
box 0 0 96 799
use nand3 g12159
timestamp 1386234893
transform 1 0 47256 0 1 -823
box 0 0 120 799
use nand2 g12262
timestamp 1386234792
transform 1 0 47376 0 1 -823
box 0 0 96 799
use nand3 g12171
timestamp 1386234893
transform 1 0 47472 0 1 -823
box 0 0 120 799
use nand3 g12172
timestamp 1386234893
transform 1 0 47592 0 1 -823
box 0 0 120 799
use and2 g12266
timestamp 1386234845
transform 1 0 47712 0 1 -823
box 0 0 120 799
use mux2 g12208
timestamp 1386235218
transform 1 0 47832 0 1 -823
box 0 0 192 799
use inv g12270
timestamp 1386238110
transform 1 0 48024 0 1 -823
box 0 0 120 799
use nor2 g12214
timestamp 1386235306
transform 1 0 48144 0 1 -823
box 0 0 120 799
use nor2 g12216
timestamp 1386235306
transform 1 0 48264 0 1 -823
box 0 0 120 799
use nand2 g12220
timestamp 1386234792
transform 1 0 48384 0 1 -823
box 0 0 96 799
use nand2 g12224
timestamp 1386234792
transform 1 0 48480 0 1 -823
box 0 0 96 799
use nand2 g12225
timestamp 1386234792
transform 1 0 48576 0 1 -823
box 0 0 96 799
use nand2 g12229
timestamp 1386234792
transform 1 0 48672 0 1 -823
box 0 0 96 799
use nand2 g12230
timestamp 1386234792
transform 1 0 48768 0 1 -823
box 0 0 96 799
use nand2 g12232
timestamp 1386234792
transform 1 0 48864 0 1 -823
box 0 0 96 799
use nand2 g12234
timestamp 1386234792
transform 1 0 48960 0 1 -823
box 0 0 96 799
use nand2 g12236
timestamp 1386234792
transform 1 0 49056 0 1 -823
box 0 0 96 799
use nand2 g12239
timestamp 1386234792
transform 1 0 49152 0 1 -823
box 0 0 96 799
use nand2 g12240
timestamp 1386234792
transform 1 0 49248 0 1 -823
box 0 0 96 799
use nand2 g12277
timestamp 1386234792
transform 1 0 49344 0 1 -823
box 0 0 96 799
use nand2 g12245
timestamp 1386234792
transform 1 0 49440 0 1 -823
box 0 0 96 799
use nand2 g12246
timestamp 1386234792
transform 1 0 49536 0 1 -823
box 0 0 96 799
use nand2 g12247
timestamp 1386234792
transform 1 0 49632 0 1 -823
box 0 0 96 799
use nor2 g12250
timestamp 1386235306
transform 1 0 49728 0 1 -823
box 0 0 120 799
use and2 g12265
timestamp 1386234845
transform 1 0 49848 0 1 -823
box 0 0 120 799
use nand2 g12268
timestamp 1386234792
transform 1 0 49968 0 1 -823
box 0 0 96 799
use nand2 g12276
timestamp 1386234792
transform 1 0 50064 0 1 -823
box 0 0 96 799
use nand2 g12238
timestamp 1386234792
transform 1 0 50160 0 1 -823
box 0 0 96 799
use nand2 g12212
timestamp 1386234792
transform 1 0 50256 0 1 -823
box 0 0 96 799
use scandtype IRQ2_reg
timestamp 1386241841
transform 1 0 50352 0 1 -823
box 0 0 624 799
use nand2 g12275
timestamp 1386234792
transform 1 0 50976 0 1 -823
box 0 0 96 799
use nand2 g12260
timestamp 1386234792
transform 1 0 51072 0 1 -823
box 0 0 96 799
use nand2 g12209
timestamp 1386234792
transform 1 0 51168 0 1 -823
box 0 0 96 799
use nand3 g12242
timestamp 1386234893
transform 1 0 51264 0 1 -823
box 0 0 120 799
use and2 g12219
timestamp 1386234845
transform 1 0 51384 0 1 -823
box 0 0 120 799
use inv g12284
timestamp 1386238110
transform 1 0 51504 0 1 -823
box 0 0 120 799
use nand2 g12241
timestamp 1386234792
transform 1 0 51624 0 1 -823
box 0 0 96 799
use nand4 g12198
timestamp 1386234936
transform 1 0 51720 0 1 -823
box 0 0 144 799
use and2 g12264
timestamp 1386234845
transform 1 0 51864 0 1 -823
box 0 0 120 799
use nand3 g12274
timestamp 1386234893
transform 1 0 51984 0 1 -823
box 0 0 120 799
use inv g12288
timestamp 1386238110
transform 1 0 52104 0 1 -823
box 0 0 120 799
use inv g12290
timestamp 1386238110
transform 1 0 52224 0 1 -823
box 0 0 120 799
use inv g12293
timestamp 1386238110
transform 1 0 52344 0 1 -823
box 0 0 120 799
use inv g12307
timestamp 1386238110
transform 1 0 52464 0 1 -823
box 0 0 120 799
use nand2 g12235
timestamp 1386234792
transform 1 0 52584 0 1 -823
box 0 0 96 799
use nor2 g12271
timestamp 1386235306
transform 1 0 52680 0 1 -823
box 0 0 120 799
use inv g12324
timestamp 1386238110
transform 1 0 52800 0 1 -823
box 0 0 120 799
use inv g12304
timestamp 1386238110
transform 1 0 52920 0 1 -823
box 0 0 120 799
use nand2 g12267
timestamp 1386234792
transform 1 0 53040 0 1 -823
box 0 0 96 799
use inv g12299
timestamp 1386238110
transform 1 0 53136 0 1 -823
box 0 0 120 799
use nand3 g12273
timestamp 1386234893
transform 1 0 53256 0 1 -823
box 0 0 120 799
use inv g12286
timestamp 1386238110
transform 1 0 53376 0 1 -823
box 0 0 120 799
use nand2 g12325
timestamp 1386234792
transform 1 0 53496 0 1 -823
box 0 0 96 799
use nand2 g12281
timestamp 1386234792
transform 1 0 53592 0 1 -823
box 0 0 96 799
use inv g12317
timestamp 1386238110
transform 1 0 53688 0 1 -823
box 0 0 120 799
use nand2 g12289
timestamp 1386234792
transform 1 0 53808 0 1 -823
box 0 0 96 799
use inv g12315
timestamp 1386238110
transform 1 0 53904 0 1 -823
box 0 0 120 799
use nand2 g12285
timestamp 1386234792
transform 1 0 54024 0 1 -823
box 0 0 96 799
use nand2 g12295
timestamp 1386234792
transform 1 0 54120 0 1 -823
box 0 0 96 799
use nand2 g12280
timestamp 1386234792
transform 1 0 54216 0 1 -823
box 0 0 96 799
use inv g12282
timestamp 1386238110
transform 1 0 54312 0 1 -823
box 0 0 120 799
use nor2 g12287
timestamp 1386235306
transform 1 0 54432 0 1 -823
box 0 0 120 799
use nor2 g12297
timestamp 1386235306
transform 1 0 54552 0 1 -823
box 0 0 120 799
use and2 g12302
timestamp 1386234845
transform 1 0 54672 0 1 -823
box 0 0 120 799
use nand2 g12308
timestamp 1386234792
transform 1 0 54792 0 1 -823
box 0 0 96 799
use nand2 g12309
timestamp 1386234792
transform 1 0 54888 0 1 -823
box 0 0 96 799
use nand2 g12312
timestamp 1386234792
transform 1 0 54984 0 1 -823
box 0 0 96 799
use inv g12322
timestamp 1386238110
transform 1 0 55080 0 1 -823
box 0 0 120 799
use nand2 g12310
timestamp 1386234792
transform 1 0 55200 0 1 -823
box 0 0 96 799
use nor2 g12330
timestamp 1386235306
transform 1 0 55296 0 1 -823
box 0 0 120 799
use nor2 g12329
timestamp 1386235306
transform 1 0 55416 0 1 -823
box 0 0 120 799
use inv g12327
timestamp 1386238110
transform 1 0 55536 0 1 -823
box 0 0 120 799
use nand2 g12300
timestamp 1386234792
transform 1 0 55656 0 1 -823
box 0 0 96 799
use nand2 g12305
timestamp 1386234792
transform 1 0 55752 0 1 -823
box 0 0 96 799
use nand2 g12303
timestamp 1386234792
transform 1 0 55848 0 1 -823
box 0 0 96 799
use scandtype IRQ1_reg
timestamp 1386241841
transform 1 0 55944 0 1 -823
box 0 0 624 799
use nand3 g12272
timestamp 1386234893
transform 1 0 56568 0 1 -823
box 0 0 120 799
use nand2 g12296
timestamp 1386234792
transform 1 0 56688 0 1 -823
box 0 0 96 799
use nand2 g12294
timestamp 1386234792
transform 1 0 56784 0 1 -823
box 0 0 96 799
use inv g12320
timestamp 1386238110
transform 1 0 56880 0 1 -823
box 0 0 120 799
use nand2 g12306
timestamp 1386234792
transform 1 0 57000 0 1 -823
box 0 0 96 799
use nand2 g12291
timestamp 1386234792
transform 1 0 57096 0 1 -823
box 0 0 96 799
use nand2 g12313
timestamp 1386234792
transform 1 0 57192 0 1 -823
box 0 0 96 799
use nand2 g12319
timestamp 1386234792
transform 1 0 57288 0 1 -823
box 0 0 96 799
use nand2 g12328
timestamp 1386234792
transform 1 0 57384 0 1 -823
box 0 0 96 799
use nor2 g12298
timestamp 1386235306
transform 1 0 57480 0 1 -823
box 0 0 120 799
use nand2 g12316
timestamp 1386234792
transform 1 0 57600 0 1 -823
box 0 0 96 799
use nor2 g12279
timestamp 1386235306
transform 1 0 57696 0 1 -823
box 0 0 120 799
use and2 g12301
timestamp 1386234845
transform 1 0 57816 0 1 -823
box 0 0 120 799
use nand2 g12314
timestamp 1386234792
transform 1 0 57936 0 1 -823
box 0 0 96 799
use nand2 g12323
timestamp 1386234792
transform 1 0 58032 0 1 -823
box 0 0 96 799
use nand2 g12321
timestamp 1386234792
transform 1 0 58128 0 1 -823
box 0 0 96 799
use nand2 g12326
timestamp 1386234792
transform 1 0 58224 0 1 -823
box 0 0 96 799
use nor2 g12283
timestamp 1386235306
transform 1 0 58320 0 1 -823
box 0 0 120 799
use nor2 g12292
timestamp 1386235306
transform 1 0 58440 0 1 -823
box 0 0 120 799
use nand2 g12318
timestamp 1386234792
transform 1 0 58560 0 1 -823
box 0 0 96 799
use and2 g12311
timestamp 1386234845
transform 1 0 58656 0 1 -823
box 0 0 120 799
use inv g12335
timestamp 1386238110
transform 1 0 58776 0 1 -823
box 0 0 120 799
use inv g12346
timestamp 1386238110
transform 1 0 58896 0 1 -823
box 0 0 120 799
use inv g12347
timestamp 1386238110
transform 1 0 59016 0 1 -823
box 0 0 120 799
use inv g12337
timestamp 1386238110
transform 1 0 59136 0 1 -823
box 0 0 120 799
use inv g12345
timestamp 1386238110
transform 1 0 59256 0 1 -823
box 0 0 120 799
use inv g12340
timestamp 1386238110
transform 1 0 59376 0 1 -823
box 0 0 120 799
use inv g12339
timestamp 1386238110
transform 1 0 59496 0 1 -823
box 0 0 120 799
use inv g12334
timestamp 1386238110
transform 1 0 59616 0 1 -823
box 0 0 120 799
use inv g12341
timestamp 1386238110
transform 1 0 59736 0 1 -823
box 0 0 120 799
use inv g12342
timestamp 1386238110
transform 1 0 59856 0 1 -823
box 0 0 120 799
<< labels >>
rlabel metal1 0 240 0 250 3 OpcodeCondIn[7]
rlabel metal1 0 480 0 490 3 OpcodeCondIn[6]
rlabel metal1 0 720 0 730 3 OpcodeCondIn[5]
rlabel metal1 0 960 0 970 3 OpcodeCondIn[4]
rlabel metal1 0 1200 0 1210 3 OpcodeCondIn[3]
rlabel metal1 0 1440 0 1450 3 OpcodeCondIn[2]
rlabel metal1 0 1680 0 1690 3 OpcodeCondIn[1]
rlabel metal1 0 1920 0 1930 3 OpcodeCondIn[0]
rlabel metal1 0 2160 0 2170 3 Flags[3]
rlabel metal1 0 2400 0 2410 3 Flags[2]
rlabel metal1 0 2640 0 2650 3 Flags[1]
rlabel metal1 0 2880 0 2890 3 Flags[0]
rlabel metal1 0 3120 0 3130 3 nWait
rlabel metal1 0 3360 0 3370 3 nIRQ
rlabel metal1 0 3600 0 3610 3 AluOp[4]
rlabel metal1 0 3840 0 3850 3 AluOp[3]
rlabel metal1 0 4080 0 4090 3 AluOp[2]
rlabel metal1 0 4320 0 4330 3 AluOp[1]
rlabel metal1 0 4560 0 4570 3 AluOp[0]
rlabel metal1 0 4800 0 4810 3 Op1Sel
rlabel metal1 0 5040 0 5050 3 AluEn
rlabel metal1 0 5280 0 5290 3 LrEn
rlabel metal1 0 5520 0 5530 3 LrWe
rlabel metal1 0 5760 0 5770 3 PcWe
rlabel metal1 0 6000 0 6010 3 PcEn
rlabel metal1 0 6240 0 6250 3 IrWe
rlabel metal1 0 6480 0 6490 3 WdSel
rlabel metal1 0 6720 0 6730 3 ImmSel
rlabel metal1 0 6960 0 6970 3 RegWe
rlabel metal1 0 7200 0 7210 3 MemEn
rlabel metal1 0 7440 0 7450 3 nWE
rlabel metal1 0 7680 0 7690 3 nOE
rlabel metal1 0 7920 0 7930 3 nME
rlabel metal1 0 8160 0 8170 3 ENB
rlabel metal1 0 8400 0 8410 3 ALE
rlabel metal1 0 8640 0 8650 3 CFlag
rlabel metal1 0 8880 0 8890 3 LrSel
rlabel metal1 0 9120 0 9130 3 AluWe
rlabel metal1 0 9360 0 9370 3 Op2Sel[1]
rlabel metal1 0 9600 0 9610 3 Op2Sel[0]
rlabel metal1 0 9840 0 9850 3 Rs1Sel[1]
rlabel metal1 0 10080 0 10090 3 Rs1Sel[0]
rlabel metal1 0 10320 0 10330 3 RwSel[1]
rlabel metal1 0 10560 0 10570 3 RwSel[0]
rlabel metal1 0 10800 0 10810 3 AluOR[1]
rlabel metal1 0 11040 0 11050 3 AluOR[0]
rlabel metal1 0 11280 0 11290 3 PcSel[2]
rlabel metal1 0 11520 0 11530 3 PcSel[1]
rlabel metal1 0 11760 0 11770 3 PcSel[0]
rlabel metal1 0 12000 0 12010 3 SysBus[15]
rlabel metal1 0 12240 0 12250 3 SysBus[14]
rlabel metal1 0 12480 0 12490 3 SysBus[13]
rlabel metal1 0 12720 0 12730 3 SysBus[12]
rlabel metal1 0 12960 0 12970 3 SysBus[11]
rlabel metal1 0 13200 0 13210 3 SysBus[10]
rlabel metal1 0 13440 0 13450 3 SysBus[9]
rlabel metal1 0 13680 0 13690 3 SysBus[8]
rlabel metal1 0 13920 0 13930 3 SysBus[7]
rlabel metal1 0 14160 0 14170 3 SysBus[6]
rlabel metal1 0 14400 0 14410 3 SysBus[5]
rlabel metal1 0 14640 0 14650 3 SysBus[4]
rlabel metal1 0 14880 0 14890 3 SysBus[3]
rlabel metal1 0 15120 0 15130 3 SysBus[2]
rlabel metal1 0 15360 0 15370 3 SysBus[1]
rlabel metal1 0 15600 0 15610 3 SysBus[0]
<< end >>
