magic
tech c035u
timestamp 1394708418
<< nwell >>
rect 1464 1428 3240 1826
rect 15048 1428 15432 1826
rect 23086 1428 23856 1826
<< pwell >>
rect 1464 1027 3240 1428
rect 15048 1034 15432 1428
rect 23086 1027 23856 1428
<< pohmic >>
rect 1464 1103 1470 1113
rect 3234 1103 3240 1113
rect 15048 1103 15054 1113
rect 15426 1103 15432 1113
rect 23086 1103 23092 1113
rect 23850 1103 23856 1113
<< nohmic >>
rect 1464 1763 1470 1773
rect 3234 1763 3240 1773
rect 15048 1763 15054 1773
rect 15426 1763 15432 1773
rect 23086 1763 23092 1773
rect 23850 1763 23856 1773
<< psubstratetap >>
rect 1470 1103 3234 1119
rect 15054 1103 15426 1119
rect 23092 1103 23850 1119
<< nsubstratetap >>
rect 1470 1757 3234 1773
rect 15054 1757 15426 1773
rect 23092 1757 23850 1773
<< metal1 >>
rect 3637 2221 6167 2231
rect 4069 2199 6143 2209
rect 4501 2177 6119 2187
rect 4933 2154 5903 2164
rect 5365 2133 5879 2143
rect 5797 2111 5855 2121
rect 4189 2007 5519 2017
rect 4237 1985 5471 1995
rect 3805 1963 5039 1973
rect 3757 1941 5087 1951
rect 3372 1919 4607 1929
rect 3325 1897 4655 1907
rect 3301 1875 3719 1885
rect 3733 1875 4151 1885
rect 4597 1875 5015 1885
rect 5029 1875 5447 1885
rect 3541 1853 3959 1863
rect 3973 1853 4391 1863
rect 4837 1853 5255 1863
rect 5269 1853 5687 1863
rect 3397 1831 3551 1841
rect 3829 1831 3983 1841
rect 4261 1831 4415 1841
rect 4693 1831 4847 1841
rect 5125 1831 5279 1841
rect 5557 1831 5711 1841
rect 1464 1809 3240 1819
rect 15048 1809 15432 1819
rect 23086 1809 23856 1819
rect 1464 1786 3240 1796
rect 15048 1786 15432 1796
rect 23086 1786 23856 1796
rect 1464 1757 1470 1773
rect 3234 1757 3240 1773
rect 1464 1748 3240 1757
rect 15048 1757 15054 1773
rect 15426 1757 15432 1773
rect 15048 1748 15432 1757
rect 23086 1757 23092 1773
rect 23850 1757 23856 1773
rect 23086 1748 23856 1757
rect 1464 1119 3240 1128
rect 1464 1103 1470 1119
rect 3234 1103 3240 1119
rect 15048 1119 15432 1128
rect 15048 1103 15054 1119
rect 15426 1103 15432 1119
rect 23086 1119 23856 1128
rect 23086 1103 23092 1119
rect 23850 1103 23856 1119
rect 1464 1080 3240 1090
rect 15048 1080 15432 1090
rect 1464 1057 3240 1067
rect 15048 1057 15432 1067
rect 1464 1034 3240 1044
rect 15048 1034 15432 1044
rect 20869 28 20903 38
rect 20917 28 20951 38
rect 20965 28 20999 38
rect 21013 28 21047 38
rect 21061 28 21095 38
rect 21109 28 21143 38
rect 21157 28 21191 38
rect 21205 28 21503 38
rect 21517 28 21551 38
rect 21565 28 21599 38
rect 21613 28 21647 38
rect 21661 28 21959 38
rect 21973 28 22007 38
rect 22021 28 22319 38
<< m2contact >>
rect 3623 2219 3637 2233
rect 6167 2219 6181 2233
rect 4055 2197 4069 2211
rect 6143 2197 6157 2211
rect 4487 2175 4501 2189
rect 6119 2175 6133 2189
rect 4919 2152 4933 2166
rect 5903 2152 5917 2166
rect 5351 2130 5365 2144
rect 5879 2130 5893 2144
rect 5783 2109 5797 2123
rect 5855 2108 5869 2122
rect 4175 2005 4189 2019
rect 5519 2005 5533 2019
rect 4223 1983 4237 1997
rect 5471 1983 5485 1997
rect 3791 1961 3805 1975
rect 5039 1961 5053 1975
rect 3743 1939 3757 1953
rect 5087 1939 5101 1953
rect 3358 1917 3372 1931
rect 4607 1917 4621 1931
rect 3311 1895 3325 1909
rect 4655 1895 4669 1909
rect 3287 1873 3301 1887
rect 3719 1873 3733 1887
rect 4151 1873 4165 1887
rect 4583 1873 4597 1887
rect 5015 1873 5029 1887
rect 5447 1873 5461 1887
rect 3527 1851 3541 1865
rect 3959 1851 3973 1865
rect 4391 1851 4405 1865
rect 4823 1851 4837 1865
rect 5255 1851 5269 1865
rect 5687 1851 5701 1865
rect 3383 1829 3397 1843
rect 3551 1829 3565 1843
rect 3815 1829 3829 1843
rect 3983 1829 3997 1843
rect 4247 1829 4261 1843
rect 4415 1829 4429 1843
rect 4679 1829 4693 1843
rect 4847 1829 4861 1843
rect 5111 1829 5125 1843
rect 5279 1829 5293 1843
rect 5543 1829 5557 1843
rect 5711 1829 5725 1843
rect 20855 26 20869 40
rect 20903 26 20917 40
rect 20951 26 20965 40
rect 20999 26 21013 40
rect 21047 26 21061 40
rect 21095 26 21109 40
rect 21143 26 21157 40
rect 21191 26 21205 40
rect 21503 25 21517 39
rect 21551 25 21565 39
rect 21599 25 21613 39
rect 21647 25 21661 39
rect 21959 26 21973 40
rect 22007 26 22021 40
rect 22319 26 22333 40
<< metal2 >>
rect 0 1826 200 2783
rect 216 1826 228 2783
rect 240 1826 252 2783
rect 264 1826 276 2783
rect 288 1826 300 2783
rect 3288 1887 3300 2783
rect 3312 1909 3324 2783
rect 3360 1931 3372 2783
rect 3288 1826 3300 1873
rect 3312 1826 3324 1895
rect 3360 1826 3372 1917
rect 3528 1865 3540 2783
rect 3384 1826 3396 1829
rect 3528 1826 3540 1851
rect 3552 1826 3564 1829
rect 3624 1826 3636 2219
rect 3744 1953 3756 2783
rect 3792 1975 3804 2783
rect 3720 1826 3732 1873
rect 3744 1826 3756 1939
rect 3792 1826 3804 1961
rect 3816 1826 3828 1829
rect 3960 1826 3972 1851
rect 3984 1826 3996 1829
rect 4056 1826 4068 2197
rect 4176 2019 4188 2783
rect 4152 1826 4164 1873
rect 4176 1826 4188 2005
rect 4224 1997 4236 2783
rect 4224 1826 4236 1983
rect 4248 1826 4260 1829
rect 4392 1826 4404 1851
rect 4416 1826 4428 1829
rect 4488 1826 4500 2175
rect 4584 1887 4596 2783
rect 4584 1826 4596 1873
rect 4608 1826 4620 1917
rect 4656 1826 4668 1895
rect 4824 1865 4836 2783
rect 4680 1826 4692 1829
rect 4824 1826 4836 1851
rect 4848 1826 4860 1829
rect 4920 1826 4932 2152
rect 5016 1826 5028 1873
rect 5040 1826 5052 1961
rect 5088 1826 5100 1939
rect 5112 1826 5124 1829
rect 5256 1826 5268 1851
rect 5280 1826 5292 1829
rect 5352 1826 5364 2130
rect 5448 1826 5460 1873
rect 5472 1826 5484 1983
rect 5520 1826 5532 2005
rect 5544 1826 5556 1829
rect 5688 1826 5700 1851
rect 5712 1826 5724 1829
rect 5784 1826 5796 2109
rect 5856 2105 5868 2108
rect 5880 2105 5892 2130
rect 5904 2105 5916 2152
rect 5954 2105 5966 2783
rect 6120 2105 6132 2175
rect 6144 2105 6156 2197
rect 6168 2105 6180 2219
rect 6264 2105 6276 2783
rect 6288 2105 6300 2783
rect 6312 2105 6324 2783
rect 15456 2002 15468 2783
rect 15576 2002 15588 2783
rect 15696 2002 15708 2783
rect 15816 2002 15828 2783
rect 15936 2002 15948 2783
rect 16056 2002 16068 2783
rect 16488 2002 16500 2783
rect 16680 2002 16692 2783
rect 16752 2002 16764 2783
rect 16848 2002 16860 2783
rect 21504 2002 21516 2783
rect 21696 2002 21708 2783
rect 21816 2002 21828 2783
rect 21936 2002 21948 2783
rect 23976 1826 24176 2783
rect 0 0 200 1027
rect 216 0 228 1027
rect 240 0 252 1027
rect 264 0 276 1027
rect 288 0 300 1027
rect 3456 1017 3468 1027
rect 3600 1017 3612 1027
rect 3456 1005 3612 1017
rect 3888 1017 3900 1027
rect 4032 1017 4044 1027
rect 3888 1005 4044 1017
rect 4320 1017 4332 1027
rect 4464 1017 4476 1027
rect 4320 1005 4476 1017
rect 4752 1017 4764 1027
rect 4896 1017 4908 1027
rect 4752 1005 4908 1017
rect 5184 1017 5196 1027
rect 5328 1017 5340 1027
rect 5184 1005 5340 1017
rect 5616 1017 5628 1027
rect 5760 1017 5772 1027
rect 5616 1005 5772 1017
rect 5904 0 5916 487
rect 6648 0 6660 487
rect 6864 0 6876 487
rect 7056 0 7068 487
rect 7800 0 7812 487
rect 8016 0 8028 487
rect 8208 0 8220 487
rect 8952 0 8964 487
rect 9168 0 9180 487
rect 9360 0 9372 487
rect 10104 0 10116 487
rect 10320 0 10332 487
rect 10512 0 10524 487
rect 11256 0 11268 487
rect 11472 0 11484 487
rect 11664 0 11676 487
rect 12408 0 12420 487
rect 12624 0 12636 487
rect 12816 0 12828 487
rect 13560 0 13572 487
rect 13776 0 13788 487
rect 13968 0 13980 487
rect 14712 0 14724 487
rect 14928 0 14940 487
rect 15504 0 15516 763
rect 15768 0 15780 763
rect 15936 0 15948 763
rect 16104 0 16116 763
rect 16128 0 16140 763
rect 16200 0 16212 763
rect 16416 0 16428 763
rect 16560 0 16572 763
rect 16896 0 16908 763
rect 17256 0 17268 763
rect 17664 0 17676 763
rect 18000 0 18012 763
rect 18312 0 18324 763
rect 18648 0 18660 763
rect 18768 0 18780 763
rect 18816 0 18828 763
rect 18984 0 18996 763
rect 20784 0 20796 763
rect 20809 0 20821 763
rect 21096 40 21108 763
rect 20856 0 20868 26
rect 20904 0 20916 26
rect 20952 0 20964 26
rect 21000 0 21012 26
rect 21048 0 21060 26
rect 21096 0 21108 26
rect 21144 0 21156 26
rect 21192 0 21204 26
rect 21432 0 21444 763
rect 21504 0 21516 25
rect 21552 0 21564 25
rect 21600 0 21612 25
rect 21648 0 21660 25
rect 21888 0 21900 763
rect 21960 0 21972 26
rect 22008 0 22020 26
rect 22248 0 22260 763
rect 22320 0 22332 26
rect 22608 0 22620 763
rect 22776 0 22788 763
rect 23016 73 23028 763
rect 23016 61 23748 73
rect 23736 0 23748 61
rect 23976 0 24176 1027
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 0 0 1 1027
box 0 0 1464 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 3240 0 1 1027
box 0 0 192 799
use tiehigh tiehigh_3
timestamp 1386086759
transform 1 0 3432 0 1 1027
box 0 0 48 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 3480 0 1 1027
box 0 0 192 799
use mux2 mux2_8
timestamp 1386235218
transform 1 0 3672 0 1 1027
box 0 0 192 799
use tiehigh tiehigh_4
timestamp 1386086759
transform 1 0 3864 0 1 1027
box 0 0 48 799
use mux2 mux2_9
timestamp 1386235218
transform 1 0 3912 0 1 1027
box 0 0 192 799
use mux2 mux2_10
timestamp 1386235218
transform 1 0 4104 0 1 1027
box 0 0 192 799
use tiehigh tiehigh_5
timestamp 1386086759
transform 1 0 4296 0 1 1027
box 0 0 48 799
use mux2 mux2_11
timestamp 1386235218
transform 1 0 4344 0 1 1027
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4536 0 1 1027
box 0 0 192 799
use tiehigh tiehigh_2
timestamp 1386086759
transform 1 0 4728 0 1 1027
box 0 0 48 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 4776 0 1 1027
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 4968 0 1 1027
box 0 0 192 799
use tiehigh tiehigh_1
timestamp 1386086759
transform 1 0 5160 0 1 1027
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 5208 0 1 1027
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 5400 0 1 1027
box 0 0 192 799
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 5592 0 1 1027
box 0 0 48 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 5640 0 1 1027
box 0 0 192 799
use regBlock_decoder regBlock_decoder_0
timestamp 1394493274
transform 1 0 5832 0 1 487
box 0 0 9216 1618
use ALUDecoder_new ALUDecoder_new_0
timestamp 1394643424
transform 1 0 15432 0 1 763
box 0 0 7654 1239
use rightend rightend_0
timestamp 1386235834
transform 1 0 23856 0 1 1027
box 0 0 320 799
<< labels >>
rlabel metal2 240 2783 252 2783 1 Test
rlabel metal2 264 2783 276 2783 1 Clock
rlabel metal2 288 2783 300 2783 1 nReset
rlabel metal2 0 2783 200 2783 5 Vdd!
rlabel metal2 4824 2783 4836 2783 5 RwSel[1]
rlabel metal2 4176 2783 4188 2783 5 Ir[8]
rlabel metal2 4224 2783 4236 2783 5 Ir[5]
rlabel metal2 3792 2783 3804 2783 5 Ir[6]
rlabel metal2 3744 2783 3756 2783 5 Ir[9]
rlabel metal2 3360 2783 3372 2783 5 Ir[7]
rlabel metal2 3312 2783 3324 2783 5 Ir[10]
rlabel metal2 3528 2783 3540 2783 5 Rs1Sel[1]
rlabel metal2 3288 2783 3300 2783 5 Rs1Sel[0]
rlabel metal2 5954 2783 5966 2783 5 RegWe
rlabel metal2 6312 2783 6324 2783 5 Ir[4]
rlabel metal2 6288 2783 6300 2783 5 Ir[3]
rlabel metal2 6264 2783 6276 2783 5 Ir[2]
rlabel metal2 4584 2783 4596 2783 5 RwSel[0]
rlabel metal2 216 2783 228 2783 5 SDO
rlabel metal2 23976 2783 24176 2783 1 GND!
rlabel metal2 5904 0 5916 0 1 Rw[0]
rlabel metal2 6648 0 6660 0 1 Rs1[0]
rlabel metal2 6864 0 6876 0 1 Rs2[0]
rlabel metal2 8016 0 8028 0 1 Rs2[1]
rlabel metal2 8208 0 8220 0 1 Rw[2]
rlabel metal2 8952 0 8964 0 1 Rs1[2]
rlabel metal2 9168 0 9180 0 1 Rs2[2]
rlabel metal2 9360 0 9372 0 1 Rw[3]
rlabel metal2 10104 0 10116 0 1 Rs1[3]
rlabel metal2 10512 0 10524 0 1 Rw[4]
rlabel metal2 11256 0 11268 0 1 Rs1[4]
rlabel metal2 11472 0 11484 0 1 Rs2[4]
rlabel metal2 11664 0 11676 0 1 Rw[5]
rlabel metal2 12408 0 12420 0 1 Rs1[5]
rlabel metal2 12624 0 12636 0 1 Rs2[5]
rlabel metal2 12816 0 12828 0 1 Rw[6]
rlabel metal2 13560 0 13572 0 1 Rs1[6]
rlabel metal2 13776 0 13788 0 1 Rs2[6]
rlabel metal2 13968 0 13980 0 1 Rw[7]
rlabel metal2 14712 0 14724 0 1 Rs1[7]
rlabel metal2 14928 0 14940 0 1 Rs2[7]
rlabel metal2 7056 0 7068 0 1 Rw[1]
rlabel metal2 7800 0 7812 0 1 Rs1[1]
rlabel metal2 10320 0 10332 0 1 Rs2[3]
rlabel metal2 23978 0 24176 0 1 GND!
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 23736 0 23748 0 1 OutEn
rlabel metal2 22320 0 22332 0 1 Sh1_R_In
rlabel metal2 22008 0 22020 0 5 Sh2B_R
rlabel metal2 21960 0 21972 0 5 Sh2A_R
rlabel metal2 21504 0 21516 0 5 Sh4Z_R
rlabel metal2 21648 0 21660 0 5 Sh4C_R
rlabel metal2 21600 0 21612 0 5 Sh4B_R
rlabel metal2 21552 0 21564 0 5 Sh4A_R
rlabel metal2 21192 0 21204 0 5 Sh8H_R
rlabel metal2 20952 0 20964 0 5 Sh8C_R
rlabel metal2 20904 0 20916 0 5 Sh8B_R
rlabel metal2 20856 0 20868 0 5 Sh8A_R
rlabel metal2 21000 0 21012 0 5 Sh8D_R
rlabel metal2 21048 0 21060 0 5 Sh8E_R
rlabel metal2 21096 0 21108 0 5 Sh8F_R
rlabel metal2 21144 0 21156 0 5 Sh8G_R
rlabel metal2 18312 0 18324 0 1 NAND
rlabel metal2 15768 0 15780 0 1 SUB
rlabel metal2 15936 0 15948 0 1 CIn_slice
rlabel metal2 16104 0 16116 0 1 LastCIn
rlabel metal2 16128 0 16140 0 1 COut
rlabel metal2 16416 0 16428 0 1 nZ
rlabel metal2 16560 0 16572 0 1 FAOut
rlabel metal2 16896 0 16908 0 1 AND
rlabel metal2 17256 0 17268 0 1 OR
rlabel metal2 17664 0 17676 0 1 XOR
rlabel metal2 18000 0 18012 0 1 NOT
rlabel metal2 18984 0 18996 0 1 ShL
rlabel metal2 18768 0 18780 0 1 ASign
rlabel metal2 18816 0 18828 0 1 ShB
rlabel metal2 18648 0 18660 0 1 NOR
rlabel metal2 21432 0 21444 0 1 Sh4
rlabel metal2 22248 0 22260 0 1 Sh1
rlabel metal2 20809 0 20821 0 1 ShR
rlabel metal2 21888 0 21900 0 1 Sh2
rlabel metal2 22608 0 22620 0 1 ShOut
rlabel metal2 22776 0 22788 0 1 LLI
rlabel metal2 15504 0 15516 0 1 ZeroA
rlabel metal2 16200 0 16212 0 1 Flags[3]
rlabel metal2 15696 2783 15708 2783 5 Ir[13]
rlabel metal2 15576 2783 15588 2783 5 Ir[14]
rlabel metal2 15456 2783 15468 2783 5 Ir[15]
rlabel metal2 15816 2783 15828 2783 5 Ir[12]
rlabel metal2 15936 2783 15948 2783 5 Ir[11]
rlabel metal2 16056 2783 16068 2783 5 CFlag
rlabel metal2 16848 2783 16860 2783 5 Flagss[0]
rlabel metal2 16752 2783 16764 2783 5 Flags[3]
rlabel metal2 16680 2783 16692 2783 5 Flags[1]
rlabel metal2 16488 2783 16500 2783 5 Flags[2]
rlabel metal2 21504 2783 21516 2783 5 Ir[3]
rlabel metal2 21696 2783 21708 2783 5 Ir[2]
rlabel metal2 21816 2783 21828 2783 5 Ir[1]
rlabel metal2 21936 2783 21948 2783 5 Ir[0]
rlabel metal2 20784 0 20796 0 1 Sh8
rlabel metal1 5829 2116 5829 2116 1 Rw0
rlabel metal1 5828 2137 5828 2137 1 Rw1
rlabel metal1 5822 2159 5822 2159 1 Rw2
rlabel metal1 5824 2181 5824 2181 1 Rs10
rlabel metal1 5824 2204 5824 2204 1 Rs11
rlabel metal1 5825 2224 5825 2224 1 Rs12
<< end >>
