magic
tech c035u
timestamp 1396314228
<< nwell >>
rect 0 556 192 954
<< pwell >>
rect 0 155 192 556
<< pohmic >>
rect 0 231 6 241
rect 186 231 192 241
<< nohmic >>
rect 0 891 6 901
rect 186 891 192 901
<< psubstratetap >>
rect 6 231 186 247
<< nsubstratetap >>
rect 6 885 186 901
<< metal1 >>
rect 0 1137 192 1147
rect 0 937 192 947
rect 0 914 192 924
rect 0 885 6 901
rect 186 885 192 901
rect 0 876 192 885
rect 0 247 192 256
rect 0 231 6 247
rect 186 231 192 247
rect 0 208 192 218
rect 0 185 192 195
rect 0 162 192 172
rect 0 140 192 150
rect 0 72 192 82
rect 0 28 192 38
<< metal2 >>
rect 48 0 60 1154
<< labels >>
rlabel metal1 0 876 0 901 1 Vdd!
rlabel metal1 0 914 0 924 1 Scan
rlabel metal1 0 937 0 947 1 ScanReturn
rlabel metal1 192 937 192 947 7 ScanReturn
rlabel metal1 0 140 0 150 3 ALUOut
rlabel metal1 192 140 192 150 7 ALUOut
rlabel metal1 192 231 192 256 7 GND!
rlabel metal1 192 208 192 218 7 Clock
rlabel metal1 192 185 192 195 7 Test
rlabel metal1 192 162 192 172 7 nReset
rlabel metal1 0 231 0 256 1 GND!
rlabel metal1 0 208 0 218 1 Clock
rlabel metal1 0 185 0 195 1 Test
rlabel metal1 0 162 0 172 1 nReset
rlabel metal1 192 876 192 901 7 Vdd!
rlabel metal1 192 914 192 924 7 Scan
rlabel metal1 0 28 0 38 3 DataIn
rlabel metal1 0 72 0 82 3 SysBus
rlabel metal1 192 28 192 38 7 DataIn
rlabel metal1 192 72 192 82 7 SysBus
rlabel metal2 48 0 60 0 1 LLI
rlabel metal2 48 1154 60 1154 5 LLI
rlabel metal1 0 1137 0 1147 3 ALUOut
rlabel metal1 192 1137 192 1147 7 ALUOut
<< end >>
