magic
tech c035u
timestamp 1396307000
<< metal1 >>
rect 0 937 2135 947
rect 1261 915 1751 925
rect 1789 915 1943 925
rect 62 893 2806 903
rect 2821 893 2951 903
rect 277 871 431 881
rect 445 871 1511 881
rect 1598 870 1895 880
rect 1981 870 2087 880
rect 2173 870 2231 880
rect 397 44 1391 54
rect 1405 44 1703 54
rect 1717 44 3095 54
<< m2contact >>
rect 2135 935 2149 949
rect 1247 913 1261 927
rect 1751 913 1765 927
rect 1775 913 1789 927
rect 1943 913 1957 927
rect 48 890 62 904
rect 2806 891 2821 905
rect 2951 891 2966 905
rect 263 869 277 883
rect 431 869 445 883
rect 1511 869 1525 883
rect 1583 868 1598 882
rect 1895 868 1909 882
rect 1967 869 1981 883
rect 2087 868 2101 882
rect 2159 868 2173 882
rect 2231 868 2245 882
rect 383 40 397 54
rect 1391 42 1405 56
rect 1703 42 1717 56
rect 3095 42 3109 56
<< metal2 >>
rect 48 865 60 890
rect 216 865 228 954
rect 264 865 276 869
rect 360 865 372 954
rect 432 865 444 869
rect 456 865 540 877
rect 576 865 588 954
rect 1248 877 1260 913
rect 1104 865 1260 877
rect 1320 865 1332 954
rect 1488 865 1500 954
rect 1512 865 1524 869
rect 1560 865 1572 954
rect 1584 865 1596 868
rect 1752 865 1764 913
rect 1776 865 1788 913
rect 1872 865 1884 954
rect 1896 865 1908 868
rect 1944 865 1956 913
rect 1968 865 1980 869
rect 2064 859 2076 954
rect 2088 865 2100 868
rect 2136 865 2148 935
rect 2160 865 2172 868
rect 2232 865 2244 868
rect 2280 865 2292 954
rect 2808 865 2820 891
rect 2952 865 2964 891
rect 3024 865 3036 954
rect 3096 865 3108 954
rect 72 56 84 66
rect 72 44 228 56
rect 216 37 228 44
rect 360 37 372 66
rect 384 54 396 66
rect 576 37 588 66
rect 1320 37 1332 66
rect 1392 56 1404 66
rect 1488 56 1500 66
rect 1680 56 1692 66
rect 1704 56 1716 66
rect 1488 44 1692 56
rect 1488 37 1500 44
rect 1872 37 1884 66
rect 2064 37 2076 66
rect 2280 37 2292 66
rect 2808 37 2820 66
rect 3024 37 3036 66
rect 3096 56 3108 66
rect 3096 37 3108 42
use halfadder halfadder_0
timestamp 1386235204
transform 1 0 0 0 1 66
box 0 0 312 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 312 0 1 66
box 0 0 192 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 504 0 1 66
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 1224 0 1 66
box 0 0 216 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 1440 0 1 66
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 1632 0 1 66
box 0 0 192 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 1824 0 1 66
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 2016 0 1 66
box 0 0 192 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 2208 0 1 66
box 0 0 720 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 2928 0 1 66
box 0 0 216 799
<< labels >>
rlabel metal1 1745 920 1745 920 1 Lr
rlabel metal1 1505 876 1505 876 1 Pc1
rlabel metal1 0 937 0 947 3 PCI_Value
rlabel metal2 216 37 228 37 1 PcIncCin
rlabel metal2 360 37 372 37 1 LrSel
rlabel metal2 576 37 588 37 1 LrWe
rlabel metal2 1320 37 1332 37 1 LrEn
rlabel metal2 1872 37 1884 37 1 PcSel[1]
rlabel metal2 1488 37 1500 37 1 PcSel[0]
rlabel metal2 2280 37 2292 37 1 PcWe
rlabel metal2 2808 37 2820 37 1 Pc
rlabel metal2 3024 37 3036 37 1 PcEn
rlabel metal2 3096 37 3108 37 1 SysBus
rlabel metal2 2064 37 2076 37 1 PcSel[2]
rlabel metal2 1320 954 1332 954 1 LrEn
rlabel metal2 576 954 588 954 1 LrWe
rlabel metal2 360 954 372 954 1 LrSel
rlabel metal2 216 954 228 954 5 PcIncCout
rlabel metal2 1872 954 1884 954 1 PcSel[1]
rlabel metal2 1560 954 1572 954 1 ALU
rlabel metal2 1488 954 1500 954 1 PcSel[0]
rlabel metal2 3024 954 3036 954 1 PcEn
rlabel metal2 2280 954 2292 954 1 PcWe
rlabel metal2 3096 954 3108 954 5 SysBus
rlabel metal2 2064 954 2076 954 5 PcSel[2]
<< end >>
