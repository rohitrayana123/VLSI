anusha                                                a n u s h a          ���J �P r o f i l e           ���J �       0 ��   � ��   ���J � x m l     