magic
tech c035u
timestamp 1394557184
<< error_ps >>
rect 901 1364 902 1366
<< nwell >>
rect -2865 941 207 1339
rect 10719 941 11103 1339
rect 18705 941 18807 1339
<< pwell >>
rect -2865 540 207 941
rect 10719 547 11103 941
rect 18705 540 18807 941
<< pohmic >>
rect -2865 616 -2859 626
rect 201 616 207 626
rect 10719 616 10725 626
rect 11097 616 11103 626
rect 18705 616 18711 626
rect 18801 616 18807 626
<< nohmic >>
rect -2865 1276 -2859 1286
rect 201 1276 207 1286
rect 10719 1276 10725 1286
rect 11097 1276 11103 1286
rect 18705 1276 18711 1286
rect 18801 1276 18807 1286
<< psubstratetap >>
rect -2859 616 201 632
rect 10725 616 11097 632
rect 18711 616 18801 632
<< nsubstratetap >>
rect -2859 1270 201 1286
rect 10725 1270 11097 1286
rect 18711 1270 18801 1286
<< metal1 >>
rect 364 1734 1838 1744
rect 556 1712 1814 1722
rect 748 1690 1790 1700
rect 988 1667 1574 1677
rect 1228 1646 1550 1656
rect 1468 1624 1526 1634
rect 676 1410 1382 1420
rect 484 1388 1142 1398
rect 293 1366 901 1376
rect 268 1344 446 1354
rect 460 1344 638 1354
rect 892 1344 1118 1354
rect 1132 1344 1358 1354
rect -2865 1322 207 1332
rect 10719 1322 11103 1332
rect 18705 1322 18807 1332
rect -2865 1299 207 1309
rect 10719 1299 11103 1309
rect 18705 1299 18807 1309
rect -2865 1270 -2859 1286
rect 201 1270 207 1286
rect -2865 1261 207 1270
rect 10719 1270 10725 1286
rect 11097 1270 11103 1286
rect 10719 1261 11103 1270
rect 18705 1270 18711 1286
rect 18801 1270 18807 1286
rect 18705 1261 18807 1270
rect -2865 632 207 641
rect -2865 616 -2859 632
rect 201 616 207 632
rect 10719 632 11103 641
rect 10719 616 10725 632
rect 11097 616 11103 632
rect 18705 632 18807 641
rect 18705 616 18711 632
rect 18801 616 18807 632
rect -2865 593 207 603
rect 10719 593 11103 603
rect -2865 570 207 580
rect 10719 570 11103 580
rect -2865 547 207 557
rect 10719 547 11103 557
<< m2contact >>
rect 350 1732 364 1746
rect 1838 1732 1852 1746
rect 542 1710 556 1724
rect 1814 1710 1828 1724
rect 734 1688 748 1702
rect 1790 1688 1804 1702
rect 974 1665 988 1679
rect 1574 1665 1588 1679
rect 1214 1643 1228 1657
rect 1550 1643 1564 1657
rect 1454 1622 1468 1636
rect 1526 1621 1540 1635
rect 662 1408 676 1422
rect 1382 1408 1396 1422
rect 470 1386 484 1400
rect 1142 1386 1156 1400
rect 279 1364 293 1378
rect 901 1364 915 1378
rect 254 1342 268 1356
rect 446 1342 460 1356
rect 638 1342 652 1356
rect 878 1342 892 1356
rect 1118 1342 1132 1356
rect 1358 1342 1372 1356
<< metal2 >>
rect -4329 1339 -4129 1795
rect -4113 1339 -4101 1795
rect -4089 1339 -4077 1795
rect -4065 1339 -4053 1795
rect -4041 1339 -4029 1795
rect 255 1356 267 1795
rect 279 1378 291 1795
rect 255 1339 267 1342
rect 279 1339 291 1364
rect 327 1339 339 1795
rect 351 1339 363 1732
rect 471 1400 483 1795
rect 447 1339 459 1342
rect 471 1339 483 1386
rect 519 1339 531 1795
rect 543 1339 555 1710
rect 663 1422 675 1795
rect 639 1339 651 1342
rect 663 1339 675 1408
rect 711 1339 723 1795
rect 735 1339 747 1688
rect 879 1356 891 1795
rect 879 1339 891 1342
rect 903 1339 915 1364
rect 975 1338 987 1665
rect 1119 1339 1131 1342
rect 1143 1338 1155 1386
rect 1215 1339 1227 1643
rect 1359 1339 1371 1342
rect 1383 1339 1395 1408
rect 1455 1339 1467 1622
rect 1527 1618 1539 1621
rect 1551 1618 1563 1643
rect 1575 1618 1587 1665
rect 1625 1618 1637 1795
rect 1791 1618 1803 1688
rect 1815 1618 1827 1710
rect 1839 1618 1851 1732
rect 1935 1618 1947 1795
rect 1959 1618 1971 1795
rect 1983 1618 1995 1795
rect 11295 1623 11307 1795
rect 11415 1623 11427 1795
rect 11535 1623 11547 1795
rect 11655 1623 11667 1795
rect 11775 1623 11787 1795
rect 12951 1623 12963 1795
rect 13383 1623 13395 1795
rect 13575 1623 13587 1795
rect 13647 1623 13659 1795
rect 13743 1623 13755 1795
rect 17415 1623 17427 1795
rect 17631 1623 17643 1795
rect 17751 1623 17763 1795
rect 17871 1623 17883 1795
rect 18255 1623 18267 1795
rect 18927 1339 19127 1795
rect -4329 0 -4129 540
rect -4113 0 -4101 540
rect -4089 0 -4077 540
rect -4065 0 -4053 540
rect -4041 0 -4029 540
rect 807 530 819 540
rect 951 530 963 540
rect 807 518 963 530
rect 1047 530 1059 540
rect 1191 530 1203 540
rect 1047 518 1203 530
rect 1287 530 1299 540
rect 1431 530 1443 540
rect 1287 518 1443 530
rect 11175 0 11187 165
rect 11439 0 11451 165
rect 11607 0 11619 165
rect 11775 0 11787 165
rect 11799 0 11811 165
rect 11871 0 11883 165
rect 12087 0 12099 165
rect 12231 0 12243 165
rect 12567 0 12579 165
rect 12927 0 12939 165
rect 13335 0 13347 165
rect 13671 0 13683 165
rect 13983 0 13995 165
rect 14319 0 14331 165
rect 14439 0 14451 165
rect 14487 0 14499 165
rect 14655 0 14667 165
rect 16455 0 16467 165
rect 16480 0 16492 165
rect 16839 0 16851 165
rect 17103 0 17115 165
rect 17559 0 17571 165
rect 17919 0 17931 165
rect 18279 0 18291 165
rect 18447 0 18459 165
rect 18687 0 18699 165
rect 18927 0 19127 540
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 -4329 0 1 540
box 0 0 1464 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 207 0 1 540
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 399 0 1 540
box 0 0 192 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 591 0 1 540
box 0 0 192 799
use tiehigh tiehigh_2
timestamp 1386086759
transform 1 0 783 0 1 540
box 0 0 48 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 831 0 1 540
box 0 0 192 799
use tiehigh tiehigh_1
timestamp 1386086759
transform 1 0 1023 0 1 540
box 0 0 48 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 1071 0 1 540
box 0 0 192 799
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 1263 0 1 540
box 0 0 48 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 1311 0 1 540
box 0 0 192 799
use regBlock_decoder regBlock_decoder_0
timestamp 1394493274
transform 1 0 1503 0 1 0
box 0 0 9216 1618
use ALUDecoder ALUDecoder_0
timestamp 1394549670
transform 1 0 11103 0 1 165
box 0 0 7602 1459
use rightend rightend_0
timestamp 1386235834
transform 1 0 18807 0 1 540
box 0 0 320 799
<< labels >>
rlabel metal2 -4113 0 -4101 0 1 SDI
rlabel metal2 -4089 0 -4077 0 1 Test
rlabel metal2 -4065 0 -4053 0 1 Clock
rlabel metal2 -4041 0 -4029 0 1 nReset
rlabel metal2 -4113 1795 -4101 1795 1 SDI
rlabel metal2 -4089 1795 -4077 1795 1 Test
rlabel metal2 -4065 1795 -4053 1795 1 Clock
rlabel metal2 -4041 1795 -4029 1795 1 nReset
rlabel metal2 -4329 1795 -4129 1795 5 Vdd!
rlabel metal2 -4329 0 -4129 0 1 Vdd!
rlabel metal2 1935 1795 1947 1795 5 Ir[2]
rlabel metal2 1959 1795 1971 1795 5 Ir[3]
rlabel metal2 1983 1795 1995 1795 5 Ir[4]
rlabel metal2 663 1795 675 1795 5 Ir[8]
rlabel metal2 471 1795 483 1795 5 Ir[9]
rlabel metal2 279 1795 291 1795 5 Ir[10]
rlabel metal2 879 1795 891 1795 5 RwSel
rlabel metal2 327 1795 339 1795 5 Ir[7]
rlabel metal2 519 1795 531 1795 5 Ir[6]
rlabel metal2 711 1795 723 1795 5 Ir[5]
rlabel metal2 255 1795 267 1795 5 Rs1Sel
rlabel metal2 1625 1795 1637 1795 5 RegWe
rlabel metal2 11295 1795 11307 1795 5 Ir[15]
rlabel metal2 11415 1795 11427 1795 5 Ir[14]
rlabel metal2 11535 1795 11547 1795 5 Ir[13]
rlabel metal2 11655 1795 11667 1795 5 Ir[12]
rlabel metal2 11775 1795 11787 1795 5 Ir[11]
rlabel metal2 12951 1795 12963 1795 5 CFlag
rlabel metal2 13383 1795 13395 1795 5 Flags[2]
rlabel metal2 13575 1795 13587 1795 5 Flags[1]
rlabel metal2 13647 1795 13659 1795 5 Flags[3]
rlabel metal2 13743 1795 13755 1795 5 Flagss[0]
rlabel metal2 17871 1795 17883 1795 5 Ir[0]
rlabel metal2 17751 1795 17763 1795 5 Ir[1]
rlabel metal2 17631 1795 17643 1795 5 Ir[2]
rlabel metal2 17415 1795 17427 1795 5 Ir[3]
rlabel metal2 18255 1795 18267 1795 5 AluEn
rlabel metal2 18929 0 19127 0 1 GND!
rlabel metal2 18927 1795 19127 1795 1 GND!
rlabel metal2 18687 0 18699 0 1 OutEn
rlabel metal2 18447 0 18459 0 1 LLI
rlabel metal2 18279 0 18291 0 1 ShOut
rlabel metal2 17559 0 17571 0 1 Sh2
rlabel metal2 16480 0 16492 0 1 ShR
rlabel metal2 17919 0 17931 0 1 Sh1
rlabel metal2 17103 0 17115 0 1 Sh4
rlabel metal2 16455 0 16467 0 1 Sh8
rlabel metal2 11175 0 11187 0 1 ZeroA
rlabel metal2 11871 0 11883 0 1 N
rlabel metal2 14319 0 14331 0 1 NOR
rlabel metal2 14487 0 14499 0 1 ShB
rlabel metal2 14439 0 14451 0 1 ASign
rlabel metal2 14655 0 14667 0 1 ShL
rlabel metal2 13671 0 13683 0 1 NOT
rlabel metal2 13335 0 13347 0 1 XOR
rlabel metal2 12927 0 12939 0 1 OR
rlabel metal2 12567 0 12579 0 1 AND
rlabel metal2 12231 0 12243 0 1 FAOut
rlabel metal2 12087 0 12099 0 1 nZ
rlabel metal2 11799 0 11811 0 1 COut
rlabel metal2 11775 0 11787 0 1 LastCIn
rlabel metal2 11607 0 11619 0 1 CIn_slice
rlabel metal2 11439 0 11451 0 1 SUB
rlabel metal2 13983 0 13995 0 1 NAND
rlabel metal2 16839 0 16851 0 1 ShInBit
<< end >>
