magic
tech c035u
timestamp 1394120169
<< metal1 >>
rect 3556 9738 9145 9748
rect 3316 9716 7990 9726
rect 3100 9694 6841 9704
rect 2884 9671 5690 9681
rect 2644 9647 4537 9657
rect 1095 9624 1934 9634
rect 2428 9625 3385 9635
rect 1804 9603 8929 9613
rect 1564 9579 7777 9589
rect 1348 9555 6624 9565
rect 1132 9531 5474 9541
rect 892 9507 4321 9517
rect 676 9486 3169 9496
rect 436 9462 2017 9472
rect 196 9439 865 9449
<< m2contact >>
rect 3542 9736 3556 9750
rect 9145 9736 9159 9750
rect 3302 9714 3316 9728
rect 7990 9714 8004 9728
rect 3086 9692 3100 9706
rect 6841 9691 6855 9705
rect 2870 9667 2884 9681
rect 5690 9669 5704 9683
rect 2630 9645 2644 9659
rect 4537 9645 4551 9659
rect 1081 9622 1095 9636
rect 1934 9623 1948 9637
rect 2414 9625 2428 9639
rect 3385 9623 3399 9637
rect 1790 9599 1804 9613
rect 8929 9601 8943 9615
rect 1550 9575 1564 9589
rect 7777 9578 7791 9592
rect 1334 9551 1348 9565
rect 6624 9554 6638 9568
rect 1118 9527 1132 9541
rect 5474 9529 5488 9543
rect 878 9507 892 9521
rect 4321 9505 4335 9519
rect 662 9485 676 9499
rect 3169 9483 3183 9497
rect 422 9460 436 9474
rect 2017 9462 2031 9476
rect 182 9439 196 9453
rect 865 9437 879 9451
<< metal2 >>
rect 87 11052 99 11121
rect 111 11052 123 11121
rect 135 11052 147 11121
rect 1839 11052 1851 11121
rect 1863 11052 1875 11121
rect 1887 11052 1899 11121
rect 183 9453 195 10098
rect 423 9474 435 10098
rect 663 9499 675 10098
rect 879 9521 891 10098
rect 866 9416 878 9437
rect 1082 9408 1094 9622
rect 1119 9541 1131 10098
rect 1335 9565 1347 10098
rect 1551 9589 1563 10098
rect 1791 9613 1803 10098
rect 1935 9637 1947 10098
rect 2018 9416 2030 9462
rect 2175 9447 2187 10098
rect 2415 9639 2427 10103
rect 2631 9659 2643 10106
rect 2871 9681 2883 10120
rect 3087 9706 3099 10083
rect 3303 9728 3315 10098
rect 3543 9750 3555 10110
rect 2175 9435 2246 9447
rect 2234 9416 2246 9435
rect 3170 9416 3182 9483
rect 3386 9369 3398 9623
rect 4322 9416 4334 9505
rect 4538 9402 4550 9645
rect 5474 9416 5486 9529
rect 5690 9401 5702 9669
rect 6626 9416 6638 9554
rect 6842 9395 6854 9691
rect 7778 9416 7790 9578
rect 7991 9354 8003 9714
rect 8930 9416 8942 9601
rect 9146 9399 9158 9736
use decoder decoder_0
timestamp 1394120018
transform 1 0 63 0 1 10098
box 0 0 1752 954
use decoder decoder_1
timestamp 1394120018
transform 1 0 1815 0 1 10098
box 0 0 1752 954
use regBlock_slice regBlock_slice_0
array 0 0 9385 0 7 1177
timestamp 1394107240
transform 1 0 0 0 1 0
box 0 0 9385 1177
<< labels >>
rlabel metal2 87 11121 99 11121 5 Rs1[0]
rlabel metal2 111 11121 123 11121 5 Rs1[1]
rlabel metal2 135 11121 147 11121 5 Rs1[2]
rlabel metal2 1839 11121 1851 11121 5 Rs2[0]
rlabel metal2 1863 11121 1875 11121 5 Rs2[1]
rlabel metal2 1887 11121 1899 11121 5 Rs2[2]
<< end >>
