../../../Design/Implementation/verilog/behavioural/control.sv