magic
tech c035u
timestamp 1398683468
<< error_ps >>
rect 251 47 263 49
rect 395 47 407 49
rect 611 47 623 49
rect 1355 47 1367 49
rect 1523 47 1535 49
rect 1907 47 1919 49
<< metal1 >>
rect 1608 15759 3247 15769
rect 0 15632 35 15642
rect 3179 15632 3247 15642
rect 0 15609 35 15619
rect 3179 15609 3247 15619
rect 0 15571 35 15596
rect 3179 15571 3247 15596
rect 0 14926 35 14951
rect 3179 14926 3247 14951
rect 0 14903 35 14913
rect 3179 14903 3247 14913
rect 0 14880 35 14890
rect 3179 14880 3247 14890
rect 0 14857 35 14867
rect 3179 14857 3247 14867
rect 3144 14801 3247 14811
rect 1608 14776 3247 14786
rect 0 14649 35 14659
rect 3179 14649 3247 14659
rect 0 14626 35 14636
rect 3179 14626 3247 14636
rect 0 14588 35 14613
rect 3179 14588 3247 14613
rect 0 13943 35 13968
rect 3179 13943 3247 13968
rect 0 13920 35 13930
rect 3179 13920 3247 13930
rect 0 13897 35 13907
rect 3179 13897 3247 13907
rect 0 13874 35 13884
rect 3179 13874 3247 13884
rect 3144 13818 3247 13828
rect 1608 13793 3247 13803
rect 0 13666 35 13676
rect 3179 13666 3247 13676
rect 0 13643 35 13653
rect 3179 13643 3247 13653
rect 0 13605 35 13630
rect 3179 13605 3247 13630
rect 0 12960 35 12985
rect 3179 12960 3247 12985
rect 0 12937 35 12947
rect 3179 12937 3247 12947
rect 0 12914 35 12924
rect 3179 12914 3247 12924
rect 0 12891 35 12901
rect 3179 12891 3247 12901
rect 3144 12835 3247 12845
rect 1608 12810 3247 12820
rect 0 12683 35 12693
rect 3179 12683 3247 12693
rect 0 12660 35 12670
rect 3179 12660 3247 12670
rect 0 12622 35 12647
rect 3179 12622 3247 12647
rect 0 11977 35 12002
rect 3179 11977 3247 12002
rect 0 11954 35 11964
rect 3179 11954 3247 11964
rect 0 11931 35 11941
rect 3179 11931 3247 11941
rect 0 11908 35 11918
rect 3179 11908 3247 11918
rect 3144 11852 3247 11862
rect 1608 11827 3247 11837
rect 0 11700 35 11710
rect 3179 11700 3247 11710
rect 0 11677 35 11687
rect 3179 11677 3247 11687
rect 0 11639 35 11664
rect 3179 11639 3247 11664
rect 0 10994 35 11019
rect 3179 10994 3247 11019
rect 0 10971 35 10981
rect 3179 10971 3247 10981
rect 0 10948 35 10958
rect 3179 10948 3247 10958
rect 0 10925 35 10935
rect 3179 10925 3247 10935
rect 3144 10869 3247 10879
rect 1608 10844 3247 10854
rect 0 10717 35 10727
rect 3179 10717 3247 10727
rect 0 10694 35 10704
rect 3179 10694 3247 10704
rect 0 10656 35 10681
rect 3179 10656 3247 10681
rect 0 10011 35 10036
rect 3179 10011 3247 10036
rect 0 9988 35 9998
rect 3179 9988 3247 9998
rect 0 9965 35 9975
rect 3179 9965 3247 9975
rect 0 9942 35 9952
rect 3179 9942 3247 9952
rect 3144 9886 3247 9896
rect 1608 9861 3247 9871
rect 0 9734 35 9744
rect 3179 9734 3247 9744
rect 0 9711 35 9721
rect 3179 9711 3247 9721
rect 0 9673 35 9698
rect 3179 9673 3247 9698
rect 0 9028 35 9053
rect 3179 9028 3247 9053
rect 0 9005 35 9015
rect 3179 9005 3247 9015
rect 0 8982 35 8992
rect 3179 8982 3247 8992
rect 0 8959 35 8969
rect 3179 8959 3247 8969
rect 3144 8903 3247 8913
rect 1608 8878 3247 8888
rect 0 8751 35 8761
rect 3179 8751 3247 8761
rect 0 8728 35 8738
rect 3179 8728 3247 8738
rect 0 8690 35 8715
rect 3179 8690 3247 8715
rect 0 8045 35 8070
rect 3179 8045 3247 8070
rect 0 8022 35 8032
rect 3179 8022 3247 8032
rect 0 7999 35 8009
rect 3179 7999 3247 8009
rect 0 7976 35 7986
rect 3179 7976 3247 7986
rect 3144 7920 3247 7930
rect 1608 7895 3247 7905
rect 0 7768 35 7778
rect 3179 7768 3247 7778
rect 0 7745 35 7755
rect 3179 7745 3247 7755
rect 0 7707 35 7732
rect 3179 7707 3247 7732
rect 0 7062 35 7087
rect 3179 7062 3247 7087
rect 0 7039 35 7049
rect 3179 7039 3247 7049
rect 0 7016 35 7026
rect 3179 7016 3247 7026
rect 0 6993 35 7003
rect 3179 6993 3247 7003
rect 3144 6937 3247 6947
rect 1608 6912 3247 6922
rect 0 6785 35 6795
rect 3179 6785 3247 6795
rect 0 6762 35 6772
rect 3179 6762 3247 6772
rect 0 6724 35 6749
rect 3179 6724 3247 6749
rect 0 6079 35 6104
rect 3179 6079 3247 6104
rect 0 6056 35 6066
rect 3179 6056 3247 6066
rect 0 6033 35 6043
rect 3179 6033 3247 6043
rect 0 6010 35 6020
rect 3179 6010 3247 6020
rect 3144 5954 3247 5964
rect 1608 5929 3247 5939
rect 0 5802 35 5812
rect 3179 5802 3247 5812
rect 0 5779 35 5789
rect 3179 5779 3247 5789
rect 0 5741 35 5766
rect 3179 5741 3247 5766
rect 0 5096 35 5121
rect 3179 5096 3247 5121
rect 0 5073 35 5083
rect 3179 5073 3247 5083
rect 0 5050 35 5060
rect 3179 5050 3247 5060
rect 0 5027 35 5037
rect 3179 5027 3247 5037
rect 3144 4971 3247 4981
rect 1608 4946 3247 4956
rect 0 4819 35 4829
rect 3179 4819 3247 4829
rect 0 4796 35 4806
rect 3179 4796 3247 4806
rect 0 4758 35 4783
rect 3179 4758 3247 4783
rect 0 4113 35 4138
rect 3179 4113 3247 4138
rect 0 4090 35 4100
rect 3179 4090 3247 4100
rect 0 4067 35 4077
rect 3179 4067 3247 4077
rect 0 4044 35 4054
rect 3179 4044 3247 4054
rect 3144 3988 3247 3998
rect 1608 3963 3247 3973
rect 0 3836 35 3846
rect 3179 3836 3247 3846
rect 0 3813 35 3823
rect 3179 3813 3247 3823
rect 0 3775 35 3800
rect 3179 3775 3247 3800
rect 0 3130 35 3155
rect 3179 3130 3247 3155
rect 0 3107 35 3117
rect 3179 3107 3247 3117
rect 0 3084 35 3094
rect 3179 3084 3247 3094
rect 0 3061 35 3071
rect 3179 3061 3247 3071
rect 3144 3005 3247 3015
rect 1608 2980 3247 2990
rect 0 2853 35 2863
rect 3179 2853 3247 2863
rect 0 2830 35 2840
rect 3179 2830 3247 2840
rect 0 2792 35 2817
rect 3179 2792 3247 2817
rect 0 2147 35 2172
rect 3179 2147 3247 2172
rect 0 2124 35 2134
rect 3179 2124 3247 2134
rect 0 2101 35 2111
rect 3179 2101 3247 2111
rect 0 2078 35 2088
rect 3179 2078 3247 2088
rect 3144 2022 3247 2032
rect 1608 1997 3247 2007
rect 0 1870 35 1880
rect 3179 1870 3247 1880
rect 0 1847 35 1857
rect 3179 1847 3247 1857
rect 0 1809 35 1834
rect 3179 1809 3247 1834
rect 0 1164 35 1189
rect 3179 1164 3247 1189
rect 0 1141 35 1151
rect 3179 1141 3247 1151
rect 0 1118 35 1128
rect 3179 1118 3247 1128
rect 0 1095 35 1105
rect 3179 1095 3247 1105
rect 3144 1039 3247 1049
rect 1608 1014 3247 1024
rect 0 887 35 897
rect 3179 887 3247 897
rect 0 864 35 874
rect 3179 864 3247 874
rect 0 826 35 851
rect 3179 826 3247 851
rect 0 181 35 206
rect 3179 181 3247 206
rect 0 158 35 168
rect 3179 158 3247 168
rect 0 135 35 145
rect 3179 135 3247 145
rect 0 112 35 122
rect 3179 112 3247 122
rect 3144 56 3247 66
<< m2contact >>
rect 1594 15755 1608 15769
rect 3130 14798 3144 14812
rect 1594 14772 1608 14786
rect 3130 13815 3144 13829
rect 1594 13789 1608 13803
rect 3130 12832 3144 12846
rect 1594 12806 1608 12820
rect 3130 11849 3144 11863
rect 1594 11823 1608 11837
rect 3130 10866 3144 10880
rect 1594 10840 1608 10854
rect 3130 9883 3144 9897
rect 1594 9857 1608 9871
rect 3130 8900 3144 8914
rect 1594 8874 1608 8888
rect 3130 7917 3144 7931
rect 1594 7891 1608 7905
rect 3130 6934 3144 6948
rect 1594 6908 1608 6922
rect 3130 5951 3144 5965
rect 1594 5925 1608 5939
rect 3130 4968 3144 4982
rect 1594 4942 1608 4956
rect 3130 3985 3144 3999
rect 1594 3959 1608 3973
rect 3130 3002 3144 3016
rect 1594 2976 1608 2990
rect 3130 2019 3144 2033
rect 1594 1993 1608 2007
rect 3130 1036 3144 1050
rect 1594 1010 1608 1024
rect 3130 53 3144 67
<< metal2 >>
rect 251 15738 263 15955
rect 395 15738 407 15955
rect 611 15738 623 15955
rect 1355 15738 1367 15955
rect 1523 15738 1535 15955
rect 1595 15738 1607 15755
rect 1907 15738 1919 15955
rect 2099 15738 2111 15955
rect 2315 15738 2327 15955
rect 3059 15738 3071 15955
rect 251 14755 263 14821
rect 395 14755 407 14821
rect 611 14755 623 14821
rect 1355 14755 1367 14821
rect 1523 14755 1535 14821
rect 1595 14755 1607 14772
rect 1907 14755 1919 14821
rect 2099 14755 2111 14821
rect 2315 14755 2327 14821
rect 2843 14795 2855 14821
rect 3059 14755 3071 14821
rect 3131 14812 3143 14821
rect 251 13772 263 13838
rect 395 13772 407 13838
rect 611 13772 623 13838
rect 1355 13772 1367 13838
rect 1523 13772 1535 13838
rect 1595 13772 1607 13789
rect 1907 13772 1919 13838
rect 2099 13772 2111 13838
rect 2315 13772 2327 13838
rect 2843 13812 2855 13838
rect 3059 13772 3071 13838
rect 3131 13829 3143 13838
rect 251 12789 263 12855
rect 395 12789 407 12855
rect 611 12789 623 12855
rect 1355 12789 1367 12855
rect 1523 12789 1535 12855
rect 1595 12789 1607 12806
rect 1907 12789 1919 12855
rect 2099 12789 2111 12855
rect 2315 12789 2327 12855
rect 2843 12829 2855 12855
rect 3059 12789 3071 12855
rect 3131 12846 3143 12855
rect 251 11806 263 11872
rect 395 11806 407 11872
rect 611 11806 623 11872
rect 1355 11806 1367 11872
rect 1523 11806 1535 11872
rect 1595 11806 1607 11823
rect 1907 11806 1919 11872
rect 2099 11806 2111 11872
rect 2315 11806 2327 11872
rect 2843 11846 2855 11872
rect 3059 11806 3071 11872
rect 3131 11863 3143 11872
rect 251 10823 263 10889
rect 395 10823 407 10889
rect 611 10823 623 10889
rect 1355 10823 1367 10889
rect 1523 10823 1535 10889
rect 1595 10823 1607 10840
rect 1907 10823 1919 10889
rect 2099 10823 2111 10889
rect 2315 10823 2327 10889
rect 2843 10863 2855 10889
rect 3059 10823 3071 10889
rect 3131 10880 3143 10889
rect 251 9840 263 9906
rect 395 9840 407 9906
rect 611 9840 623 9906
rect 1355 9840 1367 9906
rect 1523 9840 1535 9906
rect 1595 9840 1607 9857
rect 1907 9840 1919 9906
rect 2099 9840 2111 9906
rect 2315 9840 2327 9906
rect 2843 9880 2855 9906
rect 3059 9840 3071 9906
rect 3131 9897 3143 9906
rect 251 8857 263 8923
rect 395 8857 407 8923
rect 611 8857 623 8923
rect 1355 8857 1367 8923
rect 1523 8857 1535 8923
rect 1595 8857 1607 8874
rect 1907 8857 1919 8923
rect 2099 8857 2111 8923
rect 2315 8857 2327 8923
rect 2843 8897 2855 8923
rect 3059 8857 3071 8923
rect 3131 8914 3143 8923
rect 251 7874 263 7940
rect 395 7874 407 7940
rect 611 7874 623 7940
rect 1355 7874 1367 7940
rect 1523 7874 1535 7940
rect 1595 7874 1607 7891
rect 1907 7874 1919 7940
rect 2099 7874 2111 7940
rect 2315 7874 2327 7940
rect 2843 7914 2855 7940
rect 3059 7874 3071 7940
rect 3131 7931 3143 7940
rect 251 6891 263 6957
rect 395 6891 407 6957
rect 611 6891 623 6957
rect 1355 6891 1367 6957
rect 1523 6891 1535 6957
rect 1595 6891 1607 6908
rect 1907 6891 1919 6957
rect 2099 6891 2111 6957
rect 2315 6891 2327 6957
rect 2843 6931 2855 6957
rect 3059 6891 3071 6957
rect 3131 6948 3143 6957
rect 251 5908 263 5974
rect 395 5908 407 5974
rect 611 5908 623 5974
rect 1355 5908 1367 5974
rect 1523 5908 1535 5974
rect 1595 5908 1607 5925
rect 1907 5908 1919 5974
rect 2099 5908 2111 5974
rect 2315 5908 2327 5974
rect 2843 5948 2855 5974
rect 3059 5908 3071 5974
rect 3131 5965 3143 5974
rect 251 4925 263 4991
rect 395 4925 407 4991
rect 611 4925 623 4991
rect 1355 4925 1367 4991
rect 1523 4925 1535 4991
rect 1595 4925 1607 4942
rect 1907 4925 1919 4991
rect 2099 4925 2111 4991
rect 2315 4925 2327 4991
rect 2843 4965 2855 4991
rect 3059 4925 3071 4991
rect 3131 4982 3143 4991
rect 251 3942 263 4008
rect 395 3942 407 4008
rect 611 3942 623 4008
rect 1355 3942 1367 4008
rect 1523 3942 1535 4008
rect 1595 3942 1607 3959
rect 1907 3942 1919 4008
rect 2099 3942 2111 4008
rect 2315 3942 2327 4008
rect 2843 3982 2855 4008
rect 3059 3942 3071 4008
rect 3131 3999 3143 4008
rect 251 2959 263 3025
rect 395 2959 407 3025
rect 611 2959 623 3025
rect 1355 2959 1367 3025
rect 1523 2959 1535 3025
rect 1595 2959 1607 2976
rect 1907 2959 1919 3025
rect 2099 2959 2111 3025
rect 2315 2959 2327 3025
rect 2843 2999 2855 3025
rect 3059 2959 3071 3025
rect 3131 3016 3143 3025
rect 251 1976 263 2042
rect 395 1976 407 2042
rect 611 1976 623 2042
rect 1355 1976 1367 2042
rect 1523 1976 1535 2042
rect 1595 1976 1607 1993
rect 1907 1976 1919 2042
rect 2099 1976 2111 2042
rect 2315 1976 2327 2042
rect 2843 2016 2855 2042
rect 3059 1976 3071 2042
rect 3131 2033 3143 2042
rect 251 993 263 1059
rect 395 993 407 1059
rect 611 993 623 1059
rect 1355 993 1367 1059
rect 1523 993 1535 1059
rect 1595 993 1607 1010
rect 1907 993 1919 1059
rect 2099 993 2111 1059
rect 2315 993 2327 1059
rect 2843 1033 2855 1059
rect 3059 993 3071 1059
rect 3131 1050 3143 1059
rect 251 47 263 76
rect 395 47 407 76
rect 611 47 623 76
rect 1355 47 1367 76
rect 1523 47 1535 76
rect 1907 47 1919 76
rect 2099 47 2111 76
rect 2315 47 2327 76
rect 2843 47 2855 76
rect 3059 47 3071 76
rect 3131 67 3143 76
rect 251 0 263 39
rect 395 0 407 39
rect 611 0 623 39
rect 1355 0 1367 39
rect 1523 0 1535 39
rect 1907 0 1919 39
rect 2123 0 2135 39
rect 2603 0 2615 39
rect 2867 0 2879 39
use Pc_slice Pc_slice_0
array 0 0 3252 0 15 983
timestamp 1396719273
transform 1 0 35 0 1 39
box 0 37 3144 954
<< labels >>
rlabel metal2 2603 0 2615 0 1 Pc
rlabel metal2 2867 0 2879 0 1 PcEn
rlabel metal2 2123 0 2135 0 1 PcWe
rlabel metal2 1907 0 1919 0 1 PcSel[1]
rlabel metal2 1523 0 1535 0 1 PcSel[0]
rlabel metal2 1355 0 1367 0 1 LrEn
rlabel metal2 611 0 623 0 1 LrWe
rlabel metal2 395 0 407 0 1 LrSel
rlabel metal2 251 0 263 0 1 PcIncCin
rlabel metal1 3247 56 3247 66 7 SysBus[0]
rlabel metal1 3247 1039 3247 1049 7 SysBus[1]
rlabel metal1 3247 2022 3247 2032 7 SysBus[2]
rlabel metal1 3247 3005 3247 3015 7 SysBus[3]
rlabel metal1 3247 3988 3247 3998 7 SysBus[4]
rlabel metal1 3247 4971 3247 4981 7 SysBus[5]
rlabel metal1 3247 5954 3247 5964 7 SysBus[6]
rlabel metal1 3247 6937 3247 6947 7 SysBus[7]
rlabel metal1 3247 7920 3247 7930 7 SysBus[8]
rlabel metal1 3247 8903 3247 8913 7 SysBus[9]
rlabel metal1 3247 9886 3247 9896 7 SysBus[10]
rlabel metal1 3247 10869 3247 10879 7 SysBus[11]
rlabel metal1 3247 11852 3247 11862 7 SysBus[12]
rlabel metal1 3247 12835 3247 12845 7 SysBus[13]
rlabel metal1 3247 13818 3247 13828 7 SysBus[14]
rlabel metal1 3247 14801 3247 14811 7 SysBus[15]
rlabel metal1 0 112 0 122 3 nReset
rlabel metal1 0 1095 0 1105 3 nReset
rlabel metal1 0 2078 0 2088 3 nReset
rlabel metal1 0 3061 0 3071 3 nReset
rlabel metal1 0 4044 0 4054 3 nReset
rlabel metal1 0 5027 0 5037 3 nReset
rlabel metal1 0 6010 0 6020 3 nReset
rlabel metal1 0 6993 0 7003 3 nReset
rlabel metal1 0 7976 0 7986 3 nReset
rlabel metal1 0 8959 0 8969 3 nReset
rlabel metal1 0 9942 0 9952 3 nReset
rlabel metal1 0 10925 0 10935 3 nReset
rlabel metal1 0 11908 0 11918 3 nReset
rlabel metal1 0 12891 0 12901 3 nReset
rlabel metal1 0 13874 0 13884 3 nReset
rlabel metal1 0 14857 0 14867 3 nReset
rlabel metal1 0 135 0 145 3 Test
rlabel metal1 0 1118 0 1128 3 Test
rlabel metal1 0 2101 0 2111 3 Test
rlabel metal1 0 3084 0 3094 3 Test
rlabel metal1 0 4067 0 4077 3 Test
rlabel metal1 0 5050 0 5060 3 Test
rlabel metal1 0 6033 0 6043 3 Test
rlabel metal1 0 7016 0 7026 3 Test
rlabel metal1 0 7999 0 8009 3 Test
rlabel metal1 0 8982 0 8992 3 Test
rlabel metal1 0 9965 0 9975 3 Test
rlabel metal1 0 10948 0 10958 3 Test
rlabel metal1 0 11931 0 11941 3 Test
rlabel metal1 0 12914 0 12924 3 Test
rlabel metal1 0 13897 0 13907 3 Test
rlabel metal1 0 14880 0 14890 3 Test
rlabel metal1 0 158 0 168 3 Clock
rlabel metal1 0 1141 0 1151 3 Clock
rlabel metal1 0 2124 0 2134 3 Clock
rlabel metal1 0 3107 0 3117 3 Clock
rlabel metal1 0 4090 0 4100 3 Clock
rlabel metal1 0 5073 0 5083 3 Clock
rlabel metal1 0 6056 0 6066 3 Clock
rlabel metal1 0 7039 0 7049 3 Clock
rlabel metal1 0 8022 0 8032 3 Clock
rlabel metal1 0 9005 0 9015 3 Clock
rlabel metal1 0 9988 0 9998 3 Clock
rlabel metal1 0 10971 0 10981 3 Clock
rlabel metal1 0 11954 0 11964 3 Clock
rlabel metal1 0 12937 0 12947 3 Clock
rlabel metal1 0 13920 0 13930 3 Clock
rlabel metal1 0 14903 0 14913 3 Clock
rlabel metal1 0 181 0 206 3 GND!
rlabel metal1 0 1164 0 1189 3 GND!
rlabel metal1 0 2147 0 2172 3 GND!
rlabel metal1 0 3130 0 3155 3 GND!
rlabel metal1 0 4113 0 4138 3 GND!
rlabel metal1 0 5096 0 5121 3 GND!
rlabel metal1 0 6079 0 6104 3 GND!
rlabel metal1 0 7062 0 7087 3 GND!
rlabel metal1 0 8045 0 8070 3 GND!
rlabel metal1 0 9028 0 9053 3 GND!
rlabel metal1 0 10011 0 10036 3 GND!
rlabel metal1 0 10994 0 11019 3 GND!
rlabel metal1 0 11977 0 12002 3 GND!
rlabel metal1 0 12960 0 12985 3 GND!
rlabel metal1 0 13943 0 13968 3 GND!
rlabel metal1 0 14926 0 14951 3 GND!
rlabel metal1 0 887 0 897 3 ScanReturn
rlabel metal1 0 1870 0 1880 3 ScanReturn
rlabel metal1 0 2853 0 2863 3 ScanReturn
rlabel metal1 0 3836 0 3846 3 ScanReturn
rlabel metal1 0 4819 0 4829 3 ScanReturn
rlabel metal1 0 5802 0 5812 3 ScanReturn
rlabel metal1 0 6785 0 6795 3 ScanReturn
rlabel metal1 0 7768 0 7778 3 ScanReturn
rlabel metal1 0 8751 0 8761 3 ScanReturn
rlabel metal1 0 9734 0 9744 3 ScanReturn
rlabel metal1 0 10717 0 10727 3 ScanReturn
rlabel metal1 0 11700 0 11710 3 ScanReturn
rlabel metal1 0 12683 0 12693 3 ScanReturn
rlabel metal1 0 13666 0 13676 3 ScanReturn
rlabel metal1 0 14649 0 14659 3 ScanReturn
rlabel metal1 0 15632 0 15642 3 ScanReturn
rlabel metal1 0 864 0 874 3 Scan
rlabel metal1 0 1847 0 1857 3 Scan
rlabel metal1 0 2830 0 2840 3 Scan
rlabel metal1 0 3813 0 3823 3 Scan
rlabel metal1 0 4796 0 4806 3 Scan
rlabel metal1 0 5779 0 5789 3 Scan
rlabel metal1 0 6762 0 6772 3 Scan
rlabel metal1 0 7745 0 7755 3 Scan
rlabel metal1 0 8728 0 8738 3 Scan
rlabel metal1 0 9711 0 9721 3 Scan
rlabel metal1 0 10694 0 10704 3 Scan
rlabel metal1 0 11677 0 11687 3 Scan
rlabel metal1 0 12660 0 12670 3 Scan
rlabel metal1 0 13643 0 13653 3 Scan
rlabel metal1 0 14626 0 14636 3 Scan
rlabel metal1 0 15609 0 15619 3 Scan
rlabel metal1 0 826 0 851 3 Vdd!
rlabel metal1 0 1809 0 1834 3 Vdd!
rlabel metal1 0 2792 0 2817 3 Vdd!
rlabel metal1 0 3775 0 3800 3 Vdd!
rlabel metal1 0 4758 0 4783 3 Vdd!
rlabel metal1 0 5741 0 5766 3 Vdd!
rlabel metal1 0 6724 0 6749 3 Vdd!
rlabel metal1 0 7707 0 7732 3 Vdd!
rlabel metal1 0 8690 0 8715 3 Vdd!
rlabel metal1 0 9673 0 9698 3 Vdd!
rlabel metal1 0 10656 0 10681 3 Vdd!
rlabel metal1 0 11639 0 11664 3 Vdd!
rlabel metal1 0 12622 0 12647 3 Vdd!
rlabel metal1 0 13605 0 13630 3 Vdd!
rlabel metal1 0 14588 0 14613 3 Vdd!
rlabel metal1 0 15571 0 15596 3 Vdd!
rlabel metal1 3247 112 3247 122 7 nReset
rlabel metal1 3247 1095 3247 1105 7 nReset
rlabel metal1 3247 2078 3247 2088 7 nReset
rlabel metal1 3247 3061 3247 3071 7 nReset
rlabel metal1 3247 4044 3247 4054 7 nReset
rlabel metal1 3247 5027 3247 5037 7 nReset
rlabel metal1 3247 6010 3247 6020 7 nReset
rlabel metal1 3247 6993 3247 7003 7 nReset
rlabel metal1 3247 7976 3247 7986 7 nReset
rlabel metal1 3247 8959 3247 8969 7 nReset
rlabel metal1 3247 9942 3247 9952 7 nReset
rlabel metal1 3247 10925 3247 10935 7 nReset
rlabel metal1 3247 11908 3247 11918 7 nReset
rlabel metal1 3247 12891 3247 12901 7 nReset
rlabel metal1 3247 13874 3247 13884 7 nReset
rlabel metal1 3247 14857 3247 14867 7 nReset
rlabel metal1 3247 135 3247 145 7 Test
rlabel metal1 3247 1118 3247 1128 7 Test
rlabel metal1 3247 2101 3247 2111 7 Test
rlabel metal1 3247 3084 3247 3094 7 Test
rlabel metal1 3247 4067 3247 4077 7 Test
rlabel metal1 3247 5050 3247 5060 7 Test
rlabel metal1 3247 6033 3247 6043 7 Test
rlabel metal1 3247 7016 3247 7026 7 Test
rlabel metal1 3247 7999 3247 8009 7 Test
rlabel metal1 3247 8982 3247 8992 7 Test
rlabel metal1 3247 9965 3247 9975 7 Test
rlabel metal1 3247 10948 3247 10958 7 Test
rlabel metal1 3247 11931 3247 11941 7 Test
rlabel metal1 3247 12914 3247 12924 7 Test
rlabel metal1 3247 13897 3247 13907 7 Test
rlabel metal1 3247 14880 3247 14890 7 Test
rlabel metal1 3247 158 3247 168 7 Clock
rlabel metal1 3247 1141 3247 1151 7 Clock
rlabel metal1 3247 2124 3247 2134 7 Clock
rlabel metal1 3247 3107 3247 3117 7 Clock
rlabel metal1 3247 4090 3247 4100 7 Clock
rlabel metal1 3247 5073 3247 5083 7 Clock
rlabel metal1 3247 6056 3247 6066 7 Clock
rlabel metal1 3247 7039 3247 7049 7 Clock
rlabel metal1 3247 8022 3247 8032 7 Clock
rlabel metal1 3247 9005 3247 9015 7 Clock
rlabel metal1 3247 9988 3247 9998 7 Clock
rlabel metal1 3247 10971 3247 10981 7 Clock
rlabel metal1 3247 11954 3247 11964 7 Clock
rlabel metal1 3247 12937 3247 12947 7 Clock
rlabel metal1 3247 13920 3247 13930 7 Clock
rlabel metal1 3247 14903 3247 14913 7 Clock
rlabel metal1 3247 181 3247 206 7 GND!
rlabel metal1 3247 1164 3247 1189 7 GND!
rlabel metal1 3247 2147 3247 2172 7 GND!
rlabel metal1 3247 3130 3247 3155 7 GND!
rlabel metal1 3247 4113 3247 4138 7 GND!
rlabel metal1 3247 5096 3247 5121 7 GND!
rlabel metal1 3247 6079 3247 6104 7 GND!
rlabel metal1 3247 7062 3247 7087 7 GND!
rlabel metal1 3247 8045 3247 8070 7 GND!
rlabel metal1 3247 9028 3247 9053 7 GND!
rlabel metal1 3247 10011 3247 10036 7 GND!
rlabel metal1 3247 10994 3247 11019 7 GND!
rlabel metal1 3247 11977 3247 12002 7 GND!
rlabel metal1 3247 12960 3247 12985 7 GND!
rlabel metal1 3247 13943 3247 13968 7 GND!
rlabel metal1 3247 14926 3247 14951 7 GND!
rlabel metal1 3247 826 3247 851 7 Vdd!
rlabel metal1 3247 1809 3247 1834 7 Vdd!
rlabel metal1 3247 2792 3247 2817 7 Vdd!
rlabel metal1 3247 3775 3247 3800 7 Vdd!
rlabel metal1 3247 4758 3247 4783 7 Vdd!
rlabel metal1 3247 5741 3247 5766 7 Vdd!
rlabel metal1 3247 6724 3247 6749 7 Vdd!
rlabel metal1 3247 7707 3247 7732 7 Vdd!
rlabel metal1 3247 8690 3247 8715 7 Vdd!
rlabel metal1 3247 9673 3247 9698 7 Vdd!
rlabel metal1 3247 10656 3247 10681 7 Vdd!
rlabel metal1 3247 11639 3247 11664 7 Vdd!
rlabel metal1 3247 12622 3247 12647 7 Vdd!
rlabel metal1 3247 13605 3247 13630 7 Vdd!
rlabel metal1 3247 14588 3247 14613 7 Vdd!
rlabel metal1 3247 15571 3247 15596 7 Vdd!
rlabel metal1 3247 864 3247 874 7 Scan
rlabel metal1 3247 1847 3247 1857 7 Scan
rlabel metal1 3247 2830 3247 2840 7 Scan
rlabel metal1 3247 3813 3247 3823 7 Scan
rlabel metal1 3247 4796 3247 4806 7 Scan
rlabel metal1 3247 5779 3247 5789 7 Scan
rlabel metal1 3247 6762 3247 6772 7 Scan
rlabel metal1 3247 7745 3247 7755 7 Scan
rlabel metal1 3247 8728 3247 8738 7 Scan
rlabel metal1 3247 9711 3247 9721 7 Scan
rlabel metal1 3247 10694 3247 10704 7 Scan
rlabel metal1 3247 11677 3247 11687 7 Scan
rlabel metal1 3247 12660 3247 12670 7 Scan
rlabel metal1 3247 13643 3247 13653 7 Scan
rlabel metal1 3247 14626 3247 14636 7 Scan
rlabel metal1 3247 15609 3247 15619 7 Scan
rlabel metal1 3247 887 3247 897 7 ScanReturn
rlabel metal1 3247 1870 3247 1880 7 ScanReturn
rlabel metal1 3247 2853 3247 2863 7 ScanReturn
rlabel metal1 3247 3836 3247 3846 7 ScanReturn
rlabel metal1 3247 4819 3247 4829 7 ScanReturn
rlabel metal1 3247 5802 3247 5812 7 ScanReturn
rlabel metal1 3247 6785 3247 6795 7 ScanReturn
rlabel metal1 3247 7768 3247 7778 7 ScanReturn
rlabel metal1 3247 8751 3247 8761 7 ScanReturn
rlabel metal1 3247 9734 3247 9744 7 ScanReturn
rlabel metal1 3247 10717 3247 10727 7 ScanReturn
rlabel metal1 3247 11700 3247 11710 7 ScanReturn
rlabel metal1 3247 12683 3247 12693 7 ScanReturn
rlabel metal1 3247 13666 3247 13676 7 ScanReturn
rlabel metal1 3247 14649 3247 14659 7 ScanReturn
rlabel metal1 3247 15632 3247 15642 7 ScanReturn
rlabel metal1 3247 1014 3247 1024 7 ALU[0]
rlabel metal1 3247 1997 3247 2007 7 ALU[1]
rlabel metal1 3247 2980 3247 2990 7 ALU[2]
rlabel metal1 3247 3963 3247 3973 7 ALU[3]
rlabel metal1 3247 4946 3247 4956 7 ALU[4]
rlabel metal1 3247 5929 3247 5939 7 ALU[5]
rlabel metal1 3247 6912 3247 6922 7 ALU[6]
rlabel metal1 3247 7895 3247 7905 7 ALU[7]
rlabel metal1 3247 8878 3247 8888 7 ALU[8]
rlabel metal1 3247 9861 3247 9871 7 ALU[9]
rlabel metal1 3247 10844 3247 10854 7 ALU[10]
rlabel metal1 3247 11827 3247 11837 7 ALU[11]
rlabel metal1 3247 12810 3247 12820 7 ALU[12]
rlabel metal1 3247 13793 3247 13803 7 ALU[13]
rlabel metal1 3247 14776 3247 14786 7 ALU[14]
rlabel metal1 3247 15759 3247 15769 7 ALU[15]
rlabel metal2 395 15955 407 15955 5 LrSel
rlabel metal2 611 15955 623 15955 5 LrWe
rlabel metal2 1355 15955 1367 15955 5 LrEn
rlabel metal2 1523 15955 1535 15955 5 PcSel[0]
rlabel metal2 1907 15955 1919 15955 5 PcSel[1]
rlabel metal2 251 15955 263 15955 5 PcIncCout
rlabel metal2 2099 15955 2111 15955 5 PcSel[2]
rlabel metal2 2315 15955 2327 15955 5 PcWe
rlabel metal2 3059 15955 3071 15955 5 PcEn
<< end >>
