magic
tech c035u
timestamp 1398760078
<< error_s >>
rect 32520 16334 32522 16346
<< error_ps >>
rect 31458 16202 31460 16216
<< nwell >>
rect 6424 36445 36576 36490
rect 6424 6469 6469 36445
rect 36531 6469 36576 36445
rect 6424 6424 36576 6469
<< polysilicon >>
rect 6576 7624 7416 36201
rect 33998 36081 35163 36083
rect 33998 35883 35200 36081
rect 33998 35383 34198 35883
rect 33998 35183 35200 35383
rect 35000 34683 35200 35183
rect 34000 34499 35200 34683
rect 34016 34483 35200 34499
rect 34000 33883 35200 34083
rect 34000 33383 34200 33883
rect 35000 33383 35200 33883
rect 34000 33183 35200 33383
rect 34000 32499 34200 33183
rect 34016 32483 34200 32499
rect 35000 32483 35200 33183
rect 34000 31883 35200 32083
rect 34000 30499 34200 31883
rect 34500 31283 34700 31883
rect 34016 30483 34200 30499
rect 35000 30483 35200 31883
rect 34000 28683 34200 30083
rect 35000 28683 35200 30083
rect 34000 28499 35200 28683
rect 34016 28483 35200 28499
rect 34000 27883 35200 28083
rect 34000 26899 34200 27883
rect 34016 26883 34200 26899
rect 34000 26283 35200 26483
rect 34000 25783 34200 26283
rect 35000 25783 35200 26283
rect 34000 25583 35200 25783
rect 34000 24899 34200 25583
rect 34016 24883 34200 24899
rect 35000 24883 35200 25583
rect 34280 24283 34880 24483
rect 34480 24072 34680 24283
rect 34496 24056 34680 24072
rect 34480 23083 34680 24056
rect 34280 22883 34880 23083
rect 35485 22901 36191 36081
rect 35483 22877 36193 22901
rect 34201 16609 36202 22431
<< nohmic >>
rect 6429 36453 36571 36485
rect 6429 23671 6461 36453
rect 6429 23609 6450 23671
rect 6429 6461 6461 23609
rect 36539 6461 36571 36453
rect 6429 6429 36571 6461
<< polycontact >>
rect 34000 34483 34016 34499
rect 34000 32483 34016 32499
rect 34000 30483 34016 30499
rect 34000 28483 34016 28499
rect 34000 26883 34016 26899
rect 34000 24883 34016 24899
rect 34480 24056 34496 24072
<< nsubstratetap >>
rect 6450 23609 6466 23671
<< metal1 >>
rect 7363 36421 7373 36464
rect 7411 36421 7421 36464
rect 7363 36411 7421 36421
rect 7363 36171 7373 36411
rect 7363 36147 7373 36157
rect 7385 36133 7395 36171
rect 7459 35944 7469 36464
rect 10789 36451 10799 36464
rect 10843 36421 10853 36464
rect 14315 36454 14325 36482
rect 7723 36411 10853 36421
rect 7723 36397 7733 36411
rect 14371 36421 14381 36464
rect 10880 36411 14381 36421
rect 17827 36421 17837 36464
rect 17875 36448 17885 36464
rect 18019 36448 18029 36464
rect 24883 36421 24893 36464
rect 24931 36448 24941 36464
rect 25075 36448 25085 36464
rect 28411 36421 28421 36464
rect 28459 36448 28469 36464
rect 28603 36448 28613 36464
rect 31939 36424 31949 36464
rect 31987 36448 31997 36464
rect 32131 36448 32141 36464
rect 32951 36436 33736 36446
rect 17827 36411 31938 36421
rect 31963 36411 33702 36421
rect 7699 36387 7733 36397
rect 7699 36376 7709 36387
rect 31963 36397 31973 36411
rect 17888 36387 31973 36397
rect 7736 36363 10866 36373
rect 24944 36363 32937 36373
rect 7653 36336 10789 36346
rect 7653 35944 7663 36336
rect 10803 36336 14312 36346
rect 14326 36336 25063 36346
rect 25088 36339 33678 36349
rect 25053 36327 25063 36336
rect 25053 36317 31913 36327
rect 7699 35944 7709 36311
rect 7723 35944 7733 36311
rect 31903 36276 31913 36317
rect 32144 36315 33581 36325
rect 31939 36301 31949 36314
rect 31939 36291 33509 36301
rect 31903 36266 32964 36276
rect 14131 36243 33486 36253
rect 14131 36160 14141 36243
rect 32000 36219 32936 36229
rect 18019 36160 18029 36218
rect 25112 36195 33234 36205
rect 24907 36171 33258 36181
rect 24907 36160 24917 36171
rect 25280 36147 33426 36157
rect 11707 36123 33282 36133
rect 6450 35523 6509 35533
rect 6499 35509 6509 35523
rect 7459 35512 7469 35882
rect 7675 35859 8381 35869
rect 6499 35499 6522 35509
rect 7653 35485 7663 35832
rect 6443 35475 7663 35485
rect 6523 31528 6533 35447
rect 6450 31467 6498 31477
rect 6546 31439 6556 35475
rect 6450 31429 6556 31439
rect 6499 27472 6509 31394
rect 6523 27472 6533 31394
rect 6546 27472 6556 31429
rect 7459 27472 7469 35450
rect 7675 27445 7685 35859
rect 8371 35848 8381 35859
rect 11707 35848 11717 36123
rect 13099 36099 33354 36109
rect 13099 36064 13109 36099
rect 22387 36075 33461 36085
rect 22387 36064 22397 36075
rect 33451 36064 33461 36075
rect 33476 36065 33486 36243
rect 23120 36051 33402 36061
rect 33499 36061 33509 36291
rect 33571 36088 33581 36315
rect 33499 36051 33594 36061
rect 12907 36027 33498 36037
rect 12907 35968 12917 36027
rect 22123 36003 33330 36013
rect 13099 35968 13109 36002
rect 14131 35968 14141 36002
rect 18019 35968 18029 36002
rect 22123 35968 22133 36003
rect 33668 35992 33678 36339
rect 25171 35979 33522 35989
rect 25171 35968 25181 35979
rect 33692 35968 33702 36411
rect 33726 36016 33736 36436
rect 28616 35955 31986 35965
rect 32024 35955 33557 35965
rect 33547 35944 33557 35955
rect 11947 35931 33378 35941
rect 11947 35848 11957 35931
rect 33595 35941 33605 35954
rect 33595 35931 33749 35941
rect 18032 35907 33725 35917
rect 12907 35848 12917 35906
rect 13099 35848 13109 35906
rect 14131 35848 14141 35906
rect 28438 35872 28448 35896
rect 28472 35883 32890 35893
rect 28438 35862 28472 35872
rect 32880 35869 32890 35883
rect 32950 35883 33629 35893
rect 32880 35859 33605 35869
rect 6450 27435 7685 27445
rect 6433 27387 6546 27397
rect 6499 24261 6509 27362
rect 6523 24288 6533 27362
rect 6499 24251 6557 24261
rect 6523 19552 6533 24226
rect 6547 19552 6557 24251
rect 6450 19491 6509 19501
rect 6499 16285 6509 19491
rect 6523 16309 6533 19490
rect 6547 16336 6557 19490
rect 7459 16336 7469 27410
rect 7699 16360 7709 35834
rect 7482 16323 7626 16333
rect 7723 16333 7733 35834
rect 33235 33160 33245 35834
rect 33259 33160 33269 35834
rect 33283 33160 33293 35834
rect 33331 33160 33341 35834
rect 33355 33160 33365 35834
rect 33379 33160 33389 35834
rect 33403 33160 33413 35834
rect 33427 33160 33437 35834
rect 33451 33160 33461 35834
rect 33475 33160 33485 35834
rect 33499 33160 33509 35834
rect 33523 33160 33533 35834
rect 33547 33160 33557 35834
rect 33571 33160 33581 35834
rect 33595 33160 33605 35859
rect 33619 33160 33629 35883
rect 33643 33160 33653 35882
rect 33667 33160 33677 35882
rect 33691 33160 33701 35882
rect 33715 33133 33725 35907
rect 33739 35725 33749 35931
rect 33739 35715 36550 35725
rect 36499 35704 36509 35715
rect 36475 35667 36550 35677
rect 36475 35557 36485 35667
rect 36499 35560 36509 35642
rect 36451 35547 36485 35557
rect 33914 34475 33924 34499
rect 33948 34486 34000 34496
rect 33914 34465 33948 34475
rect 33211 33131 33725 33133
rect 33186 33123 33725 33131
rect 33186 33121 33221 33123
rect 33186 33061 33221 33065
rect 33691 33061 33701 33098
rect 33186 33055 33701 33061
rect 33211 33051 33701 33055
rect 33235 32056 33245 33026
rect 33259 32056 33269 33026
rect 33283 32056 33293 33026
rect 33331 32056 33341 33026
rect 33355 32056 33365 33026
rect 33379 32056 33389 33026
rect 33403 32056 33413 33026
rect 33427 32056 33437 33026
rect 33451 32056 33461 33026
rect 33475 32056 33485 33026
rect 33499 32056 33509 33026
rect 33523 32056 33533 33026
rect 33547 32056 33557 33026
rect 33571 32056 33581 33026
rect 33595 32056 33605 33026
rect 33619 32056 33629 33026
rect 33643 32056 33653 33026
rect 33667 32029 33677 33026
rect 33914 32474 33924 32498
rect 33948 32486 34000 32496
rect 33914 32464 33948 32474
rect 33211 32020 33677 32029
rect 33186 32019 33677 32020
rect 33186 32010 33221 32019
rect 33643 31957 33653 31994
rect 33211 31954 33653 31957
rect 33186 31947 33653 31954
rect 33186 31944 33221 31947
rect 33235 30928 33245 31922
rect 33259 30928 33269 31922
rect 33283 30928 33293 31922
rect 33331 30928 33341 31922
rect 33355 30928 33365 31922
rect 33379 30928 33389 31922
rect 33403 30928 33413 31922
rect 33427 30928 33437 31922
rect 33451 30928 33461 31922
rect 33475 30928 33485 31922
rect 33499 30928 33509 31922
rect 33523 30928 33533 31922
rect 33547 30928 33557 31922
rect 33571 30928 33581 31922
rect 33595 30928 33605 31922
rect 33186 30901 33221 30909
rect 33619 30901 33629 31922
rect 36451 31669 36461 35547
rect 36475 35523 36550 35533
rect 36475 31672 36485 35523
rect 36499 31693 36509 35498
rect 36499 31683 36550 31693
rect 36499 31672 36509 31683
rect 36427 31659 36461 31669
rect 36427 31552 36437 31659
rect 36451 31635 36550 31645
rect 36451 31552 36461 31635
rect 36475 31525 36485 31610
rect 36499 31528 36509 31610
rect 33186 30899 33629 30901
rect 33211 30891 33629 30899
rect 36403 31515 36485 31525
rect 33186 30833 33221 30843
rect 33211 30829 33221 30833
rect 33595 30829 33605 30866
rect 33211 30819 33605 30829
rect 33235 29824 33245 30794
rect 33259 29824 33269 30794
rect 33283 29824 33293 30794
rect 33331 29824 33341 30794
rect 33355 29824 33365 30794
rect 33379 29824 33389 30794
rect 33403 29824 33413 30794
rect 33427 29824 33437 30794
rect 33451 29824 33461 30794
rect 33475 29824 33485 30794
rect 33499 29824 33509 30794
rect 33523 29824 33533 30794
rect 33547 29824 33557 30794
rect 33186 29797 33221 29798
rect 33571 29797 33581 30794
rect 33914 30474 33924 30498
rect 33948 30486 34000 30496
rect 33914 30464 33948 30474
rect 33186 29788 33581 29797
rect 33211 29787 33581 29788
rect 33186 29725 33221 29732
rect 33547 29725 33557 29762
rect 33186 29722 33557 29725
rect 33211 29715 33557 29722
rect 33235 28720 33245 29690
rect 33259 28720 33269 29690
rect 33283 28720 33293 29690
rect 33331 28720 33341 29690
rect 33355 28720 33365 29690
rect 33379 28720 33389 29690
rect 33403 28720 33413 29690
rect 33427 28720 33437 29690
rect 33451 28720 33461 29690
rect 33475 28720 33485 29690
rect 33499 28720 33509 29690
rect 33523 28720 33533 29690
rect 36403 28693 36413 31515
rect 36475 31491 36550 31501
rect 33211 28687 36413 28693
rect 33186 28683 36413 28687
rect 33186 28677 33221 28683
rect 36427 28621 36437 31490
rect 33186 28611 36437 28621
rect 33235 27592 33245 28586
rect 33259 27592 33269 28586
rect 33283 27592 33293 28586
rect 33331 27592 33341 28586
rect 33355 27592 33365 28586
rect 33379 27592 33389 28586
rect 33403 27592 33413 28586
rect 33427 27592 33437 28586
rect 33451 27592 33461 28586
rect 33475 27592 33485 28586
rect 33499 27592 33509 28586
rect 33523 27592 33533 28586
rect 33914 28474 33924 28498
rect 33948 28486 34000 28496
rect 33914 28464 33948 28474
rect 36451 27664 36461 31490
rect 36475 27637 36485 31491
rect 36499 27661 36509 31466
rect 36499 27651 36550 27661
rect 36499 27640 36509 27651
rect 36427 27627 36485 27637
rect 33186 27566 33221 27576
rect 33211 27565 33221 27566
rect 36427 27565 36437 27627
rect 36475 27603 36550 27613
rect 33211 27555 36437 27565
rect 36451 27517 36461 27602
rect 33211 27510 36461 27517
rect 33186 27507 36461 27510
rect 33186 27500 33221 27507
rect 36475 27496 36485 27603
rect 36499 27496 36509 27578
rect 33235 26488 33245 27482
rect 33259 26488 33269 27482
rect 33283 26488 33293 27482
rect 33331 26488 33341 27482
rect 33355 26488 33365 27482
rect 33379 26488 33389 27482
rect 33403 26488 33413 27482
rect 33427 26488 33437 27482
rect 33451 26488 33461 27482
rect 33475 26488 33485 27482
rect 33499 26488 33509 27482
rect 33523 26488 33533 27482
rect 36451 27459 36550 27469
rect 33914 26873 33924 26897
rect 33948 26885 34000 26895
rect 33914 26863 33948 26873
rect 33186 26461 33221 26465
rect 36451 26461 36461 27459
rect 33186 26455 36461 26461
rect 33211 26451 36461 26455
rect 33186 26389 33221 26399
rect 36475 26389 36485 27434
rect 33211 26379 36485 26389
rect 33235 25384 33245 26354
rect 33259 25381 33269 26354
rect 33283 25408 33293 26354
rect 33331 25408 33341 26354
rect 33355 25408 33365 26354
rect 33379 25408 33389 26354
rect 33403 25408 33413 26354
rect 33427 25408 33437 26354
rect 33451 25408 33461 26354
rect 33475 25408 33485 26354
rect 33499 25408 33509 26354
rect 33523 25408 33533 26354
rect 33259 25371 33557 25381
rect 33211 25354 33269 25357
rect 33186 25347 33269 25354
rect 33186 25344 33221 25347
rect 33259 25336 33269 25347
rect 33547 25336 33557 25371
rect 33235 25309 33245 25322
rect 33235 25299 33581 25309
rect 33186 25285 33221 25288
rect 33186 25278 33245 25285
rect 33211 25275 33245 25278
rect 33235 24256 33245 25275
rect 33186 24233 33221 24243
rect 33259 24253 33269 25274
rect 33283 24280 33293 25274
rect 33331 24280 33341 25274
rect 33355 24280 33365 25274
rect 33379 24280 33389 25274
rect 33403 24280 33413 25274
rect 33427 24280 33437 25274
rect 33451 24280 33461 25274
rect 33475 24280 33485 25274
rect 33499 24280 33509 25274
rect 33523 24280 33533 25274
rect 33547 24280 33557 25274
rect 33571 24280 33581 25299
rect 33914 24874 33924 24898
rect 33948 24886 34000 24896
rect 33914 24864 33949 24874
rect 33259 24243 33605 24253
rect 33211 24229 33221 24233
rect 33595 24232 33605 24243
rect 33211 24219 33269 24229
rect 33259 24208 33269 24219
rect 33211 24177 33317 24181
rect 33186 24171 33317 24177
rect 33186 24167 33221 24171
rect 33235 23152 33245 24146
rect 33259 23152 33269 24146
rect 33283 23152 33293 24146
rect 33307 23152 33317 24171
rect 33331 23152 33341 24170
rect 33355 23152 33365 24170
rect 33379 23152 33389 24170
rect 33403 23152 33413 24170
rect 33427 23149 33437 24170
rect 33451 23176 33461 24170
rect 33475 23176 33485 24170
rect 33499 23176 33509 24170
rect 33523 23176 33533 24170
rect 33547 23176 33557 24170
rect 33571 23176 33581 24170
rect 33595 23176 33605 24170
rect 34460 24030 34470 24056
rect 34460 24020 34496 24030
rect 33427 23139 33629 23149
rect 33186 23125 33221 23132
rect 33186 23122 33437 23125
rect 33211 23115 33437 23122
rect 33427 23104 33437 23115
rect 33619 23104 33629 23139
rect 33283 23077 33293 23090
rect 33283 23067 33653 23077
rect 33186 23056 33221 23066
rect 33211 23053 33221 23056
rect 33211 23043 33293 23053
rect 33235 22048 33245 23018
rect 33259 22048 33269 23018
rect 33283 22048 33293 23043
rect 33307 22048 33317 23042
rect 33331 22048 33341 23042
rect 33355 22045 33365 23042
rect 33379 22072 33389 23042
rect 33403 22072 33413 23042
rect 33427 22072 33437 23042
rect 33451 22072 33461 23042
rect 33475 22072 33485 23042
rect 33499 22072 33509 23042
rect 33523 22072 33533 23042
rect 33547 22072 33557 23042
rect 33571 22072 33581 23042
rect 33595 22072 33605 23042
rect 33619 22072 33629 23042
rect 33643 22072 33653 23067
rect 33355 22035 33677 22045
rect 33186 22011 33365 22021
rect 33355 21976 33365 22011
rect 33379 21976 33389 22010
rect 33403 21976 33413 22010
rect 33427 21976 33437 22010
rect 33451 21973 33461 22010
rect 33667 22000 33677 22035
rect 33451 21963 33701 21973
rect 33186 21949 33221 21955
rect 33186 21945 33461 21949
rect 33211 21939 33461 21945
rect 33235 20944 33245 21914
rect 33259 20944 33269 21914
rect 33283 20944 33293 21914
rect 33307 20944 33317 21914
rect 33331 20944 33341 21914
rect 33355 20944 33365 21914
rect 33379 20944 33389 21914
rect 33403 20941 33413 21914
rect 33427 20968 33437 21914
rect 33451 20968 33461 21939
rect 33475 20968 33485 21938
rect 33499 20968 33509 21938
rect 33523 20968 33533 21938
rect 33547 20968 33557 21938
rect 33571 20968 33581 21938
rect 33595 20968 33605 21938
rect 33619 20968 33629 21938
rect 33643 20968 33653 21938
rect 33667 20968 33677 21938
rect 33691 20968 33701 21963
rect 33403 20931 33725 20941
rect 33211 20910 33413 20917
rect 33186 20907 33413 20910
rect 33186 20900 33221 20907
rect 33403 20872 33413 20907
rect 33427 20872 33437 20906
rect 33451 20872 33461 20906
rect 33475 20872 33485 20906
rect 33499 20869 33509 20906
rect 33715 20896 33725 20931
rect 33499 20859 33749 20869
rect 33211 20844 33509 20845
rect 33186 20835 33509 20844
rect 33186 20834 33221 20835
rect 33235 19816 33245 20810
rect 33259 19816 33269 20810
rect 33283 19816 33293 20810
rect 33307 19816 33317 20810
rect 33331 19813 33341 20810
rect 33355 19840 33365 20810
rect 33379 19840 33389 20810
rect 33403 19840 33413 20810
rect 33427 19840 33437 20810
rect 33451 19840 33461 20810
rect 33475 19840 33485 20810
rect 33499 19840 33509 20835
rect 33523 19840 33533 20834
rect 33547 19840 33557 20834
rect 33571 19840 33581 20834
rect 33595 19840 33605 20834
rect 33619 19840 33629 20834
rect 33643 19840 33653 20834
rect 33667 19840 33677 20834
rect 33691 19840 33701 20834
rect 33715 19840 33725 20834
rect 33739 19840 33749 20859
rect 33331 19803 33773 19813
rect 33186 19789 33221 19799
rect 33763 19792 33773 19803
rect 33211 19779 33341 19789
rect 33331 19768 33341 19779
rect 33523 19765 33533 19778
rect 33523 19755 33797 19765
rect 33211 19733 33533 19741
rect 33186 19731 33533 19733
rect 33186 19723 33221 19731
rect 33235 18712 33245 19706
rect 33259 18712 33269 19706
rect 33283 18712 33293 19706
rect 33307 18712 33317 19706
rect 33331 18712 33341 19706
rect 33355 18712 33365 19706
rect 33379 18712 33389 19706
rect 33403 18712 33413 19706
rect 33427 18712 33437 19706
rect 33451 18712 33461 19706
rect 33475 18712 33485 19706
rect 33499 18712 33509 19706
rect 33523 18712 33533 19731
rect 33547 18712 33557 19730
rect 33571 18712 33581 19730
rect 33595 18712 33605 19730
rect 33619 18712 33629 19730
rect 33643 18712 33653 19730
rect 33667 18712 33677 19730
rect 33691 18712 33701 19730
rect 33715 18712 33725 19730
rect 33739 18712 33749 19730
rect 33763 18712 33773 19730
rect 33787 18712 33797 19755
rect 33186 18685 33221 18688
rect 33186 18678 33821 18685
rect 33211 18675 33821 18678
rect 33811 18664 33821 18675
rect 33379 18637 33389 18650
rect 33379 18627 33845 18637
rect 33186 18613 33221 18622
rect 33186 18612 33389 18613
rect 33211 18603 33389 18612
rect 33235 17608 33245 18578
rect 33259 17608 33269 18578
rect 33283 17608 33293 18578
rect 33307 17608 33317 18578
rect 33331 17608 33341 18578
rect 33355 17608 33365 18578
rect 33379 17608 33389 18603
rect 33403 17608 33413 18602
rect 33427 17608 33437 18602
rect 33451 17608 33461 18602
rect 33475 17608 33485 18602
rect 33499 17608 33509 18602
rect 33523 17608 33533 18602
rect 33547 17608 33557 18602
rect 33571 17608 33581 18602
rect 33595 17608 33605 18602
rect 33619 17608 33629 18602
rect 33643 17608 33653 18602
rect 33667 17608 33677 18602
rect 33691 17608 33701 18602
rect 33715 17608 33725 18602
rect 33739 17608 33749 18602
rect 33763 17608 33773 18602
rect 33787 17608 33797 18602
rect 33811 17608 33821 18602
rect 33835 17608 33845 18627
rect 33211 17577 33869 17581
rect 33186 17571 33869 17577
rect 33186 17567 33221 17571
rect 33859 17560 33869 17571
rect 33595 17533 33605 17546
rect 33595 17523 33893 17533
rect 33186 17509 33221 17511
rect 33186 17501 33605 17509
rect 33211 17499 33605 17501
rect 33235 16480 33245 17474
rect 33259 16480 33269 17474
rect 33283 16480 33293 17474
rect 33307 16480 33317 17474
rect 33331 16480 33341 17474
rect 33355 16480 33365 17474
rect 33379 16480 33389 17474
rect 33403 16480 33413 17474
rect 33427 16477 33437 17474
rect 33451 16504 33461 17474
rect 33475 16504 33485 17474
rect 33499 16504 33509 17474
rect 33523 16504 33533 17474
rect 33547 16504 33557 17474
rect 33571 16504 33581 17474
rect 33595 16504 33605 17499
rect 33619 16504 33629 17498
rect 33643 16504 33653 17498
rect 33667 16504 33677 17498
rect 33691 16504 33701 17498
rect 33715 16504 33725 17498
rect 33739 16504 33749 17498
rect 33763 16504 33773 17498
rect 33787 16504 33797 17498
rect 33811 16504 33821 17498
rect 33835 16504 33845 17498
rect 33859 16504 33869 17498
rect 33883 16504 33893 17523
rect 33427 16467 33917 16477
rect 33186 16456 33221 16466
rect 33907 16456 33917 16467
rect 33211 16453 33221 16456
rect 33211 16443 33426 16453
rect 33416 16419 33941 16429
rect 33211 16400 33413 16405
rect 33186 16395 33413 16400
rect 33186 16390 33221 16395
rect 7650 16323 7733 16333
rect 6523 16299 7722 16309
rect 7953 16312 8519 16322
rect 33235 16312 33245 16370
rect 33259 16312 33269 16370
rect 33283 16312 33293 16370
rect 33307 16312 33317 16370
rect 33331 16312 33341 16370
rect 33355 16312 33365 16370
rect 33379 16312 33389 16370
rect 33403 16312 33413 16395
rect 33427 16312 33437 16394
rect 6499 16275 7746 16285
rect 7930 16288 8553 16298
rect 33451 16309 33461 16394
rect 33475 16336 33485 16394
rect 33499 16336 33509 16394
rect 33523 16336 33533 16394
rect 33547 16336 33557 16394
rect 33571 16336 33581 16394
rect 33595 16336 33605 16394
rect 33619 16336 33629 16394
rect 33643 16336 33653 16394
rect 33667 16336 33677 16394
rect 33691 16336 33701 16394
rect 33715 16336 33725 16394
rect 33739 16336 33749 16394
rect 33763 16336 33773 16394
rect 33787 16336 33797 16394
rect 33811 16336 33821 16394
rect 33835 16336 33845 16394
rect 33859 16336 33869 16394
rect 33883 16336 33893 16394
rect 33907 16333 33917 16394
rect 33931 16357 33941 16419
rect 33931 16347 35462 16357
rect 33907 16323 35485 16333
rect 33451 16299 35509 16309
rect 6560 16251 7440 16261
rect 7839 16266 8592 16276
rect 7472 16253 7621 16263
rect 7430 16241 7440 16251
rect 7430 16231 7596 16241
rect 7586 15646 7596 16231
rect 7611 15646 7621 16253
rect 7639 15646 7649 16248
rect 7907 16244 8626 16254
rect 7885 16220 8702 16230
rect 7815 16196 8810 16206
rect 7862 16174 8152 16184
rect 7792 16152 8122 16162
rect 7699 15646 7709 16150
rect 7723 15666 7733 16150
rect 7747 15692 7757 16150
rect 8112 16117 8122 16152
rect 8142 16139 8152 16174
rect 8377 16175 8458 16185
rect 8142 16129 8744 16139
rect 8768 16129 8888 16139
rect 8112 16107 8854 16117
rect 8878 16105 8888 16129
rect 9691 15829 9701 16298
rect 9691 15819 10362 15829
rect 10483 15829 10493 16298
rect 11035 15853 11045 16298
rect 11251 15877 11261 16298
rect 11251 15867 11274 15877
rect 11995 15877 12005 16298
rect 11298 15867 11332 15877
rect 11995 15867 12090 15877
rect 12163 15877 12173 16298
rect 12547 15901 12557 16298
rect 12739 15925 12749 16298
rect 12739 15915 12930 15925
rect 12955 15925 12965 16298
rect 13699 15949 13709 16298
rect 13699 15939 13746 15949
rect 12955 15915 13794 15925
rect 13867 15925 13877 16298
rect 32371 16285 32381 16298
rect 17134 16275 32381 16285
rect 13867 15915 14850 15925
rect 14874 15915 14944 15925
rect 17134 15905 17144 16275
rect 32556 16285 32566 16298
rect 32604 16285 32614 16298
rect 32659 16285 32669 16298
rect 32411 16275 32566 16285
rect 32587 16275 32614 16285
rect 32635 16275 32669 16285
rect 32731 16285 32741 16298
rect 32731 16275 33461 16285
rect 29803 16251 31410 16261
rect 12547 15891 15450 15901
rect 15474 15891 15519 15901
rect 17191 15890 17225 15900
rect 12163 15867 17191 15877
rect 17215 15877 17225 15890
rect 17215 15867 17243 15877
rect 11035 15843 18869 15853
rect 10483 15819 18834 15829
rect 18859 15829 18869 15843
rect 19686 15842 19720 15852
rect 18859 15819 19686 15829
rect 19710 15819 19720 15842
rect 20575 15818 20609 15828
rect 8571 15769 8581 15807
rect 8606 15795 12018 15805
rect 12104 15795 20575 15805
rect 20599 15795 20609 15818
rect 21737 15794 21771 15804
rect 8605 15771 8844 15781
rect 8868 15771 10314 15781
rect 10376 15771 17166 15781
rect 17204 15771 21737 15781
rect 21761 15771 21771 15794
rect 8567 15747 14826 15757
rect 14864 15747 21749 15757
rect 8567 15723 8734 15733
rect 8758 15723 12870 15733
rect 12944 15723 21714 15733
rect 21739 15733 21749 15747
rect 23106 15746 23140 15756
rect 21739 15723 23106 15733
rect 23130 15723 23140 15746
rect 23275 15733 23285 16250
rect 23467 15757 23477 16250
rect 23467 15747 23658 15757
rect 23707 15757 23717 16250
rect 24786 15770 24820 15780
rect 23707 15747 24786 15757
rect 24810 15749 24820 15770
rect 23275 15723 25637 15733
rect 8556 15699 8692 15709
rect 8716 15699 13722 15709
rect 13760 15699 25602 15709
rect 25627 15709 25637 15723
rect 25627 15699 25661 15709
rect 7770 15680 7836 15690
rect 8534 15675 15426 15685
rect 15464 15675 23082 15685
rect 23120 15675 25626 15685
rect 25651 15685 25661 15699
rect 27282 15698 27316 15708
rect 25651 15675 27282 15685
rect 27306 15684 27316 15698
rect 27306 15674 27340 15684
rect 7723 15656 7815 15666
rect 8534 15651 8603 15661
rect 8641 15651 13770 15661
rect 13808 15651 24762 15661
rect 24800 15651 27306 15661
rect 27330 15652 27340 15674
rect 7760 15633 7791 15643
rect 8252 15635 8458 15645
rect 8764 15627 8801 15637
rect 8825 15627 10350 15637
rect 11288 15627 20549 15637
rect 6499 15612 8286 15622
rect 6499 15496 6509 15612
rect 8300 15612 8411 15622
rect 20539 15616 20549 15627
rect 21751 15627 23621 15637
rect 23611 15616 23621 15627
rect 23672 15627 28613 15637
rect 28603 15616 28613 15627
rect 6523 15589 8262 15599
rect 6523 15469 6533 15589
rect 8276 15589 8387 15599
rect 28626 15592 28636 15618
rect 29803 15616 29813 16251
rect 31450 16251 32509 16261
rect 32587 16261 32597 16275
rect 32540 16251 32597 16261
rect 30308 16227 32154 16237
rect 30308 15616 30318 16227
rect 32540 16237 32550 16251
rect 32387 16227 32550 16237
rect 30668 16203 31436 16213
rect 30668 15616 30678 16203
rect 31458 16192 31468 16216
rect 31434 16182 31468 16192
rect 32324 16203 32397 16213
rect 32324 15616 32334 16203
rect 32348 16179 32373 16189
rect 32348 15616 32358 16179
rect 32397 16168 32407 16192
rect 32373 16158 32407 16168
rect 32635 15616 32645 16275
rect 33451 16264 33461 16275
rect 33896 16275 35533 16285
rect 33859 16261 33869 16274
rect 33859 16251 35557 16261
rect 35476 16227 35581 16237
rect 33848 16203 35605 16213
rect 33235 15637 33245 16202
rect 33259 15661 33269 16202
rect 33283 15685 33293 16202
rect 33307 15709 33317 16202
rect 33331 15733 33341 16202
rect 33355 15757 33365 16202
rect 33379 15781 33389 16202
rect 33403 15805 33413 16202
rect 33427 15829 33437 16202
rect 33451 15856 33461 16202
rect 33475 15853 33485 16202
rect 33499 15877 33509 16202
rect 33523 15901 33533 16202
rect 33547 15925 33557 16202
rect 33571 15949 33581 16202
rect 33595 15973 33605 16202
rect 33619 15997 33629 16202
rect 33643 16021 33653 16202
rect 33667 16045 33677 16202
rect 33691 16069 33701 16202
rect 33715 16093 33725 16202
rect 33739 16117 33749 16202
rect 33763 16141 33773 16202
rect 33787 16165 33797 16202
rect 33811 16189 33821 16202
rect 33811 16179 35629 16189
rect 33787 16155 35653 16165
rect 33763 16131 35677 16141
rect 33739 16107 35701 16117
rect 33715 16083 35725 16093
rect 33691 16059 35749 16069
rect 33667 16035 35773 16045
rect 33643 16011 35797 16021
rect 33619 15987 35821 15997
rect 33595 15963 35845 15973
rect 33571 15939 35869 15949
rect 33547 15915 35893 15925
rect 33523 15891 35917 15901
rect 33499 15867 35941 15877
rect 33475 15843 35965 15853
rect 33427 15819 35989 15829
rect 33403 15795 36013 15805
rect 33379 15771 36037 15781
rect 36499 15781 36509 27434
rect 36075 15771 36509 15781
rect 33355 15747 36109 15757
rect 33331 15723 36157 15733
rect 33307 15699 36402 15709
rect 33283 15675 36450 15685
rect 33259 15651 36474 15661
rect 33235 15627 36509 15637
rect 28598 15582 28636 15592
rect 36403 15544 36413 15602
rect 36451 15568 36461 15602
rect 36475 15568 36485 15602
rect 36499 15541 36509 15627
rect 36440 15531 36509 15541
rect 36076 15507 36550 15517
rect 36421 15493 36431 15507
rect 6450 15459 6533 15469
rect 6499 11413 6509 15434
rect 7700 15320 7710 15487
rect 36421 15483 36498 15493
rect 36440 15459 36550 15469
rect 36499 15421 36509 15434
rect 36210 15413 36509 15421
rect 35468 15411 36509 15413
rect 35468 15403 36220 15411
rect 35547 15375 36210 15385
rect 7757 15334 7863 15344
rect 7700 15310 7863 15320
rect 6450 11403 6509 11413
rect 7768 11319 7778 15273
rect 7792 11346 7802 15285
rect 7816 11346 7826 15285
rect 7840 11346 7850 15247
rect 35486 15179 35496 15333
rect 35510 15179 35520 15333
rect 35558 15203 35568 15333
rect 35582 15203 35592 15333
rect 35606 15203 35616 15333
rect 35630 15203 35640 15333
rect 35654 15203 35664 15333
rect 35678 15224 35688 15333
rect 35702 15251 35712 15333
rect 35726 15251 35736 15333
rect 35750 15296 35760 15333
rect 36200 15325 36210 15375
rect 36403 15352 36413 15386
rect 36451 15352 36461 15386
rect 36475 15352 36485 15386
rect 36200 15315 36550 15325
rect 35750 15286 35809 15296
rect 35750 15262 35773 15272
rect 35750 15251 35760 15262
rect 35799 15248 35809 15286
rect 35787 15238 35809 15248
rect 35678 15214 36072 15224
rect 35691 15190 35749 15200
rect 36062 15179 36072 15214
rect 35475 15142 35533 15152
rect 35475 15118 36061 15128
rect 35475 15094 35773 15104
rect 35966 15080 35976 15093
rect 35475 15070 35976 15080
rect 35475 15046 35677 15056
rect 7768 11309 7863 11319
rect 7829 11285 7863 11295
rect 7792 11269 7802 11284
rect 7792 11259 7826 11269
rect 6450 7371 7802 7381
rect 7792 7096 7802 7371
rect 7816 7096 7826 11259
rect 7840 7102 7850 11260
rect 35486 8898 35496 15021
rect 35510 8898 35520 15021
rect 35534 11485 35544 15021
rect 35558 11512 35568 15021
rect 35582 11512 35592 15021
rect 35606 11512 35616 15021
rect 35630 11512 35640 15021
rect 35654 11512 35664 15021
rect 35702 11513 35712 15045
rect 35726 11512 35736 15045
rect 35798 11512 35808 15021
rect 35822 11512 35832 15021
rect 35846 11512 35856 15021
rect 35870 11512 35880 15021
rect 35894 11512 35904 15021
rect 35918 11512 35928 15021
rect 35942 11512 35952 15021
rect 35990 11512 36000 15021
rect 36014 11512 36024 15021
rect 36038 11512 36048 15021
rect 36110 11512 36120 15117
rect 36158 11512 36168 15117
rect 36403 11512 36413 15290
rect 36451 11512 36461 15290
rect 36475 11512 36485 15290
rect 35534 11475 36550 11485
rect 36499 11464 36509 11475
rect 35558 8898 35568 11450
rect 35582 8898 35592 11450
rect 35606 8871 35616 11450
rect 35630 8874 35640 11450
rect 35654 8874 35664 11450
rect 35699 8922 35709 11451
rect 35475 8861 35616 8871
rect 35726 8872 35736 11450
rect 35798 8847 35808 11450
rect 35475 8837 35808 8847
rect 35475 8813 35653 8823
rect 35486 7237 35496 8788
rect 35510 7264 35520 8788
rect 35558 7264 35568 8788
rect 35582 7264 35592 8788
rect 35630 7264 35640 8788
rect 35726 7264 35736 8810
rect 35822 7264 35832 11450
rect 35846 7264 35856 11450
rect 35870 7264 35880 11450
rect 35894 7513 35904 11450
rect 35918 7264 35928 11450
rect 35942 7264 35952 11450
rect 35990 7264 36000 11450
rect 36014 7264 36024 11450
rect 36038 7264 36048 11450
rect 36110 7264 36120 11450
rect 36158 7264 36168 11450
rect 36403 11437 36413 11450
rect 36403 11427 36550 11437
rect 36451 7381 36461 11402
rect 36475 11293 36485 11402
rect 36499 11320 36509 11402
rect 36475 11283 36550 11293
rect 36499 7429 36509 11258
rect 36499 7419 36550 7429
rect 36499 7408 36509 7419
rect 36451 7371 36550 7381
rect 36499 7264 36509 7346
rect 35486 7227 36550 7237
rect 35510 7105 35520 7202
rect 35558 7105 35568 7202
rect 35582 7105 35592 7202
rect 35630 7105 35640 7202
rect 35726 7105 35736 7202
rect 35822 7105 35832 7202
rect 35846 7105 35856 7202
rect 7840 7092 7863 7102
rect 7315 7059 7863 7069
rect 7315 6450 7325 7059
rect 7805 7035 7850 7045
rect 35870 7054 35880 7202
rect 35475 7044 35880 7054
rect 7816 6901 7826 7010
rect 7840 6925 7850 7035
rect 35475 7020 35821 7030
rect 35475 6996 35725 7006
rect 8311 6925 8321 6938
rect 12451 6925 12461 6938
rect 7840 6915 8321 6925
rect 10987 6915 12461 6925
rect 7816 6891 8238 6901
rect 7377 6709 7421 6719
rect 7390 6687 7409 6697
rect 7411 6517 7421 6685
rect 10987 6640 10997 6915
rect 12451 6733 12461 6915
rect 14528 6915 15860 6925
rect 18056 6915 22230 6925
rect 22244 6915 25482 6925
rect 25520 6915 28590 6925
rect 28604 6915 31026 6925
rect 35582 6925 35592 6971
rect 31064 6915 35592 6925
rect 14371 6891 35557 6901
rect 14371 6760 14381 6891
rect 35630 6880 35640 6971
rect 25112 6867 25506 6877
rect 28496 6867 31050 6877
rect 32168 6867 35509 6877
rect 14515 6760 14525 6866
rect 15861 6853 15871 6866
rect 15861 6843 22206 6853
rect 35846 6853 35856 7019
rect 22220 6843 35856 6853
rect 17899 6819 35629 6829
rect 17899 6760 17909 6819
rect 35876 6805 35886 6901
rect 25496 6795 35886 6805
rect 18043 6760 18053 6794
rect 25099 6760 25109 6794
rect 35918 6781 35928 7202
rect 35942 6867 35952 7202
rect 35990 6844 36000 7202
rect 31040 6771 35928 6781
rect 12451 6723 15834 6733
rect 36014 6733 36024 7202
rect 36038 6916 36048 7202
rect 15848 6723 36024 6733
rect 14371 6640 14381 6698
rect 14515 6640 14525 6698
rect 17899 6640 17909 6698
rect 18043 6640 18053 6698
rect 24955 6651 34472 6661
rect 24955 6640 24965 6651
rect 36037 6613 36047 6831
rect 7363 6507 7421 6517
rect 7363 6450 7373 6507
rect 7411 6450 7421 6507
rect 10843 6603 36047 6613
rect 10843 6450 10853 6603
rect 32203 6579 32274 6589
rect 10987 6450 10997 6578
rect 14371 6544 14381 6578
rect 14515 6544 14525 6578
rect 17899 6544 17909 6578
rect 18043 6544 18053 6578
rect 24955 6544 24965 6578
rect 25099 6544 25109 6578
rect 28483 6544 28493 6578
rect 32203 6565 32213 6579
rect 36066 6586 36076 6854
rect 36110 6592 36120 7202
rect 36158 6593 36168 7202
rect 34551 6576 36076 6586
rect 32024 6555 32213 6565
rect 36499 6565 36509 7202
rect 32240 6555 36509 6565
rect 28640 6531 32261 6541
rect 11035 6507 32226 6517
rect 11035 6450 11045 6507
rect 14371 6450 14381 6482
rect 14515 6450 14525 6482
rect 14563 6450 14573 6507
rect 17899 6450 17909 6482
rect 18043 6450 18053 6482
rect 18091 6450 18101 6507
rect 24955 6450 24965 6482
rect 25099 6450 25109 6482
rect 25147 6450 25157 6507
rect 28483 6450 28493 6482
rect 28627 6450 28637 6482
rect 28675 6450 28685 6507
rect 32011 6450 32021 6482
rect 32155 6450 32165 6482
rect 32203 6450 32213 6507
rect 32251 6517 32261 6531
rect 32288 6531 36109 6541
rect 32251 6507 34536 6517
rect 34486 6481 36157 6491
<< m2contact >>
rect 7361 36157 7375 36171
rect 7361 36133 7375 36147
rect 10788 36437 10802 36451
rect 14313 36440 14327 36454
rect 10866 36410 10880 36424
rect 17874 36434 17888 36448
rect 18018 36434 18032 36448
rect 24930 36434 24944 36448
rect 25074 36434 25088 36448
rect 28458 36434 28472 36448
rect 28602 36434 28616 36448
rect 31986 36434 32000 36448
rect 32130 36434 32144 36448
rect 32937 36436 32951 36450
rect 31938 36410 31952 36424
rect 17874 36386 17888 36400
rect 7698 36362 7712 36376
rect 7722 36362 7736 36376
rect 10866 36362 10880 36376
rect 24930 36362 24944 36376
rect 32937 36362 32951 36376
rect 10789 36334 10803 36348
rect 14312 36334 14326 36348
rect 25074 36338 25088 36352
rect 7698 36311 7712 36325
rect 7722 36311 7736 36325
rect 31938 36314 31952 36328
rect 32130 36314 32144 36328
rect 32964 36264 32978 36278
rect 18018 36218 18032 36232
rect 31986 36218 32000 36232
rect 32936 36218 32950 36232
rect 25098 36194 25112 36208
rect 33234 36194 33248 36208
rect 33258 36170 33272 36184
rect 14130 36146 14144 36160
rect 18018 36146 18032 36160
rect 24906 36146 24920 36160
rect 25266 36146 25280 36160
rect 33426 36146 33440 36160
rect 7458 35930 7472 35944
rect 7651 35930 7665 35944
rect 7698 35930 7712 35944
rect 7722 35930 7736 35944
rect 7458 35882 7472 35896
rect 7651 35832 7665 35846
rect 6522 35498 6536 35512
rect 7458 35498 7472 35512
rect 6522 35447 6536 35461
rect 6522 31514 6536 31528
rect 6498 31465 6512 31479
rect 7458 35450 7472 35464
rect 6498 31394 6512 31408
rect 6522 31394 6536 31408
rect 6498 27458 6512 27472
rect 6522 27458 6536 27472
rect 6546 27458 6560 27472
rect 7458 27458 7472 27472
rect 33282 36122 33296 36136
rect 33354 36098 33368 36112
rect 13098 36050 13112 36064
rect 22386 36050 22400 36064
rect 23106 36050 23120 36064
rect 33402 36050 33416 36064
rect 33450 36050 33464 36064
rect 33474 36051 33488 36065
rect 33570 36074 33584 36088
rect 33594 36050 33608 36064
rect 33498 36026 33512 36040
rect 13098 36002 13112 36016
rect 14130 36002 14144 36016
rect 18018 36002 18032 36016
rect 33330 36002 33344 36016
rect 33522 35978 33536 35992
rect 33666 35978 33680 35992
rect 33724 36002 33738 36016
rect 12906 35954 12920 35968
rect 13098 35954 13112 35968
rect 14130 35954 14144 35968
rect 18018 35954 18032 35968
rect 22122 35954 22136 35968
rect 25170 35954 25184 35968
rect 28602 35954 28616 35968
rect 31986 35954 32000 35968
rect 32010 35954 32024 35968
rect 33594 35954 33608 35968
rect 33690 35954 33704 35968
rect 33378 35930 33392 35944
rect 33546 35930 33560 35944
rect 12906 35906 12920 35920
rect 13098 35906 13112 35920
rect 14130 35906 14144 35920
rect 18018 35906 18032 35920
rect 28458 35882 28472 35896
rect 32936 35882 32950 35896
rect 7698 35834 7712 35848
rect 7722 35834 7736 35848
rect 8370 35834 8384 35848
rect 11706 35834 11720 35848
rect 11946 35834 11960 35848
rect 12906 35834 12920 35848
rect 13098 35834 13112 35848
rect 14130 35834 14144 35848
rect 33234 35834 33248 35848
rect 33258 35834 33272 35848
rect 33282 35834 33296 35848
rect 33330 35834 33344 35848
rect 33354 35834 33368 35848
rect 33378 35834 33392 35848
rect 33402 35834 33416 35848
rect 33426 35834 33440 35848
rect 33450 35834 33464 35848
rect 33474 35834 33488 35848
rect 33498 35834 33512 35848
rect 33522 35834 33536 35848
rect 33546 35834 33560 35848
rect 33570 35834 33584 35848
rect 7458 27410 7472 27424
rect 6546 27385 6560 27399
rect 6498 27362 6512 27376
rect 6522 27362 6536 27376
rect 6522 24274 6536 24288
rect 6522 24226 6536 24240
rect 6522 19538 6536 19552
rect 6546 19538 6560 19552
rect 6522 19490 6536 19504
rect 6546 19490 6560 19504
rect 7697 16346 7711 16360
rect 6546 16322 6560 16336
rect 7458 16322 7472 16336
rect 7636 16322 7650 16336
rect 33642 35882 33656 35896
rect 33666 35882 33680 35896
rect 33690 35882 33704 35896
rect 33234 33146 33248 33160
rect 33258 33146 33272 33160
rect 33282 33146 33296 33160
rect 33330 33146 33344 33160
rect 33354 33146 33368 33160
rect 33378 33146 33392 33160
rect 33402 33146 33416 33160
rect 33426 33146 33440 33160
rect 33450 33146 33464 33160
rect 33474 33146 33488 33160
rect 33498 33146 33512 33160
rect 33522 33146 33536 33160
rect 33546 33146 33560 33160
rect 33570 33146 33584 33160
rect 33594 33146 33608 33160
rect 33618 33146 33632 33160
rect 33642 33146 33656 33160
rect 33666 33146 33680 33160
rect 33690 33146 33704 33160
rect 36498 35690 36512 35704
rect 36498 35642 36512 35656
rect 33934 34485 33948 34499
rect 33690 33098 33704 33112
rect 33234 33026 33248 33040
rect 33258 33026 33272 33040
rect 33282 33026 33296 33040
rect 33330 33026 33344 33040
rect 33354 33026 33368 33040
rect 33378 33026 33392 33040
rect 33402 33026 33416 33040
rect 33426 33026 33440 33040
rect 33450 33026 33464 33040
rect 33474 33026 33488 33040
rect 33498 33026 33512 33040
rect 33522 33026 33536 33040
rect 33546 33026 33560 33040
rect 33570 33026 33584 33040
rect 33594 33026 33608 33040
rect 33618 33026 33632 33040
rect 33642 33026 33656 33040
rect 33666 33026 33680 33040
rect 33234 32042 33248 32056
rect 33258 32042 33272 32056
rect 33282 32042 33296 32056
rect 33330 32042 33344 32056
rect 33354 32042 33368 32056
rect 33378 32042 33392 32056
rect 33402 32042 33416 32056
rect 33426 32042 33440 32056
rect 33450 32042 33464 32056
rect 33474 32042 33488 32056
rect 33498 32042 33512 32056
rect 33522 32042 33536 32056
rect 33546 32042 33560 32056
rect 33570 32042 33584 32056
rect 33594 32042 33608 32056
rect 33618 32042 33632 32056
rect 33642 32042 33656 32056
rect 33934 32484 33948 32498
rect 33642 31994 33656 32008
rect 33234 31922 33248 31936
rect 33258 31922 33272 31936
rect 33282 31922 33296 31936
rect 33330 31922 33344 31936
rect 33354 31922 33368 31936
rect 33378 31922 33392 31936
rect 33402 31922 33416 31936
rect 33426 31922 33440 31936
rect 33450 31922 33464 31936
rect 33474 31922 33488 31936
rect 33498 31922 33512 31936
rect 33522 31922 33536 31936
rect 33546 31922 33560 31936
rect 33570 31922 33584 31936
rect 33594 31922 33608 31936
rect 33618 31922 33632 31936
rect 33234 30914 33248 30928
rect 33258 30914 33272 30928
rect 33282 30914 33296 30928
rect 33330 30914 33344 30928
rect 33354 30914 33368 30928
rect 33378 30914 33392 30928
rect 33402 30914 33416 30928
rect 33426 30914 33440 30928
rect 33450 30914 33464 30928
rect 33474 30914 33488 30928
rect 33498 30914 33512 30928
rect 33522 30914 33536 30928
rect 33546 30914 33560 30928
rect 33570 30914 33584 30928
rect 33594 30914 33608 30928
rect 36498 35546 36512 35560
rect 36498 35498 36512 35512
rect 36474 31658 36488 31672
rect 36498 31658 36512 31672
rect 36474 31610 36488 31624
rect 36498 31610 36512 31624
rect 36426 31538 36440 31552
rect 36450 31538 36464 31552
rect 33594 30866 33608 30880
rect 33234 30794 33248 30808
rect 33258 30794 33272 30808
rect 33282 30794 33296 30808
rect 33330 30794 33344 30808
rect 33354 30794 33368 30808
rect 33378 30794 33392 30808
rect 33402 30794 33416 30808
rect 33426 30794 33440 30808
rect 33450 30794 33464 30808
rect 33474 30794 33488 30808
rect 33498 30794 33512 30808
rect 33522 30794 33536 30808
rect 33546 30794 33560 30808
rect 33570 30794 33584 30808
rect 33234 29810 33248 29824
rect 33258 29810 33272 29824
rect 33282 29810 33296 29824
rect 33330 29810 33344 29824
rect 33354 29810 33368 29824
rect 33378 29810 33392 29824
rect 33402 29810 33416 29824
rect 33426 29810 33440 29824
rect 33450 29810 33464 29824
rect 33474 29810 33488 29824
rect 33498 29810 33512 29824
rect 33522 29810 33536 29824
rect 33546 29810 33560 29824
rect 33934 30484 33948 30498
rect 33546 29762 33560 29776
rect 33234 29690 33248 29704
rect 33258 29690 33272 29704
rect 33282 29690 33296 29704
rect 33330 29690 33344 29704
rect 33354 29690 33368 29704
rect 33378 29690 33392 29704
rect 33402 29690 33416 29704
rect 33426 29690 33440 29704
rect 33450 29690 33464 29704
rect 33474 29690 33488 29704
rect 33498 29690 33512 29704
rect 33522 29690 33536 29704
rect 33234 28706 33248 28720
rect 33258 28706 33272 28720
rect 33282 28706 33296 28720
rect 33330 28706 33344 28720
rect 33354 28706 33368 28720
rect 33378 28706 33392 28720
rect 33402 28706 33416 28720
rect 33426 28706 33440 28720
rect 33450 28706 33464 28720
rect 33474 28706 33488 28720
rect 33498 28706 33512 28720
rect 33522 28706 33536 28720
rect 36498 31514 36512 31528
rect 36426 31490 36440 31504
rect 36450 31490 36464 31504
rect 33234 28586 33248 28600
rect 33258 28586 33272 28600
rect 33282 28586 33296 28600
rect 33330 28586 33344 28600
rect 33354 28586 33368 28600
rect 33378 28586 33392 28600
rect 33402 28586 33416 28600
rect 33426 28586 33440 28600
rect 33450 28586 33464 28600
rect 33474 28586 33488 28600
rect 33498 28586 33512 28600
rect 33522 28586 33536 28600
rect 33934 28484 33948 28498
rect 36450 27650 36464 27664
rect 36498 31466 36512 31480
rect 33234 27578 33248 27592
rect 33258 27578 33272 27592
rect 33282 27578 33296 27592
rect 33330 27578 33344 27592
rect 33354 27578 33368 27592
rect 33378 27578 33392 27592
rect 33402 27578 33416 27592
rect 33426 27578 33440 27592
rect 33450 27578 33464 27592
rect 33474 27578 33488 27592
rect 33498 27578 33512 27592
rect 33522 27578 33536 27592
rect 36498 27626 36512 27640
rect 36450 27602 36464 27616
rect 36498 27578 36512 27592
rect 33234 27482 33248 27496
rect 33258 27482 33272 27496
rect 33282 27482 33296 27496
rect 33330 27482 33344 27496
rect 33354 27482 33368 27496
rect 33378 27482 33392 27496
rect 33402 27482 33416 27496
rect 33426 27482 33440 27496
rect 33450 27482 33464 27496
rect 33474 27482 33488 27496
rect 33498 27482 33512 27496
rect 33522 27482 33536 27496
rect 36474 27482 36488 27496
rect 36498 27482 36512 27496
rect 33934 26883 33948 26897
rect 33234 26474 33248 26488
rect 33258 26474 33272 26488
rect 33282 26474 33296 26488
rect 33330 26474 33344 26488
rect 33354 26474 33368 26488
rect 33378 26474 33392 26488
rect 33402 26474 33416 26488
rect 33426 26474 33440 26488
rect 33450 26474 33464 26488
rect 33474 26474 33488 26488
rect 33498 26474 33512 26488
rect 33522 26474 33536 26488
rect 36474 27434 36488 27448
rect 36498 27434 36512 27448
rect 33234 26354 33248 26368
rect 33258 26354 33272 26368
rect 33282 26354 33296 26368
rect 33330 26354 33344 26368
rect 33354 26354 33368 26368
rect 33378 26354 33392 26368
rect 33402 26354 33416 26368
rect 33426 26354 33440 26368
rect 33450 26354 33464 26368
rect 33474 26354 33488 26368
rect 33498 26354 33512 26368
rect 33522 26354 33536 26368
rect 33234 25370 33248 25384
rect 33282 25394 33296 25408
rect 33330 25394 33344 25408
rect 33354 25394 33368 25408
rect 33378 25394 33392 25408
rect 33402 25394 33416 25408
rect 33426 25394 33440 25408
rect 33450 25394 33464 25408
rect 33474 25394 33488 25408
rect 33498 25394 33512 25408
rect 33522 25394 33536 25408
rect 33234 25322 33248 25336
rect 33258 25322 33272 25336
rect 33546 25322 33560 25336
rect 33258 25274 33272 25288
rect 33282 25274 33296 25288
rect 33330 25274 33344 25288
rect 33354 25274 33368 25288
rect 33378 25274 33392 25288
rect 33402 25274 33416 25288
rect 33426 25274 33440 25288
rect 33450 25274 33464 25288
rect 33474 25274 33488 25288
rect 33498 25274 33512 25288
rect 33522 25274 33536 25288
rect 33546 25274 33560 25288
rect 33234 24242 33248 24256
rect 33934 24884 33948 24898
rect 33282 24266 33296 24280
rect 33330 24266 33344 24280
rect 33354 24266 33368 24280
rect 33378 24266 33392 24280
rect 33402 24266 33416 24280
rect 33426 24266 33440 24280
rect 33450 24266 33464 24280
rect 33474 24266 33488 24280
rect 33498 24266 33512 24280
rect 33522 24266 33536 24280
rect 33546 24266 33560 24280
rect 33570 24266 33584 24280
rect 33594 24218 33608 24232
rect 33258 24194 33272 24208
rect 33234 24146 33248 24160
rect 33258 24146 33272 24160
rect 33282 24146 33296 24160
rect 33330 24170 33344 24184
rect 33354 24170 33368 24184
rect 33378 24170 33392 24184
rect 33402 24170 33416 24184
rect 33426 24170 33440 24184
rect 33450 24170 33464 24184
rect 33474 24170 33488 24184
rect 33498 24170 33512 24184
rect 33522 24170 33536 24184
rect 33546 24170 33560 24184
rect 33570 24170 33584 24184
rect 33594 24170 33608 24184
rect 33234 23138 33248 23152
rect 33258 23138 33272 23152
rect 33282 23138 33296 23152
rect 33306 23138 33320 23152
rect 33330 23138 33344 23152
rect 33354 23138 33368 23152
rect 33378 23138 33392 23152
rect 33402 23138 33416 23152
rect 34480 24040 34496 24056
rect 33450 23162 33464 23176
rect 33474 23162 33488 23176
rect 33498 23162 33512 23176
rect 33522 23162 33536 23176
rect 33546 23162 33560 23176
rect 33570 23162 33584 23176
rect 33594 23162 33608 23176
rect 33282 23090 33296 23104
rect 33426 23090 33440 23104
rect 33618 23090 33632 23104
rect 33234 23018 33248 23032
rect 33258 23018 33272 23032
rect 33306 23042 33320 23056
rect 33330 23042 33344 23056
rect 33354 23042 33368 23056
rect 33378 23042 33392 23056
rect 33402 23042 33416 23056
rect 33426 23042 33440 23056
rect 33450 23042 33464 23056
rect 33474 23042 33488 23056
rect 33498 23042 33512 23056
rect 33522 23042 33536 23056
rect 33546 23042 33560 23056
rect 33570 23042 33584 23056
rect 33594 23042 33608 23056
rect 33618 23042 33632 23056
rect 33234 22034 33248 22048
rect 33258 22034 33272 22048
rect 33282 22034 33296 22048
rect 33306 22034 33320 22048
rect 33330 22034 33344 22048
rect 33378 22058 33392 22072
rect 33402 22058 33416 22072
rect 33426 22058 33440 22072
rect 33450 22058 33464 22072
rect 33474 22058 33488 22072
rect 33498 22058 33512 22072
rect 33522 22058 33536 22072
rect 33546 22058 33560 22072
rect 33570 22058 33584 22072
rect 33594 22058 33608 22072
rect 33618 22058 33632 22072
rect 33642 22058 33656 22072
rect 33378 22010 33392 22024
rect 33402 22010 33416 22024
rect 33426 22010 33440 22024
rect 33450 22010 33464 22024
rect 33354 21962 33368 21976
rect 33378 21962 33392 21976
rect 33402 21962 33416 21976
rect 33426 21962 33440 21976
rect 33666 21986 33680 22000
rect 33234 21914 33248 21928
rect 33258 21914 33272 21928
rect 33282 21914 33296 21928
rect 33306 21914 33320 21928
rect 33330 21914 33344 21928
rect 33354 21914 33368 21928
rect 33378 21914 33392 21928
rect 33402 21914 33416 21928
rect 33426 21914 33440 21928
rect 33234 20930 33248 20944
rect 33258 20930 33272 20944
rect 33282 20930 33296 20944
rect 33306 20930 33320 20944
rect 33330 20930 33344 20944
rect 33354 20930 33368 20944
rect 33378 20930 33392 20944
rect 33474 21938 33488 21952
rect 33498 21938 33512 21952
rect 33522 21938 33536 21952
rect 33546 21938 33560 21952
rect 33570 21938 33584 21952
rect 33594 21938 33608 21952
rect 33618 21938 33632 21952
rect 33642 21938 33656 21952
rect 33666 21938 33680 21952
rect 33426 20954 33440 20968
rect 33450 20954 33464 20968
rect 33474 20954 33488 20968
rect 33498 20954 33512 20968
rect 33522 20954 33536 20968
rect 33546 20954 33560 20968
rect 33570 20954 33584 20968
rect 33594 20954 33608 20968
rect 33618 20954 33632 20968
rect 33642 20954 33656 20968
rect 33666 20954 33680 20968
rect 33690 20954 33704 20968
rect 33426 20906 33440 20920
rect 33450 20906 33464 20920
rect 33474 20906 33488 20920
rect 33498 20906 33512 20920
rect 33402 20858 33416 20872
rect 33426 20858 33440 20872
rect 33450 20858 33464 20872
rect 33474 20858 33488 20872
rect 33714 20882 33728 20896
rect 33234 20810 33248 20824
rect 33258 20810 33272 20824
rect 33282 20810 33296 20824
rect 33306 20810 33320 20824
rect 33330 20810 33344 20824
rect 33354 20810 33368 20824
rect 33378 20810 33392 20824
rect 33402 20810 33416 20824
rect 33426 20810 33440 20824
rect 33450 20810 33464 20824
rect 33474 20810 33488 20824
rect 33234 19802 33248 19816
rect 33258 19802 33272 19816
rect 33282 19802 33296 19816
rect 33306 19802 33320 19816
rect 33522 20834 33536 20848
rect 33546 20834 33560 20848
rect 33570 20834 33584 20848
rect 33594 20834 33608 20848
rect 33618 20834 33632 20848
rect 33642 20834 33656 20848
rect 33666 20834 33680 20848
rect 33690 20834 33704 20848
rect 33714 20834 33728 20848
rect 33354 19826 33368 19840
rect 33378 19826 33392 19840
rect 33402 19826 33416 19840
rect 33426 19826 33440 19840
rect 33450 19826 33464 19840
rect 33474 19826 33488 19840
rect 33498 19826 33512 19840
rect 33522 19826 33536 19840
rect 33546 19826 33560 19840
rect 33570 19826 33584 19840
rect 33594 19826 33608 19840
rect 33618 19826 33632 19840
rect 33642 19826 33656 19840
rect 33666 19826 33680 19840
rect 33690 19826 33704 19840
rect 33714 19826 33728 19840
rect 33738 19826 33752 19840
rect 33522 19778 33536 19792
rect 33762 19778 33776 19792
rect 33330 19754 33344 19768
rect 33234 19706 33248 19720
rect 33258 19706 33272 19720
rect 33282 19706 33296 19720
rect 33306 19706 33320 19720
rect 33330 19706 33344 19720
rect 33354 19706 33368 19720
rect 33378 19706 33392 19720
rect 33402 19706 33416 19720
rect 33426 19706 33440 19720
rect 33450 19706 33464 19720
rect 33474 19706 33488 19720
rect 33498 19706 33512 19720
rect 33546 19730 33560 19744
rect 33570 19730 33584 19744
rect 33594 19730 33608 19744
rect 33618 19730 33632 19744
rect 33642 19730 33656 19744
rect 33666 19730 33680 19744
rect 33690 19730 33704 19744
rect 33714 19730 33728 19744
rect 33738 19730 33752 19744
rect 33762 19730 33776 19744
rect 33234 18698 33248 18712
rect 33258 18698 33272 18712
rect 33282 18698 33296 18712
rect 33306 18698 33320 18712
rect 33330 18698 33344 18712
rect 33354 18698 33368 18712
rect 33378 18698 33392 18712
rect 33402 18698 33416 18712
rect 33426 18698 33440 18712
rect 33450 18698 33464 18712
rect 33474 18698 33488 18712
rect 33498 18698 33512 18712
rect 33522 18698 33536 18712
rect 33546 18698 33560 18712
rect 33570 18698 33584 18712
rect 33594 18698 33608 18712
rect 33618 18698 33632 18712
rect 33642 18698 33656 18712
rect 33666 18698 33680 18712
rect 33690 18698 33704 18712
rect 33714 18698 33728 18712
rect 33738 18698 33752 18712
rect 33762 18698 33776 18712
rect 33786 18698 33800 18712
rect 33378 18650 33392 18664
rect 33810 18650 33824 18664
rect 33234 18578 33248 18592
rect 33258 18578 33272 18592
rect 33282 18578 33296 18592
rect 33306 18578 33320 18592
rect 33330 18578 33344 18592
rect 33354 18578 33368 18592
rect 33402 18602 33416 18616
rect 33426 18602 33440 18616
rect 33450 18602 33464 18616
rect 33474 18602 33488 18616
rect 33498 18602 33512 18616
rect 33522 18602 33536 18616
rect 33546 18602 33560 18616
rect 33570 18602 33584 18616
rect 33594 18602 33608 18616
rect 33618 18602 33632 18616
rect 33642 18602 33656 18616
rect 33666 18602 33680 18616
rect 33690 18602 33704 18616
rect 33714 18602 33728 18616
rect 33738 18602 33752 18616
rect 33762 18602 33776 18616
rect 33786 18602 33800 18616
rect 33810 18602 33824 18616
rect 33234 17594 33248 17608
rect 33258 17594 33272 17608
rect 33282 17594 33296 17608
rect 33306 17594 33320 17608
rect 33330 17594 33344 17608
rect 33354 17594 33368 17608
rect 33378 17594 33392 17608
rect 33402 17594 33416 17608
rect 33426 17594 33440 17608
rect 33450 17594 33464 17608
rect 33474 17594 33488 17608
rect 33498 17594 33512 17608
rect 33522 17594 33536 17608
rect 33546 17594 33560 17608
rect 33570 17594 33584 17608
rect 33594 17594 33608 17608
rect 33618 17594 33632 17608
rect 33642 17594 33656 17608
rect 33666 17594 33680 17608
rect 33690 17594 33704 17608
rect 33714 17594 33728 17608
rect 33738 17594 33752 17608
rect 33762 17594 33776 17608
rect 33786 17594 33800 17608
rect 33810 17594 33824 17608
rect 33834 17594 33848 17608
rect 33594 17546 33608 17560
rect 33858 17546 33872 17560
rect 33234 17474 33248 17488
rect 33258 17474 33272 17488
rect 33282 17474 33296 17488
rect 33306 17474 33320 17488
rect 33330 17474 33344 17488
rect 33354 17474 33368 17488
rect 33378 17474 33392 17488
rect 33402 17474 33416 17488
rect 33426 17474 33440 17488
rect 33450 17474 33464 17488
rect 33474 17474 33488 17488
rect 33498 17474 33512 17488
rect 33522 17474 33536 17488
rect 33546 17474 33560 17488
rect 33570 17474 33584 17488
rect 33234 16466 33248 16480
rect 33258 16466 33272 16480
rect 33282 16466 33296 16480
rect 33306 16466 33320 16480
rect 33330 16466 33344 16480
rect 33354 16466 33368 16480
rect 33378 16466 33392 16480
rect 33402 16466 33416 16480
rect 33618 17498 33632 17512
rect 33642 17498 33656 17512
rect 33666 17498 33680 17512
rect 33690 17498 33704 17512
rect 33714 17498 33728 17512
rect 33738 17498 33752 17512
rect 33762 17498 33776 17512
rect 33786 17498 33800 17512
rect 33810 17498 33824 17512
rect 33834 17498 33848 17512
rect 33858 17498 33872 17512
rect 33450 16490 33464 16504
rect 33474 16490 33488 16504
rect 33498 16490 33512 16504
rect 33522 16490 33536 16504
rect 33546 16490 33560 16504
rect 33570 16490 33584 16504
rect 33594 16490 33608 16504
rect 33618 16490 33632 16504
rect 33642 16490 33656 16504
rect 33666 16490 33680 16504
rect 33690 16490 33704 16504
rect 33714 16490 33728 16504
rect 33738 16490 33752 16504
rect 33762 16490 33776 16504
rect 33786 16490 33800 16504
rect 33810 16490 33824 16504
rect 33834 16490 33848 16504
rect 33858 16490 33872 16504
rect 33882 16490 33896 16504
rect 33426 16442 33440 16456
rect 33906 16442 33920 16456
rect 33402 16418 33416 16432
rect 33234 16370 33248 16384
rect 33258 16370 33272 16384
rect 33282 16370 33296 16384
rect 33306 16370 33320 16384
rect 33330 16370 33344 16384
rect 33354 16370 33368 16384
rect 33378 16370 33392 16384
rect 7722 16298 7736 16312
rect 7939 16310 7953 16324
rect 8519 16310 8533 16324
rect 33426 16394 33440 16408
rect 33450 16394 33464 16408
rect 33474 16394 33488 16408
rect 33498 16394 33512 16408
rect 33522 16394 33536 16408
rect 33546 16394 33560 16408
rect 33570 16394 33584 16408
rect 33594 16394 33608 16408
rect 33618 16394 33632 16408
rect 33642 16394 33656 16408
rect 33666 16394 33680 16408
rect 33690 16394 33704 16408
rect 33714 16394 33728 16408
rect 33738 16394 33752 16408
rect 33762 16394 33776 16408
rect 33786 16394 33800 16408
rect 33810 16394 33824 16408
rect 33834 16394 33848 16408
rect 33858 16394 33872 16408
rect 33882 16394 33896 16408
rect 33906 16394 33920 16408
rect 7746 16274 7760 16288
rect 7916 16286 7930 16300
rect 8553 16286 8567 16300
rect 9690 16298 9704 16312
rect 10482 16298 10496 16312
rect 11034 16298 11048 16312
rect 11250 16298 11264 16312
rect 11994 16298 12008 16312
rect 12162 16298 12176 16312
rect 12546 16298 12560 16312
rect 12738 16298 12752 16312
rect 12954 16298 12968 16312
rect 13698 16298 13712 16312
rect 13866 16298 13880 16312
rect 32370 16298 32384 16312
rect 32555 16298 32569 16312
rect 32603 16298 32617 16312
rect 32658 16298 32672 16312
rect 32730 16298 32744 16312
rect 33234 16298 33248 16312
rect 33258 16298 33272 16312
rect 33282 16298 33296 16312
rect 33306 16298 33320 16312
rect 33330 16298 33344 16312
rect 33354 16298 33368 16312
rect 33378 16298 33392 16312
rect 33402 16298 33416 16312
rect 33426 16298 33440 16312
rect 33474 16322 33488 16336
rect 33498 16322 33512 16336
rect 33522 16322 33536 16336
rect 33546 16322 33560 16336
rect 33570 16322 33584 16336
rect 33594 16322 33608 16336
rect 33618 16322 33632 16336
rect 33642 16322 33656 16336
rect 33666 16322 33680 16336
rect 33690 16322 33704 16336
rect 33714 16322 33728 16336
rect 33738 16322 33752 16336
rect 33762 16322 33776 16336
rect 33786 16322 33800 16336
rect 33810 16322 33824 16336
rect 33834 16322 33848 16336
rect 33858 16322 33872 16336
rect 33882 16322 33896 16336
rect 35462 16346 35476 16360
rect 35485 16322 35499 16336
rect 35509 16298 35523 16312
rect 6546 16250 6560 16264
rect 7458 16251 7472 16265
rect 7825 16264 7839 16278
rect 8592 16264 8606 16278
rect 7637 16248 7651 16262
rect 7893 16242 7907 16256
rect 8626 16242 8640 16256
rect 7871 16218 7885 16232
rect 8702 16218 8716 16232
rect 7801 16196 7815 16210
rect 8810 16194 8824 16208
rect 7848 16172 7862 16186
rect 7697 16150 7711 16164
rect 7722 16150 7736 16164
rect 7746 16150 7760 16164
rect 7778 16150 7792 16164
rect 8363 16172 8377 16186
rect 8458 16172 8472 16186
rect 8744 16127 8758 16141
rect 8854 16105 8868 16119
rect 10362 15818 10376 15832
rect 11274 15866 11288 15880
rect 12090 15866 12104 15880
rect 12930 15914 12944 15928
rect 13746 15938 13760 15952
rect 13794 15914 13808 15928
rect 14850 15914 14864 15928
rect 32397 16274 32411 16288
rect 23274 16250 23288 16264
rect 23466 16250 23480 16264
rect 23706 16250 23720 16264
rect 15450 15890 15464 15904
rect 17130 15891 17144 15905
rect 17191 15866 17205 15880
rect 18834 15818 18848 15832
rect 19686 15818 19700 15832
rect 8592 15793 8606 15807
rect 12018 15793 12032 15807
rect 12090 15794 12104 15808
rect 20575 15794 20589 15808
rect 8591 15769 8605 15783
rect 8854 15768 8868 15782
rect 10314 15771 10328 15785
rect 10362 15770 10376 15784
rect 17166 15769 17180 15783
rect 17190 15770 17204 15784
rect 21737 15770 21751 15784
rect 8553 15744 8567 15758
rect 14826 15746 14840 15760
rect 14850 15746 14864 15760
rect 8553 15720 8567 15734
rect 8744 15721 8758 15735
rect 12870 15722 12884 15736
rect 12930 15722 12944 15736
rect 21714 15722 21728 15736
rect 23106 15722 23120 15736
rect 23658 15746 23672 15760
rect 24786 15746 24800 15760
rect 8702 15698 8716 15712
rect 13722 15698 13736 15712
rect 13746 15698 13760 15712
rect 25602 15698 25616 15712
rect 7746 15678 7760 15692
rect 8520 15673 8534 15687
rect 15426 15674 15440 15688
rect 15450 15674 15464 15688
rect 23082 15674 23096 15688
rect 23106 15674 23120 15688
rect 25626 15674 25640 15688
rect 27282 15674 27296 15688
rect 7815 15654 7829 15668
rect 8520 15649 8534 15663
rect 8603 15649 8617 15663
rect 8627 15649 8641 15663
rect 13770 15650 13784 15664
rect 13794 15650 13808 15664
rect 24762 15650 24776 15664
rect 24786 15650 24800 15664
rect 27306 15650 27320 15664
rect 7583 15632 7597 15646
rect 7611 15632 7625 15646
rect 7635 15632 7649 15646
rect 7698 15632 7712 15646
rect 7746 15632 7760 15646
rect 7791 15632 7805 15646
rect 8238 15633 8252 15647
rect 8458 15633 8472 15647
rect 8811 15625 8825 15639
rect 10350 15625 10364 15639
rect 11274 15626 11288 15640
rect 8286 15610 8300 15624
rect 8411 15611 8425 15625
rect 20575 15626 20589 15640
rect 21737 15626 21751 15640
rect 23658 15626 23672 15640
rect 20538 15602 20552 15616
rect 23610 15602 23624 15616
rect 28602 15602 28616 15616
rect 6498 15482 6512 15496
rect 8262 15587 8276 15601
rect 8387 15588 8401 15602
rect 31410 16250 31424 16264
rect 31436 16250 31450 16264
rect 32509 16250 32523 16264
rect 32154 16226 32168 16240
rect 32373 16226 32387 16240
rect 31436 16202 31450 16216
rect 32397 16202 32411 16216
rect 32373 16178 32387 16192
rect 33858 16274 33872 16288
rect 33882 16274 33896 16288
rect 35533 16274 35547 16288
rect 33450 16250 33464 16264
rect 35557 16250 35571 16264
rect 35462 16226 35476 16240
rect 35581 16226 35595 16240
rect 33234 16202 33248 16216
rect 33258 16202 33272 16216
rect 33282 16202 33296 16216
rect 33306 16202 33320 16216
rect 33330 16202 33344 16216
rect 33354 16202 33368 16216
rect 33378 16202 33392 16216
rect 33402 16202 33416 16216
rect 33426 16202 33440 16216
rect 33450 16202 33464 16216
rect 33474 16202 33488 16216
rect 33498 16202 33512 16216
rect 33522 16202 33536 16216
rect 33546 16202 33560 16216
rect 33570 16202 33584 16216
rect 33594 16202 33608 16216
rect 33618 16202 33632 16216
rect 33642 16202 33656 16216
rect 33666 16202 33680 16216
rect 33690 16202 33704 16216
rect 33714 16202 33728 16216
rect 33738 16202 33752 16216
rect 33762 16202 33776 16216
rect 33786 16202 33800 16216
rect 33810 16202 33824 16216
rect 33834 16202 33848 16216
rect 35605 16202 35619 16216
rect 33450 15842 33464 15856
rect 35629 16178 35643 16192
rect 35653 16154 35667 16168
rect 35677 16130 35691 16144
rect 35701 16106 35715 16120
rect 35725 16082 35739 16096
rect 35749 16058 35763 16072
rect 35773 16034 35787 16048
rect 35797 16010 35811 16024
rect 35821 15986 35835 16000
rect 35845 15962 35859 15976
rect 35869 15938 35883 15952
rect 35893 15914 35907 15928
rect 35917 15890 35931 15904
rect 35941 15866 35955 15880
rect 35965 15842 35979 15856
rect 35989 15818 36003 15832
rect 36013 15794 36027 15808
rect 36037 15770 36051 15784
rect 36061 15770 36075 15784
rect 36109 15746 36123 15760
rect 36157 15722 36171 15736
rect 36402 15697 36416 15711
rect 36450 15674 36464 15688
rect 36474 15650 36488 15664
rect 29802 15602 29816 15616
rect 30306 15602 30320 15616
rect 30666 15602 30680 15616
rect 32322 15602 32336 15616
rect 32346 15602 32360 15616
rect 32634 15602 32648 15616
rect 36402 15602 36416 15616
rect 36450 15602 36464 15616
rect 36474 15602 36488 15616
rect 36450 15554 36464 15568
rect 36474 15554 36488 15568
rect 36402 15530 36416 15544
rect 36426 15530 36440 15544
rect 36062 15505 36076 15519
rect 7698 15487 7712 15501
rect 6498 15434 6512 15448
rect 36498 15482 36512 15496
rect 36426 15458 36440 15472
rect 36498 15434 36512 15448
rect 35454 15399 35468 15413
rect 36402 15386 36416 15400
rect 36450 15386 36464 15400
rect 36474 15386 36488 15400
rect 35533 15371 35547 15385
rect 7743 15332 7757 15346
rect 7863 15333 7877 15347
rect 35485 15333 35499 15347
rect 35509 15333 35523 15347
rect 35557 15333 35571 15347
rect 35581 15333 35595 15347
rect 35605 15333 35619 15347
rect 35629 15333 35643 15347
rect 35653 15333 35667 15347
rect 35677 15333 35691 15347
rect 35701 15333 35715 15347
rect 35725 15333 35739 15347
rect 35749 15333 35763 15347
rect 7863 15309 7877 15323
rect 7766 15273 7780 15287
rect 7791 15285 7805 15299
rect 7815 15285 7829 15299
rect 7838 15247 7852 15261
rect 36402 15338 36416 15352
rect 36450 15338 36464 15352
rect 36474 15338 36488 15352
rect 36402 15290 36416 15304
rect 36450 15290 36464 15304
rect 36474 15290 36488 15304
rect 35773 15261 35787 15275
rect 35701 15237 35715 15251
rect 35725 15237 35739 15251
rect 35749 15237 35763 15251
rect 35773 15237 35787 15251
rect 35557 15189 35571 15203
rect 35581 15189 35595 15203
rect 35605 15189 35619 15203
rect 35629 15189 35643 15203
rect 35653 15189 35667 15203
rect 35677 15189 35691 15203
rect 35749 15189 35763 15203
rect 35485 15165 35499 15179
rect 35509 15165 35523 15179
rect 36061 15165 36075 15179
rect 35461 15141 35475 15155
rect 35533 15141 35547 15155
rect 35461 15117 35475 15131
rect 36061 15117 36075 15131
rect 36109 15117 36123 15131
rect 36157 15117 36171 15131
rect 35461 15093 35475 15107
rect 35773 15093 35787 15107
rect 35965 15093 35979 15107
rect 35461 15069 35475 15083
rect 35461 15045 35475 15059
rect 35677 15045 35691 15059
rect 35701 15045 35715 15059
rect 35725 15045 35739 15059
rect 35485 15021 35499 15035
rect 35509 15021 35523 15035
rect 35533 15021 35547 15035
rect 35557 15021 35571 15035
rect 35581 15021 35595 15035
rect 35605 15021 35619 15035
rect 35629 15021 35643 15035
rect 35653 15021 35667 15035
rect 7791 11332 7805 11346
rect 7815 11332 7829 11346
rect 7839 11332 7853 11346
rect 7863 11308 7877 11322
rect 7791 11284 7805 11298
rect 7815 11284 7829 11298
rect 7863 11284 7877 11298
rect 7839 11260 7853 11274
rect 35557 11498 35571 11512
rect 35581 11498 35595 11512
rect 35605 11498 35619 11512
rect 35629 11498 35643 11512
rect 35653 11498 35667 11512
rect 35700 11499 35714 11513
rect 35797 15021 35811 15035
rect 35821 15021 35835 15035
rect 35845 15021 35859 15035
rect 35869 15021 35883 15035
rect 35893 15021 35907 15035
rect 35917 15021 35931 15035
rect 35941 15021 35955 15035
rect 35989 15021 36003 15035
rect 36013 15021 36027 15035
rect 36037 15021 36051 15035
rect 35725 11498 35739 11512
rect 35797 11498 35811 11512
rect 35821 11498 35835 11512
rect 35845 11498 35859 11512
rect 35869 11498 35883 11512
rect 35893 11498 35907 11512
rect 35917 11498 35931 11512
rect 35941 11498 35955 11512
rect 35989 11498 36003 11512
rect 36013 11498 36027 11512
rect 36037 11498 36051 11512
rect 36109 11498 36123 11512
rect 36157 11498 36171 11512
rect 36402 11498 36416 11512
rect 36450 11498 36464 11512
rect 36474 11498 36488 11512
rect 35557 11450 35571 11464
rect 35581 11450 35595 11464
rect 35605 11450 35619 11464
rect 35629 11450 35643 11464
rect 35653 11450 35667 11464
rect 35699 11451 35713 11465
rect 35485 8884 35499 8898
rect 35509 8884 35523 8898
rect 35557 8884 35571 8898
rect 35581 8884 35595 8898
rect 35461 8860 35475 8874
rect 35725 11450 35739 11464
rect 35797 11450 35811 11464
rect 35821 11450 35835 11464
rect 35845 11450 35859 11464
rect 35869 11450 35883 11464
rect 35893 11450 35907 11464
rect 35917 11450 35931 11464
rect 35941 11450 35955 11464
rect 35989 11450 36003 11464
rect 36013 11450 36027 11464
rect 36037 11450 36051 11464
rect 36109 11450 36123 11464
rect 36157 11450 36171 11464
rect 36402 11450 36416 11464
rect 36498 11450 36512 11464
rect 35697 8908 35711 8922
rect 35629 8860 35643 8874
rect 35653 8860 35667 8874
rect 35725 8858 35739 8872
rect 35461 8836 35475 8850
rect 35461 8812 35475 8826
rect 35653 8812 35667 8826
rect 35725 8810 35739 8824
rect 35485 8788 35499 8802
rect 35509 8788 35523 8802
rect 35557 8788 35571 8802
rect 35581 8788 35595 8802
rect 35629 8788 35643 8802
rect 35892 7499 35906 7513
rect 36450 11402 36464 11416
rect 36474 11402 36488 11416
rect 36498 11402 36512 11416
rect 36498 11306 36512 11320
rect 36498 11258 36512 11272
rect 36498 7394 36512 7408
rect 36498 7346 36512 7360
rect 35509 7250 35523 7264
rect 35557 7250 35571 7264
rect 35581 7250 35595 7264
rect 35629 7250 35643 7264
rect 35725 7250 35739 7264
rect 35821 7250 35835 7264
rect 35845 7250 35859 7264
rect 35869 7250 35883 7264
rect 35917 7250 35931 7264
rect 35941 7250 35955 7264
rect 35989 7250 36003 7264
rect 36013 7250 36027 7264
rect 36037 7250 36051 7264
rect 36109 7250 36123 7264
rect 36157 7250 36171 7264
rect 36498 7250 36512 7264
rect 35509 7202 35523 7216
rect 35557 7202 35571 7216
rect 35581 7202 35595 7216
rect 35629 7202 35643 7216
rect 35725 7202 35739 7216
rect 35821 7202 35835 7216
rect 35845 7202 35859 7216
rect 35869 7202 35883 7216
rect 35917 7202 35931 7216
rect 35941 7202 35955 7216
rect 35989 7202 36003 7216
rect 36013 7202 36027 7216
rect 36037 7202 36051 7216
rect 36109 7202 36123 7216
rect 36157 7202 36171 7216
rect 36498 7202 36512 7216
rect 7791 7082 7805 7096
rect 7815 7082 7829 7096
rect 7863 7091 7877 7105
rect 35509 7091 35523 7105
rect 35557 7091 35571 7105
rect 35581 7091 35595 7105
rect 35629 7091 35643 7105
rect 35725 7091 35739 7105
rect 35821 7091 35835 7105
rect 35845 7091 35859 7105
rect 7863 7058 7877 7072
rect 7791 7034 7805 7048
rect 35461 7043 35475 7057
rect 7815 7010 7829 7024
rect 35461 7019 35475 7033
rect 35821 7019 35835 7033
rect 35845 7019 35859 7033
rect 35461 6995 35475 7009
rect 35725 6995 35739 7009
rect 35581 6971 35595 6985
rect 35629 6971 35643 6985
rect 8310 6938 8324 6952
rect 8238 6890 8252 6904
rect 7376 6685 7390 6699
rect 7409 6685 7423 6699
rect 14514 6914 14528 6928
rect 15860 6914 15874 6928
rect 18042 6914 18056 6928
rect 22230 6913 22244 6927
rect 25482 6914 25496 6928
rect 25506 6914 25520 6928
rect 28590 6913 28604 6927
rect 31026 6914 31040 6928
rect 31050 6914 31064 6928
rect 35557 6890 35571 6904
rect 14514 6866 14528 6880
rect 15860 6866 15874 6880
rect 25098 6866 25112 6880
rect 25506 6866 25520 6880
rect 28482 6866 28496 6880
rect 31050 6866 31064 6880
rect 32154 6866 32168 6880
rect 35509 6866 35523 6880
rect 35629 6866 35643 6880
rect 22206 6841 22220 6855
rect 35874 6901 35888 6915
rect 35629 6818 35643 6832
rect 18042 6794 18056 6808
rect 25098 6794 25112 6808
rect 25482 6794 25496 6808
rect 31026 6770 31040 6784
rect 35940 6853 35954 6867
rect 35988 6830 36002 6844
rect 14370 6746 14384 6760
rect 14514 6746 14528 6760
rect 17898 6746 17912 6760
rect 18042 6746 18056 6760
rect 25098 6746 25112 6760
rect 15834 6721 15848 6735
rect 36036 6902 36050 6916
rect 36066 6854 36080 6868
rect 36035 6831 36049 6845
rect 14370 6698 14384 6712
rect 14514 6698 14528 6712
rect 17898 6698 17912 6712
rect 18042 6698 18056 6712
rect 34472 6647 34486 6661
rect 10986 6626 11000 6640
rect 14370 6626 14384 6640
rect 14514 6626 14528 6640
rect 17898 6626 17912 6640
rect 18042 6626 18056 6640
rect 24954 6626 24968 6640
rect 10986 6578 11000 6592
rect 14370 6578 14384 6592
rect 14514 6578 14528 6592
rect 17898 6578 17912 6592
rect 18042 6578 18056 6592
rect 24954 6578 24968 6592
rect 25098 6578 25112 6592
rect 28482 6578 28496 6592
rect 32010 6554 32024 6568
rect 32274 6578 32288 6592
rect 34537 6575 34551 6589
rect 36109 6578 36123 6592
rect 36156 6579 36170 6593
rect 32226 6554 32240 6568
rect 14370 6530 14384 6544
rect 14514 6530 14528 6544
rect 17898 6530 17912 6544
rect 18042 6530 18056 6544
rect 24954 6530 24968 6544
rect 25098 6530 25112 6544
rect 28482 6530 28496 6544
rect 28626 6530 28640 6544
rect 14370 6482 14384 6496
rect 14514 6482 14528 6496
rect 17898 6482 17912 6496
rect 18042 6482 18056 6496
rect 24954 6482 24968 6496
rect 25098 6482 25112 6496
rect 28482 6482 28496 6496
rect 28626 6482 28640 6496
rect 32010 6482 32024 6496
rect 32154 6482 32168 6496
rect 32226 6506 32240 6520
rect 32274 6530 32288 6544
rect 36109 6530 36123 6544
rect 34536 6504 34550 6518
rect 34472 6479 34486 6493
rect 36157 6477 36171 6491
<< metal2 >>
rect 7699 36325 7711 36362
rect 7723 36325 7735 36362
rect 10789 36348 10801 36437
rect 10867 36376 10879 36410
rect 14313 36348 14325 36440
rect 17875 36400 17887 36434
rect 18019 36232 18031 36434
rect 24931 36376 24943 36434
rect 25075 36352 25087 36434
rect 7248 36157 7361 36171
rect 7375 36157 8348 36171
rect 7248 36147 8348 36157
rect 7248 36133 7361 36147
rect 7375 36133 8348 36147
rect 7248 35971 8348 36133
rect 13099 36016 13111 36050
rect 14131 36016 14143 36146
rect 18019 36016 18031 36146
rect 6523 35461 6535 35498
rect 6499 31408 6511 31465
rect 6523 31408 6535 31514
rect 6499 27376 6511 27458
rect 6523 27376 6535 27458
rect 6547 27399 6559 27458
rect 6523 24240 6535 24274
rect 7248 24036 7448 35971
rect 7459 35896 7471 35930
rect 7652 35846 7664 35930
rect 7699 35848 7711 35930
rect 7723 35848 7735 35930
rect 8148 35824 8348 35971
rect 12907 35920 12919 35954
rect 13099 35920 13111 35954
rect 14131 35920 14143 35954
rect 18019 35920 18031 35954
rect 8364 35834 8370 35848
rect 11700 35834 11706 35848
rect 11940 35834 11946 35848
rect 12900 35834 12906 35848
rect 13092 35834 13098 35848
rect 14126 35834 14130 35848
rect 22123 35847 22135 35954
rect 22387 35847 22399 36050
rect 23107 35847 23119 36050
rect 24907 35847 24919 36146
rect 25099 35847 25111 36194
rect 25171 35847 25183 35954
rect 25267 35847 25279 36146
rect 28459 35896 28471 36434
rect 28603 35968 28615 36434
rect 31939 36328 31951 36410
rect 31987 36277 31999 36434
rect 32131 36328 32143 36434
rect 32938 36376 32950 36436
rect 32964 36278 33948 36418
rect 31987 36265 32023 36277
rect 31987 35968 31999 36218
rect 32011 35968 32023 36265
rect 32978 36264 33948 36278
rect 32964 36218 33948 36264
rect 32937 35896 32949 36218
rect 22117 35835 22135 35847
rect 22381 35835 22399 35847
rect 23101 35835 23119 35847
rect 24900 35835 24919 35847
rect 25092 35835 25111 35847
rect 25164 35835 25183 35847
rect 25260 35835 25279 35847
rect 8364 35824 8376 35834
rect 11700 35824 11712 35834
rect 11940 35824 11952 35834
rect 12900 35824 12912 35834
rect 13092 35824 13104 35834
rect 14126 35824 14138 35834
rect 22117 35824 22129 35835
rect 22381 35824 22393 35835
rect 23101 35824 23113 35835
rect 24900 35824 24912 35835
rect 25092 35824 25104 35835
rect 25164 35824 25176 35835
rect 25260 35824 25272 35835
rect 32964 35824 33164 36218
rect 33235 35848 33247 36194
rect 33259 35848 33271 36170
rect 33283 35848 33295 36122
rect 33331 35848 33343 36002
rect 33355 35848 33367 36098
rect 33379 35848 33391 35930
rect 33403 35848 33415 36050
rect 33427 35848 33439 36146
rect 33451 35848 33463 36050
rect 33475 35848 33487 36051
rect 33499 35848 33511 36026
rect 33523 35848 33535 35978
rect 33547 35848 33559 35930
rect 33571 35848 33583 36074
rect 33595 35968 33607 36050
rect 33643 36003 33724 36015
rect 33643 35896 33655 36003
rect 33667 35896 33679 35978
rect 33691 35896 33703 35954
rect 7459 35464 7471 35498
rect 33748 34499 33948 36218
rect 36499 35656 36511 35690
rect 36499 35512 36511 35546
rect 33748 34485 33934 34499
rect 33235 33040 33247 33146
rect 33259 33040 33271 33146
rect 33283 33040 33295 33146
rect 33331 33040 33343 33146
rect 33355 33040 33367 33146
rect 33379 33040 33391 33146
rect 33403 33040 33415 33146
rect 33427 33040 33439 33146
rect 33451 33040 33463 33146
rect 33475 33040 33487 33146
rect 33499 33040 33511 33146
rect 33523 33040 33535 33146
rect 33547 33040 33559 33146
rect 33571 33040 33583 33146
rect 33595 33040 33607 33146
rect 33619 33040 33631 33146
rect 33643 33040 33655 33146
rect 33667 33040 33679 33146
rect 33691 33112 33703 33146
rect 33748 32498 33948 34485
rect 33748 32484 33934 32498
rect 33235 31936 33247 32042
rect 33259 31936 33271 32042
rect 33283 31936 33295 32042
rect 33331 31936 33343 32042
rect 33355 31936 33367 32042
rect 33379 31936 33391 32042
rect 33403 31936 33415 32042
rect 33427 31936 33439 32042
rect 33451 31936 33463 32042
rect 33475 31936 33487 32042
rect 33499 31936 33511 32042
rect 33523 31936 33535 32042
rect 33547 31936 33559 32042
rect 33571 31936 33583 32042
rect 33595 31936 33607 32042
rect 33619 31936 33631 32042
rect 33643 32008 33655 32042
rect 33235 30808 33247 30914
rect 33259 30808 33271 30914
rect 33283 30808 33295 30914
rect 33331 30808 33343 30914
rect 33355 30808 33367 30914
rect 33379 30808 33391 30914
rect 33403 30808 33415 30914
rect 33427 30808 33439 30914
rect 33451 30808 33463 30914
rect 33475 30808 33487 30914
rect 33499 30808 33511 30914
rect 33523 30808 33535 30914
rect 33547 30808 33559 30914
rect 33571 30808 33583 30914
rect 33595 30880 33607 30914
rect 33748 30498 33948 32484
rect 36475 31624 36487 31658
rect 36499 31624 36511 31658
rect 36427 31504 36439 31538
rect 36451 31504 36463 31538
rect 36499 31480 36511 31514
rect 33748 30484 33934 30498
rect 33235 29704 33247 29810
rect 33259 29704 33271 29810
rect 33283 29704 33295 29810
rect 33331 29704 33343 29810
rect 33355 29704 33367 29810
rect 33379 29704 33391 29810
rect 33403 29704 33415 29810
rect 33427 29704 33439 29810
rect 33451 29704 33463 29810
rect 33475 29704 33487 29810
rect 33499 29704 33511 29810
rect 33523 29704 33535 29810
rect 33547 29776 33559 29810
rect 33235 28600 33247 28706
rect 33259 28600 33271 28706
rect 33283 28600 33295 28706
rect 33331 28600 33343 28706
rect 33355 28600 33367 28706
rect 33379 28600 33391 28706
rect 33403 28600 33415 28706
rect 33427 28600 33439 28706
rect 33451 28600 33463 28706
rect 33475 28600 33487 28706
rect 33499 28600 33511 28706
rect 33523 28600 33535 28706
rect 33748 28498 33948 30484
rect 33748 28484 33934 28498
rect 33235 27496 33247 27578
rect 33259 27496 33271 27578
rect 33283 27496 33295 27578
rect 33331 27496 33343 27578
rect 33355 27496 33367 27578
rect 33379 27496 33391 27578
rect 33403 27496 33415 27578
rect 33427 27496 33439 27578
rect 33451 27496 33463 27578
rect 33475 27496 33487 27578
rect 33499 27496 33511 27578
rect 33523 27496 33535 27578
rect 7459 27424 7471 27458
rect 33748 26897 33948 28484
rect 36451 27616 36463 27650
rect 36499 27592 36511 27626
rect 36475 27448 36487 27482
rect 36499 27448 36511 27482
rect 33748 26883 33934 26897
rect 33235 26368 33247 26474
rect 33259 26368 33271 26474
rect 33283 26368 33295 26474
rect 33331 26368 33343 26474
rect 33355 26368 33367 26474
rect 33379 26368 33391 26474
rect 33403 26368 33415 26474
rect 33427 26368 33439 26474
rect 33451 26368 33463 26474
rect 33475 26368 33487 26474
rect 33499 26368 33511 26474
rect 33523 26368 33535 26474
rect 33235 25336 33247 25370
rect 33259 25288 33271 25322
rect 33283 25288 33295 25394
rect 33331 25288 33343 25394
rect 33355 25288 33367 25394
rect 33379 25288 33391 25394
rect 33403 25288 33415 25394
rect 33427 25288 33439 25394
rect 33451 25288 33463 25394
rect 33475 25288 33487 25394
rect 33499 25288 33511 25394
rect 33523 25288 33535 25394
rect 33547 25288 33559 25322
rect 33748 24898 33948 26883
rect 33748 24884 33934 24898
rect 33235 24160 33247 24242
rect 33259 24160 33271 24194
rect 33283 24160 33295 24266
rect 33331 24184 33343 24266
rect 33355 24184 33367 24266
rect 33379 24184 33391 24266
rect 33403 24184 33415 24266
rect 33427 24184 33439 24266
rect 33451 24184 33463 24266
rect 33475 24184 33487 24266
rect 33499 24184 33511 24266
rect 33523 24184 33535 24266
rect 33547 24184 33559 24266
rect 33571 24184 33583 24266
rect 33595 24184 33607 24218
rect 6450 23836 7448 24036
rect 33748 24056 33948 24884
rect 33748 24040 34480 24056
rect 34496 24040 36550 24056
rect 33748 23856 36550 24040
rect 34099 23492 34699 23493
rect 6450 22886 7423 23486
rect 33235 23032 33247 23138
rect 33259 23032 33271 23138
rect 33283 23104 33295 23138
rect 33307 23056 33319 23138
rect 33331 23056 33343 23138
rect 33355 23056 33367 23138
rect 33379 23056 33391 23138
rect 33403 23056 33415 23138
rect 33427 23056 33439 23090
rect 33451 23056 33463 23162
rect 33475 23056 33487 23162
rect 33499 23056 33511 23162
rect 33523 23056 33535 23162
rect 33547 23056 33559 23162
rect 33571 23056 33583 23162
rect 33595 23056 33607 23162
rect 33619 23056 33631 23090
rect 6523 19504 6535 19538
rect 6547 19504 6559 19538
rect 6547 16264 6559 16322
rect 6823 16120 7423 22886
rect 34099 22892 36552 23492
rect 33235 21928 33247 22034
rect 33259 21928 33271 22034
rect 33283 21928 33295 22034
rect 33307 21928 33319 22034
rect 33331 21928 33343 22034
rect 33379 22024 33391 22058
rect 33403 22024 33415 22058
rect 33427 22024 33439 22058
rect 33451 22024 33463 22058
rect 33355 21928 33367 21962
rect 33379 21928 33391 21962
rect 33403 21928 33415 21962
rect 33427 21928 33439 21962
rect 33475 21952 33487 22058
rect 33499 21952 33511 22058
rect 33523 21952 33535 22058
rect 33547 21952 33559 22058
rect 33571 21952 33583 22058
rect 33595 21952 33607 22058
rect 33619 21952 33631 22058
rect 33643 21952 33655 22058
rect 33667 21952 33679 21986
rect 33235 20824 33247 20930
rect 33259 20824 33271 20930
rect 33283 20824 33295 20930
rect 33307 20824 33319 20930
rect 33331 20824 33343 20930
rect 33355 20824 33367 20930
rect 33379 20824 33391 20930
rect 33427 20920 33439 20954
rect 33451 20920 33463 20954
rect 33475 20920 33487 20954
rect 33499 20920 33511 20954
rect 33403 20824 33415 20858
rect 33427 20824 33439 20858
rect 33451 20824 33463 20858
rect 33475 20824 33487 20858
rect 33523 20848 33535 20954
rect 33547 20848 33559 20954
rect 33571 20848 33583 20954
rect 33595 20848 33607 20954
rect 33619 20848 33631 20954
rect 33643 20848 33655 20954
rect 33667 20848 33679 20954
rect 33691 20848 33703 20954
rect 33715 20848 33727 20882
rect 33235 19720 33247 19802
rect 33259 19720 33271 19802
rect 33283 19720 33295 19802
rect 33307 19720 33319 19802
rect 33331 19720 33343 19754
rect 33355 19720 33367 19826
rect 33379 19720 33391 19826
rect 33403 19720 33415 19826
rect 33427 19720 33439 19826
rect 33451 19720 33463 19826
rect 33475 19720 33487 19826
rect 33499 19720 33511 19826
rect 33523 19792 33535 19826
rect 33547 19744 33559 19826
rect 33571 19744 33583 19826
rect 33595 19744 33607 19826
rect 33619 19744 33631 19826
rect 33643 19744 33655 19826
rect 33667 19744 33679 19826
rect 33691 19744 33703 19826
rect 33715 19744 33727 19826
rect 33739 19744 33751 19826
rect 33763 19744 33775 19778
rect 33235 18592 33247 18698
rect 33259 18592 33271 18698
rect 33283 18592 33295 18698
rect 33307 18592 33319 18698
rect 33331 18592 33343 18698
rect 33355 18592 33367 18698
rect 33379 18664 33391 18698
rect 33403 18616 33415 18698
rect 33427 18616 33439 18698
rect 33451 18616 33463 18698
rect 33475 18616 33487 18698
rect 33499 18616 33511 18698
rect 33523 18616 33535 18698
rect 33547 18616 33559 18698
rect 33571 18616 33583 18698
rect 33595 18616 33607 18698
rect 33619 18616 33631 18698
rect 33643 18616 33655 18698
rect 33667 18616 33679 18698
rect 33691 18616 33703 18698
rect 33715 18616 33727 18698
rect 33739 18616 33751 18698
rect 33763 18616 33775 18698
rect 33787 18616 33799 18698
rect 33811 18616 33823 18650
rect 33235 17488 33247 17594
rect 33259 17488 33271 17594
rect 33283 17488 33295 17594
rect 33307 17488 33319 17594
rect 33331 17488 33343 17594
rect 33355 17488 33367 17594
rect 33379 17488 33391 17594
rect 33403 17488 33415 17594
rect 33427 17488 33439 17594
rect 33451 17488 33463 17594
rect 33475 17488 33487 17594
rect 33499 17488 33511 17594
rect 33523 17488 33535 17594
rect 33547 17488 33559 17594
rect 33571 17488 33583 17594
rect 33595 17560 33607 17594
rect 33619 17512 33631 17594
rect 33643 17512 33655 17594
rect 33667 17512 33679 17594
rect 33691 17512 33703 17594
rect 33715 17512 33727 17594
rect 33739 17512 33751 17594
rect 33763 17512 33775 17594
rect 33787 17512 33799 17594
rect 33811 17512 33823 17594
rect 33835 17512 33847 17594
rect 33859 17512 33871 17546
rect 34099 16603 34699 22892
rect 33235 16384 33247 16466
rect 33259 16384 33271 16466
rect 33283 16384 33295 16466
rect 33307 16384 33319 16466
rect 33331 16384 33343 16466
rect 33355 16384 33367 16466
rect 33379 16384 33391 16466
rect 33403 16432 33415 16466
rect 33427 16408 33439 16442
rect 33451 16408 33463 16490
rect 33475 16408 33487 16490
rect 33499 16408 33511 16490
rect 33523 16408 33535 16490
rect 33547 16408 33559 16490
rect 33571 16408 33583 16490
rect 33595 16408 33607 16490
rect 33619 16408 33631 16490
rect 33643 16408 33655 16490
rect 33667 16408 33679 16490
rect 33691 16408 33703 16490
rect 33715 16408 33727 16490
rect 33739 16408 33751 16490
rect 33763 16408 33775 16490
rect 33787 16408 33799 16490
rect 33811 16408 33823 16490
rect 33835 16408 33847 16490
rect 33859 16408 33871 16490
rect 33883 16408 33895 16490
rect 33907 16408 33919 16442
rect 34099 16370 36389 16603
rect 7459 16265 7471 16322
rect 7637 16262 7649 16322
rect 7698 16164 7710 16346
rect 7723 16164 7735 16298
rect 7747 16164 7759 16274
rect 7779 16164 7791 16334
rect 7802 16210 7814 16334
rect 7825 16278 7837 16334
rect 7848 16321 7861 16334
rect 7849 16186 7861 16321
rect 7871 16232 7883 16334
rect 7894 16256 7906 16334
rect 7917 16300 7929 16334
rect 7940 16324 7952 16334
rect 8148 16120 8348 16334
rect 8364 16186 8376 16334
rect 6823 15720 8348 16120
rect 6823 15520 7544 15720
rect 7747 15646 7759 15678
rect 6499 15448 6511 15482
rect 7344 6885 7544 15520
rect 7584 15260 7596 15632
rect 7612 15287 7624 15632
rect 7636 15344 7648 15632
rect 7699 15501 7711 15632
rect 7636 15332 7743 15344
rect 7792 15299 7804 15632
rect 7816 15299 7828 15654
rect 8023 15429 8223 15720
rect 8239 15429 8251 15633
rect 8263 15429 8275 15587
rect 8287 15429 8299 15610
rect 8388 15602 8400 16334
rect 8412 15625 8424 16334
rect 8436 15578 8448 16334
rect 8459 15647 8471 16172
rect 8521 15687 8533 16310
rect 9684 16312 9696 16334
rect 10476 16312 10488 16334
rect 11028 16312 11040 16334
rect 11244 16312 11256 16334
rect 11988 16312 12000 16334
rect 12156 16312 12168 16334
rect 12540 16312 12552 16334
rect 12732 16312 12744 16334
rect 12948 16312 12960 16334
rect 13692 16312 13704 16334
rect 13860 16312 13872 16334
rect 9684 16298 9690 16312
rect 10476 16298 10482 16312
rect 11028 16298 11034 16312
rect 11244 16298 11250 16312
rect 11988 16298 11994 16312
rect 12156 16298 12162 16312
rect 12540 16298 12546 16312
rect 12732 16298 12738 16312
rect 12948 16298 12954 16312
rect 13692 16298 13698 16312
rect 13860 16298 13866 16312
rect 23268 16311 23280 16334
rect 23460 16311 23472 16334
rect 23700 16311 23712 16334
rect 31404 16311 31416 16334
rect 32148 16311 32160 16334
rect 32364 16312 32376 16334
rect 23268 16299 23287 16311
rect 23460 16299 23479 16311
rect 23700 16299 23719 16311
rect 31404 16299 31423 16311
rect 32148 16299 32167 16311
rect 8554 15758 8566 16286
rect 23275 16264 23287 16299
rect 23467 16264 23479 16299
rect 23707 16264 23719 16299
rect 31411 16264 31423 16299
rect 8593 15807 8605 16264
rect 8628 15663 8640 16242
rect 8703 15712 8715 16218
rect 31437 16216 31449 16250
rect 32155 16240 32167 16299
rect 32364 16298 32370 16312
rect 8745 15735 8757 16127
rect 8812 15639 8824 16194
rect 32374 16192 32386 16226
rect 32398 16216 32410 16274
rect 32510 16264 32522 16334
rect 32556 16312 32568 16334
rect 32604 16312 32616 16334
rect 32652 16312 32664 16334
rect 32724 16312 32736 16334
rect 32652 16298 32658 16312
rect 32724 16298 32730 16312
rect 32964 16146 33164 16334
rect 33235 16216 33247 16298
rect 33259 16216 33271 16298
rect 33283 16216 33295 16298
rect 33307 16216 33319 16298
rect 33331 16216 33343 16298
rect 33355 16216 33367 16298
rect 33379 16216 33391 16298
rect 33403 16216 33415 16298
rect 33427 16216 33439 16298
rect 33451 16216 33463 16250
rect 33475 16216 33487 16322
rect 33499 16216 33511 16322
rect 33523 16216 33535 16322
rect 33547 16216 33559 16322
rect 33571 16216 33583 16322
rect 33595 16216 33607 16322
rect 33619 16216 33631 16322
rect 33643 16216 33655 16322
rect 33667 16216 33679 16322
rect 33691 16216 33703 16322
rect 33715 16216 33727 16322
rect 33739 16216 33751 16322
rect 33763 16216 33775 16322
rect 33787 16216 33799 16322
rect 33811 16216 33823 16322
rect 33835 16216 33847 16322
rect 33859 16288 33871 16322
rect 33883 16288 33895 16322
rect 34099 16146 34499 16370
rect 35463 16240 35475 16346
rect 8855 15782 8867 16105
rect 32964 15947 34499 16146
rect 32964 15946 33930 15947
rect 10363 15784 10375 15818
rect 8311 15566 8448 15578
rect 8311 15429 8323 15566
rect 10315 15429 10327 15771
rect 11275 15640 11287 15866
rect 12091 15808 12103 15866
rect 10351 15429 10363 15625
rect 12019 15429 12031 15793
rect 12931 15736 12943 15914
rect 12871 15429 12883 15722
rect 13747 15712 13759 15938
rect 13723 15429 13735 15698
rect 13795 15664 13807 15914
rect 14851 15760 14863 15914
rect 13771 15615 13783 15650
rect 13771 15603 14191 15615
rect 14179 15429 14191 15603
rect 14827 15598 14839 15746
rect 15451 15688 15463 15890
rect 15427 15620 15439 15674
rect 15427 15608 15475 15620
rect 14827 15586 15439 15598
rect 15427 15429 15439 15586
rect 15463 15429 15475 15608
rect 17131 15429 17143 15891
rect 17192 15784 17204 15866
rect 17167 15429 17179 15769
rect 18835 15429 18847 15818
rect 19687 15429 19699 15818
rect 20576 15640 20588 15794
rect 20539 15429 20551 15602
rect 20575 15429 20587 15626
rect 21715 15429 21727 15722
rect 21738 15640 21750 15770
rect 23107 15688 23119 15722
rect 23083 15429 23095 15674
rect 23659 15640 23671 15746
rect 24787 15664 24799 15746
rect 23611 15429 23623 15602
rect 24763 15429 24775 15650
rect 25603 15429 25615 15698
rect 25627 15429 25639 15674
rect 27283 15429 27295 15674
rect 27307 15429 27319 15650
rect 32648 15602 32652 15616
rect 33451 15614 33463 15842
rect 34099 15747 35272 15947
rect 33451 15602 34039 15614
rect 28603 15429 28615 15602
rect 29803 15429 29815 15602
rect 30307 15429 30319 15602
rect 30667 15429 30679 15602
rect 32323 15429 32335 15602
rect 32347 15429 32359 15602
rect 32640 15464 32652 15602
rect 32640 15452 33199 15464
rect 33187 15429 33199 15452
rect 34027 15429 34039 15602
rect 35070 15573 35272 15747
rect 35071 15429 35271 15573
rect 7877 15334 7900 15346
rect 7877 15310 7900 15322
rect 7612 15275 7766 15287
rect 35455 15283 35467 15399
rect 35486 15347 35498 16322
rect 35510 15347 35522 16298
rect 35534 15385 35546 16274
rect 35558 15347 35570 16250
rect 35582 15347 35594 16226
rect 35606 15347 35618 16202
rect 35630 15347 35642 16178
rect 35654 15347 35666 16154
rect 35678 15347 35690 16130
rect 35702 15347 35714 16106
rect 35726 15347 35738 16082
rect 35750 15347 35762 16058
rect 35455 15271 35546 15283
rect 35774 15275 35786 16034
rect 7584 15248 7838 15260
rect 35429 15142 35461 15154
rect 35429 15118 35461 15130
rect 35429 15094 35461 15106
rect 35429 15070 35461 15082
rect 35429 15046 35461 15058
rect 35486 15035 35498 15165
rect 35510 15035 35522 15165
rect 35534 15155 35546 15271
rect 35534 15035 35546 15141
rect 35558 15035 35570 15189
rect 35582 15035 35594 15189
rect 35606 15035 35618 15189
rect 35630 15035 35642 15189
rect 35654 15035 35666 15189
rect 35678 15059 35690 15189
rect 35702 15059 35714 15237
rect 35726 15059 35738 15237
rect 35750 15203 35762 15237
rect 35774 15107 35786 15237
rect 35798 15035 35810 16010
rect 35822 15035 35834 15986
rect 35846 15035 35858 15962
rect 35870 15035 35882 15938
rect 35894 15035 35906 15914
rect 35918 15035 35930 15890
rect 35942 15035 35954 15866
rect 35966 15107 35978 15842
rect 35990 15035 36002 15818
rect 36014 15035 36026 15794
rect 36038 15035 36050 15770
rect 36062 15519 36074 15770
rect 36062 15131 36074 15165
rect 36110 15131 36122 15746
rect 36158 15131 36170 15722
rect 35558 11464 35570 11498
rect 35582 11464 35594 11498
rect 35606 11464 35618 11498
rect 35630 11464 35642 11498
rect 35654 11464 35666 11498
rect 35700 11465 35712 11499
rect 35726 11464 35738 11498
rect 35798 11464 35810 11498
rect 35822 11464 35834 11498
rect 35846 11464 35858 11498
rect 35870 11464 35882 11498
rect 35894 11464 35906 11498
rect 35918 11464 35930 11498
rect 35942 11464 35954 11498
rect 35990 11464 36002 11498
rect 36014 11464 36026 11498
rect 36038 11464 36050 11498
rect 36110 11464 36122 11498
rect 36158 11464 36170 11498
rect 7792 11298 7804 11332
rect 7816 11298 7828 11332
rect 7840 11274 7852 11332
rect 7877 11309 7900 11321
rect 7877 11285 7900 11297
rect 35429 8909 35697 8921
rect 35429 8861 35461 8873
rect 35429 8837 35461 8849
rect 35429 8813 35461 8825
rect 35486 8802 35498 8884
rect 35510 8802 35522 8884
rect 35558 8802 35570 8884
rect 35582 8802 35594 8884
rect 35630 8802 35642 8860
rect 35654 8826 35666 8860
rect 35726 8824 35738 8858
rect 35429 7500 35892 7512
rect 35510 7216 35522 7250
rect 35558 7216 35570 7250
rect 35582 7216 35594 7250
rect 35630 7216 35642 7250
rect 35726 7216 35738 7250
rect 35822 7216 35834 7250
rect 35846 7216 35858 7250
rect 35870 7216 35882 7250
rect 35918 7216 35930 7250
rect 35942 7216 35954 7250
rect 35990 7216 36002 7250
rect 36014 7216 36026 7250
rect 36038 7216 36050 7250
rect 36110 7216 36122 7250
rect 36158 7216 36170 7250
rect 7877 7092 7900 7104
rect 7792 7048 7804 7082
rect 7816 7024 7828 7082
rect 7863 7072 7900 7080
rect 7877 7068 7900 7072
rect 35429 7044 35461 7056
rect 35429 7020 35461 7032
rect 35429 6996 35461 7008
rect 8025 6885 8225 6985
rect 8239 6904 8251 6985
rect 8311 6952 8323 6985
rect 7344 6699 8225 6885
rect 14515 6880 14527 6914
rect 14371 6712 14383 6746
rect 14515 6712 14527 6746
rect 15835 6735 15847 6985
rect 15861 6880 15873 6914
rect 18043 6808 18055 6914
rect 22207 6855 22219 6985
rect 22231 6927 22243 6985
rect 28591 6927 28603 6985
rect 25099 6808 25111 6866
rect 25483 6808 25495 6914
rect 25507 6880 25519 6914
rect 17899 6712 17911 6746
rect 18043 6712 18055 6746
rect 7344 6685 7376 6699
rect 7390 6685 7409 6699
rect 7423 6685 8225 6699
rect 10987 6592 10999 6626
rect 14371 6592 14383 6626
rect 14515 6592 14527 6626
rect 17899 6592 17911 6626
rect 18043 6592 18055 6626
rect 24955 6592 24967 6626
rect 25099 6592 25111 6746
rect 28483 6592 28495 6866
rect 31027 6784 31039 6914
rect 31051 6880 31063 6914
rect 14371 6496 14383 6530
rect 14515 6496 14527 6530
rect 17899 6496 17911 6530
rect 18043 6496 18055 6530
rect 24955 6496 24967 6530
rect 25099 6496 25111 6530
rect 28483 6496 28495 6530
rect 28627 6496 28639 6530
rect 32011 6496 32023 6554
rect 32155 6496 32167 6866
rect 35071 6807 35271 6985
rect 35510 6880 35522 7091
rect 35558 6904 35570 7091
rect 35582 6985 35594 7091
rect 35630 6985 35642 7091
rect 35726 7009 35738 7091
rect 35822 7033 35834 7091
rect 35846 7033 35858 7091
rect 35888 6902 36036 6914
rect 35630 6832 35642 6866
rect 35954 6855 36066 6867
rect 36002 6832 36035 6844
rect 36189 6807 36389 16370
rect 36403 15616 36415 15697
rect 36451 15616 36463 15674
rect 36475 15616 36487 15650
rect 36403 15400 36415 15530
rect 36427 15472 36439 15530
rect 36451 15400 36463 15554
rect 36475 15400 36487 15554
rect 36499 15448 36511 15482
rect 36403 15304 36415 15338
rect 36451 15304 36463 15338
rect 36475 15304 36487 15338
rect 36403 11464 36415 11498
rect 36451 11416 36463 11498
rect 36475 11416 36487 11498
rect 36499 11416 36511 11450
rect 36499 11272 36511 11306
rect 36499 7360 36511 7394
rect 36499 7216 36511 7250
rect 32227 6520 32239 6554
rect 32275 6544 32287 6578
rect 34473 6493 34485 6647
rect 35071 6607 36389 6807
rect 34537 6518 34549 6575
rect 36110 6544 36122 6578
rect 36158 6491 36170 6579
<< metal4 >>
rect 6616 41276 8176 42836
rect 10142 41276 11702 42836
rect 13668 41276 15228 42836
rect 17194 41276 18754 42836
rect 20720 41276 22280 42836
rect 24246 41276 25806 42836
rect 27772 41276 29332 42836
rect 31298 41276 32858 42836
rect 34824 41276 36384 42836
rect 78 34824 1638 36384
rect 41362 34824 42922 36384
rect 78 30782 1638 32342
rect 41362 30782 42922 32342
rect 78 26740 1638 28300
rect 41362 26740 42922 28300
rect 78 22698 1638 24258
rect 41422 22758 42862 24198
rect 78 18656 1638 20216
rect 41362 18656 42922 20216
rect 78 14614 1638 16174
rect 41362 14614 42922 16174
rect 78 10572 1638 12132
rect 41362 10572 42922 12132
rect 78 6530 1638 8090
rect 41362 6530 42922 8090
rect 6616 78 8176 1638
rect 10142 78 11702 1638
rect 13668 78 15228 1638
rect 17194 78 18754 1638
rect 20720 78 22280 1638
rect 24246 78 25806 1638
rect 27772 78 29332 1638
rect 31298 78 32858 1638
rect 34824 78 36384 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 0 -1 0 42914
box 0 0 6450 6450
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 6536 1 0 36464
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 8256 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 8342 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 8428 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 8514 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 8600 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 8686 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 8772 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 8858 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 8944 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 9030 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 9116 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 9202 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 9288 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 9374 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 9460 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 9546 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 9632 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 9718 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 9804 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 9890 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 9976 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 10062 1 0 36464
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 11782 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 11868 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 11954 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 12040 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 12126 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 12212 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 12298 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 12384 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 12470 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 12556 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 12642 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 12728 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 12814 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 12900 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 12986 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 13072 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 13158 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 13244 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 13330 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 13416 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 13502 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 13588 1 0 36464
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 15308 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 15394 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 15480 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 15566 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 15652 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 15738 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 15824 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 15910 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 15996 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 16082 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 16168 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 16254 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 0 -1 16340 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 0 -1 16426 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 0 -1 16512 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 0 -1 16598 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 0 -1 16684 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 0 -1 16770 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 0 -1 16856 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 0 -1 16942 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 0 -1 17028 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 0 -1 17114 1 0 36464
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 18834 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 0 -1 18920 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 0 -1 19006 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 0 -1 19092 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 0 -1 19178 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 0 -1 19264 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 0 -1 19350 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 0 -1 19436 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 0 -1 19522 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 0 -1 19608 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 0 -1 19694 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 0 -1 19780 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 0 -1 19866 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 0 -1 19952 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 0 -1 20038 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 0 -1 20124 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 0 -1 20210 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 0 -1 20296 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 0 -1 20382 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 0 -1 20468 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 0 -1 20554 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 0 -1 20640 1 0 36464
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 22360 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 0 -1 22446 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 0 -1 22532 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 0 -1 22618 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 0 -1 22704 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 0 -1 22790 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 0 -1 22876 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 0 -1 22962 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 0 -1 23048 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 0 -1 23134 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 0 -1 23220 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 0 -1 23306 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 0 -1 23392 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 0 -1 23478 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 0 -1 23564 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 0 -1 23650 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 0 -1 23736 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 0 -1 23822 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 0 -1 23908 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 0 -1 23994 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 0 -1 24080 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 0 -1 24166 1 0 36464
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 25886 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 0 -1 25972 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 0 -1 26058 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 0 -1 26144 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 0 -1 26230 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 0 -1 26316 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 0 -1 26402 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 0 -1 26488 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 0 -1 26574 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 0 -1 26660 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 0 -1 26746 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 0 -1 26832 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 0 -1 26918 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 0 -1 27004 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 0 -1 27090 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 0 -1 27176 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 0 -1 27262 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 0 -1 27348 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 0 -1 27434 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 0 -1 27520 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 0 -1 27606 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 0 -1 27692 1 0 36464
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 29412 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 0 -1 29498 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 0 -1 29584 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 0 -1 29670 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 0 -1 29756 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 0 -1 29842 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 0 -1 29928 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 0 -1 30014 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 0 -1 30100 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 0 -1 30186 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 0 -1 30272 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 0 -1 30358 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 0 -1 30444 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 0 -1 30530 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 0 -1 30616 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 0 -1 30702 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 0 -1 30788 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 0 -1 30874 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 0 -1 30960 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 0 -1 31046 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 0 -1 31132 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 0 -1 31218 1 0 36464
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 32938 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 0 -1 33024 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 0 -1 33110 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 0 -1 33196 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 0 -1 33282 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 0 -1 33368 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 0 -1 33454 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 0 -1 33540 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 0 -1 33626 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 0 -1 33712 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 0 -1 33798 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 0 -1 33884 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 0 -1 33970 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 0 -1 34056 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 0 -1 34142 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 0 -1 34228 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 0 -1 34314 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 0 -1 34400 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 0 -1 34486 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 0 -1 34572 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 0 -1 34658 1 0 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 0 -1 34744 1 0 36464
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 36464 1 0 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 0 -1 36550 1 0 36464
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 43000 0 -1 42914
box 0 0 6450 6450
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 6450 0 -1 36464
box 0 0 6450 1720
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform -1 0 6450 0 -1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform -1 0 6450 0 -1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform -1 0 6450 0 -1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform -1 0 6450 0 -1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform -1 0 6450 0 -1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform -1 0 6450 0 -1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform -1 0 6450 0 -1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform -1 0 6450 0 -1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform -1 0 6450 0 -1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform -1 0 6450 0 -1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform -1 0 6450 0 -1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform -1 0 6450 0 -1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform -1 0 6450 0 -1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform -1 0 6450 0 -1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform -1 0 6450 0 -1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform -1 0 6450 0 -1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform -1 0 6450 0 -1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform -1 0 6450 0 -1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform -1 0 6450 0 -1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform -1 0 6450 0 -1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform -1 0 6450 0 -1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform -1 0 6450 0 -1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform -1 0 6450 0 -1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform -1 0 6450 0 -1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform -1 0 6450 0 -1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform -1 0 6450 0 -1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform -1 0 6450 0 -1 32508
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 6450 0 -1 32422
box 0 0 6450 1720
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform -1 0 6450 0 -1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform -1 0 6450 0 -1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform -1 0 6450 0 -1 30530
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform -1 0 6450 0 -1 30444
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform -1 0 6450 0 -1 30358
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform -1 0 6450 0 -1 30272
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform -1 0 6450 0 -1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform -1 0 6450 0 -1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform -1 0 6450 0 -1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform -1 0 6450 0 -1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform -1 0 6450 0 -1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform -1 0 6450 0 -1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform -1 0 6450 0 -1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform -1 0 6450 0 -1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform -1 0 6450 0 -1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform -1 0 6450 0 -1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform -1 0 6450 0 -1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform -1 0 6450 0 -1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform -1 0 6450 0 -1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform -1 0 6450 0 -1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform -1 0 6450 0 -1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform -1 0 6450 0 -1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform -1 0 6450 0 -1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform -1 0 6450 0 -1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform -1 0 6450 0 -1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform -1 0 6450 0 -1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform -1 0 6450 0 -1 28466
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 6450 0 -1 28380
box 0 0 6450 1720
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform -1 0 6450 0 -1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform -1 0 6450 0 -1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform -1 0 6450 0 -1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform -1 0 6450 0 -1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform -1 0 6450 0 -1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform -1 0 6450 0 -1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform -1 0 6450 0 -1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform -1 0 6450 0 -1 26058
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform -1 0 6450 0 -1 25972
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform -1 0 6450 0 -1 25886
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform -1 0 6450 0 -1 25800
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform -1 0 6450 0 -1 25714
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform -1 0 6450 0 -1 25628
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform -1 0 6450 0 -1 25542
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform -1 0 6450 0 -1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform -1 0 6450 0 -1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform -1 0 6450 0 -1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform -1 0 6450 0 -1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform -1 0 6450 0 -1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform -1 0 6450 0 -1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform -1 0 6450 0 -1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform -1 0 6450 0 -1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform -1 0 6450 0 -1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform -1 0 6450 0 -1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform -1 0 6450 0 -1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform -1 0 6450 0 -1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform -1 0 6450 0 -1 24424
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 6450 0 -1 24338
box 0 0 6450 1720
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform -1 0 6450 0 -1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform -1 0 6450 0 -1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform -1 0 6450 0 -1 22446
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform -1 0 6450 0 -1 22360
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform -1 0 6450 0 -1 22274
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform -1 0 6450 0 -1 22188
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform -1 0 6450 0 -1 22102
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform -1 0 6450 0 -1 22016
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform -1 0 6450 0 -1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform -1 0 6450 0 -1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform -1 0 6450 0 -1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform -1 0 6450 0 -1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform -1 0 6450 0 -1 21586
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform -1 0 6450 0 -1 21500
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform -1 0 6450 0 -1 21414
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform -1 0 6450 0 -1 21328
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform -1 0 6450 0 -1 21242
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform -1 0 6450 0 -1 21156
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform -1 0 6450 0 -1 21070
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform -1 0 6450 0 -1 20984
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform -1 0 6450 0 -1 20898
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform -1 0 6450 0 -1 20812
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform -1 0 6450 0 -1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform -1 0 6450 0 -1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform -1 0 6450 0 -1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform -1 0 6450 0 -1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform -1 0 6450 0 -1 20382
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 6450 0 -1 20296
box 0 0 6450 1720
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform -1 0 6450 0 -1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform -1 0 6450 0 -1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform -1 0 6450 0 -1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform -1 0 6450 0 -1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform -1 0 6450 0 -1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform -1 0 6450 0 -1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform -1 0 6450 0 -1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform -1 0 6450 0 -1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform -1 0 6450 0 -1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform -1 0 6450 0 -1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform -1 0 6450 0 -1 17716
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform -1 0 6450 0 -1 17630
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform -1 0 6450 0 -1 17544
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform -1 0 6450 0 -1 17458
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform -1 0 6450 0 -1 17372
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform -1 0 6450 0 -1 17286
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform -1 0 6450 0 -1 17200
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform -1 0 6450 0 -1 17114
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform -1 0 6450 0 -1 17028
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform -1 0 6450 0 -1 16942
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform -1 0 6450 0 -1 16856
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform -1 0 6450 0 -1 16770
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform -1 0 6450 0 -1 16684
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform -1 0 6450 0 -1 16598
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform -1 0 6450 0 -1 16512
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform -1 0 6450 0 -1 16426
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform -1 0 6450 0 -1 16340
box 0 0 6450 86
use datapath datapath_0
timestamp 1398693378
transform 1 0 7778 0 1 16334
box 0 0 25408 19490
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 36550 0 1 34744
box 0 0 6450 1720
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 36550 0 1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 36550 0 1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 36550 0 1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 36550 0 1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 36550 0 1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 36550 0 1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 36550 0 1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 36550 0 1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 36550 0 1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 36550 0 1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 36550 0 1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 36550 0 1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 36550 0 1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 36550 0 1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 36550 0 1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 36550 0 1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 36550 0 1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 36550 0 1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 36550 0 1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 36550 0 1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 36550 0 1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 36550 0 1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 36550 0 1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 36550 0 1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 36550 0 1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 36550 0 1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 36550 0 1 32422
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 36550 0 1 30702
box 0 0 6450 1720
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 36550 0 1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 36550 0 1 30530
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 36550 0 1 30444
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 36550 0 1 30358
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 36550 0 1 30272
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 36550 0 1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 36550 0 1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 36550 0 1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 36550 0 1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 36550 0 1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 36550 0 1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 36550 0 1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 36550 0 1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 36550 0 1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 36550 0 1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 36550 0 1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 36550 0 1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 36550 0 1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 36550 0 1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 36550 0 1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 36550 0 1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 36550 0 1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 36550 0 1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 36550 0 1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 36550 0 1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 36550 0 1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 36550 0 1 28380
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 36550 0 1 26660
box 0 0 6450 1720
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 36550 0 1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 36550 0 1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 36550 0 1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 36550 0 1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 36550 0 1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 36550 0 1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 36550 0 1 26058
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 36550 0 1 25972
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 36550 0 1 25886
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 36550 0 1 25800
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 36550 0 1 25714
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 36550 0 1 25628
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 36550 0 1 25542
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 36550 0 1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 36550 0 1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 36550 0 1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 36550 0 1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 36550 0 1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 36550 0 1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 36550 0 1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 36550 0 1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 36550 0 1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 36550 0 1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 36550 0 1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 36550 0 1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 36550 0 1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 36550 0 1 24338
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 36550 0 1 22618
box 0 0 6450 1720
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 36550 0 1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 36550 0 1 22446
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 36550 0 1 22360
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 36550 0 1 22274
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 36550 0 1 22188
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 36550 0 1 22102
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 36550 0 1 22016
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 36550 0 1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 36550 0 1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 36550 0 1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 36550 0 1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 36550 0 1 21586
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 36550 0 1 21500
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 36550 0 1 21414
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 36550 0 1 21328
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 36550 0 1 21242
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 36550 0 1 21156
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 36550 0 1 21070
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 36550 0 1 20984
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 36550 0 1 20898
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 36550 0 1 20812
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 36550 0 1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 36550 0 1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 36550 0 1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 36550 0 1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 36550 0 1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 36550 0 1 20296
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 36550 0 1 18576
box 0 0 6450 1720
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 36550 0 1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 36550 0 1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 36550 0 1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 36550 0 1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 36550 0 1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 36550 0 1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 36550 0 1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 36550 0 1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 36550 0 1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 36550 0 1 17716
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 36550 0 1 17630
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 36550 0 1 17544
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 36550 0 1 17458
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 36550 0 1 17372
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 36550 0 1 17286
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 36550 0 1 17200
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 36550 0 1 17114
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 36550 0 1 17028
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 36550 0 1 16942
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 36550 0 1 16856
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 36550 0 1 16770
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 36550 0 1 16684
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 36550 0 1 16598
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 1 0 36550 0 1 16512
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 1 0 36550 0 1 16426
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 1 0 36550 0 1 16340
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 6450 0 -1 16254
box 0 0 6450 1720
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 1 0 36550 0 1 16254
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform -1 0 6450 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform -1 0 6450 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform -1 0 6450 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform -1 0 6450 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform -1 0 6450 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform -1 0 6450 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform -1 0 6450 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform -1 0 6450 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform -1 0 6450 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform -1 0 6450 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform -1 0 6450 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform -1 0 6450 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform -1 0 6450 0 -1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform -1 0 6450 0 -1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform -1 0 6450 0 -1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform -1 0 6450 0 -1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform -1 0 6450 0 -1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform -1 0 6450 0 -1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform -1 0 6450 0 -1 12986
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform -1 0 6450 0 -1 12900
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform -1 0 6450 0 -1 12814
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform -1 0 6450 0 -1 12728
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform -1 0 6450 0 -1 12642
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform -1 0 6450 0 -1 12556
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform -1 0 6450 0 -1 12470
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform -1 0 6450 0 -1 12384
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform -1 0 6450 0 -1 12298
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 6450 0 -1 12212
box 0 0 6450 1720
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform -1 0 6450 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform -1 0 6450 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform -1 0 6450 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform -1 0 6450 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform -1 0 6450 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform -1 0 6450 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform -1 0 6450 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform -1 0 6450 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform -1 0 6450 0 -1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform -1 0 6450 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform -1 0 6450 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform -1 0 6450 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 6450 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 6450 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 6450 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 6450 0 -1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 6450 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 6450 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 6450 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 6450 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 6450 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 6450 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 6450 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 6450 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 6450 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 6450 0 -1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 6450 0 -1 8256
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 6450 0 -1 8170
box 0 0 6450 1720
use control control_0
timestamp 1398757585
transform 1 0 7900 0 1 6985
box 0 0 27529 8444
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 36550 0 1 14534
box 0 0 6450 1720
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 1 0 36550 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 1 0 36550 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 1 0 36550 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 1 0 36550 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 1 0 36550 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 1 0 36550 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 1 0 36550 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 1 0 36550 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 1 0 36550 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 1 0 36550 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 1 0 36550 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 1 0 36550 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 1 0 36550 0 1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 1 0 36550 0 1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 1 0 36550 0 1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 1 0 36550 0 1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 1 0 36550 0 1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 1 0 36550 0 1 12986
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 1 0 36550 0 1 12900
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 1 0 36550 0 1 12814
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 1 0 36550 0 1 12728
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 1 0 36550 0 1 12642
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 1 0 36550 0 1 12556
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 1 0 36550 0 1 12470
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 1 0 36550 0 1 12384
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 1 0 36550 0 1 12298
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 1 0 36550 0 1 12212
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 36550 0 1 10492
box 0 0 6450 1720
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 1 0 36550 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 1 0 36550 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 1 0 36550 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 1 0 36550 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 1 0 36550 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 1 0 36550 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 1 0 36550 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 1 0 36550 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 1 0 36550 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 1 0 36550 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 1 0 36550 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 1 0 36550 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 1 0 36550 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 1 0 36550 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 1 0 36550 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 1 0 36550 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 1 0 36550 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 1 0 36550 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 1 0 36550 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 1 0 36550 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 1 0 36550 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 1 0 36550 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 1 0 36550 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 1 0 36550 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 1 0 36550 0 1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 1 0 36550 0 1 8256
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 1 0 36550 0 1 8170
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 36550 0 1 6450
box 0 0 6450 1720
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 0 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 6450 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6536 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 8256 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 8342 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 8428 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 8514 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 8600 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8686 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8772 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8858 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8944 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 9030 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 9116 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 9202 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 9288 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 9374 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 9460 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 9546 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9632 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9718 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9804 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9890 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9976 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10062 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 11782 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 11868 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 11954 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 12040 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 12126 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 12212 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 12298 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 12384 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 12470 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 12556 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 12642 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 12728 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 12814 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12900 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12986 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 13072 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 13158 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 13244 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 13330 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 13416 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 13502 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 13588 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 15308 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 15394 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 15480 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 15566 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 15652 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 15738 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 15824 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 15910 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 15996 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 16082 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 16168 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 16254 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 16340 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 16426 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 16512 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 16598 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 16684 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 16770 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 16856 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 16942 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 17028 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 17114 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 18834 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 18920 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 19006 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 19092 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 19178 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 19264 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 19350 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 19436 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 19522 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 19608 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 19694 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 19780 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 19866 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 19952 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 20038 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 20124 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 20210 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 20296 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 20382 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 20468 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 20554 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 20640 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 22360 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 22446 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 22532 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 22618 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 22704 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 22790 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 22876 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 22962 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 23048 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 23134 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 23220 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 23306 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 23392 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 23478 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 23564 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 23650 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 23736 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 23822 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 23908 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 23994 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 24080 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 24166 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 25886 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 25972 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 26058 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 26144 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 26230 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 26316 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 26402 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 26488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 26574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 26660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 26746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 26832 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 26918 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 27004 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 27090 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 27176 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 27262 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 27348 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 27434 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 27520 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 27606 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 27692 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 29412 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 29498 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 29584 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 29670 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 29756 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 29842 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 29928 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 30014 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 30100 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 30186 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 30272 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 30358 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 30444 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 30530 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 30616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 30702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 30788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 30874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 30960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 31046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 31132 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 31218 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 32938 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 33024 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 33110 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 33196 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 33282 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 33368 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 33454 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 33540 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 33626 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 33712 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 33798 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 33884 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 33970 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 34056 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 34142 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 34228 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 34314 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 34400 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 34486 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 34572 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 34658 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 34744 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 36464 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 43000 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 6616 78 8176 1638 0 nIRQ
rlabel metal4 10142 78 11702 1638 0 Data[0]
rlabel metal4 13668 78 15228 1638 0 Data[1]
rlabel metal4 17194 78 18754 1638 0 Data[2]
rlabel metal4 20720 78 22280 1638 0 vdde!
rlabel metal4 24246 78 25806 1638 0 Data[3]
rlabel metal4 27772 78 29332 1638 0 Data[4]
rlabel metal4 31298 78 32858 1638 0 Data[5]
rlabel metal4 34824 78 36384 1638 0 gnde!
rlabel metal4 41362 6530 42922 8090 0 Data[6]
rlabel metal4 41362 10572 42922 12132 0 Data[7]
rlabel metal4 41362 14614 42922 16174 0 Data[8]
rlabel metal4 41362 18656 42922 20216 0 gnde!
rlabel metal4 41362 26740 42922 28300 0 Data[9]
rlabel metal4 41362 30782 42922 32342 0 Data[10]
rlabel metal4 41362 34824 42922 36384 0 Data[11]
rlabel metal4 34824 41276 36384 42836 0 vdde!
rlabel metal4 31298 41276 32858 42836 0 Data[12]
rlabel metal4 27772 41276 29332 42836 0 Data[13]
rlabel metal4 24246 41276 25806 42836 0 Data[14]
rlabel metal4 20720 41276 22280 42836 0 gnde!
rlabel metal4 17194 41276 18754 42836 0 Data[15]
rlabel metal4 13668 41276 15228 42836 0 ALE
rlabel metal4 10142 41276 11702 42836 0 nME
rlabel metal4 6616 41276 8176 42836 0 nWait
rlabel metal4 78 34824 1638 36384 0 nOE
rlabel metal4 78 30782 1638 32342 0 RnW
rlabel metal4 78 26740 1638 28300 0 SDO
rlabel metal4 78 22698 1638 24258 0 Vdd!
rlabel metal4 78 18656 1638 20216 0 SDI
rlabel metal4 78 14614 1638 16174 0 Test
rlabel metal4 78 10572 1638 12132 0 Clock
rlabel metal4 78 6530 1638 8090 0 nReset
<< end >>
