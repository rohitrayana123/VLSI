magic
tech c035u
timestamp 1394712986
<< metal1 >>
rect 2987 16649 3055 16659
rect 0 16517 35 16527
rect 2987 16517 3055 16527
rect 0 16494 35 16504
rect 2987 16494 3055 16504
rect 0 16456 35 16481
rect 2987 16456 3055 16481
rect 0 15811 35 15836
rect 2987 15811 3055 15836
rect 0 15788 35 15798
rect 2987 15788 3055 15798
rect 0 15765 35 15775
rect 2987 15765 3055 15775
rect 0 15742 35 15752
rect 2987 15742 3055 15752
rect 0 15713 35 15723
rect 2987 15713 3055 15723
rect 2987 15607 3055 15617
rect 0 15475 35 15485
rect 2987 15475 3055 15485
rect 0 15452 35 15462
rect 2987 15452 3055 15462
rect 0 15414 35 15439
rect 2987 15414 3055 15439
rect 0 14769 35 14794
rect 2987 14769 3055 14794
rect 0 14746 35 14756
rect 2987 14746 3055 14756
rect 0 14723 35 14733
rect 2987 14723 3055 14733
rect 0 14700 35 14710
rect 2987 14700 3055 14710
rect 0 14671 35 14681
rect 2987 14671 3055 14681
rect 2987 14565 3055 14575
rect 0 14433 35 14443
rect 2987 14433 3055 14443
rect 0 14410 35 14420
rect 2987 14410 3055 14420
rect 0 14372 35 14397
rect 2987 14372 3055 14397
rect 0 13727 35 13752
rect 2987 13727 3055 13752
rect 0 13704 35 13714
rect 2987 13704 3055 13714
rect 0 13681 35 13691
rect 2987 13681 3055 13691
rect 0 13658 35 13668
rect 2987 13658 3055 13668
rect 0 13629 35 13639
rect 2987 13629 3055 13639
rect 2987 13523 3055 13533
rect 0 13391 35 13401
rect 2987 13391 3055 13401
rect 0 13368 35 13378
rect 2987 13368 3055 13378
rect 0 13330 35 13355
rect 2987 13330 3055 13355
rect 0 12685 35 12710
rect 2987 12685 3055 12710
rect 0 12662 35 12672
rect 2987 12662 3055 12672
rect 0 12639 35 12649
rect 2987 12639 3055 12649
rect 0 12616 35 12626
rect 2987 12616 3055 12626
rect 0 12587 35 12597
rect 2987 12587 3055 12597
rect 2987 12481 3055 12491
rect 0 12349 35 12359
rect 2987 12349 3055 12359
rect 0 12326 35 12336
rect 2987 12326 3055 12336
rect 0 12288 35 12313
rect 2987 12288 3055 12313
rect 0 11643 35 11668
rect 2987 11643 3055 11668
rect 0 11620 35 11630
rect 2987 11620 3055 11630
rect 0 11597 35 11607
rect 2987 11597 3055 11607
rect 0 11574 35 11584
rect 2987 11574 3055 11584
rect 0 11545 35 11555
rect 2987 11545 3055 11555
rect 2987 11439 3055 11449
rect 0 11307 35 11317
rect 2987 11307 3055 11317
rect 0 11284 35 11294
rect 2987 11284 3055 11294
rect 0 11246 35 11271
rect 2987 11246 3055 11271
rect 0 10601 35 10626
rect 2987 10601 3055 10626
rect 0 10578 35 10588
rect 2987 10578 3055 10588
rect 0 10555 35 10565
rect 2987 10555 3055 10565
rect 0 10532 35 10542
rect 2987 10532 3055 10542
rect 0 10503 35 10513
rect 2987 10503 3055 10513
rect 2987 10397 3055 10407
rect 0 10265 35 10275
rect 2987 10265 3055 10275
rect 0 10242 35 10252
rect 2987 10242 3055 10252
rect 0 10204 35 10229
rect 2987 10204 3055 10229
rect 0 9559 35 9584
rect 2987 9559 3055 9584
rect 0 9536 35 9546
rect 2987 9536 3055 9546
rect 0 9513 35 9523
rect 2987 9513 3055 9523
rect 0 9490 35 9500
rect 2987 9490 3055 9500
rect 0 9461 35 9471
rect 2987 9461 3055 9471
rect 2987 9355 3055 9365
rect 0 9223 35 9233
rect 2987 9223 3055 9233
rect 0 9200 35 9210
rect 2987 9200 3055 9210
rect 0 9162 35 9187
rect 2987 9162 3055 9187
rect 0 8517 35 8542
rect 2987 8517 3055 8542
rect 0 8494 35 8504
rect 2987 8494 3055 8504
rect 0 8471 35 8481
rect 2987 8471 3055 8481
rect 0 8448 35 8458
rect 2987 8448 3055 8458
rect 0 8419 35 8429
rect 2987 8419 3055 8429
rect 2987 8313 3055 8323
rect 0 8181 35 8191
rect 2987 8181 3055 8191
rect 0 8158 35 8168
rect 2987 8158 3055 8168
rect 0 8120 35 8145
rect 2987 8120 3055 8145
rect 0 7475 35 7500
rect 2987 7475 3055 7500
rect 0 7452 35 7462
rect 2987 7452 3055 7462
rect 0 7429 35 7439
rect 2987 7429 3055 7439
rect 0 7406 35 7416
rect 2987 7406 3055 7416
rect 0 7377 35 7387
rect 2987 7377 3055 7387
rect 2987 7271 3055 7281
rect 0 7139 35 7149
rect 2987 7139 3055 7149
rect 0 7116 35 7126
rect 2987 7116 3055 7126
rect 0 7078 35 7103
rect 2987 7078 3055 7103
rect 0 6433 35 6458
rect 2987 6433 3055 6458
rect 0 6410 35 6420
rect 2987 6410 3055 6420
rect 0 6387 35 6397
rect 2987 6387 3055 6397
rect 0 6364 35 6374
rect 2987 6364 3055 6374
rect 0 6335 35 6345
rect 2987 6335 3055 6345
rect 2987 6229 3055 6239
rect 0 6097 35 6107
rect 2987 6097 3055 6107
rect 0 6074 35 6084
rect 2987 6074 3055 6084
rect 0 6036 35 6061
rect 2987 6036 3055 6061
rect 0 5391 35 5416
rect 2987 5391 3055 5416
rect 0 5368 35 5378
rect 2987 5368 3055 5378
rect 0 5345 35 5355
rect 2987 5345 3055 5355
rect 0 5322 35 5332
rect 2987 5322 3055 5332
rect 0 5293 35 5303
rect 2987 5293 3055 5303
rect 2987 5187 3055 5197
rect 0 5055 35 5065
rect 2987 5055 3055 5065
rect 0 5032 35 5042
rect 2987 5032 3055 5042
rect 0 4994 35 5019
rect 2987 4994 3055 5019
rect 0 4349 35 4374
rect 2987 4349 3055 4374
rect 0 4326 35 4336
rect 2987 4326 3055 4336
rect 0 4303 35 4313
rect 2987 4303 3055 4313
rect 0 4280 35 4290
rect 2987 4280 3055 4290
rect 0 4251 35 4261
rect 2987 4251 3055 4261
rect 2987 4145 3055 4155
rect 0 4013 35 4023
rect 2987 4013 3055 4023
rect 0 3990 35 4000
rect 2987 3990 3055 4000
rect 0 3952 35 3977
rect 2987 3952 3055 3977
rect 0 3307 35 3332
rect 2987 3307 3055 3332
rect 0 3284 35 3294
rect 2987 3284 3055 3294
rect 0 3261 35 3271
rect 2987 3261 3055 3271
rect 0 3238 35 3248
rect 2987 3238 3055 3248
rect 0 3209 35 3219
rect 2987 3209 3055 3219
rect 2987 3103 3055 3113
rect 0 2971 35 2981
rect 2987 2971 3055 2981
rect 0 2948 35 2958
rect 2987 2948 3055 2958
rect 0 2910 35 2935
rect 2987 2910 3055 2935
rect 0 2265 35 2290
rect 2987 2265 3055 2290
rect 0 2242 35 2252
rect 2987 2242 3055 2252
rect 0 2219 35 2229
rect 2987 2219 3055 2229
rect 0 2196 35 2206
rect 2987 2196 3055 2206
rect 0 2167 35 2177
rect 2987 2167 3055 2177
rect 2987 2061 3055 2071
rect 0 1929 35 1939
rect 2987 1929 3055 1939
rect 0 1906 35 1916
rect 2987 1906 3055 1916
rect 0 1868 35 1893
rect 2987 1868 3055 1893
rect 0 1223 35 1248
rect 2987 1223 3055 1248
rect 0 1200 35 1210
rect 2987 1200 3055 1210
rect 0 1177 35 1187
rect 2987 1177 3055 1187
rect 0 1154 35 1164
rect 2987 1154 3055 1164
rect 0 1125 35 1135
rect 2987 1125 3055 1135
rect 2987 1019 3055 1029
rect 0 887 35 897
rect 2987 887 3055 897
rect 0 864 35 874
rect 2987 864 3055 874
rect 0 826 35 851
rect 2987 826 3055 851
rect 0 181 35 206
rect 2987 181 3055 206
rect 0 158 35 168
rect 2987 158 3055 168
rect 0 135 35 145
rect 2987 135 3055 145
rect 0 112 35 122
rect 2987 112 3055 122
rect 0 83 35 93
rect 2987 83 3055 93
<< metal2 >>
rect 251 16711 263 16888
rect 395 16711 407 16888
rect 611 16711 623 16888
rect 1355 16711 1367 16888
rect 1523 16711 1535 16888
rect 1907 16711 1919 16888
rect 2123 16711 2135 16888
rect 2867 16711 2879 16888
rect 251 0 263 39
rect 395 0 407 39
rect 611 0 623 39
rect 1355 0 1367 39
rect 1523 0 1535 39
rect 1907 0 1919 39
rect 2123 0 2135 39
rect 2603 0 2615 39
rect 2867 0 2879 39
use Pc_slice Pc_slice_0
array 0 0 2952 0 15 1042
timestamp 1394709084
transform 1 0 35 0 1 39
box 0 0 2952 1042
<< labels >>
rlabel metal1 0 112 0 122 3 nReset
rlabel metal1 0 135 0 145 3 Test
rlabel metal1 0 158 0 168 3 Clock
rlabel metal1 0 181 0 206 3 GND!
rlabel metal1 0 1906 0 1916 3 Scan
rlabel metal1 0 1929 0 1939 3 ScanReturn
rlabel metal1 0 1868 0 1893 3 Vdd!
rlabel metal1 0 1223 0 1248 3 GND!
rlabel metal1 0 1154 0 1164 3 nReset
rlabel metal1 0 1177 0 1187 3 Test
rlabel metal1 0 1200 0 1210 3 Clock
rlabel metal1 0 887 0 897 3 ScanReturn
rlabel metal1 0 864 0 874 3 Scan
rlabel metal1 0 826 0 851 3 Vdd!
rlabel metal1 0 2196 0 2206 3 nReset
rlabel metal1 0 2219 0 2229 3 Test
rlabel metal1 0 2242 0 2252 3 Clock
rlabel metal1 0 2265 0 2290 3 GND!
rlabel metal1 0 2971 0 2981 3 ScanReturn
rlabel metal1 0 2948 0 2958 3 Scan
rlabel metal1 0 2910 0 2935 3 Vdd!
rlabel metal1 0 3307 0 3332 3 GND!
rlabel metal1 0 3261 0 3271 3 Test
rlabel metal1 0 3284 0 3294 3 Clock
rlabel metal1 0 3238 0 3248 3 nReset
rlabel metal1 0 4013 0 4023 3 ScanReturn
rlabel metal1 0 3990 0 4000 3 Scan
rlabel metal1 0 3952 0 3977 3 Vdd!
rlabel metal1 0 6097 0 6107 3 ScanReturn
rlabel metal1 0 6074 0 6084 3 Scan
rlabel metal1 0 6036 0 6061 3 Vdd!
rlabel metal1 0 6433 0 6458 3 GND!
rlabel metal1 0 6387 0 6397 3 Test
rlabel metal1 0 6410 0 6420 3 Clock
rlabel metal1 0 6364 0 6374 3 nReset
rlabel metal1 0 7139 0 7149 3 ScanReturn
rlabel metal1 0 7116 0 7126 3 Scan
rlabel metal1 0 7078 0 7103 3 Vdd!
rlabel metal1 0 7475 0 7500 3 GND!
rlabel metal1 0 7429 0 7439 3 Test
rlabel metal1 0 7452 0 7462 3 Clock
rlabel metal1 0 7406 0 7416 3 nReset
rlabel metal1 0 9162 0 9187 3 Vdd!
rlabel metal1 0 9200 0 9210 3 Scan
rlabel metal1 0 9223 0 9233 3 ScanReturn
rlabel metal1 0 9559 0 9584 3 GND!
rlabel metal1 0 9490 0 9500 3 nReset
rlabel metal1 0 9513 0 9523 3 Test
rlabel metal1 0 9536 0 9546 3 Clock
rlabel metal1 0 10265 0 10275 3 ScanReturn
rlabel metal1 0 10242 0 10252 3 Scan
rlabel metal1 0 10204 0 10229 3 Vdd!
rlabel metal1 0 10601 0 10626 3 GND!
rlabel metal1 0 10578 0 10588 3 Clock
rlabel metal1 0 10555 0 10565 3 Test
rlabel metal1 0 10532 0 10542 3 nReset
rlabel metal1 0 11307 0 11317 3 ScanReturn
rlabel metal1 0 11284 0 11294 3 Scan
rlabel metal1 0 11246 0 11271 3 Vdd!
rlabel metal1 0 11643 0 11668 3 GND!
rlabel metal1 0 11597 0 11607 3 Test
rlabel metal1 0 11620 0 11630 3 Clock
rlabel metal1 0 11574 0 11584 3 nReset
rlabel metal1 0 12288 0 12313 3 Vdd!
rlabel metal1 0 15811 0 15836 3 GND!
rlabel metal1 0 15742 0 15752 3 nReset
rlabel metal1 0 15765 0 15775 3 Test
rlabel metal1 0 15788 0 15798 3 Clock
rlabel metal1 0 8517 0 8542 3 GND!
rlabel metal1 0 8471 0 8481 3 Test
rlabel metal1 0 8494 0 8504 3 Clock
rlabel metal1 0 8448 0 8458 3 nReset
rlabel metal1 0 4349 0 4374 3 GND!
rlabel metal1 0 4303 0 4313 3 Test
rlabel metal1 0 4326 0 4336 3 Clock
rlabel metal1 0 4280 0 4290 3 nReset
rlabel metal1 0 4994 0 5019 3 Vdd!
rlabel metal1 0 5032 0 5042 3 Scan
rlabel metal1 0 5055 0 5065 3 ScanReturn
rlabel metal1 0 5391 0 5416 3 GND!
rlabel metal1 0 5345 0 5355 3 Test
rlabel metal1 0 5368 0 5378 3 Clock
rlabel metal1 0 5322 0 5332 3 nReset
rlabel metal1 0 12685 0 12710 3 GND!
rlabel metal1 0 12639 0 12649 3 Test
rlabel metal1 0 12662 0 12672 3 Clock
rlabel metal1 0 12616 0 12626 3 nReset
rlabel metal1 0 12326 0 12336 3 Scan
rlabel metal1 0 12349 0 12359 3 ScanReturn
rlabel metal1 0 14372 0 14397 3 Vdd!
rlabel metal1 0 14410 0 14420 3 Scan
rlabel metal1 0 14433 0 14443 3 ScanReturn
rlabel metal1 0 14700 0 14710 3 nReset
rlabel metal1 0 14723 0 14733 3 Test
rlabel metal1 0 14746 0 14756 3 Clock
rlabel metal1 0 14769 0 14794 3 GND!
rlabel metal1 0 13658 0 13668 3 nReset
rlabel metal1 0 13681 0 13691 3 Test
rlabel metal1 0 13704 0 13714 3 Clock
rlabel metal1 0 13727 0 13752 3 GND!
rlabel metal1 0 16517 0 16527 3 ScanReturn
rlabel metal1 0 16494 0 16504 3 Scan
rlabel metal1 0 16456 0 16481 3 Vdd!
rlabel metal1 0 13330 0 13355 3 Vdd!
rlabel metal1 0 13368 0 13378 3 Scan
rlabel metal1 0 13391 0 13401 3 ScanReturn
rlabel metal1 0 8181 0 8191 3 ScanReturn
rlabel metal1 0 8158 0 8168 3 Scan
rlabel metal1 0 8120 0 8145 3 Vdd!
rlabel metal1 0 15414 0 15439 3 Vdd!
rlabel metal1 0 15452 0 15462 3 Scan
rlabel metal1 0 15475 0 15485 3 ScanReturn
rlabel metal1 0 83 0 93 3 SysBus[0]
rlabel metal1 0 1125 0 1135 3 SysBus[1]
rlabel metal1 0 2167 0 2177 3 SysBus[2]
rlabel metal1 0 3209 0 3219 3 SysBus[3]
rlabel metal1 0 4251 0 4261 3 SysBus[4]
rlabel metal1 0 5293 0 5303 3 SysBus[5]
rlabel metal1 0 6335 0 6345 3 SysBus[6]
rlabel metal1 0 7377 0 7387 3 SysBus[7]
rlabel metal1 0 8419 0 8429 3 SysBus[8]
rlabel metal1 0 9461 0 9471 3 SysBus[9]
rlabel metal1 0 10503 0 10513 3 SysBus[10]
rlabel metal1 0 11545 0 11555 3 SysBus[11]
rlabel metal1 0 12587 0 12597 3 SysBus[12]
rlabel metal1 0 13629 0 13639 3 SysBus[13]
rlabel metal1 0 14671 0 14681 3 SysBus[14]
rlabel metal1 0 15713 0 15723 3 SysBus[15]
rlabel metal1 3055 12481 3055 12491 7 ALU[11]
rlabel metal1 3055 12685 3055 12710 7 GND!
rlabel metal1 3055 12662 3055 12672 7 Clock
rlabel metal1 3055 12639 3055 12649 7 Test
rlabel metal1 3055 12616 3055 12626 7 nReset
rlabel metal1 3055 12587 3055 12597 7 SysBus[12]
rlabel metal1 3055 12349 3055 12359 7 ScanReturn
rlabel metal1 3055 12326 3055 12336 7 Scan
rlabel metal1 3055 12288 3055 12313 7 Vdd!
rlabel metal1 3055 13727 3055 13752 7 GND!
rlabel metal1 3055 13704 3055 13714 7 Clock
rlabel metal1 3055 13681 3055 13691 7 Test
rlabel metal1 3055 13658 3055 13668 7 nReset
rlabel metal1 3055 13391 3055 13401 7 ScanReturn
rlabel metal1 3055 13368 3055 13378 7 Scan
rlabel metal1 3055 13330 3055 13355 7 Vdd!
rlabel metal1 3055 13523 3055 13533 7 ALU[12]
rlabel metal1 3055 13629 3055 13639 7 SysBus[13]
rlabel metal1 3055 14700 3055 14710 7 nReset
rlabel metal1 3055 14723 3055 14733 7 Test
rlabel metal1 3055 14746 3055 14756 7 Clock
rlabel metal1 3055 14769 3055 14794 7 GND!
rlabel metal1 3055 14372 3055 14397 7 Vdd!
rlabel metal1 3055 14410 3055 14420 7 Scan
rlabel metal1 3055 14433 3055 14443 7 ScanReturn
rlabel metal1 3055 15414 3055 15439 7 Vdd!
rlabel metal1 3055 15452 3055 15462 7 Scan
rlabel metal1 3055 15475 3055 15485 7 ScanReturn
rlabel metal1 3055 15742 3055 15752 7 nReset
rlabel metal1 3055 15765 3055 15775 7 Test
rlabel metal1 3055 15788 3055 15798 7 Clock
rlabel metal1 3055 15811 3055 15836 7 GND!
rlabel metal1 3055 15607 3055 15617 7 ALU[14]
rlabel metal1 3055 15713 3055 15723 7 SysBus[15]
rlabel metal1 3055 16456 3055 16481 7 Vdd!
rlabel metal1 3055 16494 3055 16504 7 Scan
rlabel metal1 3055 16517 3055 16527 7 ScanReturn
rlabel metal1 3055 16649 3055 16659 7 ALU[15]
rlabel metal1 3055 112 3055 122 7 nReset
rlabel metal1 3055 135 3055 145 7 Test
rlabel metal1 3055 158 3055 168 7 Clock
rlabel metal1 3055 181 3055 206 7 GND!
rlabel metal1 3055 83 3055 93 7 SysBus[0]
rlabel metal1 3055 1154 3055 1164 7 nReset
rlabel metal1 3055 1177 3055 1187 7 Test
rlabel metal1 3055 1200 3055 1210 7 Clock
rlabel metal1 3055 1223 3055 1248 7 GND!
rlabel metal1 3055 826 3055 851 7 Vdd!
rlabel metal1 3055 864 3055 874 7 Scan
rlabel metal1 3055 887 3055 897 7 ScanReturn
rlabel metal1 3055 1125 3055 1135 7 SysBus[1]
rlabel metal1 3055 1019 3055 1029 7 ALU[0]
rlabel metal1 3055 1929 3055 1939 7 ScanReturn
rlabel metal1 3055 1906 3055 1916 7 Scan
rlabel metal1 3055 1868 3055 1893 7 Vdd!
rlabel metal1 3055 2265 3055 2290 7 GND!
rlabel metal1 3055 2242 3055 2252 7 Clock
rlabel metal1 3055 2219 3055 2229 7 Test
rlabel metal1 3055 2196 3055 2206 7 nReset
rlabel metal1 3055 2061 3055 2071 7 ALU[1]
rlabel metal1 3055 2167 3055 2177 7 SysBus[2]
rlabel metal1 3055 3307 3055 3332 7 GND!
rlabel metal1 3055 3284 3055 3294 7 Clock
rlabel metal1 3055 3261 3055 3271 7 Test
rlabel metal1 3055 3238 3055 3248 7 nReset
rlabel metal1 3055 2971 3055 2981 7 ScanReturn
rlabel metal1 3055 2948 3055 2958 7 Scan
rlabel metal1 3055 2910 3055 2935 7 Vdd!
rlabel metal1 3055 3103 3055 3113 7 ALU[2]
rlabel metal1 3055 3209 3055 3219 7 SysBus[3]
rlabel metal1 3055 4349 3055 4374 7 GND!
rlabel metal1 3055 4326 3055 4336 7 Clock
rlabel metal1 3055 4303 3055 4313 7 Test
rlabel metal1 3055 4280 3055 4290 7 nReset
rlabel metal1 3055 4013 3055 4023 7 ScanReturn
rlabel metal1 3055 3990 3055 4000 7 Scan
rlabel metal1 3055 3952 3055 3977 7 Vdd!
rlabel metal1 3055 4145 3055 4155 7 ALU[3]
rlabel metal1 3055 4251 3055 4261 7 SysBus[4]
rlabel metal1 3055 5055 3055 5065 7 ScanReturn
rlabel metal1 3055 5032 3055 5042 7 Scan
rlabel metal1 3055 4994 3055 5019 7 Vdd!
rlabel metal1 3055 5391 3055 5416 7 GND!
rlabel metal1 3055 5368 3055 5378 7 Clock
rlabel metal1 3055 5345 3055 5355 7 Test
rlabel metal1 3055 5322 3055 5332 7 nReset
rlabel metal1 3055 5187 3055 5197 7 ALU[4]
rlabel metal1 3055 5293 3055 5303 7 SysBus[5]
rlabel metal1 3055 6097 3055 6107 7 ScanReturn
rlabel metal1 3055 6074 3055 6084 7 Scan
rlabel metal1 3055 6036 3055 6061 7 Vdd!
rlabel metal1 3055 6433 3055 6458 7 GND!
rlabel metal1 3055 6410 3055 6420 7 Clock
rlabel metal1 3055 6387 3055 6397 7 Test
rlabel metal1 3055 6364 3055 6374 7 nReset
rlabel metal1 3055 6229 3055 6239 7 ALU[5]
rlabel metal1 3055 6335 3055 6345 7 SysBus[6]
rlabel metal1 3055 7475 3055 7500 7 GND!
rlabel metal1 3055 7452 3055 7462 7 Clock
rlabel metal1 3055 7429 3055 7439 7 Test
rlabel metal1 3055 7406 3055 7416 7 nReset
rlabel metal1 3055 7139 3055 7149 7 ScanReturn
rlabel metal1 3055 7116 3055 7126 7 Scan
rlabel metal1 3055 7078 3055 7103 7 Vdd!
rlabel metal1 3055 7271 3055 7281 7 ALU[6]
rlabel metal1 3055 7377 3055 7387 7 SysBus[7]
rlabel metal1 3055 8158 3055 8168 7 Scan
rlabel metal1 3055 8120 3055 8145 7 Vdd!
rlabel metal1 3055 8181 3055 8191 7 ScanReturn
rlabel metal1 3055 8517 3055 8542 7 GND!
rlabel metal1 3055 8494 3055 8504 7 Clock
rlabel metal1 3055 8471 3055 8481 7 Test
rlabel metal1 3055 8448 3055 8458 7 nReset
rlabel metal1 3055 8313 3055 8323 7 ALU[7]
rlabel metal1 3055 8419 3055 8429 7 SysBus[8]
rlabel metal1 3055 9223 3055 9233 7 ScanReturn
rlabel metal1 3055 9200 3055 9210 7 Scan
rlabel metal1 3055 9162 3055 9187 7 Vdd!
rlabel metal1 3055 9355 3055 9365 7 ALU[8]
rlabel metal1 3055 9559 3055 9584 7 GND!
rlabel metal1 3055 9536 3055 9546 7 Clock
rlabel metal1 3055 9513 3055 9523 7 Test
rlabel metal1 3055 9490 3055 9500 7 nReset
rlabel metal1 3055 9461 3055 9471 7 SysBus[9]
rlabel metal1 3055 10204 3055 10229 7 Vdd!
rlabel metal1 3055 10242 3055 10252 7 Scan
rlabel metal1 3055 10265 3055 10275 7 ScanReturn
rlabel metal1 3055 10601 3055 10626 7 GND!
rlabel metal1 3055 10578 3055 10588 7 Clock
rlabel metal1 3055 10555 3055 10565 7 Test
rlabel metal1 3055 10532 3055 10542 7 nReset
rlabel metal1 3055 10397 3055 10407 7 ALU[9]
rlabel metal1 3055 10503 3055 10513 7 SysBus[10]
rlabel metal1 3055 11643 3055 11668 7 GND!
rlabel metal1 3055 11620 3055 11630 7 Clock
rlabel metal1 3055 11597 3055 11607 7 Test
rlabel metal1 3055 11574 3055 11584 7 nReset
rlabel metal1 3055 11307 3055 11317 7 ScanReturn
rlabel metal1 3055 11284 3055 11294 7 Scan
rlabel metal1 3055 11246 3055 11271 7 Vdd!
rlabel metal1 3055 11545 3055 11555 7 SysBus[11]
rlabel metal1 3055 11439 3055 11449 7 ALU[10]
rlabel metal1 3055 14671 3055 14681 7 SysBus[14]
rlabel metal1 3055 14565 3055 14575 7 ALU[13]
rlabel metal2 395 16888 407 16888 5 LrSel
rlabel metal2 611 16888 623 16888 5 LrWe
rlabel metal2 1355 16888 1367 16888 5 LrEn
rlabel metal2 1523 16888 1535 16888 5 PcSel[0]
rlabel metal2 1907 16888 1919 16888 5 PcSel[1]
rlabel metal2 2123 16888 2135 16888 5 PcWe
rlabel metal2 2867 16888 2879 16888 5 PcEn
rlabel metal2 251 16888 263 16888 5 PcIncCout
rlabel metal2 251 0 263 0 1 PcIncCin
rlabel metal2 395 0 407 0 1 LrSel
rlabel metal2 611 0 623 0 1 LrWe
rlabel metal2 1355 0 1367 0 1 LrEn
rlabel metal2 1523 0 1535 0 1 PcSel[0]
rlabel metal2 1907 0 1919 0 1 PcSel[1]
rlabel metal2 2123 0 2135 0 1 PcWe
rlabel metal2 2867 0 2879 0 1 PcEn
rlabel metal2 2603 0 2615 0 1 Pc
<< end >>
