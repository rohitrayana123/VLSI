magic
tech c035u
timestamp 1394308690
<< metal1 >>
rect 0 155 1469 165
rect 0 95 1469 105
<< metal2 >>
rect 5 970 205 1079
rect 221 970 233 1079
rect 245 970 257 1079
rect 269 970 281 1079
rect 293 970 305 1079
rect 5 0 205 171
rect 221 0 233 171
rect 245 0 257 171
rect 269 0 281 171
rect 293 0 305 171
use leftbuf  leftbuf_0
timestamp 1386242881
transform 1 0 5 0 1 171
box 0 0 1464 799
<< labels >>
rlabel metal2 5 0 205 0 1 Vdd!
rlabel metal2 221 0 233 0 1 SDI
rlabel metal2 245 0 257 0 1 Test
rlabel metal2 269 0 281 0 1 Clock
rlabel metal2 293 0 305 0 1 nReset
rlabel metal2 5 1079 205 1079 5 Vdd!
rlabel metal2 221 1079 233 1079 5 SDO
rlabel metal2 245 1079 257 1079 5 Test
rlabel metal2 269 1079 281 1079 5 Clock
rlabel metal2 293 1079 305 1079 5 nReset
rlabel metal1 0 95 0 105 3 SysBus
rlabel metal1 0 155 0 165 3 Ir
rlabel metal1 1469 95 1469 105 7 SysBus
rlabel metal1 1469 155 1469 165 7 Ir
<< end >>
