magic
tech c035u
timestamp 1394530846
<< metal1 >>
rect -832 17850 0 17860
rect -832 17784 0 17794
rect -832 16674 0 16684
rect -832 16608 0 16618
rect -832 15498 0 15508
rect -832 15432 0 15442
rect -832 14322 0 14332
rect -832 14256 0 14266
rect -832 13146 0 13156
rect -832 13080 0 13090
rect -832 11970 0 11980
rect -832 11904 0 11914
rect -832 10794 0 10804
rect -832 10728 0 10738
rect -832 9618 0 9628
rect -832 9552 0 9562
rect -832 8442 0 8452
rect -832 8376 0 8386
rect -832 7266 0 7276
rect -832 7200 0 7210
rect -832 6090 0 6100
rect -832 6024 0 6034
rect -832 4914 0 4924
rect -832 4848 0 4858
rect -832 3738 0 3748
rect -832 3672 0 3682
rect -832 2562 0 2572
rect -832 2496 0 2506
rect -832 1386 0 1396
rect -832 1320 0 1330
rect -832 210 0 220
rect -832 144 0 154
use slice17  slice17_0
timestamp 1394529261
transform 1 0 4334 0 1 18865
box -4329 0 18911 1795
use leftbuf_slice  leftbuf_slice_0
array 0 0 1469 0 15 1176
timestamp 1394489502
transform 1 0 0 0 1 55
box 0 -6 1469 1170
use IrAA  IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 1469 0 1 9568
box 0 -111 1008 1065
use LLIcell_U  LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1393855556
transform 1 0 22517 0 1 9568
box 0 0 192 1042
use IrBA  IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 1469 0 1 6040
box 0 -111 1008 1065
use IrBB  IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 1469 0 1 161
box 0 -112 1008 1064
use LLIcell_L  LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 22517 0 1 160
box 0 0 192 1042
use Datapath_slice  Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394491434
transform 1 0 2477 0 1 49
box 0 0 20768 1176
<< labels >>
rlabel metal1 -832 144 -832 154 3 SysBus[0]
rlabel metal1 -832 1320 -832 1330 3 SysBus[1]
rlabel metal1 -832 2496 -832 2506 3 SysBus[2]
rlabel metal1 -832 3672 -832 3682 3 SysBus[3]
rlabel metal1 -832 4848 -832 4858 3 SysBus[4]
rlabel metal1 -832 6024 -832 6034 3 SysBus[5]
rlabel metal1 -832 7200 -832 7210 3 SysBus[6]
rlabel metal1 -832 8376 -832 8386 3 SysBus[7]
rlabel metal1 -832 9552 -832 9562 3 SysBus[8]
rlabel metal1 -832 10728 -832 10738 3 SysBus[9]
rlabel metal1 -832 11904 -832 11914 3 SysBus[10]
rlabel metal1 -832 13080 -832 13090 3 SysBus[11]
rlabel metal1 -832 14256 -832 14266 3 SysBus[12]
rlabel metal1 -832 15432 -832 15442 3 SysBus[13]
rlabel metal1 -832 16608 -832 16618 3 SysBus[14]
rlabel metal1 -832 17784 -832 17794 3 SysBus[15]
rlabel metal1 -832 210 -832 220 3 Ir[0]
rlabel metal1 -832 1386 -832 1396 3 Ir[1]
rlabel metal1 -832 2562 -832 2572 3 Ir[2]
rlabel metal1 -832 3738 -832 3748 3 Ir[3]
rlabel metal1 -832 4914 -832 4924 3 Ir[4]
rlabel metal1 -832 6090 -832 6100 3 Ir[5]
rlabel metal1 -832 7266 -832 7276 3 Ir[6]
rlabel metal1 -832 8442 -832 8452 3 Ir[7]
rlabel metal1 -832 9618 -832 9628 3 Ir[8]
rlabel metal1 -832 10794 -832 10804 3 Ir[9]
rlabel metal1 -832 11970 -832 11980 3 Ir[10]
rlabel metal1 -832 13146 -832 13156 3 Ir[11]
rlabel metal1 -832 14322 -832 14332 3 Ir[12]
rlabel metal1 -832 15498 -832 15508 3 Ir[13]
rlabel metal1 -832 16674 -832 16684 3 Ir[14]
rlabel metal1 -832 17850 -832 17860 3 Ir[15]
<< end >>
