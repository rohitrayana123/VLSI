../../../Design/Implementation/verification/prog_stim.sv