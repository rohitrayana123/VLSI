magic
tech c035u
timestamp 1393699629
<< error_ps >>
rect 2303 1021 2317 1022
<< glass >>
rect -30 1201 599 1587
rect 6240 1318 7034 1423
rect 1512 1221 1656 1308
rect 3863 1019 4105 1160
rect 4607 1039 5688 1127
<< metal1 >>
rect 2677 1067 3719 1077
rect 2557 1045 3623 1055
rect 2317 1023 3431 1033
rect 2077 1002 3239 1012
rect 1957 980 3143 990
rect 709 958 1103 968
rect 2797 958 3047 968
rect 3061 958 3815 968
rect 829 936 1079 946
rect 1165 936 1320 946
rect 1381 936 1439 946
rect 2437 936 2951 946
rect 2965 936 3527 946
rect 925 914 960 924
rect 1045 914 1199 924
rect 1285 914 1415 924
rect 2197 914 2855 924
rect 2869 914 3335 924
rect 3565 914 5615 924
rect 517 892 671 902
rect 685 892 863 902
rect 877 892 2039 902
rect 2053 892 2279 902
rect 2293 892 2519 902
rect 2533 892 2759 902
rect 2773 892 3935 902
rect 3949 892 4271 902
rect 397 870 1343 880
rect 1357 870 2135 880
rect 2149 870 2255 880
rect 2269 870 2615 880
rect 2629 870 2735 880
rect 2749 870 3911 880
rect 3925 870 4151 880
rect 4165 870 4247 880
rect 4261 870 4775 880
rect 4789 870 5759 880
rect 277 848 647 858
rect 661 848 983 858
rect 997 848 1559 858
rect 1573 848 2351 858
rect 2365 848 2471 858
rect 2485 848 2591 858
rect 2605 848 2711 858
rect 2725 848 5735 858
rect 5965 848 6023 858
rect 157 826 791 836
rect 805 826 1223 836
rect 1237 826 1799 836
rect 1813 826 3887 836
rect 3973 826 4006 836
rect 4333 826 4391 836
rect 4717 826 4895 836
rect 4957 826 4991 836
rect 5101 826 5135 836
rect 5149 826 5255 836
rect 5269 826 5375 836
rect 5389 826 5495 836
rect 5557 826 5591 836
rect 5821 826 5999 836
rect 6277 826 6575 836
rect 37 804 1535 814
rect 1549 804 1679 814
rect 1693 804 1775 814
rect 1789 804 4031 814
rect 4213 804 4367 814
rect 4453 804 4487 814
rect 4837 804 4871 814
rect 4885 804 6047 814
rect 6109 804 6143 814
rect 6349 804 6383 814
rect 6613 804 6887 814
rect 85 -15 6180 -5
rect 6409 -13 6778 -3
rect 205 -37 5868 -27
rect 325 -59 5892 -49
rect 445 -81 2508 -71
rect 3120 -83 3804 -73
rect 565 -103 5916 -93
rect 1824 -123 3036 -113
rect 3072 -123 4215 -113
rect 1728 -143 3132 -133
rect 3308 -143 3468 -133
rect 3552 -143 4159 -133
rect 1563 -163 2892 -153
rect 3648 -163 6362 -153
rect 2976 -183 4669 -173
rect 1488 -203 6420 -193
rect 1632 -223 6300 -213
<< m2contact >>
rect 2663 1065 2677 1079
rect 3719 1065 3733 1079
rect 2543 1043 2557 1057
rect 3623 1043 3637 1057
rect 2303 1021 2317 1035
rect 3431 1021 3445 1035
rect 2063 1000 2077 1014
rect 3239 999 3253 1013
rect 1943 978 1957 992
rect 3143 978 3157 992
rect 695 956 709 970
rect 1103 956 1117 970
rect 2783 956 2797 970
rect 3047 956 3061 970
rect 3815 956 3829 970
rect 815 934 829 948
rect 1079 934 1093 948
rect 1151 934 1165 948
rect 1320 934 1334 948
rect 1367 934 1381 948
rect 1439 934 1453 948
rect 2423 934 2437 948
rect 2951 934 2965 948
rect 3527 934 3541 948
rect 911 912 925 926
rect 960 912 974 926
rect 1031 912 1045 926
rect 1199 912 1213 926
rect 1271 912 1285 926
rect 1415 912 1429 926
rect 2183 912 2197 926
rect 2855 912 2869 926
rect 3335 912 3349 926
rect 3551 912 3565 926
rect 5615 912 5629 926
rect 503 890 517 904
rect 671 890 685 904
rect 863 890 877 904
rect 2039 890 2053 904
rect 2279 890 2293 904
rect 2519 890 2533 904
rect 2759 890 2773 904
rect 3935 890 3949 904
rect 4271 890 4285 904
rect 383 868 397 882
rect 1343 868 1357 882
rect 2135 868 2149 882
rect 2255 868 2269 882
rect 2615 868 2629 882
rect 2735 868 2749 882
rect 3911 868 3925 882
rect 4151 868 4165 882
rect 4247 868 4261 882
rect 4775 868 4789 882
rect 5759 868 5773 882
rect 263 846 277 860
rect 647 846 661 860
rect 983 846 997 860
rect 1559 846 1573 860
rect 2351 846 2365 860
rect 2471 846 2485 860
rect 2591 846 2605 860
rect 2711 846 2725 860
rect 5735 846 5749 860
rect 5951 846 5965 860
rect 6023 846 6037 860
rect 143 824 157 838
rect 791 824 805 838
rect 1223 824 1237 838
rect 1799 824 1813 838
rect 3887 824 3901 838
rect 3959 824 3973 838
rect 4006 824 4020 838
rect 4319 824 4333 838
rect 4391 824 4405 838
rect 4703 824 4717 838
rect 4895 824 4909 838
rect 4943 824 4957 838
rect 4991 824 5005 838
rect 5087 824 5101 838
rect 5135 824 5149 838
rect 5255 824 5269 838
rect 5375 824 5389 838
rect 5495 824 5509 838
rect 5543 824 5557 838
rect 5591 824 5605 838
rect 5807 824 5821 838
rect 5999 824 6013 838
rect 6263 824 6277 838
rect 6575 824 6589 838
rect 23 802 37 816
rect 1535 802 1549 816
rect 1679 802 1693 816
rect 1775 802 1789 816
rect 4031 802 4045 816
rect 4199 802 4213 816
rect 4367 802 4381 816
rect 4439 802 4453 816
rect 4487 802 4501 816
rect 4823 802 4837 816
rect 4871 802 4885 816
rect 6047 802 6061 816
rect 6095 802 6109 816
rect 6143 802 6157 816
rect 6335 802 6349 816
rect 6383 802 6397 816
rect 6599 802 6613 816
rect 6887 802 6901 816
rect 71 -17 85 -3
rect 191 -39 205 -25
rect 311 -61 325 -47
rect 431 -83 445 -69
rect 551 -105 565 -91
<< metal2 >>
rect 24 816 36 1641
rect 144 838 156 1644
rect 264 860 276 1646
rect 384 882 396 1650
rect 504 904 516 1658
rect 24 783 36 802
rect 144 799 156 824
rect 264 799 276 846
rect 384 799 396 868
rect 504 799 516 890
rect 648 799 660 846
rect 672 799 684 890
rect 696 799 708 956
rect 792 799 804 824
rect 816 799 828 934
rect 864 799 876 890
rect 912 799 924 912
rect 960 799 972 912
rect 984 799 996 846
rect 1032 799 1044 912
rect 1080 799 1092 934
rect 1104 799 1116 956
rect 1152 799 1164 934
rect 1200 799 1212 912
rect 1224 799 1236 824
rect 1272 799 1284 912
rect 1320 799 1332 934
rect 1344 799 1356 868
rect 1368 799 1380 934
rect 1416 799 1428 912
rect 1440 799 1452 934
rect 1536 799 1548 802
rect 1560 799 1572 846
rect 1680 799 1692 802
rect 1776 799 1788 802
rect 1800 799 1812 824
rect 1944 799 1956 978
rect 2040 799 2052 890
rect 2064 799 2076 1000
rect 2136 799 2148 868
rect 2184 799 2196 912
rect 2256 799 2268 868
rect 2280 799 2292 890
rect 2304 798 2316 1021
rect 2352 799 2364 846
rect 2424 799 2436 934
rect 2472 799 2484 846
rect 2520 799 2532 890
rect 2544 798 2556 1043
rect 2592 799 2604 846
rect 2616 799 2628 868
rect 2664 798 2676 1065
rect 2712 799 2724 846
rect 2736 799 2748 868
rect 2760 797 2772 890
rect 2784 799 2796 956
rect 2856 799 2868 912
rect 2952 799 2964 934
rect 3048 799 3060 956
rect 3144 799 3156 978
rect 3240 799 3252 999
rect 3336 799 3348 912
rect 3432 799 3444 1021
rect 3528 799 3540 934
rect 3552 799 3564 912
rect 3624 799 3636 1043
rect 3720 799 3732 1065
rect 3816 799 3828 956
rect 3888 799 3900 824
rect 3912 799 3924 868
rect 3936 799 3948 890
rect 3960 799 3972 824
rect 4008 799 4020 824
rect 4032 799 4044 802
rect 4152 799 4164 868
rect 4200 799 4212 802
rect 4248 799 4260 868
rect 4272 799 4284 890
rect 4320 799 4332 824
rect 4368 799 4380 802
rect 4392 799 4404 824
rect 4440 799 4452 802
rect 4488 799 4500 802
rect 4704 759 4716 824
rect 4776 760 4788 868
rect 4824 781 4836 802
rect 4872 799 4884 802
rect 4896 799 4908 824
rect 4944 799 4956 824
rect 4992 799 5004 824
rect 5088 799 5100 824
rect 5136 798 5148 824
rect 5160 799 5172 1649
rect 5256 799 5268 824
rect 5280 799 5292 1632
rect 5376 798 5388 824
rect 5400 799 5412 1660
rect 5496 799 5508 824
rect 5520 799 5532 1653
rect 5544 799 5556 824
rect 5592 799 5604 824
rect 5616 799 5628 912
rect 5736 760 5748 846
rect 5760 755 5772 868
rect 5808 799 5820 824
rect 5952 799 5964 846
rect 6000 799 6012 824
rect 6024 799 6036 846
rect 6264 838 6276 1560
rect 6048 799 6060 802
rect 6096 796 6108 802
rect 6144 778 6156 802
rect 6264 798 6276 824
rect 6336 796 6348 802
rect 6384 796 6396 802
rect 6576 799 6588 824
rect 6600 795 6612 802
rect 6696 795 6708 1568
rect 6792 795 6804 1573
rect 6888 795 6900 802
rect 6960 799 6972 1570
rect 7008 799 7020 1569
rect 72 -3 84 0
rect 192 -25 204 12
rect 312 -47 324 0
rect 432 -69 444 0
rect 552 -91 564 0
rect 624 -16 636 15
rect 744 -104 756 15
rect 768 -59 780 0
rect 888 -60 900 0
rect 1248 -15 1260 0
rect 1488 -499 1500 0
rect 1584 -60 1596 0
rect 1563 -496 1575 -152
rect 1632 -496 1644 0
rect 1704 -36 1716 0
rect 1728 -143 1740 0
rect 1824 -123 1836 0
rect 1872 -62 1884 0
rect 1896 -80 1908 0
rect 1920 -102 1932 0
rect 1992 -62 2004 0
rect 2016 -83 2028 0
rect 2112 -60 2124 0
rect 2160 -103 2172 0
rect 2232 -59 2244 0
rect 2376 -83 2388 0
rect 2400 -101 2412 0
rect 2496 -81 2508 0
rect 2640 -108 2652 0
rect 2832 -123 2844 0
rect 2880 -163 2892 0
rect 2928 -123 2940 0
rect 2976 -183 2988 0
rect 3024 -123 3036 0
rect 3072 -123 3084 0
rect 3120 -143 3132 0
rect 3168 -559 3180 0
rect 3216 -83 3228 0
rect 3264 -571 3276 0
rect 3312 -84 3324 0
rect 3308 -564 3320 -133
rect 3360 -566 3372 0
rect 3408 -83 3420 0
rect 3456 -143 3468 0
rect 3504 -83 3516 0
rect 3552 -144 3564 0
rect 3600 -83 3612 0
rect 3648 -163 3660 0
rect 3696 -83 3708 0
rect 3744 -569 3756 0
rect 3792 -82 3804 0
rect 3840 -559 3852 0
rect 4080 -553 4092 0
rect 4128 -35 4140 0
rect 4512 -15 4524 0
rect 4536 -59 4548 0
rect 4147 -566 4159 -133
rect 4203 -564 4215 -113
rect 4584 -554 4596 15
rect 4632 -62 4644 0
rect 4656 -101 4668 0
rect 4752 -51 4764 0
rect 5016 -14 5028 0
rect 5040 -34 5052 0
rect 4657 -558 4669 -173
rect 5208 -579 5220 0
rect 5328 -572 5340 0
rect 5448 -568 5460 0
rect 5664 -553 5676 0
rect 5712 -35 5724 0
rect 5856 -37 5868 0
rect 5880 -59 5892 0
rect 5904 -103 5916 0
rect 6168 -15 6180 18
rect 6216 -569 6228 0
rect 6288 -223 6300 15
rect 6350 -581 6362 -153
rect 6408 -203 6420 3
rect 6504 -619 6516 3
rect 6768 -17 6780 3
rect 6792 -618 6804 0
rect 6960 -608 6972 18
rect 7008 -604 7020 18
use inv inv_0
timestamp 1386238110
transform 1 0 0 0 1 0
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 120 0 1 0
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 240 0 1 0
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 360 0 1 0
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 480 0 1 0
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 600 0 1 0
box 0 0 120 799
use nand3 nand3_1
timestamp 1386234893
transform 1 0 720 0 1 0
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 840 0 1 0
box 0 0 96 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 936 0 1 0
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 1056 0 1 0
box 0 0 120 799
use nand3 nand3_2
timestamp 1386234893
transform 1 0 1176 0 1 0
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1296 0 1 0
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 1392 0 1 0
box 0 0 120 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 1512 0 1 0
box 0 0 144 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 1656 0 1 0
box 0 0 96 799
use nand2 nand2_3
timestamp 1386234792
transform 1 0 1752 0 1 0
box 0 0 96 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 1848 0 1 0
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 1968 0 1 0
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 2088 0 1 0
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 2208 0 1 0
box 0 0 120 799
use nand3 nand3_8
timestamp 1386234893
transform 1 0 2328 0 1 0
box 0 0 120 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 2448 0 1 0
box 0 0 120 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 2568 0 1 0
box 0 0 120 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 2688 0 1 0
box 0 0 120 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 2808 0 1 0
box 0 0 96 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 2904 0 1 0
box 0 0 96 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 3000 0 1 0
box 0 0 96 799
use nand2 nand2_7
timestamp 1386234792
transform 1 0 3096 0 1 0
box 0 0 96 799
use nand2 nand2_8
timestamp 1386234792
transform 1 0 3192 0 1 0
box 0 0 96 799
use nand2 nand2_9
timestamp 1386234792
transform 1 0 3288 0 1 0
box 0 0 96 799
use nand2 nand2_10
timestamp 1386234792
transform 1 0 3384 0 1 0
box 0 0 96 799
use nand2 nand2_11
timestamp 1386234792
transform 1 0 3480 0 1 0
box 0 0 96 799
use nand2 nand2_12
timestamp 1386234792
transform 1 0 3576 0 1 0
box 0 0 96 799
use nand2 nand2_13
timestamp 1386234792
transform 1 0 3672 0 1 0
box 0 0 96 799
use nand2 nand2_14
timestamp 1386234792
transform 1 0 3768 0 1 0
box 0 0 96 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 3864 0 1 0
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 3984 0 1 0
box 0 0 120 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 4104 0 1 0
box 0 0 120 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 4224 0 1 0
box 0 0 120 799
use nor2 nor2_6
timestamp 1386235306
transform 1 0 4344 0 1 0
box 0 0 120 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 4464 0 1 0
box 0 0 144 799
use nor2 nor2_7
timestamp 1386235306
transform 1 0 4608 0 1 0
box 0 0 120 799
use nor2 nor2_8
timestamp 1386235306
transform 1 0 4728 0 1 0
box 0 0 120 799
use nor2 nor2_9
timestamp 1386235306
transform 1 0 4848 0 1 0
box 0 0 120 799
use nor3 nor3_2
timestamp 1386235396
transform 1 0 4968 0 1 0
box 0 0 144 799
use and2 and2_0
timestamp 1386234845
transform 1 0 5112 0 1 0
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 5232 0 1 0
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 5352 0 1 0
box 0 0 120 799
use nand2 nand2_15
timestamp 1386234792
transform 1 0 5472 0 1 0
box 0 0 96 799
use nor2 nor2_10
timestamp 1386235306
transform 1 0 5568 0 1 0
box 0 0 120 799
use nor3 nor3_3
timestamp 1386235396
transform 1 0 5688 0 1 0
box 0 0 144 799
use nor3 nor3_4
timestamp 1386235396
transform 1 0 5832 0 1 0
box 0 0 144 799
use nor3 nor3_5
timestamp 1386235396
transform 1 0 5976 0 1 0
box 0 0 144 799
use nor2 nor2_11
timestamp 1386235306
transform 1 0 6120 0 1 0
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 6240 0 1 0
box 0 0 120 799
use xor2 xor2_0
timestamp 1386237344
transform 1 0 6360 0 1 0
box 0 0 192 799
use xor2 xor2_1
timestamp 1386237344
transform 1 0 6552 0 1 0
box 0 0 192 799
use xor2 xor2_2
timestamp 1386237344
transform 1 0 6744 0 1 0
box 0 0 192 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 6936 0 1 0
box 0 0 48 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 6984 0 1 0
box 0 0 48 799
<< labels >>
rlabel metal1 104 -11 104 -11 1 nA
rlabel metal1 210 -33 210 -33 1 nB
rlabel metal1 336 -53 336 -53 1 nC
rlabel metal1 459 -78 459 -78 1 nD
rlabel metal1 579 -100 579 -100 1 nE
rlabel metal2 5093 801 5093 801 1 N
<< end >>
