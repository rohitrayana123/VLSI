magic
tech c035u
timestamp 1394528018
<< checkpaint >>
rect -5644 499 -2729 3100
rect -5629 495 -2729 499
<< nwell >>
rect -2865 941 -9 1339
rect 10503 941 11367 1339
<< pwell >>
rect -2865 540 -9 941
rect 10503 547 11367 941
<< pohmic >>
rect -2865 616 -2859 626
rect -15 616 -9 626
rect 10503 616 10509 626
rect 11361 616 11367 626
<< nohmic >>
rect -2865 1276 -2859 1286
rect -15 1276 -9 1286
rect 10503 1276 10509 1286
rect 11361 1276 11367 1286
<< psubstratetap >>
rect -2859 616 -15 632
rect 10509 616 11361 632
<< nsubstratetap >>
rect -2859 1270 -15 1286
rect 10509 1270 11361 1286
<< metal1 >>
rect 148 1734 1622 1744
rect 340 1712 1598 1722
rect 532 1690 1574 1700
rect 772 1667 1358 1677
rect 1012 1646 1334 1656
rect 1252 1624 1310 1634
rect 460 1410 1166 1420
rect 268 1388 926 1398
rect 77 1366 733 1376
rect 52 1344 230 1354
rect 244 1344 422 1354
rect 676 1344 902 1354
rect 916 1344 1142 1354
rect -2865 1322 -9 1332
rect 10503 1322 11367 1332
rect -2865 1299 -9 1309
rect 10503 1299 11367 1309
rect -2865 1270 -2859 1286
rect -15 1270 -9 1286
rect -2865 1261 -9 1270
rect 10503 1270 10509 1286
rect 11361 1270 11367 1286
rect 10503 1261 11367 1270
rect -2865 632 -9 641
rect -2865 616 -2859 632
rect -15 616 -9 632
rect 10503 632 11367 641
rect 10503 616 10509 632
rect 11361 616 11367 632
rect -2865 593 -9 603
rect 10503 593 11367 603
rect -2865 570 -9 580
rect 10503 570 11367 580
rect -2865 547 -9 557
rect 10503 547 11367 557
<< m2contact >>
rect 134 1732 148 1746
rect 1622 1732 1636 1746
rect 326 1710 340 1724
rect 1598 1710 1612 1724
rect 518 1688 532 1702
rect 1574 1688 1588 1702
rect 758 1665 772 1679
rect 1358 1665 1372 1679
rect 998 1643 1012 1657
rect 1334 1643 1348 1657
rect 1238 1622 1252 1636
rect 1310 1621 1324 1635
rect 446 1408 460 1422
rect 1166 1408 1180 1422
rect 254 1386 268 1400
rect 926 1386 940 1400
rect 63 1364 77 1378
rect 733 1364 747 1378
rect 38 1342 52 1356
rect 230 1342 244 1356
rect 422 1342 436 1356
rect 662 1342 676 1356
rect 902 1342 916 1356
rect 1142 1342 1156 1356
<< metal2 >>
rect -4329 1339 -4129 1795
rect -4113 1339 -4101 1795
rect -4089 1339 -4077 1795
rect -4065 1339 -4053 1795
rect -4041 1339 -4029 1795
rect 39 1356 51 1795
rect 63 1378 75 1795
rect 39 1339 51 1342
rect 63 1339 75 1364
rect 111 1339 123 1795
rect 135 1339 147 1732
rect 255 1400 267 1795
rect 231 1339 243 1342
rect 255 1339 267 1386
rect 303 1339 315 1795
rect 327 1339 339 1710
rect 447 1422 459 1795
rect 423 1339 435 1342
rect 447 1339 459 1408
rect 495 1339 507 1795
rect 519 1339 531 1688
rect 663 1356 675 1795
rect 663 1339 675 1342
rect 735 1339 747 1364
rect 759 1338 771 1665
rect 903 1339 915 1342
rect 927 1338 939 1386
rect 999 1339 1011 1643
rect 1143 1339 1155 1342
rect 1167 1339 1179 1408
rect 1239 1339 1251 1622
rect 1311 1618 1323 1621
rect 1335 1618 1347 1643
rect 1359 1618 1371 1665
rect 1409 1618 1421 1795
rect 1575 1618 1587 1688
rect 1599 1618 1611 1710
rect 1623 1618 1635 1732
rect 1719 1618 1731 1795
rect 1743 1618 1755 1795
rect 1767 1618 1779 1795
rect 11559 1624 11571 1795
rect 11679 1624 11691 1795
rect 11799 1624 11811 1795
rect 11919 1624 11931 1795
rect 12039 1624 12051 1795
rect 13215 1624 13227 1795
rect 13647 1624 13659 1795
rect 13839 1624 13851 1795
rect 13911 1624 13923 1795
rect 14007 1624 14019 1795
rect 17679 1624 17691 1795
rect 17895 1624 17907 1795
rect 18015 1624 18027 1795
rect 18135 1624 18147 1795
rect 18519 1624 18531 1795
rect -4329 0 -4129 540
rect -4113 0 -4101 540
rect -4089 0 -4077 540
rect -4065 0 -4053 540
rect -4041 0 -4029 540
rect 591 530 603 540
rect 735 530 747 540
rect 591 518 747 530
rect 831 530 843 540
rect 975 530 987 540
rect 831 518 987 530
rect 1071 530 1083 540
rect 1215 530 1227 540
rect 1071 518 1227 530
use leftbuf  leftbuf_1
timestamp 1386242881
transform 1 0 -4329 0 1 540
box 0 0 1464 799
use mux2  mux2_5
timestamp 1386235218
transform 1 0 -9 0 1 540
box 0 0 192 799
use mux2  mux2_4
timestamp 1386235218
transform 1 0 183 0 1 540
box 0 0 192 799
use mux2  mux2_3
timestamp 1386235218
transform 1 0 375 0 1 540
box 0 0 192 799
use tiehigh  tiehigh_2
timestamp 1386086759
transform 1 0 567 0 1 540
box 0 0 48 799
use mux2  mux2_2
timestamp 1386235218
transform 1 0 615 0 1 540
box 0 0 192 799
use tiehigh  tiehigh_1
timestamp 1386086759
transform 1 0 807 0 1 540
box 0 0 48 799
use mux2  mux2_1
timestamp 1386235218
transform 1 0 855 0 1 540
box 0 0 192 799
use tiehigh  tiehigh_0
timestamp 1386086759
transform 1 0 1047 0 1 540
box 0 0 48 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 1095 0 1 540
box 0 0 192 799
use regBlock_decoder  regBlock_decoder_0
timestamp 1394493274
transform 1 0 1287 0 1 0
box 0 0 9216 1618
use ALUDecoder  ALUDecoder_0
timestamp 1394493540
transform 1 0 11367 0 1 143
box 0 -143 7440 1481
use rightend  rightend_0
timestamp 1386235834
transform 1 0 18807 0 1 540
box 0 0 320 799
<< labels >>
rlabel metal2 -4329 0 -4129 0 1 GND!
rlabel metal2 -4113 0 -4101 0 1 SDI
rlabel metal2 -4089 0 -4077 0 1 Test
rlabel metal2 -4065 0 -4053 0 1 Clock
rlabel metal2 -4041 0 -4029 0 1 nReset
rlabel metal2 -4329 1795 -4129 1795 1 GND!
rlabel metal2 -4113 1795 -4101 1795 1 SDI
rlabel metal2 -4089 1795 -4077 1795 1 Test
rlabel metal2 -4065 1795 -4053 1795 1 Clock
rlabel metal2 -4041 1795 -4029 1795 1 nReset
rlabel metal2 1719 1795 1731 1795 5 Ir[2]
rlabel metal2 1743 1795 1755 1795 5 Ir[3]
rlabel metal2 1767 1795 1779 1795 5 Ir[4]
rlabel metal2 447 1795 459 1795 5 Ir[8]
rlabel metal2 255 1795 267 1795 5 Ir[9]
rlabel metal2 63 1795 75 1795 5 Ir[10]
rlabel metal2 663 1795 675 1795 5 RwSel
rlabel metal2 111 1795 123 1795 5 Ir[7]
rlabel metal2 303 1795 315 1795 5 Ir[6]
rlabel metal2 495 1795 507 1795 5 Ir[5]
rlabel metal2 39 1795 51 1795 5 Rs1Sel
rlabel metal2 1409 1795 1421 1795 5 RegWe
rlabel metal2 11559 1795 11571 1795 5 Ir[15]
rlabel metal2 11679 1795 11691 1795 5 Ir[14]
rlabel metal2 11799 1795 11811 1795 5 Ir[13]
rlabel metal2 11919 1795 11931 1795 5 Ir[12]
rlabel metal2 12039 1795 12051 1795 5 Ir[11]
rlabel metal2 13215 1795 13227 1795 5 CFlag
rlabel metal2 13647 1795 13659 1795 5 Flags[2]
rlabel metal2 13839 1795 13851 1795 5 Flags[1]
rlabel metal2 13911 1795 13923 1795 5 Flags[3]
rlabel metal2 14007 1795 14019 1795 5 Flagss[0]
rlabel metal2 18135 1795 18147 1795 5 Ir[0]
rlabel metal2 18015 1795 18027 1795 5 Ir[1]
rlabel metal2 17895 1795 17907 1795 5 Ir[2]
rlabel metal2 17679 1795 17691 1795 5 Ir[3]
rlabel metal2 18519 1795 18531 1795 5 AluEn
<< end >>
