magic
tech c035u
timestamp 1395340701
<< metal1 >>
rect 433 20600 14996 20610
rect 456 20576 15189 20586
rect 479 20552 15381 20562
rect 502 20528 15573 20538
rect 525 20504 15765 20514
rect 548 20480 4580 20490
rect 571 20456 5012 20466
rect 594 20432 5396 20442
rect 617 20408 4628 20418
rect 640 20384 5060 20394
rect 663 20360 5444 20370
rect 686 20336 7584 20346
rect 709 20312 7560 20322
rect 7574 20312 22772 20322
rect 732 20288 7536 20298
rect 7550 20288 22964 20298
rect 755 20264 23084 20274
rect 778 20240 23204 20250
rect 23997 18891 24189 18901
rect 3514 18780 3525 18790
rect 414 17893 419 17903
rect 433 17893 784 17903
rect 414 17861 784 17871
rect 414 17827 784 17837
rect 3477 17827 3525 17837
rect 23997 17827 24189 17837
rect 3477 17805 3525 17815
rect 23997 17715 24189 17725
rect 3514 17604 3525 17614
rect 414 16717 442 16727
rect 456 16717 784 16727
rect 414 16685 784 16695
rect 414 16651 784 16661
rect 3477 16651 3525 16661
rect 23997 16651 24189 16661
rect 3477 16629 3525 16639
rect 23997 16539 24189 16549
rect 3514 16428 3525 16438
rect 414 15541 465 15551
rect 479 15541 784 15551
rect 414 15509 784 15519
rect 414 15475 784 15485
rect 3477 15475 3525 15485
rect 23997 15475 24189 15485
rect 3477 15453 3525 15463
rect 23997 15363 24189 15373
rect 3514 15252 3525 15262
rect 414 14365 488 14375
rect 502 14365 784 14375
rect 414 14333 784 14343
rect 414 14299 784 14309
rect 3477 14299 3525 14309
rect 23997 14299 24189 14309
rect 3477 14277 3525 14287
rect 23997 14187 24189 14197
rect 3514 14076 3525 14086
rect 414 13189 511 13199
rect 525 13189 784 13199
rect 414 13157 784 13167
rect 414 13123 784 13133
rect 3477 13123 3525 13133
rect 23997 13123 24189 13133
rect 3477 13101 3525 13111
rect 23997 13011 24189 13021
rect 3514 12900 3525 12910
rect 414 12013 534 12023
rect 548 12013 784 12023
rect 414 11981 784 11991
rect 414 11947 784 11957
rect 3477 11947 3525 11957
rect 23997 11947 24189 11957
rect 3477 11925 3525 11935
rect 23997 11835 24189 11845
rect 3514 11724 3525 11734
rect 414 10837 557 10847
rect 571 10837 784 10847
rect 414 10805 784 10815
rect 414 10771 784 10781
rect 3477 10771 3525 10781
rect 23997 10771 24189 10781
rect 3477 10749 3525 10759
rect 23997 10659 24189 10669
rect 3514 10548 3525 10558
rect 414 9661 580 9671
rect 594 9661 784 9671
rect 414 9629 784 9639
rect 414 9595 784 9605
rect 3477 9595 3525 9605
rect 23997 9595 24189 9605
rect 3477 9573 3525 9583
rect 23997 9483 24189 9493
rect 3514 9372 3525 9382
rect 414 8485 603 8495
rect 617 8485 784 8495
rect 414 8453 784 8463
rect 414 8419 784 8429
rect 3477 8419 3525 8429
rect 23997 8419 24189 8429
rect 3477 8397 3525 8407
rect 23997 8307 24189 8317
rect 3514 8196 3525 8206
rect 414 7309 626 7319
rect 640 7309 784 7319
rect 414 7277 784 7287
rect 414 7243 784 7253
rect 3477 7243 3525 7253
rect 23997 7243 24189 7253
rect 3477 7221 3525 7231
rect 23997 7131 24189 7141
rect 3514 7020 3525 7030
rect 414 6133 649 6143
rect 663 6133 784 6143
rect 414 6101 784 6111
rect 414 6067 784 6077
rect 3477 6067 3525 6077
rect 23997 6067 24189 6077
rect 3477 6045 3525 6055
rect 23997 5955 24189 5965
rect 3514 5844 3525 5854
rect 414 4957 672 4967
rect 686 4957 784 4967
rect 414 4925 784 4935
rect 414 4891 784 4901
rect 3477 4891 3525 4901
rect 23997 4891 24189 4901
rect 3477 4869 3525 4879
rect 23997 4779 24189 4789
rect 3514 4668 3525 4678
rect 414 3781 695 3791
rect 709 3781 784 3791
rect 414 3749 784 3759
rect 414 3715 784 3725
rect 3477 3715 3525 3725
rect 23997 3715 24189 3725
rect 3477 3693 3525 3703
rect 23997 3603 24189 3613
rect 3514 3492 3525 3502
rect 414 2605 718 2615
rect 732 2605 784 2615
rect 414 2573 784 2583
rect 414 2539 784 2549
rect 3477 2539 3525 2549
rect 23997 2539 24189 2549
rect 3477 2517 3525 2527
rect 23997 2427 24189 2437
rect 3514 2316 3525 2326
rect 414 1429 741 1439
rect 755 1429 784 1439
rect 414 1397 784 1407
rect 414 1363 784 1373
rect 3477 1363 3525 1373
rect 23997 1363 24189 1373
rect 3477 1341 3525 1351
rect 23997 1251 24189 1261
rect 3514 1140 3525 1150
rect 414 253 764 263
rect 778 253 784 263
rect 414 221 784 231
rect 414 187 784 197
rect 3477 187 3525 197
rect 23997 187 24189 197
rect 3477 165 3525 175
rect 2474 72 17684 82
rect 17698 72 20348 82
rect 20362 72 20395 82
rect 20409 72 20444 82
rect 20458 72 20492 82
rect 20506 72 20540 82
rect 20554 72 20588 82
rect 20602 72 20636 82
rect 20650 72 20684 82
rect 20698 72 20996 82
rect 21010 72 21044 82
rect 21058 72 21091 82
rect 21105 72 21140 82
rect 21154 72 21452 82
rect 21466 72 21500 82
rect 21514 72 21884 82
rect 21898 72 25245 82
rect 989 51 3740 61
<< m2contact >>
rect 419 20598 433 20612
rect 14996 20599 15010 20613
rect 442 20574 456 20588
rect 15189 20574 15203 20588
rect 465 20550 479 20564
rect 15381 20550 15395 20564
rect 488 20526 502 20540
rect 15573 20526 15587 20540
rect 511 20502 525 20516
rect 15765 20502 15779 20517
rect 534 20478 548 20492
rect 4580 20478 4594 20492
rect 557 20454 571 20468
rect 5012 20454 5026 20468
rect 580 20430 594 20444
rect 5396 20430 5410 20444
rect 603 20406 617 20420
rect 4628 20406 4642 20420
rect 626 20382 640 20396
rect 5060 20382 5074 20396
rect 649 20358 663 20372
rect 5444 20358 5458 20372
rect 672 20334 686 20348
rect 7584 20334 7598 20348
rect 695 20310 709 20324
rect 7560 20310 7574 20324
rect 22772 20310 22786 20324
rect 718 20286 732 20300
rect 7536 20286 7550 20300
rect 22964 20285 22978 20299
rect 741 20262 755 20276
rect 23084 20262 23098 20276
rect 764 20238 778 20252
rect 23204 20238 23218 20252
rect 3500 18778 3514 18792
rect 419 17891 433 17905
rect 3500 17602 3514 17616
rect 442 16715 456 16729
rect 3500 16426 3514 16440
rect 465 15539 479 15553
rect 3500 15250 3514 15264
rect 488 14363 502 14377
rect 3500 14074 3514 14088
rect 511 13187 525 13201
rect 3500 12898 3514 12912
rect 534 12011 548 12025
rect 3500 11722 3514 11736
rect 557 10835 571 10849
rect 3500 10546 3514 10560
rect 580 9659 594 9673
rect 3500 9370 3514 9384
rect 603 8483 617 8497
rect 3500 8194 3514 8208
rect 626 7307 640 7321
rect 3500 7018 3514 7032
rect 649 6131 663 6145
rect 3500 5842 3514 5856
rect 672 4955 686 4969
rect 3500 4666 3514 4680
rect 695 3779 709 3793
rect 3500 3490 3514 3504
rect 718 2603 732 2617
rect 3500 2314 3514 2328
rect 741 1427 755 1441
rect 3500 1138 3514 1152
rect 764 251 778 265
rect 17684 70 17698 84
rect 20348 70 20362 84
rect 20395 70 20409 84
rect 20444 70 20458 84
rect 20492 70 20506 84
rect 20540 70 20554 84
rect 20588 70 20602 84
rect 20636 70 20650 84
rect 20684 70 20698 84
rect 20996 70 21010 84
rect 21044 70 21058 84
rect 21091 70 21105 84
rect 21140 70 21154 84
rect 21452 70 21466 84
rect 21500 70 21514 84
rect 21884 70 21898 84
rect 25245 70 25259 84
rect 975 49 989 63
rect 3740 48 3754 62
<< metal2 >>
rect 420 17905 432 20598
rect 443 16729 455 20574
rect 466 15553 478 20550
rect 489 14377 501 20526
rect 512 13201 524 20502
rect 535 12025 547 20478
rect 558 10849 570 20454
rect 581 9673 593 20430
rect 604 8497 616 20406
rect 627 7321 639 20382
rect 650 6145 662 20358
rect 673 4969 685 20334
rect 696 3793 708 20310
rect 719 2617 731 20286
rect 742 1441 754 20262
rect 765 265 777 20238
rect 789 20229 989 20615
rect 1005 20229 1017 20615
rect 1029 20229 1041 20615
rect 1053 20229 1065 20615
rect 1077 20229 1089 20615
rect 4557 20229 4569 20615
rect 4581 20229 4593 20478
rect 4629 20229 4641 20406
rect 4797 20229 4809 20615
rect 5013 20229 5025 20454
rect 5061 20229 5073 20382
rect 5397 20229 5409 20430
rect 5445 20229 5457 20358
rect 5757 20229 5769 20615
rect 5949 20229 5961 20615
rect 6983 20229 6995 20615
rect 7537 20229 7549 20286
rect 7561 20229 7573 20310
rect 7585 20229 7597 20334
rect 14974 20229 14986 20615
rect 14998 20229 15010 20599
rect 15190 20229 15202 20574
rect 15238 20229 15250 20615
rect 15382 20229 15394 20550
rect 15574 20229 15586 20526
rect 15766 20229 15778 20502
rect 15958 20229 15970 20615
rect 17757 20229 17769 20615
rect 17949 20229 17961 20615
rect 18021 20229 18033 20615
rect 18117 20229 18129 20615
rect 22773 20229 22785 20310
rect 22965 20229 22977 20285
rect 23085 20229 23097 20262
rect 23205 20229 23217 20238
rect 25244 20229 25444 20615
rect 24045 18885 24057 18908
rect 3501 18708 3513 18778
rect 24045 17709 24057 17843
rect 3501 17532 3513 17602
rect 24045 16533 24057 16667
rect 3501 16356 3513 16426
rect 24045 15357 24057 15491
rect 3501 15180 3513 15250
rect 24045 14181 24057 14315
rect 3501 14004 3513 14074
rect 24045 13005 24057 13139
rect 3501 12828 3513 12898
rect 24045 11829 24057 11963
rect 3501 11652 3513 11722
rect 24045 10653 24057 10787
rect 3501 10476 3513 10546
rect 24045 9477 24057 9611
rect 3501 9300 3513 9370
rect 24045 8301 24057 8435
rect 3501 8124 3513 8194
rect 24045 7125 24057 7259
rect 3501 6948 3513 7018
rect 24045 5949 24057 6083
rect 3501 5772 3513 5842
rect 24045 4773 24057 4907
rect 3501 4596 3513 4666
rect 24045 3597 24057 3731
rect 3501 3420 3513 3490
rect 24045 2421 24057 2555
rect 3501 2244 3513 2314
rect 24045 1245 24057 1379
rect 3501 1068 3513 1138
rect 789 63 989 92
rect 789 49 975 63
rect 789 43 989 49
rect 1005 43 1017 92
rect 1029 43 1041 92
rect 1053 43 1065 92
rect 1077 43 1089 92
rect 2349 43 2361 92
rect 2541 43 2553 92
rect 3333 43 3345 92
rect 3741 62 3753 92
rect 3885 43 3897 92
rect 4101 43 4113 92
rect 4845 43 4857 92
rect 5013 43 5025 92
rect 5397 43 5409 92
rect 5589 43 5601 103
rect 24045 92 24057 203
rect 5805 43 5817 92
rect 6549 43 6561 92
rect 6717 43 6729 92
rect 16125 43 16137 92
rect 16317 43 16329 92
rect 16557 43 16569 92
rect 17205 86 17217 92
rect 17397 86 17409 92
rect 17205 74 17409 86
rect 17685 84 17697 92
rect 20349 84 20361 92
rect 20397 84 20409 92
rect 20445 84 20457 92
rect 20493 84 20505 92
rect 20541 84 20553 92
rect 20589 84 20601 92
rect 20637 84 20649 92
rect 20685 84 20697 92
rect 20997 84 21009 92
rect 21045 84 21057 92
rect 21093 84 21105 92
rect 21141 84 21153 92
rect 21453 84 21465 92
rect 21501 84 21513 92
rect 21885 84 21897 92
rect 24261 43 24273 92
rect 25005 43 25017 92
rect 25245 84 25445 92
rect 25259 70 25445 84
rect 25245 43 25445 70
use slice17 slice17_0
timestamp 1395339964
transform 1 0 789 0 1 18908
box 0 0 24656 1321
use leftbuf_slice leftbuf_slice_0
array 0 0 1685 0 15 1176
timestamp 1394551156
transform 1 0 784 0 1 98
box 0 -6 1685 1170
use IrAA IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 2469 0 1 9611
box 0 -111 1008 1065
use tielow tielow_0
timestamp 1386086605
transform 1 0 3477 0 1 17909
box 0 0 48 799
use tielow tielow_1
timestamp 1386086605
transform 1 0 3477 0 1 16733
box 0 0 48 799
use tielow tielow_2
timestamp 1386086605
transform 1 0 3477 0 1 15557
box 0 0 48 799
use tielow tielow_3
timestamp 1386086605
transform 1 0 3477 0 1 14381
box 0 0 48 799
use tielow tielow_4
timestamp 1386086605
transform 1 0 3477 0 1 13205
box 0 0 48 799
use tielow tielow_5
timestamp 1386086605
transform 1 0 3477 0 1 12029
box 0 0 48 799
use tielow tielow_6
timestamp 1386086605
transform 1 0 3477 0 1 10853
box 0 0 48 799
use tielow tielow_7
timestamp 1386086605
transform 1 0 3477 0 1 9677
box 0 0 48 799
use IrBA IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 2469 0 1 6083
box 0 -111 1008 1065
use tielow tielow_8
timestamp 1386086605
transform 1 0 3477 0 1 8501
box 0 0 48 799
use tielow tielow_9
timestamp 1386086605
transform 1 0 3477 0 1 7325
box 0 0 48 799
use tielow tielow_10
timestamp 1386086605
transform 1 0 3477 0 1 6149
box 0 0 48 799
use IrBB IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 2469 0 1 204
box 0 -112 1008 1064
use tiehigh tiehigh_0
timestamp 1386086759
transform 1 0 3477 0 1 4973
box 0 0 48 799
use tielow tielow_12
timestamp 1386086605
transform 1 0 3477 0 1 3797
box 0 0 48 799
use tielow tielow_13
timestamp 1386086605
transform 1 0 3477 0 1 2621
box 0 0 48 799
use tielow tielow_14
timestamp 1386086605
transform 1 0 3477 0 1 1445
box 0 0 48 799
use tielow tielow_15
timestamp 1386086605
transform 1 0 3477 0 1 269
box 0 0 48 799
use Datapath_slice Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394725603
transform 1 0 3525 0 1 92
box 0 0 20472 1176
use LLIcell_U LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1394841956
transform 1 0 23997 0 1 9611
box 0 0 192 1042
use LLIcell_L LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23997 0 1 203
box 0 0 192 1042
use Datapath_end Datapath_end_0
array 0 0 1256 0 15 1176
timestamp 1394720841
transform 1 0 24189 0 1 92
box 0 0 1256 1176
<< labels >>
rlabel metal1 24093 1257 24093 1257 1 Aluout[0]
rlabel metal2 425 20303 425 20303 1 Ir[15]
rlabel metal2 449 20302 449 20302 1 Ir[14]
rlabel metal2 472 20302 472 20302 1 Ir[13]
rlabel metal2 495 20303 495 20303 1 Ir[12]
rlabel metal2 518 20303 518 20303 1 Ir[11]
rlabel metal2 541 20302 541 20302 1 Ir[10]
rlabel metal2 564 20303 564 20303 1 Ir[9]
rlabel metal2 587 20303 587 20303 1 Ir[8]
rlabel metal2 610 20305 610 20305 1 Ir[7]
rlabel metal2 633 20306 633 20306 1 Ir[6]
rlabel metal2 656 20307 656 20307 1 Ir[5]
rlabel metal2 679 20308 679 20308 1 Ir[4]
rlabel metal2 702 20307 702 20307 1 Ir[3]
rlabel metal2 23211 20233 23211 20233 1 Ir[0]
rlabel metal2 23090 20255 23090 20255 1 Ir[1]
rlabel metal2 22970 20280 22970 20280 1 Ir[2]
rlabel metal2 22779 20305 22779 20305 1 Ir[3]
rlabel metal2 15387 20544 15387 20544 1 Ir[13]
rlabel metal2 15580 20520 15580 20520 1 Ir[12]
rlabel metal2 15772 20495 15772 20495 1 Ir[11]
rlabel metal2 15194 20567 15194 20567 1 Ir[14]
rlabel metal2 15003 20592 15003 20592 1 Ir[15]
rlabel metal2 7541 20278 7541 20278 1 Ir[2]
rlabel metal2 7567 20302 7567 20302 1 Ir[3]
rlabel metal2 7590 20326 7590 20326 1 Ir[4]
rlabel metal2 4635 20398 4635 20398 1 Ir[7]
rlabel metal2 4586 20471 4586 20471 1 Ir[10]
rlabel metal2 5067 20375 5067 20375 1 Ir[6]
rlabel metal2 5018 20446 5018 20446 1 Ir[9]
rlabel metal2 5402 20423 5402 20423 1 Ir[8]
rlabel metal2 5452 20352 5452 20352 1 Ir[5]
rlabel metal1 414 187 414 197 3 SysBus[0]
rlabel metal1 414 1363 414 1373 3 SysBus[1]
rlabel metal1 414 2539 414 2549 3 SysBus[2]
rlabel metal1 414 3715 414 3725 3 SysBus[3]
rlabel metal1 414 4891 414 4901 3 SysBus[4]
rlabel metal1 414 6067 414 6077 3 SysBus[5]
rlabel metal1 414 7243 414 7253 3 SysBus[6]
rlabel metal1 414 8419 414 8429 3 SysBus[7]
rlabel metal1 414 9595 414 9605 3 SysBus[8]
rlabel metal1 414 10771 414 10781 3 SysBus[9]
rlabel metal1 414 11947 414 11957 3 SysBus[10]
rlabel metal1 414 13123 414 13133 3 SysBus[11]
rlabel metal1 414 14299 414 14309 3 SysBus[12]
rlabel metal1 414 15475 414 15485 3 SysBus[13]
rlabel metal1 414 16651 414 16661 3 SysBus[14]
rlabel metal1 414 17827 414 17837 3 SysBus[15]
rlabel metal1 414 253 414 263 3 Ir[0]
rlabel metal1 414 1429 414 1439 3 Ir[1]
rlabel metal1 414 2605 414 2615 3 Ir[2]
rlabel metal1 414 3781 414 3791 3 Ir[3]
rlabel metal1 414 4957 414 4967 3 Ir[4]
rlabel metal1 414 6133 414 6143 3 Ir[5]
rlabel metal1 414 7309 414 7319 3 Ir[6]
rlabel metal1 414 8485 414 8495 3 Ir[7]
rlabel metal1 414 9661 414 9671 3 Ir[8]
rlabel metal1 414 10837 414 10847 3 Ir[9]
rlabel metal1 414 12013 414 12023 3 Ir[10]
rlabel metal1 414 13189 414 13199 3 Ir[11]
rlabel metal1 414 14365 414 14375 3 Ir[12]
rlabel metal1 414 15541 414 15551 3 Ir[13]
rlabel metal1 414 16717 414 16727 3 Ir[14]
rlabel metal1 414 17893 414 17903 3 Ir[15]
rlabel metal1 414 221 414 231 3 DataIn[0]
rlabel metal1 414 17861 414 17871 3 DataIn[15]
rlabel metal1 414 16685 414 16695 3 DataIn[14]
rlabel metal1 414 15509 414 15519 3 DataIn[13]
rlabel metal1 414 14333 414 14343 3 DataIn[12]
rlabel metal1 414 13157 414 13167 3 DataIn[11]
rlabel metal1 414 11981 414 11991 3 DataIn[10]
rlabel metal1 414 10805 414 10815 3 DataIn[9]
rlabel metal1 414 9629 414 9639 3 DataIn[8]
rlabel metal1 414 8453 414 8463 3 DataIn[7]
rlabel metal1 414 7277 414 7287 3 DataIn[6]
rlabel metal1 414 6101 414 6111 3 DataIn[5]
rlabel metal1 414 4925 414 4935 3 DataIn[4]
rlabel metal1 414 3749 414 3759 3 DataIn[3]
rlabel metal1 414 2573 414 2583 3 DataIn[2]
rlabel metal1 414 1397 414 1407 3 DataIn[1]
rlabel metal2 6983 20615 6995 20615 5 RegWe
rlabel metal2 1005 20615 1017 20615 5 SDO
rlabel metal2 789 20615 989 20615 5 Vdd!
rlabel metal2 1077 20615 1089 20615 1 nReset
rlabel metal2 1053 20615 1065 20615 1 Clock
rlabel metal2 1029 20615 1041 20615 1 Test
rlabel metal2 25244 20615 25444 20615 1 GND!
rlabel metal2 18117 20615 18129 20615 5 Flags[0]
rlabel metal2 18021 20615 18033 20615 5 Flags[3]
rlabel metal2 17949 20615 17961 20615 5 Flags[1]
rlabel metal2 17757 20615 17769 20615 5 Flags[2]
rlabel metal2 15238 20615 15250 20615 5 AluOR[0]
rlabel metal2 14974 20615 14986 20615 5 AluOR[1]
rlabel metal2 15958 20615 15970 20615 5 CFlag
rlabel metal2 4557 20615 4569 20615 5 Rs1Sel[0]
rlabel metal2 4797 20615 4809 20615 5 Rs1Sel[1]
rlabel metal2 5757 20615 5769 20615 5 RwSel[0]
rlabel metal2 5949 20615 5961 20615 5 RwSel[1]
rlabel metal2 3885 43 3897 43 1 LrSel
rlabel metal2 4101 43 4113 43 1 LrWe
rlabel metal2 4845 43 4857 43 1 LrEn
rlabel metal2 5013 43 5025 43 1 PcSel[0]
rlabel metal2 5397 43 5409 43 1 PcSel[1]
rlabel metal2 24261 43 24273 43 1 AluWe
rlabel metal2 25005 43 25017 43 1 AluEn
rlabel metal2 25245 43 25445 43 1 GND!
rlabel metal2 789 43 989 43 1 Vdd!
rlabel metal2 1005 43 1017 43 1 SDI
rlabel metal2 1029 43 1041 43 1 Test
rlabel metal2 1053 43 1065 43 1 Clock
rlabel metal2 1077 43 1089 43 1 nReset
rlabel metal2 3333 43 3345 43 1 ImmSel
rlabel metal2 2541 43 2553 43 1 IrWe
rlabel metal2 2349 43 2361 43 1 MemEn
rlabel metal2 5805 43 5817 43 1 PcWe
rlabel metal2 5589 43 5601 43 1 PcSel[2]
rlabel metal2 6549 43 6561 43 1 PcEn
rlabel metal2 6717 43 6729 43 1 WdSel
rlabel metal2 16125 43 16137 43 1 Op1Sel
rlabel metal2 16317 43 16329 43 1 Op2Sel[0]
rlabel metal2 16557 43 16569 43 1 Op2Sel[1]
<< end >>
