../../../Design/Implementation/verilog/behavioural/cpu.sv