magic
tech c035u
timestamp 1396390031
<< metal1 >>
rect 0 1094 192 1104
rect 0 938 119 948
rect 0 97 71 107
rect 157 97 192 107
rect 0 29 192 39
<< m2contact >>
rect 119 936 133 950
rect 71 95 85 109
rect 143 95 157 109
<< metal2 >>
rect 48 911 60 1111
rect 120 911 132 936
rect 48 0 60 112
rect 72 109 84 112
rect 144 109 156 112
use mux2 mux2_0
timestamp 1386235218
transform 1 0 0 0 1 112
box 0 0 192 799
<< labels >>
rlabel metal1 0 97 0 107 3 LLIIn
rlabel metal1 192 97 192 107 1 ALUOut
rlabel metal1 0 938 0 948 3 B
rlabel metal2 48 1111 60 1111 5 LLI
rlabel metal1 192 1094 192 1104 7 ALUOut
rlabel metal1 0 1094 0 1104 3 ALUOut
rlabel metal1 0 29 0 39 3 SysBus
rlabel metal1 192 29 192 39 7 SysBus
rlabel metal2 48 0 60 0 1 LLI
<< end >>
