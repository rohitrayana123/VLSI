magic
tech c035u
timestamp 1398757585
<< nwell >>
rect 26595 1419 27050 1817
<< pwell >>
rect 26595 1018 27050 1419
<< pohmic >>
rect 27041 1094 27050 1104
<< nohmic >>
rect 27046 1754 27050 1764
<< psubstratetap >>
rect 26654 1329 26670 1345
rect 26780 1329 26796 1345
rect 26906 1329 26922 1345
rect 26595 1094 27041 1110
<< nsubstratetap >>
rect 26595 1748 27046 1764
<< metal1 >>
rect 15712 8420 15730 8434
rect 16876 8422 20282 8432
rect 13816 8396 13834 8410
rect 14680 8398 22766 8408
rect 2296 8374 17726 8384
rect 84 8350 23138 8360
rect 84 8326 1730 8336
rect 2008 8326 2450 8336
rect 3544 8326 7562 8336
rect 9244 8326 19154 8336
rect 19396 8326 20546 8336
rect 21916 8326 22154 8336
rect 24436 8326 25010 8336
rect 2152 8302 3554 8312
rect 3568 8302 22010 8312
rect 22024 8302 25286 8312
rect 2428 8278 7970 8288
rect 8344 8278 9266 8288
rect 9472 8278 12674 8288
rect 12880 8278 24446 8288
rect 4132 8254 7946 8264
rect 10768 8254 26126 8264
rect 27040 8254 27050 8264
rect 4216 8230 27074 8240
rect 4984 8206 8810 8216
rect 10948 8206 25778 8216
rect 5836 8182 6074 8192
rect 6280 8180 6298 8194
rect 7540 8182 9938 8192
rect 11464 8182 19406 8192
rect 20704 8180 20722 8194
rect 22408 8180 22426 8194
rect 24808 8182 27122 8192
rect 11800 8158 20930 8168
rect 27112 8158 27445 8168
rect 12652 8134 24146 8144
rect 27088 8134 27445 8144
rect 15196 8110 23402 8120
rect 27064 8110 27445 8120
rect 17716 8084 17734 8098
rect 18664 8086 27445 8096
rect 19432 8062 27098 8072
rect 27136 8062 27445 8072
rect 15832 7229 15962 7239
rect 14896 7205 14930 7215
rect 15040 7205 27002 7215
rect 14152 7181 18170 7191
rect 13240 7157 13346 7167
rect 13912 7157 14138 7167
rect 14632 7157 20294 7167
rect 13192 7133 13250 7143
rect 13816 7133 23594 7143
rect 13120 7109 24146 7119
rect 13072 7085 22250 7095
rect 13024 7061 24674 7071
rect 12976 7037 22346 7047
rect 12712 7013 14186 7023
rect 14200 7013 26234 7023
rect 12496 6989 12530 6999
rect 12664 6989 21506 6999
rect 12040 6965 12146 6975
rect 12208 6965 23978 6975
rect 11704 6941 18194 6951
rect 11368 6917 26762 6927
rect 10528 6893 21314 6903
rect 10456 6869 12938 6879
rect 13000 6869 16922 6879
rect 10384 6845 10442 6855
rect 10504 6845 10562 6855
rect 10648 6845 16442 6855
rect 10312 6821 11402 6831
rect 11608 6821 18026 6831
rect 9664 6797 17834 6807
rect 9448 6773 15050 6783
rect 15784 6773 23714 6783
rect 9376 6749 19826 6759
rect 19840 6749 22778 6759
rect 9232 6725 21290 6735
rect 9040 6701 9050 6711
rect 9184 6701 18770 6711
rect 8968 6677 17042 6687
rect 8920 6653 10802 6663
rect 10888 6653 11042 6663
rect 11104 6653 23450 6663
rect 8776 6629 13946 6639
rect 14008 6629 15986 6639
rect 8584 6605 26774 6615
rect 8464 6581 13994 6591
rect 14008 6581 23186 6591
rect 8272 6557 16130 6567
rect 16384 6557 23150 6567
rect 8224 6533 23858 6543
rect 7816 6509 18602 6519
rect 7792 6485 18722 6495
rect 20344 6485 23714 6495
rect 7768 6461 8210 6471
rect 8224 6461 8714 6471
rect 8728 6461 12626 6471
rect 12640 6461 13298 6471
rect 13312 6461 19826 6471
rect 19840 6461 22322 6471
rect 22336 6461 25202 6471
rect 25216 6461 25874 6471
rect 7528 6437 23498 6447
rect 7432 6413 15938 6423
rect 16264 6413 20330 6423
rect 7384 6389 26522 6399
rect 7312 6365 13298 6375
rect 13672 6365 13682 6375
rect 13768 6365 15746 6375
rect 15808 6365 20138 6375
rect 20152 6365 22010 6375
rect 7192 6341 12122 6351
rect 12136 6341 13394 6351
rect 13408 6341 26978 6351
rect 7096 6317 21098 6327
rect 7000 6293 8474 6303
rect 8536 6293 10394 6303
rect 10408 6293 10922 6303
rect 10936 6293 12170 6303
rect 12184 6293 15122 6303
rect 15136 6293 21074 6303
rect 21088 6293 21818 6303
rect 6904 6269 7490 6279
rect 7504 6269 21554 6279
rect 6736 6245 7346 6255
rect 7408 6245 25346 6255
rect 6712 6221 21626 6231
rect 22216 6221 22370 6231
rect 6688 6197 11834 6207
rect 11848 6197 22754 6207
rect 22768 6197 25226 6207
rect 26440 6197 26690 6207
rect 6616 6173 26426 6183
rect 6592 6149 14738 6159
rect 14752 6149 26210 6159
rect 6568 6125 9386 6135
rect 9400 6125 14690 6135
rect 14704 6125 22202 6135
rect 6376 6101 14786 6111
rect 14872 6101 25658 6111
rect 6280 6077 8426 6087
rect 8440 6077 11978 6087
rect 11992 6077 12722 6087
rect 12736 6077 15578 6087
rect 15592 6077 16586 6087
rect 16600 6077 16682 6087
rect 16696 6077 19802 6087
rect 22816 6077 23306 6087
rect 6184 6053 14666 6063
rect 14680 6053 22802 6063
rect 6016 6029 24866 6039
rect 5968 6005 13706 6015
rect 13720 6005 22826 6015
rect 5920 5981 11666 5991
rect 11800 5981 26810 5991
rect 5896 5957 23930 5967
rect 5824 5933 19082 5943
rect 19096 5933 25226 5943
rect 5800 5909 18146 5919
rect 18160 5909 18434 5919
rect 18448 5909 21530 5919
rect 21544 5909 23906 5919
rect 5728 5885 21410 5895
rect 5704 5861 9218 5871
rect 9232 5861 11330 5871
rect 11344 5861 11546 5871
rect 11560 5861 13010 5871
rect 13024 5861 13370 5871
rect 13384 5861 26570 5871
rect 5512 5837 9362 5847
rect 9376 5837 26906 5847
rect 5488 5813 9842 5823
rect 9856 5813 15434 5823
rect 15448 5813 18938 5823
rect 18952 5813 18986 5823
rect 19000 5813 20426 5823
rect 20440 5813 23942 5823
rect 26344 5813 26534 5823
rect 5464 5789 13322 5799
rect 13624 5789 18866 5799
rect 18880 5789 19730 5799
rect 19744 5789 26330 5799
rect 5344 5765 10970 5775
rect 10984 5765 13562 5775
rect 13576 5765 16442 5775
rect 16456 5765 16754 5775
rect 16768 5765 18482 5775
rect 18496 5765 21026 5775
rect 21040 5765 21842 5775
rect 21856 5765 26738 5775
rect 5056 5741 19538 5751
rect 4936 5717 22922 5727
rect 4792 5693 5978 5703
rect 5992 5693 13922 5703
rect 13936 5693 23474 5703
rect 25048 5693 26018 5703
rect 4720 5669 7898 5679
rect 7912 5669 8690 5679
rect 8704 5669 19634 5679
rect 19648 5669 20138 5679
rect 20152 5669 22922 5679
rect 22936 5669 24362 5679
rect 24376 5669 25034 5679
rect 4648 5645 15026 5655
rect 15040 5645 22514 5655
rect 22528 5645 25418 5655
rect 4552 5621 8402 5631
rect 8416 5621 10274 5631
rect 10288 5621 16562 5631
rect 16840 5621 21674 5631
rect 4504 5597 4658 5607
rect 4672 5597 10058 5607
rect 10072 5597 13202 5607
rect 13216 5597 16634 5607
rect 16648 5597 16946 5607
rect 16960 5597 22322 5607
rect 4432 5573 4946 5583
rect 4960 5573 16178 5583
rect 16192 5573 17594 5583
rect 4360 5549 8906 5559
rect 8920 5549 9986 5559
rect 10000 5549 13658 5559
rect 13672 5549 16850 5559
rect 16864 5549 19250 5559
rect 19264 5549 21050 5559
rect 21064 5549 22250 5559
rect 4240 5525 25298 5535
rect 4168 5501 10010 5511
rect 10024 5501 12626 5511
rect 12688 5501 27026 5511
rect 4144 5477 17786 5487
rect 17800 5477 23234 5487
rect 23248 5477 24170 5487
rect 4120 5453 7586 5463
rect 7600 5453 11426 5463
rect 11440 5453 12698 5463
rect 12712 5453 18626 5463
rect 18640 5453 19658 5463
rect 19672 5453 21122 5463
rect 4096 5429 18578 5439
rect 4072 5405 5810 5415
rect 5824 5405 8378 5415
rect 8392 5405 22538 5415
rect 3880 5381 22346 5391
rect 3832 5357 3890 5367
rect 3952 5357 11378 5367
rect 11392 5357 16274 5367
rect 16336 5357 20642 5367
rect 3808 5333 4010 5343
rect 4024 5333 6122 5343
rect 6136 5333 7874 5343
rect 7888 5333 8834 5343
rect 8848 5333 10298 5343
rect 10312 5333 12746 5343
rect 12760 5333 13706 5343
rect 13720 5333 18194 5343
rect 3760 5309 4274 5319
rect 4288 5309 4466 5319
rect 4480 5309 5786 5319
rect 5800 5309 6050 5319
rect 6064 5309 12026 5319
rect 12040 5309 14978 5319
rect 14992 5309 17078 5319
rect 17728 5309 17858 5319
rect 19888 5309 19994 5319
rect 3712 5285 25826 5295
rect 3592 5261 7226 5271
rect 7240 5261 9938 5271
rect 9952 5261 12098 5271
rect 12112 5261 16898 5271
rect 16912 5261 21194 5271
rect 3544 5237 7178 5247
rect 7192 5237 11114 5247
rect 11128 5237 12074 5247
rect 12088 5237 16874 5247
rect 16888 5237 26066 5247
rect 3496 5213 10610 5223
rect 10624 5213 23762 5223
rect 3376 5189 6962 5199
rect 6976 5189 13370 5199
rect 13384 5189 16202 5199
rect 16216 5189 17690 5199
rect 17704 5189 19634 5199
rect 19768 5189 19898 5199
rect 3328 5165 12314 5175
rect 12376 5165 17042 5175
rect 17056 5165 22706 5175
rect 3304 5141 18818 5151
rect 18832 5141 19946 5151
rect 19960 5141 21146 5151
rect 3256 5117 21602 5127
rect 3208 5093 17930 5103
rect 19120 5093 24914 5103
rect 3136 5069 5234 5079
rect 5296 5069 23090 5079
rect 3088 5045 20786 5055
rect 3040 5021 7538 5031
rect 7624 5021 8066 5031
rect 8080 5021 20162 5031
rect 3016 4997 10370 5007
rect 10384 4997 19874 5007
rect 20368 4997 21266 5007
rect 2920 4973 3410 4983
rect 3424 4973 4850 4983
rect 4864 4973 5402 4983
rect 5416 4973 10418 4983
rect 10432 4973 13874 4983
rect 13888 4973 23690 4983
rect 2896 4949 3770 4959
rect 3784 4949 4250 4959
rect 4264 4949 7610 4959
rect 7624 4949 10946 4959
rect 10960 4949 12554 4959
rect 12568 4949 23378 4959
rect 2872 4925 3866 4935
rect 3880 4925 4826 4935
rect 4840 4925 7850 4935
rect 7864 4925 13466 4935
rect 13480 4925 15386 4935
rect 15400 4925 15938 4935
rect 15952 4925 16826 4935
rect 16840 4925 16970 4935
rect 16984 4925 19298 4935
rect 19312 4925 19754 4935
rect 19768 4925 20834 4935
rect 20848 4925 21458 4935
rect 21472 4925 26930 4935
rect 2824 4901 16346 4911
rect 16480 4901 23810 4911
rect 2776 4877 7442 4887
rect 7456 4877 13106 4887
rect 13120 4877 17234 4887
rect 17248 4877 17882 4887
rect 17896 4877 22442 4887
rect 2704 4853 3314 4863
rect 3328 4853 7994 4863
rect 8008 4853 8138 4863
rect 8152 4853 13178 4863
rect 13192 4853 17354 4863
rect 17368 4853 23570 4863
rect 2680 4829 4634 4839
rect 4648 4829 5834 4839
rect 5848 4829 7058 4839
rect 7072 4829 9938 4839
rect 9952 4829 10850 4839
rect 10864 4829 17714 4839
rect 17728 4829 19250 4839
rect 20224 4829 20798 4839
rect 23680 4829 23738 4839
rect 2632 4805 23666 4815
rect 2584 4781 4418 4791
rect 4432 4781 14642 4791
rect 14848 4781 25130 4791
rect 2536 4757 4178 4767
rect 4192 4757 12650 4767
rect 12664 4757 16346 4767
rect 16408 4757 17162 4767
rect 18712 4757 19370 4767
rect 20032 4757 20522 4767
rect 20704 4757 20954 4767
rect 2512 4733 8954 4743
rect 8968 4733 9314 4743
rect 9328 4733 12866 4743
rect 12880 4733 14354 4743
rect 14368 4733 20114 4743
rect 20128 4733 22418 4743
rect 22432 4733 25778 4743
rect 2488 4709 7658 4719
rect 7672 4709 8930 4719
rect 8944 4709 13490 4719
rect 13504 4709 21338 4719
rect 21352 4709 22298 4719
rect 22408 4709 22454 4719
rect 23128 4709 23246 4719
rect 24328 4709 24482 4719
rect 2464 4685 3146 4695
rect 3160 4685 4730 4695
rect 4744 4685 8090 4695
rect 8104 4685 9506 4695
rect 9520 4685 11522 4695
rect 11536 4685 20066 4695
rect 20080 4685 22394 4695
rect 22408 4685 25106 4695
rect 25120 4685 25178 4695
rect 2344 4661 8114 4671
rect 8176 4661 13226 4671
rect 13432 4661 20702 4671
rect 23056 4661 23882 4671
rect 24136 4661 25442 4671
rect 2248 4637 4586 4647
rect 4600 4637 16706 4647
rect 16912 4637 17078 4647
rect 18256 4637 25730 4647
rect 2224 4613 7466 4623
rect 7480 4613 20018 4623
rect 20032 4613 25394 4623
rect 2176 4589 3170 4599
rect 3232 4589 9794 4599
rect 9976 4589 19382 4599
rect 19792 4589 20906 4599
rect 22504 4589 22730 4599
rect 22864 4589 23618 4599
rect 24016 4589 24290 4599
rect 24448 4589 24602 4599
rect 2128 4565 6146 4575
rect 6160 4565 7202 4575
rect 7216 4565 20594 4575
rect 20608 4565 24986 4575
rect 26176 4565 26450 4575
rect 2056 4541 5354 4551
rect 5368 4541 6698 4551
rect 6712 4541 11930 4551
rect 11944 4541 17330 4551
rect 17344 4541 26858 4551
rect 1960 4517 10586 4527
rect 10600 4517 24434 4527
rect 25840 4517 25874 4527
rect 26104 4517 26534 4527
rect 1912 4493 25538 4503
rect 26536 4493 27002 4503
rect 1840 4469 3962 4479
rect 3976 4469 5714 4479
rect 5728 4469 6482 4479
rect 6496 4469 6506 4479
rect 6520 4469 18122 4479
rect 18136 4469 20978 4479
rect 21064 4469 21314 4479
rect 21616 4469 21626 4479
rect 21736 4469 21914 4479
rect 21928 4469 24506 4479
rect 1816 4445 3650 4455
rect 3664 4445 9962 4455
rect 9976 4445 12242 4455
rect 12256 4445 12794 4455
rect 12808 4445 19226 4455
rect 19696 4445 24890 4455
rect 1792 4421 3674 4431
rect 3688 4421 19202 4431
rect 19216 4421 20354 4431
rect 20368 4421 24050 4431
rect 24136 4421 26642 4431
rect 1672 4397 1994 4407
rect 2008 4397 6170 4407
rect 6184 4397 8882 4407
rect 8896 4397 9890 4407
rect 9904 4397 11282 4407
rect 11296 4397 12290 4407
rect 12304 4397 13082 4407
rect 13096 4397 14114 4407
rect 14128 4397 18266 4407
rect 18280 4397 21002 4407
rect 21016 4397 23018 4407
rect 23032 4397 23906 4407
rect 23920 4397 24002 4407
rect 24016 4397 26498 4407
rect 1648 4373 6050 4383
rect 6064 4373 14882 4383
rect 15688 4373 22682 4383
rect 22768 4373 23150 4383
rect 23776 4373 23942 4383
rect 24040 4373 25610 4383
rect 26512 4373 26906 4383
rect 1624 4349 1922 4359
rect 1936 4349 3458 4359
rect 3472 4349 6074 4359
rect 6088 4349 7106 4359
rect 7120 4349 9506 4359
rect 9520 4349 13970 4359
rect 13984 4349 14234 4359
rect 14248 4349 16658 4359
rect 16672 4349 23282 4359
rect 23296 4349 24578 4359
rect 84 4325 3770 4335
rect 3784 4325 8282 4335
rect 8296 4325 9530 4335
rect 9544 4325 15986 4335
rect 16312 4325 21170 4335
rect 21184 4325 24218 4335
rect 24232 4325 24602 4335
rect 84 4301 7562 4311
rect 7696 4301 16778 4311
rect 16792 4301 26714 4311
rect 1624 4277 10994 4287
rect 11008 4277 25754 4287
rect 1648 4253 2930 4263
rect 2992 4253 6650 4263
rect 6664 4253 7922 4263
rect 7936 4253 14330 4263
rect 14344 4253 16730 4263
rect 16744 4253 20090 4263
rect 20416 4253 20546 4263
rect 20680 4253 20930 4263
rect 21352 4253 21410 4263
rect 21784 4253 22154 4263
rect 22312 4253 22538 4263
rect 22864 4253 26258 4263
rect 26272 4253 26402 4263
rect 1696 4229 4514 4239
rect 4576 4229 21482 4239
rect 22000 4229 22454 4239
rect 22960 4229 25082 4239
rect 1744 4205 13034 4215
rect 13096 4205 13106 4215
rect 13504 4205 13562 4215
rect 13792 4205 20378 4215
rect 21496 4205 21530 4215
rect 22096 4205 26186 4215
rect 1864 4181 12482 4191
rect 12568 4181 17858 4191
rect 18136 4181 18170 4191
rect 19120 4181 19154 4191
rect 19216 4181 19802 4191
rect 19960 4181 20294 4191
rect 23080 4181 23402 4191
rect 24280 4181 24794 4191
rect 2152 4157 7250 4167
rect 7264 4157 13274 4167
rect 13288 4157 18242 4167
rect 18256 4157 18962 4167
rect 18976 4157 20450 4167
rect 20464 4157 20762 4167
rect 20776 4157 21218 4167
rect 21232 4157 22154 4167
rect 22168 4157 22274 4167
rect 22288 4157 23210 4167
rect 23224 4157 26954 4167
rect 2200 4133 2594 4143
rect 2608 4133 6242 4143
rect 6256 4133 6602 4143
rect 6616 4133 6986 4143
rect 7000 4133 8618 4143
rect 8632 4133 10922 4143
rect 10936 4133 12602 4143
rect 12616 4133 14018 4143
rect 14032 4133 23786 4143
rect 23800 4133 23978 4143
rect 2344 4109 2618 4119
rect 2632 4109 5858 4119
rect 5872 4109 12722 4119
rect 12736 4109 14114 4119
rect 14128 4109 14210 4119
rect 14224 4109 15890 4119
rect 15904 4109 16418 4119
rect 16432 4109 19058 4119
rect 19072 4109 23114 4119
rect 23416 4109 24842 4119
rect 2368 4085 8306 4095
rect 8368 4085 11354 4095
rect 11368 4085 11954 4095
rect 11968 4085 24314 4095
rect 2368 4061 6890 4071
rect 6904 4061 7946 4071
rect 7960 4061 8570 4071
rect 8584 4061 13634 4071
rect 13648 4061 15842 4071
rect 15856 4061 24554 4071
rect 2392 4037 22442 4047
rect 23800 4037 24146 4047
rect 2392 4013 20186 4023
rect 20200 4013 20210 4023
rect 20464 4013 20702 4023
rect 2416 3989 2738 3999
rect 2800 3989 26570 3999
rect 2440 3965 5930 3975
rect 5944 3965 7010 3975
rect 7024 3965 11234 3975
rect 11248 3965 12050 3975
rect 12064 3965 13586 3975
rect 13600 3965 14954 3975
rect 14968 3965 15914 3975
rect 15928 3965 17162 3975
rect 17176 3965 17810 3975
rect 17824 3965 18098 3975
rect 18112 3965 19706 3975
rect 19720 3965 26354 3975
rect 2464 3941 4034 3951
rect 4048 3941 20282 3951
rect 20296 3941 26474 3951
rect 2488 3917 4370 3927
rect 4384 3917 11162 3927
rect 11176 3917 14090 3927
rect 14104 3917 16802 3927
rect 16816 3917 20042 3927
rect 20056 3917 21122 3927
rect 21136 3917 23330 3927
rect 26488 3917 26774 3927
rect 2560 3893 3434 3903
rect 3448 3893 3746 3903
rect 3760 3893 3986 3903
rect 4000 3893 7130 3903
rect 7144 3893 13730 3903
rect 13744 3893 15002 3903
rect 15016 3893 24242 3903
rect 2584 3869 19010 3879
rect 19024 3869 19610 3879
rect 19624 3869 22898 3879
rect 22912 3869 26594 3879
rect 2728 3845 10490 3855
rect 10552 3845 16058 3855
rect 16384 3845 27074 3855
rect 3112 3821 21866 3831
rect 3112 3797 5066 3807
rect 5080 3797 5138 3807
rect 5152 3797 8714 3807
rect 8728 3797 9338 3807
rect 9352 3797 16538 3807
rect 16552 3797 19850 3807
rect 19864 3797 21242 3807
rect 21256 3797 24074 3807
rect 24088 3797 24530 3807
rect 24544 3797 25946 3807
rect 3304 3773 6146 3783
rect 6160 3773 8186 3783
rect 8200 3773 8618 3783
rect 8632 3773 8858 3783
rect 8872 3773 9002 3783
rect 9016 3773 9098 3783
rect 9112 3773 10514 3783
rect 10528 3773 12386 3783
rect 12400 3773 18218 3783
rect 18232 3773 19898 3783
rect 20128 3773 21074 3783
rect 3352 3749 6434 3759
rect 6448 3749 15866 3759
rect 15880 3749 20858 3759
rect 3400 3725 6098 3735
rect 6112 3725 22562 3735
rect 3448 3701 10826 3711
rect 10840 3701 13898 3711
rect 13912 3701 20738 3711
rect 20872 3701 26882 3711
rect 3520 3677 4274 3687
rect 4288 3677 9746 3687
rect 9760 3677 12770 3687
rect 12784 3677 22706 3687
rect 3616 3653 26162 3663
rect 3616 3629 9146 3639
rect 9256 3629 27050 3639
rect 3736 3605 5666 3615
rect 5680 3605 7634 3615
rect 7648 3605 12962 3615
rect 12976 3605 13850 3615
rect 13864 3605 20498 3615
rect 20512 3605 24338 3615
rect 3808 3581 5570 3591
rect 5632 3581 20234 3591
rect 22576 3581 22826 3591
rect 3856 3557 5258 3567
rect 5272 3557 6866 3567
rect 6880 3557 12530 3567
rect 12544 3557 19346 3567
rect 19360 3557 19994 3567
rect 3952 3533 11186 3543
rect 11320 3533 19442 3543
rect 4000 3509 19322 3519
rect 4168 3485 6674 3495
rect 6688 3485 13154 3495
rect 13168 3485 21098 3495
rect 21112 3485 23186 3495
rect 23200 3485 26834 3495
rect 4192 3461 7298 3471
rect 7312 3461 24626 3471
rect 4312 3437 19562 3447
rect 4504 3413 5090 3423
rect 5176 3413 10850 3423
rect 10864 3413 18314 3423
rect 19336 3413 19382 3423
rect 4600 3389 9194 3399
rect 9304 3389 16034 3399
rect 16576 3389 25586 3399
rect 4720 3365 8738 3375
rect 8752 3365 23546 3375
rect 23560 3365 25490 3375
rect 4888 3341 10730 3351
rect 10912 3341 16610 3351
rect 16768 3341 23306 3351
rect 5008 3317 21458 3327
rect 5200 3293 11018 3303
rect 11080 3293 12074 3303
rect 12088 3293 22490 3303
rect 5368 3269 19922 3279
rect 19936 3269 25010 3279
rect 5536 3245 8090 3255
rect 8104 3245 8810 3255
rect 8824 3245 10202 3255
rect 10216 3245 14042 3255
rect 14056 3245 17018 3255
rect 17032 3245 20234 3255
rect 20248 3245 23138 3255
rect 23152 3245 25850 3255
rect 5560 3221 9650 3231
rect 9784 3221 9818 3231
rect 10072 3221 24938 3231
rect 5560 3197 22994 3207
rect 5608 3173 11882 3183
rect 11896 3173 13514 3183
rect 13528 3173 19586 3183
rect 19600 3173 21434 3183
rect 5632 3149 6770 3159
rect 6784 3149 8234 3159
rect 8248 3149 9770 3159
rect 9784 3149 11498 3159
rect 11512 3149 12506 3159
rect 12520 3149 13586 3159
rect 13600 3149 19490 3159
rect 19504 3149 25082 3159
rect 25096 3149 26450 3159
rect 5704 3125 10178 3135
rect 10240 3125 19514 3135
rect 5776 3101 17402 3111
rect 17512 3101 20882 3111
rect 5872 3077 10706 3087
rect 11008 3077 11330 3087
rect 11632 3077 23930 3087
rect 5920 3053 7034 3063
rect 7048 3053 8882 3063
rect 8896 3053 10034 3063
rect 10096 3053 24458 3063
rect 6016 3029 7034 3039
rect 7048 3029 11138 3039
rect 11224 3029 26666 3039
rect 6208 3005 6362 3015
rect 6448 3005 14258 3015
rect 14464 3005 25994 3015
rect 6208 2981 22874 2991
rect 6280 2957 12146 2967
rect 12472 2957 24722 2967
rect 6304 2933 9026 2943
rect 9088 2933 9602 2943
rect 9616 2933 13346 2943
rect 13528 2933 22586 2943
rect 6352 2909 17066 2919
rect 17200 2909 25706 2919
rect 6400 2885 23450 2895
rect 6496 2861 8978 2871
rect 8992 2861 11978 2871
rect 11992 2861 15818 2871
rect 15832 2861 20738 2871
rect 6760 2837 9434 2847
rect 9544 2837 10562 2847
rect 11104 2837 21242 2847
rect 21256 2837 22370 2847
rect 22384 2837 26042 2847
rect 6784 2813 6794 2823
rect 6856 2813 22610 2823
rect 22624 2813 23354 2823
rect 6808 2789 21386 2799
rect 22624 2789 26114 2799
rect 26128 2789 26306 2799
rect 6880 2765 20522 2775
rect 21400 2765 21506 2775
rect 6952 2741 26186 2751
rect 6952 2717 25274 2727
rect 7096 2693 7970 2703
rect 7984 2693 8642 2703
rect 8656 2693 9866 2703
rect 9880 2693 10178 2703
rect 10192 2693 11954 2703
rect 11968 2693 16010 2703
rect 16024 2693 16202 2703
rect 16216 2693 17762 2703
rect 17776 2693 22226 2703
rect 22240 2693 25514 2703
rect 7144 2669 7826 2679
rect 7840 2669 11762 2679
rect 11776 2669 13250 2679
rect 13264 2669 16994 2679
rect 17752 2669 20702 2679
rect 20716 2669 24098 2679
rect 7168 2645 17642 2655
rect 17896 2645 17906 2655
rect 7216 2621 7226 2631
rect 7288 2621 9050 2631
rect 9112 2621 14810 2631
rect 14824 2621 17474 2631
rect 7288 2597 8018 2607
rect 8032 2597 12266 2607
rect 12280 2597 14066 2607
rect 14080 2597 17378 2607
rect 17392 2597 22970 2607
rect 7360 2573 11738 2583
rect 11800 2573 22658 2583
rect 7408 2549 14138 2559
rect 14152 2549 23690 2559
rect 7432 2525 9794 2535
rect 9808 2525 24194 2535
rect 7528 2501 19274 2511
rect 7552 2477 7586 2487
rect 7744 2477 17522 2487
rect 7744 2453 9698 2463
rect 10144 2453 14162 2463
rect 14176 2453 18554 2463
rect 18568 2453 19970 2463
rect 19984 2453 20798 2463
rect 7888 2429 7898 2439
rect 7984 2429 8810 2439
rect 8824 2429 14282 2439
rect 14296 2429 21002 2439
rect 21016 2429 23738 2439
rect 23752 2429 23882 2439
rect 8056 2405 11258 2415
rect 11272 2405 17138 2415
rect 19984 2405 26282 2415
rect 26296 2405 26378 2415
rect 8296 2381 8546 2391
rect 8560 2381 12410 2391
rect 12424 2381 22034 2391
rect 8392 2357 21962 2367
rect 8416 2333 8426 2343
rect 8512 2333 9746 2343
rect 9760 2333 10418 2343
rect 10432 2333 10442 2343
rect 10456 2333 21266 2343
rect 21280 2333 21362 2343
rect 21376 2333 22130 2343
rect 22144 2333 23474 2343
rect 23488 2333 24410 2343
rect 24424 2333 24482 2343
rect 8512 2309 13538 2319
rect 13552 2309 20258 2319
rect 20272 2309 23042 2319
rect 23056 2309 23546 2319
rect 8536 2285 15698 2295
rect 15880 2285 19466 2295
rect 21976 2285 22010 2295
rect 8680 2261 17450 2271
rect 8848 2237 8906 2247
rect 8992 2237 23246 2247
rect 9160 2213 9362 2223
rect 9424 2213 13418 2223
rect 13432 2213 23018 2223
rect 9208 2189 9266 2199
rect 9328 2189 16490 2199
rect 16504 2189 23282 2199
rect 9592 2165 20474 2175
rect 9592 2141 25898 2151
rect 9640 2117 19490 2127
rect 9712 2093 9818 2103
rect 10264 2093 15962 2103
rect 16624 2093 26690 2103
rect 10600 2069 10610 2079
rect 11176 2069 11354 2079
rect 11656 2069 13682 2079
rect 13816 2069 16082 2079
rect 16096 2069 24386 2079
rect 12520 2045 22730 2055
rect 12616 2021 12698 2031
rect 12832 2021 17570 2031
rect 17584 2021 20570 2031
rect 20584 2021 20618 2031
rect 12928 1997 14930 2007
rect 14944 1997 26618 2007
rect 13120 1973 27026 1983
rect 13288 1949 13394 1959
rect 13840 1949 19058 1959
rect 19072 1949 19418 1959
rect 20632 1949 20702 1959
rect 13888 1925 13922 1935
rect 14080 1925 14186 1935
rect 14680 1925 14690 1935
rect 14920 1925 27445 1935
rect 13936 1901 15626 1911
rect 15640 1901 15914 1911
rect 15928 1901 22634 1911
rect 22648 1901 24290 1911
rect 24304 1901 24338 1911
rect 24352 1901 26258 1911
rect 14152 1877 20786 1887
rect 20800 1877 25970 1887
rect 27088 1877 27445 1887
rect 16096 1853 17978 1863
rect 17992 1853 23834 1863
rect 25984 1853 26018 1863
rect 27064 1853 27445 1863
rect 16792 1829 16922 1839
rect 17008 1829 18362 1839
rect 27040 1829 27445 1839
rect 26595 1800 27050 1810
rect 26595 1777 27050 1787
rect 27046 1748 27050 1764
rect 26595 1739 27050 1748
rect 26654 1119 26670 1329
rect 26780 1119 26796 1329
rect 26906 1119 26922 1329
rect 26595 1110 27050 1119
rect 27041 1094 27050 1110
rect 26595 1071 27050 1081
rect 26595 1048 27050 1058
rect 26595 1025 27050 1035
rect 18088 996 18290 1006
rect 18064 972 25274 982
rect 17584 948 18146 958
rect 11056 924 18962 934
rect 10960 900 18098 910
rect 19024 900 26450 910
rect 10840 876 16226 886
rect 16480 876 21746 886
rect 10648 852 15098 862
rect 15112 852 15962 862
rect 16024 852 19394 862
rect 9424 828 9890 838
rect 10120 828 21938 838
rect 9352 804 13562 814
rect 14440 804 24458 814
rect 9064 780 19346 790
rect 8776 756 12842 766
rect 13000 756 13610 766
rect 13960 756 19538 766
rect 23008 756 26282 766
rect 8440 732 26114 742
rect 8272 708 13322 718
rect 13744 708 24098 718
rect 7948 684 9698 694
rect 9880 684 21506 694
rect 21592 684 24554 694
rect 7768 660 26378 670
rect 7576 636 11258 646
rect 12376 636 14474 646
rect 14536 636 19658 646
rect 19672 636 24362 646
rect 7240 612 19178 622
rect 19480 612 20066 622
rect 21424 612 25418 622
rect 6592 588 19778 598
rect 21376 588 23498 598
rect 6400 564 13130 574
rect 13408 564 13682 574
rect 13696 564 14570 574
rect 14872 564 19586 574
rect 19744 564 20522 574
rect 20584 564 26594 574
rect 6328 540 26138 550
rect 6256 516 16682 526
rect 17272 516 27445 526
rect 5968 492 24194 502
rect 5752 468 20930 478
rect 5656 444 21314 454
rect 5512 420 22658 430
rect 4792 396 6626 406
rect 6832 396 24674 406
rect 4768 372 14378 382
rect 14920 372 21698 382
rect 4552 348 12410 358
rect 12544 348 14690 358
rect 15160 348 17810 358
rect 17824 348 24242 358
rect 4384 324 10322 334
rect 10336 324 10706 334
rect 10768 324 24506 334
rect 4336 300 26018 310
rect 3904 276 4802 286
rect 4960 276 26042 286
rect 3688 252 19418 262
rect 3640 228 12314 238
rect 14320 228 22730 238
rect 3568 204 6410 214
rect 6544 204 22058 214
rect 22072 204 23234 214
rect 2512 180 20882 190
rect 1792 156 4826 166
rect 5320 156 22826 166
rect 1672 132 9482 142
rect 10552 132 12266 142
rect 15280 132 18818 142
rect 84 108 21626 118
rect 84 84 17930 94
rect 17992 84 18410 94
rect 3544 60 20690 70
rect 26584 60 27445 70
rect 4312 36 14330 46
rect 16144 36 16322 46
rect 17296 36 25994 46
rect 26584 36 27445 46
rect 17896 12 26570 22
rect 26608 12 27445 22
<< m2contact >>
rect 15698 8420 15712 8434
rect 16862 8420 16876 8434
rect 20282 8420 20296 8434
rect 13802 8396 13816 8410
rect 14666 8396 14680 8410
rect 22766 8396 22780 8410
rect 2282 8372 2296 8386
rect 17726 8372 17740 8386
rect 70 8348 84 8362
rect 23138 8348 23152 8362
rect 70 8324 84 8338
rect 1730 8324 1744 8338
rect 1994 8324 2008 8338
rect 2450 8324 2464 8338
rect 3530 8324 3544 8338
rect 7562 8324 7576 8338
rect 9230 8324 9244 8338
rect 19154 8324 19168 8338
rect 19382 8324 19396 8338
rect 20546 8324 20560 8338
rect 21902 8324 21916 8338
rect 22154 8324 22168 8338
rect 24422 8324 24436 8338
rect 25010 8324 25024 8338
rect 2138 8300 2152 8314
rect 3554 8300 3568 8314
rect 22010 8300 22024 8314
rect 25286 8300 25300 8314
rect 2414 8276 2428 8290
rect 7970 8276 7984 8290
rect 8330 8276 8344 8290
rect 9266 8276 9280 8290
rect 9458 8276 9472 8290
rect 12674 8276 12688 8290
rect 12866 8276 12880 8290
rect 24446 8276 24460 8290
rect 4118 8252 4132 8266
rect 7946 8252 7960 8266
rect 10754 8252 10768 8266
rect 26126 8252 26140 8266
rect 27026 8252 27040 8266
rect 27050 8252 27064 8266
rect 4202 8228 4216 8242
rect 27074 8228 27088 8242
rect 4970 8204 4984 8218
rect 8810 8204 8824 8218
rect 10934 8204 10948 8218
rect 25778 8204 25792 8218
rect 5822 8180 5836 8194
rect 6074 8180 6088 8194
rect 6266 8180 6280 8194
rect 7526 8180 7540 8194
rect 9938 8180 9952 8194
rect 11450 8180 11464 8194
rect 19406 8180 19420 8194
rect 20690 8180 20704 8194
rect 22394 8180 22408 8194
rect 24794 8180 24808 8194
rect 27122 8180 27136 8194
rect 11786 8156 11800 8170
rect 20930 8156 20944 8170
rect 27098 8156 27112 8170
rect 27445 8156 27459 8170
rect 12638 8132 12652 8146
rect 24146 8132 24160 8146
rect 27074 8132 27088 8146
rect 27445 8132 27459 8146
rect 15182 8108 15196 8122
rect 23402 8108 23416 8122
rect 27050 8108 27064 8122
rect 27445 8108 27459 8122
rect 17702 8084 17716 8098
rect 18650 8084 18664 8098
rect 27445 8084 27459 8098
rect 19418 8060 19432 8074
rect 27098 8060 27112 8074
rect 27122 8060 27136 8074
rect 27445 8060 27459 8074
rect 15818 7227 15832 7241
rect 15962 7227 15976 7241
rect 14882 7203 14896 7217
rect 14930 7203 14944 7217
rect 15026 7203 15040 7217
rect 27002 7203 27016 7217
rect 14138 7179 14152 7193
rect 18170 7179 18184 7193
rect 13226 7155 13240 7169
rect 13346 7155 13360 7169
rect 13898 7155 13912 7169
rect 14138 7155 14152 7169
rect 14618 7155 14632 7169
rect 20294 7155 20308 7169
rect 13178 7131 13192 7145
rect 13250 7131 13264 7145
rect 13802 7131 13816 7145
rect 23594 7131 23608 7145
rect 13106 7107 13120 7121
rect 24146 7107 24160 7121
rect 13058 7083 13072 7097
rect 22250 7083 22264 7097
rect 13010 7059 13024 7073
rect 24674 7059 24688 7073
rect 12962 7035 12976 7049
rect 22346 7035 22360 7049
rect 12698 7011 12712 7025
rect 14186 7011 14200 7025
rect 26234 7011 26248 7025
rect 12482 6987 12496 7001
rect 12530 6987 12544 7001
rect 12650 6987 12664 7001
rect 21506 6987 21520 7001
rect 12026 6963 12040 6977
rect 12146 6963 12160 6977
rect 12194 6963 12208 6977
rect 23978 6963 23992 6977
rect 11690 6939 11704 6953
rect 18194 6939 18208 6953
rect 11354 6915 11368 6929
rect 26762 6915 26776 6929
rect 10514 6891 10528 6905
rect 21314 6891 21328 6905
rect 10442 6867 10456 6881
rect 12938 6867 12952 6881
rect 12986 6867 13000 6881
rect 16922 6867 16936 6881
rect 10370 6843 10384 6857
rect 10442 6843 10456 6857
rect 10490 6843 10504 6857
rect 10562 6843 10576 6857
rect 10634 6843 10648 6857
rect 16442 6843 16456 6857
rect 10298 6819 10312 6833
rect 11402 6819 11416 6833
rect 11594 6819 11608 6833
rect 18026 6819 18040 6833
rect 9650 6795 9664 6809
rect 17834 6795 17848 6809
rect 9434 6771 9448 6785
rect 15050 6771 15064 6785
rect 15770 6771 15784 6785
rect 23714 6771 23728 6785
rect 9362 6747 9376 6761
rect 19826 6747 19840 6761
rect 22778 6747 22792 6761
rect 9218 6723 9232 6737
rect 21290 6723 21304 6737
rect 9026 6699 9040 6713
rect 9050 6699 9064 6713
rect 9170 6699 9184 6713
rect 18770 6699 18784 6713
rect 8954 6675 8968 6689
rect 17042 6675 17056 6689
rect 8906 6651 8920 6665
rect 10802 6651 10816 6665
rect 10874 6651 10888 6665
rect 11042 6651 11056 6665
rect 11090 6651 11104 6665
rect 23450 6651 23464 6665
rect 8762 6627 8776 6641
rect 13946 6627 13960 6641
rect 13994 6627 14008 6641
rect 15986 6627 16000 6641
rect 8570 6603 8584 6617
rect 26774 6603 26788 6617
rect 8450 6579 8464 6593
rect 13994 6579 14008 6593
rect 23186 6579 23200 6593
rect 8258 6555 8272 6569
rect 16130 6555 16144 6569
rect 16370 6555 16384 6569
rect 23150 6555 23164 6569
rect 8210 6531 8224 6545
rect 23858 6531 23872 6545
rect 7802 6507 7816 6521
rect 18602 6507 18616 6521
rect 7778 6483 7792 6497
rect 18722 6483 18736 6497
rect 20330 6483 20344 6497
rect 23714 6483 23728 6497
rect 7754 6459 7768 6473
rect 8210 6459 8224 6473
rect 8714 6459 8728 6473
rect 12626 6459 12640 6473
rect 13298 6459 13312 6473
rect 19826 6459 19840 6473
rect 22322 6459 22336 6473
rect 25202 6459 25216 6473
rect 25874 6459 25888 6473
rect 7514 6435 7528 6449
rect 23498 6435 23512 6449
rect 7418 6411 7432 6425
rect 15938 6411 15952 6425
rect 16250 6411 16264 6425
rect 20330 6411 20344 6425
rect 7370 6387 7384 6401
rect 26522 6387 26536 6401
rect 7298 6363 7312 6377
rect 13298 6363 13312 6377
rect 13658 6363 13672 6377
rect 13682 6363 13696 6377
rect 13754 6363 13768 6377
rect 15746 6363 15760 6377
rect 15794 6363 15808 6377
rect 20138 6363 20152 6377
rect 22010 6363 22024 6377
rect 7178 6339 7192 6353
rect 12122 6339 12136 6353
rect 13394 6339 13408 6353
rect 26978 6339 26992 6353
rect 7082 6315 7096 6329
rect 21098 6315 21112 6329
rect 6986 6291 7000 6305
rect 8474 6291 8488 6305
rect 8522 6291 8536 6305
rect 10394 6291 10408 6305
rect 10922 6291 10936 6305
rect 12170 6291 12184 6305
rect 15122 6291 15136 6305
rect 21074 6291 21088 6305
rect 21818 6291 21832 6305
rect 6890 6267 6904 6281
rect 7490 6267 7504 6281
rect 21554 6267 21568 6281
rect 6722 6243 6736 6257
rect 7346 6243 7360 6257
rect 7394 6243 7408 6257
rect 25346 6243 25360 6257
rect 6698 6219 6712 6233
rect 21626 6219 21640 6233
rect 22202 6219 22216 6233
rect 22370 6219 22384 6233
rect 6674 6195 6688 6209
rect 11834 6195 11848 6209
rect 22754 6195 22768 6209
rect 25226 6195 25240 6209
rect 26426 6195 26440 6209
rect 26690 6195 26704 6209
rect 6602 6171 6616 6185
rect 26426 6171 26440 6185
rect 6578 6147 6592 6161
rect 14738 6147 14752 6161
rect 26210 6147 26224 6161
rect 6554 6123 6568 6137
rect 9386 6123 9400 6137
rect 14690 6123 14704 6137
rect 22202 6123 22216 6137
rect 6362 6099 6376 6113
rect 14786 6099 14800 6113
rect 14858 6099 14872 6113
rect 25658 6099 25672 6113
rect 6266 6075 6280 6089
rect 8426 6075 8440 6089
rect 11978 6075 11992 6089
rect 12722 6075 12736 6089
rect 15578 6075 15592 6089
rect 16586 6075 16600 6089
rect 16682 6075 16696 6089
rect 19802 6075 19816 6089
rect 22802 6075 22816 6089
rect 23306 6075 23320 6089
rect 6170 6051 6184 6065
rect 14666 6051 14680 6065
rect 22802 6051 22816 6065
rect 6002 6027 6016 6041
rect 24866 6027 24880 6041
rect 5954 6003 5968 6017
rect 13706 6003 13720 6017
rect 22826 6003 22840 6017
rect 5906 5979 5920 5993
rect 11666 5979 11680 5993
rect 11786 5979 11800 5993
rect 26810 5979 26824 5993
rect 5882 5955 5896 5969
rect 23930 5955 23944 5969
rect 5810 5931 5824 5945
rect 19082 5931 19096 5945
rect 25226 5931 25240 5945
rect 5786 5907 5800 5921
rect 18146 5907 18160 5921
rect 18434 5907 18448 5921
rect 21530 5907 21544 5921
rect 23906 5907 23920 5921
rect 5714 5883 5728 5897
rect 21410 5883 21424 5897
rect 5690 5859 5704 5873
rect 9218 5859 9232 5873
rect 11330 5859 11344 5873
rect 11546 5859 11560 5873
rect 13010 5859 13024 5873
rect 13370 5859 13384 5873
rect 26570 5859 26584 5873
rect 5498 5835 5512 5849
rect 9362 5835 9376 5849
rect 26906 5835 26920 5849
rect 5474 5811 5488 5825
rect 9842 5811 9856 5825
rect 15434 5811 15448 5825
rect 18938 5811 18952 5825
rect 18986 5811 19000 5825
rect 20426 5811 20440 5825
rect 23942 5811 23956 5825
rect 26330 5811 26344 5825
rect 26534 5811 26548 5825
rect 5450 5787 5464 5801
rect 13322 5787 13336 5801
rect 13610 5787 13624 5801
rect 18866 5787 18880 5801
rect 19730 5787 19744 5801
rect 26330 5787 26344 5801
rect 5330 5763 5344 5777
rect 10970 5763 10984 5777
rect 13562 5763 13576 5777
rect 16442 5763 16456 5777
rect 16754 5763 16768 5777
rect 18482 5763 18496 5777
rect 21026 5763 21040 5777
rect 21842 5763 21856 5777
rect 26738 5763 26752 5777
rect 5042 5739 5056 5753
rect 19538 5739 19552 5753
rect 4922 5715 4936 5729
rect 22922 5715 22936 5729
rect 4778 5691 4792 5705
rect 5978 5691 5992 5705
rect 13922 5691 13936 5705
rect 23474 5691 23488 5705
rect 25034 5691 25048 5705
rect 26018 5691 26032 5705
rect 4706 5667 4720 5681
rect 7898 5667 7912 5681
rect 8690 5667 8704 5681
rect 19634 5667 19648 5681
rect 20138 5667 20152 5681
rect 22922 5667 22936 5681
rect 24362 5667 24376 5681
rect 25034 5667 25048 5681
rect 4634 5643 4648 5657
rect 15026 5643 15040 5657
rect 22514 5643 22528 5657
rect 25418 5643 25432 5657
rect 4538 5619 4552 5633
rect 8402 5619 8416 5633
rect 10274 5619 10288 5633
rect 16562 5619 16576 5633
rect 16826 5619 16840 5633
rect 21674 5619 21688 5633
rect 4490 5595 4504 5609
rect 4658 5595 4672 5609
rect 10058 5595 10072 5609
rect 13202 5595 13216 5609
rect 16634 5595 16648 5609
rect 16946 5595 16960 5609
rect 22322 5595 22336 5609
rect 4418 5571 4432 5585
rect 4946 5571 4960 5585
rect 16178 5571 16192 5585
rect 17594 5571 17608 5585
rect 4346 5547 4360 5561
rect 8906 5547 8920 5561
rect 9986 5547 10000 5561
rect 13658 5547 13672 5561
rect 16850 5547 16864 5561
rect 19250 5547 19264 5561
rect 21050 5547 21064 5561
rect 22250 5547 22264 5561
rect 4226 5523 4240 5537
rect 25298 5523 25312 5537
rect 4154 5499 4168 5513
rect 10010 5499 10024 5513
rect 12626 5499 12640 5513
rect 12674 5499 12688 5513
rect 27026 5499 27040 5513
rect 4130 5475 4144 5489
rect 17786 5475 17800 5489
rect 23234 5475 23248 5489
rect 24170 5475 24184 5489
rect 4106 5451 4120 5465
rect 7586 5451 7600 5465
rect 11426 5451 11440 5465
rect 12698 5451 12712 5465
rect 18626 5451 18640 5465
rect 19658 5451 19672 5465
rect 21122 5451 21136 5465
rect 4082 5427 4096 5441
rect 18578 5427 18592 5441
rect 4058 5403 4072 5417
rect 5810 5403 5824 5417
rect 8378 5403 8392 5417
rect 22538 5403 22552 5417
rect 3866 5379 3880 5393
rect 22346 5379 22360 5393
rect 3818 5355 3832 5369
rect 3890 5355 3904 5369
rect 3938 5355 3952 5369
rect 11378 5355 11392 5369
rect 16274 5355 16288 5369
rect 16322 5355 16336 5369
rect 20642 5355 20656 5369
rect 3794 5331 3808 5345
rect 4010 5331 4024 5345
rect 6122 5331 6136 5345
rect 7874 5331 7888 5345
rect 8834 5331 8848 5345
rect 10298 5331 10312 5345
rect 12746 5331 12760 5345
rect 13706 5331 13720 5345
rect 18194 5331 18208 5345
rect 3746 5307 3760 5321
rect 4274 5307 4288 5321
rect 4466 5307 4480 5321
rect 5786 5307 5800 5321
rect 6050 5307 6064 5321
rect 12026 5307 12040 5321
rect 14978 5307 14992 5321
rect 17078 5307 17092 5321
rect 17714 5307 17728 5321
rect 17858 5307 17872 5321
rect 19874 5307 19888 5321
rect 19994 5307 20008 5321
rect 3698 5283 3712 5297
rect 25826 5283 25840 5297
rect 3578 5259 3592 5273
rect 7226 5259 7240 5273
rect 9938 5259 9952 5273
rect 12098 5259 12112 5273
rect 16898 5259 16912 5273
rect 21194 5259 21208 5273
rect 3530 5235 3544 5249
rect 7178 5235 7192 5249
rect 11114 5235 11128 5249
rect 12074 5235 12088 5249
rect 16874 5235 16888 5249
rect 26066 5235 26080 5249
rect 3482 5211 3496 5225
rect 10610 5211 10624 5225
rect 23762 5211 23776 5225
rect 3362 5187 3376 5201
rect 6962 5187 6976 5201
rect 13370 5187 13384 5201
rect 16202 5187 16216 5201
rect 17690 5187 17704 5201
rect 19634 5187 19648 5201
rect 19754 5187 19768 5201
rect 19898 5187 19912 5201
rect 3314 5163 3328 5177
rect 12314 5163 12328 5177
rect 12362 5163 12376 5177
rect 17042 5163 17056 5177
rect 22706 5163 22720 5177
rect 3290 5139 3304 5153
rect 18818 5139 18832 5153
rect 19946 5139 19960 5153
rect 21146 5139 21160 5153
rect 3242 5115 3256 5129
rect 21602 5115 21616 5129
rect 3194 5091 3208 5105
rect 17930 5091 17944 5105
rect 19106 5091 19120 5105
rect 24914 5091 24928 5105
rect 3122 5067 3136 5081
rect 5234 5067 5248 5081
rect 5282 5067 5296 5081
rect 23090 5067 23104 5081
rect 3074 5043 3088 5057
rect 20786 5043 20800 5057
rect 3026 5019 3040 5033
rect 7538 5019 7552 5033
rect 7610 5019 7624 5033
rect 8066 5019 8080 5033
rect 20162 5019 20176 5033
rect 3002 4995 3016 5009
rect 10370 4995 10384 5009
rect 19874 4995 19888 5009
rect 20354 4995 20368 5009
rect 21266 4995 21280 5009
rect 2906 4971 2920 4985
rect 3410 4971 3424 4985
rect 4850 4971 4864 4985
rect 5402 4971 5416 4985
rect 10418 4971 10432 4985
rect 13874 4971 13888 4985
rect 23690 4971 23704 4985
rect 2882 4947 2896 4961
rect 3770 4947 3784 4961
rect 4250 4947 4264 4961
rect 7610 4947 7624 4961
rect 10946 4947 10960 4961
rect 12554 4947 12568 4961
rect 23378 4947 23392 4961
rect 2858 4923 2872 4937
rect 3866 4923 3880 4937
rect 4826 4923 4840 4937
rect 7850 4923 7864 4937
rect 13466 4923 13480 4937
rect 15386 4923 15400 4937
rect 15938 4923 15952 4937
rect 16826 4923 16840 4937
rect 16970 4923 16984 4937
rect 19298 4923 19312 4937
rect 19754 4923 19768 4937
rect 20834 4923 20848 4937
rect 21458 4923 21472 4937
rect 26930 4923 26944 4937
rect 2810 4899 2824 4913
rect 16346 4899 16360 4913
rect 16466 4899 16480 4913
rect 23810 4899 23824 4913
rect 2762 4875 2776 4889
rect 7442 4875 7456 4889
rect 13106 4875 13120 4889
rect 17234 4875 17248 4889
rect 17882 4875 17896 4889
rect 22442 4875 22456 4889
rect 2690 4851 2704 4865
rect 3314 4851 3328 4865
rect 7994 4851 8008 4865
rect 8138 4851 8152 4865
rect 13178 4851 13192 4865
rect 17354 4851 17368 4865
rect 23570 4851 23584 4865
rect 2666 4827 2680 4841
rect 4634 4827 4648 4841
rect 5834 4827 5848 4841
rect 7058 4827 7072 4841
rect 9938 4827 9952 4841
rect 10850 4827 10864 4841
rect 17714 4827 17728 4841
rect 19250 4827 19264 4841
rect 20210 4827 20224 4841
rect 20798 4827 20812 4841
rect 23666 4827 23680 4841
rect 23738 4827 23752 4841
rect 2618 4803 2632 4817
rect 23666 4803 23680 4817
rect 2570 4779 2584 4793
rect 4418 4779 4432 4793
rect 14642 4779 14656 4793
rect 14834 4779 14848 4793
rect 25130 4779 25144 4793
rect 2522 4755 2536 4769
rect 4178 4755 4192 4769
rect 12650 4755 12664 4769
rect 16346 4755 16360 4769
rect 16394 4755 16408 4769
rect 17162 4755 17176 4769
rect 18698 4755 18712 4769
rect 19370 4755 19384 4769
rect 20018 4755 20032 4769
rect 20522 4755 20536 4769
rect 20690 4755 20704 4769
rect 20954 4755 20968 4769
rect 2498 4731 2512 4745
rect 8954 4731 8968 4745
rect 9314 4731 9328 4745
rect 12866 4731 12880 4745
rect 14354 4731 14368 4745
rect 20114 4731 20128 4745
rect 22418 4731 22432 4745
rect 25778 4731 25792 4745
rect 2474 4707 2488 4721
rect 7658 4707 7672 4721
rect 8930 4707 8944 4721
rect 13490 4707 13504 4721
rect 21338 4707 21352 4721
rect 22298 4707 22312 4721
rect 22394 4707 22408 4721
rect 22454 4707 22468 4721
rect 23114 4707 23128 4721
rect 23246 4707 23260 4721
rect 24314 4707 24328 4721
rect 24482 4707 24496 4721
rect 2450 4683 2464 4697
rect 3146 4683 3160 4697
rect 4730 4683 4744 4697
rect 8090 4683 8104 4697
rect 9506 4683 9520 4697
rect 11522 4683 11536 4697
rect 20066 4683 20080 4697
rect 22394 4683 22408 4697
rect 25106 4683 25120 4697
rect 25178 4683 25192 4697
rect 2330 4659 2344 4673
rect 8114 4659 8128 4673
rect 8162 4659 8176 4673
rect 13226 4659 13240 4673
rect 13418 4659 13432 4673
rect 20702 4659 20716 4673
rect 23042 4659 23056 4673
rect 23882 4659 23896 4673
rect 24122 4659 24136 4673
rect 25442 4659 25456 4673
rect 2234 4635 2248 4649
rect 4586 4635 4600 4649
rect 16706 4635 16720 4649
rect 16898 4635 16912 4649
rect 17078 4635 17092 4649
rect 18242 4635 18256 4649
rect 25730 4635 25744 4649
rect 2210 4611 2224 4625
rect 7466 4611 7480 4625
rect 20018 4611 20032 4625
rect 25394 4611 25408 4625
rect 2162 4587 2176 4601
rect 3170 4587 3184 4601
rect 3218 4587 3232 4601
rect 9794 4587 9808 4601
rect 9962 4587 9976 4601
rect 19382 4587 19396 4601
rect 19778 4587 19792 4601
rect 20906 4587 20920 4601
rect 22490 4587 22504 4601
rect 22730 4587 22744 4601
rect 22850 4587 22864 4601
rect 23618 4587 23632 4601
rect 24002 4587 24016 4601
rect 24290 4587 24304 4601
rect 24434 4587 24448 4601
rect 24602 4587 24616 4601
rect 2114 4563 2128 4577
rect 6146 4563 6160 4577
rect 7202 4563 7216 4577
rect 20594 4563 20608 4577
rect 24986 4563 25000 4577
rect 26162 4563 26176 4577
rect 26450 4563 26464 4577
rect 2042 4539 2056 4553
rect 5354 4539 5368 4553
rect 6698 4539 6712 4553
rect 11930 4539 11944 4553
rect 17330 4539 17344 4553
rect 26858 4539 26872 4553
rect 1946 4515 1960 4529
rect 10586 4515 10600 4529
rect 24434 4515 24448 4529
rect 25826 4515 25840 4529
rect 25874 4515 25888 4529
rect 26090 4515 26104 4529
rect 26534 4515 26548 4529
rect 1898 4491 1912 4505
rect 25538 4491 25552 4505
rect 26522 4491 26536 4505
rect 27002 4491 27016 4505
rect 1826 4467 1840 4481
rect 3962 4467 3976 4481
rect 5714 4467 5728 4481
rect 6482 4467 6496 4481
rect 6506 4467 6520 4481
rect 18122 4467 18136 4481
rect 20978 4467 20992 4481
rect 21050 4467 21064 4481
rect 21314 4467 21328 4481
rect 21602 4467 21616 4481
rect 21626 4467 21640 4481
rect 21722 4467 21736 4481
rect 21914 4467 21928 4481
rect 24506 4467 24520 4481
rect 1802 4443 1816 4457
rect 3650 4443 3664 4457
rect 9962 4443 9976 4457
rect 12242 4443 12256 4457
rect 12794 4443 12808 4457
rect 19226 4443 19240 4457
rect 19682 4443 19696 4457
rect 24890 4443 24904 4457
rect 1778 4419 1792 4433
rect 3674 4419 3688 4433
rect 19202 4419 19216 4433
rect 20354 4419 20368 4433
rect 24050 4419 24064 4433
rect 24122 4419 24136 4433
rect 26642 4419 26656 4433
rect 1658 4395 1672 4409
rect 1994 4395 2008 4409
rect 6170 4395 6184 4409
rect 8882 4395 8896 4409
rect 9890 4395 9904 4409
rect 11282 4395 11296 4409
rect 12290 4395 12304 4409
rect 13082 4395 13096 4409
rect 14114 4395 14128 4409
rect 18266 4395 18280 4409
rect 21002 4395 21016 4409
rect 23018 4395 23032 4409
rect 23906 4395 23920 4409
rect 24002 4395 24016 4409
rect 26498 4395 26512 4409
rect 1634 4371 1648 4385
rect 6050 4371 6064 4385
rect 14882 4371 14896 4385
rect 15674 4371 15688 4385
rect 22682 4371 22696 4385
rect 22754 4371 22768 4385
rect 23150 4371 23164 4385
rect 23762 4371 23776 4385
rect 23942 4371 23956 4385
rect 24026 4371 24040 4385
rect 25610 4371 25624 4385
rect 26498 4371 26512 4385
rect 26906 4371 26920 4385
rect 1610 4347 1624 4361
rect 1922 4347 1936 4361
rect 3458 4347 3472 4361
rect 6074 4347 6088 4361
rect 7106 4347 7120 4361
rect 9506 4347 9520 4361
rect 13970 4347 13984 4361
rect 14234 4347 14248 4361
rect 16658 4347 16672 4361
rect 23282 4347 23296 4361
rect 24578 4347 24592 4361
rect 70 4323 84 4337
rect 3770 4323 3784 4337
rect 8282 4323 8296 4337
rect 9530 4323 9544 4337
rect 15986 4323 16000 4337
rect 16298 4323 16312 4337
rect 21170 4323 21184 4337
rect 24218 4323 24232 4337
rect 24602 4323 24616 4337
rect 70 4299 84 4313
rect 7562 4299 7576 4313
rect 7682 4299 7696 4313
rect 16778 4299 16792 4313
rect 26714 4299 26728 4313
rect 1610 4275 1624 4289
rect 10994 4275 11008 4289
rect 25754 4275 25768 4289
rect 1634 4251 1648 4265
rect 2930 4251 2944 4265
rect 2978 4251 2992 4265
rect 6650 4251 6664 4265
rect 7922 4251 7936 4265
rect 14330 4251 14344 4265
rect 16730 4251 16744 4265
rect 20090 4251 20104 4265
rect 20402 4251 20416 4265
rect 20546 4251 20560 4265
rect 20666 4251 20680 4265
rect 20930 4251 20944 4265
rect 21338 4251 21352 4265
rect 21410 4251 21424 4265
rect 21770 4251 21784 4265
rect 22154 4251 22168 4265
rect 22298 4251 22312 4265
rect 22538 4251 22552 4265
rect 22850 4251 22864 4265
rect 26258 4251 26272 4265
rect 26402 4251 26416 4265
rect 1682 4227 1696 4241
rect 4514 4227 4528 4241
rect 4562 4227 4576 4241
rect 21482 4227 21496 4241
rect 21986 4227 22000 4241
rect 22454 4227 22468 4241
rect 22946 4227 22960 4241
rect 25082 4227 25096 4241
rect 1730 4203 1744 4217
rect 13034 4203 13048 4217
rect 13082 4203 13096 4217
rect 13106 4203 13120 4217
rect 13490 4203 13504 4217
rect 13562 4203 13576 4217
rect 13778 4203 13792 4217
rect 20378 4203 20392 4217
rect 21482 4203 21496 4217
rect 21530 4203 21544 4217
rect 22082 4203 22096 4217
rect 26186 4203 26200 4217
rect 1850 4179 1864 4193
rect 12482 4179 12496 4193
rect 12554 4179 12568 4193
rect 17858 4179 17872 4193
rect 18122 4179 18136 4193
rect 18170 4179 18184 4193
rect 19106 4179 19120 4193
rect 19154 4179 19168 4193
rect 19202 4179 19216 4193
rect 19802 4179 19816 4193
rect 19946 4179 19960 4193
rect 20294 4179 20308 4193
rect 23066 4179 23080 4193
rect 23402 4179 23416 4193
rect 24266 4179 24280 4193
rect 24794 4179 24808 4193
rect 2138 4155 2152 4169
rect 7250 4155 7264 4169
rect 13274 4155 13288 4169
rect 18242 4155 18256 4169
rect 18962 4155 18976 4169
rect 20450 4155 20464 4169
rect 20762 4155 20776 4169
rect 21218 4155 21232 4169
rect 22154 4155 22168 4169
rect 22274 4155 22288 4169
rect 23210 4155 23224 4169
rect 26954 4155 26968 4169
rect 2186 4131 2200 4145
rect 2594 4131 2608 4145
rect 6242 4131 6256 4145
rect 6602 4131 6616 4145
rect 6986 4131 7000 4145
rect 8618 4131 8632 4145
rect 10922 4131 10936 4145
rect 12602 4131 12616 4145
rect 14018 4131 14032 4145
rect 23786 4131 23800 4145
rect 23978 4131 23992 4145
rect 2330 4107 2344 4121
rect 2618 4107 2632 4121
rect 5858 4107 5872 4121
rect 12722 4107 12736 4121
rect 14114 4107 14128 4121
rect 14210 4107 14224 4121
rect 15890 4107 15904 4121
rect 16418 4107 16432 4121
rect 19058 4107 19072 4121
rect 23114 4107 23128 4121
rect 23402 4107 23416 4121
rect 24842 4107 24856 4121
rect 2354 4083 2368 4097
rect 8306 4083 8320 4097
rect 8354 4083 8368 4097
rect 11354 4083 11368 4097
rect 11954 4083 11968 4097
rect 24314 4083 24328 4097
rect 2354 4059 2368 4073
rect 6890 4059 6904 4073
rect 7946 4059 7960 4073
rect 8570 4059 8584 4073
rect 13634 4059 13648 4073
rect 15842 4059 15856 4073
rect 24554 4059 24568 4073
rect 2378 4035 2392 4049
rect 22442 4035 22456 4049
rect 23786 4035 23800 4049
rect 24146 4035 24160 4049
rect 2378 4011 2392 4025
rect 20186 4011 20200 4025
rect 20210 4011 20224 4025
rect 20450 4011 20464 4025
rect 20702 4011 20716 4025
rect 2402 3987 2416 4001
rect 2738 3987 2752 4001
rect 2786 3987 2800 4001
rect 26570 3987 26584 4001
rect 2426 3963 2440 3977
rect 5930 3963 5944 3977
rect 7010 3963 7024 3977
rect 11234 3963 11248 3977
rect 12050 3963 12064 3977
rect 13586 3963 13600 3977
rect 14954 3963 14968 3977
rect 15914 3963 15928 3977
rect 17162 3963 17176 3977
rect 17810 3963 17824 3977
rect 18098 3963 18112 3977
rect 19706 3963 19720 3977
rect 26354 3963 26368 3977
rect 2450 3939 2464 3953
rect 4034 3939 4048 3953
rect 20282 3939 20296 3953
rect 26474 3939 26488 3953
rect 2474 3915 2488 3929
rect 4370 3915 4384 3929
rect 11162 3915 11176 3929
rect 14090 3915 14104 3929
rect 16802 3915 16816 3929
rect 20042 3915 20056 3929
rect 21122 3915 21136 3929
rect 23330 3915 23344 3929
rect 26474 3915 26488 3929
rect 26774 3915 26788 3929
rect 2546 3891 2560 3905
rect 3434 3891 3448 3905
rect 3746 3891 3760 3905
rect 3986 3891 4000 3905
rect 7130 3891 7144 3905
rect 13730 3891 13744 3905
rect 15002 3891 15016 3905
rect 24242 3891 24256 3905
rect 2570 3867 2584 3881
rect 19010 3867 19024 3881
rect 19610 3867 19624 3881
rect 22898 3867 22912 3881
rect 26594 3867 26608 3881
rect 2714 3843 2728 3857
rect 10490 3843 10504 3857
rect 10538 3843 10552 3857
rect 16058 3843 16072 3857
rect 16370 3843 16384 3857
rect 27074 3843 27088 3857
rect 3098 3819 3112 3833
rect 21866 3819 21880 3833
rect 3098 3795 3112 3809
rect 5066 3795 5080 3809
rect 5138 3795 5152 3809
rect 8714 3795 8728 3809
rect 9338 3795 9352 3809
rect 16538 3795 16552 3809
rect 19850 3795 19864 3809
rect 21242 3795 21256 3809
rect 24074 3795 24088 3809
rect 24530 3795 24544 3809
rect 25946 3795 25960 3809
rect 3290 3771 3304 3785
rect 6146 3771 6160 3785
rect 8186 3771 8200 3785
rect 8618 3771 8632 3785
rect 8858 3771 8872 3785
rect 9002 3771 9016 3785
rect 9098 3771 9112 3785
rect 10514 3771 10528 3785
rect 12386 3771 12400 3785
rect 18218 3771 18232 3785
rect 19898 3771 19912 3785
rect 20114 3771 20128 3785
rect 21074 3771 21088 3785
rect 3338 3747 3352 3761
rect 6434 3747 6448 3761
rect 15866 3747 15880 3761
rect 20858 3747 20872 3761
rect 3386 3723 3400 3737
rect 6098 3723 6112 3737
rect 22562 3723 22576 3737
rect 3434 3699 3448 3713
rect 10826 3699 10840 3713
rect 13898 3699 13912 3713
rect 20738 3699 20752 3713
rect 20858 3699 20872 3713
rect 26882 3699 26896 3713
rect 3506 3675 3520 3689
rect 4274 3675 4288 3689
rect 9746 3675 9760 3689
rect 12770 3675 12784 3689
rect 22706 3675 22720 3689
rect 3602 3651 3616 3665
rect 26162 3651 26176 3665
rect 3602 3627 3616 3641
rect 9146 3627 9160 3641
rect 9242 3627 9256 3641
rect 27050 3627 27064 3641
rect 3722 3603 3736 3617
rect 5666 3603 5680 3617
rect 7634 3603 7648 3617
rect 12962 3603 12976 3617
rect 13850 3603 13864 3617
rect 20498 3603 20512 3617
rect 24338 3603 24352 3617
rect 3794 3579 3808 3593
rect 5570 3579 5584 3593
rect 5618 3579 5632 3593
rect 20234 3579 20248 3593
rect 22562 3579 22576 3593
rect 22826 3579 22840 3593
rect 3842 3555 3856 3569
rect 5258 3555 5272 3569
rect 6866 3555 6880 3569
rect 12530 3555 12544 3569
rect 19346 3555 19360 3569
rect 19994 3555 20008 3569
rect 3938 3531 3952 3545
rect 11186 3531 11200 3545
rect 11306 3531 11320 3545
rect 19442 3531 19456 3545
rect 3986 3507 4000 3521
rect 19322 3507 19336 3521
rect 4154 3483 4168 3497
rect 6674 3483 6688 3497
rect 13154 3483 13168 3497
rect 21098 3483 21112 3497
rect 23186 3483 23200 3497
rect 26834 3483 26848 3497
rect 4178 3459 4192 3473
rect 7298 3459 7312 3473
rect 24626 3459 24640 3473
rect 4298 3435 4312 3449
rect 19562 3435 19576 3449
rect 4490 3411 4504 3425
rect 5090 3411 5104 3425
rect 5162 3411 5176 3425
rect 10850 3411 10864 3425
rect 18314 3411 18328 3425
rect 19322 3411 19336 3425
rect 19382 3411 19396 3425
rect 4586 3387 4600 3401
rect 9194 3387 9208 3401
rect 9290 3387 9304 3401
rect 16034 3387 16048 3401
rect 16562 3387 16576 3401
rect 25586 3387 25600 3401
rect 4706 3363 4720 3377
rect 8738 3363 8752 3377
rect 23546 3363 23560 3377
rect 25490 3363 25504 3377
rect 4874 3339 4888 3353
rect 10730 3339 10744 3353
rect 10898 3339 10912 3353
rect 16610 3339 16624 3353
rect 16754 3339 16768 3353
rect 23306 3339 23320 3353
rect 4994 3315 5008 3329
rect 21458 3315 21472 3329
rect 5186 3291 5200 3305
rect 11018 3291 11032 3305
rect 11066 3291 11080 3305
rect 12074 3291 12088 3305
rect 22490 3291 22504 3305
rect 5354 3267 5368 3281
rect 19922 3267 19936 3281
rect 25010 3267 25024 3281
rect 5522 3243 5536 3257
rect 8090 3243 8104 3257
rect 8810 3243 8824 3257
rect 10202 3243 10216 3257
rect 14042 3243 14056 3257
rect 17018 3243 17032 3257
rect 20234 3243 20248 3257
rect 23138 3243 23152 3257
rect 25850 3243 25864 3257
rect 5546 3219 5560 3233
rect 9650 3219 9664 3233
rect 9770 3219 9784 3233
rect 9818 3219 9832 3233
rect 10058 3219 10072 3233
rect 24938 3219 24952 3233
rect 5546 3195 5560 3209
rect 22994 3195 23008 3209
rect 5594 3171 5608 3185
rect 11882 3171 11896 3185
rect 13514 3171 13528 3185
rect 19586 3171 19600 3185
rect 21434 3171 21448 3185
rect 5618 3147 5632 3161
rect 6770 3147 6784 3161
rect 8234 3147 8248 3161
rect 9770 3147 9784 3161
rect 11498 3147 11512 3161
rect 12506 3147 12520 3161
rect 13586 3147 13600 3161
rect 19490 3147 19504 3161
rect 25082 3147 25096 3161
rect 26450 3147 26464 3161
rect 5690 3123 5704 3137
rect 10178 3123 10192 3137
rect 10226 3123 10240 3137
rect 19514 3123 19528 3137
rect 5762 3099 5776 3113
rect 17402 3099 17416 3113
rect 17498 3099 17512 3113
rect 20882 3099 20896 3113
rect 5858 3075 5872 3089
rect 10706 3075 10720 3089
rect 10994 3075 11008 3089
rect 11330 3075 11344 3089
rect 11618 3075 11632 3089
rect 23930 3075 23944 3089
rect 5906 3051 5920 3065
rect 7034 3051 7048 3065
rect 8882 3051 8896 3065
rect 10034 3051 10048 3065
rect 10082 3051 10096 3065
rect 24458 3051 24472 3065
rect 6002 3027 6016 3041
rect 7034 3027 7048 3041
rect 11138 3027 11152 3041
rect 11210 3027 11224 3041
rect 26666 3027 26680 3041
rect 6194 3003 6208 3017
rect 6362 3003 6376 3017
rect 6434 3003 6448 3017
rect 14258 3003 14272 3017
rect 14450 3003 14464 3017
rect 25994 3003 26008 3017
rect 6194 2979 6208 2993
rect 22874 2979 22888 2993
rect 6266 2955 6280 2969
rect 12146 2955 12160 2969
rect 12458 2955 12472 2969
rect 24722 2955 24736 2969
rect 6290 2931 6304 2945
rect 9026 2931 9040 2945
rect 9074 2931 9088 2945
rect 9602 2931 9616 2945
rect 13346 2931 13360 2945
rect 13514 2931 13528 2945
rect 22586 2931 22600 2945
rect 6338 2907 6352 2921
rect 17066 2907 17080 2921
rect 17186 2907 17200 2921
rect 25706 2907 25720 2921
rect 6386 2883 6400 2897
rect 23450 2883 23464 2897
rect 6482 2859 6496 2873
rect 8978 2859 8992 2873
rect 11978 2859 11992 2873
rect 15818 2859 15832 2873
rect 20738 2859 20752 2873
rect 6746 2835 6760 2849
rect 9434 2835 9448 2849
rect 9530 2835 9544 2849
rect 10562 2835 10576 2849
rect 11090 2835 11104 2849
rect 21242 2835 21256 2849
rect 22370 2835 22384 2849
rect 26042 2835 26056 2849
rect 6770 2811 6784 2825
rect 6794 2811 6808 2825
rect 6842 2811 6856 2825
rect 22610 2811 22624 2825
rect 23354 2811 23368 2825
rect 6794 2787 6808 2801
rect 21386 2787 21400 2801
rect 22610 2787 22624 2801
rect 26114 2787 26128 2801
rect 26306 2787 26320 2801
rect 6866 2763 6880 2777
rect 20522 2763 20536 2777
rect 21386 2763 21400 2777
rect 21506 2763 21520 2777
rect 6938 2739 6952 2753
rect 26186 2739 26200 2753
rect 6938 2715 6952 2729
rect 25274 2715 25288 2729
rect 7082 2691 7096 2705
rect 7970 2691 7984 2705
rect 8642 2691 8656 2705
rect 9866 2691 9880 2705
rect 10178 2691 10192 2705
rect 11954 2691 11968 2705
rect 16010 2691 16024 2705
rect 16202 2691 16216 2705
rect 17762 2691 17776 2705
rect 22226 2691 22240 2705
rect 25514 2691 25528 2705
rect 7130 2667 7144 2681
rect 7826 2667 7840 2681
rect 11762 2667 11776 2681
rect 13250 2667 13264 2681
rect 16994 2667 17008 2681
rect 17738 2667 17752 2681
rect 20702 2667 20716 2681
rect 24098 2667 24112 2681
rect 7154 2643 7168 2657
rect 17642 2643 17656 2657
rect 17882 2643 17896 2657
rect 17906 2643 17920 2657
rect 7202 2619 7216 2633
rect 7226 2619 7240 2633
rect 7274 2619 7288 2633
rect 9050 2619 9064 2633
rect 9098 2619 9112 2633
rect 14810 2619 14824 2633
rect 17474 2619 17488 2633
rect 7274 2595 7288 2609
rect 8018 2595 8032 2609
rect 12266 2595 12280 2609
rect 14066 2595 14080 2609
rect 17378 2595 17392 2609
rect 22970 2595 22984 2609
rect 7346 2571 7360 2585
rect 11738 2571 11752 2585
rect 11786 2571 11800 2585
rect 22658 2571 22672 2585
rect 7394 2547 7408 2561
rect 14138 2547 14152 2561
rect 23690 2547 23704 2561
rect 7418 2523 7432 2537
rect 9794 2523 9808 2537
rect 24194 2523 24208 2537
rect 7514 2499 7528 2513
rect 19274 2499 19288 2513
rect 7538 2475 7552 2489
rect 7586 2475 7600 2489
rect 7730 2475 7744 2489
rect 17522 2475 17536 2489
rect 7730 2451 7744 2465
rect 9698 2451 9712 2465
rect 10130 2451 10144 2465
rect 14162 2451 14176 2465
rect 18554 2451 18568 2465
rect 19970 2451 19984 2465
rect 20798 2451 20812 2465
rect 7874 2427 7888 2441
rect 7898 2427 7912 2441
rect 7970 2427 7984 2441
rect 8810 2427 8824 2441
rect 14282 2427 14296 2441
rect 21002 2427 21016 2441
rect 23738 2427 23752 2441
rect 23882 2427 23896 2441
rect 8042 2403 8056 2417
rect 11258 2403 11272 2417
rect 17138 2403 17152 2417
rect 19970 2403 19984 2417
rect 26282 2403 26296 2417
rect 26378 2403 26392 2417
rect 8282 2379 8296 2393
rect 8546 2379 8560 2393
rect 12410 2379 12424 2393
rect 22034 2379 22048 2393
rect 8378 2355 8392 2369
rect 21962 2355 21976 2369
rect 8402 2331 8416 2345
rect 8426 2331 8440 2345
rect 8498 2331 8512 2345
rect 9746 2331 9760 2345
rect 10418 2331 10432 2345
rect 10442 2331 10456 2345
rect 21266 2331 21280 2345
rect 21362 2331 21376 2345
rect 22130 2331 22144 2345
rect 23474 2331 23488 2345
rect 24410 2331 24424 2345
rect 24482 2331 24496 2345
rect 8498 2307 8512 2321
rect 13538 2307 13552 2321
rect 20258 2307 20272 2321
rect 23042 2307 23056 2321
rect 23546 2307 23560 2321
rect 8522 2283 8536 2297
rect 15698 2283 15712 2297
rect 15866 2283 15880 2297
rect 19466 2283 19480 2297
rect 21962 2283 21976 2297
rect 22010 2283 22024 2297
rect 8666 2259 8680 2273
rect 17450 2259 17464 2273
rect 8834 2235 8848 2249
rect 8906 2235 8920 2249
rect 8978 2235 8992 2249
rect 23246 2235 23260 2249
rect 9146 2211 9160 2225
rect 9362 2211 9376 2225
rect 9410 2211 9424 2225
rect 13418 2211 13432 2225
rect 23018 2211 23032 2225
rect 9194 2187 9208 2201
rect 9266 2187 9280 2201
rect 9314 2187 9328 2201
rect 16490 2187 16504 2201
rect 23282 2187 23296 2201
rect 9578 2163 9592 2177
rect 20474 2163 20488 2177
rect 9578 2139 9592 2153
rect 25898 2139 25912 2153
rect 9626 2115 9640 2129
rect 19490 2115 19504 2129
rect 9698 2091 9712 2105
rect 9818 2091 9832 2105
rect 10250 2091 10264 2105
rect 15962 2091 15976 2105
rect 16610 2091 16624 2105
rect 26690 2091 26704 2105
rect 10586 2067 10600 2081
rect 10610 2067 10624 2081
rect 11162 2067 11176 2081
rect 11354 2067 11368 2081
rect 11642 2067 11656 2081
rect 13682 2067 13696 2081
rect 13802 2067 13816 2081
rect 16082 2067 16096 2081
rect 24386 2067 24400 2081
rect 12506 2043 12520 2057
rect 22730 2043 22744 2057
rect 12602 2019 12616 2033
rect 12698 2019 12712 2033
rect 12818 2019 12832 2033
rect 17570 2019 17584 2033
rect 20570 2019 20584 2033
rect 20618 2019 20632 2033
rect 12914 1995 12928 2009
rect 14930 1995 14944 2009
rect 26618 1995 26632 2009
rect 13106 1971 13120 1985
rect 27026 1971 27040 1985
rect 13274 1947 13288 1961
rect 13394 1947 13408 1961
rect 13826 1947 13840 1961
rect 19058 1947 19072 1961
rect 19418 1947 19432 1961
rect 20618 1947 20632 1961
rect 20702 1947 20716 1961
rect 13874 1923 13888 1937
rect 13922 1923 13936 1937
rect 14066 1923 14080 1937
rect 14186 1923 14200 1937
rect 14666 1923 14680 1937
rect 14690 1923 14704 1937
rect 14906 1923 14920 1937
rect 27445 1923 27459 1937
rect 13922 1899 13936 1913
rect 15626 1899 15640 1913
rect 15914 1899 15928 1913
rect 22634 1899 22648 1913
rect 24290 1899 24304 1913
rect 24338 1899 24352 1913
rect 26258 1899 26272 1913
rect 14138 1875 14152 1889
rect 20786 1875 20800 1889
rect 25970 1875 25984 1889
rect 27074 1875 27088 1889
rect 27445 1875 27459 1889
rect 16082 1851 16096 1865
rect 17978 1851 17992 1865
rect 23834 1851 23848 1865
rect 25970 1851 25984 1865
rect 26018 1851 26032 1865
rect 27050 1851 27064 1865
rect 27445 1851 27459 1865
rect 16778 1827 16792 1841
rect 16922 1827 16936 1841
rect 16994 1827 17008 1841
rect 18362 1827 18376 1841
rect 27026 1827 27040 1841
rect 27445 1827 27459 1841
rect 18074 994 18088 1008
rect 18290 994 18304 1008
rect 18050 970 18064 984
rect 25274 970 25288 984
rect 17570 946 17584 960
rect 18146 946 18160 960
rect 11042 922 11056 936
rect 18962 922 18976 936
rect 10946 898 10960 912
rect 18098 898 18112 912
rect 19010 898 19024 912
rect 26450 898 26464 912
rect 10826 874 10840 888
rect 16226 874 16240 888
rect 16466 874 16480 888
rect 21746 874 21760 888
rect 10634 850 10648 864
rect 15098 850 15112 864
rect 15962 850 15976 864
rect 16010 850 16024 864
rect 19394 850 19408 864
rect 9410 826 9424 840
rect 9890 826 9904 840
rect 10106 826 10120 840
rect 21938 826 21952 840
rect 9338 802 9352 816
rect 13562 802 13576 816
rect 14426 802 14440 816
rect 24458 802 24472 816
rect 9050 778 9064 792
rect 19346 778 19360 792
rect 8762 754 8776 768
rect 12842 754 12856 768
rect 12986 754 13000 768
rect 13610 754 13624 768
rect 13946 754 13960 768
rect 19538 754 19552 768
rect 22994 754 23008 768
rect 26282 754 26296 768
rect 8426 730 8440 744
rect 26114 730 26128 744
rect 8258 706 8272 720
rect 13322 706 13336 720
rect 13730 706 13744 720
rect 24098 706 24112 720
rect 7934 682 7948 696
rect 9698 682 9712 696
rect 9866 682 9880 696
rect 21506 682 21520 696
rect 21578 682 21592 696
rect 24554 682 24568 696
rect 7754 658 7768 672
rect 26378 658 26392 672
rect 7562 634 7576 648
rect 11258 634 11272 648
rect 12362 634 12376 648
rect 14474 634 14488 648
rect 14522 634 14536 648
rect 19658 634 19672 648
rect 24362 634 24376 648
rect 7226 610 7240 624
rect 19178 610 19192 624
rect 19466 610 19480 624
rect 20066 610 20080 624
rect 21410 610 21424 624
rect 25418 610 25432 624
rect 6578 586 6592 600
rect 19778 586 19792 600
rect 21362 586 21376 600
rect 23498 586 23512 600
rect 6386 562 6400 576
rect 13130 562 13144 576
rect 13394 562 13408 576
rect 13682 562 13696 576
rect 14570 562 14584 576
rect 14858 562 14872 576
rect 19586 562 19600 576
rect 19730 562 19744 576
rect 20522 562 20536 576
rect 20570 562 20584 576
rect 26594 562 26608 576
rect 6314 538 6328 552
rect 26138 538 26152 552
rect 6242 514 6256 528
rect 16682 514 16696 528
rect 17258 514 17272 528
rect 27445 514 27459 528
rect 5954 490 5968 504
rect 24194 490 24208 504
rect 5738 466 5752 480
rect 20930 466 20944 480
rect 5642 442 5656 456
rect 21314 442 21328 456
rect 5498 418 5512 432
rect 22658 418 22672 432
rect 4778 394 4792 408
rect 6626 394 6640 408
rect 6818 394 6832 408
rect 24674 394 24688 408
rect 4754 370 4768 384
rect 14378 370 14392 384
rect 14906 370 14920 384
rect 21698 370 21712 384
rect 4538 346 4552 360
rect 12410 346 12424 360
rect 12530 346 12544 360
rect 14690 346 14704 360
rect 15146 346 15160 360
rect 17810 346 17824 360
rect 24242 346 24256 360
rect 4370 322 4384 336
rect 10322 322 10336 336
rect 10706 322 10720 336
rect 10754 322 10768 336
rect 24506 322 24520 336
rect 4322 298 4336 312
rect 26018 298 26032 312
rect 3890 274 3904 288
rect 4802 274 4816 288
rect 4946 274 4960 288
rect 26042 274 26056 288
rect 3674 250 3688 264
rect 19418 250 19432 264
rect 3626 226 3640 240
rect 12314 226 12328 240
rect 14306 226 14320 240
rect 22730 226 22744 240
rect 3554 202 3568 216
rect 6410 202 6424 216
rect 6530 202 6544 216
rect 22058 202 22072 216
rect 23234 202 23248 216
rect 2498 178 2512 192
rect 20882 178 20896 192
rect 1778 154 1792 168
rect 4826 154 4840 168
rect 5306 154 5320 168
rect 22826 154 22840 168
rect 1658 130 1672 144
rect 9482 130 9496 144
rect 10538 130 10552 144
rect 12266 130 12280 144
rect 15266 130 15280 144
rect 18818 130 18832 144
rect 70 106 84 120
rect 21626 106 21640 120
rect 70 82 84 96
rect 17930 82 17944 96
rect 17978 82 17992 96
rect 18410 82 18424 96
rect 3530 58 3544 72
rect 20690 58 20704 72
rect 26570 58 26584 72
rect 27445 58 27459 72
rect 4298 34 4312 48
rect 14330 34 14344 48
rect 16130 34 16144 48
rect 16322 34 16336 48
rect 17282 34 17296 48
rect 25994 34 26008 48
rect 26570 34 26584 48
rect 27445 34 27459 48
rect 17882 10 17896 24
rect 26570 10 26584 24
rect 26594 10 26608 24
rect 27445 10 27459 24
<< metal2 >>
rect 0 8349 70 8361
rect 0 8325 70 8337
rect 123 8050 323 8444
rect 339 8050 351 8444
rect 363 8050 375 8444
rect 387 8050 399 8444
rect 411 8050 423 8444
rect 1731 8050 1743 8324
rect 1995 8050 2007 8324
rect 2139 8050 2151 8300
rect 2283 8050 2295 8372
rect 2415 8290 2427 8444
rect 2451 8338 2463 8444
rect 3531 8050 3543 8324
rect 3555 8050 3567 8300
rect 4119 8266 4131 8444
rect 4203 8050 4215 8228
rect 4971 8218 4983 8444
rect 5823 8194 5835 8444
rect 6279 8194 6291 8444
rect 7527 8194 7539 8444
rect 7563 8338 7575 8444
rect 9231 8338 9243 8444
rect 9267 8290 9279 8444
rect 6280 8180 6298 8194
rect 6075 8050 6087 8180
rect 6267 8050 6279 8180
rect 7947 8050 7959 8252
rect 7971 8050 7983 8276
rect 8331 8050 8343 8276
rect 8811 8050 8823 8204
rect 9459 8050 9471 8276
rect 9939 8050 9951 8180
rect 10755 8050 10767 8252
rect 10935 8218 10947 8444
rect 11451 8050 11463 8180
rect 11787 8170 11799 8444
rect 12639 8146 12651 8444
rect 12675 8290 12687 8444
rect 13815 8410 13827 8444
rect 13816 8396 13834 8410
rect 12867 8050 12879 8276
rect 13803 8050 13815 8396
rect 14667 8050 14679 8396
rect 15183 8122 15195 8444
rect 15711 8434 15723 8444
rect 16863 8434 16875 8444
rect 15712 8420 15730 8434
rect 15699 8050 15711 8420
rect 17703 8098 17715 8444
rect 17727 8386 17739 8444
rect 19383 8338 19395 8444
rect 17716 8084 17734 8098
rect 17715 8050 17727 8084
rect 18651 8050 18663 8084
rect 19155 8050 19167 8324
rect 19407 8194 19419 8444
rect 19419 8050 19431 8060
rect 20283 8050 20295 8420
rect 20547 8050 20559 8324
rect 20703 8194 20715 8444
rect 21903 8338 21915 8444
rect 20704 8180 20722 8194
rect 20691 8050 20703 8180
rect 20931 8050 20943 8156
rect 22011 8050 22023 8300
rect 22155 8050 22167 8324
rect 22407 8194 22419 8444
rect 22767 8410 22779 8444
rect 22408 8180 22426 8194
rect 22395 8050 22407 8180
rect 23139 8050 23151 8348
rect 24423 8338 24435 8444
rect 24447 8290 24459 8444
rect 23403 8050 23415 8108
rect 24147 8050 24159 8132
rect 24795 8050 24807 8180
rect 25011 8050 25023 8324
rect 25287 8314 25299 8444
rect 26127 8266 26139 8444
rect 25779 8050 25791 8204
rect 27027 8050 27039 8252
rect 27051 8122 27063 8252
rect 27075 8146 27087 8228
rect 27099 8074 27111 8156
rect 27123 8074 27135 8180
rect 27171 8050 27371 8444
rect 27459 8157 27529 8169
rect 27459 8133 27529 8145
rect 27459 8109 27529 8121
rect 27459 8085 27529 8097
rect 27459 8061 27529 8073
rect 0 4324 70 4336
rect 0 4300 70 4312
rect 123 1817 323 7251
rect 339 1817 351 7251
rect 363 1817 375 7251
rect 387 1817 399 7251
rect 411 1817 423 7251
rect 1611 4361 1623 7251
rect 1635 4385 1647 7251
rect 1659 4409 1671 7251
rect 1611 1817 1623 4275
rect 1635 1817 1647 4251
rect 1683 4241 1695 7251
rect 1731 4217 1743 7251
rect 1779 4433 1791 7251
rect 1803 4457 1815 7251
rect 1827 4481 1839 7251
rect 1851 4193 1863 7251
rect 1899 4505 1911 7251
rect 1923 4361 1935 7251
rect 1947 4529 1959 7251
rect 1995 4409 2007 7251
rect 2043 4553 2055 7251
rect 2115 4577 2127 7251
rect 2163 4601 2175 7251
rect 2211 4625 2223 7251
rect 2235 4649 2247 7251
rect 2331 4673 2343 7251
rect 2139 1817 2151 4155
rect 2187 1817 2199 4131
rect 2331 1817 2343 4107
rect 2355 4097 2367 7251
rect 2355 1817 2367 4059
rect 2379 4049 2391 7251
rect 2379 1817 2391 4011
rect 2403 4001 2415 7251
rect 2451 4697 2463 7251
rect 2475 4721 2487 7251
rect 2499 4745 2511 7251
rect 2523 4769 2535 7251
rect 2571 4793 2583 7251
rect 2595 4145 2607 7251
rect 2619 4817 2631 7251
rect 2667 4841 2679 7251
rect 2691 4865 2703 7251
rect 2427 1817 2439 3963
rect 2451 1817 2463 3939
rect 2475 1817 2487 3915
rect 2547 1817 2559 3891
rect 2571 1817 2583 3867
rect 2619 1817 2631 4107
rect 2715 3857 2727 7251
rect 2763 4889 2775 7251
rect 2787 4001 2799 7251
rect 2811 4913 2823 7251
rect 2859 4937 2871 7251
rect 2883 4961 2895 7251
rect 2907 4985 2919 7251
rect 2931 4265 2943 7251
rect 2979 4265 2991 7251
rect 3003 5009 3015 7251
rect 3027 5033 3039 7251
rect 3075 5057 3087 7251
rect 2739 1817 2751 3987
rect 3099 3833 3111 7251
rect 3123 5081 3135 7251
rect 3099 1817 3111 3795
rect 3147 1817 3159 4683
rect 3171 4601 3183 7251
rect 3195 5105 3207 7251
rect 3219 4601 3231 7251
rect 3243 5129 3255 7251
rect 3291 5153 3303 7251
rect 3315 5177 3327 7251
rect 3363 5201 3375 7251
rect 3411 4985 3423 7251
rect 3291 1817 3303 3771
rect 3315 1817 3327 4851
rect 3435 3905 3447 7251
rect 3459 4361 3471 7251
rect 3483 5225 3495 7251
rect 3531 5249 3543 7251
rect 3579 5273 3591 7251
rect 3339 1817 3351 3747
rect 3387 1817 3399 3723
rect 3435 1817 3447 3699
rect 3507 1817 3519 3675
rect 3603 3665 3615 7251
rect 3651 4457 3663 7251
rect 3675 4433 3687 7251
rect 3699 5297 3711 7251
rect 3747 5321 3759 7251
rect 3771 4961 3783 7251
rect 3795 5345 3807 7251
rect 3819 5369 3831 7251
rect 3867 5393 3879 7251
rect 3891 5369 3903 7251
rect 3939 5369 3951 7251
rect 3603 1817 3615 3627
rect 3723 1817 3735 3603
rect 3747 1817 3759 3891
rect 3771 1817 3783 4323
rect 3795 1817 3807 3579
rect 3843 1817 3855 3555
rect 3867 1817 3879 4923
rect 3939 1817 3951 3531
rect 3963 1817 3975 4467
rect 3987 3905 3999 7251
rect 4011 5345 4023 7251
rect 4059 5417 4071 7251
rect 4107 5465 4119 7251
rect 4131 5489 4143 7251
rect 4155 5513 4167 7251
rect 3987 1817 3999 3507
rect 4035 1817 4047 3939
rect 4083 1817 4095 5427
rect 4179 4769 4191 7251
rect 4155 1817 4167 3483
rect 4179 1817 4191 3459
rect 4227 1817 4239 5523
rect 4251 4961 4263 7251
rect 4275 5321 4287 7251
rect 4275 1817 4287 3675
rect 4299 3449 4311 7251
rect 4347 5561 4359 7251
rect 4371 3929 4383 7251
rect 4419 5585 4431 7251
rect 4467 5321 4479 7251
rect 4491 5609 4503 7251
rect 4539 5633 4551 7251
rect 4419 1817 4431 4779
rect 4587 4649 4599 7251
rect 4635 5657 4647 7251
rect 4707 5681 4719 7251
rect 4491 1817 4503 3411
rect 4515 1817 4527 4227
rect 4563 1817 4575 4227
rect 4587 1817 4599 3387
rect 4635 1817 4647 4827
rect 4659 1817 4671 5595
rect 4731 4697 4743 7251
rect 4779 5705 4791 7251
rect 4827 4937 4839 7251
rect 4851 4985 4863 7251
rect 4707 1817 4719 3363
rect 4875 3353 4887 7251
rect 4923 5729 4935 7251
rect 4947 5585 4959 7251
rect 4995 3329 5007 7251
rect 5043 5753 5055 7251
rect 5067 3809 5079 7251
rect 5091 3425 5103 7251
rect 5139 3809 5151 7251
rect 5163 3425 5175 7251
rect 5187 3305 5199 7251
rect 5235 5081 5247 7251
rect 5259 3569 5271 7251
rect 5283 5081 5295 7251
rect 5331 5777 5343 7251
rect 5355 4553 5367 7251
rect 5403 4985 5415 7251
rect 5451 5801 5463 7251
rect 5475 5825 5487 7251
rect 5499 5849 5511 7251
rect 5355 1817 5367 3267
rect 5523 1817 5535 3243
rect 5547 3233 5559 7251
rect 5571 3593 5583 7251
rect 5619 3593 5631 7251
rect 5667 3617 5679 7251
rect 5691 5873 5703 7251
rect 5715 5897 5727 7251
rect 5547 1817 5559 3195
rect 5595 1817 5607 3171
rect 5619 1817 5631 3147
rect 5691 1817 5703 3123
rect 5715 1817 5727 4467
rect 5763 3113 5775 7251
rect 5787 5921 5799 7251
rect 5811 5945 5823 7251
rect 5787 1817 5799 5307
rect 5811 1817 5823 5403
rect 5835 1817 5847 4827
rect 5859 4121 5871 7251
rect 5883 5969 5895 7251
rect 5907 5993 5919 7251
rect 5955 6017 5967 7251
rect 5979 5705 5991 7251
rect 6003 6041 6015 7251
rect 6051 5321 6063 7251
rect 5859 1817 5871 3075
rect 5907 1817 5919 3051
rect 5931 1817 5943 3963
rect 6003 1817 6015 3027
rect 6051 1817 6063 4371
rect 6075 4361 6087 7251
rect 6099 3737 6111 7251
rect 6123 1817 6135 5331
rect 6147 4577 6159 7251
rect 6171 6065 6183 7251
rect 6147 1817 6159 3771
rect 6171 1817 6183 4395
rect 6195 3017 6207 7251
rect 6243 4145 6255 7251
rect 6267 6089 6279 7251
rect 6195 1817 6207 2979
rect 6267 1817 6279 2955
rect 6291 2945 6303 7251
rect 6339 2921 6351 7251
rect 6363 6113 6375 7251
rect 6363 1817 6375 3003
rect 6387 2897 6399 7251
rect 6435 3761 6447 7251
rect 6483 4481 6495 7251
rect 6555 6137 6567 7251
rect 6579 6161 6591 7251
rect 6603 6185 6615 7251
rect 6435 1817 6447 3003
rect 6483 1817 6495 2859
rect 6507 1817 6519 4467
rect 6651 4265 6663 7251
rect 6675 6209 6687 7251
rect 6699 6233 6711 7251
rect 6603 1817 6615 4131
rect 6675 1817 6687 3483
rect 6699 1817 6711 4539
rect 6723 1817 6735 6243
rect 6747 2849 6759 7251
rect 6771 3161 6783 7251
rect 6795 2825 6807 7251
rect 6843 2825 6855 7251
rect 6867 3569 6879 7251
rect 6891 6281 6903 7251
rect 6771 1817 6783 2811
rect 6795 1817 6807 2787
rect 6867 1817 6879 2763
rect 6891 1817 6903 4059
rect 6939 2753 6951 7251
rect 6963 5201 6975 7251
rect 6987 6305 6999 7251
rect 6939 1817 6951 2715
rect 6987 1817 6999 4131
rect 7011 1817 7023 3963
rect 7035 3065 7047 7251
rect 7059 4841 7071 7251
rect 7083 6329 7095 7251
rect 7035 1817 7047 3027
rect 7083 1817 7095 2691
rect 7107 1817 7119 4347
rect 7131 3905 7143 7251
rect 7131 1817 7143 2667
rect 7155 2657 7167 7251
rect 7179 6353 7191 7251
rect 7179 1817 7191 5235
rect 7203 4577 7215 7251
rect 7227 2633 7239 5259
rect 7251 4169 7263 7251
rect 7275 2633 7287 7251
rect 7299 6377 7311 7251
rect 7347 6257 7359 7251
rect 7371 6401 7383 7251
rect 7395 6257 7407 7251
rect 7419 6425 7431 7251
rect 7443 4889 7455 7251
rect 7491 6281 7503 7251
rect 7515 6449 7527 7251
rect 7539 5033 7551 7251
rect 7203 1817 7215 2619
rect 7275 1817 7287 2595
rect 7299 1817 7311 3459
rect 7347 1817 7359 2571
rect 7395 1817 7407 2547
rect 7419 1817 7431 2523
rect 7467 1817 7479 4611
rect 7563 4313 7575 7251
rect 7515 1817 7527 2499
rect 7587 2489 7599 5451
rect 7611 5033 7623 7251
rect 7539 1817 7551 2475
rect 7611 1817 7623 4947
rect 7659 4721 7671 7251
rect 7635 1817 7647 3603
rect 7683 1817 7695 4299
rect 7731 2489 7743 7251
rect 7755 6473 7767 7251
rect 7779 6497 7791 7251
rect 7731 1817 7743 2451
rect 7803 1817 7815 6507
rect 7827 2681 7839 7251
rect 7875 5345 7887 7251
rect 7851 1817 7863 4923
rect 7899 2441 7911 5667
rect 7875 1817 7887 2427
rect 7923 1817 7935 4251
rect 7947 4073 7959 7251
rect 7971 2705 7983 7251
rect 7971 1817 7983 2427
rect 7995 1817 8007 4851
rect 8019 2609 8031 7251
rect 8067 5033 8079 7251
rect 8091 4697 8103 7251
rect 8115 4673 8127 7251
rect 8043 1817 8055 2403
rect 8091 1817 8103 3243
rect 8139 1817 8151 4851
rect 8163 4673 8175 7251
rect 8187 3785 8199 7251
rect 8211 6545 8223 7251
rect 8259 6569 8271 7251
rect 8211 1817 8223 6459
rect 8283 4337 8295 7251
rect 8379 5417 8391 7251
rect 8403 5633 8415 7251
rect 8451 6593 8463 7251
rect 8235 1817 8247 3147
rect 8283 1817 8295 2379
rect 8307 1817 8319 4083
rect 8355 1817 8367 4083
rect 8379 1817 8391 2355
rect 8427 2345 8439 6075
rect 8403 1817 8415 2331
rect 8475 1817 8487 6291
rect 8499 2345 8511 7251
rect 8523 6305 8535 7251
rect 8547 2393 8559 7251
rect 8571 6617 8583 7251
rect 8619 4145 8631 7251
rect 8499 1817 8511 2307
rect 8523 1817 8535 2283
rect 8571 1817 8583 4059
rect 8619 1817 8631 3771
rect 8643 2705 8655 7251
rect 8667 2273 8679 7251
rect 8715 6473 8727 7251
rect 8691 1817 8703 5667
rect 8715 1817 8727 3795
rect 8739 3377 8751 7251
rect 8763 6641 8775 7251
rect 8811 3257 8823 7251
rect 8835 5345 8847 7251
rect 8859 3785 8871 7251
rect 8883 4409 8895 7251
rect 8907 6665 8919 7251
rect 8955 6689 8967 7251
rect 8811 1817 8823 2427
rect 8835 1817 8847 2235
rect 8883 1817 8895 3051
rect 8907 2249 8919 5547
rect 8931 1817 8943 4707
rect 8955 1817 8967 4731
rect 8979 2873 8991 7251
rect 9003 3785 9015 7251
rect 9027 6713 9039 7251
rect 8979 1817 8991 2235
rect 9027 1817 9039 2931
rect 9051 2633 9063 6699
rect 9075 2945 9087 7251
rect 9099 3785 9111 7251
rect 9147 3641 9159 7251
rect 9099 1817 9111 2619
rect 9147 1817 9159 2211
rect 9171 1817 9183 6699
rect 9195 3401 9207 7251
rect 9219 6737 9231 7251
rect 9195 1817 9207 2187
rect 9219 1817 9231 5859
rect 9243 1817 9255 3627
rect 9267 2201 9279 7251
rect 9315 4745 9327 7251
rect 9339 3809 9351 7251
rect 9363 6761 9375 7251
rect 9291 1817 9303 3387
rect 9363 2225 9375 5835
rect 9315 1817 9327 2187
rect 9387 1817 9399 6123
rect 9411 2225 9423 7251
rect 9435 6785 9447 7251
rect 9507 4697 9519 7251
rect 9435 1817 9447 2835
rect 9507 1817 9519 4347
rect 9531 4337 9543 7251
rect 9531 1817 9543 2835
rect 9579 2177 9591 7251
rect 9579 1817 9591 2139
rect 9603 1817 9615 2931
rect 9627 2129 9639 7251
rect 9651 6809 9663 7251
rect 9651 1817 9663 3219
rect 9699 2465 9711 7251
rect 9747 3689 9759 7251
rect 9771 3233 9783 7251
rect 9795 4601 9807 7251
rect 9699 1817 9711 2091
rect 9747 1817 9759 2331
rect 9771 1817 9783 3147
rect 9795 1817 9807 2523
rect 9819 2105 9831 3219
rect 9843 1817 9855 5811
rect 9867 2705 9879 7251
rect 9891 4409 9903 7251
rect 9939 5273 9951 7251
rect 9939 1817 9951 4827
rect 9963 4601 9975 7251
rect 9963 1817 9975 4443
rect 9987 1817 9999 5547
rect 10011 1817 10023 5499
rect 10035 3065 10047 7251
rect 10059 5609 10071 7251
rect 10059 1817 10071 3219
rect 10083 3065 10095 7251
rect 10131 2465 10143 7251
rect 10179 3137 10191 7251
rect 10179 1817 10191 2691
rect 10203 1817 10215 3243
rect 10227 1817 10239 3123
rect 10251 2105 10263 7251
rect 10299 6833 10311 7251
rect 10371 6857 10383 7251
rect 10395 6305 10407 7251
rect 10275 1817 10287 5619
rect 10299 1817 10311 5331
rect 10371 1817 10383 4995
rect 10419 4985 10431 7251
rect 10443 6881 10455 7251
rect 10491 6857 10503 7251
rect 10515 6905 10527 7251
rect 10443 2345 10455 6843
rect 10539 3857 10551 7251
rect 10419 1817 10431 2331
rect 10491 1817 10503 3843
rect 10515 1817 10527 3771
rect 10563 2849 10575 6843
rect 10587 4529 10599 7251
rect 10635 6857 10647 7251
rect 10611 2081 10623 5211
rect 10707 3089 10719 7251
rect 10587 1817 10599 2067
rect 10731 1817 10743 3339
rect 10803 1817 10815 6651
rect 10827 3713 10839 7251
rect 10851 4841 10863 7251
rect 10875 6665 10887 7251
rect 10923 6305 10935 7251
rect 10947 4961 10959 7251
rect 10971 5777 10983 7251
rect 10995 4289 11007 7251
rect 11043 6665 11055 7251
rect 10851 1817 10863 3411
rect 10899 1817 10911 3339
rect 10923 1817 10935 4131
rect 11067 3305 11079 7251
rect 11091 6665 11103 7251
rect 10995 1817 11007 3075
rect 11019 1817 11031 3291
rect 11091 1817 11103 2835
rect 11115 1817 11127 5235
rect 11139 3041 11151 7251
rect 11163 3929 11175 7251
rect 11187 3545 11199 7251
rect 11235 3977 11247 7251
rect 11163 1817 11175 2067
rect 11211 1817 11223 3027
rect 11259 2417 11271 7251
rect 11283 4409 11295 7251
rect 11307 3545 11319 7251
rect 11355 6929 11367 7251
rect 11331 3089 11343 5859
rect 11379 5369 11391 7251
rect 11403 6833 11415 7251
rect 11427 5465 11439 7251
rect 11355 2081 11367 4083
rect 11499 3161 11511 7251
rect 11523 4697 11535 7251
rect 11547 5873 11559 7251
rect 11595 6833 11607 7251
rect 11619 3089 11631 7251
rect 11643 2081 11655 7251
rect 11667 5993 11679 7251
rect 11691 6953 11703 7251
rect 11739 2585 11751 7251
rect 11763 2681 11775 7251
rect 11787 5993 11799 7251
rect 11835 6209 11847 7251
rect 11883 3185 11895 7251
rect 11787 1817 11799 2571
rect 11931 1817 11943 4539
rect 11955 4097 11967 7251
rect 11979 6089 11991 7251
rect 12027 6977 12039 7251
rect 11955 1817 11967 2691
rect 11979 1817 11991 2859
rect 12027 1817 12039 5307
rect 12075 5249 12087 7251
rect 12099 5273 12111 7251
rect 12195 6977 12207 7251
rect 12051 1817 12063 3963
rect 12075 1817 12087 3291
rect 12123 1817 12135 6339
rect 12147 2969 12159 6963
rect 12171 1817 12183 6291
rect 12243 1817 12255 4443
rect 12267 2609 12279 7251
rect 12291 4409 12303 7251
rect 12315 5177 12327 7251
rect 12363 5177 12375 7251
rect 12387 1817 12399 3771
rect 12411 2393 12423 7251
rect 12483 7001 12495 7251
rect 12459 1817 12471 2955
rect 12483 1817 12495 4179
rect 12507 3161 12519 7251
rect 12531 3569 12543 6987
rect 12555 4961 12567 7251
rect 12507 1817 12519 2043
rect 12555 1817 12567 4179
rect 12603 4145 12615 7251
rect 12627 6473 12639 7251
rect 12651 7001 12663 7251
rect 12699 7025 12711 7251
rect 12723 6089 12735 7251
rect 12603 1817 12615 2019
rect 12627 1817 12639 5499
rect 12651 1817 12663 4755
rect 12675 1817 12687 5499
rect 12699 2033 12711 5451
rect 12723 1817 12735 4107
rect 12747 1817 12759 5331
rect 12771 3689 12783 7251
rect 12795 1817 12807 4443
rect 12819 2033 12831 7251
rect 12939 6881 12951 7251
rect 12963 7049 12975 7251
rect 12987 6881 12999 7251
rect 13011 7073 13023 7251
rect 13059 7097 13071 7251
rect 12867 1817 12879 4731
rect 12915 1817 12927 1995
rect 12963 1817 12975 3603
rect 13011 1817 13023 5859
rect 13083 4409 13095 7251
rect 13107 7121 13119 7251
rect 13107 4217 13119 4875
rect 13035 1817 13047 4203
rect 13083 1817 13095 4203
rect 13155 3497 13167 7251
rect 13179 7145 13191 7251
rect 13227 7169 13239 7251
rect 13107 1817 13119 1971
rect 13179 1817 13191 4851
rect 13203 1817 13215 5595
rect 13227 1817 13239 4659
rect 13251 2681 13263 7131
rect 13275 4169 13287 7251
rect 13299 6473 13311 7251
rect 13275 1817 13287 1947
rect 13299 1817 13311 6363
rect 13323 5801 13335 7251
rect 13347 2945 13359 7155
rect 13371 5873 13383 7251
rect 13371 1817 13383 5187
rect 13395 1961 13407 6339
rect 13419 4673 13431 7251
rect 13419 1817 13431 2211
rect 13467 1817 13479 4923
rect 13491 4721 13503 7251
rect 13491 1817 13503 4203
rect 13515 3185 13527 7251
rect 13515 1817 13527 2931
rect 13539 2321 13551 7251
rect 13563 4217 13575 5763
rect 13587 3977 13599 7251
rect 13611 5801 13623 7251
rect 13635 4073 13647 7251
rect 13659 6377 13671 7251
rect 13587 1817 13599 3147
rect 13659 1817 13671 5547
rect 13683 2081 13695 6363
rect 13707 6017 13719 7251
rect 13707 1817 13719 5331
rect 13731 3905 13743 7251
rect 13755 6377 13767 7251
rect 13803 7145 13815 7251
rect 13779 1817 13791 4203
rect 13851 3617 13863 7251
rect 13875 4985 13887 7251
rect 13899 7169 13911 7251
rect 13947 6641 13959 7251
rect 13803 1817 13815 2067
rect 13827 1817 13839 1947
rect 13875 1817 13887 1923
rect 13899 1817 13911 3699
rect 13923 1937 13935 5691
rect 13971 4361 13983 7251
rect 13995 6641 14007 7251
rect 13923 1817 13935 1899
rect 13995 1817 14007 6579
rect 14019 1817 14031 4131
rect 14043 3257 14055 7251
rect 14067 2609 14079 7251
rect 14091 3929 14103 7251
rect 14115 4409 14127 7251
rect 14139 7193 14151 7251
rect 14067 1817 14079 1923
rect 14115 1817 14127 4107
rect 14139 2561 14151 7155
rect 14139 1817 14151 1875
rect 14163 1817 14175 2451
rect 14187 1937 14199 7011
rect 14211 1817 14223 4107
rect 14235 1817 14247 4347
rect 14259 3017 14271 7251
rect 14619 7169 14631 7251
rect 14667 6065 14679 7251
rect 14283 1817 14295 2427
rect 14331 1817 14343 4251
rect 14355 1817 14367 4731
rect 14451 1817 14463 3003
rect 14643 1817 14655 4779
rect 14691 1937 14703 6123
rect 14667 1817 14679 1923
rect 14739 1817 14751 6147
rect 14787 1817 14799 6099
rect 14811 2633 14823 7251
rect 14835 4793 14847 7251
rect 14859 6113 14871 7251
rect 14883 7217 14895 7251
rect 14883 1817 14895 4371
rect 14907 1937 14919 7251
rect 15027 7217 15039 7251
rect 14931 2009 14943 7203
rect 14955 1817 14967 3963
rect 14979 1817 14991 5307
rect 15003 1817 15015 3891
rect 15027 1817 15039 5643
rect 15051 1817 15063 6771
rect 15123 1817 15135 6291
rect 15387 4937 15399 7251
rect 15435 5825 15447 7251
rect 15579 6089 15591 7251
rect 15627 1913 15639 7251
rect 15675 1817 15687 4371
rect 15699 2297 15711 7251
rect 15747 6377 15759 7251
rect 15771 6785 15783 7251
rect 15795 6377 15807 7251
rect 15819 7241 15831 7251
rect 15819 1817 15831 2859
rect 15843 1817 15855 4059
rect 15867 3761 15879 7251
rect 15891 4121 15903 7251
rect 15915 3977 15927 7251
rect 15939 6425 15951 7251
rect 15867 1817 15879 2283
rect 15915 1817 15927 1899
rect 15939 1817 15951 4923
rect 15963 2105 15975 7227
rect 15987 6641 15999 7251
rect 15987 1817 15999 4323
rect 16011 2705 16023 7251
rect 16035 3401 16047 7251
rect 16059 1817 16071 3843
rect 16083 2081 16095 7251
rect 16131 6569 16143 7251
rect 16083 1817 16095 1851
rect 16179 1817 16191 5571
rect 16203 5201 16215 7251
rect 16251 6425 16263 7251
rect 16323 5369 16335 7251
rect 16203 1817 16215 2691
rect 16275 1817 16287 5355
rect 16347 4913 16359 7251
rect 16371 6569 16383 7251
rect 16395 4769 16407 7251
rect 16443 6857 16455 7251
rect 16299 1817 16311 4323
rect 16347 1817 16359 4755
rect 16371 1817 16383 3843
rect 16419 1817 16431 4107
rect 16443 1817 16455 5763
rect 16467 4913 16479 7251
rect 16491 2201 16503 7251
rect 16515 1817 16527 7251
rect 16563 5633 16575 7251
rect 16587 6089 16599 7251
rect 16539 1817 16551 3795
rect 16563 1817 16575 3387
rect 16611 3353 16623 7251
rect 16611 1817 16623 2091
rect 16635 1817 16647 5595
rect 16659 4361 16671 7251
rect 16683 6089 16695 7251
rect 16707 4649 16719 7251
rect 16755 5777 16767 7251
rect 16779 4313 16791 7251
rect 16731 1817 16743 4251
rect 16803 3929 16815 7251
rect 16827 5633 16839 7251
rect 16755 1817 16767 3339
rect 16779 1817 16791 1827
rect 16827 1817 16839 4923
rect 16851 1817 16863 5547
rect 16875 5249 16887 7251
rect 16899 5273 16911 7251
rect 16899 1817 16911 4635
rect 16923 1841 16935 6867
rect 16947 5609 16959 7251
rect 16971 1817 16983 4923
rect 16995 2681 17007 7251
rect 17019 3257 17031 7251
rect 17043 6689 17055 7251
rect 16995 1817 17007 1827
rect 17043 1817 17055 5163
rect 17079 4649 17091 5307
rect 17163 4769 17175 7251
rect 17067 1817 17079 2907
rect 17139 1817 17151 2403
rect 17163 1817 17175 3963
rect 17187 1817 17199 2907
rect 17235 1817 17247 4875
rect 17331 1817 17343 4539
rect 17355 1817 17367 4851
rect 17379 1817 17391 2595
rect 17403 1817 17415 3099
rect 17451 1817 17463 2259
rect 17475 1817 17487 2619
rect 17499 1817 17511 3099
rect 17523 1817 17535 2475
rect 17571 2033 17583 7251
rect 17595 1817 17607 5571
rect 17715 5321 17727 7251
rect 17643 1817 17655 2643
rect 17691 1817 17703 5187
rect 17715 1817 17727 4827
rect 17763 2705 17775 7251
rect 17739 1817 17751 2667
rect 17787 1817 17799 5475
rect 17811 3977 17823 7251
rect 17835 1817 17847 6795
rect 17859 4193 17871 5307
rect 17883 4889 17895 7251
rect 17907 2657 17919 7251
rect 17931 5105 17943 7251
rect 17883 1817 17895 2643
rect 17979 1865 17991 7251
rect 18027 6833 18039 7251
rect 18099 3977 18111 7251
rect 18123 4481 18135 7251
rect 18147 5921 18159 7251
rect 18171 4193 18183 7179
rect 18195 6953 18207 7251
rect 18123 1817 18135 4179
rect 18195 1817 18207 5331
rect 18243 4649 18255 7251
rect 18219 1817 18231 3771
rect 18243 1817 18255 4155
rect 18267 1817 18279 4395
rect 18315 3425 18327 7251
rect 18363 1841 18375 7251
rect 18435 5921 18447 7251
rect 18483 5777 18495 7251
rect 18555 2465 18567 7251
rect 18579 5441 18591 7251
rect 18603 6521 18615 7251
rect 18627 5465 18639 7251
rect 18699 4769 18711 7251
rect 18723 6497 18735 7251
rect 18771 6713 18783 7251
rect 18819 5153 18831 7251
rect 18867 5801 18879 7251
rect 18939 5825 18951 7251
rect 18963 4169 18975 7251
rect 18987 1817 18999 5811
rect 19011 3881 19023 7251
rect 19059 4121 19071 7251
rect 19083 5945 19095 7251
rect 19107 5105 19119 7251
rect 19155 4193 19167 7251
rect 19203 4433 19215 7251
rect 19227 4457 19239 7251
rect 19251 5561 19263 7251
rect 19059 1817 19071 1947
rect 19107 1817 19119 4179
rect 19203 1817 19215 4179
rect 19251 1817 19263 4827
rect 19275 2513 19287 7251
rect 19299 1817 19311 4923
rect 19323 3521 19335 7251
rect 19347 3569 19359 7251
rect 19371 4769 19383 7251
rect 19383 3425 19395 4587
rect 19323 1817 19335 3411
rect 19419 1961 19431 7251
rect 19443 1817 19455 3531
rect 19467 2297 19479 7251
rect 19491 3161 19503 7251
rect 19515 3137 19527 7251
rect 19539 5753 19551 7251
rect 19491 1817 19503 2115
rect 19563 1817 19575 3435
rect 19587 3185 19599 7251
rect 19611 3881 19623 7251
rect 19635 5681 19647 7251
rect 19659 5465 19671 7251
rect 19635 1817 19647 5187
rect 19683 1817 19695 4443
rect 19707 3977 19719 7251
rect 19731 5801 19743 7251
rect 19755 5201 19767 7251
rect 19755 1817 19767 4923
rect 19779 4601 19791 7251
rect 19827 6761 19839 7251
rect 19803 4193 19815 6075
rect 19827 1817 19839 6459
rect 19875 5321 19887 7251
rect 19851 1817 19863 3795
rect 19875 1817 19887 4995
rect 19899 3785 19911 5187
rect 19947 5153 19959 7251
rect 19923 1817 19935 3267
rect 19947 1817 19959 4179
rect 19971 2465 19983 7251
rect 19995 3569 20007 5307
rect 20019 4769 20031 7251
rect 20067 4697 20079 7251
rect 19971 1817 19983 2403
rect 20019 1817 20031 4611
rect 20091 4265 20103 7251
rect 20115 4745 20127 7251
rect 20139 6377 20151 7251
rect 20043 1817 20055 3915
rect 20115 1817 20127 3771
rect 20139 1817 20151 5667
rect 20163 1817 20175 5019
rect 20187 4025 20199 7251
rect 20211 4841 20223 7251
rect 20211 1817 20223 4011
rect 20235 3593 20247 7251
rect 20235 1817 20247 3243
rect 20259 2321 20271 7251
rect 20295 4193 20307 7155
rect 20331 6497 20343 7251
rect 20283 1817 20295 3939
rect 20331 1817 20343 6411
rect 20355 5009 20367 7251
rect 20355 1817 20367 4419
rect 20379 4217 20391 7251
rect 20427 5825 20439 7251
rect 20403 1817 20415 4251
rect 20451 4169 20463 7251
rect 20451 1817 20463 4011
rect 20499 3617 20511 7251
rect 20523 2777 20535 4755
rect 20547 4265 20559 7251
rect 20595 4577 20607 7251
rect 20475 1817 20487 2163
rect 20619 2033 20631 7251
rect 20643 5369 20655 7251
rect 20691 4769 20703 7251
rect 20571 1817 20583 2019
rect 20619 1817 20631 1947
rect 20667 1817 20679 4251
rect 20703 4025 20715 4659
rect 20739 3713 20751 7251
rect 20763 4169 20775 7251
rect 20787 5057 20799 7251
rect 20835 4937 20847 7251
rect 20703 1961 20715 2667
rect 20739 1817 20751 2859
rect 20799 2465 20811 4827
rect 20859 3761 20871 7251
rect 20787 1817 20799 1875
rect 20859 1817 20871 3699
rect 20883 3113 20895 7251
rect 20907 1817 20919 4587
rect 20931 4265 20943 7251
rect 20955 1817 20967 4755
rect 20979 4481 20991 7251
rect 21003 4409 21015 7251
rect 21003 1817 21015 2427
rect 21027 1817 21039 5763
rect 21051 5561 21063 7251
rect 21099 6329 21111 7251
rect 21051 1817 21063 4467
rect 21075 3785 21087 6291
rect 21123 5465 21135 7251
rect 21099 1817 21111 3483
rect 21123 1817 21135 3915
rect 21147 1817 21159 5139
rect 21171 4337 21183 7251
rect 21195 1817 21207 5259
rect 21219 4169 21231 7251
rect 21243 3809 21255 7251
rect 21291 6737 21303 7251
rect 21243 1817 21255 2835
rect 21267 2345 21279 4995
rect 21315 4481 21327 6891
rect 21339 4721 21351 7251
rect 21339 1817 21351 4251
rect 21363 2345 21375 7251
rect 21387 2801 21399 7251
rect 21411 4265 21423 5883
rect 21435 3185 21447 7251
rect 21459 4937 21471 7251
rect 21483 4241 21495 7251
rect 21387 1817 21399 2763
rect 21459 1817 21471 3315
rect 21483 1817 21495 4203
rect 21507 2777 21519 6987
rect 21531 4217 21543 5907
rect 21555 1817 21567 6267
rect 21603 5129 21615 7251
rect 21627 4481 21639 6219
rect 21603 1817 21615 4467
rect 21675 1817 21687 5619
rect 21723 1817 21735 4467
rect 21771 1817 21783 4251
rect 21819 1817 21831 6291
rect 21843 1817 21855 5763
rect 21867 1817 21879 3819
rect 21915 1817 21927 4467
rect 21963 2369 21975 7251
rect 21963 1817 21975 2283
rect 21987 1817 21999 4227
rect 22011 2297 22023 6363
rect 22155 4265 22167 7251
rect 22203 6233 22215 7251
rect 22035 1817 22047 2379
rect 22083 1817 22095 4203
rect 22131 1817 22143 2331
rect 22155 1817 22167 4155
rect 22203 1817 22215 6123
rect 22227 2705 22239 7251
rect 22251 7097 22263 7251
rect 22251 1817 22263 5547
rect 22299 4721 22311 7251
rect 22323 6473 22335 7251
rect 22347 7049 22359 7251
rect 22275 1817 22287 4155
rect 22299 1817 22311 4251
rect 22323 1817 22335 5595
rect 22347 1817 22359 5379
rect 22371 2849 22383 6219
rect 22395 4721 22407 7251
rect 22443 4889 22455 7251
rect 22395 1817 22407 4683
rect 22419 1817 22431 4731
rect 22455 4241 22467 4707
rect 22491 4601 22503 7251
rect 22443 1817 22455 4035
rect 22491 1817 22503 3291
rect 22515 1817 22527 5643
rect 22539 4265 22551 5403
rect 22563 3737 22575 7251
rect 22563 1817 22575 3579
rect 22587 2945 22599 7251
rect 22611 2825 22623 7251
rect 22611 1817 22623 2787
rect 22659 2585 22671 7251
rect 22683 4385 22695 7251
rect 22707 5177 22719 7251
rect 22755 6209 22767 7251
rect 22779 6761 22791 7251
rect 22803 6089 22815 7251
rect 22635 1817 22647 1899
rect 22707 1817 22719 3675
rect 22731 2057 22743 4587
rect 22755 1817 22767 4371
rect 22803 1817 22815 6051
rect 22827 3593 22839 6003
rect 22851 4601 22863 7251
rect 22851 1817 22863 4251
rect 22875 2993 22887 7251
rect 22923 5729 22935 7251
rect 22899 1817 22911 3867
rect 22923 1817 22935 5667
rect 22947 1817 22959 4227
rect 22971 2609 22983 7251
rect 22995 3209 23007 7251
rect 23019 4409 23031 7251
rect 23043 4673 23055 7251
rect 23091 5081 23103 7251
rect 23115 4721 23127 7251
rect 23187 6593 23199 7251
rect 23151 4385 23163 6555
rect 23019 1817 23031 2211
rect 23043 1817 23055 2307
rect 23067 1817 23079 4179
rect 23211 4169 23223 7251
rect 23235 5489 23247 7251
rect 23115 1817 23127 4107
rect 23139 1817 23151 3243
rect 23187 1817 23199 3483
rect 23247 2249 23259 4707
rect 23283 4361 23295 7251
rect 23307 3353 23319 6075
rect 23331 3929 23343 7251
rect 23283 1817 23295 2187
rect 23355 1817 23367 2811
rect 23379 1817 23391 4947
rect 23403 4193 23415 7251
rect 23451 6665 23463 7251
rect 23475 5705 23487 7251
rect 23499 6449 23511 7251
rect 23403 1817 23415 4107
rect 23547 3377 23559 7251
rect 23571 4865 23583 7251
rect 23451 1817 23463 2883
rect 23475 1817 23487 2331
rect 23547 1817 23559 2307
rect 23595 1817 23607 7131
rect 23619 4601 23631 7251
rect 23667 4841 23679 7251
rect 23691 4985 23703 7251
rect 23715 6785 23727 7251
rect 23667 1817 23679 4803
rect 23691 1817 23703 2547
rect 23715 1817 23727 6483
rect 23763 5225 23775 7251
rect 23739 2441 23751 4827
rect 23763 1817 23775 4371
rect 23787 4145 23799 7251
rect 23787 1817 23799 4035
rect 23811 1817 23823 4899
rect 23835 1865 23847 7251
rect 23859 1817 23871 6531
rect 23883 4673 23895 7251
rect 23907 5921 23919 7251
rect 23931 5969 23943 7251
rect 23979 6977 23991 7251
rect 23883 1817 23895 2427
rect 23907 1817 23919 4395
rect 23943 4385 23955 5811
rect 24003 4601 24015 7251
rect 24051 4433 24063 7251
rect 23931 1817 23943 3075
rect 23979 1817 23991 4131
rect 24003 1817 24015 4395
rect 24027 1817 24039 4371
rect 24075 1817 24087 3795
rect 24099 2681 24111 7251
rect 24123 4673 24135 7251
rect 24123 1817 24135 4419
rect 24147 4049 24159 7107
rect 24171 1817 24183 5475
rect 24195 2537 24207 7251
rect 24219 1817 24231 4323
rect 24243 3905 24255 7251
rect 24315 4721 24327 7251
rect 24267 1817 24279 4179
rect 24291 1913 24303 4587
rect 24315 1817 24327 4083
rect 24339 3617 24351 7251
rect 24363 5681 24375 7251
rect 24387 2081 24399 7251
rect 24435 4601 24447 7251
rect 24339 1817 24351 1899
rect 24411 1817 24423 2331
rect 24435 1817 24447 4515
rect 24459 3065 24471 7251
rect 24483 2345 24495 4707
rect 24507 4481 24519 7251
rect 24555 4073 24567 7251
rect 24579 4361 24591 7251
rect 24603 4337 24615 4587
rect 24531 1817 24543 3795
rect 24627 3473 24639 7251
rect 24675 7073 24687 7251
rect 24723 2969 24735 7251
rect 24795 4193 24807 7251
rect 24843 4121 24855 7251
rect 24867 6041 24879 7251
rect 24891 4457 24903 7251
rect 24915 5105 24927 7251
rect 24939 3233 24951 7251
rect 24987 4577 24999 7251
rect 25011 3281 25023 7251
rect 25035 5705 25047 7251
rect 25035 1817 25047 5667
rect 25083 4241 25095 7251
rect 25107 4697 25119 7251
rect 25131 4793 25143 7251
rect 25179 4697 25191 7251
rect 25203 6473 25215 7251
rect 25227 6209 25239 7251
rect 25083 1817 25095 3147
rect 25227 1817 25239 5931
rect 25275 2729 25287 7251
rect 25299 5537 25311 7251
rect 25347 6257 25359 7251
rect 25395 4625 25407 7251
rect 25419 5657 25431 7251
rect 25443 4673 25455 7251
rect 25491 3377 25503 7251
rect 25515 2705 25527 7251
rect 25539 4505 25551 7251
rect 25587 3401 25599 7251
rect 25611 4385 25623 7251
rect 25659 6113 25671 7251
rect 25707 2921 25719 7251
rect 25731 4649 25743 7251
rect 25755 4289 25767 7251
rect 25827 5297 25839 7251
rect 25779 1817 25791 4731
rect 25827 1817 25839 4515
rect 25851 3257 25863 7251
rect 25875 4529 25887 6459
rect 25899 2153 25911 7251
rect 25947 3809 25959 7251
rect 25971 1889 25983 7251
rect 25995 3017 26007 7251
rect 26019 1865 26031 5691
rect 26043 2849 26055 7251
rect 26067 5249 26079 7251
rect 25971 1817 25983 1851
rect 26091 1817 26103 4515
rect 26115 2801 26127 7251
rect 26163 4577 26175 7251
rect 26187 4217 26199 7251
rect 26211 6161 26223 7251
rect 26163 1817 26175 3651
rect 26187 1817 26199 2739
rect 26235 1817 26247 7011
rect 26259 4265 26271 7251
rect 26283 2417 26295 7251
rect 26307 2801 26319 7251
rect 26331 5825 26343 7251
rect 26259 1817 26271 1899
rect 26331 1817 26343 5787
rect 26355 1817 26367 3963
rect 26379 2417 26391 7251
rect 26403 4265 26415 7251
rect 26427 6209 26439 7251
rect 26427 1817 26439 6171
rect 26451 3161 26463 4563
rect 26475 3953 26487 7251
rect 26499 4409 26511 7251
rect 26523 6401 26535 7251
rect 26571 5873 26583 7251
rect 26535 4529 26547 5811
rect 26475 1817 26487 3915
rect 26499 1817 26511 4371
rect 26523 1817 26535 4491
rect 26571 1817 26583 3987
rect 26595 3881 26607 7251
rect 26619 2009 26631 7251
rect 26643 4433 26655 7251
rect 26667 3041 26679 7251
rect 26691 2105 26703 6195
rect 26715 4313 26727 7251
rect 26739 5777 26751 7251
rect 26763 6929 26775 7251
rect 26775 3929 26787 6603
rect 26811 5993 26823 7251
rect 26835 3497 26847 7251
rect 26859 4553 26871 7251
rect 26883 3713 26895 7251
rect 26907 4385 26919 5835
rect 26931 4937 26943 7251
rect 26955 4169 26967 7251
rect 26979 6353 26991 7251
rect 27003 4505 27015 7203
rect 27027 5513 27039 7251
rect 27027 1841 27039 1971
rect 27051 1865 27063 3627
rect 27075 1889 27087 3843
rect 27170 1817 27370 7251
rect 27459 1924 27529 1936
rect 27459 1876 27529 1888
rect 27459 1852 27529 1864
rect 27459 1828 27529 1840
rect 0 107 70 119
rect 0 83 70 95
rect 123 0 323 1018
rect 339 0 351 1018
rect 363 0 375 1018
rect 387 0 399 1018
rect 411 0 423 1018
rect 1659 144 1671 1018
rect 1779 168 1791 1018
rect 2499 192 2511 1018
rect 3531 72 3543 1018
rect 3555 216 3567 1018
rect 3627 240 3639 1018
rect 3675 264 3687 1018
rect 3891 288 3903 1018
rect 4299 48 4311 1018
rect 4323 312 4335 1018
rect 4371 336 4383 1018
rect 4539 360 4551 1018
rect 4755 384 4767 1018
rect 4779 408 4791 1018
rect 4803 288 4815 1018
rect 4827 168 4839 1018
rect 4947 288 4959 1018
rect 5307 168 5319 1018
rect 5499 432 5511 1018
rect 5643 456 5655 1018
rect 5739 480 5751 1018
rect 5955 504 5967 1018
rect 6243 528 6255 1018
rect 6315 552 6327 1018
rect 6387 576 6399 1018
rect 6411 216 6423 1018
rect 6531 216 6543 1018
rect 6579 600 6591 1018
rect 6627 408 6639 1018
rect 6819 408 6831 1018
rect 7227 624 7239 1018
rect 7563 648 7575 1018
rect 7755 672 7767 1018
rect 8259 720 8271 1018
rect 8427 744 8439 1018
rect 8763 768 8775 1018
rect 9051 792 9063 1018
rect 9339 816 9351 1018
rect 9411 840 9423 1018
rect 7935 0 7947 682
rect 9483 144 9495 1018
rect 9699 696 9711 1018
rect 9867 696 9879 1018
rect 9891 840 9903 1018
rect 10107 840 10119 1018
rect 10323 336 10335 1018
rect 10539 144 10551 1018
rect 10635 864 10647 1018
rect 10707 336 10719 1018
rect 10755 336 10767 1018
rect 10827 888 10839 1018
rect 10947 912 10959 1018
rect 11043 936 11055 1018
rect 11259 648 11271 1018
rect 12267 144 12279 1018
rect 12315 240 12327 1018
rect 12363 648 12375 1018
rect 12411 360 12423 1018
rect 12531 360 12543 1018
rect 12843 768 12855 1018
rect 12987 768 12999 1018
rect 13131 576 13143 1018
rect 13323 720 13335 1018
rect 13395 576 13407 1018
rect 13563 816 13575 1018
rect 13611 768 13623 1018
rect 13683 576 13695 1018
rect 13731 720 13743 1018
rect 13947 768 13959 1018
rect 14379 384 14391 1018
rect 14427 816 14439 1018
rect 14475 648 14487 1018
rect 14523 648 14535 1018
rect 14571 576 14583 1018
rect 14691 360 14703 1018
rect 14859 576 14871 1018
rect 14907 384 14919 1018
rect 15099 864 15111 1018
rect 15147 360 15159 1018
rect 14307 0 14319 226
rect 15267 144 15279 1018
rect 15963 864 15975 1018
rect 16011 864 16023 1018
rect 16131 48 16143 1018
rect 16227 888 16239 1018
rect 16323 48 16335 1018
rect 16467 888 16479 1018
rect 16683 528 16695 1018
rect 17259 528 17271 1018
rect 17283 48 17295 1018
rect 17571 960 17583 1018
rect 17811 360 17823 1018
rect 14331 0 14343 34
rect 17883 24 17895 1018
rect 17931 96 17943 1018
rect 17979 96 17991 1018
rect 18051 984 18063 1018
rect 18075 1008 18087 1018
rect 18099 912 18111 1018
rect 18147 960 18159 1018
rect 18291 1008 18303 1018
rect 18411 96 18423 1018
rect 18819 144 18831 1018
rect 18963 936 18975 1018
rect 19011 912 19023 1018
rect 19179 624 19191 1018
rect 19347 792 19359 1018
rect 19395 864 19407 1018
rect 19419 264 19431 1018
rect 19467 624 19479 1018
rect 19539 768 19551 1018
rect 19587 576 19599 1018
rect 19659 648 19671 1018
rect 19731 576 19743 1018
rect 19779 600 19791 1018
rect 20067 624 20079 1018
rect 20523 576 20535 1018
rect 20571 576 20583 1018
rect 20883 192 20895 1018
rect 20931 480 20943 1018
rect 21315 456 21327 1018
rect 21363 600 21375 1018
rect 21411 624 21423 1018
rect 21507 696 21519 1018
rect 21579 696 21591 1018
rect 21627 120 21639 1018
rect 21699 384 21711 1018
rect 21747 888 21759 1018
rect 21939 840 21951 1018
rect 22059 216 22071 1018
rect 22659 432 22671 1018
rect 22731 240 22743 1018
rect 22827 168 22839 1018
rect 22995 768 23007 1018
rect 23235 216 23247 1018
rect 23499 600 23511 1018
rect 24099 720 24111 1018
rect 24195 504 24207 1018
rect 24243 360 24255 1018
rect 24363 648 24375 1018
rect 24459 816 24471 1018
rect 24507 336 24519 1018
rect 24555 696 24567 1018
rect 24675 408 24687 1018
rect 25275 984 25287 1018
rect 25419 624 25431 1018
rect 20691 0 20703 58
rect 25995 48 26007 1018
rect 26019 312 26031 1018
rect 26043 288 26055 1018
rect 26115 744 26127 1018
rect 26139 552 26151 1018
rect 26283 768 26295 1018
rect 26379 672 26391 1018
rect 26451 912 26463 1018
rect 26571 72 26583 1018
rect 26571 24 26583 34
rect 26595 24 26607 562
rect 27171 0 27371 1018
rect 27459 515 27529 527
rect 27459 59 27529 71
rect 27459 35 27529 47
rect 27459 11 27529 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7251
box 0 0 1464 799
use nand3 g8043
timestamp 1396952988
transform 1 0 1587 0 1 7251
box 0 0 120 799
use rowcrosser PcEn
timestamp 1397224710
transform 1 0 1707 0 1 7251
box 0 0 48 799
use nand3 g8112
timestamp 1396952988
transform 1 0 1755 0 1 7251
box 0 0 120 799
use nand2 g8291
timestamp 1386234792
transform 1 0 1875 0 1 7251
box 0 0 96 799
use inv g7923
timestamp 1386238110
transform 1 0 1971 0 1 7251
box 0 0 120 799
use nand2 g8060
timestamp 1386234792
transform 1 0 2091 0 1 7251
box 0 0 96 799
use and2 g7942
timestamp 1386234845
transform 1 0 2187 0 1 7251
box 0 0 120 799
use nand3 g8182
timestamp 1396952988
transform 1 0 2307 0 1 7251
box 0 0 120 799
use nand3 g8066
timestamp 1396952988
transform 1 0 2427 0 1 7251
box 0 0 120 799
use nand2 g8169
timestamp 1386234792
transform 1 0 2547 0 1 7251
box 0 0 96 799
use nand2 g7934
timestamp 1386234792
transform 1 0 2643 0 1 7251
box 0 0 96 799
use nand2 g8107
timestamp 1386234792
transform 1 0 2739 0 1 7251
box 0 0 96 799
use nand3 g8229
timestamp 1396952988
transform 1 0 2835 0 1 7251
box 0 0 120 799
use nand2 g8039
timestamp 1386234792
transform 1 0 2955 0 1 7251
box 0 0 96 799
use nand2 g7912
timestamp 1386234792
transform 1 0 3051 0 1 7251
box 0 0 96 799
use nand3 g8046
timestamp 1396952988
transform 1 0 3147 0 1 7251
box 0 0 120 799
use nor2 g8123
timestamp 1386235306
transform 1 0 3267 0 1 7251
box 0 0 120 799
use nand3 g8222
timestamp 1396952988
transform 1 0 3387 0 1 7251
box 0 0 120 799
use nand3 g8098
timestamp 1396952988
transform 1 0 3507 0 1 7251
box 0 0 120 799
use nand2 g8102
timestamp 1386234792
transform 1 0 3627 0 1 7251
box 0 0 96 799
use nand3 g8012
timestamp 1396952988
transform 1 0 3723 0 1 7251
box 0 0 120 799
use and2 g8187
timestamp 1386234845
transform 1 0 3843 0 1 7251
box 0 0 120 799
use and2 g7951
timestamp 1386234845
transform 1 0 3963 0 1 7251
box 0 0 120 799
use nand4 g8135
timestamp 1386234936
transform 1 0 4083 0 1 7251
box 0 0 144 799
use nand2 g8171
timestamp 1386234792
transform 1 0 4227 0 1 7251
box 0 0 96 799
use and2 g8154
timestamp 1386234845
transform 1 0 4323 0 1 7251
box 0 0 120 799
use and2 g8276
timestamp 1386234845
transform 1 0 4443 0 1 7251
box 0 0 120 799
use inv g8261
timestamp 1386238110
transform 1 0 4563 0 1 7251
box 0 0 120 799
use nor2 g8130
timestamp 1386235306
transform 1 0 4683 0 1 7251
box 0 0 120 799
use nand2 g8027
timestamp 1386234792
transform 1 0 4803 0 1 7251
box 0 0 96 799
use nor2 g8082
timestamp 1386235306
transform 1 0 4899 0 1 7251
box 0 0 120 799
use nand2 g8035
timestamp 1386234792
transform 1 0 5019 0 1 7251
box 0 0 96 799
use nand2 g8019
timestamp 1386234792
transform 1 0 5115 0 1 7251
box 0 0 96 799
use nand2 g8168
timestamp 1386234792
transform 1 0 5211 0 1 7251
box 0 0 96 799
use and2 g8238
timestamp 1386234845
transform 1 0 5307 0 1 7251
box 0 0 120 799
use nand2 g7989
timestamp 1386234792
transform 1 0 5427 0 1 7251
box 0 0 96 799
use and2 g8225
timestamp 1386234845
transform 1 0 5523 0 1 7251
box 0 0 120 799
use nand2 g8143
timestamp 1386234792
transform 1 0 5643 0 1 7251
box 0 0 96 799
use nand2 g8069
timestamp 1386234792
transform 1 0 5739 0 1 7251
box 0 0 96 799
use nand2 g8042
timestamp 1386234792
transform 1 0 5835 0 1 7251
box 0 0 96 799
use nand2 g8149
timestamp 1386234792
transform 1 0 5931 0 1 7251
box 0 0 96 799
use nand2 g7926
timestamp 1386234792
transform 1 0 6027 0 1 7251
box 0 0 96 799
use nand2 g8280
timestamp 1386234792
transform 1 0 6123 0 1 7251
box 0 0 96 799
use nand2 g7985
timestamp 1386234792
transform 1 0 6219 0 1 7251
box 0 0 96 799
use nand2 g8249
timestamp 1386234792
transform 1 0 6315 0 1 7251
box 0 0 96 799
use inv g8064
timestamp 1386238110
transform 1 0 6411 0 1 7251
box 0 0 120 799
use nand2 g8235
timestamp 1386234792
transform 1 0 6531 0 1 7251
box 0 0 96 799
use nand2 g7948
timestamp 1386234792
transform 1 0 6627 0 1 7251
box 0 0 96 799
use nand2 g8058
timestamp 1386234792
transform 1 0 6723 0 1 7251
box 0 0 96 799
use nand2 g8009
timestamp 1386234792
transform 1 0 6819 0 1 7251
box 0 0 96 799
use nand2 g8055
timestamp 1386234792
transform 1 0 6915 0 1 7251
box 0 0 96 799
use nand2 g7939
timestamp 1386234792
transform 1 0 7011 0 1 7251
box 0 0 96 799
use nand3 g8088
timestamp 1396952988
transform 1 0 7107 0 1 7251
box 0 0 120 799
use nand2 g7947
timestamp 1386234792
transform 1 0 7227 0 1 7251
box 0 0 96 799
use nand4 g7960
timestamp 1386234936
transform 1 0 7323 0 1 7251
box 0 0 144 799
use nand3 g8214
timestamp 1396952988
transform 1 0 7467 0 1 7251
box 0 0 120 799
use inv g8056
timestamp 1386238110
transform 1 0 7587 0 1 7251
box 0 0 120 799
use nand2 g8281
timestamp 1386234792
transform 1 0 7707 0 1 7251
box 0 0 96 799
use inv g8269
timestamp 1386238110
transform 1 0 7803 0 1 7251
box 0 0 120 799
use and2 g8183
timestamp 1386234845
transform 1 0 7923 0 1 7251
box 0 0 120 799
use nand2 g8170
timestamp 1386234792
transform 1 0 8043 0 1 7251
box 0 0 96 799
use nand2 g8124
timestamp 1386234792
transform 1 0 8139 0 1 7251
box 0 0 96 799
use and2 g8106
timestamp 1386234845
transform 1 0 8235 0 1 7251
box 0 0 120 799
use and2 g8119
timestamp 1386234845
transform 1 0 8355 0 1 7251
box 0 0 120 799
use nand3 g8275
timestamp 1396952988
transform 1 0 8475 0 1 7251
box 0 0 120 799
use nand2 g8146
timestamp 1386234792
transform 1 0 8595 0 1 7251
box 0 0 96 799
use nand2 g8127
timestamp 1386234792
transform 1 0 8691 0 1 7251
box 0 0 96 799
use nand4 g8155
timestamp 1386234936
transform 1 0 8787 0 1 7251
box 0 0 144 799
use nand3 g8033
timestamp 1396952988
transform 1 0 8931 0 1 7251
box 0 0 120 799
use and2 g7921
timestamp 1386234845
transform 1 0 9051 0 1 7251
box 0 0 120 799
use nor2 g8252
timestamp 1386235306
transform 1 0 9171 0 1 7251
box 0 0 120 799
use nand2 g7978
timestamp 1386234792
transform 1 0 9291 0 1 7251
box 0 0 96 799
use nand2 g8244
timestamp 1386234792
transform 1 0 9387 0 1 7251
box 0 0 96 799
use nor2 g7930
timestamp 1386235306
transform 1 0 9483 0 1 7251
box 0 0 120 799
use nor2 g7972
timestamp 1386235306
transform 1 0 9603 0 1 7251
box 0 0 120 799
use nand2 g8240
timestamp 1386234792
transform 1 0 9723 0 1 7251
box 0 0 96 799
use mux2 g8054
timestamp 1386235218
transform 1 0 9819 0 1 7251
box 0 0 192 799
use nand2 g8139
timestamp 1386234792
transform 1 0 10011 0 1 7251
box 0 0 96 799
use inv g8023
timestamp 1386238110
transform 1 0 10107 0 1 7251
box 0 0 120 799
use inv g8118
timestamp 1386238110
transform 1 0 10227 0 1 7251
box 0 0 120 799
use nand3 g7981
timestamp 1396952988
transform 1 0 10347 0 1 7251
box 0 0 120 799
use nand2 g8111
timestamp 1386234792
transform 1 0 10467 0 1 7251
box 0 0 96 799
use inv g8120
timestamp 1386238110
transform 1 0 10563 0 1 7251
box 0 0 120 799
use inv g8091
timestamp 1386238110
transform 1 0 10683 0 1 7251
box 0 0 120 799
use nand2 g8134
timestamp 1386234792
transform 1 0 10803 0 1 7251
box 0 0 96 799
use nand3 g8050
timestamp 1396952988
transform 1 0 10899 0 1 7251
box 0 0 120 799
use nand2 g8218
timestamp 1386234792
transform 1 0 11019 0 1 7251
box 0 0 96 799
use nand2 g7995
timestamp 1386234792
transform 1 0 11115 0 1 7251
box 0 0 96 799
use nand3 g7945
timestamp 1396952988
transform 1 0 11211 0 1 7251
box 0 0 120 799
use nand4 g8284
timestamp 1386234936
transform 1 0 11331 0 1 7251
box 0 0 144 799
use nand2 g7964
timestamp 1386234792
transform 1 0 11475 0 1 7251
box 0 0 96 799
use nand4 g8198
timestamp 1386234936
transform 1 0 11571 0 1 7251
box 0 0 144 799
use nand2 g8272
timestamp 1386234792
transform 1 0 11715 0 1 7251
box 0 0 96 799
use inv g8199
timestamp 1386238110
transform 1 0 11811 0 1 7251
box 0 0 120 799
use nor2 g8221
timestamp 1386235306
transform 1 0 11931 0 1 7251
box 0 0 120 799
use xor2 g8220
timestamp 1396952988
transform 1 0 12051 0 1 7251
box 0 0 192 799
use nand2 g8194
timestamp 1386234792
transform 1 0 12243 0 1 7251
box 0 0 96 799
use inv g8230
timestamp 1386238110
transform 1 0 12339 0 1 7251
box 0 0 120 799
use and2 g8271
timestamp 1386234845
transform 1 0 12459 0 1 7251
box 0 0 120 799
use nand2 g8004
timestamp 1386234792
transform 1 0 12579 0 1 7251
box 0 0 96 799
use and2 rm_assigns_buf_StatusReg_1
timestamp 1386234845
transform 1 0 12675 0 1 7251
box 0 0 120 799
use buffer g8074
timestamp 1386236986
transform 1 0 12795 0 1 7251
box 0 0 120 799
use nand3 g8209
timestamp 1396952988
transform 1 0 12915 0 1 7251
box 0 0 120 799
use nand2 g8103
timestamp 1386234792
transform 1 0 13035 0 1 7251
box 0 0 96 799
use and2 g8268
timestamp 1386234845
transform 1 0 13131 0 1 7251
box 0 0 120 799
use nand2 g8283
timestamp 1386234792
transform 1 0 13251 0 1 7251
box 0 0 96 799
use inv g8180
timestamp 1386238110
transform 1 0 13347 0 1 7251
box 0 0 120 799
use nand2 g8005
timestamp 1386234792
transform 1 0 13467 0 1 7251
box 0 0 96 799
use nand3 g8052
timestamp 1396952988
transform 1 0 13563 0 1 7251
box 0 0 120 799
use nand2 g8136
timestamp 1386234792
transform 1 0 13683 0 1 7251
box 0 0 96 799
use rowcrosser Op1Sel
timestamp 1397224710
transform 1 0 13779 0 1 7251
box 0 0 48 799
use nand2 g8110
timestamp 1386234792
transform 1 0 13827 0 1 7251
box 0 0 96 799
use nand2 g8153
timestamp 1386234792
transform 1 0 13923 0 1 7251
box 0 0 96 799
use nand4 StatusReg_reg_91_3_93_
timestamp 1386234936
transform 1 0 14019 0 1 7251
box 0 0 144 799
use scandtype g7922
timestamp 1386241841
transform 1 0 14163 0 1 7251
box 0 0 624 799
use nand4 stateSub_reg_91_2_93_
timestamp 1386234936
transform 1 0 14787 0 1 7251
box 0 0 144 799
use scandtype g8294
timestamp 1386241841
transform 1 0 14931 0 1 7251
box 0 0 624 799
use inv g8024
timestamp 1386238110
transform 1 0 15555 0 1 7251
box 0 0 120 799
use rowcrosser rowcrosser_0
timestamp 1397224710
transform 1 0 15675 0 1 7251
box 0 0 48 799
use nand3 g8099
timestamp 1396952988
transform 1 0 15723 0 1 7251
box 0 0 120 799
use nand3 g8057
timestamp 1396952988
transform 1 0 15843 0 1 7251
box 0 0 120 799
use nand2 g8190
timestamp 1386234792
transform 1 0 15963 0 1 7251
box 0 0 96 799
use inv g8045
timestamp 1386238110
transform 1 0 16059 0 1 7251
box 0 0 120 799
use inv g7913
timestamp 1386238110
transform 1 0 16179 0 1 7251
box 0 0 120 799
use nand3 g8018
timestamp 1396952988
transform 1 0 16299 0 1 7251
box 0 0 120 799
use nand3 g8092
timestamp 1396952988
transform 1 0 16419 0 1 7251
box 0 0 120 799
use nand2 g8277
timestamp 1386234792
transform 1 0 16539 0 1 7251
box 0 0 96 799
use nand2 g8081
timestamp 1386234792
transform 1 0 16635 0 1 7251
box 0 0 96 799
use nand3 g8243
timestamp 1396952988
transform 1 0 16731 0 1 7251
box 0 0 120 799
use nor2 g8234
timestamp 1386235306
transform 1 0 16851 0 1 7251
box 0 0 120 799
use nand2 StatusReg_reg_91_1_93_
timestamp 1386234792
transform 1 0 16971 0 1 7251
box 0 0 96 799
use scandtype g8293
timestamp 1386241841
transform 1 0 17067 0 1 7251
box 0 0 624 799
use rowcrosser AluOR_91_0_93_
timestamp 1397224710
transform 1 0 17691 0 1 7251
box 0 0 48 799
use inv g7933
timestamp 1386238110
transform 1 0 17739 0 1 7251
box 0 0 120 799
use nand2 g8028
timestamp 1386234792
transform 1 0 17859 0 1 7251
box 0 0 96 799
use inv g8213
timestamp 1386238110
transform 1 0 17955 0 1 7251
box 0 0 120 799
use nand2 g7963
timestamp 1386234792
transform 1 0 18075 0 1 7251
box 0 0 96 799
use inv g8096
timestamp 1386238110
transform 1 0 18171 0 1 7251
box 0 0 120 799
use inv g8212
timestamp 1386238110
transform 1 0 18291 0 1 7251
box 0 0 120 799
use inv g7906
timestamp 1386238110
transform 1 0 18411 0 1 7251
box 0 0 120 799
use nand4 g8015
timestamp 1386234936
transform 1 0 18531 0 1 7251
box 0 0 144 799
use and2 g8084
timestamp 1386234845
transform 1 0 18675 0 1 7251
box 0 0 120 799
use inv g8265
timestamp 1386238110
transform 1 0 18795 0 1 7251
box 0 0 120 799
use and2 g8108
timestamp 1386234845
transform 1 0 18915 0 1 7251
box 0 0 120 799
use nand2 g8049
timestamp 1386234792
transform 1 0 19035 0 1 7251
box 0 0 96 799
use rowcrosser AluEn
timestamp 1397224710
transform 1 0 19131 0 1 7251
box 0 0 48 799
use nand3 g8144
timestamp 1396952988
transform 1 0 19179 0 1 7251
box 0 0 120 799
use nand2 g8159
timestamp 1386234792
transform 1 0 19299 0 1 7251
box 0 0 96 799
use rowcrosser PcSel_91_1_93_
timestamp 1397224710
transform 1 0 19395 0 1 7251
box 0 0 48 799
use nand3 g8177
timestamp 1396952988
transform 1 0 19443 0 1 7251
box 0 0 120 799
use nand3 g7996
timestamp 1396952988
transform 1 0 19563 0 1 7251
box 0 0 120 799
use nand3 g8251
timestamp 1396952988
transform 1 0 19683 0 1 7251
box 0 0 120 799
use inv g8036
timestamp 1386238110
transform 1 0 19803 0 1 7251
box 0 0 120 799
use and2 g8226
timestamp 1386234845
transform 1 0 19923 0 1 7251
box 0 0 120 799
use nand3 g7929
timestamp 1396952988
transform 1 0 20043 0 1 7251
box 0 0 120 799
use nand4 g7979
timestamp 1386234936
transform 1 0 20163 0 1 7251
box 0 0 144 799
use nand2 g8264
timestamp 1386234792
transform 1 0 20307 0 1 7251
box 0 0 96 799
use nor2 g7924
timestamp 1386235306
transform 1 0 20403 0 1 7251
box 0 0 120 799
use rowcrosser AluWe
timestamp 1397224710
transform 1 0 20523 0 1 7251
box 0 0 48 799
use nand2 g8089
timestamp 1386234792
transform 1 0 20571 0 1 7251
box 0 0 96 799
use rowcrosser LrSel
timestamp 1397224710
transform 1 0 20667 0 1 7251
box 0 0 48 799
use nand2 g8206
timestamp 1386234792
transform 1 0 20715 0 1 7251
box 0 0 96 799
use nand2 g8237
timestamp 1386234792
transform 1 0 20811 0 1 7251
box 0 0 96 799
use rowcrosser PcSel_91_2_93_
timestamp 1397224710
transform 1 0 20907 0 1 7251
box 0 0 48 799
use and2 g8016
timestamp 1386234845
transform 1 0 20955 0 1 7251
box 0 0 120 799
use and2 g8278
timestamp 1386234845
transform 1 0 21075 0 1 7251
box 0 0 120 799
use nor2 g8181
timestamp 1386235306
transform 1 0 21195 0 1 7251
box 0 0 120 799
use nand2 g8216
timestamp 1386234792
transform 1 0 21315 0 1 7251
box 0 0 96 799
use nand2 StatusReg_reg_91_0_93_
timestamp 1386234792
transform 1 0 21411 0 1 7251
box 0 0 96 799
use scandtype g8253
timestamp 1386241841
transform 1 0 21507 0 1 7251
box 0 0 624 799
use rowcrosser MemEn
timestamp 1397224710
transform 1 0 22131 0 1 7251
box 0 0 48 799
use nand2 g8186
timestamp 1386234792
transform 1 0 22179 0 1 7251
box 0 0 96 799
use nand2 g7946
timestamp 1386234792
transform 1 0 22275 0 1 7251
box 0 0 96 799
use rowcrosser nME
timestamp 1397224710
transform 1 0 22371 0 1 7251
box 0 0 48 799
use inv g8090
timestamp 1386238110
transform 1 0 22419 0 1 7251
box 0 0 120 799
use nand2 g8195
timestamp 1386234792
transform 1 0 22539 0 1 7251
box 0 0 96 799
use nand2 g8223
timestamp 1386234792
transform 1 0 22635 0 1 7251
box 0 0 96 799
use nand2 g8077
timestamp 1386234792
transform 1 0 22731 0 1 7251
box 0 0 96 799
use nor2 g8133
timestamp 1386235306
transform 1 0 22827 0 1 7251
box 0 0 120 799
use nand3 g7971
timestamp 1396952988
transform 1 0 22947 0 1 7251
box 0 0 120 799
use nand2 g8041
timestamp 1386234792
transform 1 0 23067 0 1 7251
box 0 0 96 799
use nand2 g8289
timestamp 1386234792
transform 1 0 23163 0 1 7251
box 0 0 96 799
use inv g8002
timestamp 1386238110
transform 1 0 23259 0 1 7251
box 0 0 120 799
use rowcrosser Op2Sel_91_0_93_
timestamp 1397224710
transform 1 0 23379 0 1 7251
box 0 0 48 799
use nand2 g8128
timestamp 1386234792
transform 1 0 23427 0 1 7251
box 0 0 96 799
use and2 g8100
timestamp 1386234845
transform 1 0 23523 0 1 7251
box 0 0 120 799
use nand2 g8029
timestamp 1386234792
transform 1 0 23643 0 1 7251
box 0 0 96 799
use nor2 g8117
timestamp 1386235306
transform 1 0 23739 0 1 7251
box 0 0 120 799
use nand2 g8167
timestamp 1386234792
transform 1 0 23859 0 1 7251
box 0 0 96 799
use and2 g7982
timestamp 1386234845
transform 1 0 23955 0 1 7251
box 0 0 120 799
use nand2 g8227
timestamp 1386234792
transform 1 0 24075 0 1 7251
box 0 0 96 799
use inv g8191
timestamp 1386238110
transform 1 0 24171 0 1 7251
box 0 0 120 799
use nand3 g7975
timestamp 1396952988
transform 1 0 24291 0 1 7251
box 0 0 120 799
use and2 g8270
timestamp 1386234845
transform 1 0 24411 0 1 7251
box 0 0 120 799
use and2 g8073
timestamp 1386234845
transform 1 0 24531 0 1 7251
box 0 0 120 799
use inv g7967
timestamp 1386238110
transform 1 0 24651 0 1 7251
box 0 0 120 799
use rowcrosser PcSel_91_0_93_
timestamp 1397224710
transform 1 0 24771 0 1 7251
box 0 0 48 799
use nand4 g7925
timestamp 1386234936
transform 1 0 24819 0 1 7251
box 0 0 144 799
use nand2 g8163
timestamp 1386234792
transform 1 0 24963 0 1 7251
box 0 0 96 799
use nand2 g8273
timestamp 1386234792
transform 1 0 25059 0 1 7251
box 0 0 96 799
use nand2 g7969
timestamp 1386234792
transform 1 0 25155 0 1 7251
box 0 0 96 799
use nor2 g8051
timestamp 1386235306
transform 1 0 25251 0 1 7251
box 0 0 120 799
use nand2 g8147
timestamp 1386234792
transform 1 0 25371 0 1 7251
box 0 0 96 799
use nand2 g7955
timestamp 1386234792
transform 1 0 25467 0 1 7251
box 0 0 96 799
use and2 g7928
timestamp 1386234845
transform 1 0 25563 0 1 7251
box 0 0 120 799
use nand3 g8030
timestamp 1396952988
transform 1 0 25683 0 1 7251
box 0 0 120 799
use nor2 g8217
timestamp 1386235306
transform 1 0 25803 0 1 7251
box 0 0 120 799
use nand2 g8248
timestamp 1386234792
transform 1 0 25923 0 1 7251
box 0 0 96 799
use and2 g8114
timestamp 1386234845
transform 1 0 26019 0 1 7251
box 0 0 120 799
use nand2 g8174
timestamp 1386234792
transform 1 0 26139 0 1 7251
box 0 0 96 799
use nand3 g8241
timestamp 1396952988
transform 1 0 26235 0 1 7251
box 0 0 120 799
use nand2 g8067
timestamp 1386234792
transform 1 0 26355 0 1 7251
box 0 0 96 799
use nand2 g7990
timestamp 1386234792
transform 1 0 26451 0 1 7251
box 0 0 96 799
use nand4 g8158
timestamp 1386234936
transform 1 0 26547 0 1 7251
box 0 0 144 799
use nand2 g8063
timestamp 1386234792
transform 1 0 26691 0 1 7251
box 0 0 96 799
use nand3 g8257
timestamp 1396952988
transform 1 0 26787 0 1 7251
box 0 0 120 799
use nand2 ENB
timestamp 1386234792
transform 1 0 26907 0 1 7251
box 0 0 96 799
use rowcrosser RwSel_91_1_93_
timestamp 1397224710
transform 1 0 27003 0 1 7251
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27051 0 1 7251
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 1018
box 0 0 1464 799
use nand2 stateSub_reg_91_0_93_
timestamp 1386234792
transform 1 0 1587 0 1 1018
box 0 0 96 799
use scandtype g8150
timestamp 1386241841
transform 1 0 1683 0 1 1018
box 0 0 624 799
use nand2 g8020
timestamp 1386234792
transform 1 0 2307 0 1 1018
box 0 0 96 799
use nand3 g8178
timestamp 1396952988
transform 1 0 2403 0 1 1018
box 0 0 120 799
use and2 state_reg_91_1_93_
timestamp 1386234845
transform 1 0 2523 0 1 1018
box 0 0 120 799
use scandtype g8250
timestamp 1386241841
transform 1 0 2643 0 1 1018
box 0 0 624 799
use nand2 g8148
timestamp 1386234792
transform 1 0 3267 0 1 1018
box 0 0 96 799
use inv g7976
timestamp 1386238110
transform 1 0 3363 0 1 1018
box 0 0 120 799
use nand2 g7993
timestamp 1386234792
transform 1 0 3483 0 1 1018
box 0 0 96 799
use nor2 g8196
timestamp 1386235306
transform 1 0 3579 0 1 1018
box 0 0 120 799
use nand3 g8211
timestamp 1396952988
transform 1 0 3699 0 1 1018
box 0 0 120 799
use nand2 g8175
timestamp 1386234792
transform 1 0 3819 0 1 1018
box 0 0 96 799
use nand2 g8078
timestamp 1386234792
transform 1 0 3915 0 1 1018
box 0 0 96 799
use inv g8093
timestamp 1386238110
transform 1 0 4011 0 1 1018
box 0 0 120 799
use and2 g7974
timestamp 1386234845
transform 1 0 4131 0 1 1018
box 0 0 120 799
use nand2 g8104
timestamp 1386234792
transform 1 0 4251 0 1 1018
box 0 0 96 799
use inv g7940
timestamp 1386238110
transform 1 0 4347 0 1 1018
box 0 0 120 799
use nand4 g8160
timestamp 1386234936
transform 1 0 4467 0 1 1018
box 0 0 144 799
use nor2 g8076
timestamp 1386235306
transform 1 0 4611 0 1 1018
box 0 0 120 799
use nand3 StatusReg_reg_91_2_93_
timestamp 1396952988
transform 1 0 4731 0 1 1018
box 0 0 120 799
use scandtype g8161
timestamp 1386241841
transform 1 0 4851 0 1 1018
box 0 0 624 799
use nand2 g8224
timestamp 1386234792
transform 1 0 5475 0 1 1018
box 0 0 96 799
use nand2 g8094
timestamp 1386234792
transform 1 0 5571 0 1 1018
box 0 0 96 799
use nand2 g8121
timestamp 1386234792
transform 1 0 5667 0 1 1018
box 0 0 96 799
use nand3 g8037
timestamp 1396952988
transform 1 0 5763 0 1 1018
box 0 0 120 799
use nand2 g8266
timestamp 1386234792
transform 1 0 5883 0 1 1018
box 0 0 96 799
use inv g8189
timestamp 1386238110
transform 1 0 5979 0 1 1018
box 0 0 120 799
use nand3 g8125
timestamp 1396952988
transform 1 0 6099 0 1 1018
box 0 0 120 799
use nor2 g7915
timestamp 1386235306
transform 1 0 6219 0 1 1018
box 0 0 120 799
use nand3 g8232
timestamp 1396952988
transform 1 0 6339 0 1 1018
box 0 0 120 799
use nand2 g8152
timestamp 1386234792
transform 1 0 6459 0 1 1018
box 0 0 96 799
use nand2 g8080
timestamp 1386234792
transform 1 0 6555 0 1 1018
box 0 0 96 799
use nand2 g7937
timestamp 1386234792
transform 1 0 6651 0 1 1018
box 0 0 96 799
use nand2 g7997
timestamp 1386234792
transform 1 0 6747 0 1 1018
box 0 0 96 799
use nor2 g8267
timestamp 1386235306
transform 1 0 6843 0 1 1018
box 0 0 120 799
use nand2 g8282
timestamp 1386234792
transform 1 0 6963 0 1 1018
box 0 0 96 799
use nand2 g8274
timestamp 1386234792
transform 1 0 7059 0 1 1018
box 0 0 96 799
use nand2 g8236
timestamp 1386234792
transform 1 0 7155 0 1 1018
box 0 0 96 799
use nor2 g8101
timestamp 1386235306
transform 1 0 7251 0 1 1018
box 0 0 120 799
use nor2 g8011
timestamp 1386235306
transform 1 0 7371 0 1 1018
box 0 0 120 799
use nand2 g8185
timestamp 1386234792
transform 1 0 7491 0 1 1018
box 0 0 96 799
use and2 g7927
timestamp 1386234845
transform 1 0 7587 0 1 1018
box 0 0 120 799
use and2 g8255
timestamp 1386234845
transform 1 0 7707 0 1 1018
box 0 0 120 799
use and2 g8086
timestamp 1386234845
transform 1 0 7827 0 1 1018
box 0 0 120 799
use and2 g8301
timestamp 1386234845
transform 1 0 7947 0 1 1018
box 0 0 120 799
use inv g7962
timestamp 1386238110
transform 1 0 8067 0 1 1018
box 0 0 120 799
use nand4 g8192
timestamp 1386234936
transform 1 0 8187 0 1 1018
box 0 0 144 799
use nand3 g7988
timestamp 1396952988
transform 1 0 8331 0 1 1018
box 0 0 120 799
use nand2 g8292
timestamp 1386234792
transform 1 0 8451 0 1 1018
box 0 0 96 799
use inv g8254
timestamp 1386238110
transform 1 0 8547 0 1 1018
box 0 0 120 799
use and2 g8116
timestamp 1386234845
transform 1 0 8667 0 1 1018
box 0 0 120 799
use and2 g8166
timestamp 1386234845
transform 1 0 8787 0 1 1018
box 0 0 120 799
use nand2 g8145
timestamp 1386234792
transform 1 0 8907 0 1 1018
box 0 0 96 799
use and2 g7907
timestamp 1386234845
transform 1 0 9003 0 1 1018
box 0 0 120 799
use nand4 g8001
timestamp 1386234936
transform 1 0 9123 0 1 1018
box 0 0 144 799
use nand2 g7959
timestamp 1386234792
transform 1 0 9267 0 1 1018
box 0 0 96 799
use nand2 g8014
timestamp 1386234792
transform 1 0 9363 0 1 1018
box 0 0 96 799
use nand2 g7998
timestamp 1386234792
transform 1 0 9459 0 1 1018
box 0 0 96 799
use nor2 g8228
timestamp 1386235306
transform 1 0 9555 0 1 1018
box 0 0 120 799
use rowcrosser Flags_91_0_93_
timestamp 1397224710
transform 1 0 9675 0 1 1018
box 0 0 48 799
use nand2 g7987
timestamp 1386234792
transform 1 0 9723 0 1 1018
box 0 0 96 799
use nand2 g8072
timestamp 1386234792
transform 1 0 9819 0 1 1018
box 0 0 96 799
use nand3 g7966
timestamp 1396952988
transform 1 0 9915 0 1 1018
box 0 0 120 799
use inv g8279
timestamp 1386238110
transform 1 0 10035 0 1 1018
box 0 0 120 799
use nand2 g8105
timestamp 1386234792
transform 1 0 10155 0 1 1018
box 0 0 96 799
use nand2 g8259
timestamp 1386234792
transform 1 0 10251 0 1 1018
box 0 0 96 799
use inv g8129
timestamp 1386238110
transform 1 0 10347 0 1 1018
box 0 0 120 799
use nand2 g8122
timestamp 1386234792
transform 1 0 10467 0 1 1018
box 0 0 96 799
use inv g8059
timestamp 1386238110
transform 1 0 10563 0 1 1018
box 0 0 120 799
use nand2 g8097
timestamp 1386234792
transform 1 0 10683 0 1 1018
box 0 0 96 799
use nand2 g8062
timestamp 1386234792
transform 1 0 10779 0 1 1018
box 0 0 96 799
use nand2 g8025
timestamp 1386234792
transform 1 0 10875 0 1 1018
box 0 0 96 799
use nand2 g8247
timestamp 1386234792
transform 1 0 10971 0 1 1018
box 0 0 96 799
use nor2 IntStatus_reg
timestamp 1386235306
transform 1 0 11067 0 1 1018
box 0 0 120 799
use scanreg g8263
timestamp 1386241447
transform 1 0 11187 0 1 1018
box 0 0 720 799
use nand2 g8131
timestamp 1386234792
transform 1 0 11907 0 1 1018
box 0 0 96 799
use nand2 g8256
timestamp 1386234792
transform 1 0 12003 0 1 1018
box 0 0 96 799
use inv g8087
timestamp 1386238110
transform 1 0 12099 0 1 1018
box 0 0 120 799
use and2 g7970
timestamp 1386234845
transform 1 0 12219 0 1 1018
box 0 0 120 799
use nand2 g7932
timestamp 1386234792
transform 1 0 12339 0 1 1018
box 0 0 96 799
use nand4 g7991
timestamp 1386234936
transform 1 0 12435 0 1 1018
box 0 0 144 799
use nand3 g8137
timestamp 1396952988
transform 1 0 12579 0 1 1018
box 0 0 120 799
use and2 g8201
timestamp 1386234845
transform 1 0 12699 0 1 1018
box 0 0 120 799
use nor2 g7952
timestamp 1386235306
transform 1 0 12819 0 1 1018
box 0 0 120 799
use nand3 g7936
timestamp 1396952988
transform 1 0 12939 0 1 1018
box 0 0 120 799
use nand2 g8207
timestamp 1386234792
transform 1 0 13059 0 1 1018
box 0 0 96 799
use nand2 g8044
timestamp 1386234792
transform 1 0 13155 0 1 1018
box 0 0 96 799
use nand2 g8006
timestamp 1386234792
transform 1 0 13251 0 1 1018
box 0 0 96 799
use nand2 g8173
timestamp 1386234792
transform 1 0 13347 0 1 1018
box 0 0 96 799
use nand2 g7983
timestamp 1386234792
transform 1 0 13443 0 1 1018
box 0 0 96 799
use nand2 g8157
timestamp 1386234792
transform 1 0 13539 0 1 1018
box 0 0 96 799
use nand3 g7956
timestamp 1396952988
transform 1 0 13635 0 1 1018
box 0 0 120 799
use nand2 g8040
timestamp 1386234792
transform 1 0 13755 0 1 1018
box 0 0 96 799
use nand3 g8068
timestamp 1396952988
transform 1 0 13851 0 1 1018
box 0 0 120 799
use and2 g8140
timestamp 1386234845
transform 1 0 13971 0 1 1018
box 0 0 120 799
use nand2 g8141
timestamp 1386234792
transform 1 0 14091 0 1 1018
box 0 0 96 799
use and2 g8210
timestamp 1386234845
transform 1 0 14187 0 1 1018
box 0 0 120 799
use nand2 g8003
timestamp 1386234792
transform 1 0 14307 0 1 1018
box 0 0 96 799
use nand2 g8203
timestamp 1386234792
transform 1 0 14403 0 1 1018
box 0 0 96 799
use inv g8065
timestamp 1386238110
transform 1 0 14499 0 1 1018
box 0 0 120 799
use nand2 g8113
timestamp 1386234792
transform 1 0 14619 0 1 1018
box 0 0 96 799
use inv g7977
timestamp 1386238110
transform 1 0 14715 0 1 1018
box 0 0 120 799
use nand2 g8070
timestamp 1386234792
transform 1 0 14835 0 1 1018
box 0 0 96 799
use nand4 g8038
timestamp 1386234936
transform 1 0 14931 0 1 1018
box 0 0 144 799
use nand2 IRQ2_reg
timestamp 1386234792
transform 1 0 15075 0 1 1018
box 0 0 96 799
use scandtype g8233
timestamp 1386241841
transform 1 0 15171 0 1 1018
box 0 0 624 799
use nand2 g7980
timestamp 1386234792
transform 1 0 15795 0 1 1018
box 0 0 96 799
use nand4 g7954
timestamp 1386234936
transform 1 0 15891 0 1 1018
box 0 0 144 799
use nor2 g8151
timestamp 1386235306
transform 1 0 16035 0 1 1018
box 0 0 120 799
use nand2 g7920
timestamp 1386234792
transform 1 0 16155 0 1 1018
box 0 0 96 799
use nand4 g8138
timestamp 1386234936
transform 1 0 16251 0 1 1018
box 0 0 144 799
use nand2 g7968
timestamp 1386234792
transform 1 0 16395 0 1 1018
box 0 0 96 799
use nand2 g8188
timestamp 1386234792
transform 1 0 16491 0 1 1018
box 0 0 96 799
use and2 g8176
timestamp 1386234845
transform 1 0 16587 0 1 1018
box 0 0 120 799
use nand2 g8172
timestamp 1386234792
transform 1 0 16707 0 1 1018
box 0 0 96 799
use and2 g8026
timestamp 1386234845
transform 1 0 16803 0 1 1018
box 0 0 120 799
use mux2 g8031
timestamp 1386235218
transform 1 0 16923 0 1 1018
box 0 0 192 799
use nand2 g7935
timestamp 1386234792
transform 1 0 17115 0 1 1018
box 0 0 96 799
use nand2 g8162
timestamp 1386234792
transform 1 0 17211 0 1 1018
box 0 0 96 799
use nand3 g8095
timestamp 1396952988
transform 1 0 17307 0 1 1018
box 0 0 120 799
use nand3 g7950
timestamp 1396952988
transform 1 0 17427 0 1 1018
box 0 0 120 799
use nor2 g8008
timestamp 1386235306
transform 1 0 17547 0 1 1018
box 0 0 120 799
use nand2 g8013
timestamp 1386234792
transform 1 0 17667 0 1 1018
box 0 0 96 799
use nand2 g8299
timestamp 1386234792
transform 1 0 17763 0 1 1018
box 0 0 96 799
use rowcrosser Flags_91_1_93_
timestamp 1397224710
transform 1 0 17859 0 1 1018
box 0 0 48 799
use inv g7984
timestamp 1386238110
transform 1 0 17907 0 1 1018
box 0 0 120 799
use nand4 g8126
timestamp 1386234936
transform 1 0 18027 0 1 1018
box 0 0 144 799
use nand4 IRQ1_reg
timestamp 1386234936
transform 1 0 18171 0 1 1018
box 0 0 144 799
use scandtype g7986
timestamp 1386241841
transform 1 0 18315 0 1 1018
box 0 0 624 799
use nand2 rm_assigns_buf_MemEn
timestamp 1386234792
transform 1 0 18939 0 1 1018
box 0 0 96 799
use buffer g8205
timestamp 1386236986
transform 1 0 19035 0 1 1018
box 0 0 120 799
use nor2 g8164
timestamp 1386235306
transform 1 0 19155 0 1 1018
box 0 0 120 799
use nand2 g7949
timestamp 1386234792
transform 1 0 19275 0 1 1018
box 0 0 96 799
use nand4 g8017
timestamp 1386234936
transform 1 0 19371 0 1 1018
box 0 0 144 799
use nand2 g8010
timestamp 1386234792
transform 1 0 19515 0 1 1018
box 0 0 96 799
use nand2 g8165
timestamp 1386234792
transform 1 0 19611 0 1 1018
box 0 0 96 799
use nand2 g8260
timestamp 1386234792
transform 1 0 19707 0 1 1018
box 0 0 96 799
use nand2 g8245
timestamp 1386234792
transform 1 0 19803 0 1 1018
box 0 0 96 799
use nand2 g8034
timestamp 1386234792
transform 1 0 19899 0 1 1018
box 0 0 96 799
use nand2 g8215
timestamp 1386234792
transform 1 0 19995 0 1 1018
box 0 0 96 799
use nand2 g8079
timestamp 1386234792
transform 1 0 20091 0 1 1018
box 0 0 96 799
use nor2 g7999
timestamp 1386235306
transform 1 0 20187 0 1 1018
box 0 0 120 799
use nor2 g8239
timestamp 1386235306
transform 1 0 20307 0 1 1018
box 0 0 120 799
use nor2 g8007
timestamp 1386235306
transform 1 0 20427 0 1 1018
box 0 0 120 799
use rowcrosser g8197
timestamp 1397224710
transform 1 0 20547 0 1 1018
box 0 0 48 799
use inv g8262
timestamp 1386238110
transform 1 0 20595 0 1 1018
box 0 0 120 799
use inv g7965
timestamp 1386238110
transform 1 0 20715 0 1 1018
box 0 0 120 799
use nand4 g8109
timestamp 1386234936
transform 1 0 20835 0 1 1018
box 0 0 144 799
use nand2 g8085
timestamp 1386234792
transform 1 0 20979 0 1 1018
box 0 0 96 799
use nand2 g8298
timestamp 1386234792
transform 1 0 21075 0 1 1018
box 0 0 96 799
use inv g7944
timestamp 1386238110
transform 1 0 21171 0 1 1018
box 0 0 120 799
use nand4 g8021
timestamp 1386234936
transform 1 0 21291 0 1 1018
box 0 0 144 799
use nand2 g7961
timestamp 1386234792
transform 1 0 21435 0 1 1018
box 0 0 96 799
use nand3 g7931
timestamp 1396952988
transform 1 0 21531 0 1 1018
box 0 0 120 799
use nand4 g8184
timestamp 1386234936
transform 1 0 21651 0 1 1018
box 0 0 144 799
use nand2 g7938
timestamp 1386234792
transform 1 0 21795 0 1 1018
box 0 0 96 799
use nand3 g8132
timestamp 1396952988
transform 1 0 21891 0 1 1018
box 0 0 120 799
use nand2 g8219
timestamp 1386234792
transform 1 0 22011 0 1 1018
box 0 0 96 799
use and2 g8061
timestamp 1386234845
transform 1 0 22107 0 1 1018
box 0 0 120 799
use nand4 g8258
timestamp 1386234936
transform 1 0 22227 0 1 1018
box 0 0 144 799
use nand2 g8115
timestamp 1386234792
transform 1 0 22371 0 1 1018
box 0 0 96 799
use nor2 g8202
timestamp 1386235306
transform 1 0 22467 0 1 1018
box 0 0 120 799
use nand2 g7973
timestamp 1386234792
transform 1 0 22587 0 1 1018
box 0 0 96 799
use nand2 g8246
timestamp 1386234792
transform 1 0 22683 0 1 1018
box 0 0 96 799
use nand2 g8208
timestamp 1386234792
transform 1 0 22779 0 1 1018
box 0 0 96 799
use nand2 g7958
timestamp 1386234792
transform 1 0 22875 0 1 1018
box 0 0 96 799
use nand3 g8156
timestamp 1396952988
transform 1 0 22971 0 1 1018
box 0 0 120 799
use and2 g8231
timestamp 1386234845
transform 1 0 23091 0 1 1018
box 0 0 120 799
use inv g8047
timestamp 1386238110
transform 1 0 23211 0 1 1018
box 0 0 120 799
use nand2 g7957
timestamp 1386234792
transform 1 0 23331 0 1 1018
box 0 0 96 799
use nand2 g8179
timestamp 1386234792
transform 1 0 23427 0 1 1018
box 0 0 96 799
use inv g8022
timestamp 1386238110
transform 1 0 23523 0 1 1018
box 0 0 120 799
use nand2 g8193
timestamp 1386234792
transform 1 0 23643 0 1 1018
box 0 0 96 799
use nand2 g8071
timestamp 1386234792
transform 1 0 23739 0 1 1018
box 0 0 96 799
use nand3 g8285
timestamp 1396952988
transform 1 0 23835 0 1 1018
box 0 0 120 799
use nand2 g8083
timestamp 1386234792
transform 1 0 23955 0 1 1018
box 0 0 96 799
use nand2 g7953
timestamp 1386234792
transform 1 0 24051 0 1 1018
box 0 0 96 799
use nand4 g8204
timestamp 1386234936
transform 1 0 24147 0 1 1018
box 0 0 144 799
use nand2 g8053
timestamp 1386234792
transform 1 0 24291 0 1 1018
box 0 0 96 799
use nand2 g8000
timestamp 1386234792
transform 1 0 24387 0 1 1018
box 0 0 96 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 24483 0 1 1018
box 0 0 96 799
use scandtype g8142
timestamp 1386241841
transform 1 0 24579 0 1 1018
box 0 0 624 799
use inv stateSub_reg_91_1_93_
timestamp 1386238110
transform 1 0 25203 0 1 1018
box 0 0 120 799
use scandtype g7914
timestamp 1386241841
transform 1 0 25323 0 1 1018
box 0 0 624 799
use nand3 g8075
timestamp 1396952988
transform 1 0 25947 0 1 1018
box 0 0 120 799
use nand4 g7994
timestamp 1386234936
transform 1 0 26067 0 1 1018
box 0 0 144 799
use nand2 g8032
timestamp 1386234792
transform 1 0 26211 0 1 1018
box 0 0 96 799
use nand2 g7941
timestamp 1386234792
transform 1 0 26307 0 1 1018
box 0 0 96 799
use nand4 SysBus_91_0_93_
timestamp 1386234936
transform 1 0 26403 0 1 1018
box 0 0 144 799
use rowcrosser CFlag
timestamp 1397224710
transform 1 0 26547 0 1 1018
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27050 0 1 1018
box 0 0 320 799
<< labels >>
rlabel m2contact 27081 3850 27081 3850 6 Rs1Sel[1]
rlabel m2contact 27081 1882 27081 1882 6 Rs1Sel[1]
rlabel m2contact 27057 3634 27057 3634 6 Rs1Sel[0]
rlabel m2contact 27057 1858 27057 1858 6 Rs1Sel[0]
rlabel m2contact 27033 1978 27033 1978 6 Flags[3]
rlabel m2contact 27033 1834 27033 1834 6 Flags[3]
rlabel m2contact 27033 5506 27033 5506 6 AluOR[0]
rlabel m2contact 27009 7210 27009 7210 6 n_350
rlabel m2contact 27009 4498 27009 4498 6 n_350
rlabel m2contact 26985 6346 26985 6346 6 n_128
rlabel m2contact 26961 4162 26961 4162 6 n_182
rlabel m2contact 26937 4930 26937 4930 6 n_235
rlabel m2contact 26913 5842 26913 5842 6 n_349
rlabel m2contact 26913 4378 26913 4378 6 n_349
rlabel m2contact 26889 3706 26889 3706 6 n_228
rlabel m2contact 26865 4546 26865 4546 6 n_186
rlabel m2contact 26841 3490 26841 3490 6 n_187
rlabel m2contact 26817 5986 26817 5986 6 n_60
rlabel m2contact 26781 6610 26781 6610 6 n_136
rlabel m2contact 26781 3922 26781 3922 6 n_136
rlabel m2contact 26769 6922 26769 6922 6 n_118
rlabel m2contact 26745 5770 26745 5770 6 n_141
rlabel m2contact 26721 4306 26721 4306 6 n_117
rlabel m2contact 26697 6202 26697 6202 6 n_41
rlabel m2contact 26697 2098 26697 2098 6 n_41
rlabel m2contact 26673 3034 26673 3034 6 n_226
rlabel m2contact 26649 4426 26649 4426 6 n_140
rlabel m2contact 26625 2002 26625 2002 6 n_225
rlabel m2contact 26601 3874 26601 3874 6 n_101
rlabel m2contact 26577 5866 26577 5866 6 n_325
rlabel m2contact 26577 3994 26577 3994 6 Flags[1]
rlabel m2contact 26541 5818 26541 5818 6 n_63
rlabel m2contact 26541 4522 26541 4522 6 n_63
rlabel m2contact 26529 4498 26529 4498 6 n_350
rlabel m2contact 26529 6394 26529 6394 6 n_256
rlabel m2contact 26505 4378 26505 4378 6 n_349
rlabel m2contact 26505 4402 26505 4402 6 OpcodeCondIn[6]
rlabel m2contact 26481 3922 26481 3922 6 n_136
rlabel m2contact 26481 3946 26481 3946 6 n_255
rlabel m2contact 26457 4570 26457 4570 6 state[0]
rlabel m2contact 26457 3154 26457 3154 6 state[0]
rlabel m2contact 26433 6202 26433 6202 6 n_41
rlabel m2contact 26433 6178 26433 6178 6 n_227
rlabel m2contact 26409 4258 26409 4258 6 n_39
rlabel m2contact 26385 2410 26385 2410 6 n_40
rlabel m2contact 26361 3970 26361 3970 6 n_293
rlabel m2contact 26337 5818 26337 5818 6 n_63
rlabel m2contact 26337 5794 26337 5794 6 n_292
rlabel m2contact 26313 2794 26313 2794 6 n_48
rlabel m2contact 26289 2410 26289 2410 6 n_40
rlabel m2contact 26265 4258 26265 4258 6 n_39
rlabel m2contact 26265 1906 26265 1906 6 n_236
rlabel m2contact 26241 7018 26241 7018 6 n_280
rlabel m2contact 26217 6154 26217 6154 6 n_176
rlabel m2contact 26193 4210 26193 4210 6 n_122
rlabel m2contact 26193 2746 26193 2746 6 n_166
rlabel m2contact 26169 4570 26169 4570 6 state[0]
rlabel m2contact 26169 3658 26169 3658 6 n_16
rlabel m2contact 26121 2794 26121 2794 6 n_48
rlabel m2contact 26097 4522 26097 4522 6 n_63
rlabel m2contact 26073 5242 26073 5242 6 OpcodeCondIn[0]
rlabel m2contact 26049 2842 26049 2842 6 n_20
rlabel m2contact 26025 5698 26025 5698 6 n_370
rlabel m2contact 26025 1858 26025 1858 6 n_370
rlabel m2contact 26001 3010 26001 3010 6 n_72
rlabel m2contact 25977 1858 25977 1858 6 n_370
rlabel m2contact 25977 1882 25977 1882 6 n_71
rlabel m2contact 25953 3802 25953 3802 6 n_251
rlabel m2contact 25905 2146 25905 2146 6 n_250
rlabel m2contact 25881 6466 25881 6466 6 stateSub[1]
rlabel m2contact 25881 4522 25881 4522 6 stateSub[1]
rlabel m2contact 25857 3250 25857 3250 6 OpcodeCondIn[4]
rlabel m2contact 25833 4522 25833 4522 6 stateSub[1]
rlabel m2contact 25833 5290 25833 5290 6 n_192
rlabel m2contact 25785 4738 25785 4738 6 n_103
rlabel m2contact 25761 4282 25761 4282 6 n_200
rlabel m2contact 25737 4642 25737 4642 6 n_352
rlabel m2contact 25713 2914 25713 2914 6 n_249
rlabel m2contact 25665 6106 25665 6106 6 n_289
rlabel m2contact 25617 4378 25617 4378 6 n_7
rlabel m2contact 25593 3394 25593 3394 6 n_252
rlabel m2contact 25545 4498 25545 4498 6 n_91
rlabel m2contact 25521 2698 25521 2698 6 OpcodeCondIn[7]
rlabel m2contact 25497 3370 25497 3370 6 n_92
rlabel m2contact 25449 4666 25449 4666 6 n_233
rlabel m2contact 25425 5650 25425 5650 6 n_158
rlabel m2contact 25401 4618 25401 4618 6 n_244
rlabel m2contact 25353 6250 25353 6250 6 n_321
rlabel m2contact 25305 5530 25305 5530 6 n_173
rlabel m2contact 25281 2722 25281 2722 6 n_302
rlabel m2contact 25233 6202 25233 6202 6 n_44
rlabel m2contact 25233 5938 25233 5938 6 n_111
rlabel m2contact 25209 6466 25209 6466 6 stateSub[1]
rlabel m2contact 25185 4690 25185 4690 6 state[1]
rlabel m2contact 25137 4786 25137 4786 6 n_83
rlabel m2contact 25113 4690 25113 4690 6 state[1]
rlabel m2contact 25089 4234 25089 4234 6 n_55
rlabel m2contact 25089 3154 25089 3154 6 state[0]
rlabel m2contact 25041 5698 25041 5698 6 n_370
rlabel m2contact 25041 5674 25041 5674 6 n_68
rlabel m2contact 25017 3274 25017 3274 6 StatusReg[2]
rlabel m2contact 24993 4570 24993 4570 6 n_371
rlabel m2contact 24945 3226 24945 3226 6 n_333
rlabel m2contact 24921 5098 24921 5098 6 n_139
rlabel m2contact 24897 4450 24897 4450 6 n_288
rlabel m2contact 24873 6034 24873 6034 6 n_208
rlabel m2contact 24849 4114 24849 4114 6 n_203
rlabel m2contact 24801 4186 24801 4186 6 RwSel[1]
rlabel m2contact 24729 2962 24729 2962 6 n_254
rlabel m2contact 24681 7066 24681 7066 6 n_222
rlabel m2contact 24633 3466 24633 3466 6 n_25
rlabel m2contact 24609 4594 24609 4594 6 n_338
rlabel m2contact 24609 4330 24609 4330 6 n_338
rlabel m2contact 24585 4354 24585 4354 6 OpcodeCondIn[3]
rlabel m2contact 24561 4066 24561 4066 6 OpcodeCondIn[5]
rlabel m2contact 24537 3802 24537 3802 6 n_251
rlabel m2contact 24513 4474 24513 4474 6 n_358
rlabel m2contact 24489 4714 24489 4714 6 n_318
rlabel m2contact 24489 2338 24489 2338 6 n_318
rlabel m2contact 24465 3058 24465 3058 6 n_232
rlabel m2contact 24441 4594 24441 4594 6 n_338
rlabel m2contact 24441 4522 24441 4522 6 n_137
rlabel m2contact 24417 2338 24417 2338 6 n_318
rlabel m2contact 24393 2074 24393 2074 6 n_77
rlabel m2contact 24369 5674 24369 5674 6 n_68
rlabel m2contact 24345 1906 24345 1906 6 n_236
rlabel m2contact 24345 3610 24345 3610 6 n_133
rlabel m2contact 24321 4714 24321 4714 6 n_318
rlabel m2contact 24321 4090 24321 4090 6 n_30
rlabel m2contact 24297 4594 24297 4594 6 n_236
rlabel m2contact 24297 1906 24297 1906 6 n_236
rlabel m2contact 24273 4186 24273 4186 6 RwSel[1]
rlabel m2contact 24249 3898 24249 3898 6 n_195
rlabel m2contact 24225 4330 24225 4330 6 n_338
rlabel m2contact 24201 2530 24201 2530 6 n_86
rlabel m2contact 24177 5482 24177 5482 6 n_298
rlabel m2contact 24153 7114 24153 7114 6 n_35
rlabel m2contact 24153 4042 24153 4042 6 n_35
rlabel m2contact 24129 4426 24129 4426 6 n_140
rlabel m2contact 24129 4666 24129 4666 6 n_233
rlabel m2contact 24105 2674 24105 2674 6 n_313
rlabel m2contact 24081 3802 24081 3802 6 n_251
rlabel m2contact 24057 4426 24057 4426 6 n_206
rlabel m2contact 24033 4378 24033 4378 6 n_7
rlabel m2contact 24009 4594 24009 4594 6 n_236
rlabel m2contact 24009 4402 24009 4402 6 OpcodeCondIn[6]
rlabel m2contact 23985 6970 23985 6970 6 n_21
rlabel m2contact 23985 4138 23985 4138 6 stateSub[0]
rlabel m2contact 23949 5818 23949 5818 6 stateSub[2]
rlabel m2contact 23949 4378 23949 4378 6 stateSub[2]
rlabel m2contact 23937 3082 23937 3082 6 n_223
rlabel m2contact 23937 5962 23937 5962 6 n_157
rlabel m2contact 23913 5914 23913 5914 6 n_156
rlabel m2contact 23913 4402 23913 4402 6 OpcodeCondIn[6]
rlabel m2contact 23889 4666 23889 4666 6 n_121
rlabel m2contact 23889 2434 23889 2434 6 n_190
rlabel m2contact 23865 6538 23865 6538 6 n_64
rlabel m2contact 23841 1858 23841 1858 6 n_214
rlabel m2contact 23817 4906 23817 4906 6 n_76
rlabel m2contact 23793 4042 23793 4042 6 n_35
rlabel m2contact 23793 4138 23793 4138 6 stateSub[0]
rlabel m2contact 23769 4378 23769 4378 6 stateSub[2]
rlabel m2contact 23769 5218 23769 5218 6 n_152
rlabel m2contact 23745 4834 23745 4834 6 n_190
rlabel m2contact 23745 2434 23745 2434 6 n_190
rlabel m2contact 23721 6490 23721 6490 6 n_286
rlabel m2contact 23721 6778 23721 6778 6 n_191
rlabel m2contact 23697 2554 23697 2554 6 n_180
rlabel m2contact 23697 4978 23697 4978 6 n_160
rlabel m2contact 23673 4834 23673 4834 6 n_190
rlabel m2contact 23673 4810 23673 4810 6 n_258
rlabel m2contact 23625 4594 23625 4594 6 n_96
rlabel m2contact 23601 7138 23601 7138 6 PcSel[2]
rlabel m2contact 23577 4858 23577 4858 6 n_95
rlabel m2contact 23553 2314 23553 2314 6 n_340
rlabel m2contact 23553 3370 23553 3370 6 n_92
rlabel m2contact 23505 6442 23505 6442 6 n_300
rlabel m2contact 23481 2338 23481 2338 6 n_318
rlabel m2contact 23481 5698 23481 5698 6 n_210
rlabel m2contact 23457 6658 23457 6658 6 n_234
rlabel m2contact 23457 2890 23457 2890 6 n_317
rlabel m2contact 23409 4114 23409 4114 6 n_203
rlabel m2contact 23409 4186 23409 4186 6 PcSel[1]
rlabel m2contact 23385 4954 23385 4954 6 n_161
rlabel m2contact 23361 2818 23361 2818 6 n_202
rlabel m2contact 23337 3922 23337 3922 6 n_243
rlabel m2contact 23313 6082 23313 6082 6 n_51
rlabel m2contact 23313 3346 23313 3346 6 n_51
rlabel m2contact 23289 2194 23289 2194 6 n_171
rlabel m2contact 23289 4354 23289 4354 6 OpcodeCondIn[3]
rlabel m2contact 23253 4714 23253 4714 6 n_105
rlabel m2contact 23253 2242 23253 2242 6 n_105
rlabel m2contact 23241 5482 23241 5482 6 n_298
rlabel m2contact 23217 4162 23217 4162 6 n_182
rlabel m2contact 23193 6586 23193 6586 6 n_209
rlabel m2contact 23193 3490 23193 3490 6 n_187
rlabel m2contact 23157 6562 23157 6562 6 n_310
rlabel m2contact 23157 4378 23157 4378 6 n_310
rlabel m2contact 23145 3250 23145 3250 6 OpcodeCondIn[4]
rlabel m2contact 23121 4714 23121 4714 6 n_105
rlabel m2contact 23121 4114 23121 4114 6 n_150
rlabel m2contact 23097 5074 23097 5074 6 n_287
rlabel m2contact 23073 4186 23073 4186 6 PcSel[1]
rlabel m2contact 23049 4666 23049 4666 6 n_121
rlabel m2contact 23049 2314 23049 2314 6 n_340
rlabel m2contact 23025 2218 23025 2218 6 n_328
rlabel m2contact 23025 4402 23025 4402 6 OpcodeCondIn[6]
rlabel m2contact 23001 3202 23001 3202 6 n_84
rlabel m2contact 22977 2602 22977 2602 6 n_37
rlabel m2contact 22953 4234 22953 4234 6 n_55
rlabel m2contact 22929 5722 22929 5722 6 n_127
rlabel m2contact 22929 5674 22929 5674 6 n_68
rlabel m2contact 22905 3874 22905 3874 6 n_101
rlabel m2contact 22881 2986 22881 2986 6 n_32
rlabel m2contact 22857 4258 22857 4258 6 n_39
rlabel m2contact 22857 4594 22857 4594 6 n_96
rlabel m2contact 22833 6010 22833 6010 6 n_196
rlabel m2contact 22833 3586 22833 3586 6 n_196
rlabel m2contact 22809 6082 22809 6082 6 n_51
rlabel m2contact 22809 6058 22809 6058 6 StatusReg[3]
rlabel m2contact 22785 6754 22785 6754 6 n_27
rlabel m2contact 22761 4378 22761 4378 6 n_310
rlabel m2contact 22761 6202 22761 6202 6 n_44
rlabel m2contact 22737 4594 22737 4594 6 n_361
rlabel m2contact 22737 2050 22737 2050 6 n_361
rlabel m2contact 22713 5170 22713 5170 6 n_89
rlabel m2contact 22713 3682 22713 3682 6 n_309
rlabel m2contact 22689 4378 22689 4378 6 IRQ2
rlabel m2contact 22665 2578 22665 2578 6 IntStatus
rlabel m2contact 22641 1906 22641 1906 6 n_236
rlabel m2contact 22617 2794 22617 2794 6 n_48
rlabel m2contact 22617 2818 22617 2818 6 n_202
rlabel m2contact 22593 2938 22593 2938 6 n_102
rlabel m2contact 22569 3586 22569 3586 6 n_196
rlabel m2contact 22569 3730 22569 3730 6 n_130
rlabel m2contact 22545 5410 22545 5410 6 n_164
rlabel m2contact 22545 4258 22545 4258 6 n_164
rlabel m2contact 22521 5650 22521 5650 6 n_158
rlabel m2contact 22497 4594 22497 4594 6 n_361
rlabel m2contact 22497 3298 22497 3298 6 n_159
rlabel m2contact 22461 4714 22461 4714 6 AluEn
rlabel m2contact 22461 4234 22461 4234 6 AluEn
rlabel m2contact 22449 4882 22449 4882 6 n_365
rlabel m2contact 22449 4042 22449 4042 6 n_17
rlabel m2contact 22425 4738 22425 4738 6 n_103
rlabel m2contact 22401 4714 22401 4714 6 AluEn
rlabel m2contact 22401 4690 22401 4690 6 state[1]
rlabel m2contact 22377 6226 22377 6226 6 n_20
rlabel m2contact 22377 2842 22377 2842 6 n_20
rlabel m2contact 22353 7042 22353 7042 6 n_98
rlabel m2contact 22353 5386 22353 5386 6 n_168
rlabel m2contact 22329 6466 22329 6466 6 stateSub[1]
rlabel m2contact 22329 5602 22329 5602 6 n_167
rlabel m2contact 22305 4258 22305 4258 6 n_164
rlabel m2contact 22305 4714 22305 4714 6 n_104
rlabel m2contact 22281 4162 22281 4162 6 n_182
rlabel m2contact 22257 7090 22257 7090 6 n_19
rlabel m2contact 22257 5554 22257 5554 6 n_198
rlabel m2contact 22233 2698 22233 2698 6 OpcodeCondIn[7]
rlabel m2contact 22209 6226 22209 6226 6 n_20
rlabel m2contact 22209 6130 22209 6130 6 n_259
rlabel m2contact 22161 4258 22161 4258 6 AluWe
rlabel m2contact 22161 4162 22161 4162 6 n_182
rlabel m2contact 22137 2338 22137 2338 6 n_318
rlabel m2contact 22089 4210 22089 4210 6 n_122
rlabel m2contact 22041 2386 22041 2386 6 n_135
rlabel m2contact 22017 6370 22017 6370 6 n_270
rlabel m2contact 22017 2290 22017 2290 6 n_270
rlabel m2contact 21993 4234 21993 4234 6 AluEn
rlabel m2contact 21969 2290 21969 2290 6 n_270
rlabel m2contact 21969 2362 21969 2362 6 n_400
rlabel m2contact 21921 4474 21921 4474 6 n_358
rlabel m2contact 21873 3826 21873 3826 6 n_99
rlabel m2contact 21849 5770 21849 5770 6 n_141
rlabel m2contact 21825 6298 21825 6298 6 n_154
rlabel m2contact 21777 4258 21777 4258 6 AluWe
rlabel m2contact 21729 4474 21729 4474 6 n_358
rlabel m2contact 21681 5626 21681 5626 6 n_142
rlabel m2contact 21633 6226 21633 6226 6 n_45
rlabel m2contact 21633 4474 21633 4474 6 n_45
rlabel m2contact 21609 4474 21609 4474 6 n_45
rlabel m2contact 21609 5122 21609 5122 6 n_381
rlabel m2contact 21561 6274 21561 6274 6 n_323
rlabel m2contact 21537 5914 21537 5914 6 n_156
rlabel m2contact 21537 4210 21537 4210 6 n_156
rlabel m2contact 21513 6994 21513 6994 6 n_8
rlabel m2contact 21513 2770 21513 2770 6 n_8
rlabel m2contact 21489 4210 21489 4210 6 n_156
rlabel m2contact 21489 4234 21489 4234 6 n_52
rlabel m2contact 21465 3322 21465 3322 6 n_148
rlabel m2contact 21465 4930 21465 4930 6 n_235
rlabel m2contact 21441 3178 21441 3178 6 n_62
rlabel m2contact 21417 5890 21417 5890 6 n_50
rlabel m2contact 21417 4258 21417 4258 6 n_50
rlabel m2contact 21393 2770 21393 2770 6 n_8
rlabel m2contact 21393 2794 21393 2794 6 n_100
rlabel m2contact 21369 2338 21369 2338 6 n_318
rlabel m2contact 21345 4258 21345 4258 6 n_50
rlabel m2contact 21345 4714 21345 4714 6 n_104
rlabel m2contact 21321 6898 21321 6898 6 n_178
rlabel m2contact 21321 4474 21321 4474 6 n_178
rlabel m2contact 21297 6730 21297 6730 6 n_11
rlabel m2contact 21273 5002 21273 5002 6 n_318
rlabel m2contact 21273 2338 21273 2338 6 n_318
rlabel m2contact 21249 2842 21249 2842 6 n_20
rlabel m2contact 21249 3802 21249 3802 6 n_251
rlabel m2contact 21225 4162 21225 4162 6 n_182
rlabel m2contact 21201 5266 21201 5266 6 OpcodeCondIn[1]
rlabel m2contact 21177 4330 21177 4330 6 n_338
rlabel m2contact 21153 5146 21153 5146 6 n_238
rlabel m2contact 21129 5458 21129 5458 6 n_344
rlabel m2contact 21129 3922 21129 3922 6 n_243
rlabel m2contact 21105 6322 21105 6322 6 n_262
rlabel m2contact 21105 3490 21105 3490 6 n_187
rlabel m2contact 21081 6298 21081 6298 6 n_154
rlabel m2contact 21081 3778 21081 3778 6 n_154
rlabel m2contact 21057 4474 21057 4474 6 n_178
rlabel m2contact 21057 5554 21057 5554 6 n_198
rlabel m2contact 21033 5770 21033 5770 6 n_141
rlabel m2contact 21009 2434 21009 2434 6 n_190
rlabel m2contact 21009 4402 21009 4402 6 OpcodeCondIn[6]
rlabel m2contact 20985 4474 20985 4474 6 n_204
rlabel m2contact 20961 4762 20961 4762 6 Op2Sel[0]
rlabel m2contact 20937 4258 20937 4258 6 LrSel
rlabel m2contact 20913 4594 20913 4594 6 n_303
rlabel m2contact 20889 3106 20889 3106 6 n_57
rlabel m2contact 20865 3706 20865 3706 6 n_228
rlabel m2contact 20865 3754 20865 3754 6 n_56
rlabel m2contact 20841 4930 20841 4930 6 n_235
rlabel m2contact 20805 4834 20805 4834 6 n_356
rlabel m2contact 20805 2458 20805 2458 6 n_356
rlabel m2contact 20793 1882 20793 1882 6 n_71
rlabel m2contact 20793 5050 20793 5050 6 n_184
rlabel m2contact 20769 4162 20769 4162 6 n_182
rlabel m2contact 20745 2866 20745 2866 6 n_66
rlabel m2contact 20745 3706 20745 3706 6 n_183
rlabel m2contact 20709 2674 20709 2674 6 n_313
rlabel m2contact 20709 1954 20709 1954 6 n_313
rlabel m2contact 20709 4666 20709 4666 6 n_14
rlabel m2contact 20709 4018 20709 4018 6 n_14
rlabel m2contact 20697 4762 20697 4762 6 Op2Sel[0]
rlabel m2contact 20673 4258 20673 4258 6 LrSel
rlabel m2contact 20649 5362 20649 5362 6 n_372
rlabel m2contact 20625 1954 20625 1954 6 n_313
rlabel m2contact 20625 2026 20625 2026 6 CFlag
rlabel m2contact 20601 4570 20601 4570 6 n_371
rlabel m2contact 20577 2026 20577 2026 6 CFlag
rlabel m2contact 20553 4258 20553 4258 6 Op1Sel
rlabel m2contact 20529 4762 20529 4762 6 n_242
rlabel m2contact 20529 2770 20529 2770 6 n_242
rlabel m2contact 20505 3610 20505 3610 6 n_133
rlabel m2contact 20481 2170 20481 2170 6 n_6
rlabel m2contact 20457 4018 20457 4018 6 n_14
rlabel m2contact 20457 4162 20457 4162 6 n_182
rlabel m2contact 20433 5818 20433 5818 6 stateSub[2]
rlabel m2contact 20409 4258 20409 4258 6 Op1Sel
rlabel m2contact 20385 4210 20385 4210 6 n_319
rlabel m2contact 20361 5002 20361 5002 6 n_318
rlabel m2contact 20361 4426 20361 4426 6 n_206
rlabel m2contact 20337 6490 20337 6490 6 n_286
rlabel m2contact 20337 6418 20337 6418 6 n_264
rlabel m2contact 20301 7162 20301 7162 6 n_399
rlabel m2contact 20301 4186 20301 4186 6 n_399
rlabel m2contact 20289 3946 20289 3946 6 n_255
rlabel m2contact 20265 2314 20265 2314 6 n_340
rlabel m2contact 20241 3586 20241 3586 6 n_332
rlabel m2contact 20241 3250 20241 3250 6 OpcodeCondIn[4]
rlabel m2contact 20217 4834 20217 4834 6 n_356
rlabel m2contact 20217 4018 20217 4018 6 n_189
rlabel m2contact 20193 4018 20193 4018 6 n_189
rlabel m2contact 20169 5026 20169 5026 6 n_88
rlabel m2contact 20145 6370 20145 6370 6 n_270
rlabel m2contact 20145 5674 20145 5674 6 n_68
rlabel m2contact 20121 3778 20121 3778 6 n_154
rlabel m2contact 20121 4738 20121 4738 6 n_103
rlabel m2contact 20097 4258 20097 4258 6 n_61
rlabel m2contact 20073 4690 20073 4690 6 state[1]
rlabel m2contact 20049 3922 20049 3922 6 n_243
rlabel m2contact 20025 4762 20025 4762 6 n_242
rlabel m2contact 20025 4618 20025 4618 6 n_244
rlabel m2contact 20001 5314 20001 5314 6 n_231
rlabel m2contact 20001 3562 20001 3562 6 n_231
rlabel m2contact 19977 2410 19977 2410 6 n_40
rlabel m2contact 19977 2458 19977 2458 6 n_356
rlabel m2contact 19953 4186 19953 4186 6 n_399
rlabel m2contact 19953 5146 19953 5146 6 n_238
rlabel m2contact 19929 3274 19929 3274 6 StatusReg[2]
rlabel m2contact 19905 5194 19905 5194 6 n_266
rlabel m2contact 19905 3778 19905 3778 6 n_266
rlabel m2contact 19881 5314 19881 5314 6 n_231
rlabel m2contact 19881 5002 19881 5002 6 n_28
rlabel m2contact 19857 3802 19857 3802 6 n_251
rlabel m2contact 19833 6754 19833 6754 6 n_27
rlabel m2contact 19833 6466 19833 6466 6 stateSub[1]
rlabel m2contact 19809 6082 19809 6082 6 OpcodeCondIn[2]
rlabel m2contact 19809 4186 19809 4186 6 OpcodeCondIn[2]
rlabel m2contact 19785 4594 19785 4594 6 n_303
rlabel m2contact 19761 5194 19761 5194 6 n_266
rlabel m2contact 19761 4930 19761 4930 6 n_235
rlabel m2contact 19737 5794 19737 5794 6 n_292
rlabel m2contact 19713 3970 19713 3970 6 n_293
rlabel m2contact 19689 4450 19689 4450 6 n_288
rlabel m2contact 19665 5458 19665 5458 6 n_344
rlabel m2contact 19641 5674 19641 5674 6 n_68
rlabel m2contact 19641 5194 19641 5194 6 n_291
rlabel m2contact 19617 3874 19617 3874 6 n_101
rlabel m2contact 19593 3178 19593 3178 6 n_62
rlabel m2contact 19569 3442 19569 3442 6 n_120
rlabel m2contact 19545 5746 19545 5746 6 n_85
rlabel m2contact 19521 3130 19521 3130 6 n_10
rlabel m2contact 19497 2122 19497 2122 6 n_347
rlabel m2contact 19497 3154 19497 3154 6 state[0]
rlabel m2contact 19473 2290 19473 2290 6 n_46
rlabel m2contact 19449 3538 19449 3538 6 n_279
rlabel m2contact 19425 1954 19425 1954 6 ENB
rlabel m2contact 19389 4594 19389 4594 6 n_12
rlabel m2contact 19389 3418 19389 3418 6 n_12
rlabel m2contact 19377 4762 19377 4762 6 n_110
rlabel m2contact 19353 3562 19353 3562 6 n_231
rlabel m2contact 19329 3418 19329 3418 6 n_12
rlabel m2contact 19329 3514 19329 3514 6 n_81
rlabel m2contact 19305 4930 19305 4930 6 n_235
rlabel m2contact 19281 2506 19281 2506 6 n_199
rlabel m2contact 19257 5554 19257 5554 6 n_198
rlabel m2contact 19257 4834 19257 4834 6 n_261
rlabel m2contact 19233 4450 19233 4450 6 n_205
rlabel m2contact 19209 4186 19209 4186 6 OpcodeCondIn[2]
rlabel m2contact 19209 4426 19209 4426 6 n_206
rlabel m2contact 19161 4186 19161 4186 6 MemEn
rlabel m2contact 19113 4186 19113 4186 6 MemEn
rlabel m2contact 19113 5098 19113 5098 6 n_139
rlabel m2contact 19089 5938 19089 5938 6 n_111
rlabel m2contact 19065 1954 19065 1954 6 ENB
rlabel m2contact 19065 4114 19065 4114 6 n_150
rlabel m2contact 19017 3874 19017 3874 6 n_101
rlabel m2contact 18993 5818 18993 5818 6 stateSub[2]
rlabel m2contact 18969 4162 18969 4162 6 n_182
rlabel m2contact 18945 5818 18945 5818 6 stateSub[2]
rlabel m2contact 18873 5794 18873 5794 6 n_292
rlabel m2contact 18825 5146 18825 5146 6 n_238
rlabel m2contact 18777 6706 18777 6706 6 n_217
rlabel m2contact 18729 6490 18729 6490 6 n_170
rlabel m2contact 18705 4762 18705 4762 6 n_110
rlabel m2contact 18633 5458 18633 5458 6 n_344
rlabel m2contact 18609 6514 18609 6514 6 n_368
rlabel m2contact 18585 5434 18585 5434 6 n_221
rlabel m2contact 18561 2458 18561 2458 6 n_356
rlabel m2contact 18489 5770 18489 5770 6 n_141
rlabel m2contact 18441 5914 18441 5914 6 n_156
rlabel m2contact 18369 1834 18369 1834 6 n_194
rlabel m2contact 18321 3418 18321 3418 6 n_193
rlabel m2contact 18273 4402 18273 4402 6 OpcodeCondIn[6]
rlabel m2contact 18249 4642 18249 4642 6 n_352
rlabel m2contact 18249 4162 18249 4162 6 n_182
rlabel m2contact 18225 3778 18225 3778 6 n_266
rlabel m2contact 18201 6946 18201 6946 6 n_334
rlabel m2contact 18201 5338 18201 5338 6 n_132
rlabel m2contact 18177 7186 18177 7186 6 n_38
rlabel m2contact 18177 4186 18177 4186 6 n_38
rlabel m2contact 18153 5914 18153 5914 6 n_156
rlabel m2contact 18129 4186 18129 4186 6 n_38
rlabel m2contact 18129 4474 18129 4474 6 n_204
rlabel m2contact 18105 3970 18105 3970 6 n_293
rlabel m2contact 18033 6826 18033 6826 6 n_215
rlabel m2contact 17985 1858 17985 1858 6 n_214
rlabel m2contact 17937 5098 17937 5098 6 n_367
rlabel m2contact 17913 2650 17913 2650 6 Flags[0]
rlabel m2contact 17889 2650 17889 2650 6 Flags[0]
rlabel m2contact 17889 4882 17889 4882 6 n_365
rlabel m2contact 17865 5314 17865 5314 6 PcEn
rlabel m2contact 17865 4186 17865 4186 6 PcEn
rlabel m2contact 17841 6802 17841 6802 6 n_276
rlabel m2contact 17817 3970 17817 3970 6 n_293
rlabel m2contact 17793 5482 17793 5482 6 n_298
rlabel m2contact 17769 2698 17769 2698 6 OpcodeCondIn[7]
rlabel m2contact 17745 2674 17745 2674 6 n_313
rlabel m2contact 17721 5314 17721 5314 6 PcEn
rlabel m2contact 17721 4834 17721 4834 6 n_261
rlabel m2contact 17697 5194 17697 5194 6 n_291
rlabel m2contact 17649 2650 17649 2650 6 n_322
rlabel m2contact 17601 5578 17601 5578 6 n_147
rlabel m2contact 17577 2026 17577 2026 6 CFlag
rlabel m2contact 17529 2482 17529 2482 6 n_124
rlabel m2contact 17505 3106 17505 3106 6 n_57
rlabel m2contact 17481 2626 17481 2626 6 n_123
rlabel m2contact 17457 2266 17457 2266 6 n_5
rlabel m2contact 17409 3106 17409 3106 6 n_34
rlabel m2contact 17385 2602 17385 2602 6 n_37
rlabel m2contact 17361 4858 17361 4858 6 n_95
rlabel m2contact 17337 4546 17337 4546 6 n_186
rlabel m2contact 17241 4882 17241 4882 6 n_365
rlabel m2contact 17193 2914 17193 2914 6 n_249
rlabel m2contact 17169 4762 17169 4762 6 n_380
rlabel m2contact 17169 3970 17169 3970 6 n_293
rlabel m2contact 17145 2410 17145 2410 6 n_248
rlabel m2contact 17085 5314 17085 5314 6 n_143
rlabel m2contact 17085 4642 17085 4642 6 n_143
rlabel m2contact 17073 2914 17073 2914 6 n_268
rlabel m2contact 17049 5170 17049 5170 6 n_89
rlabel m2contact 17049 6682 17049 6682 6 n_24
rlabel m2contact 17025 3250 17025 3250 6 OpcodeCondIn[4]
rlabel m2contact 17001 1834 17001 1834 6 n_194
rlabel m2contact 17001 2674 17001 2674 6 n_59
rlabel m2contact 16977 4930 16977 4930 6 n_235
rlabel m2contact 16953 5602 16953 5602 6 n_167
rlabel m2contact 16929 6874 16929 6874 6 n_80
rlabel m2contact 16929 1834 16929 1834 6 n_80
rlabel m2contact 16905 4642 16905 4642 6 n_143
rlabel m2contact 16905 5266 16905 5266 6 OpcodeCondIn[1]
rlabel m2contact 16881 5242 16881 5242 6 OpcodeCondIn[0]
rlabel m2contact 16857 5554 16857 5554 6 n_198
rlabel m2contact 16833 5626 16833 5626 6 n_142
rlabel m2contact 16833 4930 16833 4930 6 n_235
rlabel m2contact 16809 3922 16809 3922 6 n_243
rlabel m2contact 16785 1834 16785 1834 6 n_80
rlabel m2contact 16785 4306 16785 4306 6 n_117
rlabel m2contact 16761 3346 16761 3346 6 n_51
rlabel m2contact 16761 5770 16761 5770 6 n_141
rlabel m2contact 16737 4258 16737 4258 6 n_61
rlabel m2contact 16713 4642 16713 4642 6 n_13
rlabel m2contact 16689 6082 16689 6082 6 OpcodeCondIn[2]
rlabel m2contact 16665 4354 16665 4354 6 OpcodeCondIn[3]
rlabel m2contact 16641 5602 16641 5602 6 n_167
rlabel m2contact 16617 2098 16617 2098 6 n_41
rlabel m2contact 16617 3346 16617 3346 6 n_146
rlabel m2contact 16593 6082 16593 6082 6 OpcodeCondIn[2]
rlabel m2contact 16569 3394 16569 3394 6 n_252
rlabel m2contact 16569 5626 16569 5626 6 n_163
rlabel m2contact 16545 3802 16545 3802 6 n_251
rlabel metal2 16521 6634 16521 6634 6 n_172
rlabel m2contact 16497 2194 16497 2194 6 n_171
rlabel m2contact 16473 4906 16473 4906 6 n_76
rlabel m2contact 16449 6850 16449 6850 6 n_138
rlabel m2contact 16449 5770 16449 5770 6 n_141
rlabel m2contact 16425 4114 16425 4114 6 n_150
rlabel m2contact 16401 4762 16401 4762 6 n_380
rlabel m2contact 16377 3850 16377 3850 6 Rs1Sel[1]
rlabel m2contact 16377 6562 16377 6562 6 n_310
rlabel m2contact 16353 4906 16353 4906 6 n_366
rlabel m2contact 16353 4762 16353 4762 6 n_297
rlabel m2contact 16329 5362 16329 5362 6 n_372
rlabel m2contact 16305 4330 16305 4330 6 n_338
rlabel m2contact 16281 5362 16281 5362 6 n_345
rlabel m2contact 16257 6418 16257 6418 6 n_264
rlabel m2contact 16209 2698 16209 2698 6 OpcodeCondIn[7]
rlabel m2contact 16209 5194 16209 5194 6 n_291
rlabel m2contact 16185 5578 16185 5578 6 n_147
rlabel m2contact 16137 6562 16137 6562 6 n_78
rlabel m2contact 16089 1858 16089 1858 6 n_214
rlabel m2contact 16089 2074 16089 2074 6 n_77
rlabel m2contact 16065 3850 16065 3850 6 n_305
rlabel m2contact 16041 3394 16041 3394 6 n_169
rlabel m2contact 16017 2698 16017 2698 6 OpcodeCondIn[7]
rlabel m2contact 15993 6634 15993 6634 6 n_125
rlabel m2contact 15993 4330 15993 4330 6 nWait
rlabel m2contact 15969 7234 15969 7234 6 n_271
rlabel m2contact 15969 2098 15969 2098 6 n_271
rlabel m2contact 15945 6418 15945 6418 6 n_151
rlabel m2contact 15945 4930 15945 4930 6 n_235
rlabel m2contact 15921 1906 15921 1906 6 n_236
rlabel m2contact 15921 3970 15921 3970 6 n_293
rlabel m2contact 15897 4114 15897 4114 6 n_150
rlabel m2contact 15873 2290 15873 2290 6 n_46
rlabel m2contact 15873 3754 15873 3754 6 n_56
rlabel m2contact 15849 4066 15849 4066 6 OpcodeCondIn[5]
rlabel m2contact 15825 7234 15825 7234 6 n_271
rlabel m2contact 15825 2866 15825 2866 6 n_66
rlabel m2contact 15801 6370 15801 6370 6 n_270
rlabel m2contact 15777 6778 15777 6778 6 n_191
rlabel m2contact 15753 6370 15753 6370 6 n_197
rlabel m2contact 15705 2290 15705 2290 6 PcSel[0]
rlabel m2contact 15681 4378 15681 4378 6 IRQ2
rlabel m2contact 15633 1906 15633 1906 6 n_236
rlabel m2contact 15585 6082 15585 6082 6 OpcodeCondIn[2]
rlabel m2contact 15441 5818 15441 5818 6 stateSub[2]
rlabel m2contact 15393 4930 15393 4930 6 n_235
rlabel m2contact 15129 6298 15129 6298 6 n_154
rlabel m2contact 15057 6778 15057 6778 6 n_144
rlabel m2contact 15033 7210 15033 7210 6 n_350
rlabel m2contact 15033 5650 15033 5650 6 n_158
rlabel m2contact 15009 3898 15009 3898 6 n_195
rlabel m2contact 14985 5314 14985 5314 6 n_143
rlabel m2contact 14961 3970 14961 3970 6 n_293
rlabel m2contact 14937 7210 14937 7210 6 n_225
rlabel m2contact 14937 2002 14937 2002 6 n_225
rlabel m2contact 14913 1930 14913 1930 6 RwSel[0]
rlabel m2contact 14889 7210 14889 7210 6 n_225
rlabel m2contact 14889 4378 14889 4378 6 n_74
rlabel m2contact 14865 6106 14865 6106 6 n_289
rlabel m2contact 14841 4786 14841 4786 6 n_83
rlabel m2contact 14817 2626 14817 2626 6 n_123
rlabel m2contact 14793 6106 14793 6106 6 n_177
rlabel m2contact 14745 6154 14745 6154 6 n_176
rlabel m2contact 14697 6130 14697 6130 6 n_259
rlabel m2contact 14697 1930 14697 1930 6 n_259
rlabel m2contact 14673 1930 14673 1930 6 n_259
rlabel m2contact 14673 6058 14673 6058 6 StatusReg[3]
rlabel m2contact 14649 4786 14649 4786 6 n_257
rlabel m2contact 14625 7162 14625 7162 6 n_399
rlabel m2contact 14457 3010 14457 3010 6 n_72
rlabel m2contact 14361 4738 14361 4738 6 n_103
rlabel m2contact 14337 4258 14337 4258 6 n_61
rlabel m2contact 14289 2434 14289 2434 6 n_190
rlabel m2contact 14265 3010 14265 3010 6 n_382
rlabel m2contact 14241 4354 14241 4354 6 OpcodeCondIn[3]
rlabel m2contact 14217 4114 14217 4114 6 n_150
rlabel m2contact 14193 7018 14193 7018 6 n_280
rlabel m2contact 14193 1930 14193 1930 6 n_280
rlabel m2contact 14169 2458 14169 2458 6 n_356
rlabel m2contact 14145 1882 14145 1882 6 n_71
rlabel m2contact 14145 7186 14145 7186 6 n_38
rlabel m2contact 14145 7162 14145 7162 6 n_180
rlabel m2contact 14145 2554 14145 2554 6 n_180
rlabel m2contact 14121 4114 14121 4114 6 n_150
rlabel m2contact 14121 4402 14121 4402 6 OpcodeCondIn[6]
rlabel m2contact 14097 3922 14097 3922 6 n_243
rlabel m2contact 14073 1930 14073 1930 6 n_280
rlabel m2contact 14073 2602 14073 2602 6 n_37
rlabel m2contact 14049 3250 14049 3250 6 OpcodeCondIn[4]
rlabel m2contact 14025 4138 14025 4138 6 stateSub[0]
rlabel m2contact 14001 6634 14001 6634 6 n_125
rlabel m2contact 14001 6586 14001 6586 6 n_209
rlabel m2contact 13977 4354 13977 4354 4 OpcodeCondIn[3]
rlabel m2contact 13953 6634 13953 6634 4 n_93
rlabel m2contact 13929 1906 13929 1906 4 n_236
rlabel m2contact 13929 5698 13929 5698 4 n_210
rlabel m2contact 13929 1930 13929 1930 4 n_210
rlabel m2contact 13905 7162 13905 7162 4 n_180
rlabel m2contact 13905 3706 13905 3706 4 n_183
rlabel m2contact 13881 1930 13881 1930 4 n_210
rlabel m2contact 13881 4978 13881 4978 4 n_160
rlabel m2contact 13857 3610 13857 3610 4 n_133
rlabel m2contact 13833 1954 13833 1954 4 ENB
rlabel m2contact 13809 2074 13809 2074 4 n_77
rlabel m2contact 13809 7138 13809 7138 4 PcSel[2]
rlabel m2contact 13785 4210 13785 4210 4 n_319
rlabel m2contact 13761 6370 13761 6370 4 n_197
rlabel m2contact 13737 3898 13737 3898 4 n_195
rlabel m2contact 13713 6010 13713 6010 4 n_196
rlabel m2contact 13713 5338 13713 5338 4 n_132
rlabel m2contact 13689 6370 13689 6370 4 n_294
rlabel m2contact 13689 2074 13689 2074 4 n_294
rlabel m2contact 13665 6370 13665 6370 4 n_294
rlabel m2contact 13665 5554 13665 5554 4 n_198
rlabel m2contact 13641 4066 13641 4066 4 OpcodeCondIn[5]
rlabel m2contact 13617 5794 13617 5794 4 n_292
rlabel m2contact 13593 3154 13593 3154 4 state[0]
rlabel m2contact 13593 3970 13593 3970 4 n_293
rlabel m2contact 13569 5770 13569 5770 4 n_141
rlabel m2contact 13569 4210 13569 4210 4 n_141
rlabel m2contact 13545 2314 13545 2314 4 n_340
rlabel m2contact 13521 2938 13521 2938 4 n_102
rlabel m2contact 13521 3178 13521 3178 4 n_62
rlabel m2contact 13497 4210 13497 4210 4 n_141
rlabel m2contact 13497 4714 13497 4714 4 n_104
rlabel m2contact 13473 4930 13473 4930 4 n_235
rlabel m2contact 13425 4666 13425 4666 4 n_14
rlabel m2contact 13425 2218 13425 2218 4 n_328
rlabel m2contact 13401 6346 13401 6346 4 n_128
rlabel m2contact 13401 1954 13401 1954 4 n_128
rlabel m2contact 13377 5866 13377 5866 4 n_325
rlabel m2contact 13377 5194 13377 5194 4 n_291
rlabel m2contact 13353 7162 13353 7162 4 n_246
rlabel m2contact 13353 2938 13353 2938 4 n_246
rlabel m2contact 13329 5794 13329 5794 4 n_15
rlabel m2contact 13305 6466 13305 6466 4 stateSub[1]
rlabel m2contact 13305 6370 13305 6370 4 n_97
rlabel m2contact 13281 1954 13281 1954 4 n_128
rlabel m2contact 13281 4162 13281 4162 4 n_182
rlabel m2contact 13257 7138 13257 7138 4 n_59
rlabel m2contact 13257 2674 13257 2674 4 n_59
rlabel m2contact 13233 7162 13233 7162 4 n_246
rlabel m2contact 13233 4666 13233 4666 4 n_23
rlabel m2contact 13209 5602 13209 5602 4 n_167
rlabel m2contact 13185 7138 13185 7138 4 n_59
rlabel m2contact 13185 4858 13185 4858 4 n_95
rlabel m2contact 13161 3490 13161 3490 4 n_187
rlabel m2contact 13113 7114 13113 7114 4 n_35
rlabel m2contact 13113 1978 13113 1978 4 Flags[3]
rlabel m2contact 13113 4882 13113 4882 4 n_365
rlabel m2contact 13113 4210 13113 4210 4 n_365
rlabel m2contact 13089 4210 13089 4210 4 n_365
rlabel m2contact 13089 4402 13089 4402 4 OpcodeCondIn[6]
rlabel m2contact 13065 7090 13065 7090 4 n_19
rlabel m2contact 13041 4210 13041 4210 4 nME
rlabel m2contact 13017 7066 13017 7066 4 n_222
rlabel m2contact 13017 5866 13017 5866 4 n_325
rlabel m2contact 12993 6874 12993 6874 4 n_80
rlabel m2contact 12969 7042 12969 7042 4 n_98
rlabel m2contact 12969 3610 12969 3610 4 n_133
rlabel m2contact 12945 6874 12945 6874 4 n_155
rlabel m2contact 12921 2002 12921 2002 4 n_225
rlabel m2contact 12873 4738 12873 4738 4 n_103
rlabel m2contact 12825 2026 12825 2026 4 CFlag
rlabel m2contact 12801 4450 12801 4450 4 n_205
rlabel m2contact 12777 3682 12777 3682 4 n_309
rlabel m2contact 12753 5338 12753 5338 4 n_132
rlabel m2contact 12729 6082 12729 6082 4 OpcodeCondIn[2]
rlabel m2contact 12729 4114 12729 4114 4 n_150
rlabel m2contact 12705 7018 12705 7018 4 n_280
rlabel m2contact 12705 5458 12705 5458 4 n_344
rlabel m2contact 12705 2026 12705 2026 4 n_344
rlabel m2contact 12681 5506 12681 5506 4 AluOR[0]
rlabel m2contact 12657 6994 12657 6994 4 n_8
rlabel m2contact 12657 4762 12657 4762 4 n_297
rlabel m2contact 12633 6466 12633 6466 4 stateSub[1]
rlabel m2contact 12633 5506 12633 5506 4 n_295
rlabel m2contact 12609 2026 12609 2026 4 n_344
rlabel m2contact 12609 4138 12609 4138 4 stateSub[0]
rlabel m2contact 12561 4186 12561 4186 4 PcEn
rlabel m2contact 12561 4954 12561 4954 4 n_161
rlabel m2contact 12537 6994 12537 6994 4 n_231
rlabel m2contact 12537 3562 12537 3562 4 n_231
rlabel m2contact 12513 2050 12513 2050 4 n_361
rlabel m2contact 12513 3154 12513 3154 4 state[0]
rlabel m2contact 12489 6994 12489 6994 4 n_231
rlabel m2contact 12489 4186 12489 4186 4 n_207
rlabel m2contact 12465 2962 12465 2962 4 n_254
rlabel m2contact 12417 2386 12417 2386 4 n_135
rlabel m2contact 12393 3778 12393 3778 4 n_266
rlabel m2contact 12369 5170 12369 5170 4 n_89
rlabel m2contact 12321 5170 12321 5170 4 n_29
rlabel m2contact 12297 4402 12297 4402 4 OpcodeCondIn[6]
rlabel m2contact 12273 2602 12273 2602 4 n_37
rlabel m2contact 12249 4450 12249 4450 4 n_205
rlabel m2contact 12201 6970 12201 6970 4 n_21
rlabel m2contact 12177 6298 12177 6298 4 n_154
rlabel m2contact 12153 6970 12153 6970 4 n_31
rlabel m2contact 12153 2962 12153 2962 4 n_31
rlabel m2contact 12129 6346 12129 6346 4 n_128
rlabel m2contact 12105 5266 12105 5266 4 OpcodeCondIn[1]
rlabel m2contact 12081 3298 12081 3298 4 n_159
rlabel m2contact 12081 5242 12081 5242 4 OpcodeCondIn[0]
rlabel m2contact 12057 3970 12057 3970 4 n_293
rlabel m2contact 12033 6970 12033 6970 4 n_31
rlabel m2contact 12033 5314 12033 5314 4 n_143
rlabel m2contact 11985 2866 11985 2866 4 n_66
rlabel m2contact 11985 6082 11985 6082 4 OpcodeCondIn[2]
rlabel m2contact 11961 4090 11961 4090 4 n_30
rlabel m2contact 11961 2698 11961 2698 4 OpcodeCondIn[7]
rlabel m2contact 11937 4546 11937 4546 4 n_186
rlabel m2contact 11889 3178 11889 3178 4 n_62
rlabel m2contact 11841 6202 11841 6202 4 n_44
rlabel m2contact 11793 2578 11793 2578 4 IntStatus
rlabel m2contact 11793 5986 11793 5986 4 n_60
rlabel m2contact 11769 2674 11769 2674 4 n_59
rlabel m2contact 11745 2578 11745 2578 4 n_26
rlabel m2contact 11697 6946 11697 6946 4 n_334
rlabel m2contact 11673 5986 11673 5986 4 n_224
rlabel m2contact 11649 2074 11649 2074 4 n_294
rlabel m2contact 11625 3082 11625 3082 4 n_223
rlabel m2contact 11601 6826 11601 6826 4 n_215
rlabel m2contact 11553 5866 11553 5866 4 n_325
rlabel m2contact 11529 4690 11529 4690 4 state[1]
rlabel m2contact 11505 3154 11505 3154 4 state[0]
rlabel m2contact 11433 5458 11433 5458 4 n_344
rlabel m2contact 11409 6826 11409 6826 4 n_285
rlabel m2contact 11385 5362 11385 5362 4 n_345
rlabel m2contact 11361 6922 11361 6922 4 n_118
rlabel m2contact 11361 4090 11361 4090 4 n_30
rlabel m2contact 11361 2074 11361 2074 4 n_30
rlabel m2contact 11337 5866 11337 5866 4 n_325
rlabel m2contact 11337 3082 11337 3082 4 n_325
rlabel m2contact 11313 3538 11313 3538 4 n_279
rlabel m2contact 11289 4402 11289 4402 4 OpcodeCondIn[6]
rlabel m2contact 11265 2410 11265 2410 4 n_248
rlabel m2contact 11241 3970 11241 3970 4 n_293
rlabel m2contact 11217 3034 11217 3034 4 n_226
rlabel m2contact 11193 3538 11193 3538 4 n_36
rlabel m2contact 11169 2074 11169 2074 4 n_30
rlabel m2contact 11169 3922 11169 3922 4 n_243
rlabel m2contact 11145 3034 11145 3034 4 n_22
rlabel m2contact 11121 5242 11121 5242 4 OpcodeCondIn[0]
rlabel m2contact 11097 2842 11097 2842 4 n_20
rlabel m2contact 11097 6658 11097 6658 4 n_234
rlabel m2contact 11073 3298 11073 3298 4 n_159
rlabel m2contact 11049 6658 11049 6658 4 n_181
rlabel m2contact 11025 3298 11025 3298 4 n_213
rlabel m2contact 11001 3082 11001 3082 4 n_325
rlabel m2contact 11001 4282 11001 4282 4 n_200
rlabel m2contact 10977 5770 10977 5770 4 n_141
rlabel m2contact 10953 4954 10953 4954 4 n_161
rlabel m2contact 10929 6298 10929 6298 4 n_154
rlabel m2contact 10929 4138 10929 4138 4 stateSub[0]
rlabel m2contact 10905 3346 10905 3346 4 n_146
rlabel m2contact 10881 6658 10881 6658 4 n_181
rlabel m2contact 10857 3418 10857 3418 4 n_193
rlabel m2contact 10857 4834 10857 4834 4 n_261
rlabel m2contact 10833 3706 10833 3706 4 n_183
rlabel m2contact 10809 6658 10809 6658 4 n_69
rlabel m2contact 10737 3346 10737 3346 4 n_134
rlabel m2contact 10713 3082 10713 3082 4 n_153
rlabel m2contact 10641 6850 10641 6850 4 n_138
rlabel m2contact 10617 5218 10617 5218 4 n_152
rlabel m2contact 10617 2074 10617 2074 4 n_152
rlabel m2contact 10593 2074 10593 2074 4 n_152
rlabel m2contact 10593 4522 10593 4522 4 n_137
rlabel m2contact 10569 6850 10569 6850 4 n_274
rlabel m2contact 10569 2842 10569 2842 4 n_274
rlabel m2contact 10545 3850 10545 3850 4 n_305
rlabel m2contact 10521 6898 10521 6898 4 n_178
rlabel m2contact 10521 3778 10521 3778 4 n_266
rlabel m2contact 10497 6850 10497 6850 4 n_274
rlabel m2contact 10497 3850 10497 3850 4 n_65
rlabel m2contact 10449 6874 10449 6874 4 n_155
rlabel m2contact 10449 6850 10449 6850 4 n_318
rlabel m2contact 10449 2338 10449 2338 4 n_318
rlabel m2contact 10425 2338 10425 2338 4 n_318
rlabel m2contact 10425 4978 10425 4978 4 n_160
rlabel m2contact 10401 6298 10401 6298 4 n_154
rlabel m2contact 10377 6850 10377 6850 4 n_318
rlabel m2contact 10377 5002 10377 5002 4 n_28
rlabel m2contact 10305 6826 10305 6826 4 n_285
rlabel m2contact 10305 5338 10305 5338 4 n_132
rlabel m2contact 10281 5626 10281 5626 4 n_163
rlabel m2contact 10257 2098 10257 2098 4 n_271
rlabel m2contact 10233 3130 10233 3130 4 n_10
rlabel m2contact 10209 3250 10209 3250 4 OpcodeCondIn[4]
rlabel m2contact 10185 2698 10185 2698 4 OpcodeCondIn[7]
rlabel m2contact 10185 3130 10185 3130 4 n_149
rlabel m2contact 10137 2458 10137 2458 4 n_356
rlabel m2contact 10089 3058 10089 3058 4 n_232
rlabel m2contact 10065 3226 10065 3226 4 n_333
rlabel m2contact 10065 5602 10065 5602 4 n_167
rlabel m2contact 10041 3058 10041 3058 4 n_240
rlabel m2contact 10017 5506 10017 5506 4 n_295
rlabel m2contact 9993 5554 9993 5554 4 n_198
rlabel m2contact 9969 4594 9969 4594 4 n_12
rlabel m2contact 9969 4450 9969 4450 4 n_205
rlabel m2contact 9945 5266 9945 5266 4 OpcodeCondIn[1]
rlabel m2contact 9945 4834 9945 4834 4 n_261
rlabel m2contact 9897 4402 9897 4402 4 OpcodeCondIn[6]
rlabel m2contact 9873 2698 9873 2698 4 OpcodeCondIn[7]
rlabel m2contact 9849 5818 9849 5818 4 stateSub[2]
rlabel m2contact 9825 3226 9825 3226 4 SysBus[0]
rlabel m2contact 9825 2098 9825 2098 4 SysBus[0]
rlabel m2contact 9801 2530 9801 2530 4 n_86
rlabel m2contact 9801 4594 9801 4594 4 n_311
rlabel m2contact 9777 3226 9777 3226 4 SysBus[0]
rlabel m2contact 9777 3154 9777 3154 4 state[0]
rlabel m2contact 9753 2338 9753 2338 4 n_318
rlabel m2contact 9753 3682 9753 3682 4 n_309
rlabel m2contact 9705 2098 9705 2098 4 SysBus[0]
rlabel m2contact 9705 2458 9705 2458 4 n_355
rlabel m2contact 9657 6802 9657 6802 4 n_276
rlabel m2contact 9657 3226 9657 3226 4 n_301
rlabel m2contact 9633 2122 9633 2122 4 n_347
rlabel m2contact 9609 2938 9609 2938 4 n_246
rlabel m2contact 9585 2146 9585 2146 4 n_250
rlabel m2contact 9585 2170 9585 2170 4 n_6
rlabel m2contact 9537 2842 9537 2842 4 n_274
rlabel m2contact 9537 4330 9537 4330 4 nWait
rlabel m2contact 9513 4690 9513 4690 4 state[1]
rlabel m2contact 9513 4354 9513 4354 4 OpcodeCondIn[3]
rlabel m2contact 9441 6778 9441 6778 4 n_144
rlabel m2contact 9441 2842 9441 2842 4 n_312
rlabel m2contact 9417 2218 9417 2218 4 n_328
rlabel m2contact 9393 6130 9393 6130 4 n_259
rlabel m2contact 9369 6754 9369 6754 4 n_27
rlabel m2contact 9369 5842 9369 5842 4 n_349
rlabel m2contact 9369 2218 9369 2218 4 n_349
rlabel m2contact 9345 3802 9345 3802 4 n_251
rlabel m2contact 9321 2194 9321 2194 4 n_171
rlabel m2contact 9321 4738 9321 4738 4 n_103
rlabel m2contact 9297 3394 9297 3394 4 n_169
rlabel m2contact 9273 2194 9273 2194 4 n_353
rlabel m2contact 9249 3634 9249 3634 4 Rs1Sel[0]
rlabel m2contact 9225 6730 9225 6730 4 n_11
rlabel m2contact 9225 5866 9225 5866 4 n_325
rlabel m2contact 9201 2194 9201 2194 4 n_353
rlabel m2contact 9201 3394 9201 3394 4 n_320
rlabel m2contact 9177 6706 9177 6706 4 n_217
rlabel m2contact 9153 2218 9153 2218 4 n_349
rlabel m2contact 9153 3634 9153 3634 4 n_247
rlabel m2contact 9105 2626 9105 2626 4 n_123
rlabel m2contact 9105 3778 9105 3778 4 n_266
rlabel m2contact 9081 2938 9081 2938 4 n_246
rlabel m2contact 9057 6706 9057 6706 4 n_67
rlabel m2contact 9057 2626 9057 2626 4 n_67
rlabel m2contact 9033 6706 9033 6706 4 n_67
rlabel m2contact 9033 2938 9033 2938 4 n_9
rlabel m2contact 9009 3778 9009 3778 4 n_266
rlabel m2contact 8985 2242 8985 2242 4 n_105
rlabel m2contact 8985 2866 8985 2866 4 n_66
rlabel m2contact 8961 6682 8961 6682 4 n_24
rlabel m2contact 8961 4738 8961 4738 4 n_103
rlabel m2contact 8937 4714 8937 4714 4 n_104
rlabel m2contact 8913 6658 8913 6658 4 n_69
rlabel m2contact 8913 5554 8913 5554 4 n_198
rlabel m2contact 8913 2242 8913 2242 4 n_198
rlabel m2contact 8889 3058 8889 3058 4 n_240
rlabel m2contact 8889 4402 8889 4402 4 OpcodeCondIn[6]
rlabel m2contact 8865 3778 8865 3778 4 n_266
rlabel m2contact 8841 2242 8841 2242 4 n_198
rlabel m2contact 8841 5338 8841 5338 4 n_132
rlabel m2contact 8817 2434 8817 2434 4 n_190
rlabel m2contact 8817 3250 8817 3250 4 OpcodeCondIn[4]
rlabel m2contact 8769 6634 8769 6634 4 n_93
rlabel m2contact 8745 3370 8745 3370 4 n_92
rlabel m2contact 8721 6466 8721 6466 4 stateSub[1]
rlabel m2contact 8721 3802 8721 3802 4 n_251
rlabel m2contact 8697 5674 8697 5674 4 n_68
rlabel m2contact 8673 2266 8673 2266 4 n_5
rlabel m2contact 8649 2698 8649 2698 4 OpcodeCondIn[7]
rlabel m2contact 8625 3778 8625 3778 4 n_266
rlabel m2contact 8625 4138 8625 4138 4 stateSub[0]
rlabel m2contact 8577 6610 8577 6610 4 n_136
rlabel m2contact 8577 4066 8577 4066 4 OpcodeCondIn[5]
rlabel m2contact 8553 2386 8553 2386 4 n_135
rlabel m2contact 8529 2290 8529 2290 4 PcSel[0]
rlabel m2contact 8529 6298 8529 6298 4 n_154
rlabel m2contact 8505 2314 8505 2314 4 n_340
rlabel m2contact 8505 2338 8505 2338 4 n_318
rlabel m2contact 8481 6298 8481 6298 4 n_290
rlabel m2contact 8457 6586 8457 6586 4 n_209
rlabel m2contact 8433 6082 8433 6082 4 OpcodeCondIn[2]
rlabel m2contact 8433 2338 8433 2338 4 OpcodeCondIn[2]
rlabel m2contact 8409 2338 8409 2338 4 OpcodeCondIn[2]
rlabel m2contact 8409 5626 8409 5626 4 n_163
rlabel m2contact 8385 2362 8385 2362 4 n_400
rlabel m2contact 8385 5410 8385 5410 4 n_164
rlabel m2contact 8361 4090 8361 4090 4 n_30
rlabel m2contact 8313 4090 8313 4090 4 n_174
rlabel m2contact 8289 2386 8289 2386 4 n_135
rlabel m2contact 8289 4330 8289 4330 4 nWait
rlabel m2contact 8265 6562 8265 6562 4 n_78
rlabel m2contact 8241 3154 8241 3154 4 state[0]
rlabel m2contact 8217 6538 8217 6538 4 n_64
rlabel m2contact 8217 6466 8217 6466 4 stateSub[1]
rlabel m2contact 8193 3778 8193 3778 4 n_266
rlabel m2contact 8169 4666 8169 4666 4 n_23
rlabel m2contact 8145 4858 8145 4858 4 n_95
rlabel m2contact 8121 4666 8121 4666 4 n_90
rlabel m2contact 8097 3250 8097 3250 4 OpcodeCondIn[4]
rlabel m2contact 8097 4690 8097 4690 4 state[1]
rlabel m2contact 8073 5026 8073 5026 4 n_88
rlabel m2contact 8049 2410 8049 2410 4 n_248
rlabel m2contact 8025 2602 8025 2602 4 n_37
rlabel m2contact 8001 4858 8001 4858 4 n_95
rlabel m2contact 7977 2434 7977 2434 4 n_190
rlabel m2contact 7977 2698 7977 2698 4 OpcodeCondIn[7]
rlabel m2contact 7953 4066 7953 4066 4 OpcodeCondIn[5]
rlabel m2contact 7929 4258 7929 4258 4 n_61
rlabel m2contact 7905 5674 7905 5674 4 n_68
rlabel m2contact 7905 2434 7905 2434 4 n_68
rlabel m2contact 7881 2434 7881 2434 4 n_68
rlabel m2contact 7881 5338 7881 5338 4 n_132
rlabel m2contact 7857 4930 7857 4930 4 n_235
rlabel m2contact 7833 2674 7833 2674 4 n_59
rlabel m2contact 7809 6514 7809 6514 4 n_368
rlabel m2contact 7785 6490 7785 6490 4 n_170
rlabel m2contact 7761 6466 7761 6466 4 stateSub[1]
rlabel m2contact 7737 2458 7737 2458 4 n_355
rlabel m2contact 7737 2482 7737 2482 4 n_124
rlabel m2contact 7689 4306 7689 4306 4 n_117
rlabel m2contact 7665 4714 7665 4714 4 n_104
rlabel m2contact 7641 3610 7641 3610 4 n_133
rlabel m2contact 7617 5026 7617 5026 4 n_88
rlabel m2contact 7617 4954 7617 4954 4 n_161
rlabel m2contact 7593 5458 7593 5458 4 n_344
rlabel m2contact 7593 2482 7593 2482 4 n_344
rlabel m2contact 7569 4306 7569 4306 4 nOE
rlabel m2contact 7545 2482 7545 2482 4 n_344
rlabel m2contact 7545 5026 7545 5026 4 n_47
rlabel m2contact 7521 2506 7521 2506 4 n_199
rlabel m2contact 7521 6442 7521 6442 4 n_300
rlabel m2contact 7497 6274 7497 6274 4 n_323
rlabel m2contact 7473 4618 7473 4618 4 n_244
rlabel m2contact 7449 4882 7449 4882 4 n_365
rlabel m2contact 7425 2530 7425 2530 4 n_86
rlabel m2contact 7425 6418 7425 6418 4 n_151
rlabel m2contact 7401 2554 7401 2554 4 n_180
rlabel m2contact 7401 6250 7401 6250 4 n_321
rlabel m2contact 7377 6394 7377 6394 4 n_256
rlabel m2contact 7353 2578 7353 2578 4 n_26
rlabel m2contact 7353 6250 7353 6250 4 n_188
rlabel m2contact 7305 6370 7305 6370 4 n_97
rlabel m2contact 7305 3466 7305 3466 4 n_25
rlabel m2contact 7281 2602 7281 2602 4 n_37
rlabel m2contact 7281 2626 7281 2626 4 n_67
rlabel m2contact 7257 4162 7257 4162 4 n_182
rlabel m2contact 7233 5266 7233 5266 4 OpcodeCondIn[1]
rlabel m2contact 7233 2626 7233 2626 4 OpcodeCondIn[1]
rlabel m2contact 7209 2626 7209 2626 4 OpcodeCondIn[1]
rlabel m2contact 7209 4570 7209 4570 4 n_371
rlabel m2contact 7185 6346 7185 6346 4 n_128
rlabel m2contact 7185 5242 7185 5242 4 OpcodeCondIn[0]
rlabel m2contact 7161 2650 7161 2650 4 n_322
rlabel m2contact 7137 2674 7137 2674 4 n_59
rlabel m2contact 7137 3898 7137 3898 4 n_195
rlabel m2contact 7113 4354 7113 4354 4 OpcodeCondIn[3]
rlabel m2contact 7089 2698 7089 2698 4 OpcodeCondIn[7]
rlabel m2contact 7089 6322 7089 6322 4 n_262
rlabel m2contact 7065 4834 7065 4834 4 n_261
rlabel m2contact 7041 3034 7041 3034 4 n_22
rlabel m2contact 7041 3058 7041 3058 4 n_240
rlabel m2contact 7017 3970 7017 3970 4 n_293
rlabel m2contact 6993 6298 6993 6298 4 n_290
rlabel m2contact 6993 4138 6993 4138 4 stateSub[0]
rlabel m2contact 6969 5194 6969 5194 4 n_291
rlabel m2contact 6945 2722 6945 2722 4 n_302
rlabel m2contact 6945 2746 6945 2746 4 n_166
rlabel m2contact 6897 6274 6897 6274 4 n_323
rlabel m2contact 6897 4066 6897 4066 4 OpcodeCondIn[5]
rlabel m2contact 6873 2770 6873 2770 4 n_242
rlabel m2contact 6873 3562 6873 3562 4 n_231
rlabel m2contact 6849 2818 6849 2818 4 n_202
rlabel m2contact 6801 2794 6801 2794 4 n_100
rlabel m2contact 6801 2818 6801 2818 4 n_348
rlabel m2contact 6777 2818 6777 2818 4 n_348
rlabel m2contact 6777 3154 6777 3154 4 state[0]
rlabel m2contact 6753 2842 6753 2842 4 n_312
rlabel m2contact 6729 6250 6729 6250 4 n_188
rlabel m2contact 6705 6226 6705 6226 4 n_45
rlabel m2contact 6705 4546 6705 4546 4 n_186
rlabel m2contact 6681 6202 6681 6202 4 n_44
rlabel m2contact 6681 3490 6681 3490 4 n_187
rlabel m2contact 6657 4258 6657 4258 4 n_61
rlabel m2contact 6609 6178 6609 6178 4 n_227
rlabel m2contact 6609 4138 6609 4138 4 stateSub[0]
rlabel m2contact 6585 6154 6585 6154 4 n_176
rlabel m2contact 6561 6130 6561 6130 4 n_259
rlabel m2contact 6513 4474 6513 4474 4 n_204
rlabel m2contact 6489 2866 6489 2866 4 n_66
rlabel m2contact 6489 4474 6489 4474 4 n_204
rlabel m2contact 6441 3010 6441 3010 4 n_382
rlabel m2contact 6441 3754 6441 3754 4 n_56
rlabel m2contact 6393 2890 6393 2890 4 n_317
rlabel m2contact 6369 6106 6369 6106 4 n_177
rlabel m2contact 6369 3010 6369 3010 4 n_369
rlabel m2contact 6345 2914 6345 2914 4 n_268
rlabel m2contact 6297 2938 6297 2938 4 n_9
rlabel m2contact 6273 2962 6273 2962 4 n_31
rlabel m2contact 6273 6082 6273 6082 4 OpcodeCondIn[2]
rlabel m2contact 6249 4138 6249 4138 4 stateSub[0]
rlabel m2contact 6201 2986 6201 2986 4 n_32
rlabel m2contact 6201 3010 6201 3010 4 n_369
rlabel m2contact 6177 6058 6177 6058 4 StatusReg[3]
rlabel m2contact 6177 4402 6177 4402 4 OpcodeCondIn[6]
rlabel m2contact 6153 3778 6153 3778 4 n_266
rlabel m2contact 6153 4570 6153 4570 4 n_371
rlabel m2contact 6129 5338 6129 5338 4 n_132
rlabel m2contact 6105 3730 6105 3730 4 n_130
rlabel m2contact 6081 4354 6081 4354 4 OpcodeCondIn[3]
rlabel m2contact 6057 5314 6057 5314 4 n_143
rlabel m2contact 6057 4378 6057 4378 4 n_74
rlabel m2contact 6009 3034 6009 3034 4 n_22
rlabel m2contact 6009 6034 6009 6034 4 n_208
rlabel m2contact 5985 5698 5985 5698 4 n_210
rlabel m2contact 5961 6010 5961 6010 4 n_196
rlabel m2contact 5937 3970 5937 3970 4 n_293
rlabel m2contact 5913 3058 5913 3058 4 n_240
rlabel m2contact 5913 5986 5913 5986 4 n_224
rlabel m2contact 5889 5962 5889 5962 4 n_157
rlabel m2contact 5865 3082 5865 3082 4 n_153
rlabel m2contact 5865 4114 5865 4114 4 n_150
rlabel m2contact 5841 4834 5841 4834 4 n_261
rlabel m2contact 5817 5938 5817 5938 4 n_111
rlabel m2contact 5817 5410 5817 5410 4 n_164
rlabel m2contact 5793 5914 5793 5914 4 n_156
rlabel m2contact 5793 5314 5793 5314 4 n_143
rlabel m2contact 5769 3106 5769 3106 4 n_34
rlabel m2contact 5721 5890 5721 5890 4 n_50
rlabel m2contact 5721 4474 5721 4474 4 n_204
rlabel m2contact 5697 3130 5697 3130 4 n_149
rlabel m2contact 5697 5866 5697 5866 4 n_325
rlabel m2contact 5673 3610 5673 3610 4 n_133
rlabel m2contact 5625 3154 5625 3154 4 state[0]
rlabel m2contact 5625 3586 5625 3586 4 n_332
rlabel m2contact 5601 3178 5601 3178 4 n_62
rlabel m2contact 5577 3586 5577 3586 4 n_115
rlabel m2contact 5553 3202 5553 3202 4 n_84
rlabel m2contact 5553 3226 5553 3226 4 n_301
rlabel m2contact 5529 3250 5529 3250 4 OpcodeCondIn[4]
rlabel m2contact 5505 5842 5505 5842 4 n_349
rlabel m2contact 5481 5818 5481 5818 4 stateSub[2]
rlabel m2contact 5457 5794 5457 5794 4 n_15
rlabel m2contact 5409 4978 5409 4978 4 n_160
rlabel m2contact 5361 3274 5361 3274 4 StatusReg[2]
rlabel m2contact 5361 4546 5361 4546 4 n_186
rlabel m2contact 5337 5770 5337 5770 4 n_141
rlabel m2contact 5289 5074 5289 5074 4 n_287
rlabel m2contact 5265 3562 5265 3562 4 n_231
rlabel m2contact 5241 5074 5241 5074 4 n_239
rlabel m2contact 5193 3298 5193 3298 4 n_213
rlabel m2contact 5169 3418 5169 3418 4 n_193
rlabel m2contact 5145 3802 5145 3802 4 n_251
rlabel m2contact 5097 3418 5097 3418 4 n_114
rlabel m2contact 5073 3802 5073 3802 4 n_251
rlabel m2contact 5049 5746 5049 5746 4 n_85
rlabel m2contact 5001 3322 5001 3322 4 n_148
rlabel m2contact 4953 5578 4953 5578 4 n_147
rlabel m2contact 4929 5722 4929 5722 4 n_127
rlabel m2contact 4881 3346 4881 3346 4 n_134
rlabel m2contact 4857 4978 4857 4978 4 n_160
rlabel m2contact 4833 4930 4833 4930 4 n_235
rlabel m2contact 4785 5698 4785 5698 4 n_210
rlabel m2contact 4737 4690 4737 4690 4 state[1]
rlabel m2contact 4713 3370 4713 3370 4 n_92
rlabel m2contact 4713 5674 4713 5674 4 n_68
rlabel m2contact 4665 5602 4665 5602 4 n_167
rlabel m2contact 4641 5650 4641 5650 4 n_158
rlabel m2contact 4641 4834 4641 4834 4 n_261
rlabel m2contact 4593 3394 4593 3394 4 n_320
rlabel m2contact 4593 4642 4593 4642 4 n_13
rlabel m2contact 4569 4234 4569 4234 4 n_52
rlabel m2contact 4545 5626 4545 5626 4 n_163
rlabel m2contact 4521 4234 4521 4234 4 n_75
rlabel m2contact 4497 3418 4497 3418 4 n_114
rlabel m2contact 4497 5602 4497 5602 4 n_167
rlabel m2contact 4473 5314 4473 5314 4 n_143
rlabel m2contact 4425 5578 4425 5578 4 n_147
rlabel m2contact 4425 4786 4425 4786 4 n_257
rlabel m2contact 4377 3922 4377 3922 4 n_243
rlabel m2contact 4353 5554 4353 5554 4 n_198
rlabel m2contact 4305 3442 4305 3442 4 n_120
rlabel m2contact 4281 5314 4281 5314 4 n_143
rlabel m2contact 4281 3682 4281 3682 4 n_309
rlabel m2contact 4257 4954 4257 4954 4 n_161
rlabel m2contact 4233 5530 4233 5530 4 n_173
rlabel m2contact 4185 3466 4185 3466 4 n_25
rlabel m2contact 4185 4762 4185 4762 4 n_297
rlabel m2contact 4161 3490 4161 3490 4 n_187
rlabel m2contact 4161 5506 4161 5506 4 n_295
rlabel m2contact 4137 5482 4137 5482 4 n_298
rlabel m2contact 4113 5458 4113 5458 4 n_344
rlabel m2contact 4089 5434 4089 5434 4 n_221
rlabel m2contact 4065 5410 4065 5410 4 n_164
rlabel m2contact 4041 3946 4041 3946 4 n_255
rlabel m2contact 4017 5338 4017 5338 4 n_132
rlabel m2contact 3993 3514 3993 3514 4 n_81
rlabel m2contact 3993 3898 3993 3898 4 n_195
rlabel m2contact 3969 4474 3969 4474 4 n_204
rlabel m2contact 3945 3538 3945 3538 4 n_36
rlabel m2contact 3945 5362 3945 5362 4 n_345
rlabel m2contact 3897 5362 3897 5362 4 n_126
rlabel m2contact 3873 5386 3873 5386 4 n_168
rlabel m2contact 3873 4930 3873 4930 4 n_235
rlabel m2contact 3849 3562 3849 3562 4 n_231
rlabel m2contact 3825 5362 3825 5362 4 n_126
rlabel m2contact 3801 3586 3801 3586 4 n_115
rlabel m2contact 3801 5338 3801 5338 4 n_132
rlabel m2contact 3777 4954 3777 4954 4 n_161
rlabel m2contact 3777 4330 3777 4330 4 nWait
rlabel m2contact 3753 5314 3753 5314 4 n_143
rlabel m2contact 3753 3898 3753 3898 4 n_195
rlabel m2contact 3729 3610 3729 3610 4 n_133
rlabel m2contact 3705 5290 3705 5290 4 n_192
rlabel m2contact 3681 4426 3681 4426 4 n_206
rlabel m2contact 3657 4450 3657 4450 4 n_205
rlabel m2contact 3609 3634 3609 3634 4 n_247
rlabel m2contact 3609 3658 3609 3658 4 n_16
rlabel m2contact 3585 5266 3585 5266 4 OpcodeCondIn[1]
rlabel m2contact 3537 5242 3537 5242 4 OpcodeCondIn[0]
rlabel m2contact 3513 3682 3513 3682 4 n_309
rlabel m2contact 3489 5218 3489 5218 4 n_152
rlabel m2contact 3465 4354 3465 4354 4 OpcodeCondIn[3]
rlabel m2contact 3441 3706 3441 3706 4 n_183
rlabel m2contact 3441 3898 3441 3898 4 n_195
rlabel m2contact 3417 4978 3417 4978 4 n_160
rlabel m2contact 3393 3730 3393 3730 4 n_130
rlabel m2contact 3369 5194 3369 5194 4 n_291
rlabel m2contact 3345 3754 3345 3754 4 n_56
rlabel m2contact 3321 5170 3321 5170 4 n_29
rlabel m2contact 3321 4858 3321 4858 4 n_95
rlabel m2contact 3297 3778 3297 3778 4 n_266
rlabel m2contact 3297 5146 3297 5146 4 n_238
rlabel m2contact 3249 5122 3249 5122 4 n_381
rlabel m2contact 3225 4594 3225 4594 4 n_311
rlabel m2contact 3201 5098 3201 5098 4 n_367
rlabel m2contact 3177 4594 3177 4594 4 n_376
rlabel m2contact 3153 4690 3153 4690 4 state[1]
rlabel m2contact 3129 5074 3129 5074 4 n_239
rlabel m2contact 3105 3802 3105 3802 4 n_251
rlabel m2contact 3105 3826 3105 3826 4 n_99
rlabel m2contact 3081 5050 3081 5050 4 n_184
rlabel m2contact 3033 5026 3033 5026 4 n_47
rlabel m2contact 3009 5002 3009 5002 4 n_28
rlabel m2contact 2985 4258 2985 4258 4 n_61
rlabel m2contact 2937 4258 2937 4258 4 n_162
rlabel m2contact 2913 4978 2913 4978 4 n_160
rlabel m2contact 2889 4954 2889 4954 4 n_161
rlabel m2contact 2865 4930 2865 4930 4 n_235
rlabel m2contact 2817 4906 2817 4906 4 n_366
rlabel m2contact 2793 3994 2793 3994 4 Flags[1]
rlabel m2contact 2769 4882 2769 4882 4 n_365
rlabel m2contact 2745 3994 2745 3994 4 n_282
rlabel m2contact 2721 3850 2721 3850 4 n_65
rlabel m2contact 2697 4858 2697 4858 4 n_95
rlabel m2contact 2673 4834 2673 4834 4 n_261
rlabel m2contact 2625 4810 2625 4810 4 n_258
rlabel m2contact 2625 4114 2625 4114 4 n_150
rlabel m2contact 2601 4138 2601 4138 4 stateSub[0]
rlabel m2contact 2577 3874 2577 3874 4 n_101
rlabel m2contact 2577 4786 2577 4786 4 n_257
rlabel m2contact 2553 3898 2553 3898 4 n_195
rlabel m2contact 2529 4762 2529 4762 4 n_297
rlabel m2contact 2505 4738 2505 4738 4 n_103
rlabel m2contact 2481 3922 2481 3922 4 n_243
rlabel m2contact 2481 4714 2481 4714 4 n_104
rlabel m2contact 2457 3946 2457 3946 4 n_255
rlabel m2contact 2457 4690 2457 4690 4 state[1]
rlabel m2contact 2433 3970 2433 3970 4 n_293
rlabel m2contact 2409 3994 2409 3994 4 n_282
rlabel m2contact 2385 4018 2385 4018 4 n_189
rlabel m2contact 2385 4042 2385 4042 4 n_17
rlabel m2contact 2361 4066 2361 4066 4 OpcodeCondIn[5]
rlabel m2contact 2361 4090 2361 4090 4 n_174
rlabel m2contact 2337 4114 2337 4114 4 n_150
rlabel m2contact 2337 4666 2337 4666 4 n_90
rlabel m2contact 2241 4642 2241 4642 4 n_13
rlabel m2contact 2217 4618 2217 4618 4 n_244
rlabel m2contact 2193 4138 2193 4138 4 stateSub[0]
rlabel m2contact 2169 4594 2169 4594 4 n_376
rlabel m2contact 2145 4162 2145 4162 4 n_182
rlabel m2contact 2121 4570 2121 4570 4 n_371
rlabel m2contact 2049 4546 2049 4546 4 n_186
rlabel m2contact 2001 4402 2001 4402 4 OpcodeCondIn[6]
rlabel m2contact 1953 4522 1953 4522 4 n_137
rlabel m2contact 1929 4354 1929 4354 4 OpcodeCondIn[3]
rlabel m2contact 1905 4498 1905 4498 4 n_91
rlabel m2contact 1857 4186 1857 4186 4 n_207
rlabel m2contact 1833 4474 1833 4474 4 n_204
rlabel m2contact 1809 4450 1809 4450 4 n_205
rlabel m2contact 1785 4426 1785 4426 4 n_206
rlabel m2contact 1737 4210 1737 4210 4 nME
rlabel m2contact 1689 4234 1689 4234 4 n_75
rlabel m2contact 1665 4402 1665 4402 4 OpcodeCondIn[6]
rlabel m2contact 1641 4258 1641 4258 4 n_162
rlabel m2contact 1641 4378 1641 4378 4 n_74
rlabel m2contact 1617 4282 1617 4282 4 n_200
rlabel m2contact 1617 4354 1617 4354 4 OpcodeCondIn[3]
rlabel m2contact 27129 8187 27129 8187 6 RwSel[1]
rlabel m2contact 27129 8067 27129 8067 6 RwSel[1]
rlabel m2contact 27105 8163 27105 8163 6 ENB
rlabel m2contact 27105 8067 27105 8067 6 ENB
rlabel m2contact 27081 8235 27081 8235 6 AluOR[1]
rlabel m2contact 27081 8139 27081 8139 6 AluOR[1]
rlabel m2contact 27057 8259 27057 8259 6 AluOR[0]
rlabel m2contact 27057 8115 27057 8115 6 AluOR[0]
rlabel m2contact 27033 8259 27033 8259 6 AluOR[0]
rlabel m2contact 26133 8259 26133 8259 6 StatusRegEn
rlabel m2contact 25785 8211 25785 8211 6 ImmSel
rlabel m2contact 25293 8307 25293 8307 6 StatusReg[0]
rlabel m2contact 25017 8331 25017 8331 6 StatusReg[2]
rlabel m2contact 24801 8187 24801 8187 6 RwSel[1]
rlabel m2contact 24453 8283 24453 8283 6 StatusReg[1]
rlabel m2contact 24429 8331 24429 8331 6 StatusReg[2]
rlabel m2contact 24153 8139 24153 8139 6 LrWe
rlabel m2contact 23409 8115 23409 8115 6 PcSel[1]
rlabel m2contact 23145 8355 23145 8355 6 ALE
rlabel m2contact 22773 8403 22773 8403 6 StatusReg[3]
rlabel metal2 22419 8187 22419 8187 6 AluEn
rlabel m2contact 22401 8187 22401 8187 6 AluEn
rlabel m2contact 22161 8331 22161 8331 6 AluWe
rlabel m2contact 22017 8307 22017 8307 6 StatusReg[0]
rlabel m2contact 21909 8331 21909 8331 6 AluWe
rlabel m2contact 20937 8163 20937 8163 6 LrSel
rlabel metal2 20715 8187 20715 8187 6 Op2Sel[0]
rlabel m2contact 20697 8187 20697 8187 6 Op2Sel[0]
rlabel m2contact 20553 8331 20553 8331 6 Op1Sel
rlabel m2contact 20289 8427 20289 8427 6 PcWe
rlabel m2contact 19425 8067 19425 8067 6 ENB
rlabel m2contact 19413 8187 19413 8187 6 Op2Sel[1]
rlabel m2contact 19389 8331 19389 8331 6 Op1Sel
rlabel m2contact 19161 8331 19161 8331 6 MemEn
rlabel m2contact 18657 8091 18657 8091 6 RegWe
rlabel m2contact 17733 8379 17733 8379 6 WdSel
rlabel metal2 17727 8091 17727 8091 6 PcEn
rlabel m2contact 17709 8091 17709 8091 6 PcEn
rlabel m2contact 16869 8427 16869 8427 6 PcWe
rlabel metal2 15723 8427 15723 8427 6 PcSel[0]
rlabel m2contact 15705 8427 15705 8427 6 PcSel[0]
rlabel m2contact 15189 8115 15189 8115 6 PcSel[1]
rlabel m2contact 14673 8403 14673 8403 6 StatusReg[3]
rlabel metal2 13827 8403 13827 8403 4 PcSel[2]
rlabel m2contact 13809 8403 13809 8403 4 PcSel[2]
rlabel m2contact 12873 8283 12873 8283 4 StatusReg[1]
rlabel m2contact 12681 8283 12681 8283 4 LrEn
rlabel m2contact 12645 8139 12645 8139 4 LrWe
rlabel m2contact 11793 8163 11793 8163 4 LrSel
rlabel m2contact 11457 8187 11457 8187 4 Op2Sel[1]
rlabel m2contact 10941 8211 10941 8211 4 ImmSel
rlabel m2contact 10761 8259 10761 8259 4 StatusRegEn
rlabel m2contact 9945 8187 9945 8187 4 OpcodeCondIn[1]
rlabel m2contact 9465 8283 9465 8283 4 LrEn
rlabel m2contact 9273 8283 9273 8283 4 IrWe
rlabel m2contact 9237 8331 9237 8331 4 MemEn
rlabel m2contact 8817 8211 8817 8211 4 OpcodeCondIn[4]
rlabel m2contact 8337 8283 8337 8283 4 IrWe
rlabel m2contact 7977 8283 7977 8283 4 OpcodeCondIn[7]
rlabel m2contact 7953 8259 7953 8259 4 OpcodeCondIn[5]
rlabel m2contact 7569 8331 7569 8331 4 OpcodeCondIn[0]
rlabel m2contact 7533 8187 7533 8187 4 OpcodeCondIn[1]
rlabel metal2 6291 8187 6291 8187 4 OpcodeCondIn[2]
rlabel m2contact 6273 8187 6273 8187 4 OpcodeCondIn[2]
rlabel m2contact 6081 8187 6081 8187 4 OpcodeCondIn[3]
rlabel m2contact 5829 8187 5829 8187 4 OpcodeCondIn[3]
rlabel m2contact 4977 8211 4977 8211 4 OpcodeCondIn[4]
rlabel m2contact 4209 8235 4209 8235 4 AluOR[1]
rlabel m2contact 4125 8259 4125 8259 4 OpcodeCondIn[5]
rlabel m2contact 3561 8307 3561 8307 4 StatusReg[0]
rlabel m2contact 3537 8331 3537 8331 4 OpcodeCondIn[0]
rlabel m2contact 2457 8331 2457 8331 4 OpcodeCondIn[6]
rlabel m2contact 2421 8283 2421 8283 4 OpcodeCondIn[7]
rlabel m2contact 2289 8379 2289 8379 4 WdSel
rlabel m2contact 2145 8307 2145 8307 4 StatusReg[0]
rlabel m2contact 2001 8331 2001 8331 4 OpcodeCondIn[6]
rlabel m2contact 1737 8331 1737 8331 4 nME
rlabel m2contact 26601 569 26601 569 8 CFlag
rlabel m2contact 26601 17 26601 17 8 CFlag
rlabel m2contact 26577 65 26577 65 8 Flags[1]
rlabel m2contact 26577 41 26577 41 8 Flags[0]
rlabel m2contact 26577 17 26577 17 8 Flags[0]
rlabel metal2 26577 545 26577 545 8 Flags[1]
rlabel m2contact 26457 905 26457 905 6 n_316
rlabel m2contact 26385 665 26385 665 8 n_265
rlabel m2contact 26289 761 26289 761 8 n_281
rlabel m2contact 26145 545 26145 545 8 n_113
rlabel m2contact 26121 737 26121 737 8 n_43
rlabel m2contact 26049 281 26049 281 8 n_378
rlabel m2contact 26025 305 26025 305 8 n_308
rlabel m2contact 26001 41 26001 41 8 n_364
rlabel m2contact 25425 617 25425 617 8 n_362
rlabel m2contact 25281 977 25281 977 6 n_112
rlabel m2contact 24681 401 24681 401 8 n_354
rlabel m2contact 24561 689 24561 689 8 n_278
rlabel m2contact 24513 329 24513 329 8 n_230
rlabel m2contact 24465 809 24465 809 6 n_145
rlabel m2contact 24369 641 24369 641 8 n_58
rlabel m2contact 24249 353 24249 353 8 n_275
rlabel m2contact 24201 497 24201 497 8 n_241
rlabel m2contact 24105 713 24105 713 8 n_107
rlabel m2contact 23505 593 23505 593 8 n_335
rlabel m2contact 23241 209 23241 209 8 n_87
rlabel m2contact 23001 761 23001 761 8 n_281
rlabel m2contact 22833 161 22833 161 8 n_401
rlabel m2contact 22737 233 22737 233 8 SysBus[1]
rlabel m2contact 22665 425 22665 425 8 n_49
rlabel m2contact 22065 209 22065 209 8 n_87
rlabel m2contact 21945 833 21945 833 6 n_351
rlabel m2contact 21753 881 21753 881 6 n_131
rlabel m2contact 21705 377 21705 377 8 n_306
rlabel m2contact 21633 113 21633 113 8 nWE
rlabel m2contact 21585 689 21585 689 8 n_278
rlabel m2contact 21513 689 21513 689 8 n_216
rlabel m2contact 21417 617 21417 617 8 n_362
rlabel m2contact 21369 593 21369 593 8 n_335
rlabel m2contact 21321 449 21321 449 8 n_53
rlabel m2contact 20937 473 20937 473 8 n_218
rlabel m2contact 20889 185 20889 185 8 n_272
rlabel m2contact 20697 65 20697 65 8 SysBus[3]
rlabel m2contact 20577 569 20577 569 8 CFlag
rlabel m2contact 20529 569 20529 569 8 n_42
rlabel m2contact 20073 617 20073 617 8 n_245
rlabel m2contact 19785 593 19785 593 8 n_82
rlabel m2contact 19737 569 19737 569 8 n_42
rlabel m2contact 19665 641 19665 641 8 n_58
rlabel m2contact 19593 569 19593 569 8 n_273
rlabel m2contact 19545 761 19545 761 8 n_211
rlabel m2contact 19473 617 19473 617 8 n_245
rlabel m2contact 19425 257 19425 257 8 n_304
rlabel m2contact 19401 857 19401 857 6 n_237
rlabel m2contact 19353 785 19353 785 8 n_33
rlabel m2contact 19185 617 19185 617 8 n_4
rlabel m2contact 19017 905 19017 905 6 n_316
rlabel m2contact 18969 929 18969 929 6 n_269
rlabel m2contact 18825 137 18825 137 8 IRQ1
rlabel m2contact 18417 89 18417 89 8 n_3
rlabel m2contact 18297 1001 18297 1001 6 n_70
rlabel m2contact 18153 953 18153 953 6 n_284
rlabel m2contact 18105 905 18105 905 6 n_229
rlabel m2contact 18081 1001 18081 1001 6 n_70
rlabel m2contact 18057 977 18057 977 6 n_112
rlabel m2contact 17985 89 17985 89 8 n_3
rlabel m2contact 17937 89 17937 89 8 nIRQ
rlabel m2contact 17889 17 17889 17 8 Flags[0]
rlabel m2contact 17817 353 17817 353 8 n_275
rlabel m2contact 17577 953 17577 953 6 n_284
rlabel m2contact 17289 41 17289 41 8 n_364
rlabel m2contact 17265 521 17265 521 8 Flags[2]
rlabel m2contact 16689 521 16689 521 8 n_79
rlabel m2contact 16473 881 16473 881 6 n_131
rlabel m2contact 16329 41 16329 41 8 n_336
rlabel m2contact 16233 881 16233 881 6 n_119
rlabel m2contact 16137 41 16137 41 8 n_336
rlabel m2contact 16017 857 16017 857 6 n_237
rlabel m2contact 15969 857 15969 857 6 n_212
rlabel m2contact 15273 137 15273 137 8 IRQ1
rlabel m2contact 15153 353 15153 353 8 n_275
rlabel m2contact 15105 857 15105 857 6 n_212
rlabel m2contact 14913 377 14913 377 8 n_306
rlabel m2contact 14865 569 14865 569 8 n_273
rlabel m2contact 14697 353 14697 353 8 n_260
rlabel m2contact 14577 569 14577 569 8 n_106
rlabel m2contact 14529 641 14529 641 8 n_58
rlabel m2contact 14481 641 14481 641 8 n_219
rlabel m2contact 14433 809 14433 809 6 n_145
rlabel m2contact 14385 377 14385 377 8 n_54
rlabel m2contact 14337 41 14337 41 8 SysBus[2]
rlabel m2contact 14313 233 14313 233 8 SysBus[1]
rlabel m2contact 13953 761 13953 761 2 n_211
rlabel m2contact 13737 713 13737 713 2 n_107
rlabel m2contact 13689 569 13689 569 2 n_106
rlabel m2contact 13617 761 13617 761 2 n_263
rlabel m2contact 13569 809 13569 809 4 n_220
rlabel m2contact 13401 569 13401 569 2 n_106
rlabel m2contact 13329 713 13329 713 2 n_129
rlabel m2contact 13137 569 13137 569 2 n_363
rlabel m2contact 12993 761 12993 761 2 n_263
rlabel m2contact 12849 761 12849 761 2 n_18
rlabel m2contact 12537 353 12537 353 2 n_260
rlabel m2contact 12417 353 12417 353 2 n_267
rlabel m2contact 12369 641 12369 641 2 n_219
rlabel m2contact 12321 233 12321 233 2 n_185
rlabel m2contact 12273 137 12273 137 2 n_94
rlabel m2contact 11265 641 11265 641 2 n_277
rlabel m2contact 11049 929 11049 929 4 n_269
rlabel m2contact 10953 905 10953 905 4 n_229
rlabel m2contact 10833 881 10833 881 4 n_119
rlabel m2contact 10761 329 10761 329 2 n_230
rlabel m2contact 10713 329 10713 329 2 n_179
rlabel m2contact 10641 857 10641 857 4 n_212
rlabel m2contact 10545 137 10545 137 2 n_94
rlabel m2contact 10329 329 10329 329 2 n_179
rlabel m2contact 10113 833 10113 833 4 n_351
rlabel m2contact 9897 833 9897 833 4 n_283
rlabel m2contact 9873 689 9873 689 2 n_216
rlabel m2contact 9705 689 9705 689 2 SysBus[0]
rlabel m2contact 9489 137 9489 137 2 n_201
rlabel m2contact 9417 833 9417 833 4 n_283
rlabel m2contact 9345 809 9345 809 4 n_220
rlabel m2contact 9057 785 9057 785 2 n_33
rlabel m2contact 8769 761 8769 761 2 n_18
rlabel m2contact 8433 737 8433 737 2 n_43
rlabel m2contact 8265 713 8265 713 2 n_129
rlabel m2contact 7941 689 7941 689 2 SysBus[0]
rlabel m2contact 7761 665 7761 665 2 n_265
rlabel m2contact 7569 641 7569 641 2 n_277
rlabel m2contact 7233 617 7233 617 2 n_4
rlabel m2contact 6825 401 6825 401 2 n_354
rlabel m2contact 6633 401 6633 401 2 n_108
rlabel m2contact 6585 593 6585 593 2 n_82
rlabel m2contact 6537 209 6537 209 2 n_87
rlabel m2contact 6417 209 6417 209 2 n_307
rlabel m2contact 6393 569 6393 569 2 n_363
rlabel m2contact 6321 545 6321 545 2 n_113
rlabel m2contact 6249 521 6249 521 2 n_79
rlabel m2contact 5961 497 5961 497 2 n_241
rlabel m2contact 5745 473 5745 473 2 n_218
rlabel m2contact 5649 449 5649 449 2 n_53
rlabel m2contact 5505 425 5505 425 2 n_49
rlabel m2contact 5313 161 5313 161 2 n_401
rlabel m2contact 4953 281 4953 281 2 n_378
rlabel m2contact 4833 161 4833 161 2 n_165
rlabel m2contact 4809 281 4809 281 2 n_73
rlabel m2contact 4785 401 4785 401 2 n_108
rlabel m2contact 4761 377 4761 377 2 n_54
rlabel m2contact 4545 353 4545 353 2 n_267
rlabel m2contact 4377 329 4377 329 2 n_179
rlabel m2contact 4329 305 4329 305 2 n_308
rlabel m2contact 4305 41 4305 41 2 SysBus[2]
rlabel m2contact 3897 281 3897 281 2 n_73
rlabel m2contact 3681 257 3681 257 2 n_304
rlabel m2contact 3633 233 3633 233 2 n_185
rlabel m2contact 3561 209 3561 209 2 n_307
rlabel m2contact 3537 65 3537 65 2 SysBus[3]
rlabel m2contact 2505 185 2505 185 2 n_272
rlabel m2contact 1785 161 1785 161 2 n_165
rlabel m2contact 1665 137 1665 137 2 n_201
rlabel metal2 26127 8444 26139 8444 6 StatusRegEn
rlabel metal2 25287 8444 25299 8444 6 StatusReg[0]
rlabel metal2 24447 8444 24459 8444 6 StatusReg[1]
rlabel metal2 24423 8444 24435 8444 6 StatusReg[2]
rlabel metal2 22767 8444 22779 8444 6 StatusReg[3]
rlabel metal2 22407 8444 22419 8444 6 AluEn
rlabel metal2 21903 8444 21915 8444 6 AluWe
rlabel metal2 20703 8444 20715 8444 6 Op2Sel[0]
rlabel metal2 19407 8444 19419 8444 6 Op2Sel[1]
rlabel metal2 19383 8444 19395 8444 6 Op1Sel
rlabel metal2 17727 8444 17739 8444 6 WdSel
rlabel metal2 17703 8444 17715 8444 6 PcEn
rlabel metal2 16863 8444 16875 8444 6 PcWe
rlabel metal2 15711 8444 15723 8444 6 PcSel[0]
rlabel metal2 15183 8444 15195 8444 6 PcSel[1]
rlabel metal2 13815 8444 13827 8444 4 PcSel[2]
rlabel metal2 12675 8444 12687 8444 4 LrEn
rlabel metal2 12639 8444 12651 8444 4 LrWe
rlabel metal2 11787 8444 11799 8444 4 LrSel
rlabel metal2 10935 8444 10947 8444 4 ImmSel
rlabel metal2 9267 8444 9279 8444 4 IrWe
rlabel metal2 9231 8444 9243 8444 4 MemEn
rlabel metal2 7563 8444 7575 8444 4 OpcodeCondIn[0]
rlabel metal2 7527 8444 7539 8444 4 OpcodeCondIn[1]
rlabel metal2 6279 8444 6291 8444 4 OpcodeCondIn[2]
rlabel metal2 5823 8444 5835 8444 4 OpcodeCondIn[3]
rlabel metal2 4971 8444 4983 8444 4 OpcodeCondIn[4]
rlabel metal2 4119 8444 4131 8444 4 OpcodeCondIn[5]
rlabel metal2 2451 8444 2463 8444 4 OpcodeCondIn[6]
rlabel metal2 2415 8444 2427 8444 4 OpcodeCondIn[7]
rlabel metal2 20691 0 20703 0 8 SysBus[3]
rlabel metal2 14331 0 14343 0 8 SysBus[2]
rlabel metal2 14307 0 14319 0 8 SysBus[1]
rlabel metal2 7935 0 7947 0 2 SysBus[0]
rlabel metal2 0 107 0 119 2 nWE
rlabel metal2 0 83 0 95 2 nIRQ
rlabel metal2 0 4324 0 4336 4 nWait
rlabel metal2 0 4300 0 4312 4 nOE
rlabel metal2 0 8349 0 8361 4 ALE
rlabel metal2 0 8325 0 8337 4 nME
rlabel metal2 27529 515 27529 527 8 Flags[2]
rlabel metal2 27529 59 27529 71 8 Flags[1]
rlabel metal2 27529 35 27529 47 8 Flags[0]
rlabel metal2 27529 11 27529 23 8 CFlag
rlabel metal2 27529 1924 27529 1936 6 RwSel[0]
rlabel metal2 27529 1876 27529 1888 6 Rs1Sel[1]
rlabel metal2 27529 1852 27529 1864 6 Rs1Sel[0]
rlabel metal2 27529 1828 27529 1840 6 Flags[3]
rlabel metal2 27529 8157 27529 8169 6 ENB
rlabel metal2 27529 8133 27529 8145 6 AluOR[1]
rlabel metal2 27529 8109 27529 8121 6 AluOR[0]
rlabel metal2 27529 8085 27529 8097 6 RegWe
rlabel metal2 27529 8061 27529 8073 6 RwSel[1]
rlabel metal2 27171 0 27371 0 1 GND!
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 123 8444 323 8444 5 Vdd!
rlabel metal2 339 8444 351 8444 5 SDO
rlabel metal2 363 8444 375 8444 5 Test
rlabel metal2 387 8444 399 8444 5 Clock
rlabel metal2 411 8444 423 8444 5 nReset
rlabel metal2 27171 8444 27371 8444 5 GND!
<< end >>
