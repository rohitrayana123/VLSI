magic
tech c035u
timestamp 1395748630
<< metal1 >>
rect 7440 41410 7450 41452
rect 7488 41410 7498 41452
rect 7440 41400 7498 41410
rect 6450 40416 6514 40426
rect 6504 40402 6514 40416
rect 7440 40405 7450 41400
rect 7536 40405 7546 41452
rect 11472 41437 11482 41452
rect 11520 41410 11530 41452
rect 15600 41437 15610 41452
rect 11400 41400 11530 41410
rect 11400 41386 11410 41400
rect 15648 41410 15658 41452
rect 19728 41410 19738 41452
rect 19776 41437 19786 41452
rect 19920 41437 19930 41452
rect 27984 41410 27994 41452
rect 28032 41437 28042 41452
rect 28176 41437 28186 41452
rect 32112 41410 32122 41452
rect 32160 41437 32170 41452
rect 32304 41437 32314 41452
rect 36240 41410 36250 41452
rect 11557 41400 15658 41410
rect 15672 41400 36274 41410
rect 11376 41376 11410 41386
rect 11376 41365 11386 41376
rect 15672 41386 15682 41400
rect 36264 41389 36274 41400
rect 36288 41389 36298 41452
rect 36432 41437 36442 41452
rect 36312 41400 36935 41410
rect 36312 41389 36322 41400
rect 11437 41376 15682 41386
rect 19789 41376 36239 41386
rect 36336 41376 36970 41386
rect 11400 41352 11471 41362
rect 11400 41338 11410 41352
rect 11485 41352 15599 41362
rect 36336 41362 36346 41376
rect 28045 41352 36346 41362
rect 36360 41352 36911 41362
rect 11352 41328 11410 41338
rect 11448 41328 11543 41338
rect 6504 40392 6527 40402
rect 11352 40378 11362 41328
rect 11448 41314 11458 41328
rect 11400 41304 11458 41314
rect 6450 40368 11362 40378
rect 6504 35722 6514 40368
rect 6528 35749 6538 40343
rect 7440 37378 7450 40343
rect 7536 37405 7546 40343
rect 11376 37405 11386 41303
rect 11400 37405 11410 41304
rect 11424 37405 11434 41279
rect 15600 37573 15610 41351
rect 19920 37693 19930 41351
rect 36360 41338 36370 41352
rect 36960 41362 36970 41376
rect 36960 41352 36994 41362
rect 28189 41328 36370 41338
rect 36733 41328 36959 41338
rect 36984 41338 36994 41352
rect 36984 41328 37018 41338
rect 37008 41317 37018 41328
rect 36277 41304 36994 41314
rect 32160 37693 32170 41303
rect 32304 37693 32314 41303
rect 36240 41290 36250 41303
rect 36240 41280 36311 41290
rect 36984 41290 36994 41304
rect 36984 41280 37042 41290
rect 36432 41266 36442 41279
rect 36432 41256 36994 41266
rect 36288 37690 36298 41255
rect 36720 37693 36730 41231
rect 36912 37693 36922 41231
rect 36288 37680 36311 37690
rect 36936 37690 36946 41231
rect 36960 37717 36970 41231
rect 36984 37717 36994 41256
rect 37008 37714 37018 41255
rect 37032 40642 37042 41280
rect 37032 40632 41538 40642
rect 41472 40618 41482 40632
rect 41448 40608 41482 40618
rect 41448 40474 41458 40608
rect 41472 40584 41538 40594
rect 41472 40477 41482 40584
rect 41424 40464 41458 40474
rect 37008 37704 37031 37714
rect 36936 37680 37055 37690
rect 18024 37656 37079 37666
rect 18024 37573 18034 37656
rect 36301 37632 36767 37642
rect 36925 37632 37103 37642
rect 19920 37573 19930 37631
rect 28981 37608 37007 37618
rect 37093 37608 37127 37618
rect 28776 37584 37162 37594
rect 28776 37573 28786 37584
rect 37152 37573 37162 37584
rect 29149 37560 37079 37570
rect 15576 37536 36946 37546
rect 7440 37368 11458 37378
rect 6504 35712 6562 35722
rect 6450 35688 6514 35698
rect 6504 35677 6514 35688
rect 6552 35650 6562 35712
rect 6450 35640 6562 35650
rect 6504 30997 6514 35615
rect 6528 30997 6538 35615
rect 6552 30994 6562 35640
rect 6552 30984 6586 30994
rect 6450 30960 6562 30970
rect 6552 30949 6562 30960
rect 6576 30922 6586 30984
rect 6450 30912 6586 30922
rect 6504 26317 6514 30887
rect 6528 26317 6538 30887
rect 6552 26314 6562 30887
rect 6552 26304 6586 26314
rect 6450 26280 6562 26290
rect 6504 21685 6514 26255
rect 6528 21685 6538 26255
rect 6552 21685 6562 26280
rect 6576 21685 6586 26304
rect 6450 21648 6610 21658
rect 6504 16957 6514 21623
rect 6528 16957 6538 21623
rect 6552 16957 6562 21623
rect 6576 16954 6586 21623
rect 6600 16981 6610 21648
rect 6576 16944 6634 16954
rect 6450 16920 6586 16930
rect 6504 12229 6514 16895
rect 6528 15850 6538 16895
rect 6552 15874 6562 16895
rect 6576 15898 6586 16920
rect 6600 16546 6610 16919
rect 6624 16594 6634 16944
rect 7536 16621 7546 37343
rect 11424 37330 11434 37343
rect 11365 37320 11434 37330
rect 11328 37296 11375 37306
rect 11328 16621 11338 37296
rect 11448 37306 11458 37368
rect 11448 37296 11903 37306
rect 11376 37272 12034 37282
rect 11352 16621 11362 37271
rect 11376 16621 11386 37272
rect 12024 37261 12034 37272
rect 15576 37261 15586 37536
rect 36936 37525 36946 37536
rect 36997 37536 37175 37546
rect 16968 37512 36911 37522
rect 15600 37282 15610 37511
rect 16968 37477 16978 37512
rect 36960 37522 36970 37535
rect 36960 37512 37199 37522
rect 26256 37488 36983 37498
rect 26256 37477 26266 37488
rect 37189 37488 37234 37498
rect 37224 37477 37234 37488
rect 26989 37464 37175 37474
rect 16776 37440 36959 37450
rect 16776 37381 16786 37440
rect 37045 37440 37271 37450
rect 25992 37416 37031 37426
rect 16968 37381 16978 37415
rect 18024 37381 18034 37415
rect 19920 37381 19930 37415
rect 25992 37381 26002 37416
rect 37069 37416 37295 37426
rect 29040 37392 37055 37402
rect 29040 37381 29050 37392
rect 37117 37392 37330 37402
rect 37320 37381 37330 37392
rect 32317 37368 36287 37378
rect 36325 37368 37258 37378
rect 37248 37357 37258 37368
rect 15816 37344 37103 37354
rect 15816 37309 15826 37344
rect 37272 37354 37282 37367
rect 37272 37344 37343 37354
rect 19933 37320 37367 37330
rect 32173 37296 36754 37306
rect 15600 37272 36719 37282
rect 36744 37282 36754 37296
rect 36781 37296 37271 37306
rect 37309 37296 37402 37306
rect 36744 37272 37306 37282
rect 36720 37261 36730 37271
rect 11400 16621 11410 37247
rect 36912 34477 36922 37247
rect 36936 34477 36946 37247
rect 36960 34477 36970 37247
rect 36984 34477 36994 37247
rect 37008 34477 37018 37247
rect 37032 34477 37042 37247
rect 37056 34477 37066 37247
rect 37080 34477 37090 37247
rect 37104 34477 37114 37247
rect 37128 34477 37138 37247
rect 37152 34477 37162 37247
rect 37176 34477 37186 37247
rect 37200 34477 37210 37247
rect 37224 34477 37234 37247
rect 37248 34477 37258 37247
rect 37272 34477 37282 37247
rect 37296 34477 37306 37272
rect 37320 34477 37330 37271
rect 37344 34477 37354 37271
rect 37368 34477 37378 37271
rect 37392 34450 37402 37296
rect 41424 35914 41434 40464
rect 41448 40440 41538 40450
rect 41448 35941 41458 40440
rect 41472 35941 41482 40415
rect 41424 35904 41538 35914
rect 41424 35893 41434 35904
rect 41400 35856 41538 35866
rect 41400 35773 41410 35856
rect 41424 35746 41434 35831
rect 41448 35749 41458 35831
rect 41472 35749 41482 35831
rect 36888 34444 37402 34450
rect 36858 34440 37402 34444
rect 41376 35736 41434 35746
rect 36858 34434 36898 34440
rect 37368 34378 37378 34415
rect 36858 34368 37378 34378
rect 36912 33301 36922 34343
rect 36936 33301 36946 34343
rect 36960 33301 36970 34343
rect 36984 33301 36994 34343
rect 37008 33301 37018 34343
rect 37032 33301 37042 34343
rect 37056 33301 37066 34343
rect 37080 33301 37090 34343
rect 37104 33301 37114 34343
rect 37128 33301 37138 34343
rect 37152 33301 37162 34343
rect 37176 33301 37186 34343
rect 37200 33301 37210 34343
rect 37224 33301 37234 34343
rect 37248 33301 37258 34343
rect 37272 33301 37282 34343
rect 37296 33301 37306 34343
rect 37320 33301 37330 34343
rect 37344 33274 37354 34343
rect 36888 33268 37354 33274
rect 36858 33264 37354 33268
rect 36858 33258 36898 33264
rect 37320 33202 37330 33239
rect 36858 33192 37330 33202
rect 36912 32125 36922 33167
rect 36936 32125 36946 33167
rect 36960 32125 36970 33167
rect 36984 32125 36994 33167
rect 37008 32125 37018 33167
rect 37032 32125 37042 33167
rect 37056 32125 37066 33167
rect 37080 32125 37090 33167
rect 37104 32125 37114 33167
rect 37128 32125 37138 33167
rect 37152 32125 37162 33167
rect 37176 32125 37186 33167
rect 37200 32125 37210 33167
rect 37224 32125 37234 33167
rect 37248 32125 37258 33167
rect 37272 32125 37282 33167
rect 37296 32098 37306 33167
rect 36888 32092 37306 32098
rect 36858 32088 37306 32092
rect 36858 32082 36898 32088
rect 37272 32026 37282 32063
rect 36858 32016 37282 32026
rect 36912 30949 36922 31991
rect 36936 30949 36946 31991
rect 36960 30949 36970 31991
rect 36984 30949 36994 31991
rect 37008 30949 37018 31991
rect 37032 30949 37042 31991
rect 37056 30949 37066 31991
rect 37080 30949 37090 31991
rect 37104 30949 37114 31991
rect 37128 30949 37138 31991
rect 37152 30949 37162 31991
rect 37176 30949 37186 31991
rect 37200 30949 37210 31991
rect 37224 30949 37234 31991
rect 37248 30922 37258 31991
rect 41376 31186 41386 35736
rect 41424 35712 41538 35722
rect 41400 31213 41410 35711
rect 41424 31213 41434 35712
rect 41448 31213 41458 35687
rect 41472 31213 41482 35687
rect 41376 31176 41538 31186
rect 41376 31152 41447 31162
rect 41376 31045 41386 31152
rect 41448 31128 41538 31138
rect 41400 31045 41410 31127
rect 41424 31045 41434 31127
rect 41448 31045 41458 31128
rect 41472 31018 41482 31103
rect 36888 30916 37258 30922
rect 36858 30912 37258 30916
rect 41352 31008 41482 31018
rect 36858 30906 36898 30912
rect 37224 30850 37234 30887
rect 36858 30840 37234 30850
rect 36912 29773 36922 30815
rect 36936 29773 36946 30815
rect 36960 29773 36970 30815
rect 36984 29773 36994 30815
rect 37008 29773 37018 30815
rect 37032 29773 37042 30815
rect 37056 29773 37066 30815
rect 37080 29773 37090 30815
rect 37104 29773 37114 30815
rect 37128 29773 37138 30815
rect 37152 29773 37162 30815
rect 37176 29773 37186 30815
rect 37200 29773 37210 30815
rect 41352 29746 41362 31008
rect 41472 30984 41538 30994
rect 36888 29740 41362 29746
rect 36858 29736 41362 29740
rect 36858 29730 36898 29736
rect 41376 29674 41386 30983
rect 36858 29664 41386 29674
rect 36912 28597 36922 29639
rect 36936 28597 36946 29639
rect 36960 28597 36970 29639
rect 36984 28597 36994 29639
rect 37008 28597 37018 29639
rect 37032 28597 37042 29639
rect 37056 28597 37066 29639
rect 37080 28597 37090 29639
rect 37104 28597 37114 29639
rect 37128 28597 37138 29639
rect 37152 28597 37162 29639
rect 37176 28597 37186 29639
rect 37200 28597 37210 29639
rect 41400 28570 41410 30983
rect 36888 28564 41410 28570
rect 36858 28560 41410 28564
rect 36858 28554 36898 28560
rect 41424 28498 41434 30983
rect 36858 28488 41434 28498
rect 36912 27421 36922 28463
rect 36936 27421 36946 28463
rect 36960 27421 36970 28463
rect 36984 27421 36994 28463
rect 37008 27421 37018 28463
rect 37032 27421 37042 28463
rect 37056 27421 37066 28463
rect 37080 27421 37090 28463
rect 37104 27421 37114 28463
rect 37128 27421 37138 28463
rect 37152 27421 37162 28463
rect 37176 27421 37186 28463
rect 37200 27421 37210 28463
rect 41448 27394 41458 30983
rect 36888 27388 41458 27394
rect 36858 27384 41458 27388
rect 36858 27378 36898 27384
rect 41472 27322 41482 30984
rect 36858 27312 41482 27322
rect 36912 26245 36922 27287
rect 36936 26242 36946 27287
rect 36960 26269 36970 27287
rect 36984 26269 36994 27287
rect 37008 26269 37018 27287
rect 37032 26269 37042 27287
rect 37056 26269 37066 27287
rect 37080 26269 37090 27287
rect 37104 26269 37114 27287
rect 37128 26269 37138 27287
rect 37152 26269 37162 27287
rect 37176 26269 37186 27287
rect 37200 26314 37210 27287
rect 37200 26304 41495 26314
rect 36936 26232 37210 26242
rect 36888 26212 36946 26218
rect 36858 26208 36946 26212
rect 36858 26202 36898 26208
rect 36936 26173 36946 26208
rect 36960 26173 36970 26207
rect 36984 26173 36994 26207
rect 37008 26173 37018 26207
rect 37032 26173 37042 26207
rect 37056 26173 37066 26207
rect 37080 26173 37090 26207
rect 37104 26173 37114 26207
rect 37128 26170 37138 26207
rect 37200 26197 37210 26232
rect 37128 26160 37234 26170
rect 36858 26136 37138 26146
rect 36912 25069 36922 26111
rect 36936 25069 36946 26111
rect 36960 25069 36970 26111
rect 36984 25066 36994 26111
rect 37008 25093 37018 26111
rect 37032 25093 37042 26111
rect 37056 25093 37066 26111
rect 37080 25093 37090 26111
rect 37104 25093 37114 26111
rect 37128 25093 37138 26136
rect 37152 25093 37162 26135
rect 37176 25093 37186 26135
rect 37200 25093 37210 26135
rect 37224 25093 37234 26160
rect 36984 25056 37258 25066
rect 36888 25036 36994 25042
rect 36858 25032 36994 25036
rect 36858 25026 36898 25032
rect 36984 25021 36994 25032
rect 37248 25021 37258 25056
rect 36936 24994 36946 25007
rect 36936 24984 37282 24994
rect 36858 24960 36946 24970
rect 36912 23893 36922 24935
rect 36936 23893 36946 24960
rect 36960 23890 36970 24959
rect 36984 23917 36994 24959
rect 37008 23917 37018 24959
rect 37032 23917 37042 24959
rect 37056 23917 37066 24959
rect 37080 23917 37090 24959
rect 37104 23917 37114 24959
rect 37128 23917 37138 24959
rect 37152 23917 37162 24959
rect 37176 23917 37186 24959
rect 37200 23917 37210 24959
rect 37224 23917 37234 24959
rect 37248 23917 37258 24959
rect 37272 23917 37282 24984
rect 36960 23880 37306 23890
rect 36888 23860 36970 23866
rect 36858 23856 36970 23860
rect 36858 23850 36898 23856
rect 36960 23821 36970 23856
rect 36984 23821 36994 23855
rect 37008 23818 37018 23855
rect 37296 23845 37306 23880
rect 37008 23808 37330 23818
rect 36858 23784 37018 23794
rect 36912 22717 36922 23759
rect 36936 22717 36946 23759
rect 36960 22717 36970 23759
rect 36984 22717 36994 23759
rect 37008 22717 37018 23784
rect 37032 22717 37042 23783
rect 37056 22714 37066 23783
rect 37080 22741 37090 23783
rect 37104 22741 37114 23783
rect 37128 22741 37138 23783
rect 37152 22741 37162 23783
rect 37176 22741 37186 23783
rect 37200 22741 37210 23783
rect 37224 22741 37234 23783
rect 37248 22741 37258 23783
rect 37272 22741 37282 23783
rect 37296 22741 37306 23783
rect 37320 22741 37330 23808
rect 37056 22704 37354 22714
rect 36888 22684 37066 22690
rect 36858 22680 37066 22684
rect 36858 22674 36898 22680
rect 37056 22645 37066 22680
rect 37080 22642 37090 22679
rect 37344 22669 37354 22704
rect 37080 22632 37378 22642
rect 36858 22608 37090 22618
rect 36912 21541 36922 22583
rect 36936 21541 36946 22583
rect 36960 21541 36970 22583
rect 36984 21541 36994 22583
rect 37008 21541 37018 22583
rect 37032 21541 37042 22583
rect 37056 21541 37066 22583
rect 37080 21541 37090 22608
rect 37104 21538 37114 22607
rect 37128 21565 37138 22607
rect 37152 21565 37162 22607
rect 37176 21565 37186 22607
rect 37200 21565 37210 22607
rect 37224 21565 37234 22607
rect 37248 21565 37258 22607
rect 37272 21565 37282 22607
rect 37296 21565 37306 22607
rect 37320 21565 37330 22607
rect 37344 21565 37354 22607
rect 37368 21565 37378 22632
rect 37104 21528 37402 21538
rect 36888 21508 37114 21514
rect 36858 21504 37114 21508
rect 36858 21498 36898 21504
rect 37104 21493 37114 21504
rect 37392 21493 37402 21528
rect 36912 21466 36922 21479
rect 36912 21456 37426 21466
rect 36858 21432 36922 21442
rect 36912 20365 36922 21432
rect 36936 20365 36946 21431
rect 36960 20365 36970 21431
rect 36984 20365 36994 21431
rect 37008 20365 37018 21431
rect 37032 20365 37042 21431
rect 37056 20365 37066 21431
rect 37080 20365 37090 21431
rect 37104 20365 37114 21431
rect 37128 20365 37138 21431
rect 37152 20365 37162 21431
rect 37176 20365 37186 21431
rect 37200 20365 37210 21431
rect 37224 20365 37234 21431
rect 37248 20365 37258 21431
rect 37272 20362 37282 21431
rect 37296 20389 37306 21431
rect 37320 20389 37330 21431
rect 37344 20389 37354 21431
rect 37368 20389 37378 21431
rect 37392 20389 37402 21431
rect 37416 20389 37426 21456
rect 37272 20352 37450 20362
rect 36888 20332 37282 20338
rect 36858 20328 37282 20332
rect 36858 20322 36898 20328
rect 37272 20317 37282 20328
rect 37440 20317 37450 20352
rect 37176 20290 37186 20303
rect 37176 20280 37474 20290
rect 36858 20256 37186 20266
rect 36912 19189 36922 20231
rect 36936 19189 36946 20231
rect 36960 19189 36970 20231
rect 36984 19189 36994 20231
rect 37008 19189 37018 20231
rect 37032 19189 37042 20231
rect 37056 19186 37066 20231
rect 37080 19213 37090 20231
rect 37104 19213 37114 20231
rect 37128 19213 37138 20231
rect 37152 19213 37162 20231
rect 37176 19213 37186 20256
rect 37200 19213 37210 20255
rect 37224 19213 37234 20255
rect 37248 19213 37258 20255
rect 37272 19213 37282 20255
rect 37296 19213 37306 20255
rect 37320 19213 37330 20255
rect 37344 19213 37354 20255
rect 37368 19213 37378 20255
rect 37392 19213 37402 20255
rect 37416 19213 37426 20255
rect 37440 19213 37450 20255
rect 37464 19213 37474 20280
rect 37056 19176 37498 19186
rect 36888 19156 37066 19162
rect 36858 19152 37066 19156
rect 36858 19146 36898 19152
rect 37056 19141 37066 19152
rect 37488 19141 37498 19176
rect 37032 19114 37042 19127
rect 37032 19104 37522 19114
rect 36858 19080 37042 19090
rect 36912 18010 36922 19055
rect 36936 18037 36946 19055
rect 36960 18037 36970 19055
rect 36984 18037 36994 19055
rect 37008 18037 37018 19055
rect 37032 18037 37042 19080
rect 37056 18037 37066 19079
rect 37080 18037 37090 19079
rect 37104 18037 37114 19079
rect 37128 18037 37138 19079
rect 37152 18037 37162 19079
rect 37176 18037 37186 19079
rect 37200 18037 37210 19079
rect 37224 18037 37234 19079
rect 37248 18037 37258 19079
rect 37272 18037 37282 19079
rect 37296 18037 37306 19079
rect 37320 18037 37330 19079
rect 37344 18037 37354 19079
rect 37368 18037 37378 19079
rect 37392 18037 37402 19079
rect 37416 18037 37426 19079
rect 37440 18037 37450 19079
rect 37464 18037 37474 19079
rect 37488 18037 37498 19079
rect 37512 18037 37522 19104
rect 36912 18000 37546 18010
rect 36888 17980 36922 17986
rect 36858 17976 36922 17980
rect 36858 17970 36898 17976
rect 36912 17941 36922 17976
rect 36936 17941 36946 17975
rect 36960 17941 36970 17975
rect 36984 17941 36994 17975
rect 37008 17941 37018 17975
rect 37032 17941 37042 17975
rect 37056 17941 37066 17975
rect 37080 17941 37090 17975
rect 37104 17941 37114 17975
rect 37128 17941 37138 17975
rect 37152 17941 37162 17975
rect 37176 17941 37186 17975
rect 37200 17941 37210 17975
rect 37224 17941 37234 17975
rect 37248 17941 37258 17975
rect 37272 17941 37282 17975
rect 37296 17941 37306 17975
rect 37320 17941 37330 17975
rect 37344 17941 37354 17975
rect 37368 17941 37378 17975
rect 37392 17941 37402 17975
rect 37416 17941 37426 17975
rect 37440 17938 37450 17975
rect 37536 17965 37546 18000
rect 37440 17928 37570 17938
rect 36858 17904 37450 17914
rect 36912 16837 36922 17879
rect 36936 16837 36946 17879
rect 36960 16837 36970 17879
rect 36984 16837 36994 17879
rect 37008 16837 37018 17879
rect 37032 16837 37042 17879
rect 37056 16837 37066 17879
rect 37080 16837 37090 17879
rect 37104 16837 37114 17879
rect 37128 16834 37138 17879
rect 37152 16861 37162 17879
rect 37176 16861 37186 17879
rect 37200 16861 37210 17879
rect 37224 16861 37234 17879
rect 37248 16861 37258 17879
rect 37272 16861 37282 17879
rect 37296 16861 37306 17879
rect 37320 16861 37330 17879
rect 37344 16861 37354 17879
rect 37368 16861 37378 17879
rect 37392 16861 37402 17879
rect 37416 16861 37426 17879
rect 37440 16861 37450 17904
rect 37464 16861 37474 17903
rect 37488 16861 37498 17903
rect 37512 16861 37522 17903
rect 37536 16861 37546 17903
rect 37560 16930 37570 17928
rect 41472 16968 41538 16978
rect 41472 16957 41482 16968
rect 37560 16920 41538 16930
rect 37128 16824 37570 16834
rect 36888 16804 37138 16810
rect 36858 16800 37138 16804
rect 36858 16794 36898 16800
rect 37128 16789 37138 16800
rect 37560 16786 37570 16824
rect 41472 16813 41482 16895
rect 37560 16776 41538 16786
rect 37032 16762 37042 16775
rect 37032 16752 37570 16762
rect 36858 16728 37042 16738
rect 36912 16621 36922 16703
rect 36936 16621 36946 16703
rect 36960 16621 36970 16703
rect 36984 16621 36994 16703
rect 37008 16618 37018 16703
rect 37032 16645 37042 16728
rect 37056 16645 37066 16727
rect 37080 16645 37090 16727
rect 37104 16645 37114 16727
rect 37128 16645 37138 16727
rect 37152 16645 37162 16727
rect 37176 16645 37186 16727
rect 37200 16645 37210 16727
rect 37224 16645 37234 16727
rect 37248 16645 37258 16727
rect 37272 16645 37282 16727
rect 37296 16645 37306 16727
rect 37320 16645 37330 16727
rect 37344 16645 37354 16727
rect 37368 16645 37378 16727
rect 37392 16645 37402 16727
rect 37416 16645 37426 16727
rect 37440 16645 37450 16727
rect 37464 16645 37474 16727
rect 37488 16645 37498 16727
rect 37512 16645 37522 16727
rect 37536 16645 37546 16727
rect 37560 16645 37570 16752
rect 37008 16608 37594 16618
rect 11904 16594 11914 16607
rect 6624 16584 11434 16594
rect 11424 16573 11434 16584
rect 11640 16584 11914 16594
rect 11640 16573 11650 16584
rect 12109 16594 12119 16607
rect 11941 16584 12119 16594
rect 11664 16560 12035 16570
rect 11664 16546 11674 16560
rect 12060 16546 12070 16559
rect 6600 16536 11674 16546
rect 11750 16536 12070 16546
rect 7536 15925 7546 16511
rect 11328 16018 11338 16511
rect 11293 16008 11338 16018
rect 11352 15994 11362 16511
rect 11269 15984 11362 15994
rect 11376 15970 11386 16511
rect 11400 15973 11410 16511
rect 11424 15973 11434 16511
rect 11245 15960 11386 15970
rect 11451 15970 11461 16511
rect 11472 15994 11482 16484
rect 11497 16018 11507 16511
rect 11520 16042 11530 16484
rect 11544 16066 11554 16511
rect 11568 16090 11578 16484
rect 11591 16114 11601 16511
rect 11612 16138 11622 16484
rect 11640 16165 11650 16511
rect 11750 16141 11760 16536
rect 12084 16522 12094 16559
rect 11774 16512 12094 16522
rect 11774 16141 11784 16512
rect 11798 16488 11927 16498
rect 11798 16141 11808 16488
rect 11612 16128 11663 16138
rect 11591 16104 11831 16114
rect 11568 16080 11855 16090
rect 11544 16056 11879 16066
rect 13368 16066 13378 16607
rect 13560 16090 13570 16607
rect 13560 16080 13847 16090
rect 14352 16090 14362 16607
rect 14352 16080 14711 16090
rect 14904 16090 14914 16607
rect 15120 16114 15130 16607
rect 15120 16104 15575 16114
rect 15864 16114 15874 16607
rect 16032 16138 16042 16607
rect 16416 16165 16426 16607
rect 16608 16162 16618 16607
rect 16824 16186 16834 16607
rect 16824 16176 16991 16186
rect 17568 16186 17578 16607
rect 17736 16210 17746 16607
rect 17736 16200 18167 16210
rect 17568 16176 18191 16186
rect 16608 16152 19895 16162
rect 16032 16128 20759 16138
rect 15864 16104 21191 16114
rect 14904 16080 22127 16090
rect 13368 16056 20735 16066
rect 20773 16056 22895 16066
rect 11520 16032 16967 16042
rect 17005 16032 23927 16042
rect 11497 16008 18143 16018
rect 18181 16008 24239 16018
rect 11472 15984 18167 15994
rect 18205 15984 25823 15994
rect 27144 15973 27154 16607
rect 11451 15960 19871 15970
rect 19909 15960 26783 15970
rect 27336 15970 27346 16607
rect 27576 15994 27586 16607
rect 35280 16594 35290 16607
rect 32760 16584 35290 16594
rect 27576 15984 27671 15994
rect 32760 15973 32770 16584
rect 35319 16584 36239 16594
rect 36301 16584 37018 16594
rect 37008 16573 37018 16584
rect 37584 16573 37594 16608
rect 33600 16560 36023 16570
rect 33600 15973 33610 16560
rect 36048 16560 36311 16570
rect 36048 16546 36058 16560
rect 35282 16536 36058 16546
rect 35282 15973 35292 16536
rect 36181 16536 36287 16546
rect 36384 16546 36394 16559
rect 36384 16536 37618 16546
rect 36168 16512 36215 16522
rect 35306 15973 35316 16511
rect 36168 15973 36178 16512
rect 36253 16512 36263 16522
rect 37608 16522 37618 16536
rect 37608 16512 38591 16522
rect 36720 16498 36730 16511
rect 36720 16488 38855 16498
rect 37597 16464 39167 16474
rect 36912 15973 36922 16463
rect 36936 15973 36946 16463
rect 36960 15973 36970 16463
rect 36984 15973 36994 16463
rect 37008 15973 37018 16463
rect 27336 15960 28511 15970
rect 11197 15936 11279 15946
rect 37032 15946 37042 16463
rect 11317 15936 37042 15946
rect 37056 15946 37066 16463
rect 37080 15970 37090 16463
rect 37104 15994 37114 16463
rect 37128 16018 37138 16463
rect 37152 16042 37162 16463
rect 37176 16066 37186 16463
rect 37200 16090 37210 16463
rect 37224 16114 37234 16463
rect 37248 16138 37258 16463
rect 37272 16162 37282 16463
rect 37296 16186 37306 16463
rect 37320 16210 37330 16463
rect 37344 16234 37354 16463
rect 37368 16258 37378 16463
rect 37392 16282 37402 16463
rect 37416 16306 37426 16463
rect 37440 16330 37450 16463
rect 37464 16354 37474 16463
rect 37488 16378 37498 16463
rect 37512 16402 37522 16463
rect 37536 16426 37546 16463
rect 37560 16450 37570 16463
rect 37560 16440 39191 16450
rect 37536 16416 39215 16426
rect 37512 16392 39239 16402
rect 37488 16368 39263 16378
rect 37464 16344 39287 16354
rect 37440 16320 39311 16330
rect 37416 16296 39335 16306
rect 37392 16272 39359 16282
rect 37368 16248 39383 16258
rect 37344 16224 39407 16234
rect 37320 16200 39431 16210
rect 37296 16176 39455 16186
rect 37272 16152 39479 16162
rect 37248 16128 39503 16138
rect 37224 16104 39527 16114
rect 37200 16080 39551 16090
rect 37176 16056 39575 16066
rect 37152 16032 39647 16042
rect 37128 16008 39671 16018
rect 37104 15984 39695 15994
rect 37080 15960 39743 15970
rect 37056 15936 39791 15946
rect 11149 15912 11399 15922
rect 11437 15912 11725 15922
rect 11893 15912 16391 15922
rect 16429 15912 26759 15922
rect 27157 15912 30193 15922
rect 36997 15912 41375 15922
rect 6576 15888 11749 15898
rect 11856 15898 11866 15911
rect 11856 15888 15551 15898
rect 15589 15888 23903 15898
rect 23941 15888 27647 15898
rect 27685 15888 30218 15898
rect 6552 15864 7463 15874
rect 7477 15864 11591 15874
rect 11605 15864 11639 15874
rect 11677 15864 13823 15874
rect 13861 15864 21167 15874
rect 21205 15864 24215 15874
rect 24253 15864 28487 15874
rect 28525 15864 31607 15874
rect 6528 15840 11290 15850
rect 7464 12229 7474 15815
rect 7536 12229 7546 15815
rect 11136 15684 11146 15815
rect 11184 15709 11194 15815
rect 11232 15709 11242 15815
rect 11256 15709 11266 15815
rect 11280 15709 11290 15840
rect 11328 15840 11773 15850
rect 11304 15709 11314 15839
rect 11328 15709 11338 15840
rect 11845 15840 14698 15850
rect 14688 15829 14698 15840
rect 14725 15840 22114 15850
rect 22104 15829 22114 15840
rect 22141 15840 22882 15850
rect 22872 15829 22882 15840
rect 22909 15840 25810 15850
rect 25800 15829 25810 15840
rect 25837 15840 30181 15850
rect 30171 15829 30181 15840
rect 30232 15840 31906 15850
rect 31896 15829 31906 15840
rect 32760 15829 32770 15911
rect 33600 15829 33610 15911
rect 36168 15829 36178 15911
rect 36912 15850 36922 15911
rect 36936 15874 36946 15911
rect 36960 15898 36970 15911
rect 36960 15888 41423 15898
rect 36936 15864 41447 15874
rect 41472 15850 41482 16751
rect 36912 15840 39610 15850
rect 11136 15674 11351 15684
rect 11197 15650 11351 15660
rect 11232 12229 11242 15623
rect 11256 12229 11266 15623
rect 11280 12229 11290 15623
rect 11304 12229 11314 15623
rect 11328 12202 11338 15623
rect 39168 15615 39178 15815
rect 39192 15615 39202 15815
rect 39216 15615 39226 15815
rect 39240 15615 39250 15815
rect 39264 15615 39274 15815
rect 39288 15588 39298 15815
rect 39312 15591 39322 15815
rect 39336 15591 39346 15815
rect 39360 15591 39370 15815
rect 39384 15591 39394 15815
rect 39157 15578 39298 15588
rect 39408 15564 39418 15815
rect 39432 15567 39442 15815
rect 39456 15567 39466 15815
rect 39480 15567 39490 15815
rect 39504 15567 39514 15815
rect 39528 15567 39538 15815
rect 39552 15567 39562 15815
rect 39576 15567 39586 15815
rect 39600 15567 39610 15840
rect 39624 15840 41482 15850
rect 39624 15567 39634 15840
rect 39157 15554 39418 15564
rect 39648 15540 39658 15815
rect 39157 15530 39658 15540
rect 39157 15506 39431 15516
rect 39157 15482 39383 15492
rect 6450 12192 11338 12202
rect 6504 7666 6514 12167
rect 7464 7693 7474 12167
rect 7536 11587 7546 12167
rect 11232 11612 11242 12167
rect 11256 11612 11266 12167
rect 11280 11612 11290 12167
rect 11304 11612 11314 12167
rect 7536 11577 11351 11587
rect 11293 11553 11351 11563
rect 11232 7693 11242 11543
rect 11256 7693 11266 11543
rect 11304 7693 11314 11519
rect 39168 10501 39178 15457
rect 39192 10501 39202 15457
rect 39216 10501 39226 15457
rect 39240 10501 39250 15457
rect 39264 10501 39274 15457
rect 39312 10501 39322 15457
rect 39336 10501 39346 15457
rect 39360 10501 39370 15457
rect 39456 10501 39466 15505
rect 39480 10501 39490 15505
rect 39504 10501 39514 15505
rect 39528 10501 39538 15505
rect 39552 10474 39562 15505
rect 39157 10464 39562 10474
rect 39168 9261 39178 10439
rect 39192 9261 39202 10439
rect 39216 9261 39226 10439
rect 39240 9261 39250 10439
rect 39264 9261 39274 10439
rect 39312 9261 39322 10439
rect 39336 9261 39346 10439
rect 39360 9235 39370 10439
rect 39157 9225 39370 9235
rect 39456 9211 39466 10439
rect 39157 9201 39466 9211
rect 39157 9177 39335 9187
rect 39168 8053 39178 9143
rect 39192 8053 39202 9143
rect 39216 8053 39226 9143
rect 39240 8053 39250 9143
rect 39264 8053 39274 9143
rect 39312 8053 39322 9143
rect 39480 8053 39490 10439
rect 39504 8053 39514 10439
rect 39528 8026 39538 10439
rect 39157 8016 39538 8026
rect 39168 7693 39178 7991
rect 39192 7693 39202 7991
rect 39216 7693 39226 7991
rect 39240 7693 39250 7991
rect 39264 7693 39274 7991
rect 39312 7693 39322 7991
rect 39480 7693 39490 7991
rect 6504 7656 11351 7666
rect 39504 7658 39514 7991
rect 39157 7648 39514 7658
rect 39576 7645 39586 15505
rect 39600 7645 39610 15505
rect 7464 7501 7474 7631
rect 11232 7525 11242 7631
rect 11256 7525 11266 7631
rect 11304 7573 11314 7631
rect 39157 7624 39239 7634
rect 39624 7610 39634 15505
rect 39157 7600 39634 7610
rect 11808 7546 11818 7559
rect 11280 7536 11818 7546
rect 11832 7536 19367 7546
rect 11280 7498 11290 7536
rect 11208 7488 11290 7498
rect 11352 7512 11735 7522
rect 11208 7474 11218 7488
rect 6450 7464 11218 7474
rect 11352 7474 11362 7512
rect 11832 7522 11842 7536
rect 19392 7536 22559 7546
rect 19392 7522 19402 7536
rect 39192 7546 39202 7568
rect 22584 7536 39202 7546
rect 22584 7522 22594 7536
rect 11760 7512 11842 7522
rect 15816 7512 19402 7522
rect 19800 7512 22594 7522
rect 22608 7512 25823 7522
rect 11760 7498 11770 7512
rect 11245 7464 11362 7474
rect 11688 7488 11770 7498
rect 7464 6565 7474 7439
rect 11256 6562 11266 7439
rect 11304 6589 11314 7439
rect 11328 6589 11338 7439
rect 11256 6552 11362 6562
rect 7440 6528 11327 6538
rect 7440 6514 7450 6528
rect 11352 6538 11362 6552
rect 11688 6541 11698 7488
rect 15816 7453 15826 7512
rect 19368 7450 19378 7487
rect 19800 7477 19810 7512
rect 22608 7498 22618 7512
rect 28200 7512 35303 7522
rect 19944 7488 22618 7498
rect 19944 7477 19954 7488
rect 25824 7477 25834 7511
rect 28200 7477 28210 7512
rect 35317 7512 36455 7522
rect 39216 7522 39226 7568
rect 36480 7512 39226 7522
rect 39240 7522 39250 7600
rect 39672 7549 39682 15815
rect 39696 7549 39706 15815
rect 39744 7549 39754 15815
rect 39792 7549 39802 15815
rect 41376 12202 41386 15815
rect 41424 12229 41434 15815
rect 41448 12229 41458 15815
rect 41472 12250 41482 15840
rect 41472 12240 41538 12250
rect 41376 12192 41538 12202
rect 41424 7549 41434 12167
rect 41448 12058 41458 12167
rect 41448 12048 41538 12058
rect 39240 7512 41538 7522
rect 36480 7498 36490 7512
rect 41472 7501 41482 7512
rect 32184 7488 36490 7498
rect 32184 7477 32194 7488
rect 36517 7488 39479 7498
rect 36493 7464 39263 7474
rect 39672 7450 39682 7487
rect 19368 7440 39682 7450
rect 15672 7416 39311 7426
rect 15672 6541 15682 7416
rect 36469 7392 36503 7402
rect 39181 7392 39191 7402
rect 15816 6541 15826 7391
rect 19800 6541 19810 7391
rect 19944 6541 19954 7391
rect 22560 7378 22570 7391
rect 39600 7378 39610 7415
rect 39696 7381 39706 7487
rect 39744 7381 39754 7487
rect 22560 7368 39610 7378
rect 36469 7344 36479 7354
rect 39792 7354 39802 7487
rect 41424 7474 41434 7487
rect 41424 7464 41538 7474
rect 41472 7357 41482 7439
rect 39168 7344 39802 7354
rect 25824 7330 25834 7343
rect 39168 7330 39178 7344
rect 25824 7320 39178 7330
rect 39205 7320 41538 7330
rect 28200 6565 28210 7295
rect 32184 6565 32194 7295
rect 36456 6613 36466 7295
rect 39576 6637 39586 7295
rect 39696 6637 39706 7295
rect 39744 6637 39754 7295
rect 41472 6610 41482 7295
rect 36517 6600 41482 6610
rect 36325 6576 36551 6586
rect 39696 6562 39706 6575
rect 32341 6552 39706 6562
rect 11352 6528 11578 6538
rect 7416 6504 7450 6514
rect 7416 6450 7426 6504
rect 7477 6504 7522 6514
rect 7464 6450 7474 6503
rect 7512 6450 7522 6504
rect 11568 6514 11578 6528
rect 28069 6528 36538 6538
rect 11317 6504 11554 6514
rect 11568 6504 36503 6514
rect 11544 6450 11554 6504
rect 11688 6450 11698 6479
rect 11736 6450 11746 6504
rect 15672 6450 15682 6479
rect 15816 6450 15826 6479
rect 15864 6450 15874 6504
rect 19800 6450 19810 6479
rect 19944 6450 19954 6479
rect 19992 6450 20002 6504
rect 28056 6450 28066 6479
rect 28200 6450 28210 6479
rect 28248 6450 28258 6504
rect 32184 6450 32194 6479
rect 32328 6450 32338 6479
rect 32376 6450 32386 6504
rect 36528 6514 36538 6528
rect 39744 6538 39754 6575
rect 36565 6528 39754 6538
rect 36528 6504 39575 6514
rect 36312 6450 36322 6479
rect 36456 6450 36466 6479
rect 36504 6450 36514 6503
<< m2contact >>
rect 11471 41423 11485 41437
rect 15599 41423 15613 41437
rect 11543 41399 11557 41413
rect 19775 41423 19789 41437
rect 19919 41423 19933 41437
rect 28031 41423 28045 41437
rect 28175 41423 28189 41437
rect 32159 41423 32173 41437
rect 32303 41423 32317 41437
rect 11423 41375 11437 41389
rect 36431 41423 36445 41437
rect 36935 41399 36949 41413
rect 19775 41375 19789 41389
rect 36239 41375 36253 41389
rect 36263 41375 36277 41389
rect 36287 41375 36301 41389
rect 36311 41375 36325 41389
rect 11375 41351 11389 41365
rect 11471 41351 11485 41365
rect 15599 41351 15613 41365
rect 19919 41351 19933 41365
rect 28031 41351 28045 41365
rect 6527 40391 6541 40405
rect 7439 40391 7453 40405
rect 7535 40391 7549 40405
rect 11375 41303 11389 41317
rect 11543 41327 11557 41341
rect 6527 40343 6541 40357
rect 7439 40343 7453 40357
rect 7535 40343 7549 40357
rect 11423 41279 11437 41293
rect 28175 41327 28189 41341
rect 36911 41351 36925 41365
rect 36719 41327 36733 41341
rect 36959 41327 36973 41341
rect 32159 41303 32173 41317
rect 32303 41303 32317 41317
rect 36239 41303 36253 41317
rect 36263 41303 36277 41317
rect 36311 41279 36325 41293
rect 36431 41279 36445 41293
rect 37007 41303 37021 41317
rect 36287 41255 36301 41269
rect 19919 37679 19933 37693
rect 32159 37679 32173 37693
rect 32303 37679 32317 37693
rect 36719 41231 36733 41245
rect 36911 41231 36925 41245
rect 36935 41231 36949 41245
rect 36959 41231 36973 41245
rect 36311 37679 36325 37693
rect 36719 37679 36733 37693
rect 36911 37679 36925 37693
rect 37007 41255 37021 41269
rect 36959 37703 36973 37717
rect 36983 37703 36997 37717
rect 37031 37703 37045 37717
rect 37055 37679 37069 37693
rect 37079 37655 37093 37669
rect 19919 37631 19933 37645
rect 36287 37631 36301 37645
rect 36767 37631 36781 37645
rect 36911 37631 36925 37645
rect 37103 37631 37117 37645
rect 28967 37607 28981 37621
rect 37007 37607 37021 37621
rect 37079 37607 37093 37621
rect 37127 37607 37141 37621
rect 15599 37559 15613 37573
rect 18023 37559 18037 37573
rect 19919 37559 19933 37573
rect 28775 37559 28789 37573
rect 29135 37559 29149 37573
rect 37079 37559 37093 37573
rect 37151 37559 37165 37573
rect 7535 37391 7549 37405
rect 11375 37391 11389 37405
rect 11399 37391 11413 37405
rect 11423 37391 11437 37405
rect 7535 37343 7549 37357
rect 11423 37343 11437 37357
rect 6527 35735 6541 35749
rect 6503 35663 6517 35677
rect 6503 35615 6517 35629
rect 6527 35615 6541 35629
rect 6503 30983 6517 30997
rect 6527 30983 6541 30997
rect 6551 30935 6565 30949
rect 6503 30887 6517 30901
rect 6527 30887 6541 30901
rect 6551 30887 6565 30901
rect 6503 26303 6517 26317
rect 6527 26303 6541 26317
rect 6503 26255 6517 26269
rect 6527 26255 6541 26269
rect 6503 21671 6517 21685
rect 6527 21671 6541 21685
rect 6551 21671 6565 21685
rect 6575 21671 6589 21685
rect 6503 21623 6517 21637
rect 6527 21623 6541 21637
rect 6551 21623 6565 21637
rect 6575 21623 6589 21637
rect 6503 16943 6517 16957
rect 6527 16943 6541 16957
rect 6551 16943 6565 16957
rect 6599 16967 6613 16981
rect 6503 16895 6517 16909
rect 6527 16895 6541 16909
rect 6551 16895 6565 16909
rect 6599 16919 6613 16933
rect 11351 37319 11365 37333
rect 11375 37295 11389 37309
rect 11903 37295 11917 37309
rect 11351 37271 11365 37285
rect 36959 37535 36973 37549
rect 36983 37535 36997 37549
rect 37175 37535 37189 37549
rect 15599 37511 15613 37525
rect 36911 37511 36925 37525
rect 36935 37511 36949 37525
rect 37199 37511 37213 37525
rect 36983 37487 36997 37501
rect 37175 37487 37189 37501
rect 16967 37463 16981 37477
rect 26255 37463 26269 37477
rect 26975 37463 26989 37477
rect 37175 37463 37189 37477
rect 37223 37463 37237 37477
rect 36959 37439 36973 37453
rect 37031 37439 37045 37453
rect 37271 37439 37285 37453
rect 16967 37415 16981 37429
rect 18023 37415 18037 37429
rect 19919 37415 19933 37429
rect 37031 37415 37045 37429
rect 37055 37415 37069 37429
rect 37295 37415 37309 37429
rect 37055 37391 37069 37405
rect 37103 37391 37117 37405
rect 16775 37367 16789 37381
rect 16967 37367 16981 37381
rect 18023 37367 18037 37381
rect 19919 37367 19933 37381
rect 25991 37367 26005 37381
rect 29039 37367 29053 37381
rect 32303 37367 32317 37381
rect 36287 37367 36301 37381
rect 36311 37367 36325 37381
rect 37271 37367 37285 37381
rect 37319 37367 37333 37381
rect 37103 37343 37117 37357
rect 37247 37343 37261 37357
rect 37343 37343 37357 37357
rect 19919 37319 19933 37333
rect 37367 37319 37381 37333
rect 15815 37295 15829 37309
rect 32159 37295 32173 37309
rect 36719 37271 36733 37285
rect 36767 37295 36781 37309
rect 37271 37295 37285 37309
rect 37295 37295 37309 37309
rect 11399 37247 11413 37261
rect 12023 37247 12037 37261
rect 15575 37247 15589 37261
rect 36719 37247 36733 37261
rect 36911 37247 36925 37261
rect 36935 37247 36949 37261
rect 36959 37247 36973 37261
rect 36983 37247 36997 37261
rect 37007 37247 37021 37261
rect 37031 37247 37045 37261
rect 37055 37247 37069 37261
rect 37079 37247 37093 37261
rect 37103 37247 37117 37261
rect 37127 37247 37141 37261
rect 37151 37247 37165 37261
rect 37175 37247 37189 37261
rect 37199 37247 37213 37261
rect 37223 37247 37237 37261
rect 37247 37247 37261 37261
rect 37271 37247 37285 37261
rect 37319 37271 37333 37285
rect 37343 37271 37357 37285
rect 37367 37271 37381 37285
rect 36911 34463 36925 34477
rect 36935 34463 36949 34477
rect 36959 34463 36973 34477
rect 36983 34463 36997 34477
rect 37007 34463 37021 34477
rect 37031 34463 37045 34477
rect 37055 34463 37069 34477
rect 37079 34463 37093 34477
rect 37103 34463 37117 34477
rect 37127 34463 37141 34477
rect 37151 34463 37165 34477
rect 37175 34463 37189 34477
rect 37199 34463 37213 34477
rect 37223 34463 37237 34477
rect 37247 34463 37261 34477
rect 37271 34463 37285 34477
rect 37295 34463 37309 34477
rect 37319 34463 37333 34477
rect 37343 34463 37357 34477
rect 37367 34463 37381 34477
rect 41471 40463 41485 40477
rect 41471 40415 41485 40429
rect 41447 35927 41461 35941
rect 41471 35927 41485 35941
rect 41423 35879 41437 35893
rect 41423 35831 41437 35845
rect 41447 35831 41461 35845
rect 41471 35831 41485 35845
rect 41399 35759 41413 35773
rect 37367 34415 37381 34429
rect 36911 34343 36925 34357
rect 36935 34343 36949 34357
rect 36959 34343 36973 34357
rect 36983 34343 36997 34357
rect 37007 34343 37021 34357
rect 37031 34343 37045 34357
rect 37055 34343 37069 34357
rect 37079 34343 37093 34357
rect 37103 34343 37117 34357
rect 37127 34343 37141 34357
rect 37151 34343 37165 34357
rect 37175 34343 37189 34357
rect 37199 34343 37213 34357
rect 37223 34343 37237 34357
rect 37247 34343 37261 34357
rect 37271 34343 37285 34357
rect 37295 34343 37309 34357
rect 37319 34343 37333 34357
rect 37343 34343 37357 34357
rect 36911 33287 36925 33301
rect 36935 33287 36949 33301
rect 36959 33287 36973 33301
rect 36983 33287 36997 33301
rect 37007 33287 37021 33301
rect 37031 33287 37045 33301
rect 37055 33287 37069 33301
rect 37079 33287 37093 33301
rect 37103 33287 37117 33301
rect 37127 33287 37141 33301
rect 37151 33287 37165 33301
rect 37175 33287 37189 33301
rect 37199 33287 37213 33301
rect 37223 33287 37237 33301
rect 37247 33287 37261 33301
rect 37271 33287 37285 33301
rect 37295 33287 37309 33301
rect 37319 33287 37333 33301
rect 37319 33239 37333 33253
rect 36911 33167 36925 33181
rect 36935 33167 36949 33181
rect 36959 33167 36973 33181
rect 36983 33167 36997 33181
rect 37007 33167 37021 33181
rect 37031 33167 37045 33181
rect 37055 33167 37069 33181
rect 37079 33167 37093 33181
rect 37103 33167 37117 33181
rect 37127 33167 37141 33181
rect 37151 33167 37165 33181
rect 37175 33167 37189 33181
rect 37199 33167 37213 33181
rect 37223 33167 37237 33181
rect 37247 33167 37261 33181
rect 37271 33167 37285 33181
rect 37295 33167 37309 33181
rect 36911 32111 36925 32125
rect 36935 32111 36949 32125
rect 36959 32111 36973 32125
rect 36983 32111 36997 32125
rect 37007 32111 37021 32125
rect 37031 32111 37045 32125
rect 37055 32111 37069 32125
rect 37079 32111 37093 32125
rect 37103 32111 37117 32125
rect 37127 32111 37141 32125
rect 37151 32111 37165 32125
rect 37175 32111 37189 32125
rect 37199 32111 37213 32125
rect 37223 32111 37237 32125
rect 37247 32111 37261 32125
rect 37271 32111 37285 32125
rect 37271 32063 37285 32077
rect 36911 31991 36925 32005
rect 36935 31991 36949 32005
rect 36959 31991 36973 32005
rect 36983 31991 36997 32005
rect 37007 31991 37021 32005
rect 37031 31991 37045 32005
rect 37055 31991 37069 32005
rect 37079 31991 37093 32005
rect 37103 31991 37117 32005
rect 37127 31991 37141 32005
rect 37151 31991 37165 32005
rect 37175 31991 37189 32005
rect 37199 31991 37213 32005
rect 37223 31991 37237 32005
rect 37247 31991 37261 32005
rect 36911 30935 36925 30949
rect 36935 30935 36949 30949
rect 36959 30935 36973 30949
rect 36983 30935 36997 30949
rect 37007 30935 37021 30949
rect 37031 30935 37045 30949
rect 37055 30935 37069 30949
rect 37079 30935 37093 30949
rect 37103 30935 37117 30949
rect 37127 30935 37141 30949
rect 37151 30935 37165 30949
rect 37175 30935 37189 30949
rect 37199 30935 37213 30949
rect 37223 30935 37237 30949
rect 41447 35735 41461 35749
rect 41471 35735 41485 35749
rect 41399 35711 41413 35725
rect 41447 35687 41461 35701
rect 41471 35687 41485 35701
rect 41399 31199 41413 31213
rect 41423 31199 41437 31213
rect 41447 31199 41461 31213
rect 41471 31199 41485 31213
rect 41447 31151 41461 31165
rect 41399 31127 41413 31141
rect 41423 31127 41437 31141
rect 41471 31103 41485 31117
rect 41375 31031 41389 31045
rect 41399 31031 41413 31045
rect 41423 31031 41437 31045
rect 41447 31031 41461 31045
rect 37223 30887 37237 30901
rect 36911 30815 36925 30829
rect 36935 30815 36949 30829
rect 36959 30815 36973 30829
rect 36983 30815 36997 30829
rect 37007 30815 37021 30829
rect 37031 30815 37045 30829
rect 37055 30815 37069 30829
rect 37079 30815 37093 30829
rect 37103 30815 37117 30829
rect 37127 30815 37141 30829
rect 37151 30815 37165 30829
rect 37175 30815 37189 30829
rect 37199 30815 37213 30829
rect 36911 29759 36925 29773
rect 36935 29759 36949 29773
rect 36959 29759 36973 29773
rect 36983 29759 36997 29773
rect 37007 29759 37021 29773
rect 37031 29759 37045 29773
rect 37055 29759 37069 29773
rect 37079 29759 37093 29773
rect 37103 29759 37117 29773
rect 37127 29759 37141 29773
rect 37151 29759 37165 29773
rect 37175 29759 37189 29773
rect 37199 29759 37213 29773
rect 41375 30983 41389 30997
rect 41399 30983 41413 30997
rect 41423 30983 41437 30997
rect 41447 30983 41461 30997
rect 36911 29639 36925 29653
rect 36935 29639 36949 29653
rect 36959 29639 36973 29653
rect 36983 29639 36997 29653
rect 37007 29639 37021 29653
rect 37031 29639 37045 29653
rect 37055 29639 37069 29653
rect 37079 29639 37093 29653
rect 37103 29639 37117 29653
rect 37127 29639 37141 29653
rect 37151 29639 37165 29653
rect 37175 29639 37189 29653
rect 37199 29639 37213 29653
rect 36911 28583 36925 28597
rect 36935 28583 36949 28597
rect 36959 28583 36973 28597
rect 36983 28583 36997 28597
rect 37007 28583 37021 28597
rect 37031 28583 37045 28597
rect 37055 28583 37069 28597
rect 37079 28583 37093 28597
rect 37103 28583 37117 28597
rect 37127 28583 37141 28597
rect 37151 28583 37165 28597
rect 37175 28583 37189 28597
rect 37199 28583 37213 28597
rect 36911 28463 36925 28477
rect 36935 28463 36949 28477
rect 36959 28463 36973 28477
rect 36983 28463 36997 28477
rect 37007 28463 37021 28477
rect 37031 28463 37045 28477
rect 37055 28463 37069 28477
rect 37079 28463 37093 28477
rect 37103 28463 37117 28477
rect 37127 28463 37141 28477
rect 37151 28463 37165 28477
rect 37175 28463 37189 28477
rect 37199 28463 37213 28477
rect 36911 27407 36925 27421
rect 36935 27407 36949 27421
rect 36959 27407 36973 27421
rect 36983 27407 36997 27421
rect 37007 27407 37021 27421
rect 37031 27407 37045 27421
rect 37055 27407 37069 27421
rect 37079 27407 37093 27421
rect 37103 27407 37117 27421
rect 37127 27407 37141 27421
rect 37151 27407 37165 27421
rect 37175 27407 37189 27421
rect 37199 27407 37213 27421
rect 36911 27287 36925 27301
rect 36935 27287 36949 27301
rect 36959 27287 36973 27301
rect 36983 27287 36997 27301
rect 37007 27287 37021 27301
rect 37031 27287 37045 27301
rect 37055 27287 37069 27301
rect 37079 27287 37093 27301
rect 37103 27287 37117 27301
rect 37127 27287 37141 27301
rect 37151 27287 37165 27301
rect 37175 27287 37189 27301
rect 37199 27287 37213 27301
rect 36911 26231 36925 26245
rect 41495 26303 41509 26317
rect 36959 26255 36973 26269
rect 36983 26255 36997 26269
rect 37007 26255 37021 26269
rect 37031 26255 37045 26269
rect 37055 26255 37069 26269
rect 37079 26255 37093 26269
rect 37103 26255 37117 26269
rect 37127 26255 37141 26269
rect 37151 26255 37165 26269
rect 37175 26255 37189 26269
rect 36959 26207 36973 26221
rect 36983 26207 36997 26221
rect 37007 26207 37021 26221
rect 37031 26207 37045 26221
rect 37055 26207 37069 26221
rect 37079 26207 37093 26221
rect 37103 26207 37117 26221
rect 37127 26207 37141 26221
rect 36935 26159 36949 26173
rect 36959 26159 36973 26173
rect 36983 26159 36997 26173
rect 37007 26159 37021 26173
rect 37031 26159 37045 26173
rect 37055 26159 37069 26173
rect 37079 26159 37093 26173
rect 37103 26159 37117 26173
rect 37199 26183 37213 26197
rect 36911 26111 36925 26125
rect 36935 26111 36949 26125
rect 36959 26111 36973 26125
rect 36983 26111 36997 26125
rect 37007 26111 37021 26125
rect 37031 26111 37045 26125
rect 37055 26111 37069 26125
rect 37079 26111 37093 26125
rect 37103 26111 37117 26125
rect 36911 25055 36925 25069
rect 36935 25055 36949 25069
rect 36959 25055 36973 25069
rect 37151 26135 37165 26149
rect 37175 26135 37189 26149
rect 37199 26135 37213 26149
rect 37007 25079 37021 25093
rect 37031 25079 37045 25093
rect 37055 25079 37069 25093
rect 37079 25079 37093 25093
rect 37103 25079 37117 25093
rect 37127 25079 37141 25093
rect 37151 25079 37165 25093
rect 37175 25079 37189 25093
rect 37199 25079 37213 25093
rect 37223 25079 37237 25093
rect 36935 25007 36949 25021
rect 36983 25007 36997 25021
rect 37247 25007 37261 25021
rect 36911 24935 36925 24949
rect 36959 24959 36973 24973
rect 36983 24959 36997 24973
rect 37007 24959 37021 24973
rect 37031 24959 37045 24973
rect 37055 24959 37069 24973
rect 37079 24959 37093 24973
rect 37103 24959 37117 24973
rect 37127 24959 37141 24973
rect 37151 24959 37165 24973
rect 37175 24959 37189 24973
rect 37199 24959 37213 24973
rect 37223 24959 37237 24973
rect 37247 24959 37261 24973
rect 36911 23879 36925 23893
rect 36935 23879 36949 23893
rect 36983 23903 36997 23917
rect 37007 23903 37021 23917
rect 37031 23903 37045 23917
rect 37055 23903 37069 23917
rect 37079 23903 37093 23917
rect 37103 23903 37117 23917
rect 37127 23903 37141 23917
rect 37151 23903 37165 23917
rect 37175 23903 37189 23917
rect 37199 23903 37213 23917
rect 37223 23903 37237 23917
rect 37247 23903 37261 23917
rect 37271 23903 37285 23917
rect 36983 23855 36997 23869
rect 37007 23855 37021 23869
rect 36959 23807 36973 23821
rect 36983 23807 36997 23821
rect 37295 23831 37309 23845
rect 36911 23759 36925 23773
rect 36935 23759 36949 23773
rect 36959 23759 36973 23773
rect 36983 23759 36997 23773
rect 37031 23783 37045 23797
rect 37055 23783 37069 23797
rect 37079 23783 37093 23797
rect 37103 23783 37117 23797
rect 37127 23783 37141 23797
rect 37151 23783 37165 23797
rect 37175 23783 37189 23797
rect 37199 23783 37213 23797
rect 37223 23783 37237 23797
rect 37247 23783 37261 23797
rect 37271 23783 37285 23797
rect 37295 23783 37309 23797
rect 36911 22703 36925 22717
rect 36935 22703 36949 22717
rect 36959 22703 36973 22717
rect 36983 22703 36997 22717
rect 37007 22703 37021 22717
rect 37031 22703 37045 22717
rect 37079 22727 37093 22741
rect 37103 22727 37117 22741
rect 37127 22727 37141 22741
rect 37151 22727 37165 22741
rect 37175 22727 37189 22741
rect 37199 22727 37213 22741
rect 37223 22727 37237 22741
rect 37247 22727 37261 22741
rect 37271 22727 37285 22741
rect 37295 22727 37309 22741
rect 37319 22727 37333 22741
rect 37079 22679 37093 22693
rect 37055 22631 37069 22645
rect 37343 22655 37357 22669
rect 36911 22583 36925 22597
rect 36935 22583 36949 22597
rect 36959 22583 36973 22597
rect 36983 22583 36997 22597
rect 37007 22583 37021 22597
rect 37031 22583 37045 22597
rect 37055 22583 37069 22597
rect 37103 22607 37117 22621
rect 37127 22607 37141 22621
rect 37151 22607 37165 22621
rect 37175 22607 37189 22621
rect 37199 22607 37213 22621
rect 37223 22607 37237 22621
rect 37247 22607 37261 22621
rect 37271 22607 37285 22621
rect 37295 22607 37309 22621
rect 37319 22607 37333 22621
rect 37343 22607 37357 22621
rect 36911 21527 36925 21541
rect 36935 21527 36949 21541
rect 36959 21527 36973 21541
rect 36983 21527 36997 21541
rect 37007 21527 37021 21541
rect 37031 21527 37045 21541
rect 37055 21527 37069 21541
rect 37079 21527 37093 21541
rect 37127 21551 37141 21565
rect 37151 21551 37165 21565
rect 37175 21551 37189 21565
rect 37199 21551 37213 21565
rect 37223 21551 37237 21565
rect 37247 21551 37261 21565
rect 37271 21551 37285 21565
rect 37295 21551 37309 21565
rect 37319 21551 37333 21565
rect 37343 21551 37357 21565
rect 37367 21551 37381 21565
rect 36911 21479 36925 21493
rect 37103 21479 37117 21493
rect 37391 21479 37405 21493
rect 36935 21431 36949 21445
rect 36959 21431 36973 21445
rect 36983 21431 36997 21445
rect 37007 21431 37021 21445
rect 37031 21431 37045 21445
rect 37055 21431 37069 21445
rect 37079 21431 37093 21445
rect 37103 21431 37117 21445
rect 37127 21431 37141 21445
rect 37151 21431 37165 21445
rect 37175 21431 37189 21445
rect 37199 21431 37213 21445
rect 37223 21431 37237 21445
rect 37247 21431 37261 21445
rect 37271 21431 37285 21445
rect 37295 21431 37309 21445
rect 37319 21431 37333 21445
rect 37343 21431 37357 21445
rect 37367 21431 37381 21445
rect 37391 21431 37405 21445
rect 36911 20351 36925 20365
rect 36935 20351 36949 20365
rect 36959 20351 36973 20365
rect 36983 20351 36997 20365
rect 37007 20351 37021 20365
rect 37031 20351 37045 20365
rect 37055 20351 37069 20365
rect 37079 20351 37093 20365
rect 37103 20351 37117 20365
rect 37127 20351 37141 20365
rect 37151 20351 37165 20365
rect 37175 20351 37189 20365
rect 37199 20351 37213 20365
rect 37223 20351 37237 20365
rect 37247 20351 37261 20365
rect 37295 20375 37309 20389
rect 37319 20375 37333 20389
rect 37343 20375 37357 20389
rect 37367 20375 37381 20389
rect 37391 20375 37405 20389
rect 37415 20375 37429 20389
rect 37175 20303 37189 20317
rect 37271 20303 37285 20317
rect 37439 20303 37453 20317
rect 36911 20231 36925 20245
rect 36935 20231 36949 20245
rect 36959 20231 36973 20245
rect 36983 20231 36997 20245
rect 37007 20231 37021 20245
rect 37031 20231 37045 20245
rect 37055 20231 37069 20245
rect 37079 20231 37093 20245
rect 37103 20231 37117 20245
rect 37127 20231 37141 20245
rect 37151 20231 37165 20245
rect 36911 19175 36925 19189
rect 36935 19175 36949 19189
rect 36959 19175 36973 19189
rect 36983 19175 36997 19189
rect 37007 19175 37021 19189
rect 37031 19175 37045 19189
rect 37199 20255 37213 20269
rect 37223 20255 37237 20269
rect 37247 20255 37261 20269
rect 37271 20255 37285 20269
rect 37295 20255 37309 20269
rect 37319 20255 37333 20269
rect 37343 20255 37357 20269
rect 37367 20255 37381 20269
rect 37391 20255 37405 20269
rect 37415 20255 37429 20269
rect 37439 20255 37453 20269
rect 37079 19199 37093 19213
rect 37103 19199 37117 19213
rect 37127 19199 37141 19213
rect 37151 19199 37165 19213
rect 37175 19199 37189 19213
rect 37199 19199 37213 19213
rect 37223 19199 37237 19213
rect 37247 19199 37261 19213
rect 37271 19199 37285 19213
rect 37295 19199 37309 19213
rect 37319 19199 37333 19213
rect 37343 19199 37357 19213
rect 37367 19199 37381 19213
rect 37391 19199 37405 19213
rect 37415 19199 37429 19213
rect 37439 19199 37453 19213
rect 37463 19199 37477 19213
rect 37031 19127 37045 19141
rect 37055 19127 37069 19141
rect 37487 19127 37501 19141
rect 36911 19055 36925 19069
rect 36935 19055 36949 19069
rect 36959 19055 36973 19069
rect 36983 19055 36997 19069
rect 37007 19055 37021 19069
rect 37055 19079 37069 19093
rect 37079 19079 37093 19093
rect 37103 19079 37117 19093
rect 37127 19079 37141 19093
rect 37151 19079 37165 19093
rect 37175 19079 37189 19093
rect 37199 19079 37213 19093
rect 37223 19079 37237 19093
rect 37247 19079 37261 19093
rect 37271 19079 37285 19093
rect 37295 19079 37309 19093
rect 37319 19079 37333 19093
rect 37343 19079 37357 19093
rect 37367 19079 37381 19093
rect 37391 19079 37405 19093
rect 37415 19079 37429 19093
rect 37439 19079 37453 19093
rect 37463 19079 37477 19093
rect 37487 19079 37501 19093
rect 36935 18023 36949 18037
rect 36959 18023 36973 18037
rect 36983 18023 36997 18037
rect 37007 18023 37021 18037
rect 37031 18023 37045 18037
rect 37055 18023 37069 18037
rect 37079 18023 37093 18037
rect 37103 18023 37117 18037
rect 37127 18023 37141 18037
rect 37151 18023 37165 18037
rect 37175 18023 37189 18037
rect 37199 18023 37213 18037
rect 37223 18023 37237 18037
rect 37247 18023 37261 18037
rect 37271 18023 37285 18037
rect 37295 18023 37309 18037
rect 37319 18023 37333 18037
rect 37343 18023 37357 18037
rect 37367 18023 37381 18037
rect 37391 18023 37405 18037
rect 37415 18023 37429 18037
rect 37439 18023 37453 18037
rect 37463 18023 37477 18037
rect 37487 18023 37501 18037
rect 37511 18023 37525 18037
rect 36935 17975 36949 17989
rect 36959 17975 36973 17989
rect 36983 17975 36997 17989
rect 37007 17975 37021 17989
rect 37031 17975 37045 17989
rect 37055 17975 37069 17989
rect 37079 17975 37093 17989
rect 37103 17975 37117 17989
rect 37127 17975 37141 17989
rect 37151 17975 37165 17989
rect 37175 17975 37189 17989
rect 37199 17975 37213 17989
rect 37223 17975 37237 17989
rect 37247 17975 37261 17989
rect 37271 17975 37285 17989
rect 37295 17975 37309 17989
rect 37319 17975 37333 17989
rect 37343 17975 37357 17989
rect 37367 17975 37381 17989
rect 37391 17975 37405 17989
rect 37415 17975 37429 17989
rect 37439 17975 37453 17989
rect 36911 17927 36925 17941
rect 36935 17927 36949 17941
rect 36959 17927 36973 17941
rect 36983 17927 36997 17941
rect 37007 17927 37021 17941
rect 37031 17927 37045 17941
rect 37055 17927 37069 17941
rect 37079 17927 37093 17941
rect 37103 17927 37117 17941
rect 37127 17927 37141 17941
rect 37151 17927 37165 17941
rect 37175 17927 37189 17941
rect 37199 17927 37213 17941
rect 37223 17927 37237 17941
rect 37247 17927 37261 17941
rect 37271 17927 37285 17941
rect 37295 17927 37309 17941
rect 37319 17927 37333 17941
rect 37343 17927 37357 17941
rect 37367 17927 37381 17941
rect 37391 17927 37405 17941
rect 37415 17927 37429 17941
rect 37535 17951 37549 17965
rect 36911 17879 36925 17893
rect 36935 17879 36949 17893
rect 36959 17879 36973 17893
rect 36983 17879 36997 17893
rect 37007 17879 37021 17893
rect 37031 17879 37045 17893
rect 37055 17879 37069 17893
rect 37079 17879 37093 17893
rect 37103 17879 37117 17893
rect 37127 17879 37141 17893
rect 37151 17879 37165 17893
rect 37175 17879 37189 17893
rect 37199 17879 37213 17893
rect 37223 17879 37237 17893
rect 37247 17879 37261 17893
rect 37271 17879 37285 17893
rect 37295 17879 37309 17893
rect 37319 17879 37333 17893
rect 37343 17879 37357 17893
rect 37367 17879 37381 17893
rect 37391 17879 37405 17893
rect 37415 17879 37429 17893
rect 36911 16823 36925 16837
rect 36935 16823 36949 16837
rect 36959 16823 36973 16837
rect 36983 16823 36997 16837
rect 37007 16823 37021 16837
rect 37031 16823 37045 16837
rect 37055 16823 37069 16837
rect 37079 16823 37093 16837
rect 37103 16823 37117 16837
rect 37463 17903 37477 17917
rect 37487 17903 37501 17917
rect 37511 17903 37525 17917
rect 37535 17903 37549 17917
rect 41471 16943 41485 16957
rect 41471 16895 41485 16909
rect 37151 16847 37165 16861
rect 37175 16847 37189 16861
rect 37199 16847 37213 16861
rect 37223 16847 37237 16861
rect 37247 16847 37261 16861
rect 37271 16847 37285 16861
rect 37295 16847 37309 16861
rect 37319 16847 37333 16861
rect 37343 16847 37357 16861
rect 37367 16847 37381 16861
rect 37391 16847 37405 16861
rect 37415 16847 37429 16861
rect 37439 16847 37453 16861
rect 37463 16847 37477 16861
rect 37487 16847 37501 16861
rect 37511 16847 37525 16861
rect 37535 16847 37549 16861
rect 37031 16775 37045 16789
rect 37127 16775 37141 16789
rect 41471 16799 41485 16813
rect 36911 16703 36925 16717
rect 36935 16703 36949 16717
rect 36959 16703 36973 16717
rect 36983 16703 36997 16717
rect 37007 16703 37021 16717
rect 7535 16607 7549 16621
rect 11327 16607 11341 16621
rect 11351 16607 11365 16621
rect 11375 16607 11389 16621
rect 11399 16607 11413 16621
rect 11903 16607 11917 16621
rect 12107 16607 12121 16621
rect 13367 16607 13381 16621
rect 13559 16607 13573 16621
rect 14351 16607 14365 16621
rect 14903 16607 14917 16621
rect 15119 16607 15133 16621
rect 15863 16607 15877 16621
rect 16031 16607 16045 16621
rect 16415 16607 16429 16621
rect 16607 16607 16621 16621
rect 16823 16607 16837 16621
rect 17567 16607 17581 16621
rect 17735 16607 17749 16621
rect 27143 16607 27157 16621
rect 27335 16607 27349 16621
rect 27575 16607 27589 16621
rect 35279 16607 35293 16621
rect 36911 16607 36925 16621
rect 36935 16607 36949 16621
rect 36959 16607 36973 16621
rect 36983 16607 36997 16621
rect 37055 16727 37069 16741
rect 37079 16727 37093 16741
rect 37103 16727 37117 16741
rect 37127 16727 37141 16741
rect 37151 16727 37165 16741
rect 37175 16727 37189 16741
rect 37199 16727 37213 16741
rect 37223 16727 37237 16741
rect 37247 16727 37261 16741
rect 37271 16727 37285 16741
rect 37295 16727 37309 16741
rect 37319 16727 37333 16741
rect 37343 16727 37357 16741
rect 37367 16727 37381 16741
rect 37391 16727 37405 16741
rect 37415 16727 37429 16741
rect 37439 16727 37453 16741
rect 37463 16727 37477 16741
rect 37487 16727 37501 16741
rect 37511 16727 37525 16741
rect 37535 16727 37549 16741
rect 41471 16751 41485 16765
rect 37031 16631 37045 16645
rect 37055 16631 37069 16645
rect 37079 16631 37093 16645
rect 37103 16631 37117 16645
rect 37127 16631 37141 16645
rect 37151 16631 37165 16645
rect 37175 16631 37189 16645
rect 37199 16631 37213 16645
rect 37223 16631 37237 16645
rect 37247 16631 37261 16645
rect 37271 16631 37285 16645
rect 37295 16631 37309 16645
rect 37319 16631 37333 16645
rect 37343 16631 37357 16645
rect 37367 16631 37381 16645
rect 37391 16631 37405 16645
rect 37415 16631 37429 16645
rect 37439 16631 37453 16645
rect 37463 16631 37477 16645
rect 37487 16631 37501 16645
rect 37511 16631 37525 16645
rect 37535 16631 37549 16645
rect 37559 16631 37573 16645
rect 11927 16583 11941 16597
rect 11423 16559 11437 16573
rect 11639 16559 11653 16573
rect 12035 16559 12049 16573
rect 12059 16559 12073 16573
rect 12083 16559 12097 16573
rect 7535 16511 7549 16525
rect 11327 16511 11341 16525
rect 11351 16511 11365 16525
rect 11375 16511 11389 16525
rect 11399 16511 11413 16525
rect 11423 16511 11437 16525
rect 11450 16511 11464 16525
rect 11496 16511 11510 16525
rect 11542 16511 11556 16525
rect 11588 16511 11602 16525
rect 11639 16511 11653 16525
rect 11279 16007 11293 16021
rect 11255 15983 11269 15997
rect 11231 15959 11245 15973
rect 11399 15959 11413 15973
rect 11423 15959 11437 15973
rect 11472 16484 11486 16498
rect 11519 16484 11533 16498
rect 11565 16484 11579 16498
rect 11611 16484 11625 16498
rect 11639 16151 11653 16165
rect 11927 16487 11941 16501
rect 11663 16127 11677 16141
rect 11749 16127 11763 16141
rect 11773 16127 11787 16141
rect 11797 16127 11811 16141
rect 11831 16103 11845 16117
rect 11855 16079 11869 16093
rect 11879 16055 11893 16069
rect 13847 16079 13861 16093
rect 14711 16079 14725 16093
rect 15575 16103 15589 16117
rect 16415 16151 16429 16165
rect 16991 16175 17005 16189
rect 18167 16199 18181 16213
rect 18191 16175 18205 16189
rect 19895 16151 19909 16165
rect 20759 16127 20773 16141
rect 21191 16103 21205 16117
rect 22127 16079 22141 16093
rect 20735 16055 20749 16069
rect 20759 16055 20773 16069
rect 22895 16055 22909 16069
rect 16967 16031 16981 16045
rect 16991 16031 17005 16045
rect 23927 16031 23941 16045
rect 18143 16007 18157 16021
rect 18167 16007 18181 16021
rect 24239 16007 24253 16021
rect 18167 15983 18181 15997
rect 18191 15983 18205 15997
rect 25823 15983 25837 15997
rect 19871 15959 19885 15973
rect 19895 15959 19909 15973
rect 26783 15959 26797 15973
rect 27143 15959 27157 15973
rect 27671 15983 27685 15997
rect 35305 16583 35319 16597
rect 36239 16583 36253 16597
rect 36263 16583 36277 16597
rect 36287 16583 36301 16597
rect 36023 16559 36037 16573
rect 36311 16559 36325 16573
rect 36383 16559 36397 16573
rect 37007 16559 37021 16573
rect 37583 16559 37597 16573
rect 36167 16535 36181 16549
rect 36287 16535 36301 16549
rect 35305 16511 35319 16525
rect 36215 16511 36229 16525
rect 36239 16511 36253 16525
rect 36263 16511 36277 16525
rect 36719 16511 36733 16525
rect 38591 16511 38605 16525
rect 38855 16487 38869 16501
rect 36911 16463 36925 16477
rect 36935 16463 36949 16477
rect 36959 16463 36973 16477
rect 36983 16463 36997 16477
rect 37007 16463 37021 16477
rect 37031 16463 37045 16477
rect 37055 16463 37069 16477
rect 37079 16463 37093 16477
rect 37103 16463 37117 16477
rect 37127 16463 37141 16477
rect 37151 16463 37165 16477
rect 37175 16463 37189 16477
rect 37199 16463 37213 16477
rect 37223 16463 37237 16477
rect 37247 16463 37261 16477
rect 37271 16463 37285 16477
rect 37295 16463 37309 16477
rect 37319 16463 37333 16477
rect 37343 16463 37357 16477
rect 37367 16463 37381 16477
rect 37391 16463 37405 16477
rect 37415 16463 37429 16477
rect 37439 16463 37453 16477
rect 37463 16463 37477 16477
rect 37487 16463 37501 16477
rect 37511 16463 37525 16477
rect 37535 16463 37549 16477
rect 37559 16463 37573 16477
rect 37583 16463 37597 16477
rect 39167 16463 39181 16477
rect 28511 15959 28525 15973
rect 32759 15959 32773 15973
rect 33599 15959 33613 15973
rect 35281 15959 35295 15973
rect 35305 15959 35319 15973
rect 36167 15959 36181 15973
rect 36911 15959 36925 15973
rect 36935 15959 36949 15973
rect 36959 15959 36973 15973
rect 36983 15959 36997 15973
rect 37007 15959 37021 15973
rect 11183 15935 11197 15949
rect 11279 15935 11293 15949
rect 11303 15935 11317 15949
rect 39191 16439 39205 16453
rect 39215 16415 39229 16429
rect 39239 16391 39253 16405
rect 39263 16367 39277 16381
rect 39287 16343 39301 16357
rect 39311 16319 39325 16333
rect 39335 16295 39349 16309
rect 39359 16271 39373 16285
rect 39383 16247 39397 16261
rect 39407 16223 39421 16237
rect 39431 16199 39445 16213
rect 39455 16175 39469 16189
rect 39479 16151 39493 16165
rect 39503 16127 39517 16141
rect 39527 16103 39541 16117
rect 39551 16079 39565 16093
rect 39575 16055 39589 16069
rect 39647 16031 39661 16045
rect 39671 16007 39685 16021
rect 39695 15983 39709 15997
rect 39743 15959 39757 15973
rect 39791 15935 39805 15949
rect 7535 15911 7549 15925
rect 11135 15911 11149 15925
rect 11399 15911 11413 15925
rect 11423 15911 11437 15925
rect 11725 15911 11739 15925
rect 11855 15911 11869 15925
rect 11879 15911 11893 15925
rect 16391 15911 16405 15925
rect 16415 15911 16429 15925
rect 26759 15911 26773 15925
rect 27143 15911 27157 15925
rect 30193 15911 30207 15925
rect 32759 15911 32773 15925
rect 33599 15911 33613 15925
rect 36167 15911 36181 15925
rect 36911 15911 36925 15925
rect 36935 15911 36949 15925
rect 36959 15911 36973 15925
rect 36983 15911 36997 15925
rect 41375 15911 41389 15925
rect 11749 15887 11763 15901
rect 15551 15887 15565 15901
rect 15575 15887 15589 15901
rect 23903 15887 23917 15901
rect 23927 15887 23941 15901
rect 27647 15887 27661 15901
rect 27671 15887 27685 15901
rect 30218 15887 30232 15901
rect 7463 15863 7477 15877
rect 11591 15863 11605 15877
rect 11639 15863 11653 15877
rect 11663 15863 11677 15877
rect 13823 15863 13837 15877
rect 13847 15863 13861 15877
rect 21167 15863 21181 15877
rect 21191 15863 21205 15877
rect 24215 15863 24229 15877
rect 24239 15863 24253 15877
rect 28487 15863 28501 15877
rect 28511 15863 28525 15877
rect 31607 15863 31621 15877
rect 7463 15815 7477 15829
rect 7535 15815 7549 15829
rect 11135 15815 11149 15829
rect 11183 15815 11197 15829
rect 11231 15815 11245 15829
rect 11255 15815 11269 15829
rect 11303 15839 11317 15853
rect 11773 15839 11787 15853
rect 11831 15839 11845 15853
rect 14711 15839 14725 15853
rect 22127 15839 22141 15853
rect 22895 15839 22909 15853
rect 25823 15839 25837 15853
rect 30218 15839 30232 15853
rect 41423 15887 41437 15901
rect 41447 15863 41461 15877
rect 14687 15815 14701 15829
rect 22103 15815 22117 15829
rect 22871 15815 22885 15829
rect 25799 15815 25813 15829
rect 30169 15815 30183 15829
rect 31895 15815 31909 15829
rect 32759 15815 32773 15829
rect 33599 15815 33613 15829
rect 36167 15815 36181 15829
rect 39167 15815 39181 15829
rect 39191 15815 39205 15829
rect 39215 15815 39229 15829
rect 39239 15815 39253 15829
rect 39263 15815 39277 15829
rect 39287 15815 39301 15829
rect 39311 15815 39325 15829
rect 39335 15815 39349 15829
rect 39359 15815 39373 15829
rect 39383 15815 39397 15829
rect 39407 15815 39421 15829
rect 39431 15815 39445 15829
rect 39455 15815 39469 15829
rect 39479 15815 39493 15829
rect 39503 15815 39517 15829
rect 39527 15815 39541 15829
rect 39551 15815 39565 15829
rect 39575 15815 39589 15829
rect 11183 15695 11197 15709
rect 11231 15695 11245 15709
rect 11255 15695 11269 15709
rect 11279 15695 11293 15709
rect 11303 15695 11317 15709
rect 11327 15695 11341 15709
rect 11351 15673 11365 15687
rect 11183 15649 11197 15663
rect 11351 15649 11365 15663
rect 11231 15623 11245 15637
rect 11255 15623 11269 15637
rect 11279 15623 11293 15637
rect 11303 15623 11317 15637
rect 11327 15623 11341 15637
rect 6503 12215 6517 12229
rect 7463 12215 7477 12229
rect 7535 12215 7549 12229
rect 11231 12215 11245 12229
rect 11255 12215 11269 12229
rect 11279 12215 11293 12229
rect 11303 12215 11317 12229
rect 39167 15601 39181 15615
rect 39191 15601 39205 15615
rect 39215 15601 39229 15615
rect 39239 15601 39253 15615
rect 39263 15601 39277 15615
rect 39143 15577 39157 15591
rect 39311 15577 39325 15591
rect 39335 15577 39349 15591
rect 39359 15577 39373 15591
rect 39383 15577 39397 15591
rect 39143 15553 39157 15567
rect 39647 15815 39661 15829
rect 39671 15815 39685 15829
rect 39695 15815 39709 15829
rect 39743 15815 39757 15829
rect 39791 15815 39805 15829
rect 41375 15815 41389 15829
rect 41423 15815 41437 15829
rect 41447 15815 41461 15829
rect 39431 15553 39445 15567
rect 39455 15553 39469 15567
rect 39479 15553 39493 15567
rect 39503 15553 39517 15567
rect 39527 15553 39541 15567
rect 39551 15553 39565 15567
rect 39575 15553 39589 15567
rect 39599 15553 39613 15567
rect 39623 15553 39637 15567
rect 39143 15529 39157 15543
rect 39143 15505 39157 15519
rect 39431 15505 39445 15519
rect 39455 15505 39469 15519
rect 39479 15505 39493 15519
rect 39503 15505 39517 15519
rect 39527 15505 39541 15519
rect 39551 15505 39565 15519
rect 39575 15505 39589 15519
rect 39599 15505 39613 15519
rect 39623 15505 39637 15519
rect 39143 15481 39157 15495
rect 39383 15481 39397 15495
rect 39167 15457 39181 15471
rect 39191 15457 39205 15471
rect 39215 15457 39229 15471
rect 39239 15457 39253 15471
rect 39263 15457 39277 15471
rect 39311 15457 39325 15471
rect 39335 15457 39349 15471
rect 39359 15457 39373 15471
rect 6503 12167 6517 12181
rect 7463 12167 7477 12181
rect 7535 12167 7549 12181
rect 11231 12167 11245 12181
rect 11255 12167 11269 12181
rect 11279 12167 11293 12181
rect 11303 12167 11317 12181
rect 11231 11598 11245 11612
rect 11255 11598 11269 11612
rect 11279 11598 11293 11612
rect 11303 11598 11317 11612
rect 11351 11576 11365 11590
rect 11231 11543 11245 11557
rect 11255 11543 11269 11557
rect 11279 11552 11293 11566
rect 11351 11552 11365 11566
rect 11303 11519 11317 11533
rect 39167 10487 39181 10501
rect 39191 10487 39205 10501
rect 39215 10487 39229 10501
rect 39239 10487 39253 10501
rect 39263 10487 39277 10501
rect 39311 10487 39325 10501
rect 39335 10487 39349 10501
rect 39359 10487 39373 10501
rect 39455 10487 39469 10501
rect 39479 10487 39493 10501
rect 39503 10487 39517 10501
rect 39527 10487 39541 10501
rect 39143 10463 39157 10477
rect 39167 10439 39181 10453
rect 39191 10439 39205 10453
rect 39215 10439 39229 10453
rect 39239 10439 39253 10453
rect 39263 10439 39277 10453
rect 39311 10439 39325 10453
rect 39335 10439 39349 10453
rect 39359 10439 39373 10453
rect 39455 10439 39469 10453
rect 39479 10439 39493 10453
rect 39503 10439 39517 10453
rect 39527 10439 39541 10453
rect 39167 9247 39181 9261
rect 39191 9247 39205 9261
rect 39215 9247 39229 9261
rect 39239 9247 39253 9261
rect 39263 9247 39277 9261
rect 39311 9247 39325 9261
rect 39335 9247 39349 9261
rect 39143 9224 39157 9238
rect 39143 9200 39157 9214
rect 39143 9176 39157 9190
rect 39335 9175 39349 9189
rect 39167 9143 39181 9157
rect 39191 9143 39205 9157
rect 39215 9143 39229 9157
rect 39239 9143 39253 9157
rect 39263 9143 39277 9157
rect 39311 9143 39325 9157
rect 39167 8039 39181 8053
rect 39191 8039 39205 8053
rect 39215 8039 39229 8053
rect 39239 8039 39253 8053
rect 39263 8039 39277 8053
rect 39311 8039 39325 8053
rect 39479 8039 39493 8053
rect 39503 8039 39517 8053
rect 39143 8015 39157 8029
rect 39167 7991 39181 8005
rect 39191 7991 39205 8005
rect 39215 7991 39229 8005
rect 39239 7991 39253 8005
rect 39263 7991 39277 8005
rect 39311 7991 39325 8005
rect 39479 7991 39493 8005
rect 39503 7991 39517 8005
rect 7463 7679 7477 7693
rect 11231 7679 11245 7693
rect 11255 7679 11269 7693
rect 11303 7679 11317 7693
rect 39167 7679 39181 7693
rect 39191 7679 39205 7693
rect 39215 7679 39229 7693
rect 39239 7679 39253 7693
rect 39263 7679 39277 7693
rect 39311 7679 39325 7693
rect 39479 7679 39493 7693
rect 11351 7655 11365 7669
rect 39143 7647 39157 7661
rect 7463 7631 7477 7645
rect 11231 7631 11245 7645
rect 11255 7631 11269 7645
rect 11303 7631 11317 7645
rect 39143 7623 39157 7637
rect 39239 7623 39253 7637
rect 39575 7631 39589 7645
rect 39599 7631 39613 7645
rect 39143 7599 39157 7613
rect 11303 7559 11317 7573
rect 11807 7559 11821 7573
rect 39191 7568 39205 7582
rect 39215 7568 39229 7582
rect 11231 7511 11245 7525
rect 11255 7511 11269 7525
rect 7463 7487 7477 7501
rect 11231 7463 11245 7477
rect 11735 7511 11749 7525
rect 19367 7535 19381 7549
rect 22559 7535 22573 7549
rect 7463 7439 7477 7453
rect 11255 7439 11269 7453
rect 11303 7439 11317 7453
rect 11327 7439 11341 7453
rect 7463 6551 7477 6565
rect 11303 6575 11317 6589
rect 11327 6575 11341 6589
rect 11327 6527 11341 6541
rect 19367 7487 19381 7501
rect 15815 7439 15829 7453
rect 25823 7511 25837 7525
rect 35303 7511 35317 7525
rect 36455 7511 36469 7525
rect 41423 12215 41437 12229
rect 41447 12215 41461 12229
rect 41423 12167 41437 12181
rect 41447 12167 41461 12181
rect 39671 7535 39685 7549
rect 39695 7535 39709 7549
rect 39743 7535 39757 7549
rect 39791 7535 39805 7549
rect 41423 7535 41437 7549
rect 36503 7487 36517 7501
rect 39479 7487 39493 7501
rect 39671 7487 39685 7501
rect 39695 7487 39709 7501
rect 39743 7487 39757 7501
rect 39791 7487 39805 7501
rect 41423 7487 41437 7501
rect 41471 7487 41485 7501
rect 19799 7463 19813 7477
rect 19943 7463 19957 7477
rect 25823 7463 25837 7477
rect 28199 7463 28213 7477
rect 32183 7463 32197 7477
rect 36479 7463 36493 7477
rect 39263 7463 39277 7477
rect 39311 7415 39325 7429
rect 39599 7415 39613 7429
rect 15815 7391 15829 7405
rect 19799 7391 19813 7405
rect 19943 7391 19957 7405
rect 22559 7391 22573 7405
rect 36455 7391 36469 7405
rect 36503 7391 36517 7405
rect 39167 7391 39181 7405
rect 39191 7391 39205 7405
rect 39695 7367 39709 7381
rect 39743 7367 39757 7381
rect 25823 7343 25837 7357
rect 36455 7343 36469 7357
rect 36479 7343 36493 7357
rect 41471 7439 41485 7453
rect 41471 7343 41485 7357
rect 39191 7319 39205 7333
rect 28199 7295 28213 7309
rect 32183 7295 32197 7309
rect 36455 7295 36469 7309
rect 39575 7295 39589 7309
rect 39695 7295 39709 7309
rect 39743 7295 39757 7309
rect 41471 7295 41485 7309
rect 39575 6623 39589 6637
rect 39695 6623 39709 6637
rect 39743 6623 39757 6637
rect 36455 6599 36469 6613
rect 36503 6599 36517 6613
rect 36311 6575 36325 6589
rect 36551 6575 36565 6589
rect 39695 6575 39709 6589
rect 39743 6575 39757 6589
rect 28199 6551 28213 6565
rect 32183 6551 32197 6565
rect 32327 6551 32341 6565
rect 7463 6503 7477 6517
rect 11303 6503 11317 6517
rect 11687 6527 11701 6541
rect 15671 6527 15685 6541
rect 15815 6527 15829 6541
rect 19799 6527 19813 6541
rect 19943 6527 19957 6541
rect 28055 6527 28069 6541
rect 11687 6479 11701 6493
rect 15671 6479 15685 6493
rect 15815 6479 15829 6493
rect 19799 6479 19813 6493
rect 19943 6479 19957 6493
rect 28055 6479 28069 6493
rect 28199 6479 28213 6493
rect 32183 6479 32197 6493
rect 32327 6479 32341 6493
rect 36503 6503 36517 6517
rect 36551 6527 36565 6541
rect 39575 6503 39589 6517
rect 36311 6479 36325 6493
rect 36455 6479 36469 6493
<< metal2 >>
rect 11376 41317 11388 41351
rect 11424 41293 11436 41375
rect 11472 41365 11484 41423
rect 11544 41341 11556 41399
rect 15600 41365 15612 41423
rect 19776 41389 19788 41423
rect 19920 41365 19932 41423
rect 28032 41365 28044 41423
rect 28176 41341 28188 41423
rect 32160 41317 32172 41423
rect 32304 41317 32316 41423
rect 36240 41317 36252 41375
rect 36264 41317 36276 41375
rect 36288 41269 36300 41375
rect 36312 41293 36324 41375
rect 36432 41293 36444 41423
rect 36720 41245 36732 41327
rect 36912 41245 36924 41351
rect 36936 41245 36948 41399
rect 36960 41245 36972 41327
rect 37008 41269 37020 41303
rect 41472 40429 41484 40463
rect 6528 40357 6540 40391
rect 7440 40357 7452 40391
rect 7536 40357 7548 40391
rect 19920 37645 19932 37679
rect 15600 37525 15612 37559
rect 16968 37429 16980 37463
rect 18024 37429 18036 37559
rect 19920 37429 19932 37559
rect 7536 37357 7548 37391
rect 11352 37285 11364 37319
rect 11376 37309 11388 37391
rect 11400 37261 11412 37391
rect 11424 37357 11436 37391
rect 11904 37222 11916 37295
rect 12037 37247 12048 37261
rect 15589 37247 15600 37261
rect 15816 37260 15828 37295
rect 16776 37260 16788 37367
rect 16968 37260 16980 37367
rect 18024 37260 18036 37367
rect 19920 37333 19932 37367
rect 15816 37248 15840 37260
rect 16776 37248 16800 37260
rect 16968 37248 16992 37260
rect 12036 37222 12048 37247
rect 15588 37222 15600 37247
rect 15828 37222 15840 37248
rect 16788 37222 16800 37248
rect 16980 37222 16992 37248
rect 18014 37248 18036 37260
rect 25992 37260 26004 37367
rect 26256 37260 26268 37463
rect 26976 37260 26988 37463
rect 28776 37260 28788 37559
rect 28968 37260 28980 37607
rect 29040 37260 29052 37367
rect 29136 37260 29148 37559
rect 32160 37309 32172 37679
rect 32304 37381 32316 37679
rect 36288 37381 36300 37631
rect 36312 37381 36324 37679
rect 36720 37285 36732 37679
rect 36912 37645 36924 37679
rect 36768 37309 36780 37631
rect 36960 37549 36972 37703
rect 36984 37549 36996 37703
rect 36912 37261 36924 37511
rect 36936 37261 36948 37511
rect 36960 37261 36972 37439
rect 36984 37261 36996 37487
rect 37008 37261 37020 37607
rect 37032 37453 37044 37703
rect 37056 37429 37068 37679
rect 37080 37621 37092 37655
rect 37032 37261 37044 37415
rect 37056 37261 37068 37391
rect 37080 37261 37092 37559
rect 37104 37405 37116 37631
rect 37104 37261 37116 37343
rect 37128 37261 37140 37607
rect 37152 37261 37164 37559
rect 37176 37501 37188 37535
rect 37176 37261 37188 37463
rect 37200 37261 37212 37511
rect 37224 37261 37236 37463
rect 37272 37381 37284 37439
rect 37248 37261 37260 37343
rect 37296 37309 37308 37415
rect 37272 37261 37284 37295
rect 37320 37285 37332 37367
rect 37344 37285 37356 37343
rect 37368 37285 37380 37319
rect 25992 37248 26017 37260
rect 26256 37248 26281 37260
rect 26976 37248 27001 37260
rect 28776 37248 28800 37260
rect 28968 37248 28992 37260
rect 29040 37248 29064 37260
rect 29136 37248 29160 37260
rect 18014 37222 18026 37248
rect 26005 37222 26017 37248
rect 26269 37222 26281 37248
rect 26989 37222 27001 37248
rect 28788 37222 28800 37248
rect 28980 37222 28992 37248
rect 29052 37222 29064 37248
rect 29148 37222 29160 37248
rect 36720 37222 36732 37247
rect 41424 35845 41436 35879
rect 41448 35845 41460 35927
rect 41472 35845 41484 35927
rect 6504 35629 6516 35663
rect 6528 35629 6540 35735
rect 41400 35725 41412 35759
rect 41448 35701 41460 35735
rect 41472 35701 41484 35735
rect 36912 34357 36924 34463
rect 36936 34357 36948 34463
rect 36960 34357 36972 34463
rect 36984 34357 36996 34463
rect 37008 34357 37020 34463
rect 37032 34357 37044 34463
rect 37056 34357 37068 34463
rect 37080 34357 37092 34463
rect 37104 34357 37116 34463
rect 37128 34357 37140 34463
rect 37152 34357 37164 34463
rect 37176 34357 37188 34463
rect 37200 34357 37212 34463
rect 37224 34357 37236 34463
rect 37248 34357 37260 34463
rect 37272 34357 37284 34463
rect 37296 34357 37308 34463
rect 37320 34357 37332 34463
rect 37344 34357 37356 34463
rect 37368 34429 37380 34463
rect 36912 33181 36924 33287
rect 36936 33181 36948 33287
rect 36960 33181 36972 33287
rect 36984 33181 36996 33287
rect 37008 33181 37020 33287
rect 37032 33181 37044 33287
rect 37056 33181 37068 33287
rect 37080 33181 37092 33287
rect 37104 33181 37116 33287
rect 37128 33181 37140 33287
rect 37152 33181 37164 33287
rect 37176 33181 37188 33287
rect 37200 33181 37212 33287
rect 37224 33181 37236 33287
rect 37248 33181 37260 33287
rect 37272 33181 37284 33287
rect 37296 33181 37308 33287
rect 37320 33253 37332 33287
rect 36912 32005 36924 32111
rect 36936 32005 36948 32111
rect 36960 32005 36972 32111
rect 36984 32005 36996 32111
rect 37008 32005 37020 32111
rect 37032 32005 37044 32111
rect 37056 32005 37068 32111
rect 37080 32005 37092 32111
rect 37104 32005 37116 32111
rect 37128 32005 37140 32111
rect 37152 32005 37164 32111
rect 37176 32005 37188 32111
rect 37200 32005 37212 32111
rect 37224 32005 37236 32111
rect 37248 32005 37260 32111
rect 37272 32077 37284 32111
rect 41400 31141 41412 31199
rect 41424 31141 41436 31199
rect 41448 31165 41460 31199
rect 41472 31117 41484 31199
rect 41376 30997 41388 31031
rect 41400 30997 41412 31031
rect 41424 30997 41436 31031
rect 41448 30997 41460 31031
rect 6504 30901 6516 30983
rect 6528 30901 6540 30983
rect 6552 30901 6564 30935
rect 36912 30829 36924 30935
rect 36936 30829 36948 30935
rect 36960 30829 36972 30935
rect 36984 30829 36996 30935
rect 37008 30829 37020 30935
rect 37032 30829 37044 30935
rect 37056 30829 37068 30935
rect 37080 30829 37092 30935
rect 37104 30829 37116 30935
rect 37128 30829 37140 30935
rect 37152 30829 37164 30935
rect 37176 30829 37188 30935
rect 37200 30829 37212 30935
rect 37224 30901 37236 30935
rect 36912 29653 36924 29759
rect 36936 29653 36948 29759
rect 36960 29653 36972 29759
rect 36984 29653 36996 29759
rect 37008 29653 37020 29759
rect 37032 29653 37044 29759
rect 37056 29653 37068 29759
rect 37080 29653 37092 29759
rect 37104 29653 37116 29759
rect 37128 29653 37140 29759
rect 37152 29653 37164 29759
rect 37176 29653 37188 29759
rect 37200 29653 37212 29759
rect 36912 28477 36924 28583
rect 36936 28477 36948 28583
rect 36960 28477 36972 28583
rect 36984 28477 36996 28583
rect 37008 28477 37020 28583
rect 37032 28477 37044 28583
rect 37056 28477 37068 28583
rect 37080 28477 37092 28583
rect 37104 28477 37116 28583
rect 37128 28477 37140 28583
rect 37152 28477 37164 28583
rect 37176 28477 37188 28583
rect 37200 28477 37212 28583
rect 36912 27301 36924 27407
rect 36936 27301 36948 27407
rect 36960 27301 36972 27407
rect 36984 27301 36996 27407
rect 37008 27301 37020 27407
rect 37032 27301 37044 27407
rect 37056 27301 37068 27407
rect 37080 27301 37092 27407
rect 37104 27301 37116 27407
rect 37128 27301 37140 27407
rect 37152 27301 37164 27407
rect 37176 27301 37188 27407
rect 37200 27301 37212 27407
rect 41509 26304 41538 26316
rect 6504 26269 6516 26303
rect 6528 26269 6540 26303
rect 36912 26125 36924 26231
rect 36960 26221 36972 26255
rect 36984 26221 36996 26255
rect 37008 26221 37020 26255
rect 37032 26221 37044 26255
rect 37056 26221 37068 26255
rect 37080 26221 37092 26255
rect 37104 26221 37116 26255
rect 37128 26221 37140 26255
rect 36936 26125 36948 26159
rect 36960 26125 36972 26159
rect 36984 26125 36996 26159
rect 37008 26125 37020 26159
rect 37032 26125 37044 26159
rect 37056 26125 37068 26159
rect 37080 26125 37092 26159
rect 37104 26125 37116 26159
rect 37152 26149 37164 26255
rect 37176 26149 37188 26255
rect 37200 26149 37212 26183
rect 36912 24949 36924 25055
rect 36936 25021 36948 25055
rect 36960 24973 36972 25055
rect 36984 24973 36996 25007
rect 37008 24973 37020 25079
rect 37032 24973 37044 25079
rect 37056 24973 37068 25079
rect 37080 24973 37092 25079
rect 37104 24973 37116 25079
rect 37128 24973 37140 25079
rect 37152 24973 37164 25079
rect 37176 24973 37188 25079
rect 37200 24973 37212 25079
rect 37224 24973 37236 25079
rect 37248 24973 37260 25007
rect 36912 23773 36924 23879
rect 36936 23773 36948 23879
rect 36984 23869 36996 23903
rect 37008 23869 37020 23903
rect 36960 23773 36972 23807
rect 36984 23773 36996 23807
rect 37032 23797 37044 23903
rect 37056 23797 37068 23903
rect 37080 23797 37092 23903
rect 37104 23797 37116 23903
rect 37128 23797 37140 23903
rect 37152 23797 37164 23903
rect 37176 23797 37188 23903
rect 37200 23797 37212 23903
rect 37224 23797 37236 23903
rect 37248 23797 37260 23903
rect 37272 23797 37284 23903
rect 37296 23797 37308 23831
rect 36912 22597 36924 22703
rect 36936 22597 36948 22703
rect 36960 22597 36972 22703
rect 36984 22597 36996 22703
rect 37008 22597 37020 22703
rect 37032 22597 37044 22703
rect 37080 22693 37092 22727
rect 37056 22597 37068 22631
rect 37104 22621 37116 22727
rect 37128 22621 37140 22727
rect 37152 22621 37164 22727
rect 37176 22621 37188 22727
rect 37200 22621 37212 22727
rect 37224 22621 37236 22727
rect 37248 22621 37260 22727
rect 37272 22621 37284 22727
rect 37296 22621 37308 22727
rect 37320 22621 37332 22727
rect 37344 22621 37356 22655
rect 6504 21637 6516 21671
rect 6528 21637 6540 21671
rect 6552 21637 6564 21671
rect 6576 21637 6588 21671
rect 36912 21493 36924 21527
rect 36936 21445 36948 21527
rect 36960 21445 36972 21527
rect 36984 21445 36996 21527
rect 37008 21445 37020 21527
rect 37032 21445 37044 21527
rect 37056 21445 37068 21527
rect 37080 21445 37092 21527
rect 37104 21445 37116 21479
rect 37128 21445 37140 21551
rect 37152 21445 37164 21551
rect 37176 21445 37188 21551
rect 37200 21445 37212 21551
rect 37224 21445 37236 21551
rect 37248 21445 37260 21551
rect 37272 21445 37284 21551
rect 37296 21445 37308 21551
rect 37320 21445 37332 21551
rect 37344 21445 37356 21551
rect 37368 21445 37380 21551
rect 37392 21445 37404 21479
rect 36912 20245 36924 20351
rect 36936 20245 36948 20351
rect 36960 20245 36972 20351
rect 36984 20245 36996 20351
rect 37008 20245 37020 20351
rect 37032 20245 37044 20351
rect 37056 20245 37068 20351
rect 37080 20245 37092 20351
rect 37104 20245 37116 20351
rect 37128 20245 37140 20351
rect 37152 20245 37164 20351
rect 37176 20317 37188 20351
rect 37200 20269 37212 20351
rect 37224 20269 37236 20351
rect 37248 20269 37260 20351
rect 37272 20269 37284 20303
rect 37296 20269 37308 20375
rect 37320 20269 37332 20375
rect 37344 20269 37356 20375
rect 37368 20269 37380 20375
rect 37392 20269 37404 20375
rect 37416 20269 37428 20375
rect 37440 20269 37452 20303
rect 36912 19069 36924 19175
rect 36936 19069 36948 19175
rect 36960 19069 36972 19175
rect 36984 19069 36996 19175
rect 37008 19069 37020 19175
rect 37032 19141 37044 19175
rect 37056 19093 37068 19127
rect 37080 19093 37092 19199
rect 37104 19093 37116 19199
rect 37128 19093 37140 19199
rect 37152 19093 37164 19199
rect 37176 19093 37188 19199
rect 37200 19093 37212 19199
rect 37224 19093 37236 19199
rect 37248 19093 37260 19199
rect 37272 19093 37284 19199
rect 37296 19093 37308 19199
rect 37320 19093 37332 19199
rect 37344 19093 37356 19199
rect 37368 19093 37380 19199
rect 37392 19093 37404 19199
rect 37416 19093 37428 19199
rect 37440 19093 37452 19199
rect 37464 19093 37476 19199
rect 37488 19093 37500 19127
rect 36936 17989 36948 18023
rect 36960 17989 36972 18023
rect 36984 17989 36996 18023
rect 37008 17989 37020 18023
rect 37032 17989 37044 18023
rect 37056 17989 37068 18023
rect 37080 17989 37092 18023
rect 37104 17989 37116 18023
rect 37128 17989 37140 18023
rect 37152 17989 37164 18023
rect 37176 17989 37188 18023
rect 37200 17989 37212 18023
rect 37224 17989 37236 18023
rect 37248 17989 37260 18023
rect 37272 17989 37284 18023
rect 37296 17989 37308 18023
rect 37320 17989 37332 18023
rect 37344 17989 37356 18023
rect 37368 17989 37380 18023
rect 37392 17989 37404 18023
rect 37416 17989 37428 18023
rect 37440 17989 37452 18023
rect 36912 17893 36924 17927
rect 36936 17893 36948 17927
rect 36960 17893 36972 17927
rect 36984 17893 36996 17927
rect 37008 17893 37020 17927
rect 37032 17893 37044 17927
rect 37056 17893 37068 17927
rect 37080 17893 37092 17927
rect 37104 17893 37116 17927
rect 37128 17893 37140 17927
rect 37152 17893 37164 17927
rect 37176 17893 37188 17927
rect 37200 17893 37212 17927
rect 37224 17893 37236 17927
rect 37248 17893 37260 17927
rect 37272 17893 37284 17927
rect 37296 17893 37308 17927
rect 37320 17893 37332 17927
rect 37344 17893 37356 17927
rect 37368 17893 37380 17927
rect 37392 17893 37404 17927
rect 37416 17893 37428 17927
rect 37464 17917 37476 18023
rect 37488 17917 37500 18023
rect 37512 17917 37524 18023
rect 37536 17917 37548 17951
rect 6504 16909 6516 16943
rect 6528 16909 6540 16943
rect 6552 16909 6564 16943
rect 6600 16933 6612 16967
rect 41472 16909 41484 16943
rect 36912 16717 36924 16823
rect 36936 16717 36948 16823
rect 36960 16717 36972 16823
rect 36984 16717 36996 16823
rect 37008 16717 37020 16823
rect 37032 16789 37044 16823
rect 37056 16741 37068 16823
rect 37080 16741 37092 16823
rect 37104 16741 37116 16823
rect 37128 16741 37140 16775
rect 37152 16741 37164 16847
rect 37176 16741 37188 16847
rect 37200 16741 37212 16847
rect 37224 16741 37236 16847
rect 37248 16741 37260 16847
rect 37272 16741 37284 16847
rect 37296 16741 37308 16847
rect 37320 16741 37332 16847
rect 37344 16741 37356 16847
rect 37368 16741 37380 16847
rect 37392 16741 37404 16847
rect 37416 16741 37428 16847
rect 37440 16741 37452 16847
rect 37464 16741 37476 16847
rect 37488 16741 37500 16847
rect 37512 16741 37524 16847
rect 37536 16741 37548 16847
rect 41472 16765 41484 16799
rect 7536 16525 7548 16607
rect 11328 16525 11340 16607
rect 11352 16525 11364 16607
rect 11376 16525 11388 16607
rect 11400 16525 11412 16607
rect 11424 16525 11436 16559
rect 11451 16525 11463 16650
rect 11474 16498 11486 16650
rect 11497 16525 11509 16650
rect 11520 16498 11532 16650
rect 11543 16525 11555 16650
rect 11566 16498 11578 16650
rect 11589 16525 11601 16650
rect 11612 16498 11624 16650
rect 11904 16621 11916 16650
rect 11640 16525 11652 16559
rect 11928 16501 11940 16583
rect 12036 16573 12048 16650
rect 12060 16573 12072 16650
rect 12084 16573 12096 16650
rect 12108 16621 12120 16650
rect 13380 16621 13392 16650
rect 13572 16621 13584 16650
rect 14364 16621 14376 16650
rect 14916 16621 14928 16650
rect 15132 16621 15144 16650
rect 15876 16621 15888 16650
rect 16044 16621 16056 16650
rect 16428 16621 16440 16650
rect 16620 16621 16632 16650
rect 16836 16621 16848 16650
rect 17580 16621 17592 16650
rect 17748 16621 17760 16650
rect 27156 16621 27168 16650
rect 27348 16621 27360 16650
rect 27588 16621 27600 16650
rect 35292 16621 35304 16650
rect 13381 16607 13392 16621
rect 13573 16607 13584 16621
rect 14365 16607 14376 16621
rect 14917 16607 14928 16621
rect 15133 16607 15144 16621
rect 15877 16607 15888 16621
rect 16045 16607 16056 16621
rect 16429 16607 16440 16621
rect 16621 16607 16632 16621
rect 16837 16607 16848 16621
rect 17581 16607 17592 16621
rect 17749 16607 17760 16621
rect 27157 16607 27168 16621
rect 27349 16607 27360 16621
rect 27589 16607 27600 16621
rect 35293 16607 35304 16621
rect 36036 16620 36048 16650
rect 36180 16620 36192 16650
rect 36228 16620 36240 16650
rect 36276 16620 36288 16650
rect 36324 16620 36336 16650
rect 36396 16620 36408 16650
rect 36024 16608 36048 16620
rect 36168 16608 36192 16620
rect 36216 16608 36240 16620
rect 36264 16608 36288 16620
rect 36312 16608 36336 16620
rect 36384 16608 36408 16620
rect 35306 16525 35318 16583
rect 36024 16573 36036 16608
rect 36168 16549 36180 16608
rect 36216 16525 36228 16608
rect 36264 16597 36276 16608
rect 36240 16525 36252 16583
rect 36264 16525 36276 16583
rect 36288 16549 36300 16583
rect 36312 16573 36324 16608
rect 36384 16573 36396 16608
rect 36720 16525 36732 16650
rect 36912 16477 36924 16607
rect 36936 16477 36948 16607
rect 36960 16477 36972 16607
rect 36984 16477 36996 16607
rect 37008 16477 37020 16559
rect 37032 16477 37044 16631
rect 37056 16477 37068 16631
rect 37080 16477 37092 16631
rect 37104 16477 37116 16631
rect 37128 16477 37140 16631
rect 37152 16477 37164 16631
rect 37176 16477 37188 16631
rect 37200 16477 37212 16631
rect 37224 16477 37236 16631
rect 37248 16477 37260 16631
rect 37272 16477 37284 16631
rect 37296 16477 37308 16631
rect 37320 16477 37332 16631
rect 37344 16477 37356 16631
rect 37368 16477 37380 16631
rect 37392 16477 37404 16631
rect 37416 16477 37428 16631
rect 37440 16477 37452 16631
rect 37464 16477 37476 16631
rect 37488 16477 37500 16631
rect 37512 16477 37524 16631
rect 37536 16477 37548 16631
rect 37560 16477 37572 16631
rect 37584 16477 37596 16559
rect 7464 15829 7476 15863
rect 7536 15829 7548 15911
rect 11136 15829 11148 15911
rect 11184 15829 11196 15935
rect 11232 15829 11244 15959
rect 11256 15829 11268 15983
rect 11280 15949 11292 16007
rect 11304 15853 11316 15935
rect 11400 15925 11412 15959
rect 11424 15925 11436 15959
rect 11640 15877 11652 16151
rect 11664 15877 11676 16127
rect 11592 15793 11604 15863
rect 11726 15793 11738 15911
rect 11750 15901 11762 16127
rect 11750 15793 11762 15887
rect 11774 15853 11786 16127
rect 11774 15793 11786 15839
rect 11798 15793 11810 16127
rect 11832 15853 11844 16103
rect 11856 15925 11868 16079
rect 11880 15925 11892 16055
rect 13848 15877 13860 16079
rect 13824 15828 13836 15863
rect 14712 15853 14724 16079
rect 15576 15901 15588 16103
rect 16416 15925 16428 16151
rect 16992 16045 17004 16175
rect 13814 15816 13836 15828
rect 13814 15793 13826 15816
rect 14678 15815 14687 15829
rect 15552 15828 15564 15887
rect 15542 15816 15564 15828
rect 16392 15828 16404 15911
rect 16968 15828 16980 16031
rect 18168 16021 18180 16199
rect 18144 15828 18156 16007
rect 18192 15997 18204 16175
rect 16392 15816 16406 15828
rect 16968 15816 16982 15828
rect 14678 15793 14690 15815
rect 15542 15793 15554 15816
rect 16394 15793 16406 15816
rect 16970 15793 16982 15816
rect 18134 15816 18156 15828
rect 18168 15828 18180 15983
rect 19896 15973 19908 16151
rect 20760 16069 20772 16127
rect 19872 15828 19884 15959
rect 20736 15828 20748 16055
rect 21192 15877 21204 16103
rect 18168 15816 18182 15828
rect 18134 15793 18146 15816
rect 18170 15793 18182 15816
rect 19862 15816 19884 15828
rect 20726 15816 20748 15828
rect 21168 15828 21180 15863
rect 22128 15853 22140 16079
rect 22896 15853 22908 16055
rect 23928 15901 23940 16031
rect 21168 15816 21182 15828
rect 19862 15793 19874 15816
rect 20726 15793 20738 15816
rect 21170 15793 21182 15816
rect 22117 15815 22118 15829
rect 22885 15815 22886 15829
rect 23904 15828 23916 15887
rect 24240 15877 24252 16007
rect 24216 15828 24228 15863
rect 25824 15853 25836 15983
rect 23904 15816 23918 15828
rect 24216 15816 24230 15828
rect 22106 15793 22118 15815
rect 22874 15793 22886 15815
rect 23906 15793 23918 15816
rect 24218 15793 24230 15816
rect 25813 15815 25814 15829
rect 26760 15828 26772 15911
rect 26784 15828 26796 15959
rect 27144 15925 27156 15959
rect 27672 15901 27684 15983
rect 27648 15828 27660 15887
rect 28512 15877 28524 15959
rect 32760 15925 32772 15959
rect 33600 15925 33612 15959
rect 26760 15816 26774 15828
rect 26784 15816 26798 15828
rect 25802 15793 25814 15815
rect 26762 15793 26774 15816
rect 26786 15793 26798 15816
rect 27638 15816 27660 15828
rect 28488 15828 28500 15863
rect 28488 15816 28502 15828
rect 27638 15793 27650 15816
rect 28490 15793 28502 15816
rect 30170 15793 30182 15815
rect 30194 15793 30206 15911
rect 30219 15853 30231 15887
rect 31608 15828 31620 15863
rect 31608 15816 31622 15828
rect 31610 15793 31622 15816
rect 31909 15815 31910 15829
rect 31898 15793 31910 15815
rect 32750 15815 32759 15829
rect 33613 15815 33614 15829
rect 32750 15793 32762 15815
rect 33602 15793 33614 15815
rect 35282 15793 35294 15959
rect 35306 15793 35318 15959
rect 36168 15925 36180 15959
rect 36912 15925 36924 15959
rect 36936 15925 36948 15959
rect 36960 15925 36972 15959
rect 36984 15925 36996 15959
rect 36158 15815 36167 15829
rect 37008 15828 37020 15959
rect 38592 15828 38604 16511
rect 37008 15816 37022 15828
rect 38592 15816 38606 15828
rect 36158 15793 36170 15815
rect 37010 15793 37022 15816
rect 38594 15793 38606 15816
rect 38856 15793 38868 16487
rect 39168 15829 39180 16463
rect 39192 15829 39204 16439
rect 39216 15829 39228 16415
rect 39240 15829 39252 16391
rect 39264 15829 39276 16367
rect 39288 15829 39300 16343
rect 39312 15829 39324 16319
rect 39336 15829 39348 16295
rect 39360 15829 39372 16271
rect 39384 15829 39396 16247
rect 39408 15829 39420 16223
rect 39432 15829 39444 16199
rect 39456 15829 39468 16175
rect 39480 15829 39492 16151
rect 39504 15829 39516 16127
rect 39528 15829 39540 16103
rect 39552 15829 39564 16079
rect 39576 15829 39588 16055
rect 39648 15829 39660 16031
rect 39672 15829 39684 16007
rect 39696 15829 39708 15983
rect 39744 15829 39756 15959
rect 39792 15829 39804 15935
rect 41376 15829 41388 15911
rect 41424 15829 41436 15887
rect 41448 15829 41460 15863
rect 11184 15663 11196 15695
rect 11232 15637 11244 15695
rect 11256 15637 11268 15695
rect 11280 15637 11292 15695
rect 11304 15637 11316 15695
rect 11328 15637 11340 15695
rect 11365 15674 11387 15686
rect 11365 15650 11387 15662
rect 39122 15578 39143 15590
rect 39122 15554 39143 15566
rect 39122 15530 39143 15542
rect 39122 15506 39143 15518
rect 39122 15482 39143 15494
rect 39168 15471 39180 15601
rect 39192 15471 39204 15601
rect 39216 15471 39228 15601
rect 39240 15471 39252 15601
rect 39264 15471 39276 15601
rect 39312 15471 39324 15577
rect 39336 15471 39348 15577
rect 39360 15471 39372 15577
rect 39384 15495 39396 15577
rect 39432 15519 39444 15553
rect 39456 15519 39468 15553
rect 39480 15519 39492 15553
rect 39504 15519 39516 15553
rect 39528 15519 39540 15553
rect 39552 15519 39564 15553
rect 39576 15519 39588 15553
rect 39600 15519 39612 15553
rect 39624 15519 39636 15553
rect 6504 12181 6516 12215
rect 7464 12181 7476 12215
rect 7536 12181 7548 12215
rect 11232 12181 11244 12215
rect 11256 12181 11268 12215
rect 11280 12181 11292 12215
rect 11304 12181 11316 12215
rect 41424 12181 41436 12215
rect 41448 12181 41460 12215
rect 11232 11557 11244 11598
rect 11256 11557 11268 11598
rect 11280 11566 11292 11598
rect 11304 11533 11316 11598
rect 11365 11577 11387 11589
rect 11365 11553 11387 11565
rect 39122 10477 39157 10485
rect 39122 10473 39143 10477
rect 39168 10453 39180 10487
rect 39192 10453 39204 10487
rect 39216 10453 39228 10487
rect 39240 10453 39252 10487
rect 39264 10453 39276 10487
rect 39312 10453 39324 10487
rect 39336 10453 39348 10487
rect 39360 10453 39372 10487
rect 39456 10453 39468 10487
rect 39480 10453 39492 10487
rect 39504 10453 39516 10487
rect 39528 10453 39540 10487
rect 39122 9225 39143 9237
rect 39122 9201 39143 9213
rect 39122 9177 39143 9189
rect 39168 9157 39180 9247
rect 39192 9157 39204 9247
rect 39216 9157 39228 9247
rect 39240 9157 39252 9247
rect 39264 9157 39276 9247
rect 39312 9157 39324 9247
rect 39336 9189 39348 9247
rect 39122 8015 39143 8020
rect 39122 8008 39157 8015
rect 39168 8005 39180 8039
rect 39192 8005 39204 8039
rect 39216 8005 39228 8039
rect 39240 8005 39252 8039
rect 39264 8005 39276 8039
rect 39312 8005 39324 8039
rect 39480 8005 39492 8039
rect 39504 8005 39516 8039
rect 7464 7645 7476 7679
rect 11232 7645 11244 7679
rect 11256 7645 11268 7679
rect 11304 7645 11316 7679
rect 11365 7655 11387 7660
rect 11351 7648 11387 7655
rect 39122 7648 39143 7660
rect 11328 7624 11387 7636
rect 39122 7624 39143 7636
rect 7464 7453 7476 7487
rect 11232 7477 11244 7511
rect 11256 7453 11268 7511
rect 11304 7453 11316 7559
rect 11328 7453 11340 7624
rect 39122 7600 39143 7612
rect 11726 7572 11738 7589
rect 11798 7573 11810 7589
rect 11726 7560 11748 7572
rect 11736 7525 11748 7560
rect 11798 7559 11807 7573
rect 19370 7572 19382 7589
rect 22562 7572 22574 7589
rect 19368 7560 19382 7572
rect 22560 7560 22574 7572
rect 25814 7572 25826 7589
rect 35306 7572 35318 7589
rect 25814 7560 25836 7572
rect 19368 7549 19380 7560
rect 22560 7549 22572 7560
rect 19368 7501 19380 7535
rect 15816 7405 15828 7439
rect 19800 7405 19812 7463
rect 19944 7405 19956 7463
rect 22560 7405 22572 7535
rect 25824 7525 25836 7560
rect 35304 7560 35318 7572
rect 35304 7525 35316 7560
rect 25824 7357 25836 7463
rect 28200 7309 28212 7463
rect 32184 7309 32196 7463
rect 36456 7405 36468 7511
rect 36480 7357 36492 7463
rect 36504 7405 36516 7487
rect 39168 7405 39180 7679
rect 39192 7582 39204 7679
rect 39216 7582 39228 7679
rect 39240 7637 39252 7679
rect 39264 7477 39276 7679
rect 39312 7429 39324 7679
rect 39480 7501 39492 7679
rect 36456 7309 36468 7343
rect 39192 7333 39204 7391
rect 39576 7309 39588 7631
rect 39600 7429 39612 7631
rect 39672 7501 39684 7535
rect 39696 7501 39708 7535
rect 39744 7501 39756 7535
rect 39792 7501 39804 7535
rect 41424 7501 41436 7535
rect 41472 7453 41484 7487
rect 39696 7309 39708 7367
rect 39744 7309 39756 7367
rect 41472 7309 41484 7343
rect 7464 6517 7476 6551
rect 11304 6517 11316 6575
rect 11328 6541 11340 6575
rect 11688 6493 11700 6527
rect 15672 6493 15684 6527
rect 15816 6493 15828 6527
rect 19800 6493 19812 6527
rect 19944 6493 19956 6527
rect 28056 6493 28068 6527
rect 28200 6493 28212 6551
rect 32184 6493 32196 6551
rect 32328 6493 32340 6551
rect 36312 6493 36324 6575
rect 36456 6493 36468 6599
rect 36504 6517 36516 6599
rect 36552 6541 36564 6575
rect 39576 6517 39588 6623
rect 39696 6589 39708 6623
rect 39744 6589 39756 6623
<< metal4 >>
rect 6702 46264 8262 47824
rect 10830 46264 12390 47824
rect 14958 46264 16518 47824
rect 19086 46264 20646 47824
rect 23214 46264 24774 47824
rect 27342 46264 28902 47824
rect 31470 46264 33030 47824
rect 35598 46264 37158 47824
rect 39726 46264 41286 47824
rect 78 39726 1638 41286
rect 46350 39726 47910 41286
rect 78 34996 1638 36556
rect 46350 34996 47910 36556
rect 78 30266 1638 31826
rect 46350 30266 47910 31826
rect 78 25536 1638 27096
rect 46350 25536 47910 27096
rect 78 20806 1638 22366
rect 46350 20806 47910 22366
rect 78 16076 1638 17636
rect 46350 16076 47910 17636
rect 78 11346 1638 12906
rect 46350 11346 47910 12906
rect 78 6616 1638 8176
rect 46350 6616 47910 8176
rect 6702 78 8262 1638
rect 10830 78 12390 1638
rect 14958 78 16518 1638
rect 19086 78 20646 1638
rect 23214 78 24774 1638
rect 27342 78 28902 1638
rect 31470 78 33030 1638
rect 35598 78 37158 1638
rect 39726 78 41286 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 0 -1 0 47902
box 0 0 6450 6450
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform 0 -1 6536 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform 0 -1 6622 1 0 41452
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 8342 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform 0 -1 8428 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform 0 -1 8514 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform 0 -1 8600 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform 0 -1 8686 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform 0 -1 8772 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform 0 -1 8858 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform 0 -1 8944 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform 0 -1 9030 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform 0 -1 9116 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform 0 -1 9202 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform 0 -1 9288 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform 0 -1 9374 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform 0 -1 9460 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform 0 -1 9546 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform 0 -1 9632 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform 0 -1 9718 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform 0 -1 9804 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform 0 -1 9890 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform 0 -1 9976 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform 0 -1 10062 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform 0 -1 10148 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform 0 -1 10234 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform 0 -1 10320 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform 0 -1 10406 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform 0 -1 10492 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform 0 -1 10578 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform 0 -1 10664 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform 0 -1 10750 1 0 41452
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 12470 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform 0 -1 12556 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform 0 -1 12642 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform 0 -1 12728 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform 0 -1 12814 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform 0 -1 12900 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform 0 -1 12986 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform 0 -1 13072 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform 0 -1 13158 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform 0 -1 13244 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform 0 -1 13330 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform 0 -1 13416 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform 0 -1 13502 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform 0 -1 13588 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform 0 -1 13674 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform 0 -1 13760 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform 0 -1 13846 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform 0 -1 13932 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform 0 -1 14018 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform 0 -1 14104 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform 0 -1 14190 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform 0 -1 14276 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform 0 -1 14362 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform 0 -1 14448 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform 0 -1 14534 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform 0 -1 14620 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform 0 -1 14706 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform 0 -1 14792 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform 0 -1 14878 1 0 41452
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 16598 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform 0 -1 16684 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform 0 -1 16770 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform 0 -1 16856 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform 0 -1 16942 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform 0 -1 17028 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform 0 -1 17114 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform 0 -1 17200 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform 0 -1 17286 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform 0 -1 17372 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform 0 -1 17458 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform 0 -1 17544 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform 0 -1 17630 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform 0 -1 17716 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform 0 -1 17802 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform 0 -1 17888 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform 0 -1 17974 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform 0 -1 18060 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform 0 -1 18146 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform 0 -1 18232 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform 0 -1 18318 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform 0 -1 18404 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform 0 -1 18490 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform 0 -1 18576 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform 0 -1 18662 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform 0 -1 18748 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform 0 -1 18834 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform 0 -1 18920 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform 0 -1 19006 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 20726 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform 0 -1 20812 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform 0 -1 20898 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform 0 -1 20984 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform 0 -1 21070 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform 0 -1 21156 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform 0 -1 21242 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform 0 -1 21328 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform 0 -1 21414 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform 0 -1 21500 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform 0 -1 21586 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform 0 -1 21672 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform 0 -1 21758 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform 0 -1 21844 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform 0 -1 21930 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform 0 -1 22016 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform 0 -1 22102 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform 0 -1 22188 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform 0 -1 22274 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform 0 -1 22360 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform 0 -1 22446 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform 0 -1 22532 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform 0 -1 22618 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform 0 -1 22704 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform 0 -1 22790 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform 0 -1 22876 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform 0 -1 22962 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform 0 -1 23048 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform 0 -1 23134 1 0 41452
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 24854 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform 0 -1 24940 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform 0 -1 25026 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform 0 -1 25112 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform 0 -1 25198 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform 0 -1 25284 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform 0 -1 25370 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform 0 -1 25456 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform 0 -1 25542 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform 0 -1 25628 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform 0 -1 25714 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform 0 -1 25800 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform 0 -1 25886 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform 0 -1 25972 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform 0 -1 26058 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform 0 -1 26144 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform 0 -1 26230 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform 0 -1 26316 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform 0 -1 26402 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform 0 -1 26488 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform 0 -1 26574 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform 0 -1 26660 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform 0 -1 26746 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform 0 -1 26832 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform 0 -1 26918 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform 0 -1 27004 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 27090 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 27176 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 27262 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 28982 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 29068 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 29154 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 29240 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 29326 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 29412 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 29498 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 29584 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 29670 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 29756 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 29842 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 29928 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 30014 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 30100 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 30186 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 30272 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 30358 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 30444 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 0 -1 30530 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 0 -1 30616 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 0 -1 30702 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 0 -1 30788 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 0 -1 30874 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 0 -1 30960 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 0 -1 31046 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 0 -1 31132 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 0 -1 31218 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 0 -1 31304 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 0 -1 31390 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 33110 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 0 -1 33196 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 0 -1 33282 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 0 -1 33368 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 0 -1 33454 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 33540 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 33626 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 33712 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 33798 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 33884 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 33970 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 34056 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 34142 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 34228 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 34314 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 34400 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 34486 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 34572 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 34658 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 34744 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 34830 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 34916 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 35002 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 35088 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 35174 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 35260 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 35346 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 35432 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 35518 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 37238 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 37324 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 37410 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 37496 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 37582 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 37668 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 37754 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 37840 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 37926 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 38012 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 38098 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 38184 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 38270 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 38356 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 38442 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 38528 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 38614 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 38700 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 38786 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 38872 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 38958 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 39044 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 39130 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 39216 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 39302 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 39388 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 39474 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 39560 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 39646 1 0 41452
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 41366 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 41452 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 41538 1 0 41452
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 47988 0 -1 47902
box 0 0 6450 6450
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 6450 0 -1 41452
box 0 0 6450 86
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 6450 0 -1 41366
box 0 0 6450 1720
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 6450 0 -1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 6450 0 -1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 6450 0 -1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 6450 0 -1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 6450 0 -1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 6450 0 -1 39216
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 6450 0 -1 39130
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 6450 0 -1 39044
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 6450 0 -1 38958
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 6450 0 -1 38872
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 6450 0 -1 38786
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 6450 0 -1 38700
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 6450 0 -1 38614
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 6450 0 -1 38528
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform -1 0 6450 0 -1 38442
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform -1 0 6450 0 -1 38356
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform -1 0 6450 0 -1 38270
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform -1 0 6450 0 -1 38184
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform -1 0 6450 0 -1 38098
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform -1 0 6450 0 -1 38012
box 0 0 6450 86
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform -1 0 6450 0 -1 37926
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform -1 0 6450 0 -1 37840
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform -1 0 6450 0 -1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform -1 0 6450 0 -1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform -1 0 6450 0 -1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform -1 0 6450 0 -1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform -1 0 6450 0 -1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform -1 0 6450 0 -1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform -1 0 6450 0 -1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 1 0 41538 0 1 41366
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 41538 0 1 39646
box 0 0 6450 1720
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 1 0 41538 0 1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 1 0 41538 0 1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 1 0 41538 0 1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 1 0 41538 0 1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 1 0 41538 0 1 39216
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 1 0 41538 0 1 39130
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 1 0 41538 0 1 39044
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 1 0 41538 0 1 38958
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 1 0 41538 0 1 38872
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 1 0 41538 0 1 38786
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 1 0 41538 0 1 38700
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 1 0 41538 0 1 38614
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 1 0 41538 0 1 38528
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 1 0 41538 0 1 38442
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 1 0 41538 0 1 38356
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 1 0 41538 0 1 38270
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 1 0 41538 0 1 38184
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 1 0 41538 0 1 38098
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 1 0 41538 0 1 38012
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 1 0 41538 0 1 37926
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 1 0 41538 0 1 37840
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 1 0 41538 0 1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 1 0 41538 0 1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 1 0 41538 0 1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 1 0 41538 0 1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 1 0 41538 0 1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 1 0 41538 0 1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 1 0 41538 0 1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform -1 0 6450 0 -1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform -1 0 6450 0 -1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform -1 0 6450 0 -1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform -1 0 6450 0 -1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform -1 0 6450 0 -1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform -1 0 6450 0 -1 36722
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 6450 0 -1 36636
box 0 0 6450 1720
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform -1 0 6450 0 -1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform -1 0 6450 0 -1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform -1 0 6450 0 -1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform -1 0 6450 0 -1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform -1 0 6450 0 -1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform -1 0 6450 0 -1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform -1 0 6450 0 -1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform -1 0 6450 0 -1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform -1 0 6450 0 -1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform -1 0 6450 0 -1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform -1 0 6450 0 -1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform -1 0 6450 0 -1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform -1 0 6450 0 -1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform -1 0 6450 0 -1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform -1 0 6450 0 -1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform -1 0 6450 0 -1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform -1 0 6450 0 -1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform -1 0 6450 0 -1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform -1 0 6450 0 -1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform -1 0 6450 0 -1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform -1 0 6450 0 -1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform -1 0 6450 0 -1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform -1 0 6450 0 -1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform -1 0 6450 0 -1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform -1 0 6450 0 -1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform -1 0 6450 0 -1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform -1 0 6450 0 -1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform -1 0 6450 0 -1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform -1 0 6450 0 -1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform -1 0 6450 0 -1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform -1 0 6450 0 -1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform -1 0 6450 0 -1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform -1 0 6450 0 -1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform -1 0 6450 0 -1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform -1 0 6450 0 -1 31992
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 6450 0 -1 31906
box 0 0 6450 1720
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform -1 0 6450 0 -1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform -1 0 6450 0 -1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform -1 0 6450 0 -1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform -1 0 6450 0 -1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform -1 0 6450 0 -1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform -1 0 6450 0 -1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform -1 0 6450 0 -1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform -1 0 6450 0 -1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform -1 0 6450 0 -1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform -1 0 6450 0 -1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform -1 0 6450 0 -1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform -1 0 6450 0 -1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform -1 0 6450 0 -1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform -1 0 6450 0 -1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_788
timestamp 1300117811
transform -1 0 6450 0 -1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_789
timestamp 1300117811
transform -1 0 6450 0 -1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_790
timestamp 1300117811
transform -1 0 6450 0 -1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_791
timestamp 1300117811
transform -1 0 6450 0 -1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_792
timestamp 1300117811
transform -1 0 6450 0 -1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_793
timestamp 1300117811
transform -1 0 6450 0 -1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_794
timestamp 1300117811
transform -1 0 6450 0 -1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_795
timestamp 1300117811
transform -1 0 6450 0 -1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_796
timestamp 1300117811
transform -1 0 6450 0 -1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_797
timestamp 1300117811
transform -1 0 6450 0 -1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_798
timestamp 1300117811
transform -1 0 6450 0 -1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_799
timestamp 1300117811
transform -1 0 6450 0 -1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_800
timestamp 1300117811
transform -1 0 6450 0 -1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_801
timestamp 1300117811
transform -1 0 6450 0 -1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_802
timestamp 1300117811
transform -1 0 6450 0 -1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_803
timestamp 1300117811
transform -1 0 6450 0 -1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_804
timestamp 1300117811
transform -1 0 6450 0 -1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_805
timestamp 1300117811
transform -1 0 6450 0 -1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_806
timestamp 1300117811
transform -1 0 6450 0 -1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_807
timestamp 1300117811
transform -1 0 6450 0 -1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_808
timestamp 1300117811
transform -1 0 6450 0 -1 27262
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 6450 0 -1 27176
box 0 0 6450 1720
use fillpp_mt fillpp_mt_809
timestamp 1300117811
transform -1 0 6450 0 -1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_810
timestamp 1300117811
transform -1 0 6450 0 -1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_811
timestamp 1300117811
transform -1 0 6450 0 -1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_812
timestamp 1300117811
transform -1 0 6450 0 -1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_813
timestamp 1300117811
transform -1 0 6450 0 -1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_814
timestamp 1300117811
transform -1 0 6450 0 -1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_815
timestamp 1300117811
transform -1 0 6450 0 -1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_816
timestamp 1300117811
transform -1 0 6450 0 -1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_817
timestamp 1300117811
transform -1 0 6450 0 -1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_818
timestamp 1300117811
transform -1 0 6450 0 -1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_819
timestamp 1300117811
transform -1 0 6450 0 -1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_820
timestamp 1300117811
transform -1 0 6450 0 -1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_821
timestamp 1300117811
transform -1 0 6450 0 -1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_822
timestamp 1300117811
transform -1 0 6450 0 -1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_823
timestamp 1300117811
transform -1 0 6450 0 -1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_824
timestamp 1300117811
transform -1 0 6450 0 -1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_825
timestamp 1300117811
transform -1 0 6450 0 -1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_826
timestamp 1300117811
transform -1 0 6450 0 -1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_827
timestamp 1300117811
transform -1 0 6450 0 -1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_828
timestamp 1300117811
transform -1 0 6450 0 -1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_829
timestamp 1300117811
transform -1 0 6450 0 -1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_830
timestamp 1300117811
transform -1 0 6450 0 -1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_831
timestamp 1300117811
transform -1 0 6450 0 -1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_832
timestamp 1300117811
transform -1 0 6450 0 -1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_833
timestamp 1300117811
transform -1 0 6450 0 -1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_834
timestamp 1300117811
transform -1 0 6450 0 -1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_835
timestamp 1300117811
transform -1 0 6450 0 -1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_836
timestamp 1300117811
transform -1 0 6450 0 -1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_837
timestamp 1300117811
transform -1 0 6450 0 -1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_838
timestamp 1300117811
transform -1 0 6450 0 -1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_839
timestamp 1300117811
transform -1 0 6450 0 -1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_840
timestamp 1300117811
transform -1 0 6450 0 -1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_841
timestamp 1300117811
transform -1 0 6450 0 -1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_842
timestamp 1300117811
transform -1 0 6450 0 -1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_843
timestamp 1300117811
transform -1 0 6450 0 -1 22532
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 6450 0 -1 22446
box 0 0 6450 1720
use fillpp_mt fillpp_mt_844
timestamp 1300117811
transform -1 0 6450 0 -1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_845
timestamp 1300117811
transform -1 0 6450 0 -1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_846
timestamp 1300117811
transform -1 0 6450 0 -1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_847
timestamp 1300117811
transform -1 0 6450 0 -1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_848
timestamp 1300117811
transform -1 0 6450 0 -1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_849
timestamp 1300117811
transform -1 0 6450 0 -1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_850
timestamp 1300117811
transform -1 0 6450 0 -1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_851
timestamp 1300117811
transform -1 0 6450 0 -1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_852
timestamp 1300117811
transform -1 0 6450 0 -1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_853
timestamp 1300117811
transform -1 0 6450 0 -1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_854
timestamp 1300117811
transform -1 0 6450 0 -1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_855
timestamp 1300117811
transform -1 0 6450 0 -1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_856
timestamp 1300117811
transform -1 0 6450 0 -1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_857
timestamp 1300117811
transform -1 0 6450 0 -1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_858
timestamp 1300117811
transform -1 0 6450 0 -1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_859
timestamp 1300117811
transform -1 0 6450 0 -1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_860
timestamp 1300117811
transform -1 0 6450 0 -1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_861
timestamp 1300117811
transform -1 0 6450 0 -1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_862
timestamp 1300117811
transform -1 0 6450 0 -1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_863
timestamp 1300117811
transform -1 0 6450 0 -1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_864
timestamp 1300117811
transform -1 0 6450 0 -1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_865
timestamp 1300117811
transform -1 0 6450 0 -1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_866
timestamp 1300117811
transform -1 0 6450 0 -1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_867
timestamp 1300117811
transform -1 0 6450 0 -1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_868
timestamp 1300117811
transform -1 0 6450 0 -1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_869
timestamp 1300117811
transform -1 0 6450 0 -1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_870
timestamp 1300117811
transform -1 0 6450 0 -1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_871
timestamp 1300117811
transform -1 0 6450 0 -1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_872
timestamp 1300117811
transform -1 0 6450 0 -1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_873
timestamp 1300117811
transform -1 0 6450 0 -1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_874
timestamp 1300117811
transform -1 0 6450 0 -1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_875
timestamp 1300117811
transform -1 0 6450 0 -1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_876
timestamp 1300117811
transform -1 0 6450 0 -1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_877
timestamp 1300117811
transform -1 0 6450 0 -1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_878
timestamp 1300117811
transform -1 0 6450 0 -1 17802
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 6450 0 -1 17716
box 0 0 6450 1720
use datapath datapath_0
timestamp 1395690245
transform 1 0 11450 0 1 16650
box 0 0 25408 20572
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 1 0 41538 0 1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 1 0 41538 0 1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 1 0 41538 0 1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 1 0 41538 0 1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 1 0 41538 0 1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 1 0 41538 0 1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 1 0 41538 0 1 36636
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 41538 0 1 34916
box 0 0 6450 1720
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 1 0 41538 0 1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 1 0 41538 0 1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 1 0 41538 0 1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 1 0 41538 0 1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 1 0 41538 0 1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 1 0 41538 0 1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 1 0 41538 0 1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 1 0 41538 0 1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 1 0 41538 0 1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 1 0 41538 0 1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 1 0 41538 0 1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 1 0 41538 0 1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 1 0 41538 0 1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 1 0 41538 0 1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 1 0 41538 0 1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 1 0 41538 0 1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 1 0 41538 0 1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 1 0 41538 0 1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 1 0 41538 0 1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 1 0 41538 0 1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 1 0 41538 0 1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 1 0 41538 0 1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 1 0 41538 0 1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 1 0 41538 0 1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 1 0 41538 0 1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 1 0 41538 0 1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 1 0 41538 0 1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 1 0 41538 0 1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 1 0 41538 0 1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 1 0 41538 0 1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 1 0 41538 0 1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 1 0 41538 0 1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 1 0 41538 0 1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 1 0 41538 0 1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 1 0 41538 0 1 31906
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 41538 0 1 30186
box 0 0 6450 1720
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 1 0 41538 0 1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 1 0 41538 0 1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 1 0 41538 0 1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 1 0 41538 0 1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 1 0 41538 0 1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 1 0 41538 0 1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 1 0 41538 0 1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 1 0 41538 0 1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 1 0 41538 0 1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 1 0 41538 0 1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 41538 0 1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 41538 0 1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 41538 0 1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 41538 0 1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 41538 0 1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 41538 0 1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 41538 0 1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 41538 0 1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 41538 0 1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 41538 0 1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 41538 0 1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 41538 0 1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 41538 0 1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 41538 0 1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 41538 0 1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 41538 0 1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 41538 0 1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 41538 0 1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 41538 0 1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 41538 0 1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 41538 0 1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 41538 0 1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 41538 0 1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 41538 0 1 27262
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 41538 0 1 27176
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 41538 0 1 25456
box 0 0 6450 1720
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 41538 0 1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 41538 0 1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 41538 0 1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 41538 0 1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 41538 0 1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 41538 0 1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 41538 0 1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 41538 0 1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 41538 0 1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 41538 0 1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 41538 0 1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 41538 0 1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 41538 0 1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 41538 0 1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 41538 0 1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 41538 0 1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 41538 0 1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 41538 0 1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 41538 0 1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 41538 0 1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 41538 0 1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 41538 0 1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 41538 0 1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 41538 0 1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 41538 0 1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 41538 0 1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 41538 0 1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 41538 0 1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 41538 0 1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 41538 0 1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 41538 0 1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 41538 0 1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 41538 0 1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 41538 0 1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 41538 0 1 22446
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 41538 0 1 20726
box 0 0 6450 1720
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 41538 0 1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 41538 0 1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 41538 0 1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 41538 0 1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 41538 0 1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 41538 0 1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 41538 0 1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 41538 0 1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 41538 0 1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 41538 0 1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 41538 0 1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 41538 0 1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 41538 0 1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 41538 0 1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 41538 0 1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 41538 0 1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 41538 0 1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 41538 0 1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 41538 0 1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 41538 0 1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 41538 0 1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 41538 0 1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 41538 0 1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 41538 0 1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 41538 0 1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 41538 0 1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 41538 0 1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 41538 0 1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 41538 0 1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 41538 0 1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 41538 0 1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 41538 0 1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 41538 0 1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 41538 0 1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 41538 0 1 17716
box 0 0 6450 86
use fillpp_mt fillpp_mt_879
timestamp 1300117811
transform -1 0 6450 0 -1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_880
timestamp 1300117811
transform -1 0 6450 0 -1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_881
timestamp 1300117811
transform -1 0 6450 0 -1 15824
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 41538 0 1 15996
box 0 0 6450 1720
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 41538 0 1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 41538 0 1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_882
timestamp 1300117811
transform -1 0 6450 0 -1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_883
timestamp 1300117811
transform -1 0 6450 0 -1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_884
timestamp 1300117811
transform -1 0 6450 0 -1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_885
timestamp 1300117811
transform -1 0 6450 0 -1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_886
timestamp 1300117811
transform -1 0 6450 0 -1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_887
timestamp 1300117811
transform -1 0 6450 0 -1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_888
timestamp 1300117811
transform -1 0 6450 0 -1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_889
timestamp 1300117811
transform -1 0 6450 0 -1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_890
timestamp 1300117811
transform -1 0 6450 0 -1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_891
timestamp 1300117811
transform -1 0 6450 0 -1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_892
timestamp 1300117811
transform -1 0 6450 0 -1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_893
timestamp 1300117811
transform -1 0 6450 0 -1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_894
timestamp 1300117811
transform -1 0 6450 0 -1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_895
timestamp 1300117811
transform -1 0 6450 0 -1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_896
timestamp 1300117811
transform -1 0 6450 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_897
timestamp 1300117811
transform -1 0 6450 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_898
timestamp 1300117811
transform -1 0 6450 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_899
timestamp 1300117811
transform -1 0 6450 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_900
timestamp 1300117811
transform -1 0 6450 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_901
timestamp 1300117811
transform -1 0 6450 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_902
timestamp 1300117811
transform -1 0 6450 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_903
timestamp 1300117811
transform -1 0 6450 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_904
timestamp 1300117811
transform -1 0 6450 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_905
timestamp 1300117811
transform -1 0 6450 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_906
timestamp 1300117811
transform -1 0 6450 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_907
timestamp 1300117811
transform -1 0 6450 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_908
timestamp 1300117811
transform -1 0 6450 0 -1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_909
timestamp 1300117811
transform -1 0 6450 0 -1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_910
timestamp 1300117811
transform -1 0 6450 0 -1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_911
timestamp 1300117811
transform -1 0 6450 0 -1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_912
timestamp 1300117811
transform -1 0 6450 0 -1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_913
timestamp 1300117811
transform -1 0 6450 0 -1 13072
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 6450 0 -1 12986
box 0 0 6450 1720
use fillpp_mt fillpp_mt_914
timestamp 1300117811
transform -1 0 6450 0 -1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_915
timestamp 1300117811
transform -1 0 6450 0 -1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_916
timestamp 1300117811
transform -1 0 6450 0 -1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_917
timestamp 1300117811
transform -1 0 6450 0 -1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_918
timestamp 1300117811
transform -1 0 6450 0 -1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_919
timestamp 1300117811
transform -1 0 6450 0 -1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_920
timestamp 1300117811
transform -1 0 6450 0 -1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_921
timestamp 1300117811
transform -1 0 6450 0 -1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_922
timestamp 1300117811
transform -1 0 6450 0 -1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_923
timestamp 1300117811
transform -1 0 6450 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_924
timestamp 1300117811
transform -1 0 6450 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_925
timestamp 1300117811
transform -1 0 6450 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_926
timestamp 1300117811
transform -1 0 6450 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_927
timestamp 1300117811
transform -1 0 6450 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_928
timestamp 1300117811
transform -1 0 6450 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_929
timestamp 1300117811
transform -1 0 6450 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_930
timestamp 1300117811
transform -1 0 6450 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_931
timestamp 1300117811
transform -1 0 6450 0 -1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_932
timestamp 1300117811
transform -1 0 6450 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_933
timestamp 1300117811
transform -1 0 6450 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_934
timestamp 1300117811
transform -1 0 6450 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_935
timestamp 1300117811
transform -1 0 6450 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_936
timestamp 1300117811
transform -1 0 6450 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_937
timestamp 1300117811
transform -1 0 6450 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_938
timestamp 1300117811
transform -1 0 6450 0 -1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_939
timestamp 1300117811
transform -1 0 6450 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_940
timestamp 1300117811
transform -1 0 6450 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_941
timestamp 1300117811
transform -1 0 6450 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_942
timestamp 1300117811
transform -1 0 6450 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_943
timestamp 1300117811
transform -1 0 6450 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_944
timestamp 1300117811
transform -1 0 6450 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_945
timestamp 1300117811
transform -1 0 6450 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_946
timestamp 1300117811
transform -1 0 6450 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_947
timestamp 1300117811
transform -1 0 6450 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_948
timestamp 1300117811
transform -1 0 6450 0 -1 8342
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 6450 0 -1 8256
box 0 0 6450 1720
use control control_0
timestamp 1395747878
transform 1 0 11387 0 1 7589
box 0 0 27735 8204
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 41538 0 1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 41538 0 1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 41538 0 1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 41538 0 1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 41538 0 1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 41538 0 1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 41538 0 1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 41538 0 1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 41538 0 1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 41538 0 1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 41538 0 1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 41538 0 1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 41538 0 1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 41538 0 1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 41538 0 1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 41538 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 41538 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 41538 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 41538 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 41538 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 41538 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 41538 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 41538 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 41538 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 41538 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 41538 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 41538 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 41538 0 1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 41538 0 1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 41538 0 1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 41538 0 1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 41538 0 1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 41538 0 1 12986
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 41538 0 1 11266
box 0 0 6450 1720
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 41538 0 1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 41538 0 1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 41538 0 1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 41538 0 1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 41538 0 1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 41538 0 1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 41538 0 1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 41538 0 1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 41538 0 1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 41538 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 41538 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 41538 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 41538 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 41538 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 41538 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 41538 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 41538 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 41538 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 41538 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 41538 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 41538 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 41538 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 41538 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 41538 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 41538 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 41538 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 41538 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 41538 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 41538 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 41538 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 41538 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 41538 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 41538 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 41538 0 1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 41538 0 1 8256
box 0 0 6450 86
use fillpp_mt fillpp_mt_949
timestamp 1300117811
transform -1 0 6450 0 -1 6536
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 41538 0 1 6536
box 0 0 6450 1720
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 41538 0 1 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 0 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 6450 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 6536 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6622 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 8342 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 8428 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 8514 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 8600 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8686 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8772 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8858 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8944 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 9030 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 9116 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 9202 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 9288 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 9374 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 9460 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 9546 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9632 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9718 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9804 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9890 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9976 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 10062 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 10148 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 10234 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 10320 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 10406 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 10492 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 10578 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 10664 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10750 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 12470 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 12556 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 12642 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 12728 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 12814 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12900 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12986 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 13072 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 13158 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 13244 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 13330 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 13416 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 13502 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 13588 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 13674 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 13760 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 13846 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 13932 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 14018 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 14104 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 14190 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 14276 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 14362 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 14448 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 14534 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 14620 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 14706 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 14792 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 14878 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 16598 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 16684 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 16770 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 16856 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 16942 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 17028 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 17114 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 17200 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 17286 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 17372 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 17458 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 17544 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 17630 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 17716 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 17802 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 17888 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 17974 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 18060 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 18146 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 18232 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 18318 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 18404 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 18490 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 18576 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 18662 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 18748 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 18834 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 18920 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 19006 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 20726 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 20812 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 20898 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 20984 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 21070 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 21156 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 21242 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 21328 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 21414 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 21500 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 21586 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 21672 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 21758 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 21844 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 21930 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 22016 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 22102 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 22188 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 22274 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 22360 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 22446 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 22532 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 22618 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 22704 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 22790 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 22876 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 22962 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 23048 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 23134 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 24854 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 24940 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 25026 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 25112 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 25198 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 25284 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 25370 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 25456 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 25542 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 25628 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 25714 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 25800 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 25886 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 25972 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 26058 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 26144 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 26230 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 26316 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 26402 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 26488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 26574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 26660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 26746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 26832 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 26918 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 27004 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 27090 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 27176 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 27262 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 28982 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 29068 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 29154 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 29240 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 29326 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 29412 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 29498 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 29584 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 29670 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 29756 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 29842 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 29928 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 30014 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 30100 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 30186 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 30272 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 30358 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 30444 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 30530 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 30616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 30702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 30788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 30874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 30960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 31046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 31132 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 31218 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 31304 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 31390 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 0 1 33110 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 0 1 33196 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 0 1 33282 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 0 1 33368 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 0 1 33454 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 0 1 33540 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 0 1 33626 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 0 1 33712 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 0 1 33798 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 0 1 33884 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 0 1 33970 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 0 1 34056 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 0 1 34142 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 0 1 34228 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 0 1 34314 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 0 1 34400 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 0 1 34486 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 0 1 34572 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 0 1 34658 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 0 1 34744 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 0 1 34830 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 0 1 34916 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 0 1 35002 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 0 1 35088 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 0 1 35174 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 0 1 35260 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 0 1 35346 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 0 1 35432 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 35518 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 0 1 37238 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 0 1 37324 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 0 1 37410 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 0 1 37496 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 0 1 37582 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 0 1 37668 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 0 1 37754 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 0 1 37840 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 0 1 37926 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 0 1 38012 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 0 1 38098 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 0 1 38184 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 0 1 38270 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 0 1 38356 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 0 1 38442 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 0 1 38528 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 0 1 38614 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 0 1 38700 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 0 1 38786 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 0 1 38872 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 0 1 38958 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 0 1 39044 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 0 1 39130 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 0 1 39216 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 0 1 39302 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 0 1 39388 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 0 1 39474 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 0 1 39560 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 39646 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 0 1 41366 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 0 1 41452 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 47988 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 6702 78 8262 1638 0 nIRQ
rlabel metal4 10830 78 12390 1638 0 Data[0]
rlabel metal4 14958 78 16518 1638 0 Data[1]
rlabel metal4 19086 78 20646 1638 0 Data[2]
rlabel metal4 23214 78 24774 1638 0 vdde!
rlabel metal4 27342 78 28902 1638 0 Data[3]
rlabel metal4 31470 78 33030 1638 0 Data[4]
rlabel metal4 35598 78 37158 1638 0 Data[5]
rlabel metal4 39726 78 41286 1638 0 gnde!
rlabel metal4 46350 6616 47910 8176 0 Data[6]
rlabel metal4 46350 11346 47910 12906 0 Data[7]
rlabel metal4 46350 16076 47910 17636 0 Data[8]
rlabel metal4 46350 20806 47910 22366 0 gnde!
rlabel metal4 46350 25536 47910 27096 0 GND!
rlabel metal4 46350 30266 47910 31826 0 Data[9]
rlabel metal4 46350 34996 47910 36556 0 Data[10]
rlabel metal4 46350 39726 47910 41286 0 Data[11]
rlabel metal4 39726 46264 41286 47824 0 vdde!
rlabel metal4 35598 46264 37158 47824 0 Data[12]
rlabel metal4 31470 46264 33030 47824 0 Data[13]
rlabel metal4 27342 46264 28902 47824 0 Data[14]
rlabel metal4 23214 46264 24774 47824 0 gnde!
rlabel metal4 19086 46264 20646 47824 0 Data[15]
rlabel metal4 14958 46264 16518 47824 0 ALE
rlabel metal4 10830 46264 12390 47824 0 nME
rlabel metal4 6702 46264 8262 47824 0 nWait
rlabel metal4 78 39726 1638 41286 0 nOE
rlabel metal4 78 34996 1638 36556 0 RnW
rlabel metal4 78 30266 1638 31826 0 SDO
rlabel metal4 78 25536 1638 27096 0 Vdd!
rlabel metal4 78 20806 1638 22366 0 SDI
rlabel metal4 78 16076 1638 17636 0 Test
rlabel metal4 78 11346 1638 12906 0 Clock
rlabel metal4 78 6616 1638 8176 0 nReset
<< end >>
