magic
tech c035u
timestamp 1394128586
<< error_s >>
rect 4065 2045 4079 2050
rect 6788 423 6806 821
rect 6788 22 6812 423
use ALUDecoder ALUDecoder_0
timestamp 1394128449
transform 1 0 130 0 1 2040
box -130 0 7234 1481
use ALUSlice ALUSlice_1
timestamp 1394120777
transform 1 0 0 0 1 998
box 0 0 6788 1042
use LLIcell_U LLIcell_U_0
timestamp 1393855556
transform 1 0 6788 0 1 998
box 0 0 192 1042
use ALUSlice ALUSlice_0
timestamp 1394120777
transform 1 0 0 0 1 -44
box 0 0 6788 1042
use LLIcell_L LLIcell_L_0
timestamp 1393855517
transform 1 0 6788 0 1 -44
box 0 0 192 1042
<< end >>
