magic
tech c035u
timestamp 1396906989
<< metal1 >>
rect 21120 39730 21130 39773
rect 21168 39730 21178 39773
rect 21120 39720 21178 39730
rect 21120 39226 21130 39720
rect 21216 39253 21226 39773
rect 24552 39757 24562 39773
rect 24600 39730 24610 39773
rect 28080 39757 28090 39773
rect 21480 39720 24610 39730
rect 21480 39706 21490 39720
rect 28128 39730 28138 39773
rect 24637 39720 28138 39730
rect 31584 39730 31594 39773
rect 31632 39757 31642 39773
rect 31776 39757 31786 39773
rect 38640 39730 38650 39773
rect 38688 39757 38698 39773
rect 38832 39757 38842 39773
rect 42168 39730 42178 39773
rect 42216 39757 42226 39773
rect 42360 39757 42370 39773
rect 45696 39733 45706 39773
rect 45744 39757 45754 39773
rect 45888 39757 45898 39773
rect 31584 39720 45695 39730
rect 45720 39720 47050 39730
rect 21456 39696 21490 39706
rect 21456 39685 21466 39696
rect 21517 39696 24551 39706
rect 24565 39696 28079 39706
rect 45720 39706 45730 39720
rect 31645 39696 45730 39706
rect 46837 39696 47015 39706
rect 47040 39706 47050 39720
rect 47040 39696 47074 39706
rect 21493 39672 24623 39682
rect 21432 39648 21503 39658
rect 21432 39253 21442 39648
rect 21456 39253 21466 39623
rect 21480 39253 21490 39623
rect 28080 39589 28090 39695
rect 38701 39672 47039 39682
rect 47064 39682 47074 39696
rect 47064 39672 47087 39682
rect 31776 39589 31786 39671
rect 38845 39648 47122 39658
rect 47112 39634 47122 39648
rect 45901 39624 47074 39634
rect 47112 39624 47135 39634
rect 42216 39589 42226 39623
rect 42360 39589 42370 39623
rect 45696 39610 45706 39623
rect 47064 39610 47074 39624
rect 45696 39600 47002 39610
rect 47064 39600 47159 39610
rect 45757 39576 45767 39586
rect 46992 39586 47002 39600
rect 46992 39576 47207 39586
rect 27888 39552 47002 39562
rect 27888 39469 27898 39552
rect 45757 39528 46871 39538
rect 46992 39538 47002 39552
rect 47053 39552 47231 39562
rect 46992 39528 47255 39538
rect 28080 39469 28090 39527
rect 31776 39469 31786 39527
rect 38869 39504 47111 39514
rect 47149 39504 47290 39514
rect 38664 39480 47194 39490
rect 38664 39469 38674 39480
rect 47184 39469 47194 39480
rect 39037 39456 47135 39466
rect 47280 39466 47290 39504
rect 47280 39456 47314 39466
rect 25464 39432 47290 39442
rect 21120 39216 21514 39226
rect 21408 39192 21431 39202
rect 20207 38832 20266 38842
rect 20256 38818 20266 38832
rect 21216 38821 21226 39191
rect 20256 38808 20279 38818
rect 21408 38794 21418 39192
rect 21504 39202 21514 39216
rect 21504 39192 22007 39202
rect 20207 38784 21418 38794
rect 21432 39168 22138 39178
rect 20256 34810 20266 38784
rect 20280 34837 20290 38759
rect 20256 34800 20314 34810
rect 20207 34776 20266 34786
rect 20256 34765 20266 34776
rect 20304 34738 20314 34800
rect 20207 34728 20314 34738
rect 20256 30781 20266 34703
rect 20280 30781 20290 34703
rect 20304 30781 20314 34728
rect 21216 30781 21226 38759
rect 21432 30754 21442 39168
rect 22128 39157 22138 39168
rect 25464 39157 25474 39432
rect 47280 39421 47290 39432
rect 47304 39421 47314 39456
rect 26856 39408 47074 39418
rect 26856 39373 26866 39408
rect 47064 39397 47074 39408
rect 36144 39384 47039 39394
rect 36144 39373 36154 39384
rect 47160 39394 47170 39407
rect 47160 39384 47327 39394
rect 36877 39360 47159 39370
rect 47221 39360 47351 39370
rect 26664 39336 46991 39346
rect 26664 39277 26674 39336
rect 47101 39336 47375 39346
rect 35880 39312 47207 39322
rect 26856 39277 26866 39311
rect 27888 39277 27898 39311
rect 28080 39277 28090 39311
rect 31776 39277 31786 39311
rect 35880 39277 35890 39312
rect 47245 39312 47399 39322
rect 38928 39288 47231 39298
rect 38928 39277 38938 39288
rect 47317 39288 47423 39298
rect 42373 39264 45743 39274
rect 45781 39264 47314 39274
rect 47304 39253 47314 39264
rect 47389 39264 47447 39274
rect 25704 39240 47087 39250
rect 25704 39157 25714 39240
rect 47352 39250 47362 39263
rect 47352 39240 47506 39250
rect 31789 39216 47482 39226
rect 26664 39157 26674 39215
rect 26856 39157 26866 39215
rect 27888 39157 27898 39215
rect 28080 39178 28090 39215
rect 42229 39192 46858 39202
rect 28080 39168 46823 39178
rect 46848 39178 46858 39192
rect 46885 39192 47386 39202
rect 46848 39168 47362 39178
rect 46824 39157 46834 39167
rect 20207 30744 21442 30754
rect 20304 30706 20314 30719
rect 20207 30696 20314 30706
rect 20256 26794 20266 30671
rect 20280 26821 20290 30671
rect 20256 26784 20314 26794
rect 20207 26760 20266 26770
rect 20256 22834 20266 26760
rect 20280 22861 20290 26759
rect 20304 22861 20314 26784
rect 20256 22824 20338 22834
rect 20207 22800 20266 22810
rect 20256 18805 20266 22800
rect 20280 19618 20290 22799
rect 20304 19645 20314 22799
rect 20328 19642 20338 22824
rect 21216 19645 21226 30719
rect 21456 19666 21466 39143
rect 21445 19656 21466 19666
rect 20328 19632 21119 19642
rect 21480 19642 21490 39143
rect 46992 36469 47002 39143
rect 47016 36469 47026 39143
rect 47040 36469 47050 39143
rect 47064 36469 47074 39143
rect 47088 36469 47098 39143
rect 47112 36469 47122 39143
rect 47136 36469 47146 39143
rect 47160 36469 47170 39143
rect 47184 36469 47194 39143
rect 47208 36469 47218 39143
rect 47232 36469 47242 39143
rect 47256 36469 47266 39143
rect 47280 36469 47290 39143
rect 47304 36469 47314 39143
rect 47328 36469 47338 39143
rect 47352 36469 47362 39168
rect 47376 36469 47386 39192
rect 47400 36469 47410 39191
rect 47424 36469 47434 39191
rect 47448 36469 47458 39191
rect 47472 36442 47482 39216
rect 47496 39034 47506 39240
rect 47496 39024 50307 39034
rect 50256 39013 50266 39024
rect 50232 38976 50307 38986
rect 50232 38866 50242 38976
rect 50256 38869 50266 38951
rect 46968 36440 47482 36442
rect 46943 36432 47482 36440
rect 50208 38856 50242 38866
rect 46943 36430 46978 36432
rect 46943 36370 46978 36374
rect 47448 36370 47458 36407
rect 46943 36364 47458 36370
rect 46968 36360 47458 36364
rect 46992 35365 47002 36335
rect 47016 35365 47026 36335
rect 47040 35365 47050 36335
rect 47064 35365 47074 36335
rect 47088 35365 47098 36335
rect 47112 35365 47122 36335
rect 47136 35365 47146 36335
rect 47160 35365 47170 36335
rect 47184 35365 47194 36335
rect 47208 35365 47218 36335
rect 47232 35365 47242 36335
rect 47256 35365 47266 36335
rect 47280 35365 47290 36335
rect 47304 35365 47314 36335
rect 47328 35365 47338 36335
rect 47352 35365 47362 36335
rect 47376 35365 47386 36335
rect 47400 35365 47410 36335
rect 47424 35338 47434 36335
rect 46968 35329 47434 35338
rect 46943 35328 47434 35329
rect 46943 35319 46978 35328
rect 47400 35266 47410 35303
rect 46968 35263 47410 35266
rect 46943 35256 47410 35263
rect 46943 35253 46978 35256
rect 46992 34237 47002 35231
rect 47016 34237 47026 35231
rect 47040 34237 47050 35231
rect 47064 34237 47074 35231
rect 47088 34237 47098 35231
rect 47112 34237 47122 35231
rect 47136 34237 47146 35231
rect 47160 34237 47170 35231
rect 47184 34237 47194 35231
rect 47208 34237 47218 35231
rect 47232 34237 47242 35231
rect 47256 34237 47266 35231
rect 47280 34237 47290 35231
rect 47304 34237 47314 35231
rect 47328 34237 47338 35231
rect 47352 34237 47362 35231
rect 46943 34210 46978 34218
rect 47376 34210 47386 35231
rect 50208 34978 50218 38856
rect 50232 38832 50307 38842
rect 50232 34981 50242 38832
rect 50256 35002 50266 38807
rect 50256 34992 50307 35002
rect 50256 34981 50266 34992
rect 50184 34968 50218 34978
rect 50184 34861 50194 34968
rect 50208 34944 50307 34954
rect 50208 34861 50218 34944
rect 50232 34834 50242 34919
rect 50256 34837 50266 34919
rect 46943 34208 47386 34210
rect 46968 34200 47386 34208
rect 50160 34824 50242 34834
rect 46943 34142 46978 34152
rect 46968 34138 46978 34142
rect 47352 34138 47362 34175
rect 46968 34128 47362 34138
rect 46992 33133 47002 34103
rect 47016 33133 47026 34103
rect 47040 33133 47050 34103
rect 47064 33133 47074 34103
rect 47088 33133 47098 34103
rect 47112 33133 47122 34103
rect 47136 33133 47146 34103
rect 47160 33133 47170 34103
rect 47184 33133 47194 34103
rect 47208 33133 47218 34103
rect 47232 33133 47242 34103
rect 47256 33133 47266 34103
rect 47280 33133 47290 34103
rect 47304 33133 47314 34103
rect 46943 33106 46978 33107
rect 47328 33106 47338 34103
rect 46943 33097 47338 33106
rect 46968 33096 47338 33097
rect 46943 33034 46978 33041
rect 47304 33034 47314 33071
rect 46943 33031 47314 33034
rect 46968 33024 47314 33031
rect 46992 32029 47002 32999
rect 47016 32029 47026 32999
rect 47040 32029 47050 32999
rect 47064 32029 47074 32999
rect 47088 32029 47098 32999
rect 47112 32029 47122 32999
rect 47136 32029 47146 32999
rect 47160 32029 47170 32999
rect 47184 32029 47194 32999
rect 47208 32029 47218 32999
rect 47232 32029 47242 32999
rect 47256 32029 47266 32999
rect 47280 32029 47290 32999
rect 50160 32002 50170 34824
rect 50232 34800 50307 34810
rect 46968 31996 50170 32002
rect 46943 31992 50170 31996
rect 46943 31986 46978 31992
rect 50184 31930 50194 34799
rect 46943 31920 50194 31930
rect 46992 30901 47002 31895
rect 47016 30901 47026 31895
rect 47040 30901 47050 31895
rect 47064 30901 47074 31895
rect 47088 30901 47098 31895
rect 47112 30901 47122 31895
rect 47136 30901 47146 31895
rect 47160 30901 47170 31895
rect 47184 30901 47194 31895
rect 47208 30901 47218 31895
rect 47232 30901 47242 31895
rect 47256 30901 47266 31895
rect 47280 30901 47290 31895
rect 50208 30973 50218 34799
rect 50232 30946 50242 34800
rect 50256 30970 50266 34775
rect 50256 30960 50307 30970
rect 50256 30949 50266 30960
rect 50184 30936 50242 30946
rect 46943 30875 46978 30885
rect 46968 30874 46978 30875
rect 50184 30874 50194 30936
rect 50232 30912 50307 30922
rect 46968 30864 50194 30874
rect 50208 30826 50218 30911
rect 46968 30819 50218 30826
rect 46943 30816 50218 30819
rect 46943 30809 46978 30816
rect 50232 30805 50242 30912
rect 50256 30805 50266 30887
rect 46992 29797 47002 30791
rect 47016 29797 47026 30791
rect 47040 29797 47050 30791
rect 47064 29797 47074 30791
rect 47088 29797 47098 30791
rect 47112 29797 47122 30791
rect 47136 29797 47146 30791
rect 47160 29797 47170 30791
rect 47184 29797 47194 30791
rect 47208 29797 47218 30791
rect 47232 29797 47242 30791
rect 47256 29797 47266 30791
rect 47280 29797 47290 30791
rect 50208 30768 50307 30778
rect 46943 29770 46978 29774
rect 50208 29770 50218 30768
rect 46943 29764 50218 29770
rect 46968 29760 50218 29764
rect 46943 29698 46978 29708
rect 50232 29698 50242 30743
rect 46968 29688 50242 29698
rect 46992 28693 47002 29663
rect 47016 28693 47026 29663
rect 47040 28693 47050 29663
rect 47064 28693 47074 29663
rect 47088 28693 47098 29663
rect 47112 28693 47122 29663
rect 47136 28693 47146 29663
rect 47160 28693 47170 29663
rect 47184 28693 47194 29663
rect 47208 28693 47218 29663
rect 47232 28693 47242 29663
rect 47256 28690 47266 29663
rect 47280 28717 47290 29663
rect 47256 28680 47314 28690
rect 46968 28663 47266 28666
rect 46943 28656 47266 28663
rect 46943 28653 46978 28656
rect 47256 28618 47266 28656
rect 47304 28645 47314 28680
rect 47256 28608 47338 28618
rect 46943 28594 46978 28597
rect 46943 28587 47266 28594
rect 46968 28584 47266 28587
rect 46992 27565 47002 28559
rect 47016 27565 47026 28559
rect 46943 27542 46978 27552
rect 47040 27562 47050 28559
rect 47064 27589 47074 28559
rect 47088 27589 47098 28559
rect 47112 27589 47122 28559
rect 47136 27589 47146 28559
rect 47160 27589 47170 28559
rect 47184 27589 47194 28559
rect 47208 27589 47218 28559
rect 47232 27589 47242 28559
rect 47256 27589 47266 28584
rect 47280 27589 47290 28583
rect 47304 27589 47314 28583
rect 47328 27589 47338 28608
rect 47040 27552 47362 27562
rect 46968 27538 46978 27542
rect 47352 27541 47362 27552
rect 46968 27528 47039 27538
rect 47029 27504 47386 27514
rect 46968 27486 47026 27490
rect 46943 27480 47026 27486
rect 46943 27476 46978 27480
rect 46992 26461 47002 27455
rect 47016 26461 47026 27480
rect 47040 26461 47050 27479
rect 47064 26458 47074 27479
rect 47088 26485 47098 27479
rect 47112 26485 47122 27479
rect 47136 26485 47146 27479
rect 47160 26485 47170 27479
rect 47184 26485 47194 27479
rect 47208 26485 47218 27479
rect 47232 26485 47242 27479
rect 47256 26485 47266 27479
rect 47280 26485 47290 27479
rect 47304 26485 47314 27479
rect 47328 26485 47338 27479
rect 47352 26485 47362 27479
rect 47376 26794 47386 27504
rect 50256 26821 50266 30743
rect 47376 26784 50279 26794
rect 47064 26448 47386 26458
rect 46943 26434 46978 26441
rect 46943 26431 47074 26434
rect 46968 26424 47074 26431
rect 47064 26413 47074 26424
rect 47376 26413 47386 26448
rect 46992 26386 47002 26399
rect 46992 26376 47410 26386
rect 46943 26365 46978 26375
rect 46968 26362 46978 26365
rect 46968 26352 47002 26362
rect 46992 25357 47002 26352
rect 47016 25357 47026 26351
rect 47040 25357 47050 26351
rect 47064 25357 47074 26351
rect 47088 25357 47098 26351
rect 47112 25354 47122 26351
rect 47136 25381 47146 26351
rect 47160 25381 47170 26351
rect 47184 25381 47194 26351
rect 47208 25381 47218 26351
rect 47232 25381 47242 26351
rect 47256 25381 47266 26351
rect 47280 25381 47290 26351
rect 47304 25381 47314 26351
rect 47328 25381 47338 26351
rect 47352 25381 47362 26351
rect 47376 25381 47386 26351
rect 47400 25381 47410 26376
rect 47112 25344 47434 25354
rect 46943 25320 47122 25330
rect 47112 25285 47122 25320
rect 47136 25285 47146 25319
rect 47160 25285 47170 25319
rect 47184 25285 47194 25319
rect 47208 25285 47218 25319
rect 47232 25282 47242 25319
rect 47424 25309 47434 25344
rect 47232 25272 47458 25282
rect 46943 25258 46978 25264
rect 46943 25254 47242 25258
rect 46968 25248 47242 25254
rect 46992 24253 47002 25223
rect 47016 24253 47026 25223
rect 47040 24253 47050 25223
rect 47064 24253 47074 25223
rect 47088 24253 47098 25223
rect 47112 24253 47122 25223
rect 47136 24253 47146 25223
rect 47160 24253 47170 25223
rect 47184 24253 47194 25223
rect 47208 24253 47218 25223
rect 47232 24253 47242 25248
rect 47256 24250 47266 25247
rect 47280 24277 47290 25247
rect 47304 24277 47314 25247
rect 47328 24277 47338 25247
rect 47352 24277 47362 25247
rect 47376 24277 47386 25247
rect 47400 24277 47410 25247
rect 47424 24277 47434 25247
rect 47448 24277 47458 25272
rect 47256 24240 47482 24250
rect 46968 24219 47266 24226
rect 46943 24216 47266 24219
rect 46943 24209 46978 24216
rect 47256 24205 47266 24216
rect 47472 24205 47482 24240
rect 47136 24178 47146 24191
rect 47136 24168 47506 24178
rect 46968 24153 47146 24154
rect 46943 24144 47146 24153
rect 46943 24143 46978 24144
rect 46992 23125 47002 24119
rect 47016 23125 47026 24119
rect 47040 23125 47050 24119
rect 47064 23125 47074 24119
rect 47088 23122 47098 24119
rect 47112 23149 47122 24119
rect 47136 23149 47146 24144
rect 47160 23149 47170 24143
rect 47184 23149 47194 24143
rect 47208 23149 47218 24143
rect 47232 23149 47242 24143
rect 47256 23149 47266 24143
rect 47280 23149 47290 24143
rect 47304 23149 47314 24143
rect 47328 23149 47338 24143
rect 47352 23149 47362 24143
rect 47376 23149 47386 24143
rect 47400 23149 47410 24143
rect 47424 23149 47434 24143
rect 47448 23149 47458 24143
rect 47472 23149 47482 24143
rect 47496 23149 47506 24168
rect 47088 23112 47530 23122
rect 46943 23098 46978 23108
rect 47520 23101 47530 23112
rect 46968 23088 47098 23098
rect 47088 23077 47098 23088
rect 47376 23074 47386 23087
rect 47376 23064 47554 23074
rect 46968 23042 47386 23050
rect 46943 23040 47386 23042
rect 46943 23032 46978 23040
rect 46992 22021 47002 23015
rect 47016 22021 47026 23015
rect 47040 22021 47050 23015
rect 47064 22021 47074 23015
rect 47088 22021 47098 23015
rect 47112 22021 47122 23015
rect 47136 22021 47146 23015
rect 47160 22021 47170 23015
rect 47184 22021 47194 23015
rect 47208 22021 47218 23015
rect 47232 22018 47242 23015
rect 47256 22045 47266 23015
rect 47280 22045 47290 23015
rect 47304 22045 47314 23015
rect 47328 22045 47338 23015
rect 47352 22045 47362 23015
rect 47376 22045 47386 23040
rect 47400 22045 47410 23039
rect 47424 22045 47434 23039
rect 47448 22045 47458 23039
rect 47472 22045 47482 23039
rect 47496 22045 47506 23039
rect 47520 22045 47530 23039
rect 47544 22045 47554 23064
rect 47232 22008 47578 22018
rect 46943 21994 46978 21997
rect 46943 21987 47242 21994
rect 46968 21984 47242 21987
rect 47232 21973 47242 21984
rect 47568 21973 47578 22008
rect 47160 21946 47170 21959
rect 47160 21936 47602 21946
rect 46943 21922 46978 21931
rect 46943 21921 47170 21922
rect 46968 21912 47170 21921
rect 46992 20917 47002 21887
rect 47016 20917 47026 21887
rect 47040 20917 47050 21887
rect 47064 20917 47074 21887
rect 47088 20917 47098 21887
rect 47112 20917 47122 21887
rect 47136 20917 47146 21887
rect 47160 20917 47170 21912
rect 47184 20917 47194 21911
rect 47208 20917 47218 21911
rect 47232 20917 47242 21911
rect 47256 20917 47266 21911
rect 47280 20917 47290 21911
rect 47304 20917 47314 21911
rect 47328 20917 47338 21911
rect 47352 20917 47362 21911
rect 47376 20917 47386 21911
rect 47400 20917 47410 21911
rect 47424 20917 47434 21911
rect 47448 20917 47458 21911
rect 47472 20917 47482 21911
rect 47496 20917 47506 21911
rect 47520 20917 47530 21911
rect 47544 20917 47554 21911
rect 47568 20914 47578 21911
rect 47592 20941 47602 21936
rect 47568 20904 47626 20914
rect 46968 20886 47578 20890
rect 46943 20880 47578 20886
rect 46943 20876 46978 20880
rect 47568 20869 47578 20880
rect 47616 20869 47626 20904
rect 47208 20842 47218 20855
rect 47208 20832 47650 20842
rect 46943 20818 46978 20820
rect 46943 20810 47218 20818
rect 46968 20808 47218 20810
rect 46992 19789 47002 20783
rect 47016 19789 47026 20783
rect 47040 19789 47050 20783
rect 47064 19789 47074 20783
rect 47088 19789 47098 20783
rect 47112 19789 47122 20783
rect 47136 19789 47146 20783
rect 47160 19789 47170 20783
rect 47184 19789 47194 20783
rect 47208 19789 47218 20808
rect 47232 19789 47242 20807
rect 47256 19786 47266 20807
rect 47280 19813 47290 20807
rect 47304 19813 47314 20807
rect 47328 19813 47338 20807
rect 47352 19813 47362 20807
rect 47376 19813 47386 20807
rect 47400 19813 47410 20807
rect 47424 19813 47434 20807
rect 47448 19813 47458 20807
rect 47472 19813 47482 20807
rect 47496 19813 47506 20807
rect 47520 19813 47530 20807
rect 47544 19813 47554 20807
rect 47568 19813 47578 20807
rect 47592 19813 47602 20807
rect 47616 19813 47626 20807
rect 47640 19813 47650 20832
rect 47256 19776 47674 19786
rect 46943 19765 46978 19775
rect 47664 19765 47674 19776
rect 46968 19762 46978 19765
rect 46968 19752 47255 19762
rect 47245 19728 47698 19738
rect 46968 19709 47242 19714
rect 46943 19704 47242 19709
rect 46943 19699 46978 19704
rect 21397 19632 21490 19642
rect 46992 19621 47002 19679
rect 47016 19621 47026 19679
rect 47040 19621 47050 19679
rect 20280 19608 21490 19618
rect 20207 18768 20290 18778
rect 20256 14749 20266 18743
rect 20280 18370 20290 18768
rect 20304 18397 20314 19583
rect 21120 19498 21130 19583
rect 21216 19525 21226 19583
rect 21384 19525 21394 19583
rect 21432 19525 21442 19583
rect 21480 19525 21490 19608
rect 47064 19618 47074 19679
rect 47088 19645 47098 19679
rect 47112 19645 47122 19679
rect 47136 19645 47146 19679
rect 47160 19645 47170 19679
rect 47184 19645 47194 19679
rect 47208 19645 47218 19679
rect 47232 19645 47242 19704
rect 47256 19645 47266 19703
rect 47280 19645 47290 19703
rect 47304 19645 47314 19703
rect 47328 19645 47338 19703
rect 47352 19645 47362 19703
rect 47376 19645 47386 19703
rect 47400 19645 47410 19703
rect 47424 19645 47434 19703
rect 47448 19645 47458 19703
rect 47472 19645 47482 19703
rect 47496 19645 47506 19703
rect 47520 19645 47530 19703
rect 47544 19645 47554 19703
rect 47568 19645 47578 19703
rect 47592 19645 47602 19703
rect 47616 19645 47626 19703
rect 47640 19645 47650 19703
rect 47664 19645 47674 19703
rect 47688 19645 47698 19728
rect 47064 19608 47722 19618
rect 21584 19594 21594 19607
rect 21584 19584 21762 19594
rect 21752 19573 21762 19584
rect 21651 19546 21661 19559
rect 21651 19536 21786 19546
rect 21776 19525 21786 19536
rect 22008 19498 22018 19607
rect 21120 19488 22018 19498
rect 21216 18397 21226 19463
rect 21384 18397 21394 19463
rect 21432 18397 21442 19463
rect 21480 18397 21490 19463
rect 21536 18490 21546 19463
rect 21560 18517 21570 19424
rect 21604 18538 21614 19463
rect 21628 18590 21638 19463
rect 21680 18671 21690 19463
rect 21673 18661 21690 18671
rect 21704 18634 21714 19463
rect 21648 18624 21714 18634
rect 21648 18565 21658 18624
rect 21728 18610 21738 19488
rect 21752 18613 21762 19463
rect 21776 18613 21786 19463
rect 22008 18613 22018 19488
rect 23448 18613 23458 19607
rect 24240 18613 24250 19607
rect 24792 18613 24802 19607
rect 25008 18613 25018 19607
rect 25752 18613 25762 19607
rect 21696 18600 21738 18610
rect 21672 18565 21682 18599
rect 21696 18565 21706 18600
rect 25920 18610 25930 19607
rect 26304 18634 26314 19607
rect 26496 18658 26506 19607
rect 26712 18682 26722 19607
rect 26712 18672 26783 18682
rect 27456 18682 27466 19607
rect 27624 18709 27634 19607
rect 46128 19594 46138 19607
rect 46272 19594 46282 19607
rect 31008 19584 46138 19594
rect 46152 19584 46282 19594
rect 27456 18672 27671 18682
rect 26496 18648 29327 18658
rect 31008 18637 31018 19584
rect 42864 19560 45167 19570
rect 26304 18624 30191 18634
rect 37032 18613 37042 19559
rect 37224 18613 37234 19559
rect 37464 18613 37474 19559
rect 42864 18613 42874 19560
rect 46152 19570 46162 19584
rect 46368 19594 46378 19607
rect 46309 19584 46378 19594
rect 46416 19594 46426 19607
rect 46416 19584 47074 19594
rect 47064 19573 47074 19584
rect 47712 19573 47722 19608
rect 45205 19560 46162 19570
rect 46206 19560 46319 19570
rect 43704 19536 45911 19546
rect 43704 18613 43714 19536
rect 44544 19512 45191 19522
rect 44544 18613 44554 19512
rect 46206 18613 46216 19560
rect 46230 19536 46295 19546
rect 46230 18613 46240 19536
rect 46488 19546 46498 19559
rect 46488 19536 47746 19546
rect 47736 19522 47746 19536
rect 47736 19512 47770 19522
rect 46824 19498 46834 19511
rect 46824 19488 47746 19498
rect 46992 18613 47002 19463
rect 47016 18613 47026 19463
rect 47040 18613 47050 19463
rect 47064 18613 47074 19463
rect 47088 18613 47098 19463
rect 47112 18613 47122 19463
rect 47136 18613 47146 19463
rect 47160 18613 47170 19463
rect 47184 18613 47194 19463
rect 47208 18613 47218 19463
rect 47232 18613 47242 19463
rect 25920 18600 31895 18610
rect 47256 18586 47266 19463
rect 21720 18576 47266 18586
rect 47280 18586 47290 19463
rect 47304 18610 47314 19463
rect 47328 18634 47338 19463
rect 47352 18658 47362 19463
rect 47376 18682 47386 19463
rect 47400 18706 47410 19463
rect 47424 18730 47434 19463
rect 47448 18754 47458 19463
rect 47472 18778 47482 19463
rect 47496 18802 47506 19463
rect 47520 18826 47530 19463
rect 47544 18850 47554 19463
rect 47568 18874 47578 19463
rect 47592 18898 47602 19463
rect 47616 18922 47626 19463
rect 47640 18946 47650 19463
rect 47664 18970 47674 19463
rect 47688 18994 47698 19463
rect 47712 19018 47722 19463
rect 47736 19042 47746 19488
rect 47760 19066 47770 19512
rect 47760 19056 47903 19066
rect 47736 19032 49127 19042
rect 47712 19008 49415 19018
rect 47688 18984 49439 18994
rect 47664 18960 49463 18970
rect 47640 18936 49487 18946
rect 47616 18912 49511 18922
rect 47592 18888 49535 18898
rect 47568 18864 49559 18874
rect 47544 18840 49583 18850
rect 47520 18816 49607 18826
rect 50256 18826 50266 26759
rect 50256 18816 50307 18826
rect 50256 18805 50266 18816
rect 47496 18792 49631 18802
rect 47472 18768 50307 18778
rect 47448 18744 49655 18754
rect 47424 18720 49679 18730
rect 47400 18696 49703 18706
rect 47376 18672 49727 18682
rect 50256 18661 50266 18743
rect 47352 18648 49751 18658
rect 47328 18624 50307 18634
rect 47304 18600 49775 18610
rect 47280 18576 49799 18586
rect 21720 18565 21730 18576
rect 21787 18552 22223 18562
rect 25021 18552 25103 18562
rect 25765 18552 32735 18562
rect 47245 18552 49823 18562
rect 21604 18528 22247 18538
rect 23448 18538 23458 18551
rect 23448 18528 24215 18538
rect 24240 18538 24250 18551
rect 24240 18528 24263 18538
rect 24792 18538 24802 18551
rect 24792 18528 33575 18538
rect 21763 18504 25079 18514
rect 25117 18504 33599 18514
rect 21536 18480 24191 18490
rect 24229 18480 31871 18490
rect 31909 18480 35303 18490
rect 21685 18456 29303 18466
rect 29341 18456 36124 18466
rect 21560 18397 21570 18455
rect 21624 18418 21634 18455
rect 21685 18432 22168 18442
rect 22261 18432 26759 18442
rect 26797 18432 36172 18442
rect 37032 18442 37042 18551
rect 37224 18466 37234 18551
rect 37464 18490 37474 18551
rect 37464 18480 37823 18490
rect 37224 18456 38495 18466
rect 37032 18432 39431 18442
rect 21624 18408 27599 18418
rect 27637 18408 40319 18418
rect 21661 18384 30167 18394
rect 30205 18384 36148 18394
rect 36186 18384 38471 18394
rect 38509 18384 41074 18394
rect 20280 18360 22144 18370
rect 22237 18360 27647 18370
rect 27685 18360 39407 18370
rect 39445 18360 41039 18370
rect 41064 18370 41074 18384
rect 41064 18360 41578 18370
rect 21573 18336 24250 18346
rect 20304 14749 20314 18335
rect 21216 14749 21226 18335
rect 21384 18221 21394 18335
rect 21432 18253 21442 18335
rect 21480 18253 21490 18335
rect 24240 18325 24250 18336
rect 24277 18336 32722 18346
rect 32712 18325 32722 18336
rect 32749 18336 35290 18346
rect 35280 18325 35290 18336
rect 35317 18336 37810 18346
rect 37800 18325 37810 18336
rect 41568 18346 41578 18360
rect 37837 18336 41554 18346
rect 41568 18336 42034 18346
rect 41544 18325 41554 18336
rect 42024 18325 42034 18336
rect 42864 18325 42874 18551
rect 43704 18325 43714 18551
rect 44544 18325 44554 18551
rect 46205 18325 46215 18551
rect 46229 18325 46239 18551
rect 46992 18346 47002 18551
rect 47016 18370 47026 18551
rect 47040 18394 47050 18551
rect 47064 18421 47074 18551
rect 47088 18418 47098 18551
rect 47112 18442 47122 18551
rect 47136 18466 47146 18551
rect 47160 18490 47170 18551
rect 47184 18514 47194 18551
rect 47208 18538 47218 18551
rect 47208 18528 49847 18538
rect 50256 18538 50266 18599
rect 49885 18528 50266 18538
rect 47184 18504 49895 18514
rect 47160 18480 49919 18490
rect 47136 18456 49943 18466
rect 47112 18432 49991 18442
rect 47088 18408 50039 18418
rect 47040 18384 50159 18394
rect 47016 18360 50207 18370
rect 46992 18336 50266 18346
rect 21672 18253 21682 18311
rect 21696 18253 21706 18311
rect 21720 18253 21730 18311
rect 21384 18211 21743 18221
rect 21445 18187 21743 18197
rect 21480 14749 21490 18162
rect 21672 14722 21682 18162
rect 20207 14712 21682 14722
rect 20256 10717 20266 14687
rect 20207 10680 20290 10690
rect 20256 10186 20266 10655
rect 20280 10234 20290 10680
rect 20304 10387 20314 14687
rect 21216 14124 21226 14687
rect 21480 14151 21490 14687
rect 21696 14151 21706 18162
rect 21720 14151 21730 18162
rect 49416 18152 49426 18311
rect 49440 18152 49450 18311
rect 49464 18152 49474 18311
rect 49488 18173 49498 18311
rect 49512 18200 49522 18311
rect 49536 18200 49546 18311
rect 49560 18200 49570 18311
rect 49584 18200 49594 18311
rect 49608 18200 49618 18311
rect 49632 18200 49642 18311
rect 49656 18200 49666 18311
rect 49680 18200 49690 18311
rect 49704 18200 49714 18311
rect 49728 18200 49738 18311
rect 49752 18200 49762 18311
rect 49776 18200 49786 18311
rect 49800 18200 49810 18311
rect 49824 18200 49834 18311
rect 49848 18200 49858 18311
rect 49872 18200 49882 18311
rect 49896 18200 49906 18311
rect 49920 18200 49930 18311
rect 49944 18200 49954 18311
rect 49488 18163 49978 18173
rect 49488 18139 49871 18149
rect 49488 18128 49498 18139
rect 49405 18115 49487 18125
rect 49968 18125 49978 18163
rect 49872 18115 49978 18125
rect 49872 18101 49882 18115
rect 49405 18091 49882 18101
rect 49405 18067 49751 18077
rect 49776 18053 49786 18066
rect 49405 18043 49786 18053
rect 49405 18019 49583 18029
rect 49416 17101 49426 17994
rect 49440 17101 49450 17994
rect 49464 17101 49474 17994
rect 49488 17101 49498 17994
rect 49512 17101 49522 17994
rect 49536 17101 49546 17994
rect 49560 17101 49570 17994
rect 49608 17101 49618 18018
rect 49632 17101 49642 18018
rect 49656 17101 49666 18018
rect 49680 17101 49690 18018
rect 49704 17074 49714 18018
rect 49405 17064 49714 17074
rect 21216 14114 21743 14124
rect 21493 14090 21743 14100
rect 21696 10414 21706 14063
rect 21720 10414 21730 14063
rect 49416 13285 49426 17039
rect 49440 13285 49450 17039
rect 49464 13285 49474 17039
rect 49488 14794 49498 17039
rect 49512 14821 49522 17039
rect 49536 14821 49546 17039
rect 49560 14821 49570 17039
rect 49608 14821 49618 17039
rect 49632 14821 49642 17039
rect 49656 14821 49666 17039
rect 49680 14821 49690 17039
rect 49728 14821 49738 18018
rect 49800 14821 49810 18066
rect 49824 14821 49834 18066
rect 49848 14821 49858 18066
rect 49896 14821 49906 18090
rect 49920 14821 49930 18090
rect 49944 14821 49954 18090
rect 49992 14821 50002 18311
rect 50040 14821 50050 18311
rect 50160 14821 50170 18311
rect 50208 14821 50218 18311
rect 50256 14818 50266 18336
rect 50245 14808 50266 14818
rect 49488 14784 50307 14794
rect 50184 14770 50194 14784
rect 50184 14760 50255 14770
rect 49512 13285 49522 14759
rect 49536 13285 49546 14759
rect 49560 13285 49570 14759
rect 49608 13258 49618 14759
rect 49405 13248 49618 13258
rect 49416 11919 49426 13223
rect 49440 11919 49450 13223
rect 49464 11919 49474 13223
rect 49512 11919 49522 13223
rect 49536 11919 49546 13223
rect 49560 11919 49570 13223
rect 49632 11919 49642 14759
rect 49656 11919 49666 14759
rect 49680 11919 49690 14759
rect 49728 11919 49738 14759
rect 49800 11892 49810 14759
rect 49405 11882 49810 11892
rect 49405 11858 49655 11868
rect 49416 10749 49426 11833
rect 49440 10749 49450 11833
rect 49464 10749 49474 11833
rect 49512 10749 49522 11833
rect 49536 10749 49546 11833
rect 49560 10749 49570 11833
rect 49632 10749 49642 11833
rect 49680 10749 49690 11857
rect 49728 10749 49738 11857
rect 49824 10749 49834 14759
rect 49848 10749 49858 14759
rect 49896 10722 49906 14759
rect 49405 10712 49906 10722
rect 49405 10688 49679 10698
rect 49416 10546 49426 10663
rect 49440 10573 49450 10663
rect 49464 10573 49474 10663
rect 49512 10573 49522 10663
rect 49536 10573 49546 10663
rect 49560 10573 49570 10663
rect 49632 10573 49642 10663
rect 49728 10573 49738 10687
rect 49824 10573 49834 10687
rect 49848 10573 49858 10687
rect 49920 10573 49930 14759
rect 49944 10573 49954 14759
rect 49992 10573 50002 14759
rect 50040 10573 50050 14759
rect 50160 14602 50170 14759
rect 50221 14736 50307 14746
rect 50232 14629 50242 14711
rect 50256 14629 50266 14711
rect 50160 14592 50307 14602
rect 50232 10690 50242 14567
rect 50256 10738 50266 14567
rect 50256 10728 50307 10738
rect 50256 10717 50266 10728
rect 50232 10680 50307 10690
rect 50256 10573 50266 10655
rect 49416 10536 50307 10546
rect 20304 10377 21743 10387
rect 21672 10353 21743 10363
rect 21672 10261 21682 10353
rect 49440 10365 49450 10511
rect 49464 10365 49474 10511
rect 49512 10365 49522 10511
rect 49536 10365 49546 10511
rect 49560 10365 49570 10511
rect 49632 10338 49642 10511
rect 49405 10328 49642 10338
rect 21696 10261 21706 10319
rect 21720 10261 21730 10319
rect 49405 10304 49535 10314
rect 22200 10234 22210 10247
rect 20280 10224 22210 10234
rect 24744 10224 29735 10234
rect 21744 10200 22127 10210
rect 21744 10186 21754 10200
rect 20256 10176 21754 10186
rect 21672 9850 21682 10151
rect 21096 9840 21682 9850
rect 21096 9826 21106 9840
rect 21696 9826 21706 10151
rect 21072 9816 21106 9826
rect 21120 9816 21706 9826
rect 21720 9826 21730 10151
rect 21720 9816 24610 9826
rect 21072 9759 21082 9816
rect 21120 9759 21130 9816
rect 21168 9759 21178 9816
rect 24600 9759 24610 9816
rect 24744 9759 24754 10224
rect 29773 10224 32903 10234
rect 32941 10224 39215 10234
rect 39253 10224 45935 10234
rect 49464 10234 49474 10279
rect 49512 10237 49522 10279
rect 45973 10224 49474 10234
rect 49560 10210 49570 10303
rect 28128 10200 49570 10210
rect 28128 9853 28138 10200
rect 49728 10189 49738 10511
rect 49824 10189 49834 10511
rect 28272 10176 29759 10186
rect 28272 9853 28282 10176
rect 31800 10176 32927 10186
rect 31800 10165 31810 10176
rect 38869 10176 39239 10186
rect 42253 10176 45959 10186
rect 45997 10176 49511 10186
rect 49848 10162 49858 10511
rect 32917 10152 49858 10162
rect 29736 10042 29746 10151
rect 31656 10128 49439 10138
rect 31656 10069 31666 10128
rect 49920 10114 49930 10511
rect 39229 10104 49930 10114
rect 31800 10069 31810 10103
rect 38856 10069 38866 10103
rect 45912 10080 45983 10090
rect 45912 10069 45922 10080
rect 46008 10080 46727 10090
rect 46008 10066 46018 10080
rect 46741 10080 49727 10090
rect 45949 10056 46018 10066
rect 49824 10042 49834 10079
rect 29736 10032 49834 10042
rect 31656 9853 31666 10007
rect 31800 9853 31810 10007
rect 38856 9877 38866 10007
rect 42240 9877 42250 10007
rect 45912 9949 45922 10007
rect 49944 9949 49954 10511
rect 49992 9922 50002 10511
rect 45768 9912 50002 9922
rect 45768 9901 45778 9912
rect 50040 9901 50050 10511
rect 45960 9888 46007 9898
rect 45960 9874 45970 9888
rect 42397 9864 45970 9874
rect 50256 9874 50266 10511
rect 45997 9864 50266 9874
rect 38725 9840 50039 9850
rect 24792 9816 45983 9826
rect 24792 9759 24802 9816
rect 28128 9759 28138 9791
rect 28272 9759 28282 9791
rect 28320 9759 28330 9816
rect 31656 9759 31666 9791
rect 31800 9759 31810 9791
rect 31848 9759 31858 9816
rect 38712 9759 38722 9791
rect 38856 9759 38866 9791
rect 38904 9759 38914 9816
rect 42240 9759 42250 9791
rect 42384 9759 42394 9791
rect 42432 9759 42442 9816
rect 45768 9759 45778 9791
rect 45912 9759 45922 9791
rect 45960 9759 45970 9816
rect 46021 9816 49943 9826
<< m2contact >>
rect 24551 39743 24565 39757
rect 28079 39743 28093 39757
rect 24623 39719 24637 39733
rect 31631 39743 31645 39757
rect 31775 39743 31789 39757
rect 38687 39743 38701 39757
rect 38831 39743 38845 39757
rect 42215 39743 42229 39757
rect 42359 39743 42373 39757
rect 45743 39743 45757 39757
rect 45887 39743 45901 39757
rect 45695 39719 45709 39733
rect 21503 39695 21517 39709
rect 24551 39695 24565 39709
rect 28079 39695 28093 39709
rect 31631 39695 31645 39709
rect 46823 39695 46837 39709
rect 47015 39695 47029 39709
rect 21455 39671 21469 39685
rect 21479 39671 21493 39685
rect 24623 39671 24637 39685
rect 21503 39647 21517 39661
rect 21455 39623 21469 39637
rect 21479 39623 21493 39637
rect 31775 39671 31789 39685
rect 38687 39671 38701 39685
rect 47039 39671 47053 39685
rect 47087 39671 47101 39685
rect 38831 39647 38845 39661
rect 42215 39623 42229 39637
rect 42359 39623 42373 39637
rect 45695 39623 45709 39637
rect 45887 39623 45901 39637
rect 47135 39623 47149 39637
rect 28079 39575 28093 39589
rect 31775 39575 31789 39589
rect 42215 39575 42229 39589
rect 42359 39575 42373 39589
rect 45743 39575 45757 39589
rect 45767 39575 45781 39589
rect 47159 39599 47173 39613
rect 47207 39575 47221 39589
rect 28079 39527 28093 39541
rect 31775 39527 31789 39541
rect 45743 39527 45757 39541
rect 46871 39527 46885 39541
rect 47039 39551 47053 39565
rect 47231 39551 47245 39565
rect 47255 39527 47269 39541
rect 38855 39503 38869 39517
rect 47111 39503 47125 39517
rect 47135 39503 47149 39517
rect 27887 39455 27901 39469
rect 28079 39455 28093 39469
rect 31775 39455 31789 39469
rect 38663 39455 38677 39469
rect 39023 39455 39037 39469
rect 47135 39455 47149 39469
rect 47183 39455 47197 39469
rect 21215 39239 21229 39253
rect 21431 39239 21445 39253
rect 21455 39239 21469 39253
rect 21479 39239 21493 39253
rect 21215 39191 21229 39205
rect 20279 38807 20293 38821
rect 21215 38807 21229 38821
rect 21431 39191 21445 39205
rect 22007 39191 22021 39205
rect 20279 38759 20293 38773
rect 21215 38759 21229 38773
rect 20279 34823 20293 34837
rect 20255 34751 20269 34765
rect 20255 34703 20269 34717
rect 20279 34703 20293 34717
rect 20255 30767 20269 30781
rect 20279 30767 20293 30781
rect 20303 30767 20317 30781
rect 21215 30767 21229 30781
rect 47159 39407 47173 39421
rect 47279 39407 47293 39421
rect 47303 39407 47317 39421
rect 47039 39383 47053 39397
rect 47063 39383 47077 39397
rect 47327 39383 47341 39397
rect 26855 39359 26869 39373
rect 36143 39359 36157 39373
rect 36863 39359 36877 39373
rect 47159 39359 47173 39373
rect 47207 39359 47221 39373
rect 47351 39359 47365 39373
rect 46991 39335 47005 39349
rect 47087 39335 47101 39349
rect 47375 39335 47389 39349
rect 26855 39311 26869 39325
rect 27887 39311 27901 39325
rect 28079 39311 28093 39325
rect 31775 39311 31789 39325
rect 47207 39311 47221 39325
rect 47231 39311 47245 39325
rect 47399 39311 47413 39325
rect 47231 39287 47245 39301
rect 47303 39287 47317 39301
rect 47423 39287 47437 39301
rect 26663 39263 26677 39277
rect 26855 39263 26869 39277
rect 27887 39263 27901 39277
rect 28079 39263 28093 39277
rect 31775 39263 31789 39277
rect 35879 39263 35893 39277
rect 38927 39263 38941 39277
rect 42359 39263 42373 39277
rect 45743 39263 45757 39277
rect 45767 39263 45781 39277
rect 47351 39263 47365 39277
rect 47375 39263 47389 39277
rect 47447 39263 47461 39277
rect 47087 39239 47101 39253
rect 47303 39239 47317 39253
rect 26663 39215 26677 39229
rect 26855 39215 26869 39229
rect 27887 39215 27901 39229
rect 28079 39215 28093 39229
rect 31775 39215 31789 39229
rect 42215 39191 42229 39205
rect 46823 39167 46837 39181
rect 46871 39191 46885 39205
rect 21455 39143 21469 39157
rect 21479 39143 21493 39157
rect 22127 39143 22141 39157
rect 25463 39143 25477 39157
rect 25703 39143 25717 39157
rect 26663 39143 26677 39157
rect 26855 39143 26869 39157
rect 27887 39143 27901 39157
rect 46823 39143 46837 39157
rect 46991 39143 47005 39157
rect 47015 39143 47029 39157
rect 47039 39143 47053 39157
rect 47063 39143 47077 39157
rect 47087 39143 47101 39157
rect 47111 39143 47125 39157
rect 47135 39143 47149 39157
rect 47159 39143 47173 39157
rect 47183 39143 47197 39157
rect 47207 39143 47221 39157
rect 47231 39143 47245 39157
rect 47255 39143 47269 39157
rect 47279 39143 47293 39157
rect 47303 39143 47317 39157
rect 47327 39143 47341 39157
rect 20303 30719 20317 30733
rect 21215 30719 21229 30733
rect 20255 30671 20269 30685
rect 20279 30671 20293 30685
rect 20279 26807 20293 26821
rect 20279 26759 20293 26773
rect 20279 22847 20293 22861
rect 20303 22847 20317 22861
rect 20279 22799 20293 22813
rect 20303 22799 20317 22813
rect 20303 19631 20317 19645
rect 21431 19655 21445 19669
rect 21119 19631 21133 19645
rect 21215 19631 21229 19645
rect 21383 19631 21397 19645
rect 47399 39191 47413 39205
rect 47423 39191 47437 39205
rect 47447 39191 47461 39205
rect 46991 36455 47005 36469
rect 47015 36455 47029 36469
rect 47039 36455 47053 36469
rect 47063 36455 47077 36469
rect 47087 36455 47101 36469
rect 47111 36455 47125 36469
rect 47135 36455 47149 36469
rect 47159 36455 47173 36469
rect 47183 36455 47197 36469
rect 47207 36455 47221 36469
rect 47231 36455 47245 36469
rect 47255 36455 47269 36469
rect 47279 36455 47293 36469
rect 47303 36455 47317 36469
rect 47327 36455 47341 36469
rect 47351 36455 47365 36469
rect 47375 36455 47389 36469
rect 47399 36455 47413 36469
rect 47423 36455 47437 36469
rect 47447 36455 47461 36469
rect 50255 38999 50269 39013
rect 50255 38951 50269 38965
rect 47447 36407 47461 36421
rect 46991 36335 47005 36349
rect 47015 36335 47029 36349
rect 47039 36335 47053 36349
rect 47063 36335 47077 36349
rect 47087 36335 47101 36349
rect 47111 36335 47125 36349
rect 47135 36335 47149 36349
rect 47159 36335 47173 36349
rect 47183 36335 47197 36349
rect 47207 36335 47221 36349
rect 47231 36335 47245 36349
rect 47255 36335 47269 36349
rect 47279 36335 47293 36349
rect 47303 36335 47317 36349
rect 47327 36335 47341 36349
rect 47351 36335 47365 36349
rect 47375 36335 47389 36349
rect 47399 36335 47413 36349
rect 47423 36335 47437 36349
rect 46991 35351 47005 35365
rect 47015 35351 47029 35365
rect 47039 35351 47053 35365
rect 47063 35351 47077 35365
rect 47087 35351 47101 35365
rect 47111 35351 47125 35365
rect 47135 35351 47149 35365
rect 47159 35351 47173 35365
rect 47183 35351 47197 35365
rect 47207 35351 47221 35365
rect 47231 35351 47245 35365
rect 47255 35351 47269 35365
rect 47279 35351 47293 35365
rect 47303 35351 47317 35365
rect 47327 35351 47341 35365
rect 47351 35351 47365 35365
rect 47375 35351 47389 35365
rect 47399 35351 47413 35365
rect 47399 35303 47413 35317
rect 46991 35231 47005 35245
rect 47015 35231 47029 35245
rect 47039 35231 47053 35245
rect 47063 35231 47077 35245
rect 47087 35231 47101 35245
rect 47111 35231 47125 35245
rect 47135 35231 47149 35245
rect 47159 35231 47173 35245
rect 47183 35231 47197 35245
rect 47207 35231 47221 35245
rect 47231 35231 47245 35245
rect 47255 35231 47269 35245
rect 47279 35231 47293 35245
rect 47303 35231 47317 35245
rect 47327 35231 47341 35245
rect 47351 35231 47365 35245
rect 47375 35231 47389 35245
rect 46991 34223 47005 34237
rect 47015 34223 47029 34237
rect 47039 34223 47053 34237
rect 47063 34223 47077 34237
rect 47087 34223 47101 34237
rect 47111 34223 47125 34237
rect 47135 34223 47149 34237
rect 47159 34223 47173 34237
rect 47183 34223 47197 34237
rect 47207 34223 47221 34237
rect 47231 34223 47245 34237
rect 47255 34223 47269 34237
rect 47279 34223 47293 34237
rect 47303 34223 47317 34237
rect 47327 34223 47341 34237
rect 47351 34223 47365 34237
rect 50255 38855 50269 38869
rect 50255 38807 50269 38821
rect 50231 34967 50245 34981
rect 50255 34967 50269 34981
rect 50231 34919 50245 34933
rect 50255 34919 50269 34933
rect 50183 34847 50197 34861
rect 50207 34847 50221 34861
rect 47351 34175 47365 34189
rect 46991 34103 47005 34117
rect 47015 34103 47029 34117
rect 47039 34103 47053 34117
rect 47063 34103 47077 34117
rect 47087 34103 47101 34117
rect 47111 34103 47125 34117
rect 47135 34103 47149 34117
rect 47159 34103 47173 34117
rect 47183 34103 47197 34117
rect 47207 34103 47221 34117
rect 47231 34103 47245 34117
rect 47255 34103 47269 34117
rect 47279 34103 47293 34117
rect 47303 34103 47317 34117
rect 47327 34103 47341 34117
rect 46991 33119 47005 33133
rect 47015 33119 47029 33133
rect 47039 33119 47053 33133
rect 47063 33119 47077 33133
rect 47087 33119 47101 33133
rect 47111 33119 47125 33133
rect 47135 33119 47149 33133
rect 47159 33119 47173 33133
rect 47183 33119 47197 33133
rect 47207 33119 47221 33133
rect 47231 33119 47245 33133
rect 47255 33119 47269 33133
rect 47279 33119 47293 33133
rect 47303 33119 47317 33133
rect 47303 33071 47317 33085
rect 46991 32999 47005 33013
rect 47015 32999 47029 33013
rect 47039 32999 47053 33013
rect 47063 32999 47077 33013
rect 47087 32999 47101 33013
rect 47111 32999 47125 33013
rect 47135 32999 47149 33013
rect 47159 32999 47173 33013
rect 47183 32999 47197 33013
rect 47207 32999 47221 33013
rect 47231 32999 47245 33013
rect 47255 32999 47269 33013
rect 47279 32999 47293 33013
rect 46991 32015 47005 32029
rect 47015 32015 47029 32029
rect 47039 32015 47053 32029
rect 47063 32015 47077 32029
rect 47087 32015 47101 32029
rect 47111 32015 47125 32029
rect 47135 32015 47149 32029
rect 47159 32015 47173 32029
rect 47183 32015 47197 32029
rect 47207 32015 47221 32029
rect 47231 32015 47245 32029
rect 47255 32015 47269 32029
rect 47279 32015 47293 32029
rect 50255 34823 50269 34837
rect 50183 34799 50197 34813
rect 50207 34799 50221 34813
rect 46991 31895 47005 31909
rect 47015 31895 47029 31909
rect 47039 31895 47053 31909
rect 47063 31895 47077 31909
rect 47087 31895 47101 31909
rect 47111 31895 47125 31909
rect 47135 31895 47149 31909
rect 47159 31895 47173 31909
rect 47183 31895 47197 31909
rect 47207 31895 47221 31909
rect 47231 31895 47245 31909
rect 47255 31895 47269 31909
rect 47279 31895 47293 31909
rect 50207 30959 50221 30973
rect 50255 34775 50269 34789
rect 46991 30887 47005 30901
rect 47015 30887 47029 30901
rect 47039 30887 47053 30901
rect 47063 30887 47077 30901
rect 47087 30887 47101 30901
rect 47111 30887 47125 30901
rect 47135 30887 47149 30901
rect 47159 30887 47173 30901
rect 47183 30887 47197 30901
rect 47207 30887 47221 30901
rect 47231 30887 47245 30901
rect 47255 30887 47269 30901
rect 47279 30887 47293 30901
rect 50255 30935 50269 30949
rect 50207 30911 50221 30925
rect 50255 30887 50269 30901
rect 46991 30791 47005 30805
rect 47015 30791 47029 30805
rect 47039 30791 47053 30805
rect 47063 30791 47077 30805
rect 47087 30791 47101 30805
rect 47111 30791 47125 30805
rect 47135 30791 47149 30805
rect 47159 30791 47173 30805
rect 47183 30791 47197 30805
rect 47207 30791 47221 30805
rect 47231 30791 47245 30805
rect 47255 30791 47269 30805
rect 47279 30791 47293 30805
rect 50231 30791 50245 30805
rect 50255 30791 50269 30805
rect 46991 29783 47005 29797
rect 47015 29783 47029 29797
rect 47039 29783 47053 29797
rect 47063 29783 47077 29797
rect 47087 29783 47101 29797
rect 47111 29783 47125 29797
rect 47135 29783 47149 29797
rect 47159 29783 47173 29797
rect 47183 29783 47197 29797
rect 47207 29783 47221 29797
rect 47231 29783 47245 29797
rect 47255 29783 47269 29797
rect 47279 29783 47293 29797
rect 50231 30743 50245 30757
rect 50255 30743 50269 30757
rect 46991 29663 47005 29677
rect 47015 29663 47029 29677
rect 47039 29663 47053 29677
rect 47063 29663 47077 29677
rect 47087 29663 47101 29677
rect 47111 29663 47125 29677
rect 47135 29663 47149 29677
rect 47159 29663 47173 29677
rect 47183 29663 47197 29677
rect 47207 29663 47221 29677
rect 47231 29663 47245 29677
rect 47255 29663 47269 29677
rect 47279 29663 47293 29677
rect 46991 28679 47005 28693
rect 47015 28679 47029 28693
rect 47039 28679 47053 28693
rect 47063 28679 47077 28693
rect 47087 28679 47101 28693
rect 47111 28679 47125 28693
rect 47135 28679 47149 28693
rect 47159 28679 47173 28693
rect 47183 28679 47197 28693
rect 47207 28679 47221 28693
rect 47231 28679 47245 28693
rect 47279 28703 47293 28717
rect 47303 28631 47317 28645
rect 46991 28559 47005 28573
rect 47015 28559 47029 28573
rect 47039 28559 47053 28573
rect 47063 28559 47077 28573
rect 47087 28559 47101 28573
rect 47111 28559 47125 28573
rect 47135 28559 47149 28573
rect 47159 28559 47173 28573
rect 47183 28559 47197 28573
rect 47207 28559 47221 28573
rect 47231 28559 47245 28573
rect 46991 27551 47005 27565
rect 47015 27551 47029 27565
rect 47279 28583 47293 28597
rect 47303 28583 47317 28597
rect 47063 27575 47077 27589
rect 47087 27575 47101 27589
rect 47111 27575 47125 27589
rect 47135 27575 47149 27589
rect 47159 27575 47173 27589
rect 47183 27575 47197 27589
rect 47207 27575 47221 27589
rect 47231 27575 47245 27589
rect 47255 27575 47269 27589
rect 47279 27575 47293 27589
rect 47303 27575 47317 27589
rect 47327 27575 47341 27589
rect 47039 27527 47053 27541
rect 47351 27527 47365 27541
rect 47015 27503 47029 27517
rect 46991 27455 47005 27469
rect 47039 27479 47053 27493
rect 47063 27479 47077 27493
rect 47087 27479 47101 27493
rect 47111 27479 47125 27493
rect 47135 27479 47149 27493
rect 47159 27479 47173 27493
rect 47183 27479 47197 27493
rect 47207 27479 47221 27493
rect 47231 27479 47245 27493
rect 47255 27479 47269 27493
rect 47279 27479 47293 27493
rect 47303 27479 47317 27493
rect 47327 27479 47341 27493
rect 47351 27479 47365 27493
rect 46991 26447 47005 26461
rect 47015 26447 47029 26461
rect 47039 26447 47053 26461
rect 50255 26807 50269 26821
rect 50279 26783 50293 26797
rect 50255 26759 50269 26773
rect 47087 26471 47101 26485
rect 47111 26471 47125 26485
rect 47135 26471 47149 26485
rect 47159 26471 47173 26485
rect 47183 26471 47197 26485
rect 47207 26471 47221 26485
rect 47231 26471 47245 26485
rect 47255 26471 47269 26485
rect 47279 26471 47293 26485
rect 47303 26471 47317 26485
rect 47327 26471 47341 26485
rect 47351 26471 47365 26485
rect 46991 26399 47005 26413
rect 47063 26399 47077 26413
rect 47375 26399 47389 26413
rect 47015 26351 47029 26365
rect 47039 26351 47053 26365
rect 47063 26351 47077 26365
rect 47087 26351 47101 26365
rect 47111 26351 47125 26365
rect 47135 26351 47149 26365
rect 47159 26351 47173 26365
rect 47183 26351 47197 26365
rect 47207 26351 47221 26365
rect 47231 26351 47245 26365
rect 47255 26351 47269 26365
rect 47279 26351 47293 26365
rect 47303 26351 47317 26365
rect 47327 26351 47341 26365
rect 47351 26351 47365 26365
rect 47375 26351 47389 26365
rect 46991 25343 47005 25357
rect 47015 25343 47029 25357
rect 47039 25343 47053 25357
rect 47063 25343 47077 25357
rect 47087 25343 47101 25357
rect 47135 25367 47149 25381
rect 47159 25367 47173 25381
rect 47183 25367 47197 25381
rect 47207 25367 47221 25381
rect 47231 25367 47245 25381
rect 47255 25367 47269 25381
rect 47279 25367 47293 25381
rect 47303 25367 47317 25381
rect 47327 25367 47341 25381
rect 47351 25367 47365 25381
rect 47375 25367 47389 25381
rect 47399 25367 47413 25381
rect 47135 25319 47149 25333
rect 47159 25319 47173 25333
rect 47183 25319 47197 25333
rect 47207 25319 47221 25333
rect 47231 25319 47245 25333
rect 47111 25271 47125 25285
rect 47135 25271 47149 25285
rect 47159 25271 47173 25285
rect 47183 25271 47197 25285
rect 47207 25271 47221 25285
rect 47423 25295 47437 25309
rect 46991 25223 47005 25237
rect 47015 25223 47029 25237
rect 47039 25223 47053 25237
rect 47063 25223 47077 25237
rect 47087 25223 47101 25237
rect 47111 25223 47125 25237
rect 47135 25223 47149 25237
rect 47159 25223 47173 25237
rect 47183 25223 47197 25237
rect 47207 25223 47221 25237
rect 47255 25247 47269 25261
rect 47279 25247 47293 25261
rect 47303 25247 47317 25261
rect 47327 25247 47341 25261
rect 47351 25247 47365 25261
rect 47375 25247 47389 25261
rect 47399 25247 47413 25261
rect 47423 25247 47437 25261
rect 46991 24239 47005 24253
rect 47015 24239 47029 24253
rect 47039 24239 47053 24253
rect 47063 24239 47077 24253
rect 47087 24239 47101 24253
rect 47111 24239 47125 24253
rect 47135 24239 47149 24253
rect 47159 24239 47173 24253
rect 47183 24239 47197 24253
rect 47207 24239 47221 24253
rect 47231 24239 47245 24253
rect 47279 24263 47293 24277
rect 47303 24263 47317 24277
rect 47327 24263 47341 24277
rect 47351 24263 47365 24277
rect 47375 24263 47389 24277
rect 47399 24263 47413 24277
rect 47423 24263 47437 24277
rect 47447 24263 47461 24277
rect 47135 24191 47149 24205
rect 47255 24191 47269 24205
rect 47471 24191 47485 24205
rect 46991 24119 47005 24133
rect 47015 24119 47029 24133
rect 47039 24119 47053 24133
rect 47063 24119 47077 24133
rect 47087 24119 47101 24133
rect 47111 24119 47125 24133
rect 46991 23111 47005 23125
rect 47015 23111 47029 23125
rect 47039 23111 47053 23125
rect 47063 23111 47077 23125
rect 47159 24143 47173 24157
rect 47183 24143 47197 24157
rect 47207 24143 47221 24157
rect 47231 24143 47245 24157
rect 47255 24143 47269 24157
rect 47279 24143 47293 24157
rect 47303 24143 47317 24157
rect 47327 24143 47341 24157
rect 47351 24143 47365 24157
rect 47375 24143 47389 24157
rect 47399 24143 47413 24157
rect 47423 24143 47437 24157
rect 47447 24143 47461 24157
rect 47471 24143 47485 24157
rect 47111 23135 47125 23149
rect 47135 23135 47149 23149
rect 47159 23135 47173 23149
rect 47183 23135 47197 23149
rect 47207 23135 47221 23149
rect 47231 23135 47245 23149
rect 47255 23135 47269 23149
rect 47279 23135 47293 23149
rect 47303 23135 47317 23149
rect 47327 23135 47341 23149
rect 47351 23135 47365 23149
rect 47375 23135 47389 23149
rect 47399 23135 47413 23149
rect 47423 23135 47437 23149
rect 47447 23135 47461 23149
rect 47471 23135 47485 23149
rect 47495 23135 47509 23149
rect 47375 23087 47389 23101
rect 47519 23087 47533 23101
rect 47087 23063 47101 23077
rect 46991 23015 47005 23029
rect 47015 23015 47029 23029
rect 47039 23015 47053 23029
rect 47063 23015 47077 23029
rect 47087 23015 47101 23029
rect 47111 23015 47125 23029
rect 47135 23015 47149 23029
rect 47159 23015 47173 23029
rect 47183 23015 47197 23029
rect 47207 23015 47221 23029
rect 47231 23015 47245 23029
rect 47255 23015 47269 23029
rect 47279 23015 47293 23029
rect 47303 23015 47317 23029
rect 47327 23015 47341 23029
rect 47351 23015 47365 23029
rect 46991 22007 47005 22021
rect 47015 22007 47029 22021
rect 47039 22007 47053 22021
rect 47063 22007 47077 22021
rect 47087 22007 47101 22021
rect 47111 22007 47125 22021
rect 47135 22007 47149 22021
rect 47159 22007 47173 22021
rect 47183 22007 47197 22021
rect 47207 22007 47221 22021
rect 47399 23039 47413 23053
rect 47423 23039 47437 23053
rect 47447 23039 47461 23053
rect 47471 23039 47485 23053
rect 47495 23039 47509 23053
rect 47519 23039 47533 23053
rect 47255 22031 47269 22045
rect 47279 22031 47293 22045
rect 47303 22031 47317 22045
rect 47327 22031 47341 22045
rect 47351 22031 47365 22045
rect 47375 22031 47389 22045
rect 47399 22031 47413 22045
rect 47423 22031 47437 22045
rect 47447 22031 47461 22045
rect 47471 22031 47485 22045
rect 47495 22031 47509 22045
rect 47519 22031 47533 22045
rect 47543 22031 47557 22045
rect 47159 21959 47173 21973
rect 47231 21959 47245 21973
rect 47567 21959 47581 21973
rect 46991 21887 47005 21901
rect 47015 21887 47029 21901
rect 47039 21887 47053 21901
rect 47063 21887 47077 21901
rect 47087 21887 47101 21901
rect 47111 21887 47125 21901
rect 47135 21887 47149 21901
rect 47183 21911 47197 21925
rect 47207 21911 47221 21925
rect 47231 21911 47245 21925
rect 47255 21911 47269 21925
rect 47279 21911 47293 21925
rect 47303 21911 47317 21925
rect 47327 21911 47341 21925
rect 47351 21911 47365 21925
rect 47375 21911 47389 21925
rect 47399 21911 47413 21925
rect 47423 21911 47437 21925
rect 47447 21911 47461 21925
rect 47471 21911 47485 21925
rect 47495 21911 47509 21925
rect 47519 21911 47533 21925
rect 47543 21911 47557 21925
rect 47567 21911 47581 21925
rect 46991 20903 47005 20917
rect 47015 20903 47029 20917
rect 47039 20903 47053 20917
rect 47063 20903 47077 20917
rect 47087 20903 47101 20917
rect 47111 20903 47125 20917
rect 47135 20903 47149 20917
rect 47159 20903 47173 20917
rect 47183 20903 47197 20917
rect 47207 20903 47221 20917
rect 47231 20903 47245 20917
rect 47255 20903 47269 20917
rect 47279 20903 47293 20917
rect 47303 20903 47317 20917
rect 47327 20903 47341 20917
rect 47351 20903 47365 20917
rect 47375 20903 47389 20917
rect 47399 20903 47413 20917
rect 47423 20903 47437 20917
rect 47447 20903 47461 20917
rect 47471 20903 47485 20917
rect 47495 20903 47509 20917
rect 47519 20903 47533 20917
rect 47543 20903 47557 20917
rect 47591 20927 47605 20941
rect 47207 20855 47221 20869
rect 47567 20855 47581 20869
rect 47615 20855 47629 20869
rect 46991 20783 47005 20797
rect 47015 20783 47029 20797
rect 47039 20783 47053 20797
rect 47063 20783 47077 20797
rect 47087 20783 47101 20797
rect 47111 20783 47125 20797
rect 47135 20783 47149 20797
rect 47159 20783 47173 20797
rect 47183 20783 47197 20797
rect 47231 20807 47245 20821
rect 47255 20807 47269 20821
rect 47279 20807 47293 20821
rect 47303 20807 47317 20821
rect 47327 20807 47341 20821
rect 47351 20807 47365 20821
rect 47375 20807 47389 20821
rect 47399 20807 47413 20821
rect 47423 20807 47437 20821
rect 47447 20807 47461 20821
rect 47471 20807 47485 20821
rect 47495 20807 47509 20821
rect 47519 20807 47533 20821
rect 47543 20807 47557 20821
rect 47567 20807 47581 20821
rect 47591 20807 47605 20821
rect 47615 20807 47629 20821
rect 46991 19775 47005 19789
rect 47015 19775 47029 19789
rect 47039 19775 47053 19789
rect 47063 19775 47077 19789
rect 47087 19775 47101 19789
rect 47111 19775 47125 19789
rect 47135 19775 47149 19789
rect 47159 19775 47173 19789
rect 47183 19775 47197 19789
rect 47207 19775 47221 19789
rect 47231 19775 47245 19789
rect 47279 19799 47293 19813
rect 47303 19799 47317 19813
rect 47327 19799 47341 19813
rect 47351 19799 47365 19813
rect 47375 19799 47389 19813
rect 47399 19799 47413 19813
rect 47423 19799 47437 19813
rect 47447 19799 47461 19813
rect 47471 19799 47485 19813
rect 47495 19799 47509 19813
rect 47519 19799 47533 19813
rect 47543 19799 47557 19813
rect 47567 19799 47581 19813
rect 47591 19799 47605 19813
rect 47615 19799 47629 19813
rect 47639 19799 47653 19813
rect 47255 19751 47269 19765
rect 47663 19751 47677 19765
rect 47231 19727 47245 19741
rect 46991 19679 47005 19693
rect 47015 19679 47029 19693
rect 47039 19679 47053 19693
rect 47063 19679 47077 19693
rect 47087 19679 47101 19693
rect 47111 19679 47125 19693
rect 47135 19679 47149 19693
rect 47159 19679 47173 19693
rect 47183 19679 47197 19693
rect 47207 19679 47221 19693
rect 20303 19583 20317 19597
rect 21119 19583 21133 19597
rect 21215 19583 21229 19597
rect 21383 19583 21397 19597
rect 21431 19583 21445 19597
rect 20255 18791 20269 18805
rect 20255 18743 20269 18757
rect 21581 19607 21595 19621
rect 22007 19607 22021 19621
rect 23447 19607 23461 19621
rect 24239 19607 24253 19621
rect 24791 19607 24805 19621
rect 25007 19607 25021 19621
rect 25751 19607 25765 19621
rect 25919 19607 25933 19621
rect 26303 19607 26317 19621
rect 26495 19607 26509 19621
rect 26711 19607 26725 19621
rect 27455 19607 27469 19621
rect 27623 19607 27637 19621
rect 46127 19607 46141 19621
rect 46271 19607 46285 19621
rect 46367 19607 46381 19621
rect 46415 19607 46429 19621
rect 46991 19607 47005 19621
rect 47015 19607 47029 19621
rect 47039 19607 47053 19621
rect 47255 19703 47269 19717
rect 47279 19703 47293 19717
rect 47303 19703 47317 19717
rect 47327 19703 47341 19717
rect 47351 19703 47365 19717
rect 47375 19703 47389 19717
rect 47399 19703 47413 19717
rect 47423 19703 47437 19717
rect 47447 19703 47461 19717
rect 47471 19703 47485 19717
rect 47495 19703 47509 19717
rect 47519 19703 47533 19717
rect 47543 19703 47557 19717
rect 47567 19703 47581 19717
rect 47591 19703 47605 19717
rect 47615 19703 47629 19717
rect 47639 19703 47653 19717
rect 47663 19703 47677 19717
rect 47087 19631 47101 19645
rect 47111 19631 47125 19645
rect 47135 19631 47149 19645
rect 47159 19631 47173 19645
rect 47183 19631 47197 19645
rect 47207 19631 47221 19645
rect 47231 19631 47245 19645
rect 47255 19631 47269 19645
rect 47279 19631 47293 19645
rect 47303 19631 47317 19645
rect 47327 19631 47341 19645
rect 47351 19631 47365 19645
rect 47375 19631 47389 19645
rect 47399 19631 47413 19645
rect 47423 19631 47437 19645
rect 47447 19631 47461 19645
rect 47471 19631 47485 19645
rect 47495 19631 47509 19645
rect 47519 19631 47533 19645
rect 47543 19631 47557 19645
rect 47567 19631 47581 19645
rect 47591 19631 47605 19645
rect 47615 19631 47629 19645
rect 47639 19631 47653 19645
rect 47663 19631 47677 19645
rect 47687 19631 47701 19645
rect 21650 19559 21664 19573
rect 21751 19559 21765 19573
rect 21215 19511 21229 19525
rect 21383 19511 21397 19525
rect 21431 19511 21445 19525
rect 21479 19511 21493 19525
rect 21775 19511 21789 19525
rect 21215 19463 21229 19477
rect 21383 19463 21397 19477
rect 21431 19463 21445 19477
rect 21479 19463 21493 19477
rect 21535 19463 21549 19477
rect 21603 19463 21617 19477
rect 21627 19463 21641 19477
rect 21679 19463 21693 19477
rect 21703 19463 21717 19477
rect 21558 19424 21572 19438
rect 21671 18647 21685 18661
rect 21624 18576 21638 18590
rect 21671 18599 21685 18613
rect 21751 19463 21765 19477
rect 21775 19463 21789 19477
rect 21749 18599 21763 18613
rect 21773 18599 21787 18613
rect 22007 18599 22021 18613
rect 23447 18599 23461 18613
rect 24239 18599 24253 18613
rect 24791 18599 24805 18613
rect 25007 18599 25021 18613
rect 25751 18599 25765 18613
rect 26783 18671 26797 18685
rect 27623 18695 27637 18709
rect 27671 18671 27685 18685
rect 29327 18647 29341 18661
rect 37031 19559 37045 19573
rect 37223 19559 37237 19573
rect 37463 19559 37477 19573
rect 30191 18623 30205 18637
rect 31007 18623 31021 18637
rect 45167 19559 45181 19573
rect 45191 19559 45205 19573
rect 46295 19583 46309 19597
rect 45911 19535 45925 19549
rect 45191 19511 45205 19525
rect 46319 19559 46333 19573
rect 46487 19559 46501 19573
rect 47063 19559 47077 19573
rect 47711 19559 47725 19573
rect 46295 19535 46309 19549
rect 46823 19511 46837 19525
rect 46991 19463 47005 19477
rect 47015 19463 47029 19477
rect 47039 19463 47053 19477
rect 47063 19463 47077 19477
rect 47087 19463 47101 19477
rect 47111 19463 47125 19477
rect 47135 19463 47149 19477
rect 47159 19463 47173 19477
rect 47183 19463 47197 19477
rect 47207 19463 47221 19477
rect 47231 19463 47245 19477
rect 47255 19463 47269 19477
rect 47279 19463 47293 19477
rect 47303 19463 47317 19477
rect 47327 19463 47341 19477
rect 47351 19463 47365 19477
rect 47375 19463 47389 19477
rect 47399 19463 47413 19477
rect 47423 19463 47437 19477
rect 47447 19463 47461 19477
rect 47471 19463 47485 19477
rect 47495 19463 47509 19477
rect 47519 19463 47533 19477
rect 47543 19463 47557 19477
rect 47567 19463 47581 19477
rect 47591 19463 47605 19477
rect 47615 19463 47629 19477
rect 47639 19463 47653 19477
rect 47663 19463 47677 19477
rect 47687 19463 47701 19477
rect 47711 19463 47725 19477
rect 31895 18599 31909 18613
rect 37031 18599 37045 18613
rect 37223 18599 37237 18613
rect 37463 18599 37477 18613
rect 42863 18599 42877 18613
rect 43703 18599 43717 18613
rect 44543 18599 44557 18613
rect 46204 18599 46218 18613
rect 46228 18599 46242 18613
rect 46991 18599 47005 18613
rect 47015 18599 47029 18613
rect 47039 18599 47053 18613
rect 47063 18599 47077 18613
rect 47087 18599 47101 18613
rect 47111 18599 47125 18613
rect 47135 18599 47149 18613
rect 47159 18599 47173 18613
rect 47183 18599 47197 18613
rect 47207 18599 47221 18613
rect 47231 18599 47245 18613
rect 47903 19055 47917 19069
rect 49127 19031 49141 19045
rect 49415 19007 49429 19021
rect 49439 18983 49453 18997
rect 49463 18959 49477 18973
rect 49487 18935 49501 18949
rect 49511 18911 49525 18925
rect 49535 18887 49549 18901
rect 49559 18863 49573 18877
rect 49583 18839 49597 18853
rect 49607 18815 49621 18829
rect 49631 18791 49645 18805
rect 50255 18791 50269 18805
rect 49655 18743 49669 18757
rect 50255 18743 50269 18757
rect 49679 18719 49693 18733
rect 49703 18695 49717 18709
rect 49727 18671 49741 18685
rect 49751 18647 49765 18661
rect 50255 18647 50269 18661
rect 49775 18599 49789 18613
rect 50255 18599 50269 18613
rect 49799 18575 49813 18589
rect 21647 18551 21661 18565
rect 21671 18551 21685 18565
rect 21695 18551 21709 18565
rect 21719 18551 21733 18565
rect 21773 18551 21787 18565
rect 22223 18551 22237 18565
rect 23447 18551 23461 18565
rect 24239 18551 24253 18565
rect 24791 18551 24805 18565
rect 25007 18551 25021 18565
rect 25103 18551 25117 18565
rect 25751 18551 25765 18565
rect 32735 18551 32749 18565
rect 37031 18551 37045 18565
rect 37223 18551 37237 18565
rect 37463 18551 37477 18565
rect 42863 18551 42877 18565
rect 43703 18551 43717 18565
rect 44543 18551 44557 18565
rect 46204 18551 46218 18565
rect 46228 18551 46242 18565
rect 46991 18551 47005 18565
rect 47015 18551 47029 18565
rect 47039 18551 47053 18565
rect 47063 18551 47077 18565
rect 47087 18551 47101 18565
rect 47111 18551 47125 18565
rect 47135 18551 47149 18565
rect 47159 18551 47173 18565
rect 47183 18551 47197 18565
rect 47207 18551 47221 18565
rect 47231 18551 47245 18565
rect 49823 18551 49837 18565
rect 22247 18527 22261 18541
rect 24215 18527 24229 18541
rect 24263 18527 24277 18541
rect 33575 18527 33589 18541
rect 21559 18503 21573 18517
rect 21749 18503 21763 18517
rect 25079 18503 25093 18517
rect 25103 18503 25117 18517
rect 33599 18503 33613 18517
rect 24191 18479 24205 18493
rect 24215 18479 24229 18493
rect 31871 18479 31885 18493
rect 31895 18479 31909 18493
rect 35303 18479 35317 18493
rect 21559 18455 21573 18469
rect 21623 18455 21637 18469
rect 21671 18455 21685 18469
rect 29303 18455 29317 18469
rect 29327 18455 29341 18469
rect 36124 18455 36138 18469
rect 21671 18431 21685 18445
rect 22168 18431 22182 18445
rect 22247 18431 22261 18445
rect 26759 18431 26773 18445
rect 26783 18431 26797 18445
rect 36172 18431 36186 18445
rect 37823 18479 37837 18493
rect 38495 18455 38509 18469
rect 39431 18431 39445 18445
rect 27599 18407 27613 18421
rect 27623 18407 27637 18421
rect 40319 18407 40333 18421
rect 20303 18383 20317 18397
rect 21215 18383 21229 18397
rect 21383 18383 21397 18397
rect 21431 18383 21445 18397
rect 21479 18383 21493 18397
rect 21559 18383 21573 18397
rect 21647 18383 21661 18397
rect 30167 18383 30181 18397
rect 30191 18383 30205 18397
rect 36148 18383 36162 18397
rect 36172 18383 36186 18397
rect 38471 18383 38485 18397
rect 38495 18383 38509 18397
rect 22144 18359 22158 18373
rect 22223 18359 22237 18373
rect 27647 18359 27661 18373
rect 27671 18359 27685 18373
rect 39407 18359 39421 18373
rect 39431 18359 39445 18373
rect 41039 18359 41053 18373
rect 20303 18335 20317 18349
rect 21215 18335 21229 18349
rect 21383 18335 21397 18349
rect 21431 18335 21445 18349
rect 21479 18335 21493 18349
rect 21559 18335 21573 18349
rect 24263 18335 24277 18349
rect 32735 18335 32749 18349
rect 35303 18335 35317 18349
rect 37823 18335 37837 18349
rect 47063 18407 47077 18421
rect 49847 18527 49861 18541
rect 49871 18527 49885 18541
rect 49895 18503 49909 18517
rect 49919 18479 49933 18493
rect 49943 18455 49957 18469
rect 49991 18431 50005 18445
rect 50039 18407 50053 18421
rect 50159 18383 50173 18397
rect 50207 18359 50221 18373
rect 21671 18311 21685 18325
rect 21695 18311 21709 18325
rect 21719 18311 21733 18325
rect 24239 18311 24253 18325
rect 32711 18311 32725 18325
rect 35279 18311 35293 18325
rect 37799 18311 37813 18325
rect 41543 18311 41557 18325
rect 42023 18311 42037 18325
rect 42863 18311 42877 18325
rect 43703 18311 43717 18325
rect 44543 18311 44557 18325
rect 46204 18311 46218 18325
rect 46228 18311 46242 18325
rect 49415 18311 49429 18325
rect 49439 18311 49453 18325
rect 49463 18311 49477 18325
rect 49487 18311 49501 18325
rect 49511 18311 49525 18325
rect 49535 18311 49549 18325
rect 49559 18311 49573 18325
rect 49583 18311 49597 18325
rect 49607 18311 49621 18325
rect 49631 18311 49645 18325
rect 49655 18311 49669 18325
rect 49679 18311 49693 18325
rect 49703 18311 49717 18325
rect 49727 18311 49741 18325
rect 49751 18311 49765 18325
rect 49775 18311 49789 18325
rect 49799 18311 49813 18325
rect 49823 18311 49837 18325
rect 49847 18311 49861 18325
rect 49871 18311 49885 18325
rect 49895 18311 49909 18325
rect 49919 18311 49933 18325
rect 49943 18311 49957 18325
rect 49991 18311 50005 18325
rect 50039 18311 50053 18325
rect 50159 18311 50173 18325
rect 50207 18311 50221 18325
rect 21431 18239 21445 18253
rect 21479 18239 21493 18253
rect 21671 18239 21685 18253
rect 21695 18239 21709 18253
rect 21719 18239 21733 18253
rect 21743 18210 21757 18224
rect 21431 18186 21445 18200
rect 21743 18186 21757 18200
rect 21479 18162 21493 18176
rect 21671 18162 21685 18176
rect 21695 18162 21709 18176
rect 21719 18162 21733 18176
rect 20255 14735 20269 14749
rect 20303 14735 20317 14749
rect 21215 14735 21229 14749
rect 21479 14735 21493 14749
rect 20255 14687 20269 14701
rect 20303 14687 20317 14701
rect 21215 14687 21229 14701
rect 21479 14687 21493 14701
rect 20255 10703 20269 10717
rect 20255 10655 20269 10669
rect 49511 18186 49525 18200
rect 49535 18186 49549 18200
rect 49559 18186 49573 18200
rect 49583 18186 49597 18200
rect 49607 18186 49621 18200
rect 49631 18186 49645 18200
rect 49655 18186 49669 18200
rect 49679 18186 49693 18200
rect 49703 18186 49717 18200
rect 49727 18186 49741 18200
rect 49751 18186 49765 18200
rect 49775 18186 49789 18200
rect 49799 18186 49813 18200
rect 49823 18186 49837 18200
rect 49847 18186 49861 18200
rect 49871 18186 49885 18200
rect 49895 18186 49909 18200
rect 49919 18186 49933 18200
rect 49943 18186 49957 18200
rect 49415 18138 49429 18152
rect 49439 18138 49453 18152
rect 49463 18138 49477 18152
rect 49871 18138 49885 18152
rect 49391 18114 49405 18128
rect 49487 18114 49501 18128
rect 49391 18090 49405 18104
rect 49895 18090 49909 18104
rect 49919 18090 49933 18104
rect 49943 18090 49957 18104
rect 49391 18066 49405 18080
rect 49751 18066 49765 18080
rect 49775 18066 49789 18080
rect 49799 18066 49813 18080
rect 49823 18066 49837 18080
rect 49847 18066 49861 18080
rect 49391 18042 49405 18056
rect 49391 18018 49405 18032
rect 49583 18018 49597 18032
rect 49607 18018 49621 18032
rect 49631 18018 49645 18032
rect 49655 18018 49669 18032
rect 49679 18018 49693 18032
rect 49703 18018 49717 18032
rect 49727 18018 49741 18032
rect 49415 17994 49429 18008
rect 49439 17994 49453 18008
rect 49463 17994 49477 18008
rect 49487 17994 49501 18008
rect 49511 17994 49525 18008
rect 49535 17994 49549 18008
rect 49559 17994 49573 18008
rect 49415 17087 49429 17101
rect 49439 17087 49453 17101
rect 49463 17087 49477 17101
rect 49487 17087 49501 17101
rect 49511 17087 49525 17101
rect 49535 17087 49549 17101
rect 49559 17087 49573 17101
rect 49607 17087 49621 17101
rect 49631 17087 49645 17101
rect 49655 17087 49669 17101
rect 49679 17087 49693 17101
rect 49391 17063 49405 17077
rect 49415 17039 49429 17053
rect 49439 17039 49453 17053
rect 49463 17039 49477 17053
rect 49487 17039 49501 17053
rect 49511 17039 49525 17053
rect 49535 17039 49549 17053
rect 49559 17039 49573 17053
rect 49607 17039 49621 17053
rect 49631 17039 49645 17053
rect 49655 17039 49669 17053
rect 49679 17039 49693 17053
rect 21479 14137 21493 14151
rect 21695 14137 21709 14151
rect 21719 14137 21733 14151
rect 21743 14113 21757 14127
rect 21479 14089 21493 14103
rect 21743 14089 21757 14103
rect 21695 14063 21709 14077
rect 21719 14063 21733 14077
rect 49511 14807 49525 14821
rect 49535 14807 49549 14821
rect 49559 14807 49573 14821
rect 49607 14807 49621 14821
rect 49631 14807 49645 14821
rect 49655 14807 49669 14821
rect 49679 14807 49693 14821
rect 49727 14807 49741 14821
rect 49799 14807 49813 14821
rect 49823 14807 49837 14821
rect 49847 14807 49861 14821
rect 49895 14807 49909 14821
rect 49919 14807 49933 14821
rect 49943 14807 49957 14821
rect 49991 14807 50005 14821
rect 50039 14807 50053 14821
rect 50159 14807 50173 14821
rect 50207 14807 50221 14821
rect 50231 14807 50245 14821
rect 49511 14759 49525 14773
rect 49535 14759 49549 14773
rect 49559 14759 49573 14773
rect 49607 14759 49621 14773
rect 49631 14759 49645 14773
rect 49655 14759 49669 14773
rect 49679 14759 49693 14773
rect 49727 14759 49741 14773
rect 49799 14759 49813 14773
rect 49823 14759 49837 14773
rect 49847 14759 49861 14773
rect 49895 14759 49909 14773
rect 49919 14759 49933 14773
rect 49943 14759 49957 14773
rect 49991 14759 50005 14773
rect 50039 14759 50053 14773
rect 50159 14759 50173 14773
rect 50255 14759 50269 14773
rect 49415 13271 49429 13285
rect 49439 13271 49453 13285
rect 49463 13271 49477 13285
rect 49511 13271 49525 13285
rect 49535 13271 49549 13285
rect 49559 13271 49573 13285
rect 49391 13247 49405 13261
rect 49415 13223 49429 13237
rect 49439 13223 49453 13237
rect 49463 13223 49477 13237
rect 49511 13223 49525 13237
rect 49535 13223 49549 13237
rect 49559 13223 49573 13237
rect 49415 11905 49429 11919
rect 49439 11905 49453 11919
rect 49463 11905 49477 11919
rect 49511 11905 49525 11919
rect 49535 11905 49549 11919
rect 49559 11905 49573 11919
rect 49631 11905 49645 11919
rect 49655 11905 49669 11919
rect 49679 11905 49693 11919
rect 49727 11905 49741 11919
rect 49391 11881 49405 11895
rect 49391 11857 49405 11871
rect 49655 11857 49669 11871
rect 49679 11857 49693 11871
rect 49727 11857 49741 11871
rect 49415 11833 49429 11847
rect 49439 11833 49453 11847
rect 49463 11833 49477 11847
rect 49511 11833 49525 11847
rect 49535 11833 49549 11847
rect 49559 11833 49573 11847
rect 49631 11833 49645 11847
rect 49415 10735 49429 10749
rect 49439 10735 49453 10749
rect 49463 10735 49477 10749
rect 49511 10735 49525 10749
rect 49535 10735 49549 10749
rect 49559 10735 49573 10749
rect 49631 10735 49645 10749
rect 49679 10735 49693 10749
rect 49727 10735 49741 10749
rect 49823 10735 49837 10749
rect 49847 10735 49861 10749
rect 49391 10711 49405 10725
rect 49391 10687 49405 10701
rect 49679 10687 49693 10701
rect 49727 10687 49741 10701
rect 49823 10687 49837 10701
rect 49847 10687 49861 10701
rect 49415 10663 49429 10677
rect 49439 10663 49453 10677
rect 49463 10663 49477 10677
rect 49511 10663 49525 10677
rect 49535 10663 49549 10677
rect 49559 10663 49573 10677
rect 49631 10663 49645 10677
rect 50207 14735 50221 14749
rect 50231 14711 50245 14725
rect 50255 14711 50269 14725
rect 50231 14615 50245 14629
rect 50255 14615 50269 14629
rect 50231 14567 50245 14581
rect 50255 14567 50269 14581
rect 50255 10703 50269 10717
rect 50255 10655 50269 10669
rect 49439 10559 49453 10573
rect 49463 10559 49477 10573
rect 49511 10559 49525 10573
rect 49535 10559 49549 10573
rect 49559 10559 49573 10573
rect 49631 10559 49645 10573
rect 49727 10559 49741 10573
rect 49823 10559 49837 10573
rect 49847 10559 49861 10573
rect 49919 10559 49933 10573
rect 49943 10559 49957 10573
rect 49991 10559 50005 10573
rect 50039 10559 50053 10573
rect 50255 10559 50269 10573
rect 49439 10511 49453 10525
rect 49463 10511 49477 10525
rect 49511 10511 49525 10525
rect 49535 10511 49549 10525
rect 49559 10511 49573 10525
rect 49631 10511 49645 10525
rect 49727 10511 49741 10525
rect 49823 10511 49837 10525
rect 49847 10511 49861 10525
rect 49919 10511 49933 10525
rect 49943 10511 49957 10525
rect 49991 10511 50005 10525
rect 50039 10511 50053 10525
rect 50255 10511 50269 10525
rect 21695 10400 21709 10414
rect 21719 10400 21733 10414
rect 21743 10376 21757 10390
rect 21743 10352 21757 10366
rect 49439 10351 49453 10365
rect 49463 10351 49477 10365
rect 49511 10351 49525 10365
rect 49535 10351 49549 10365
rect 49559 10351 49573 10365
rect 21695 10319 21709 10333
rect 21719 10319 21733 10333
rect 49391 10327 49405 10341
rect 49391 10303 49405 10317
rect 49535 10303 49549 10317
rect 49559 10303 49573 10317
rect 49463 10279 49477 10293
rect 49511 10279 49525 10293
rect 21671 10247 21685 10261
rect 21695 10247 21709 10261
rect 21719 10247 21733 10261
rect 22199 10247 22213 10261
rect 22127 10199 22141 10213
rect 21671 10151 21685 10165
rect 21695 10151 21709 10165
rect 21719 10151 21733 10165
rect 29735 10223 29749 10237
rect 29759 10223 29773 10237
rect 32903 10223 32917 10237
rect 32927 10223 32941 10237
rect 39215 10223 39229 10237
rect 39239 10223 39253 10237
rect 45935 10223 45949 10237
rect 45959 10223 45973 10237
rect 49511 10223 49525 10237
rect 29759 10175 29773 10189
rect 32927 10175 32941 10189
rect 38855 10175 38869 10189
rect 39239 10175 39253 10189
rect 42239 10175 42253 10189
rect 45959 10175 45973 10189
rect 45983 10175 45997 10189
rect 49511 10175 49525 10189
rect 49727 10175 49741 10189
rect 49823 10175 49837 10189
rect 29735 10151 29749 10165
rect 31799 10151 31813 10165
rect 32903 10151 32917 10165
rect 49439 10127 49453 10141
rect 31799 10103 31813 10117
rect 38855 10103 38869 10117
rect 39215 10103 39229 10117
rect 45983 10079 45997 10093
rect 31655 10055 31669 10069
rect 31799 10055 31813 10069
rect 38855 10055 38869 10069
rect 45911 10055 45925 10069
rect 45935 10055 45949 10069
rect 46727 10079 46741 10093
rect 49727 10079 49741 10093
rect 49823 10079 49837 10093
rect 31655 10007 31669 10021
rect 31799 10007 31813 10021
rect 38855 10007 38869 10021
rect 42239 10007 42253 10021
rect 45911 10007 45925 10021
rect 45911 9935 45925 9949
rect 49943 9935 49957 9949
rect 45767 9887 45781 9901
rect 38855 9863 38869 9877
rect 42239 9863 42253 9877
rect 42383 9863 42397 9877
rect 46007 9887 46021 9901
rect 50039 9887 50053 9901
rect 45983 9863 45997 9877
rect 28127 9839 28141 9853
rect 28271 9839 28285 9853
rect 31655 9839 31669 9853
rect 31799 9839 31813 9853
rect 38711 9839 38725 9853
rect 50039 9839 50053 9853
rect 28127 9791 28141 9805
rect 28271 9791 28285 9805
rect 31655 9791 31669 9805
rect 31799 9791 31813 9805
rect 38711 9791 38725 9805
rect 38855 9791 38869 9805
rect 42239 9791 42253 9805
rect 42383 9791 42397 9805
rect 45767 9791 45781 9805
rect 45911 9791 45925 9805
rect 45983 9815 45997 9829
rect 46007 9815 46021 9829
rect 49943 9815 49957 9829
<< metal2 >>
rect 24552 39709 24564 39743
rect 21456 39637 21468 39671
rect 21480 39637 21492 39671
rect 21504 39661 21516 39695
rect 24624 39685 24636 39719
rect 28080 39709 28092 39743
rect 31632 39709 31644 39743
rect 31776 39685 31788 39743
rect 38688 39685 38700 39743
rect 38832 39661 38844 39743
rect 42216 39637 42228 39743
rect 42360 39637 42372 39743
rect 45696 39637 45708 39719
rect 45744 39589 45756 39743
rect 45888 39637 45900 39743
rect 28080 39541 28092 39575
rect 31776 39541 31788 39575
rect 26856 39325 26868 39359
rect 27888 39325 27900 39455
rect 28080 39325 28092 39455
rect 31776 39325 31788 39455
rect 21216 39205 21228 39239
rect 21432 39205 21444 39239
rect 21456 39157 21468 39239
rect 21480 39157 21492 39239
rect 26664 39229 26676 39263
rect 26856 39229 26868 39263
rect 27888 39229 27900 39263
rect 28080 39229 28092 39263
rect 31776 39229 31788 39263
rect 22008 39133 22020 39191
rect 22121 39143 22127 39157
rect 25457 39143 25463 39157
rect 25697 39143 25703 39157
rect 26657 39143 26663 39157
rect 26849 39143 26855 39157
rect 27883 39143 27887 39157
rect 35880 39156 35892 39263
rect 36144 39156 36156 39359
rect 36864 39156 36876 39359
rect 38664 39156 38676 39455
rect 38856 39156 38868 39503
rect 38928 39156 38940 39263
rect 39024 39156 39036 39455
rect 42216 39205 42228 39575
rect 42360 39277 42372 39575
rect 45744 39277 45756 39527
rect 45768 39277 45780 39575
rect 46824 39181 46836 39695
rect 46872 39205 46884 39527
rect 46992 39157 47004 39335
rect 47016 39157 47028 39695
rect 47040 39565 47052 39671
rect 47040 39157 47052 39383
rect 47064 39157 47076 39383
rect 47088 39349 47100 39671
rect 47136 39517 47148 39623
rect 47088 39157 47100 39239
rect 47112 39157 47124 39503
rect 47136 39157 47148 39455
rect 47160 39421 47172 39599
rect 47160 39157 47172 39359
rect 47184 39157 47196 39455
rect 47208 39373 47220 39575
rect 47232 39325 47244 39551
rect 47208 39157 47220 39311
rect 47232 39157 47244 39287
rect 47256 39157 47268 39527
rect 47280 39157 47292 39407
rect 47304 39301 47316 39407
rect 47304 39157 47316 39239
rect 47328 39157 47340 39383
rect 47352 39277 47364 39359
rect 47376 39277 47388 39335
rect 47400 39205 47412 39311
rect 47424 39205 47436 39287
rect 47448 39205 47460 39263
rect 35874 39144 35892 39156
rect 36138 39144 36156 39156
rect 36858 39144 36876 39156
rect 38657 39144 38676 39156
rect 38849 39144 38868 39156
rect 38921 39144 38940 39156
rect 39017 39144 39036 39156
rect 22121 39133 22133 39143
rect 25457 39133 25469 39143
rect 25697 39133 25709 39143
rect 26657 39133 26669 39143
rect 26849 39133 26861 39143
rect 27883 39133 27895 39143
rect 35874 39133 35886 39144
rect 36138 39133 36150 39144
rect 36858 39133 36870 39144
rect 38657 39133 38669 39144
rect 38849 39133 38861 39144
rect 38921 39133 38933 39144
rect 39017 39133 39029 39144
rect 46824 39133 46836 39143
rect 50256 38965 50268 38999
rect 50256 38821 50268 38855
rect 20280 38773 20292 38807
rect 21216 38773 21228 38807
rect 46992 36349 47004 36455
rect 47016 36349 47028 36455
rect 47040 36349 47052 36455
rect 47064 36349 47076 36455
rect 47088 36349 47100 36455
rect 47112 36349 47124 36455
rect 47136 36349 47148 36455
rect 47160 36349 47172 36455
rect 47184 36349 47196 36455
rect 47208 36349 47220 36455
rect 47232 36349 47244 36455
rect 47256 36349 47268 36455
rect 47280 36349 47292 36455
rect 47304 36349 47316 36455
rect 47328 36349 47340 36455
rect 47352 36349 47364 36455
rect 47376 36349 47388 36455
rect 47400 36349 47412 36455
rect 47424 36349 47436 36455
rect 47448 36421 47460 36455
rect 46992 35245 47004 35351
rect 47016 35245 47028 35351
rect 47040 35245 47052 35351
rect 47064 35245 47076 35351
rect 47088 35245 47100 35351
rect 47112 35245 47124 35351
rect 47136 35245 47148 35351
rect 47160 35245 47172 35351
rect 47184 35245 47196 35351
rect 47208 35245 47220 35351
rect 47232 35245 47244 35351
rect 47256 35245 47268 35351
rect 47280 35245 47292 35351
rect 47304 35245 47316 35351
rect 47328 35245 47340 35351
rect 47352 35245 47364 35351
rect 47376 35245 47388 35351
rect 47400 35317 47412 35351
rect 50232 34933 50244 34967
rect 50256 34933 50268 34967
rect 20256 34717 20268 34751
rect 20280 34717 20292 34823
rect 50184 34813 50196 34847
rect 50208 34813 50220 34847
rect 50256 34789 50268 34823
rect 46992 34117 47004 34223
rect 47016 34117 47028 34223
rect 47040 34117 47052 34223
rect 47064 34117 47076 34223
rect 47088 34117 47100 34223
rect 47112 34117 47124 34223
rect 47136 34117 47148 34223
rect 47160 34117 47172 34223
rect 47184 34117 47196 34223
rect 47208 34117 47220 34223
rect 47232 34117 47244 34223
rect 47256 34117 47268 34223
rect 47280 34117 47292 34223
rect 47304 34117 47316 34223
rect 47328 34117 47340 34223
rect 47352 34189 47364 34223
rect 46992 33013 47004 33119
rect 47016 33013 47028 33119
rect 47040 33013 47052 33119
rect 47064 33013 47076 33119
rect 47088 33013 47100 33119
rect 47112 33013 47124 33119
rect 47136 33013 47148 33119
rect 47160 33013 47172 33119
rect 47184 33013 47196 33119
rect 47208 33013 47220 33119
rect 47232 33013 47244 33119
rect 47256 33013 47268 33119
rect 47280 33013 47292 33119
rect 47304 33085 47316 33119
rect 46992 31909 47004 32015
rect 47016 31909 47028 32015
rect 47040 31909 47052 32015
rect 47064 31909 47076 32015
rect 47088 31909 47100 32015
rect 47112 31909 47124 32015
rect 47136 31909 47148 32015
rect 47160 31909 47172 32015
rect 47184 31909 47196 32015
rect 47208 31909 47220 32015
rect 47232 31909 47244 32015
rect 47256 31909 47268 32015
rect 47280 31909 47292 32015
rect 50208 30925 50220 30959
rect 50256 30901 50268 30935
rect 46992 30805 47004 30887
rect 47016 30805 47028 30887
rect 47040 30805 47052 30887
rect 47064 30805 47076 30887
rect 47088 30805 47100 30887
rect 47112 30805 47124 30887
rect 47136 30805 47148 30887
rect 47160 30805 47172 30887
rect 47184 30805 47196 30887
rect 47208 30805 47220 30887
rect 47232 30805 47244 30887
rect 47256 30805 47268 30887
rect 47280 30805 47292 30887
rect 20256 30685 20268 30767
rect 20280 30685 20292 30767
rect 20304 30733 20316 30767
rect 21216 30733 21228 30767
rect 50232 30757 50244 30791
rect 50256 30757 50268 30791
rect 46992 29677 47004 29783
rect 47016 29677 47028 29783
rect 47040 29677 47052 29783
rect 47064 29677 47076 29783
rect 47088 29677 47100 29783
rect 47112 29677 47124 29783
rect 47136 29677 47148 29783
rect 47160 29677 47172 29783
rect 47184 29677 47196 29783
rect 47208 29677 47220 29783
rect 47232 29677 47244 29783
rect 47256 29677 47268 29783
rect 47280 29677 47292 29783
rect 46992 28573 47004 28679
rect 47016 28573 47028 28679
rect 47040 28573 47052 28679
rect 47064 28573 47076 28679
rect 47088 28573 47100 28679
rect 47112 28573 47124 28679
rect 47136 28573 47148 28679
rect 47160 28573 47172 28679
rect 47184 28573 47196 28679
rect 47208 28573 47220 28679
rect 47232 28573 47244 28679
rect 47280 28597 47292 28703
rect 47304 28597 47316 28631
rect 46992 27469 47004 27551
rect 47016 27517 47028 27551
rect 47040 27493 47052 27527
rect 47064 27493 47076 27575
rect 47088 27493 47100 27575
rect 47112 27493 47124 27575
rect 47136 27493 47148 27575
rect 47160 27493 47172 27575
rect 47184 27493 47196 27575
rect 47208 27493 47220 27575
rect 47232 27493 47244 27575
rect 47256 27493 47268 27575
rect 47280 27493 47292 27575
rect 47304 27493 47316 27575
rect 47328 27493 47340 27575
rect 47352 27493 47364 27527
rect 20280 26773 20292 26807
rect 50256 26773 50268 26807
rect 50293 26784 50307 26796
rect 46992 26413 47004 26447
rect 47016 26365 47028 26447
rect 47040 26365 47052 26447
rect 47064 26365 47076 26399
rect 47088 26365 47100 26471
rect 47112 26365 47124 26471
rect 47136 26365 47148 26471
rect 47160 26365 47172 26471
rect 47184 26365 47196 26471
rect 47208 26365 47220 26471
rect 47232 26365 47244 26471
rect 47256 26365 47268 26471
rect 47280 26365 47292 26471
rect 47304 26365 47316 26471
rect 47328 26365 47340 26471
rect 47352 26365 47364 26471
rect 47376 26365 47388 26399
rect 46992 25237 47004 25343
rect 47016 25237 47028 25343
rect 47040 25237 47052 25343
rect 47064 25237 47076 25343
rect 47088 25237 47100 25343
rect 47136 25333 47148 25367
rect 47160 25333 47172 25367
rect 47184 25333 47196 25367
rect 47208 25333 47220 25367
rect 47232 25333 47244 25367
rect 47112 25237 47124 25271
rect 47136 25237 47148 25271
rect 47160 25237 47172 25271
rect 47184 25237 47196 25271
rect 47208 25237 47220 25271
rect 47256 25261 47268 25367
rect 47280 25261 47292 25367
rect 47304 25261 47316 25367
rect 47328 25261 47340 25367
rect 47352 25261 47364 25367
rect 47376 25261 47388 25367
rect 47400 25261 47412 25367
rect 47424 25261 47436 25295
rect 46992 24133 47004 24239
rect 47016 24133 47028 24239
rect 47040 24133 47052 24239
rect 47064 24133 47076 24239
rect 47088 24133 47100 24239
rect 47112 24133 47124 24239
rect 47136 24205 47148 24239
rect 47160 24157 47172 24239
rect 47184 24157 47196 24239
rect 47208 24157 47220 24239
rect 47232 24157 47244 24239
rect 47256 24157 47268 24191
rect 47280 24157 47292 24263
rect 47304 24157 47316 24263
rect 47328 24157 47340 24263
rect 47352 24157 47364 24263
rect 47376 24157 47388 24263
rect 47400 24157 47412 24263
rect 47424 24157 47436 24263
rect 47448 24157 47460 24263
rect 47472 24157 47484 24191
rect 46992 23029 47004 23111
rect 47016 23029 47028 23111
rect 47040 23029 47052 23111
rect 47064 23029 47076 23111
rect 47088 23029 47100 23063
rect 47112 23029 47124 23135
rect 47136 23029 47148 23135
rect 47160 23029 47172 23135
rect 47184 23029 47196 23135
rect 47208 23029 47220 23135
rect 47232 23029 47244 23135
rect 47256 23029 47268 23135
rect 47280 23029 47292 23135
rect 47304 23029 47316 23135
rect 47328 23029 47340 23135
rect 47352 23029 47364 23135
rect 47376 23101 47388 23135
rect 47400 23053 47412 23135
rect 47424 23053 47436 23135
rect 47448 23053 47460 23135
rect 47472 23053 47484 23135
rect 47496 23053 47508 23135
rect 47520 23053 47532 23087
rect 20280 22813 20292 22847
rect 20304 22813 20316 22847
rect 46992 21901 47004 22007
rect 47016 21901 47028 22007
rect 47040 21901 47052 22007
rect 47064 21901 47076 22007
rect 47088 21901 47100 22007
rect 47112 21901 47124 22007
rect 47136 21901 47148 22007
rect 47160 21973 47172 22007
rect 47184 21925 47196 22007
rect 47208 21925 47220 22007
rect 47232 21925 47244 21959
rect 47256 21925 47268 22031
rect 47280 21925 47292 22031
rect 47304 21925 47316 22031
rect 47328 21925 47340 22031
rect 47352 21925 47364 22031
rect 47376 21925 47388 22031
rect 47400 21925 47412 22031
rect 47424 21925 47436 22031
rect 47448 21925 47460 22031
rect 47472 21925 47484 22031
rect 47496 21925 47508 22031
rect 47520 21925 47532 22031
rect 47544 21925 47556 22031
rect 47568 21925 47580 21959
rect 46992 20797 47004 20903
rect 47016 20797 47028 20903
rect 47040 20797 47052 20903
rect 47064 20797 47076 20903
rect 47088 20797 47100 20903
rect 47112 20797 47124 20903
rect 47136 20797 47148 20903
rect 47160 20797 47172 20903
rect 47184 20797 47196 20903
rect 47208 20869 47220 20903
rect 47232 20821 47244 20903
rect 47256 20821 47268 20903
rect 47280 20821 47292 20903
rect 47304 20821 47316 20903
rect 47328 20821 47340 20903
rect 47352 20821 47364 20903
rect 47376 20821 47388 20903
rect 47400 20821 47412 20903
rect 47424 20821 47436 20903
rect 47448 20821 47460 20903
rect 47472 20821 47484 20903
rect 47496 20821 47508 20903
rect 47520 20821 47532 20903
rect 47544 20821 47556 20903
rect 47568 20821 47580 20855
rect 47592 20821 47604 20927
rect 47616 20821 47628 20855
rect 46992 19693 47004 19775
rect 47016 19693 47028 19775
rect 47040 19693 47052 19775
rect 47064 19693 47076 19775
rect 47088 19693 47100 19775
rect 47112 19693 47124 19775
rect 47136 19693 47148 19775
rect 47160 19693 47172 19775
rect 47184 19693 47196 19775
rect 47208 19693 47220 19775
rect 47232 19741 47244 19775
rect 47256 19717 47268 19751
rect 47280 19717 47292 19799
rect 47304 19717 47316 19799
rect 47328 19717 47340 19799
rect 47352 19717 47364 19799
rect 47376 19717 47388 19799
rect 47400 19717 47412 19799
rect 47424 19717 47436 19799
rect 47448 19717 47460 19799
rect 47472 19717 47484 19799
rect 47496 19717 47508 19799
rect 47520 19717 47532 19799
rect 47544 19717 47556 19799
rect 47568 19717 47580 19799
rect 47592 19717 47604 19799
rect 47616 19717 47628 19799
rect 47640 19717 47652 19799
rect 47664 19717 47676 19751
rect 20304 19597 20316 19631
rect 21120 19597 21132 19631
rect 21216 19597 21228 19631
rect 21384 19597 21396 19631
rect 21432 19597 21444 19655
rect 21216 19477 21228 19511
rect 21384 19477 21396 19511
rect 21432 19477 21444 19511
rect 21480 19477 21492 19511
rect 21536 19477 21548 19643
rect 21559 19438 21571 19643
rect 21582 19621 21594 19643
rect 21605 19477 21617 19643
rect 21628 19477 21640 19643
rect 21651 19573 21663 19643
rect 21674 19608 21686 19643
rect 21697 19633 21709 19643
rect 21697 19621 21716 19633
rect 22008 19621 22020 19643
rect 21674 19595 21692 19608
rect 21680 19477 21692 19595
rect 21704 19477 21716 19621
rect 21752 19477 21764 19559
rect 21776 19477 21788 19511
rect 20256 18757 20268 18791
rect 21672 18613 21684 18647
rect 21560 18469 21572 18503
rect 21624 18469 21636 18576
rect 21648 18397 21660 18551
rect 21672 18469 21684 18551
rect 20304 18349 20316 18383
rect 21216 18349 21228 18383
rect 21384 18349 21396 18383
rect 21432 18349 21444 18383
rect 21480 18349 21492 18383
rect 21560 18349 21572 18383
rect 21672 18325 21684 18431
rect 21696 18325 21708 18551
rect 21720 18325 21732 18551
rect 21750 18517 21762 18599
rect 21774 18565 21786 18599
rect 22008 18282 22020 18599
rect 22121 18282 22133 19643
rect 22145 18373 22157 19643
rect 22169 18445 22181 19643
rect 22145 18282 22157 18359
rect 22169 18282 22181 18431
rect 22193 18282 22205 19643
rect 23441 19621 23453 19643
rect 24233 19621 24245 19643
rect 24785 19621 24797 19643
rect 25001 19621 25013 19643
rect 25745 19621 25757 19643
rect 25913 19621 25925 19643
rect 26297 19621 26309 19643
rect 26489 19621 26501 19643
rect 26705 19621 26717 19643
rect 27449 19621 27461 19643
rect 27617 19621 27629 19643
rect 23441 19607 23447 19621
rect 24233 19607 24239 19621
rect 24785 19607 24791 19621
rect 25001 19607 25007 19621
rect 25745 19607 25751 19621
rect 25913 19607 25919 19621
rect 26297 19607 26303 19621
rect 26489 19607 26495 19621
rect 26705 19607 26711 19621
rect 27449 19607 27455 19621
rect 27617 19607 27623 19621
rect 37025 19620 37037 19643
rect 37217 19620 37229 19643
rect 37457 19620 37469 19643
rect 45161 19620 45173 19643
rect 45905 19620 45917 19643
rect 46121 19621 46133 19643
rect 46265 19621 46277 19643
rect 37025 19608 37044 19620
rect 37217 19608 37236 19620
rect 37457 19608 37476 19620
rect 45161 19608 45180 19620
rect 45905 19608 45924 19620
rect 37032 19573 37044 19608
rect 37224 19573 37236 19608
rect 37464 19573 37476 19608
rect 45168 19573 45180 19608
rect 45192 19525 45204 19559
rect 45912 19549 45924 19608
rect 46121 19607 46127 19621
rect 46265 19607 46271 19621
rect 46313 19620 46325 19643
rect 46361 19621 46373 19643
rect 46409 19621 46421 19643
rect 46313 19608 46332 19620
rect 46296 19549 46308 19583
rect 46320 19573 46332 19608
rect 46361 19607 46367 19621
rect 46409 19607 46415 19621
rect 46481 19620 46493 19643
rect 46481 19608 46500 19620
rect 46488 19573 46500 19608
rect 46824 19525 46836 19643
rect 46992 19477 47004 19607
rect 47016 19477 47028 19607
rect 47040 19477 47052 19607
rect 47064 19477 47076 19559
rect 47088 19477 47100 19631
rect 47112 19477 47124 19631
rect 47136 19477 47148 19631
rect 47160 19477 47172 19631
rect 47184 19477 47196 19631
rect 47208 19477 47220 19631
rect 47232 19477 47244 19631
rect 47256 19477 47268 19631
rect 47280 19477 47292 19631
rect 47304 19477 47316 19631
rect 47328 19477 47340 19631
rect 47352 19477 47364 19631
rect 47376 19477 47388 19631
rect 47400 19477 47412 19631
rect 47424 19477 47436 19631
rect 47448 19477 47460 19631
rect 47472 19477 47484 19631
rect 47496 19477 47508 19631
rect 47520 19477 47532 19631
rect 47544 19477 47556 19631
rect 47568 19477 47580 19631
rect 47592 19477 47604 19631
rect 47616 19477 47628 19631
rect 47640 19477 47652 19631
rect 47664 19477 47676 19631
rect 47688 19477 47700 19631
rect 47712 19477 47724 19559
rect 23448 18565 23460 18599
rect 24240 18565 24252 18599
rect 24792 18565 24804 18599
rect 25008 18565 25020 18599
rect 25752 18565 25764 18599
rect 22224 18373 22236 18551
rect 22248 18445 22260 18527
rect 24216 18493 24228 18527
rect 24192 18324 24204 18479
rect 24264 18349 24276 18527
rect 25104 18517 25116 18551
rect 24192 18312 24209 18324
rect 24197 18282 24209 18312
rect 24233 18311 24239 18325
rect 25080 18324 25092 18503
rect 26784 18445 26796 18671
rect 26760 18324 26772 18431
rect 27624 18421 27636 18695
rect 25080 18312 25097 18324
rect 24233 18282 24245 18311
rect 25085 18282 25097 18312
rect 26753 18312 26772 18324
rect 27600 18324 27612 18407
rect 27672 18373 27684 18671
rect 29328 18469 29340 18647
rect 27648 18324 27660 18359
rect 27600 18312 27617 18324
rect 26753 18282 26765 18312
rect 27605 18282 27617 18312
rect 27641 18312 27660 18324
rect 29304 18324 29316 18455
rect 30192 18397 30204 18623
rect 30168 18324 30180 18383
rect 29304 18312 29321 18324
rect 27641 18282 27653 18312
rect 29309 18282 29321 18312
rect 30161 18312 30180 18324
rect 31008 18324 31020 18623
rect 31896 18493 31908 18599
rect 37032 18565 37044 18599
rect 37224 18565 37236 18599
rect 37464 18565 37476 18599
rect 42864 18565 42876 18599
rect 43704 18565 43716 18599
rect 44544 18565 44556 18599
rect 46205 18565 46217 18599
rect 46229 18565 46241 18599
rect 46992 18565 47004 18599
rect 47016 18565 47028 18599
rect 47040 18565 47052 18599
rect 47064 18565 47076 18599
rect 47088 18565 47100 18599
rect 47112 18565 47124 18599
rect 47136 18565 47148 18599
rect 47160 18565 47172 18599
rect 47184 18565 47196 18599
rect 47208 18565 47220 18599
rect 47232 18565 47244 18599
rect 31872 18324 31884 18479
rect 32736 18349 32748 18551
rect 31008 18312 31025 18324
rect 30161 18282 30173 18312
rect 31013 18282 31025 18312
rect 31865 18312 31884 18324
rect 31865 18282 31877 18312
rect 32725 18311 32729 18325
rect 33576 18324 33588 18527
rect 32717 18282 32729 18311
rect 33569 18312 33588 18324
rect 33600 18324 33612 18503
rect 35304 18349 35316 18479
rect 33600 18312 33617 18324
rect 33569 18282 33581 18312
rect 33605 18282 33617 18312
rect 35273 18311 35279 18325
rect 35273 18282 35285 18311
rect 36125 18282 36137 18455
rect 36173 18397 36185 18431
rect 36149 18282 36161 18383
rect 37824 18349 37836 18479
rect 38496 18397 38508 18455
rect 37813 18311 37817 18325
rect 38472 18324 38484 18383
rect 39432 18373 39444 18431
rect 39408 18324 39420 18359
rect 40320 18324 40332 18407
rect 41040 18324 41052 18359
rect 38472 18312 38489 18324
rect 39408 18312 39425 18324
rect 40320 18312 40337 18324
rect 41040 18312 41057 18324
rect 37805 18282 37817 18311
rect 38477 18282 38489 18312
rect 39413 18282 39425 18312
rect 40325 18282 40337 18312
rect 41045 18282 41057 18312
rect 41557 18311 41561 18325
rect 42037 18311 42041 18325
rect 42877 18311 42881 18325
rect 43717 18311 43721 18325
rect 44557 18311 44561 18325
rect 47064 18324 47076 18407
rect 47904 18324 47916 19055
rect 47064 18312 47081 18324
rect 47904 18312 47921 18324
rect 41549 18282 41561 18311
rect 42029 18282 42041 18311
rect 42869 18282 42881 18311
rect 43709 18282 43721 18311
rect 44549 18282 44561 18311
rect 46205 18282 46217 18311
rect 46229 18282 46241 18311
rect 47069 18282 47081 18312
rect 47909 18282 47921 18312
rect 49128 18282 49140 19031
rect 49416 18325 49428 19007
rect 49440 18325 49452 18983
rect 49464 18325 49476 18959
rect 49488 18325 49500 18935
rect 49512 18325 49524 18911
rect 49536 18325 49548 18887
rect 49560 18325 49572 18863
rect 49584 18325 49596 18839
rect 49608 18325 49620 18815
rect 49632 18325 49644 18791
rect 50256 18757 50268 18791
rect 49656 18325 49668 18743
rect 49680 18325 49692 18719
rect 49704 18325 49716 18695
rect 49728 18325 49740 18671
rect 49752 18325 49764 18647
rect 50256 18613 50268 18647
rect 49776 18325 49788 18599
rect 49800 18325 49812 18575
rect 49824 18325 49836 18551
rect 49848 18325 49860 18527
rect 49872 18325 49884 18527
rect 49896 18325 49908 18503
rect 49920 18325 49932 18479
rect 49944 18325 49956 18455
rect 49992 18325 50004 18431
rect 50040 18325 50052 18407
rect 50160 18325 50172 18383
rect 50208 18325 50220 18359
rect 21432 18200 21444 18239
rect 21480 18176 21492 18239
rect 21672 18176 21684 18239
rect 21696 18176 21708 18239
rect 21720 18176 21732 18239
rect 21757 18211 21782 18223
rect 21757 18187 21782 18199
rect 49359 18115 49391 18127
rect 49359 18091 49391 18103
rect 49359 18067 49391 18079
rect 49359 18043 49391 18055
rect 49359 18019 49391 18031
rect 49416 18008 49428 18138
rect 49440 18008 49452 18138
rect 49464 18008 49476 18138
rect 49488 18008 49500 18114
rect 49512 18008 49524 18186
rect 49536 18008 49548 18186
rect 49560 18008 49572 18186
rect 49584 18032 49596 18186
rect 49608 18032 49620 18186
rect 49632 18032 49644 18186
rect 49656 18032 49668 18186
rect 49680 18032 49692 18186
rect 49704 18032 49716 18186
rect 49728 18032 49740 18186
rect 49752 18080 49764 18186
rect 49776 18080 49788 18186
rect 49800 18080 49812 18186
rect 49824 18080 49836 18186
rect 49848 18080 49860 18186
rect 49872 18152 49884 18186
rect 49896 18104 49908 18186
rect 49920 18104 49932 18186
rect 49944 18104 49956 18186
rect 49359 17077 49405 17078
rect 49359 17066 49391 17077
rect 49416 17053 49428 17087
rect 49440 17053 49452 17087
rect 49464 17053 49476 17087
rect 49488 17053 49500 17087
rect 49512 17053 49524 17087
rect 49536 17053 49548 17087
rect 49560 17053 49572 17087
rect 49608 17053 49620 17087
rect 49632 17053 49644 17087
rect 49656 17053 49668 17087
rect 49680 17053 49692 17087
rect 49512 14773 49524 14807
rect 49536 14773 49548 14807
rect 49560 14773 49572 14807
rect 49608 14773 49620 14807
rect 49632 14773 49644 14807
rect 49656 14773 49668 14807
rect 49680 14773 49692 14807
rect 49728 14773 49740 14807
rect 49800 14773 49812 14807
rect 49824 14773 49836 14807
rect 49848 14773 49860 14807
rect 49896 14773 49908 14807
rect 49920 14773 49932 14807
rect 49944 14773 49956 14807
rect 49992 14773 50004 14807
rect 50040 14773 50052 14807
rect 50160 14773 50172 14807
rect 50208 14749 50220 14807
rect 20256 14701 20268 14735
rect 20304 14701 20316 14735
rect 21216 14701 21228 14735
rect 21480 14701 21492 14735
rect 50232 14725 50244 14807
rect 50256 14725 50268 14759
rect 50232 14581 50244 14615
rect 50256 14581 50268 14615
rect 21480 14103 21492 14137
rect 21696 14077 21708 14137
rect 21720 14077 21732 14137
rect 21757 14114 21782 14126
rect 21757 14090 21782 14102
rect 49359 13261 49405 13262
rect 49359 13250 49391 13261
rect 49416 13237 49428 13271
rect 49440 13237 49452 13271
rect 49464 13237 49476 13271
rect 49512 13237 49524 13271
rect 49536 13237 49548 13271
rect 49560 13237 49572 13271
rect 49359 11882 49391 11894
rect 49359 11858 49391 11870
rect 49416 11847 49428 11905
rect 49440 11847 49452 11905
rect 49464 11847 49476 11905
rect 49512 11847 49524 11905
rect 49536 11847 49548 11905
rect 49560 11847 49572 11905
rect 49632 11847 49644 11905
rect 49656 11871 49668 11905
rect 49680 11871 49692 11905
rect 49728 11871 49740 11905
rect 49359 10713 49391 10725
rect 20256 10669 20268 10703
rect 49359 10689 49391 10701
rect 49416 10677 49428 10735
rect 49440 10677 49452 10735
rect 49464 10677 49476 10735
rect 49512 10677 49524 10735
rect 49536 10677 49548 10735
rect 49560 10677 49572 10735
rect 49632 10677 49644 10735
rect 49680 10701 49692 10735
rect 49728 10701 49740 10735
rect 49824 10701 49836 10735
rect 49848 10701 49860 10735
rect 50256 10669 50268 10703
rect 49440 10525 49452 10559
rect 49464 10525 49476 10559
rect 49512 10525 49524 10559
rect 49536 10525 49548 10559
rect 49560 10525 49572 10559
rect 49632 10525 49644 10559
rect 49728 10525 49740 10559
rect 49824 10525 49836 10559
rect 49848 10525 49860 10559
rect 49920 10525 49932 10559
rect 49944 10525 49956 10559
rect 49992 10525 50004 10559
rect 50040 10525 50052 10559
rect 50256 10525 50268 10559
rect 21696 10333 21708 10400
rect 21720 10333 21732 10400
rect 21757 10377 21782 10389
rect 21757 10353 21782 10365
rect 49359 10329 49391 10341
rect 49359 10305 49391 10317
rect 22121 10260 22133 10294
rect 22193 10261 22205 10294
rect 22121 10248 22140 10260
rect 21672 10165 21684 10247
rect 21696 10165 21708 10247
rect 21720 10165 21732 10247
rect 22128 10213 22140 10248
rect 22193 10247 22199 10261
rect 29729 10260 29741 10294
rect 32909 10260 32921 10294
rect 39221 10260 39233 10294
rect 46733 10260 46745 10294
rect 29729 10248 29748 10260
rect 29736 10237 29748 10248
rect 32904 10248 32921 10260
rect 39216 10248 39233 10260
rect 46728 10248 46745 10260
rect 32904 10237 32916 10248
rect 39216 10237 39228 10248
rect 29736 10165 29748 10223
rect 29760 10189 29772 10223
rect 32904 10165 32916 10223
rect 32928 10189 32940 10223
rect 31800 10117 31812 10151
rect 38856 10117 38868 10175
rect 39216 10117 39228 10223
rect 39240 10189 39252 10223
rect 31656 10021 31668 10055
rect 31800 10021 31812 10055
rect 38856 10021 38868 10055
rect 42240 10021 42252 10175
rect 45936 10069 45948 10223
rect 45960 10189 45972 10223
rect 45984 10093 45996 10175
rect 46728 10093 46740 10248
rect 49440 10141 49452 10351
rect 49464 10293 49476 10351
rect 49512 10293 49524 10351
rect 49536 10317 49548 10351
rect 49560 10317 49572 10351
rect 49512 10189 49524 10223
rect 49728 10093 49740 10175
rect 49824 10093 49836 10175
rect 45912 10021 45924 10055
rect 28128 9805 28140 9839
rect 28272 9805 28284 9839
rect 31656 9805 31668 9839
rect 31800 9805 31812 9839
rect 38712 9805 38724 9839
rect 38856 9805 38868 9863
rect 42240 9805 42252 9863
rect 42384 9805 42396 9863
rect 45768 9805 45780 9887
rect 45912 9805 45924 9935
rect 45984 9829 45996 9863
rect 46008 9829 46020 9887
rect 49944 9829 49956 9935
rect 50040 9853 50052 9887
<< metal4 >>
rect 20373 44585 21933 46145
rect 23899 44585 25459 46145
rect 27425 44585 28985 46145
rect 30951 44585 32511 46145
rect 34477 44585 36037 46145
rect 38003 44585 39563 46145
rect 41529 44585 43089 46145
rect 45055 44585 46615 46145
rect 48581 44585 50141 46145
rect 13835 38133 15395 39693
rect 55119 38133 56679 39693
rect 13835 34091 15395 35651
rect 55119 34091 56679 35651
rect 13835 30049 15395 31609
rect 55119 30049 56679 31609
rect 13835 26007 15395 27567
rect 55119 26007 56679 27567
rect 13835 21965 15395 23525
rect 55119 21965 56679 23525
rect 13835 17923 15395 19483
rect 55119 17923 56679 19483
rect 13835 13881 15395 15441
rect 55119 13881 56679 15441
rect 13835 9839 15395 11399
rect 55119 9839 56679 11399
rect 20373 3387 21933 4947
rect 23899 3387 25459 4947
rect 27425 3387 28985 4947
rect 30951 3387 32511 4947
rect 34477 3387 36037 4947
rect 38003 3387 39563 4947
rect 41529 3387 43089 4947
rect 45055 3387 46615 4947
rect 48581 3387 50141 4947
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 13757 -1 0 46223
box 0 0 6450 6450
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 20293 1 0 39773
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 22013 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 22099 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 22185 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 22271 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 22357 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 22443 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 22529 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 22615 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 22701 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 22787 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 22873 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 22959 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 23045 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 23131 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 23217 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 23303 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 23389 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 23475 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 23561 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 23647 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 23733 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 23819 1 0 39773
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 25539 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 25625 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 25711 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 25797 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 25883 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 25969 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 26055 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 26141 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 26227 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 26313 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 26399 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 26485 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 26571 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 26657 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 26743 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 26829 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 26915 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 27001 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 27087 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 27173 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 27259 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 27345 1 0 39773
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 29065 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 29151 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 29237 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 29323 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 29409 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 29495 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 29581 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 29667 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 29753 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 29839 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 29925 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 30011 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 0 -1 30097 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 0 -1 30183 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 0 -1 30269 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 0 -1 30355 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 0 -1 30441 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 0 -1 30527 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 0 -1 30613 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 0 -1 30699 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 0 -1 30785 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 0 -1 30871 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 32591 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 0 -1 32677 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 0 -1 32763 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 0 -1 32849 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 0 -1 32935 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 0 -1 33021 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 0 -1 33107 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 0 -1 33193 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 0 -1 33279 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 0 -1 33365 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 0 -1 33451 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 0 -1 33537 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 0 -1 33623 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 0 -1 33709 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 0 -1 33795 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 0 -1 33881 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 0 -1 33967 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 0 -1 34053 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 0 -1 34139 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 0 -1 34225 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 0 -1 34311 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 0 -1 34397 1 0 39773
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 36117 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 0 -1 36203 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 0 -1 36289 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 0 -1 36375 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 0 -1 36461 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 0 -1 36547 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 0 -1 36633 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 0 -1 36719 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 0 -1 36805 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 0 -1 36891 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 0 -1 36977 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 0 -1 37063 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 0 -1 37149 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 0 -1 37235 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 0 -1 37321 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 0 -1 37407 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 0 -1 37493 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 0 -1 37579 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 0 -1 37665 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 0 -1 37751 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 0 -1 37837 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 0 -1 37923 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 39643 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 0 -1 39729 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 0 -1 39815 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 0 -1 39901 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 0 -1 39987 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 0 -1 40073 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 0 -1 40159 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 0 -1 40245 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 0 -1 40331 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 0 -1 40417 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 0 -1 40503 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 0 -1 40589 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 0 -1 40675 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 0 -1 40761 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 0 -1 40847 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 0 -1 40933 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 0 -1 41019 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 0 -1 41105 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 0 -1 41191 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 0 -1 41277 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 0 -1 41363 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 0 -1 41449 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 43169 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 0 -1 43255 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 0 -1 43341 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 0 -1 43427 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 0 -1 43513 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 0 -1 43599 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 0 -1 43685 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 0 -1 43771 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 0 -1 43857 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 0 -1 43943 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 0 -1 44029 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 0 -1 44115 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 0 -1 44201 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 0 -1 44287 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 0 -1 44373 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 0 -1 44459 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 0 -1 44545 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 0 -1 44631 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 0 -1 44717 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 0 -1 44803 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 0 -1 44889 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 0 -1 44975 1 0 39773
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 46695 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 0 -1 46781 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 0 -1 46867 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 0 -1 46953 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 0 -1 47039 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 0 -1 47125 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 0 -1 47211 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 0 -1 47297 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 0 -1 47383 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 0 -1 47469 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 0 -1 47555 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 0 -1 47641 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 0 -1 47727 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 0 -1 47813 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 0 -1 47899 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 0 -1 47985 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 0 -1 48071 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 0 -1 48157 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 0 -1 48243 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 0 -1 48329 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 0 -1 48415 1 0 39773
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 0 -1 48501 1 0 39773
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 50221 1 0 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 0 -1 50307 1 0 39773
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 56757 0 -1 46223
box 0 0 6450 6450
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 20207 0 -1 39773
box 0 0 6450 1720
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform -1 0 20207 0 -1 38053
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform -1 0 20207 0 -1 37967
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform -1 0 20207 0 -1 37881
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform -1 0 20207 0 -1 37795
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform -1 0 20207 0 -1 37709
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform -1 0 20207 0 -1 37623
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform -1 0 20207 0 -1 37537
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform -1 0 20207 0 -1 37451
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform -1 0 20207 0 -1 37365
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform -1 0 20207 0 -1 37279
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform -1 0 20207 0 -1 37193
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform -1 0 20207 0 -1 37107
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform -1 0 20207 0 -1 37021
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform -1 0 20207 0 -1 36935
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform -1 0 20207 0 -1 36849
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform -1 0 20207 0 -1 36763
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform -1 0 20207 0 -1 36677
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform -1 0 20207 0 -1 36591
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform -1 0 20207 0 -1 36505
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform -1 0 20207 0 -1 36419
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform -1 0 20207 0 -1 36333
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform -1 0 20207 0 -1 36247
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform -1 0 20207 0 -1 36161
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform -1 0 20207 0 -1 36075
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform -1 0 20207 0 -1 35989
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform -1 0 20207 0 -1 35903
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform -1 0 20207 0 -1 35817
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 20207 0 -1 35731
box 0 0 6450 1720
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform -1 0 20207 0 -1 34011
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform -1 0 20207 0 -1 33925
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform -1 0 20207 0 -1 33839
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform -1 0 20207 0 -1 33753
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform -1 0 20207 0 -1 33667
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform -1 0 20207 0 -1 33581
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform -1 0 20207 0 -1 33495
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform -1 0 20207 0 -1 33409
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform -1 0 20207 0 -1 33323
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform -1 0 20207 0 -1 33237
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform -1 0 20207 0 -1 33151
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform -1 0 20207 0 -1 33065
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform -1 0 20207 0 -1 32979
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform -1 0 20207 0 -1 32893
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform -1 0 20207 0 -1 32807
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform -1 0 20207 0 -1 32721
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform -1 0 20207 0 -1 32635
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform -1 0 20207 0 -1 32549
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform -1 0 20207 0 -1 32463
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform -1 0 20207 0 -1 32377
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform -1 0 20207 0 -1 32291
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform -1 0 20207 0 -1 32205
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform -1 0 20207 0 -1 32119
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform -1 0 20207 0 -1 32033
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform -1 0 20207 0 -1 31947
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform -1 0 20207 0 -1 31861
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform -1 0 20207 0 -1 31775
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 20207 0 -1 31689
box 0 0 6450 1720
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform -1 0 20207 0 -1 29969
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform -1 0 20207 0 -1 29883
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform -1 0 20207 0 -1 29797
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform -1 0 20207 0 -1 29711
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform -1 0 20207 0 -1 29625
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform -1 0 20207 0 -1 29539
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform -1 0 20207 0 -1 29453
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform -1 0 20207 0 -1 29367
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform -1 0 20207 0 -1 29281
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform -1 0 20207 0 -1 29195
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform -1 0 20207 0 -1 29109
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform -1 0 20207 0 -1 29023
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform -1 0 20207 0 -1 28937
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform -1 0 20207 0 -1 28851
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform -1 0 20207 0 -1 28765
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform -1 0 20207 0 -1 28679
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform -1 0 20207 0 -1 28593
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform -1 0 20207 0 -1 28507
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform -1 0 20207 0 -1 28421
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform -1 0 20207 0 -1 28335
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform -1 0 20207 0 -1 28249
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform -1 0 20207 0 -1 28163
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform -1 0 20207 0 -1 28077
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform -1 0 20207 0 -1 27991
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform -1 0 20207 0 -1 27905
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform -1 0 20207 0 -1 27819
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform -1 0 20207 0 -1 27733
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 20207 0 -1 27647
box 0 0 6450 1720
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform -1 0 20207 0 -1 25927
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform -1 0 20207 0 -1 25841
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform -1 0 20207 0 -1 25755
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform -1 0 20207 0 -1 25669
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform -1 0 20207 0 -1 25583
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform -1 0 20207 0 -1 25497
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform -1 0 20207 0 -1 25411
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform -1 0 20207 0 -1 25325
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform -1 0 20207 0 -1 25239
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform -1 0 20207 0 -1 25153
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform -1 0 20207 0 -1 25067
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform -1 0 20207 0 -1 24981
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform -1 0 20207 0 -1 24895
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform -1 0 20207 0 -1 24809
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform -1 0 20207 0 -1 24723
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform -1 0 20207 0 -1 24637
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform -1 0 20207 0 -1 24551
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform -1 0 20207 0 -1 24465
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform -1 0 20207 0 -1 24379
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform -1 0 20207 0 -1 24293
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform -1 0 20207 0 -1 24207
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform -1 0 20207 0 -1 24121
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform -1 0 20207 0 -1 24035
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform -1 0 20207 0 -1 23949
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform -1 0 20207 0 -1 23863
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform -1 0 20207 0 -1 23777
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform -1 0 20207 0 -1 23691
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 20207 0 -1 23605
box 0 0 6450 1720
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform -1 0 20207 0 -1 21885
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform -1 0 20207 0 -1 21799
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform -1 0 20207 0 -1 21713
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform -1 0 20207 0 -1 21627
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform -1 0 20207 0 -1 21541
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform -1 0 20207 0 -1 21455
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform -1 0 20207 0 -1 21369
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform -1 0 20207 0 -1 21283
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform -1 0 20207 0 -1 21197
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform -1 0 20207 0 -1 21111
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform -1 0 20207 0 -1 21025
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform -1 0 20207 0 -1 20939
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform -1 0 20207 0 -1 20853
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform -1 0 20207 0 -1 20767
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform -1 0 20207 0 -1 20681
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform -1 0 20207 0 -1 20595
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform -1 0 20207 0 -1 20509
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform -1 0 20207 0 -1 20423
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform -1 0 20207 0 -1 20337
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform -1 0 20207 0 -1 20251
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform -1 0 20207 0 -1 20165
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform -1 0 20207 0 -1 20079
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform -1 0 20207 0 -1 19993
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform -1 0 20207 0 -1 19907
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform -1 0 20207 0 -1 19821
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform -1 0 20207 0 -1 19735
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform -1 0 20207 0 -1 19649
box 0 0 6450 86
use datapath datapath_0
timestamp 1396719273
transform 1 0 21535 0 1 19643
box 0 0 25408 19490
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 50307 0 1 38053
box 0 0 6450 1720
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 50307 0 1 37967
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 50307 0 1 37881
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 50307 0 1 37795
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 50307 0 1 37709
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 50307 0 1 37623
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 50307 0 1 37537
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 50307 0 1 37451
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 50307 0 1 37365
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 50307 0 1 37279
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 50307 0 1 37193
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 50307 0 1 37107
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 50307 0 1 37021
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 50307 0 1 36935
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 50307 0 1 36849
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 50307 0 1 36763
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 50307 0 1 36677
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 50307 0 1 36591
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 50307 0 1 36505
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 50307 0 1 36419
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 50307 0 1 36333
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 50307 0 1 36247
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 50307 0 1 36161
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 50307 0 1 36075
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 50307 0 1 35989
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 50307 0 1 35903
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 50307 0 1 35817
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 50307 0 1 35731
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 50307 0 1 34011
box 0 0 6450 1720
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 50307 0 1 33925
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 50307 0 1 33839
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 50307 0 1 33753
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 50307 0 1 33667
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 50307 0 1 33581
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 50307 0 1 33495
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 50307 0 1 33409
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 50307 0 1 33323
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 50307 0 1 33237
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 50307 0 1 33151
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 50307 0 1 33065
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 50307 0 1 32979
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 50307 0 1 32893
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 50307 0 1 32807
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 50307 0 1 32721
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 50307 0 1 32635
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 50307 0 1 32549
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 50307 0 1 32463
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 50307 0 1 32377
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 50307 0 1 32291
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 50307 0 1 32205
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 50307 0 1 32119
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 50307 0 1 32033
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 50307 0 1 31947
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 50307 0 1 31861
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 50307 0 1 31775
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 50307 0 1 31689
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 50307 0 1 29969
box 0 0 6450 1720
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 50307 0 1 29883
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 50307 0 1 29797
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 50307 0 1 29711
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 50307 0 1 29625
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 50307 0 1 29539
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 50307 0 1 29453
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 50307 0 1 29367
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 50307 0 1 29281
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 50307 0 1 29195
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 50307 0 1 29109
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 50307 0 1 29023
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 50307 0 1 28937
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 50307 0 1 28851
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 50307 0 1 28765
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 50307 0 1 28679
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 50307 0 1 28593
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 50307 0 1 28507
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 50307 0 1 28421
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 50307 0 1 28335
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 50307 0 1 28249
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 50307 0 1 28163
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 50307 0 1 28077
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 50307 0 1 27991
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 50307 0 1 27905
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 50307 0 1 27819
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 50307 0 1 27733
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 50307 0 1 27647
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 50307 0 1 25927
box 0 0 6450 1720
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 50307 0 1 25841
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 50307 0 1 25755
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 50307 0 1 25669
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 50307 0 1 25583
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 50307 0 1 25497
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 50307 0 1 25411
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 50307 0 1 25325
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 50307 0 1 25239
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 50307 0 1 25153
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 50307 0 1 25067
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 50307 0 1 24981
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 50307 0 1 24895
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 50307 0 1 24809
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 50307 0 1 24723
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 50307 0 1 24637
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 50307 0 1 24551
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 50307 0 1 24465
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 50307 0 1 24379
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 50307 0 1 24293
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 50307 0 1 24207
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 50307 0 1 24121
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 50307 0 1 24035
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 50307 0 1 23949
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 50307 0 1 23863
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 50307 0 1 23777
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 50307 0 1 23691
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 50307 0 1 23605
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 50307 0 1 21885
box 0 0 6450 1720
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 50307 0 1 21799
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 50307 0 1 21713
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 50307 0 1 21627
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 50307 0 1 21541
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 50307 0 1 21455
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 50307 0 1 21369
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 50307 0 1 21283
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 50307 0 1 21197
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 50307 0 1 21111
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 50307 0 1 21025
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 50307 0 1 20939
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 50307 0 1 20853
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 50307 0 1 20767
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 50307 0 1 20681
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 50307 0 1 20595
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 50307 0 1 20509
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 50307 0 1 20423
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 50307 0 1 20337
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 50307 0 1 20251
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 50307 0 1 20165
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 50307 0 1 20079
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 50307 0 1 19993
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 50307 0 1 19907
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 1 0 50307 0 1 19821
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 1 0 50307 0 1 19735
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 1 0 50307 0 1 19649
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 20207 0 -1 19563
box 0 0 6450 1720
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 1 0 50307 0 1 19563
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform -1 0 20207 0 -1 17843
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform -1 0 20207 0 -1 17757
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform -1 0 20207 0 -1 17671
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform -1 0 20207 0 -1 17585
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform -1 0 20207 0 -1 17499
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform -1 0 20207 0 -1 17413
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform -1 0 20207 0 -1 17327
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform -1 0 20207 0 -1 17241
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform -1 0 20207 0 -1 17155
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform -1 0 20207 0 -1 17069
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform -1 0 20207 0 -1 16983
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform -1 0 20207 0 -1 16897
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform -1 0 20207 0 -1 16811
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform -1 0 20207 0 -1 16725
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform -1 0 20207 0 -1 16639
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform -1 0 20207 0 -1 16553
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform -1 0 20207 0 -1 16467
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform -1 0 20207 0 -1 16381
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform -1 0 20207 0 -1 16295
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform -1 0 20207 0 -1 16209
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform -1 0 20207 0 -1 16123
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform -1 0 20207 0 -1 16037
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform -1 0 20207 0 -1 15951
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform -1 0 20207 0 -1 15865
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform -1 0 20207 0 -1 15779
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform -1 0 20207 0 -1 15693
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform -1 0 20207 0 -1 15607
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 20207 0 -1 15521
box 0 0 6450 1720
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform -1 0 20207 0 -1 13801
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform -1 0 20207 0 -1 13715
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform -1 0 20207 0 -1 13629
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform -1 0 20207 0 -1 13543
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform -1 0 20207 0 -1 13457
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform -1 0 20207 0 -1 13371
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform -1 0 20207 0 -1 13285
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform -1 0 20207 0 -1 13199
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform -1 0 20207 0 -1 13113
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform -1 0 20207 0 -1 13027
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform -1 0 20207 0 -1 12941
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform -1 0 20207 0 -1 12855
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 20207 0 -1 12769
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 20207 0 -1 12683
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 20207 0 -1 12597
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 20207 0 -1 12511
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 20207 0 -1 12425
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 20207 0 -1 12339
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 20207 0 -1 12253
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 20207 0 -1 12167
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 20207 0 -1 12081
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 20207 0 -1 11995
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 20207 0 -1 11909
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 20207 0 -1 11823
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 20207 0 -1 11737
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 20207 0 -1 11651
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 20207 0 -1 11565
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 20207 0 -1 11479
box 0 0 6450 1720
use control control_0
timestamp 1396906397
transform 1 0 21782 0 1 10294
box 0 0 27577 7988
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 50307 0 1 17843
box 0 0 6450 1720
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 1 0 50307 0 1 17757
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 1 0 50307 0 1 17671
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 1 0 50307 0 1 17585
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 1 0 50307 0 1 17499
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 1 0 50307 0 1 17413
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 1 0 50307 0 1 17327
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 1 0 50307 0 1 17241
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 1 0 50307 0 1 17155
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 1 0 50307 0 1 17069
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 1 0 50307 0 1 16983
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 1 0 50307 0 1 16897
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 1 0 50307 0 1 16811
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 1 0 50307 0 1 16725
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 1 0 50307 0 1 16639
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 1 0 50307 0 1 16553
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 1 0 50307 0 1 16467
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 1 0 50307 0 1 16381
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 1 0 50307 0 1 16295
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 1 0 50307 0 1 16209
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 1 0 50307 0 1 16123
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 1 0 50307 0 1 16037
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 1 0 50307 0 1 15951
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 1 0 50307 0 1 15865
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 1 0 50307 0 1 15779
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 1 0 50307 0 1 15693
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 1 0 50307 0 1 15607
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 1 0 50307 0 1 15521
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 50307 0 1 13801
box 0 0 6450 1720
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 1 0 50307 0 1 13715
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 1 0 50307 0 1 13629
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 1 0 50307 0 1 13543
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 1 0 50307 0 1 13457
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 1 0 50307 0 1 13371
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 1 0 50307 0 1 13285
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 1 0 50307 0 1 13199
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 1 0 50307 0 1 13113
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 1 0 50307 0 1 13027
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 1 0 50307 0 1 12941
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 1 0 50307 0 1 12855
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 1 0 50307 0 1 12769
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 1 0 50307 0 1 12683
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 1 0 50307 0 1 12597
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 1 0 50307 0 1 12511
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 1 0 50307 0 1 12425
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 1 0 50307 0 1 12339
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 1 0 50307 0 1 12253
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 1 0 50307 0 1 12167
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 1 0 50307 0 1 12081
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 1 0 50307 0 1 11995
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 1 0 50307 0 1 11909
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 1 0 50307 0 1 11823
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 1 0 50307 0 1 11737
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 1 0 50307 0 1 11651
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 1 0 50307 0 1 11565
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 1 0 50307 0 1 11479
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 50307 0 1 9759
box 0 0 6450 1720
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 13757 0 1 3309
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 20207 -1 0 9759
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 20293 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 22013 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 22099 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 22185 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 22271 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 22357 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 22443 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 22529 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 22615 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 22701 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 22787 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 22873 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 22959 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 23045 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 23131 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 23217 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 23303 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 23389 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 23475 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 23561 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 23647 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 23733 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 23819 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 25539 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 25625 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 25711 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 25797 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 25883 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 25969 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 26055 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 26141 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 26227 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 26313 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 26399 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 26485 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 26571 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 26657 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 26743 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 26829 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 26915 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 27001 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 27087 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 27173 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 27259 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 27345 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 29065 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 29151 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 29237 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 29323 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 29409 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 29495 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 29581 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 29667 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 29753 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 29839 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 29925 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 30011 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 30097 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 30183 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 30269 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 30355 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 30441 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 30527 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 30613 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 30699 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 30785 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 30871 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 32591 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 32677 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 32763 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 32849 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 32935 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 33021 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 33107 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 33193 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 33279 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 33365 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 33451 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 33537 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 33623 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 33709 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 33795 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 33881 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 33967 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 34053 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 34139 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 34225 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 34311 -1 0 9759
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 34397 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 36117 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 36203 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 36289 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 36375 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 36461 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 36547 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 36633 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 36719 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 36805 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 36891 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 36977 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 37063 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 37149 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 37235 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 37321 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 37407 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 37493 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 37579 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 37665 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 37751 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 37837 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 37923 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 39643 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 39729 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 39815 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 39901 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 39987 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 40073 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 40159 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 40245 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 40331 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 40417 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 40503 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 40589 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 40675 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 40761 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 40847 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 40933 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 41019 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 41105 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 41191 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 41277 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 41363 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 41449 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 43169 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 43255 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 43341 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 43427 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 43513 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 43599 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 43685 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 43771 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 43857 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 43943 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 44029 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 44115 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 44201 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 44287 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 44373 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 44459 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 44545 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 44631 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 44717 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 44803 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 44889 -1 0 9759
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 44975 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 46695 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 46781 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 46867 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 46953 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 47039 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 47125 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 47211 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 47297 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 47383 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 47469 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 47555 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 47641 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 47727 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 47813 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 47899 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 47985 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 48071 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 48157 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 48243 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 48329 -1 0 9759
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 48415 -1 0 9759
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 48501 -1 0 9759
box 0 0 6450 1720
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 50221 -1 0 9759
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 56757 1 0 3309
box 0 0 6450 6450
<< labels >>
rlabel metal4 20373 3387 21933 4947 0 nIRQ
rlabel metal4 23899 3387 25459 4947 0 Data[0]
rlabel metal4 27425 3387 28985 4947 0 Data[1]
rlabel metal4 30951 3387 32511 4947 0 Data[2]
rlabel metal4 34477 3387 36037 4947 0 vdde!
rlabel metal4 38003 3387 39563 4947 0 Data[3]
rlabel metal4 41529 3387 43089 4947 0 Data[4]
rlabel metal4 45055 3387 46615 4947 0 Data[5]
rlabel metal4 48581 3387 50141 4947 0 gnde!
rlabel metal4 55119 9839 56679 11399 0 Data[6]
rlabel metal4 55119 13881 56679 15441 0 Data[7]
rlabel metal4 55119 17923 56679 19483 0 Data[8]
rlabel metal4 55119 21965 56679 23525 0 gnde!
rlabel metal4 55119 26007 56679 27567 0 GND!
rlabel metal4 55119 30049 56679 31609 0 Data[9]
rlabel metal4 55119 34091 56679 35651 0 Data[10]
rlabel metal4 55119 38133 56679 39693 0 Data[11]
rlabel metal4 48581 44585 50141 46145 0 vdde!
rlabel metal4 45055 44585 46615 46145 0 Data[12]
rlabel metal4 41529 44585 43089 46145 0 Data[13]
rlabel metal4 38003 44585 39563 46145 0 Data[14]
rlabel metal4 34477 44585 36037 46145 0 gnde!
rlabel metal4 30951 44585 32511 46145 0 Data[15]
rlabel metal4 27425 44585 28985 46145 0 ALE
rlabel metal4 23899 44585 25459 46145 0 nME
rlabel metal4 20373 44585 21933 46145 0 nWait
rlabel metal4 13835 38133 15395 39693 0 nOE
rlabel metal4 13835 34091 15395 35651 0 RnW
rlabel metal4 13835 30049 15395 31609 0 SDO
rlabel metal4 13835 26007 15395 27567 0 Vdd!
rlabel metal4 13835 21965 15395 23525 0 SDI
rlabel metal4 13835 17923 15395 19483 0 Test
rlabel metal4 13835 13881 15395 15441 0 Clock
rlabel metal4 13835 9839 15395 11399 0 nReset
<< end >>
