magic
tech c035u
timestamp 1397219778
<< metal1 >>
rect 1539 1082 1549 1106
rect 1573 1094 3215 1104
rect 3229 1094 20472 1104
rect 1539 1072 1575 1082
rect 12552 965 12623 975
rect 12552 943 12863 953
rect 12901 944 13055 954
rect 13141 938 13176 948
rect 12709 916 13176 926
rect 12973 84 13103 94
rect 2821 65 12671 75
rect 0 29 3095 39
rect 3109 29 3263 39
rect 3277 29 20472 39
rect 0 7 12815 17
<< m2contact >>
rect 1559 1092 1573 1106
rect 3215 1092 3229 1106
rect 12623 963 12637 977
rect 12863 941 12877 955
rect 12887 940 12901 954
rect 13055 942 13069 956
rect 13127 936 13141 950
rect 12695 914 12709 928
rect 12959 80 12973 94
rect 13103 82 13117 96
rect 2807 64 2821 78
rect 12671 63 12685 77
rect 3095 27 3109 41
rect 3263 27 3277 41
rect 12815 5 12829 19
<< metal2 >>
rect 216 1000 228 1111
rect 360 1000 372 1111
rect 576 1000 588 1111
rect 1320 1000 1332 1111
rect 1488 1000 1500 1111
rect 1560 1000 1572 1092
rect 1872 1000 1884 1111
rect 2064 1000 2076 1111
rect 2280 1000 2292 1111
rect 3024 1000 3036 1111
rect 3192 911 3204 1111
rect 3216 911 3228 1092
rect 3288 982 3372 994
rect 3408 982 3420 1111
rect 4152 982 4164 1111
rect 4368 982 4380 1111
rect 4560 982 4572 1111
rect 5304 982 5316 1111
rect 5520 982 5532 1111
rect 5712 982 5724 1111
rect 6456 982 6468 1111
rect 6672 982 6684 1111
rect 6864 982 6876 1111
rect 7608 982 7620 1111
rect 7824 982 7836 1111
rect 8016 982 8028 1111
rect 8760 982 8772 1111
rect 8976 982 8988 1111
rect 9168 982 9180 1111
rect 9912 982 9924 1111
rect 10128 982 10140 1111
rect 10320 982 10332 1111
rect 11064 982 11076 1111
rect 11280 982 11292 1111
rect 11472 982 11484 1111
rect 12216 982 12228 1111
rect 12432 982 12444 1111
rect 3288 911 3300 982
rect 12600 911 12612 1111
rect 12624 911 12636 963
rect 12696 911 12708 914
rect 12792 911 12804 1111
rect 12864 911 12876 941
rect 12888 911 12900 940
rect 13032 911 13044 1111
rect 13248 1088 13260 1111
rect 13512 1088 13524 1111
rect 13680 1088 13692 1111
rect 13848 1088 13860 1111
rect 13872 1088 13884 1111
rect 13944 1088 13956 1111
rect 14160 1088 14172 1111
rect 14304 1088 14316 1111
rect 14640 1088 14652 1111
rect 15000 1088 15012 1111
rect 15408 1088 15420 1111
rect 15744 1088 15756 1111
rect 16056 1088 16068 1111
rect 16392 1088 16404 1111
rect 16512 1088 16524 1111
rect 16560 1088 16572 1111
rect 16728 1088 16740 1111
rect 16824 1088 16836 1111
rect 16872 1088 16884 1111
rect 16920 1088 16932 1111
rect 16968 1088 16980 1111
rect 17016 1088 17028 1111
rect 17064 1088 17076 1111
rect 17112 1088 17124 1111
rect 17160 1088 17172 1111
rect 17472 1088 17484 1111
rect 17520 1088 17532 1111
rect 17568 1088 17580 1111
rect 17616 1088 17628 1111
rect 17928 1088 17940 1111
rect 17976 1088 17988 1111
rect 18360 1088 18372 1111
rect 18528 1088 18540 1111
rect 18553 1088 18565 1111
rect 18600 1088 18612 1111
rect 18648 1088 18660 1111
rect 18696 1088 18708 1111
rect 18744 1088 18756 1111
rect 18792 1088 18804 1111
rect 18840 1088 18852 1111
rect 18888 1088 18900 1111
rect 18936 1088 18948 1111
rect 19176 1088 19188 1111
rect 19248 1088 19260 1111
rect 19296 1088 19308 1111
rect 19344 1088 19356 1111
rect 19392 1088 19404 1111
rect 19632 1088 19644 1111
rect 19704 1088 19716 1111
rect 19752 1088 19764 1111
rect 19992 1088 20004 1111
rect 20064 1088 20076 1111
rect 20352 1088 20364 1111
rect 13056 911 13068 942
rect 13128 911 13140 936
rect 216 0 228 83
rect 360 0 372 83
rect 576 0 588 83
rect 1320 0 1332 83
rect 1488 0 1500 83
rect 1872 0 1884 83
rect 2064 0 2076 83
rect 2280 0 2292 83
rect 2808 78 2820 83
rect 3024 0 3036 83
rect 3096 41 3108 83
rect 3192 0 3204 112
rect 3264 41 3276 112
rect 3408 0 3420 88
rect 4152 0 4164 88
rect 4368 0 4380 88
rect 4560 0 4572 88
rect 5304 0 5316 88
rect 5520 0 5532 88
rect 5712 0 5724 88
rect 6456 0 6468 88
rect 6672 0 6684 88
rect 6864 0 6876 88
rect 7608 0 7620 88
rect 7824 0 7836 88
rect 8016 0 8028 88
rect 8760 0 8772 88
rect 8976 0 8988 88
rect 9168 0 9180 88
rect 9912 0 9924 88
rect 10128 0 10140 88
rect 10320 0 10332 88
rect 11064 0 11076 88
rect 11280 0 11292 88
rect 11472 0 11484 88
rect 12216 0 12228 88
rect 12432 0 12444 88
rect 12600 0 12612 112
rect 12672 77 12684 112
rect 12696 100 12708 112
rect 12792 0 12804 112
rect 12816 19 12828 112
rect 12960 94 12972 112
rect 13032 0 13044 112
rect 13104 96 13116 112
rect 13128 100 13140 112
rect 13248 0 13260 46
rect 13512 0 13524 46
rect 13680 0 13692 46
rect 13872 0 13884 46
rect 14160 0 14172 46
rect 14304 0 14316 46
rect 14640 0 14652 46
rect 15000 0 15012 46
rect 15408 0 15420 46
rect 15744 0 15756 46
rect 16056 0 16068 46
rect 16392 0 16404 46
rect 16560 0 16572 46
rect 16728 0 16740 46
rect 16824 0 16836 46
rect 16872 0 16884 46
rect 16920 0 16932 46
rect 16968 0 16980 46
rect 17016 0 17028 46
rect 17064 0 17076 46
rect 17112 0 17124 46
rect 17160 0 17172 46
rect 17472 0 17484 46
rect 17520 0 17532 46
rect 17568 0 17580 46
rect 17616 0 17628 46
rect 17928 0 17940 46
rect 17976 0 17988 46
rect 18360 0 18372 46
rect 18528 0 18540 46
rect 18553 0 18565 46
rect 18600 0 18612 46
rect 18648 0 18660 46
rect 18696 0 18708 46
rect 18744 0 18756 46
rect 18792 0 18804 46
rect 18840 0 18852 46
rect 18888 0 18900 46
rect 18936 0 18948 46
rect 19176 0 19188 46
rect 19248 0 19260 46
rect 19296 0 19308 46
rect 19344 0 19356 46
rect 19392 0 19404 46
rect 19632 0 19644 46
rect 19704 0 19716 46
rect 19752 0 19764 46
rect 19992 0 20004 46
rect 20064 0 20076 46
rect 20352 0 20364 46
use Pc_slice Pc_slice_0
timestamp 1396719273
transform 1 0 0 0 1 46
box 0 37 3144 954
use mux2 mux2_0
timestamp 1386235218
transform 1 0 3144 0 1 112
box 0 0 192 799
use regBlock_slice regBlock_slice_0
timestamp 1396393625
transform 1 0 3336 0 1 67
box 0 21 9216 915
use mux2 mux2_1
timestamp 1386235218
transform 1 0 12552 0 1 112
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 12744 0 1 112
box 0 0 192 799
use tielow tielow_0
timestamp 1386086605
transform 1 0 12936 0 1 112
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 12984 0 1 112
box 0 0 192 799
use ALUSlice ALUSlice_0
timestamp 1397052528
transform 1 0 13176 0 1 46
box 0 0 7296 1042
<< labels >>
rlabel metal2 12792 1111 12804 1111 5 Op2Sel[0]
rlabel metal2 13032 1111 13044 1111 5 Op2Sel[1]
rlabel metal2 20064 1111 20076 1111 5 Sh1_R_in
rlabel metal2 16824 1111 16836 1111 5 Sh8Z_L
rlabel metal2 17160 1111 17172 1111 5 Sh8G_L
rlabel metal2 17064 1111 17076 1111 5 Sh8E_L
rlabel metal2 17112 1111 17124 1111 5 Sh8F_L
rlabel metal2 16920 1111 16932 1111 5 Sh8B_L
rlabel metal2 17016 1111 17028 1111 5 Sh8D_L
rlabel metal2 16968 1111 16980 1111 5 Sh8C_L
rlabel metal2 16872 1111 16884 1111 5 Sh8A_L
rlabel metal1 20472 1094 20472 1104 7 AluOut
rlabel metal2 16512 1111 16524 1111 5 A
rlabel metal2 18360 1111 18372 1111 5 Sh1_L_Out
rlabel metal2 18528 1111 18540 1111 5 Sh8
rlabel metal2 18696 1111 18708 1111 5 Sh8C_R
rlabel metal2 18648 1111 18660 1111 5 Sh8B_R
rlabel metal2 18600 1111 18612 1111 5 Sh8A_R
rlabel metal2 17616 1111 17628 1111 5 Sh4C_L
rlabel metal2 17568 1111 17580 1111 5 Sh4B_L
rlabel metal2 17976 1111 17988 1111 5 Sh2B_L
rlabel metal2 17928 1111 17940 1111 5 Sh2A_L
rlabel metal2 18553 1111 18565 1111 5 ShR
rlabel metal2 17520 1111 17532 1111 5 Sh4A_L
rlabel metal2 17472 1111 17484 1111 5 Sh4Z_L
rlabel metal2 19248 1111 19260 1111 5 Sh4Z_R
rlabel metal2 19992 1111 20004 1111 5 Sh1
rlabel metal2 19632 1111 19644 1111 5 Sh2
rlabel metal2 20352 1111 20364 1111 5 ShOut
rlabel metal2 19752 1111 19764 1111 5 Sh2B_R
rlabel metal2 19704 1111 19716 1111 5 Sh2A_R
rlabel metal2 19392 1111 19404 1111 5 Sh4C_R
rlabel metal2 19344 1111 19356 1111 5 Sh4B_R
rlabel metal2 19296 1111 19308 1111 5 Sh4A_R
rlabel metal2 19176 1111 19188 1111 5 Sh4
rlabel metal2 18744 1111 18756 1111 5 Sh8D_R
rlabel metal2 18792 1111 18804 1111 5 Sh8E_R
rlabel metal2 18840 1111 18852 1111 5 Sh8F_R
rlabel metal2 18888 1111 18900 1111 5 Sh8G_R
rlabel metal2 18936 1111 18948 1111 5 Sh8H_R
rlabel metal2 13248 1111 13260 1111 5 ZeroA
rlabel metal2 13680 1111 13692 1111 5 CIn
rlabel metal2 13944 1111 13956 1111 5 Sum
rlabel metal2 13872 1111 13884 1111 5 COut
rlabel metal2 16560 1111 16572 1111 5 ShB
rlabel metal2 16392 1111 16404 1111 5 NOR
rlabel metal2 16056 1111 16068 1111 5 NAND
rlabel metal2 15744 1111 15756 1111 5 NOT
rlabel metal2 15408 1111 15420 1111 5 XOR
rlabel metal2 15000 1111 15012 1111 5 OR
rlabel metal2 14640 1111 14652 1111 5 AND
rlabel metal2 13512 1111 13524 1111 5 SUB
rlabel metal2 14160 1111 14172 1111 5 nZ
rlabel metal2 14304 1111 14316 1111 5 FAOut
rlabel metal2 16728 1111 16740 1111 5 ShL
rlabel metal2 13848 1111 13860 1111 5 CIn_Slice
rlabel metal1 12942 1099 12942 1099 6 AluOut
rlabel metal2 12600 1111 12612 1111 5 Op1Sel
rlabel metal2 3192 1111 3204 1111 5 WdSel
rlabel metal2 3408 1111 3420 1111 5 Rw[0]
rlabel metal2 4152 1111 4164 1111 5 Rs1[0]
rlabel metal2 4368 1111 4380 1111 5 Rs2[0]
rlabel metal2 4560 1111 4572 1111 5 Rw[1]
rlabel metal2 5304 1111 5316 1111 5 Rs1[1]
rlabel metal2 5520 1111 5532 1111 5 Rs2[1]
rlabel metal2 5712 1111 5724 1111 5 Rw[2]
rlabel metal2 6456 1111 6468 1111 5 Rs1[2]
rlabel metal2 6672 1111 6684 1111 5 Rs2[2]
rlabel metal2 6864 1111 6876 1111 5 Rw[3]
rlabel metal2 7608 1111 7620 1111 5 Rs1[3]
rlabel metal2 7824 1111 7836 1111 5 Rs2[3]
rlabel metal2 8016 1111 8028 1111 5 Rw[4]
rlabel metal2 8760 1111 8772 1111 5 Rs1[4]
rlabel metal2 8976 1111 8988 1111 5 Rs2[4]
rlabel metal2 9168 1111 9180 1111 5 Rw[5]
rlabel metal2 10128 1111 10140 1111 5 Rs2[5]
rlabel metal2 9912 1111 9924 1111 5 Rs1[5]
rlabel metal2 10320 1111 10332 1111 5 Rw[6]
rlabel metal2 11064 1111 11076 1111 5 Rs1[6]
rlabel metal2 11280 1111 11292 1111 5 Rs2[6]
rlabel metal2 11472 1111 11484 1111 5 Rw[7]
rlabel metal2 12216 1111 12228 1111 5 Rs1[7]
rlabel metal2 12432 1111 12444 1111 5 Rs2[7]
rlabel metal2 3024 1111 3036 1111 5 PcEn
rlabel metal2 1872 1111 1884 1111 5 PcSel[1]
rlabel metal2 1488 1111 1500 1111 5 PcSel[0]
rlabel metal2 1320 1111 1332 1111 5 LrEn
rlabel metal2 576 1111 588 1111 5 LrWe
rlabel metal2 360 1111 372 1111 5 LrSel
rlabel metal2 216 1111 228 1111 5 PcIncCout
rlabel metal2 2280 1111 2292 1111 5 PcWe
rlabel metal2 2064 1111 2076 1111 5 PcSel[2]
rlabel metal1 12577 970 12577 970 1 Rd1
rlabel metal1 12579 948 12579 948 1 Rd2
rlabel metal2 3294 988 3294 988 1 WData
rlabel metal1 20472 29 20472 39 7 SysBus
rlabel metal1 12925 33 12925 33 1 SysBus
rlabel metal1 12544 34 12544 34 1 SysBus
rlabel metal1 3288 34 3288 34 1 SysBus
rlabel metal1 0 29 0 39 1 SysBus
rlabel metal2 13032 0 13044 0 1 Op2Sel[1]
rlabel metal2 17112 0 17124 0 1 Sh8G_L
rlabel metal2 17064 0 17076 0 1 Sh8F_L
rlabel metal2 17016 0 17028 0 1 Sh8E_L
rlabel metal2 16968 0 16980 0 1 Sh8D_L
rlabel metal2 18360 0 18372 0 1 Sh1_L_In
rlabel metal2 18600 0 18612 0 1 Sh8Z_R
rlabel metal2 18648 0 18660 0 1 Sh8A_R
rlabel metal2 18696 0 18708 0 1 Sh8B_R
rlabel metal2 17616 0 17628 0 1 Sh4D_L
rlabel metal2 17568 0 17580 0 1 Sh4C_L
rlabel metal2 17520 0 17532 0 1 Sh4B_L
rlabel metal2 17976 0 17988 0 1 Sh2C_L
rlabel metal2 17928 0 17940 0 1 Sh2B_L
rlabel metal2 18553 0 18565 0 1 ShR
rlabel metal2 18528 0 18540 0 1 Sh8
rlabel metal2 17472 0 17484 0 1 Sh4A_L
rlabel metal2 17160 0 17172 0 1 Sh8H_L
rlabel metal2 20064 0 20076 0 1 Sh1_R_Out
rlabel metal2 19752 0 19764 0 1 Sh2A_R
rlabel metal2 19704 0 19716 0 1 Sh2Z_R
rlabel metal2 19296 0 19308 0 1 Sh4Z_R
rlabel metal2 19344 0 19356 0 1 Sh4A_R
rlabel metal2 19392 0 19404 0 1 Sh4B_R
rlabel metal2 20352 0 20364 0 1 ShOut
rlabel metal2 19632 0 19644 0 1 Sh2
rlabel metal2 19992 0 20004 0 1 Sh1
rlabel metal2 19176 0 19188 0 1 Sh4
rlabel metal2 18744 0 18756 0 1 Sh8C_R
rlabel metal2 18792 0 18804 0 1 Sh8D_R
rlabel metal2 18840 0 18852 0 1 Sh8E_R
rlabel metal2 18888 0 18900 0 1 Sh8F_R
rlabel metal2 18936 0 18948 0 1 Sh8G_R
rlabel metal2 16824 0 16836 0 1 Sh8A_L
rlabel metal2 16920 0 16932 0 1 Sh8C_L
rlabel metal2 16872 0 16884 0 1 Sh8B_L
rlabel metal2 13248 0 13260 0 1 ZeroA
rlabel metal2 14304 0 14316 0 1 FAOut
rlabel metal2 13680 0 13692 0 1 CIn
rlabel metal2 14640 0 14652 0 1 AND
rlabel metal2 15000 0 15012 0 1 OR
rlabel metal2 15408 0 15420 0 1 XOR
rlabel metal2 15744 0 15756 0 1 NOT
rlabel metal2 16056 0 16068 0 1 NAND
rlabel metal2 16392 0 16404 0 1 NOR
rlabel metal2 16728 0 16740 0 1 ShL
rlabel metal2 16560 0 16572 0 1 ShB
rlabel metal2 13512 0 13524 0 1 SUB
rlabel metal2 14160 0 14172 0 1 nZ_prev
rlabel metal2 13872 0 13884 0 1 CIn_Slice
rlabel metal2 12792 0 12804 0 1 Op2Sel[0]
rlabel metal2 12600 0 12612 0 1 Op1Sel
rlabel metal2 4368 0 4380 0 1 Rs2[0]
rlabel metal2 3408 0 3420 0 1 Rw[0]
rlabel metal2 12432 0 12444 0 1 Rs2[7]
rlabel metal2 12216 0 12228 0 1 Rs1[7]
rlabel metal2 11472 0 11484 0 1 Rw[7]
rlabel metal2 11280 0 11292 0 1 Rs2[6]
rlabel metal2 11064 0 11076 0 1 Rs1[6]
rlabel metal2 10320 0 10332 0 1 Rw[6]
rlabel metal2 10128 0 10140 0 1 Rs2[5]
rlabel metal2 9912 0 9924 0 1 Rs1[5]
rlabel metal2 9168 0 9180 0 1 Rw[5]
rlabel metal2 8976 0 8988 0 1 Rs2[4]
rlabel metal2 8760 0 8772 0 1 Rs1[4]
rlabel metal2 8016 0 8028 0 1 Rw[4]
rlabel metal2 7824 0 7836 0 1 Rs2[3]
rlabel metal2 7608 0 7620 0 1 Rs1[3]
rlabel metal2 6864 0 6876 0 1 Rw[3]
rlabel metal2 6672 0 6684 0 1 Rs2[2]
rlabel metal2 6456 0 6468 0 1 Rs1[2]
rlabel metal2 5712 0 5724 0 1 Rw[2]
rlabel metal2 5520 0 5532 0 1 Rs2[1]
rlabel metal2 5304 0 5316 0 1 Rs1[1]
rlabel metal2 4560 0 4572 0 1 Rw[1]
rlabel metal2 4152 0 4164 0 1 Rs1[0]
rlabel metal2 3192 0 3204 0 1 WdSel
rlabel metal2 3024 0 3036 0 1 PcEn
rlabel metal2 2280 0 2292 0 1 PcWe
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 2064 0 2076 0 1 PcSel[2]
rlabel metal2 19248 0 19260 0 1 Sh4Y_R
rlabel metal1 12546 70 12546 70 1 Pc
rlabel metal1 12545 12 12545 12 1 Imm
rlabel metal1 0 7 0 17 1 Imm
rlabel metal2 12702 105 12702 105 1 A
rlabel metal2 13134 105 13134 105 1 B
<< end >>
