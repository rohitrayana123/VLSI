magic
tech c035u
timestamp 1394477235
<< checkpaint >>
rect -1228 1340 2176 2371
rect -1300 1338 2176 1340
rect -1300 -1318 2308 1338
rect -1228 -1340 2308 -1318
rect -1228 -1411 2176 -1340
<< metal1 >>
rect 805 892 935 902
rect 757 870 887 880
rect 0 50 599 60
rect 0 -16 23 -6
rect 37 -16 1008 -6
rect 973 -38 1008 -28
<< m2contact >>
rect 791 890 805 904
rect 935 890 949 904
rect 743 868 757 882
rect 887 868 901 882
rect 599 48 613 62
rect 23 -18 37 -4
rect 959 -40 973 -26
<< metal2 >>
rect 72 865 84 1065
rect 744 882 756 1065
rect 792 904 804 1065
rect 744 865 756 868
rect 792 865 804 890
rect 864 865 876 1065
rect 888 865 900 868
rect 936 865 948 890
rect 24 -4 36 66
rect 72 -111 84 66
rect 600 62 612 66
rect 744 -111 756 66
rect 792 -111 804 66
rect 864 -111 876 66
rect 960 -26 972 66
use scanreg  scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 66
box 0 0 720 799
use rowcrosser  rowcrosser_0
timestamp 1386086759
transform 1 0 720 0 1 66
box 0 0 48 799
use rowcrosser  rowcrosser_1
timestamp 1386086759
transform 1 0 768 0 1 66
box 0 0 48 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 816 0 1 66
box 0 0 192 799
<< labels >>
rlabel metal1 0 50 0 60 3 Ir
rlabel metal1 1008 -38 1008 -28 7 Imm
rlabel metal1 1008 -16 1008 -6 7 SysBus
rlabel metal1 0 -16 0 -6 3 SysBus
rlabel metal2 72 -111 84 -111 1 IrWe
rlabel metal2 744 -111 756 -111 1 Ext0
rlabel metal2 792 -111 804 -111 1 Ext1
rlabel metal2 864 -111 876 -111 1 ImmSel
rlabel metal2 864 1065 876 1065 5 ImmSel
rlabel metal2 792 1065 804 1065 5 Ext1
rlabel metal2 744 1065 756 1065 5 Ext0
rlabel metal2 72 1065 84 1065 5 IrWe
<< end >>
