magic
tech c035u
timestamp 1394562612
<< metal1 >>
rect 481 21074 16460 21084
rect 16474 21074 23884 21084
rect 504 21050 16580 21060
rect 16594 21050 23884 21060
rect 527 21026 16700 21036
rect 16714 21026 23884 21036
rect 550 21002 16820 21012
rect 16834 21002 23884 21012
rect 573 20978 16940 20988
rect 16954 20978 23884 20988
rect 596 20954 4148 20964
rect 4162 20954 23884 20964
rect 619 20930 4580 20940
rect 4594 20930 23884 20940
rect 642 20906 5012 20916
rect 5026 20906 23884 20916
rect 665 20882 4196 20892
rect 4210 20882 23884 20892
rect 688 20858 4628 20868
rect 4642 20858 23884 20868
rect 711 20834 5060 20844
rect 5074 20834 23884 20844
rect 734 20810 7148 20820
rect 7162 20810 23884 20820
rect 757 20786 7124 20796
rect 7138 20786 22580 20796
rect 22594 20786 23884 20796
rect 780 20762 7100 20772
rect 7114 20762 22796 20772
rect 22810 20762 23884 20772
rect 803 20738 22916 20748
rect 22930 20738 23884 20748
rect 826 20714 23036 20724
rect 23050 20714 23884 20724
rect 0 17893 467 17903
rect 481 17893 832 17903
rect 0 17861 832 17871
rect 0 17827 832 17837
rect 0 16717 490 16727
rect 504 16717 832 16727
rect 0 16685 832 16695
rect 0 16651 832 16661
rect 0 15541 513 15551
rect 527 15541 832 15551
rect 0 15509 832 15519
rect 0 15475 832 15485
rect 0 14365 536 14375
rect 550 14365 832 14375
rect 0 14333 832 14343
rect 0 14299 832 14309
rect 0 13189 559 13199
rect 573 13189 832 13199
rect 0 13157 832 13167
rect 0 13123 832 13133
rect 0 12013 582 12023
rect 596 12013 832 12023
rect 0 11981 832 11991
rect 0 11947 832 11957
rect 0 10837 605 10847
rect 619 10837 832 10847
rect 0 10805 832 10815
rect 0 10771 832 10781
rect 0 9661 628 9671
rect 642 9661 832 9671
rect 0 9629 832 9639
rect 0 9595 832 9605
rect 0 8485 651 8495
rect 665 8485 832 8495
rect 0 8453 832 8463
rect 0 8419 832 8429
rect 0 7309 674 7319
rect 688 7309 832 7319
rect 0 7277 832 7287
rect 0 7243 832 7253
rect 0 6133 697 6143
rect 711 6133 832 6143
rect 0 6101 832 6111
rect 0 6067 832 6077
rect 0 4957 720 4967
rect 734 4957 832 4967
rect 0 4925 832 4935
rect 0 4891 832 4901
rect 0 3781 743 3791
rect 757 3781 832 3791
rect 0 3749 832 3759
rect 0 3715 832 3725
rect 0 2605 766 2615
rect 780 2605 832 2615
rect 0 2573 832 2583
rect 0 2539 832 2549
rect 0 1429 789 1439
rect 803 1429 832 1439
rect 0 1397 832 1407
rect 0 1363 832 1373
rect 0 253 812 263
rect 826 253 832 263
rect 0 221 832 231
rect 0 187 832 197
rect 2522 72 3740 82
rect 3754 72 17252 82
rect 17266 72 19916 82
rect 19930 72 19963 82
rect 19977 72 20012 82
rect 20026 72 20060 82
rect 20074 72 20108 82
rect 20122 72 20156 82
rect 20170 72 20204 82
rect 20218 72 20252 82
rect 20266 72 20564 82
rect 20578 72 20612 82
rect 20626 72 20659 82
rect 20673 72 20708 82
rect 20722 72 21020 82
rect 21034 72 21068 82
rect 21082 72 21452 82
rect 21466 72 24093 82
<< m2contact >>
rect 467 21072 481 21086
rect 16460 21073 16474 21087
rect 490 21048 504 21062
rect 16580 21048 16594 21062
rect 513 21024 527 21038
rect 16700 21024 16714 21038
rect 536 21000 550 21014
rect 16820 21000 16834 21014
rect 559 20976 573 20990
rect 16940 20976 16954 20990
rect 582 20952 596 20966
rect 4148 20952 4162 20966
rect 605 20928 619 20942
rect 4580 20928 4594 20942
rect 628 20904 642 20918
rect 5012 20904 5026 20918
rect 651 20880 665 20894
rect 4196 20880 4210 20894
rect 674 20856 688 20870
rect 4628 20856 4642 20870
rect 697 20832 711 20846
rect 5060 20832 5074 20846
rect 720 20808 734 20822
rect 7148 20808 7162 20822
rect 743 20784 757 20798
rect 7124 20784 7138 20798
rect 22580 20784 22594 20798
rect 766 20760 780 20774
rect 7100 20760 7114 20774
rect 22796 20759 22810 20773
rect 789 20736 803 20750
rect 22916 20736 22930 20750
rect 812 20712 826 20726
rect 23036 20712 23050 20726
rect 467 17891 481 17905
rect 490 16715 504 16729
rect 513 15539 527 15553
rect 536 14363 550 14377
rect 559 13187 573 13201
rect 582 12011 596 12025
rect 605 10835 619 10849
rect 628 9659 642 9673
rect 651 8483 665 8497
rect 674 7307 688 7321
rect 697 6131 711 6145
rect 720 4955 734 4969
rect 743 3779 757 3793
rect 766 2603 780 2617
rect 789 1427 803 1441
rect 812 251 826 265
rect 3740 70 3754 84
rect 17252 70 17266 84
rect 19916 70 19930 84
rect 19963 70 19977 84
rect 20012 70 20026 84
rect 20060 70 20074 84
rect 20108 70 20122 84
rect 20156 70 20170 84
rect 20204 70 20218 84
rect 20252 70 20266 84
rect 20564 70 20578 84
rect 20612 70 20626 84
rect 20659 70 20673 84
rect 20708 70 20722 84
rect 21020 70 21034 84
rect 21068 70 21082 84
rect 21452 70 21466 84
rect 24093 70 24107 84
<< metal2 >>
rect 468 17905 480 21072
rect 491 16729 503 21048
rect 514 15553 526 21024
rect 537 14377 549 21000
rect 560 13201 572 20976
rect 583 12025 595 20952
rect 606 10849 618 20928
rect 629 9673 641 20904
rect 652 8497 664 20880
rect 675 7321 687 20856
rect 698 6145 710 20832
rect 721 4969 733 20808
rect 744 3793 756 20784
rect 767 2617 779 20760
rect 790 1441 802 20736
rect 813 265 825 20712
rect 837 20703 1037 21230
rect 1053 20703 1065 21230
rect 1077 20703 1089 21230
rect 1101 20703 1113 21230
rect 1125 20703 1137 21230
rect 4125 20703 4137 21230
rect 4149 20703 4161 20952
rect 4197 20703 4209 20880
rect 4365 20703 4377 21230
rect 4581 20703 4593 20928
rect 4629 20703 4641 20856
rect 5013 20703 5025 20904
rect 5061 20703 5073 20832
rect 5421 20703 5433 21230
rect 5661 20703 5673 21230
rect 6791 20703 6803 21230
rect 7101 20703 7113 20760
rect 7125 20703 7137 20784
rect 7149 20703 7161 20808
rect 16461 20703 16473 21073
rect 16581 20703 16593 21048
rect 16701 20703 16713 21024
rect 16821 20703 16833 21000
rect 16941 20703 16953 20976
rect 18117 20703 18129 21230
rect 18549 20703 18561 21230
rect 18741 20703 18753 21230
rect 18813 20703 18825 21230
rect 18909 20703 18921 21230
rect 22581 20703 22593 20784
rect 22797 20703 22809 20759
rect 22917 20703 22929 20736
rect 23037 20703 23049 20712
rect 23421 20703 23433 21230
rect 24093 20703 24293 21230
rect 837 0 1037 92
rect 1053 0 1065 92
rect 1077 0 1089 92
rect 1101 0 1113 92
rect 1125 0 1137 92
rect 2397 0 2409 92
rect 2589 0 2601 92
rect 3381 0 3393 92
rect 3741 84 3753 92
rect 3885 0 3897 92
rect 4101 0 4113 92
rect 4845 0 4857 92
rect 5013 0 5025 92
rect 5397 0 5409 92
rect 5613 0 5625 92
rect 6357 0 6369 92
rect 6525 0 6537 92
rect 15933 0 15945 92
rect 16125 0 16137 92
rect 16773 83 16785 92
rect 16965 83 16977 92
rect 17253 84 17265 92
rect 19917 84 19929 92
rect 19965 84 19977 92
rect 20013 84 20025 92
rect 20061 84 20073 92
rect 20109 84 20121 92
rect 20157 84 20169 92
rect 20205 84 20217 92
rect 20253 84 20265 92
rect 20565 84 20577 92
rect 20613 84 20625 92
rect 20661 84 20673 92
rect 20709 84 20721 92
rect 21021 84 21033 92
rect 21069 84 21081 92
rect 21453 84 21465 92
rect 16773 71 16977 83
rect 23853 0 23865 92
rect 24093 84 24293 92
rect 24107 70 24293 84
rect 24093 0 24293 70
use slice17 slice17_0
timestamp 1394562424
transform 1 0 837 0 1 18908
box 0 0 23456 1795
use leftbuf_slice leftbuf_slice_0
array 0 0 1685 0 15 1176
timestamp 1394551156
transform 1 0 832 0 1 98
box 0 -6 1685 1170
use IrAA IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 2517 0 1 9611
box 0 -111 1008 1065
use LLIcell_U LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1393855556
transform 1 0 23565 0 1 9611
box 0 0 192 1042
use IrBA IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 2517 0 1 6083
box 0 -111 1008 1065
use IrBB IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 2517 0 1 204
box 0 -112 1008 1064
use LLIcell_L LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23565 0 1 203
box 0 0 192 1042
use Datapath_slice Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394556877
transform 1 0 3525 0 1 92
box 0 0 20768 1176
<< labels >>
rlabel metal1 0 187 0 197 3 SysBus[0]
rlabel metal1 0 1363 0 1373 3 SysBus[1]
rlabel metal1 0 2539 0 2549 3 SysBus[2]
rlabel metal1 0 3715 0 3725 3 SysBus[3]
rlabel metal1 0 4891 0 4901 3 SysBus[4]
rlabel metal1 0 6067 0 6077 3 SysBus[5]
rlabel metal1 0 7243 0 7253 3 SysBus[6]
rlabel metal1 0 8419 0 8429 3 SysBus[7]
rlabel metal1 0 9595 0 9605 3 SysBus[8]
rlabel metal1 0 10771 0 10781 3 SysBus[9]
rlabel metal1 0 11947 0 11957 3 SysBus[10]
rlabel metal1 0 13123 0 13133 3 SysBus[11]
rlabel metal1 0 14299 0 14309 3 SysBus[12]
rlabel metal1 0 15475 0 15485 3 SysBus[13]
rlabel metal1 0 16651 0 16661 3 SysBus[14]
rlabel metal1 0 17827 0 17837 3 SysBus[15]
rlabel metal1 0 253 0 263 3 Ir[0]
rlabel metal1 0 1429 0 1439 3 Ir[1]
rlabel metal1 0 2605 0 2615 3 Ir[2]
rlabel metal1 0 3781 0 3791 3 Ir[3]
rlabel metal1 0 4957 0 4967 3 Ir[4]
rlabel metal1 0 6133 0 6143 3 Ir[5]
rlabel metal1 0 7309 0 7319 3 Ir[6]
rlabel metal1 0 8485 0 8495 3 Ir[7]
rlabel metal1 0 9661 0 9671 3 Ir[8]
rlabel metal1 0 10837 0 10847 3 Ir[9]
rlabel metal1 0 12013 0 12023 3 Ir[10]
rlabel metal1 0 13189 0 13199 3 Ir[11]
rlabel metal1 0 14365 0 14375 3 Ir[12]
rlabel metal1 0 15541 0 15551 3 Ir[13]
rlabel metal1 0 16717 0 16727 3 Ir[14]
rlabel metal1 0 17893 0 17903 3 Ir[15]
rlabel metal2 837 0 1037 0 1 Vdd!
rlabel metal2 1053 0 1065 0 1 SDI
rlabel metal2 1077 0 1089 0 1 Test
rlabel metal2 1101 0 1113 0 1 Clock
rlabel metal2 1125 0 1137 0 1 nReset
rlabel metal2 750 20781 750 20781 1 Ir[3]
rlabel metal2 727 20782 727 20782 1 Ir[4]
rlabel metal2 704 20781 704 20781 1 Ir[5]
rlabel metal2 681 20780 681 20780 1 Ir[6]
rlabel metal2 658 20779 658 20779 1 Ir[7]
rlabel metal2 635 20777 635 20777 1 Ir[8]
rlabel metal2 612 20777 612 20777 1 Ir[9]
rlabel metal2 589 20776 589 20776 1 Ir[10]
rlabel metal2 566 20777 566 20777 1 Ir[11]
rlabel metal2 543 20777 543 20777 1 Ir[12]
rlabel metal2 520 20776 520 20776 1 Ir[13]
rlabel metal2 497 20776 497 20776 1 Ir[14]
rlabel metal2 473 20777 473 20777 1 Ir[15]
rlabel metal2 1053 21230 1065 21230 1 SDI
rlabel metal2 1077 21230 1089 21230 1 Test
rlabel metal2 1101 21230 1113 21230 1 Clock
rlabel metal2 1125 21230 1137 21230 1 nReset
rlabel metal2 837 21230 1037 21230 5 Vdd!
rlabel metal2 3885 0 3897 0 1 LrSel
rlabel metal2 4101 0 4113 0 1 LrWe
rlabel metal2 4845 0 4857 0 1 LrEn
rlabel metal2 5013 0 5025 0 1 PcSel[0]
rlabel metal2 5397 0 5409 0 1 PcSel[1]
rlabel metal2 5613 0 5625 0 1 PcWe
rlabel metal2 6357 0 6369 0 1 PcEn
rlabel metal2 6525 0 6537 0 1 WdSel
rlabel metal2 16125 0 16137 0 1 Op2Sel
rlabel metal2 15933 0 15945 0 1 Op1Sel
rlabel metal2 24093 0 24293 0 1 GND!
rlabel metal2 23853 0 23865 0 1 AluEn
rlabel metal2 3381 0 3393 0 1 ImmSel
rlabel metal2 2589 0 2601 0 1 IrWe
rlabel metal2 6791 21230 6803 21230 5 RegWe
rlabel metal2 18117 21230 18129 21230 5 CFlag
rlabel metal2 18549 21230 18561 21230 5 Flags[2]
rlabel metal2 18741 21230 18753 21230 5 Flags[1]
rlabel metal2 18813 21230 18825 21230 5 Flags[3]
rlabel metal2 23421 21230 23433 21230 5 AluEn
rlabel metal2 24093 21230 24293 21230 1 GND!
rlabel metal2 18909 21230 18921 21230 5 Flags[0]
rlabel metal2 7105 20752 7105 20752 1 Ir[2]
rlabel metal2 7131 20776 7131 20776 1 Ir[3]
rlabel metal2 7154 20800 7154 20800 1 Ir[4]
rlabel metal2 16466 21066 16466 21066 1 Ir[15]
rlabel metal2 16585 21041 16585 21041 1 Ir[14]
rlabel metal2 16706 21018 16706 21018 1 Ir[13]
rlabel metal2 16827 20994 16827 20994 1 Ir[12]
rlabel metal2 16947 20969 16947 20969 1 Ir[11]
rlabel metal2 22587 20779 22587 20779 1 Ir[3]
rlabel metal2 22802 20754 22802 20754 1 Ir[2]
rlabel metal2 22922 20729 22922 20729 1 Ir[1]
rlabel metal2 23043 20707 23043 20707 1 Ir[0]
rlabel metal1 0 221 0 231 3 DataIn[0]
rlabel metal1 0 17861 0 17871 3 DataIn[15]
rlabel metal1 0 16685 0 16695 3 DataIn[14]
rlabel metal1 0 15509 0 15519 3 DataIn[13]
rlabel metal1 0 14333 0 14343 3 DataIn[12]
rlabel metal1 0 13157 0 13167 3 DataIn[11]
rlabel metal1 0 11981 0 11991 3 DataIn[10]
rlabel metal1 0 10805 0 10815 3 DataIn[9]
rlabel metal1 0 9629 0 9639 3 DataIn[8]
rlabel metal1 0 8453 0 8463 3 DataIn[7]
rlabel metal1 0 7277 0 7287 3 DataIn[6]
rlabel metal1 0 6101 0 6111 3 DataIn[5]
rlabel metal1 0 4925 0 4935 3 DataIn[4]
rlabel metal1 0 3749 0 3759 3 DataIn[3]
rlabel metal1 0 2573 0 2583 3 DataIn[2]
rlabel metal1 0 1397 0 1407 3 DataIn[1]
rlabel metal2 2397 0 2409 0 1 MemEn
rlabel metal2 4125 21230 4137 21230 5 Rs1Sel[0]
rlabel metal2 4365 21230 4377 21230 5 Rs1Sel[1]
rlabel metal1 4606 20959 4606 20959 1 Ir[10]
rlabel metal2 5421 21230 5433 21230 5 RwSel[0]
rlabel metal2 5661 21230 5673 21230 5 RwSel[1]
rlabel metal2 4154 20945 4154 20945 1 Ir[10]
rlabel metal2 4203 20872 4203 20872 1 Ir[7]
rlabel metal2 4586 20920 4586 20920 1 Ir[9]
rlabel metal2 4635 20849 4635 20849 1 Ir[6]
rlabel metal2 5018 20897 5018 20897 1 Ir[8]
rlabel metal2 5068 20826 5068 20826 1 Ir[5]
<< end >>
