magic
tech c035u
timestamp 1394841956
<< nwell >>
rect 0 467 192 865
<< pwell >>
rect 0 66 192 467
<< pohmic >>
rect 0 142 6 152
rect 186 142 192 152
<< nohmic >>
rect 0 802 6 812
rect 186 802 192 812
<< psubstratetap >>
rect 6 142 186 158
<< nsubstratetap >>
rect 6 796 186 812
<< metal1 >>
rect 0 848 192 858
rect 0 825 192 835
rect 0 796 6 812
rect 186 796 192 812
rect 0 787 192 796
rect 0 158 192 167
rect 0 142 6 158
rect 186 142 192 158
rect 0 119 192 129
rect 0 96 192 106
rect 0 73 192 83
rect 0 51 192 61
<< metal2 >>
rect 48 0 60 1042
<< labels >>
rlabel metal2 48 0 60 0 1 LLI
rlabel metal1 0 787 0 812 1 Vdd!
rlabel metal1 0 825 0 835 1 Scan
rlabel metal1 0 848 0 858 1 ScanReturn
rlabel metal1 192 848 192 858 7 ScanReturn
rlabel metal2 48 1042 60 1042 5 LLI
rlabel metal1 0 51 0 61 3 ALUOut
rlabel metal1 192 51 192 61 7 ALUOut
rlabel metal1 192 142 192 167 7 GND!
rlabel metal1 192 119 192 129 7 Clock
rlabel metal1 192 96 192 106 7 Test
rlabel metal1 192 73 192 83 7 nReset
rlabel metal1 0 142 0 167 1 GND!
rlabel metal1 0 119 0 129 1 Clock
rlabel metal1 0 96 0 106 1 Test
rlabel metal1 0 73 0 83 1 nReset
rlabel metal1 192 787 192 812 7 Vdd!
rlabel metal1 192 825 192 835 7 Scan
<< end >>
