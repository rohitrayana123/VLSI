magic
tech c035u
timestamp 1394841445
<< nwell >>
rect 1464 958 3480 1356
rect 15288 958 15912 1356
rect 23566 958 24336 1356
<< pwell >>
rect 1464 557 3480 958
rect 15288 564 15912 958
rect 23566 557 24336 958
<< pohmic >>
rect 1464 633 1470 643
rect 3474 633 3480 643
rect 15288 633 15294 643
rect 15906 633 15912 643
rect 23566 633 23572 643
rect 24330 633 24336 643
<< nohmic >>
rect 1464 1293 1470 1303
rect 3474 1293 3480 1303
rect 15288 1293 15294 1303
rect 15906 1293 15912 1303
rect 23566 1293 23572 1303
rect 24330 1293 24336 1303
<< psubstratetap >>
rect 1470 633 3474 649
rect 15294 633 15906 649
rect 23572 633 24330 649
<< nsubstratetap >>
rect 1470 1287 3474 1303
rect 15294 1287 15906 1303
rect 23572 1287 24330 1303
<< metal1 >>
rect 3877 1751 6407 1761
rect 13501 1757 16535 1767
rect 4309 1729 6383 1739
rect 13309 1735 16415 1745
rect 4741 1707 6359 1717
rect 13117 1713 16295 1723
rect 5173 1684 6143 1694
rect 12925 1691 16175 1701
rect 5605 1663 6119 1673
rect 12733 1669 16055 1679
rect 6037 1641 6095 1651
rect 12541 1647 15935 1657
rect 4429 1537 5759 1547
rect 4477 1515 5711 1525
rect 4045 1493 5279 1503
rect 3997 1471 5327 1481
rect 3612 1449 4847 1459
rect 3565 1427 4895 1437
rect 3541 1405 3959 1415
rect 3973 1405 4391 1415
rect 4837 1405 5255 1415
rect 5269 1405 5687 1415
rect 3781 1383 4199 1393
rect 4213 1383 4631 1393
rect 5077 1383 5495 1393
rect 5509 1383 5927 1393
rect 3637 1361 3791 1371
rect 4069 1361 4223 1371
rect 4501 1361 4655 1371
rect 4933 1361 5087 1371
rect 5365 1361 5519 1371
rect 5797 1361 5951 1371
rect 1464 1339 3480 1349
rect 15288 1339 15912 1349
rect 23566 1339 24336 1349
rect 1464 1316 3480 1326
rect 15288 1316 15912 1326
rect 23566 1316 24336 1326
rect 1464 1287 1470 1303
rect 3474 1287 3480 1303
rect 1464 1278 3480 1287
rect 15288 1287 15294 1303
rect 15906 1287 15912 1303
rect 15288 1278 15912 1287
rect 23566 1287 23572 1303
rect 24330 1287 24336 1303
rect 23566 1278 24336 1287
rect 1464 649 3480 658
rect 1464 633 1470 649
rect 3474 633 3480 649
rect 15288 649 15912 658
rect 15288 633 15294 649
rect 15906 633 15912 649
rect 23566 649 24336 658
rect 23566 633 23572 649
rect 24330 633 24336 649
rect 1464 610 3480 620
rect 15288 610 15912 620
rect 1464 587 3480 597
rect 15288 587 15912 597
rect 1464 564 3480 574
rect 15288 564 15912 574
rect 21349 28 21383 38
rect 21397 28 21431 38
rect 21445 28 21479 38
rect 21493 28 21527 38
rect 21541 28 21575 38
rect 21589 28 21623 38
rect 21637 28 21671 38
rect 21685 28 21983 38
rect 21997 28 22031 38
rect 22045 28 22079 38
rect 22093 28 22127 38
rect 22141 28 22439 38
rect 22453 28 22487 38
rect 22501 28 22799 38
<< m2contact >>
rect 3863 1749 3877 1763
rect 6407 1749 6421 1763
rect 13487 1756 13501 1770
rect 16535 1755 16549 1769
rect 4295 1727 4309 1741
rect 6383 1727 6397 1741
rect 13295 1733 13309 1747
rect 16415 1733 16429 1747
rect 4727 1705 4741 1719
rect 6359 1705 6373 1719
rect 13103 1711 13117 1725
rect 16295 1711 16309 1725
rect 5159 1682 5173 1696
rect 6143 1682 6157 1696
rect 12911 1689 12925 1703
rect 16175 1689 16189 1703
rect 5591 1660 5605 1674
rect 6119 1660 6133 1674
rect 12719 1667 12733 1681
rect 16055 1667 16069 1681
rect 6023 1639 6037 1653
rect 6095 1638 6109 1652
rect 12527 1645 12541 1659
rect 15935 1645 15949 1659
rect 4415 1535 4429 1549
rect 5759 1535 5773 1549
rect 4463 1513 4477 1527
rect 5711 1513 5725 1527
rect 4031 1491 4045 1505
rect 5279 1491 5293 1505
rect 3983 1469 3997 1483
rect 5327 1469 5341 1483
rect 3598 1447 3612 1461
rect 4847 1447 4861 1461
rect 3551 1425 3565 1439
rect 4895 1425 4909 1439
rect 3527 1403 3541 1417
rect 3959 1403 3973 1417
rect 4391 1403 4405 1417
rect 4823 1403 4837 1417
rect 5255 1403 5269 1417
rect 5687 1403 5701 1417
rect 3767 1381 3781 1395
rect 4199 1381 4213 1395
rect 4631 1381 4645 1395
rect 5063 1381 5077 1395
rect 5495 1381 5509 1395
rect 5927 1381 5941 1395
rect 3623 1359 3637 1373
rect 3791 1359 3805 1373
rect 4055 1359 4069 1373
rect 4223 1359 4237 1373
rect 4487 1359 4501 1373
rect 4655 1359 4669 1373
rect 4919 1359 4933 1373
rect 5087 1359 5101 1373
rect 5351 1359 5365 1373
rect 5519 1359 5533 1373
rect 5783 1359 5797 1373
rect 5951 1359 5965 1373
rect 21335 26 21349 40
rect 21383 26 21397 40
rect 21431 26 21445 40
rect 21479 26 21493 40
rect 21527 26 21541 40
rect 21575 26 21589 40
rect 21623 26 21637 40
rect 21671 26 21685 40
rect 21983 25 21997 39
rect 22031 25 22045 39
rect 22079 25 22093 39
rect 22127 25 22141 39
rect 22439 26 22453 40
rect 22487 26 22501 40
rect 22799 26 22813 40
<< metal2 >>
rect 0 1356 200 1793
rect 216 1356 228 1793
rect 240 1356 252 1793
rect 264 1356 276 1793
rect 288 1356 300 1793
rect 3528 1417 3540 1793
rect 3552 1439 3564 1793
rect 3600 1461 3612 1793
rect 3528 1356 3540 1403
rect 3552 1356 3564 1425
rect 3600 1356 3612 1447
rect 3768 1395 3780 1793
rect 3624 1356 3636 1359
rect 3768 1356 3780 1381
rect 3792 1356 3804 1359
rect 3864 1356 3876 1749
rect 3984 1483 3996 1793
rect 4032 1505 4044 1793
rect 3960 1356 3972 1403
rect 3984 1356 3996 1469
rect 4032 1356 4044 1491
rect 4056 1356 4068 1359
rect 4200 1356 4212 1381
rect 4224 1356 4236 1359
rect 4296 1356 4308 1727
rect 4416 1549 4428 1793
rect 4392 1356 4404 1403
rect 4416 1356 4428 1535
rect 4464 1527 4476 1793
rect 4464 1356 4476 1513
rect 4488 1356 4500 1359
rect 4632 1356 4644 1381
rect 4656 1356 4668 1359
rect 4728 1356 4740 1705
rect 4824 1417 4836 1793
rect 4824 1356 4836 1403
rect 4848 1356 4860 1447
rect 4896 1356 4908 1425
rect 5064 1395 5076 1793
rect 4920 1356 4932 1359
rect 5064 1356 5076 1381
rect 5088 1356 5100 1359
rect 5160 1356 5172 1682
rect 5256 1356 5268 1403
rect 5280 1356 5292 1491
rect 5328 1356 5340 1469
rect 5352 1356 5364 1359
rect 5496 1356 5508 1381
rect 5520 1356 5532 1359
rect 5592 1356 5604 1660
rect 5688 1356 5700 1403
rect 5712 1356 5724 1513
rect 5760 1356 5772 1535
rect 5784 1356 5796 1359
rect 5928 1356 5940 1381
rect 5952 1356 5964 1359
rect 6024 1356 6036 1639
rect 6096 1635 6108 1638
rect 6120 1635 6132 1660
rect 6144 1635 6156 1682
rect 6194 1635 6206 1793
rect 6360 1635 6372 1705
rect 6384 1635 6396 1727
rect 6408 1635 6420 1749
rect 6504 1635 6516 1793
rect 6528 1635 6540 1793
rect 6552 1635 6564 1793
rect 12432 1635 12444 1793
rect 12456 1635 12468 1793
rect 12528 1635 12540 1645
rect 12648 1635 12660 1793
rect 12696 1635 12708 1793
rect 12720 1635 12732 1667
rect 12840 1635 12852 1793
rect 12912 1635 12924 1689
rect 13032 1635 13044 1793
rect 13104 1635 13116 1711
rect 13224 1635 13236 1793
rect 13296 1635 13308 1733
rect 13416 1635 13428 1793
rect 13488 1635 13500 1756
rect 15936 1529 15948 1645
rect 16056 1527 16068 1667
rect 16176 1532 16188 1689
rect 16296 1532 16308 1711
rect 16416 1532 16428 1733
rect 16536 1531 16548 1755
rect 16968 1532 16980 1793
rect 17160 1532 17172 1793
rect 17232 1532 17244 1793
rect 17328 1532 17340 1793
rect 21984 1532 21996 1793
rect 22176 1532 22188 1793
rect 22296 1532 22308 1793
rect 22416 1532 22428 1793
rect 24456 1356 24656 1793
rect 0 0 200 557
rect 216 0 228 557
rect 240 0 252 557
rect 264 0 276 557
rect 288 0 300 557
rect 3696 547 3708 557
rect 3840 547 3852 557
rect 3696 535 3852 547
rect 4128 547 4140 557
rect 4272 547 4284 557
rect 4128 535 4284 547
rect 4560 547 4572 557
rect 4704 547 4716 557
rect 4560 535 4716 547
rect 4992 547 5004 557
rect 5136 547 5148 557
rect 4992 535 5148 547
rect 5424 547 5436 557
rect 5568 547 5580 557
rect 5424 535 5580 547
rect 5856 547 5868 557
rect 6000 547 6012 557
rect 5856 535 6012 547
rect 6144 0 6156 17
rect 6888 0 6900 17
rect 7104 0 7116 17
rect 7296 0 7308 17
rect 8040 0 8052 17
rect 8256 0 8268 17
rect 8448 0 8460 17
rect 9192 0 9204 17
rect 9408 0 9420 17
rect 9600 0 9612 17
rect 10344 0 10356 17
rect 10560 0 10572 17
rect 10752 0 10764 17
rect 11496 0 11508 17
rect 11712 0 11724 17
rect 11904 0 11916 17
rect 12648 0 12660 17
rect 12864 0 12876 17
rect 13056 0 13068 17
rect 13800 0 13812 17
rect 14016 0 14028 17
rect 14208 0 14220 17
rect 14952 0 14964 17
rect 15168 0 15180 17
rect 15984 0 15996 293
rect 16248 0 16260 293
rect 16416 0 16428 293
rect 16584 0 16596 293
rect 16608 0 16620 293
rect 16680 0 16692 293
rect 16896 0 16908 293
rect 17040 0 17052 293
rect 17376 0 17388 293
rect 17736 0 17748 293
rect 18144 0 18156 293
rect 18480 0 18492 293
rect 18792 0 18804 293
rect 19128 0 19140 293
rect 19248 0 19260 293
rect 19296 0 19308 293
rect 19464 0 19476 293
rect 21264 0 21276 293
rect 21289 0 21301 293
rect 21576 40 21588 293
rect 21336 0 21348 26
rect 21384 0 21396 26
rect 21432 0 21444 26
rect 21480 0 21492 26
rect 21528 0 21540 26
rect 21576 0 21588 26
rect 21624 0 21636 26
rect 21672 0 21684 26
rect 21912 0 21924 293
rect 21984 0 21996 25
rect 22032 0 22044 25
rect 22080 0 22092 25
rect 22128 0 22140 25
rect 22368 0 22380 293
rect 22440 0 22452 26
rect 22488 0 22500 26
rect 22728 0 22740 293
rect 22800 0 22812 26
rect 23088 0 23100 293
rect 23256 0 23268 293
rect 23496 73 23508 293
rect 23496 61 24228 73
rect 24216 0 24228 61
rect 24456 0 24656 557
use leftbuf  leftbuf_1
timestamp 1386242881
transform 1 0 0 0 1 557
box 0 0 1464 799
use mux2  mux2_6
timestamp 1386235218
transform 1 0 3480 0 1 557
box 0 0 192 799
use tiehigh  tiehigh_3
timestamp 1386086759
transform 1 0 3672 0 1 557
box 0 0 48 799
use mux2  mux2_7
timestamp 1386235218
transform 1 0 3720 0 1 557
box 0 0 192 799
use mux2  mux2_8
timestamp 1386235218
transform 1 0 3912 0 1 557
box 0 0 192 799
use tiehigh  tiehigh_4
timestamp 1386086759
transform 1 0 4104 0 1 557
box 0 0 48 799
use mux2  mux2_9
timestamp 1386235218
transform 1 0 4152 0 1 557
box 0 0 192 799
use mux2  mux2_10
timestamp 1386235218
transform 1 0 4344 0 1 557
box 0 0 192 799
use tiehigh  tiehigh_5
timestamp 1386086759
transform 1 0 4536 0 1 557
box 0 0 48 799
use mux2  mux2_11
timestamp 1386235218
transform 1 0 4584 0 1 557
box 0 0 192 799
use mux2  mux2_4
timestamp 1386235218
transform 1 0 4776 0 1 557
box 0 0 192 799
use tiehigh  tiehigh_2
timestamp 1386086759
transform 1 0 4968 0 1 557
box 0 0 48 799
use mux2  mux2_5
timestamp 1386235218
transform 1 0 5016 0 1 557
box 0 0 192 799
use mux2  mux2_2
timestamp 1386235218
transform 1 0 5208 0 1 557
box 0 0 192 799
use tiehigh  tiehigh_1
timestamp 1386086759
transform 1 0 5400 0 1 557
box 0 0 48 799
use mux2  mux2_3
timestamp 1386235218
transform 1 0 5448 0 1 557
box 0 0 192 799
use mux2  mux2_1
timestamp 1386235218
transform 1 0 5640 0 1 557
box 0 0 192 799
use tiehigh  tiehigh_0
timestamp 1386086759
transform 1 0 5832 0 1 557
box 0 0 48 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 5880 0 1 557
box 0 0 192 799
use regBlock_decoder  regBlock_decoder_0
timestamp 1394802642
transform 1 0 6072 0 1 17
box 0 0 9216 1618
use ALUDecoder_new  ALUDecoder_new_0
timestamp 1394841445
transform 1 0 15912 0 1 293
box 0 0 7656 1239
use rightend  rightend_0
timestamp 1386235834
transform 1 0 24336 0 1 557
box 0 0 320 799
<< labels >>
rlabel metal1 6069 1646 6069 1646 1 Rw0
rlabel metal1 6068 1667 6068 1667 1 Rw1
rlabel metal1 6062 1689 6062 1689 1 Rw2
rlabel metal1 6064 1711 6064 1711 1 Rs10
rlabel metal1 6064 1734 6064 1734 1 Rs11
rlabel metal1 6065 1754 6065 1754 1 Rs12
rlabel metal2 21264 0 21276 0 1 Sh8
rlabel metal2 16680 0 16692 0 1 Flags[3]
rlabel metal2 15984 0 15996 0 1 ZeroA
rlabel metal2 23256 0 23268 0 1 LLI
rlabel metal2 23088 0 23100 0 1 ShOut
rlabel metal2 22368 0 22380 0 1 Sh2
rlabel metal2 21289 0 21301 0 1 ShR
rlabel metal2 22728 0 22740 0 1 Sh1
rlabel metal2 21912 0 21924 0 1 Sh4
rlabel metal2 19128 0 19140 0 1 NOR
rlabel metal2 19296 0 19308 0 1 ShB
rlabel metal2 19248 0 19260 0 1 ASign
rlabel metal2 19464 0 19476 0 1 ShL
rlabel metal2 18480 0 18492 0 1 NOT
rlabel metal2 18144 0 18156 0 1 XOR
rlabel metal2 17736 0 17748 0 1 OR
rlabel metal2 17376 0 17388 0 1 AND
rlabel metal2 17040 0 17052 0 1 FAOut
rlabel metal2 16896 0 16908 0 1 nZ
rlabel metal2 16608 0 16620 0 1 COut
rlabel metal2 16584 0 16596 0 1 LastCIn
rlabel metal2 16416 0 16428 0 1 CIn_slice
rlabel metal2 16248 0 16260 0 1 SUB
rlabel metal2 18792 0 18804 0 1 NAND
rlabel metal2 21624 0 21636 0 5 Sh8G_R
rlabel metal2 21576 0 21588 0 5 Sh8F_R
rlabel metal2 21528 0 21540 0 5 Sh8E_R
rlabel metal2 21480 0 21492 0 5 Sh8D_R
rlabel metal2 21336 0 21348 0 5 Sh8A_R
rlabel metal2 21384 0 21396 0 5 Sh8B_R
rlabel metal2 21432 0 21444 0 5 Sh8C_R
rlabel metal2 21672 0 21684 0 5 Sh8H_R
rlabel metal2 22032 0 22044 0 5 Sh4A_R
rlabel metal2 22080 0 22092 0 5 Sh4B_R
rlabel metal2 22128 0 22140 0 5 Sh4C_R
rlabel metal2 21984 0 21996 0 5 Sh4Z_R
rlabel metal2 22440 0 22452 0 5 Sh2A_R
rlabel metal2 22488 0 22500 0 5 Sh2B_R
rlabel metal2 22800 0 22812 0 1 Sh1_R_In
rlabel metal2 24216 0 24228 0 1 OutEn
rlabel metal2 24458 0 24656 0 1 GND!
rlabel metal2 6144 0 6156 0 1 Rw[0]
rlabel metal2 6888 0 6900 0 1 Rs1[0]
rlabel metal2 7104 0 7116 0 1 Rs2[0]
rlabel metal2 8256 0 8268 0 1 Rs2[1]
rlabel metal2 8448 0 8460 0 1 Rw[2]
rlabel metal2 9192 0 9204 0 1 Rs1[2]
rlabel metal2 9408 0 9420 0 1 Rs2[2]
rlabel metal2 9600 0 9612 0 1 Rw[3]
rlabel metal2 10344 0 10356 0 1 Rs1[3]
rlabel metal2 10752 0 10764 0 1 Rw[4]
rlabel metal2 11496 0 11508 0 1 Rs1[4]
rlabel metal2 11712 0 11724 0 1 Rs2[4]
rlabel metal2 11904 0 11916 0 1 Rw[5]
rlabel metal2 12648 0 12660 0 1 Rs1[5]
rlabel metal2 12864 0 12876 0 1 Rs2[5]
rlabel metal2 13056 0 13068 0 1 Rw[6]
rlabel metal2 13800 0 13812 0 1 Rs1[6]
rlabel metal2 14016 0 14028 0 1 Rs2[6]
rlabel metal2 14208 0 14220 0 1 Rw[7]
rlabel metal2 14952 0 14964 0 1 Rs1[7]
rlabel metal2 15168 0 15180 0 1 Rs2[7]
rlabel metal2 7296 0 7308 0 1 Rw[1]
rlabel metal2 8040 0 8052 0 1 Rs1[1]
rlabel metal2 10560 0 10572 0 1 Rs2[3]
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 5064 1793 5076 1793 5 RwSel[1]
rlabel metal2 4416 1793 4428 1793 5 Ir[8]
rlabel metal2 4464 1793 4476 1793 5 Ir[5]
rlabel metal2 4032 1793 4044 1793 5 Ir[6]
rlabel metal2 3984 1793 3996 1793 5 Ir[9]
rlabel metal2 3600 1793 3612 1793 5 Ir[7]
rlabel metal2 3552 1793 3564 1793 5 Ir[10]
rlabel metal2 3768 1793 3780 1793 5 Rs1Sel[1]
rlabel metal2 3528 1793 3540 1793 5 Rs1Sel[0]
rlabel metal2 6194 1793 6206 1793 5 RegWe
rlabel metal2 6552 1793 6564 1793 5 Ir[4]
rlabel metal2 6528 1793 6540 1793 5 Ir[3]
rlabel metal2 6504 1793 6516 1793 5 Ir[2]
rlabel metal2 4824 1793 4836 1793 5 RwSel[0]
rlabel metal2 240 1793 252 1793 1 Test
rlabel metal2 264 1793 276 1793 1 Clock
rlabel metal2 288 1793 300 1793 1 nReset
rlabel metal2 0 1793 200 1793 5 Vdd!
rlabel metal2 216 1793 228 1793 5 SDO
rlabel metal2 24456 1793 24656 1793 1 GND!
rlabel metal2 17328 1793 17340 1793 5 Flagss[0]
rlabel metal2 17232 1793 17244 1793 5 Flags[3]
rlabel metal2 17160 1793 17172 1793 5 Flags[1]
rlabel metal2 16968 1793 16980 1793 5 Flags[2]
rlabel metal2 21984 1793 21996 1793 5 Ir[3]
rlabel metal2 22176 1793 22188 1793 5 Ir[2]
rlabel metal2 22296 1793 22308 1793 5 Ir[1]
rlabel metal2 22416 1793 22428 1793 5 Ir[0]
rlabel metal2 12432 1793 12444 1793 1 AluOR[1]
rlabel metal2 12456 1793 12468 1793 5 Ir[15]
rlabel metal2 12648 1793 12660 1793 5 Ir[14]
rlabel metal2 12696 1793 12708 1793 1 AluOR[0]
rlabel metal2 12840 1793 12852 1793 5 Ir[13]
rlabel metal2 13032 1793 13044 1793 5 Ir[12]
rlabel metal2 13224 1793 13236 1793 5 Ir[11]
rlabel metal2 13416 1793 13428 1793 5 Cin
<< end >>
