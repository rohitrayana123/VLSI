magic
tech c035u
timestamp 1394190327
<< metal1 >>
rect 0 16206 48 16216
rect 0 16168 48 16193
rect 0 15523 48 15548
rect 0 15500 48 15510
rect 0 15477 48 15487
rect 0 15454 48 15464
rect 0 15422 48 15432
rect 0 15402 48 15412
rect 1056 15402 1121 15412
rect 0 15183 48 15193
rect 0 15145 48 15170
rect 0 14500 48 14525
rect 0 14477 48 14487
rect 0 14454 48 14464
rect 0 14431 48 14441
rect 0 14399 48 14409
rect 0 14379 48 14389
rect 1056 14379 1121 14389
rect 0 14160 48 14170
rect 0 14122 48 14147
rect 0 13477 48 13502
rect 0 13454 48 13464
rect 0 13431 48 13441
rect 0 13408 48 13418
rect 0 13376 48 13386
rect 0 13356 48 13366
rect 1056 13356 1121 13366
rect 0 13137 48 13147
rect 0 13099 48 13124
rect 0 12454 48 12479
rect 0 12431 48 12441
rect 0 12408 48 12418
rect 0 12385 48 12395
rect 0 12353 48 12363
rect 0 12333 48 12343
rect 1056 12333 1121 12343
rect 0 12114 48 12124
rect 0 12076 48 12101
rect 0 11431 48 11456
rect 0 11408 48 11418
rect 0 11385 48 11395
rect 0 11362 48 11372
rect 0 11330 48 11340
rect 0 11310 48 11320
rect 1056 11310 1121 11320
rect 0 11091 48 11101
rect 0 11053 48 11078
rect 0 10408 48 10433
rect 0 10385 48 10395
rect 0 10362 48 10372
rect 0 10339 48 10349
rect 0 10307 48 10317
rect 0 10287 48 10297
rect 1056 10287 1121 10297
rect 0 10068 48 10078
rect 0 10030 48 10055
rect 0 9385 48 9410
rect 0 9362 48 9372
rect 0 9339 48 9349
rect 0 9316 48 9326
rect 0 9284 48 9294
rect 0 9264 48 9274
rect 1056 9264 1121 9274
rect 0 9045 48 9055
rect 0 9007 48 9032
rect 0 8362 48 8387
rect 0 8339 48 8349
rect 0 8316 48 8326
rect 0 8293 48 8303
rect 0 8261 48 8271
rect 0 8241 48 8251
rect 1056 8241 1121 8251
rect 0 8022 48 8032
rect 0 7984 48 8009
rect 0 7339 48 7364
rect 0 7316 48 7326
rect 0 7293 48 7303
rect 0 7270 48 7280
rect 0 7238 48 7248
rect 0 7218 48 7228
rect 1056 7218 1121 7228
rect 0 6999 48 7009
rect 0 6961 48 6986
rect 0 6316 48 6341
rect 0 6293 48 6303
rect 0 6270 48 6280
rect 0 6247 48 6257
rect 0 6215 48 6225
rect 0 6195 48 6205
rect 1056 6195 1121 6205
rect 0 5976 48 5986
rect 0 5938 48 5963
rect 0 5293 48 5318
rect 0 5270 48 5280
rect 0 5247 48 5257
rect 0 5224 48 5234
rect 0 5192 48 5202
rect 0 5172 48 5182
rect 1056 5172 1121 5182
rect 0 4953 48 4963
rect 0 4915 48 4940
rect 0 4270 48 4295
rect 0 4247 48 4257
rect 0 4224 48 4234
rect 0 4201 48 4211
rect 0 4169 48 4179
rect 0 4149 48 4159
rect 1056 4149 1121 4159
rect 0 3930 48 3940
rect 0 3892 48 3917
rect 0 3247 48 3272
rect 0 3224 48 3234
rect 0 3201 48 3211
rect 0 3178 48 3188
rect 0 3146 48 3156
rect 0 3126 48 3136
rect 1056 3126 1121 3136
rect 0 2907 48 2917
rect 0 2869 48 2894
rect 0 2224 48 2249
rect 0 2201 48 2211
rect 0 2178 48 2188
rect 0 2155 48 2165
rect 0 2123 48 2133
rect 0 2103 48 2113
rect 1056 2103 1121 2113
rect 0 1884 48 1894
rect 0 1846 48 1871
rect 0 1201 48 1226
rect 0 1178 48 1188
rect 0 1155 48 1165
rect 0 1132 48 1142
rect 0 1100 48 1110
rect 0 1080 48 1090
rect 1056 1080 1121 1090
rect 0 861 48 871
rect 0 823 48 848
rect 0 178 48 203
rect 0 155 48 165
rect 0 132 48 142
rect 0 109 48 119
rect 0 77 48 87
rect 0 57 48 67
rect 1056 57 1121 67
<< metal2 >>
rect 120 16368 132 16419
rect 912 16368 924 16419
use IrAA IrAA_0
array 0 0 1008 0 7 1023
timestamp 1394146470
transform 1 0 48 0 1 8184
box 0 0 1008 1023
use IrBA IrBA_0
array 0 0 1008 0 2 1023
timestamp 1394190290
transform 1 0 48 0 1 5115
box 0 0 1008 1023
use IrBB IrBB_0
array 0 0 1008 0 4 1023
timestamp 1394190216
transform 1 0 48 0 1 0
box 0 0 1008 1023
<< labels >>
rlabel metal1 0 823 0 848 3 Vdd!
rlabel metal1 0 178 0 203 3 GND!
rlabel metal1 0 155 0 165 3 Clock
rlabel metal1 0 132 0 142 3 Test
rlabel metal1 0 109 0 119 3 nReset
rlabel metal1 0 77 0 87 3 IrIn[0]
rlabel metal1 0 57 0 67 3 Ir[0]
rlabel metal1 0 861 0 871 3 SDI
rlabel metal1 0 1132 0 1142 3 nReset
rlabel metal1 0 1155 0 1165 3 Test
rlabel metal1 0 1178 0 1188 3 Clock
rlabel metal1 0 1201 0 1226 3 GND!
rlabel metal1 0 1846 0 1871 3 Vdd!
rlabel metal1 0 1884 0 1894 3 SDI
rlabel metal1 0 15454 0 15464 3 nReset
rlabel metal1 0 15477 0 15487 3 Test
rlabel metal1 0 15500 0 15510 3 Clock
rlabel metal1 0 15523 0 15548 3 GND!
rlabel metal1 0 16168 0 16193 3 Vdd!
rlabel metal1 0 16206 0 16216 3 SDI
rlabel metal1 0 14431 0 14441 3 nReset
rlabel metal1 0 14454 0 14464 3 Test
rlabel metal1 0 14477 0 14487 3 Clock
rlabel metal1 0 14500 0 14525 3 GND!
rlabel metal1 0 15145 0 15170 3 Vdd!
rlabel metal1 0 15183 0 15193 3 SDI
rlabel metal1 0 13408 0 13418 3 nReset
rlabel metal1 0 13431 0 13441 3 Test
rlabel metal1 0 13454 0 13464 3 Clock
rlabel metal1 0 13477 0 13502 3 GND!
rlabel metal1 0 14122 0 14147 3 Vdd!
rlabel metal1 0 14160 0 14170 3 SDI
rlabel metal1 0 11362 0 11372 3 nReset
rlabel metal1 0 11385 0 11395 3 Test
rlabel metal1 0 11408 0 11418 3 Clock
rlabel metal1 0 11431 0 11456 3 GND!
rlabel metal1 0 12076 0 12101 3 Vdd!
rlabel metal1 0 12114 0 12124 3 SDI
rlabel metal1 0 10339 0 10349 3 nReset
rlabel metal1 0 10362 0 10372 3 Test
rlabel metal1 0 10385 0 10395 3 Clock
rlabel metal1 0 10408 0 10433 3 GND!
rlabel metal1 0 11053 0 11078 3 Vdd!
rlabel metal1 0 11091 0 11101 3 SDI
rlabel metal1 0 9316 0 9326 3 nReset
rlabel metal1 0 9339 0 9349 3 Test
rlabel metal1 0 9362 0 9372 3 Clock
rlabel metal1 0 9385 0 9410 3 GND!
rlabel metal1 0 10030 0 10055 3 Vdd!
rlabel metal1 0 10068 0 10078 3 SDI
rlabel metal1 0 8293 0 8303 3 nReset
rlabel metal1 0 8316 0 8326 3 Test
rlabel metal1 0 8339 0 8349 3 Clock
rlabel metal1 0 8362 0 8387 3 GND!
rlabel metal1 0 9007 0 9032 3 Vdd!
rlabel metal1 0 9045 0 9055 3 SDI
rlabel metal1 0 7270 0 7280 3 nReset
rlabel metal1 0 7293 0 7303 3 Test
rlabel metal1 0 7316 0 7326 3 Clock
rlabel metal1 0 7339 0 7364 3 GND!
rlabel metal1 0 7984 0 8009 3 Vdd!
rlabel metal1 0 8022 0 8032 3 SDI
rlabel metal1 0 6247 0 6257 3 nReset
rlabel metal1 0 6270 0 6280 3 Test
rlabel metal1 0 6293 0 6303 3 Clock
rlabel metal1 0 6316 0 6341 3 GND!
rlabel metal1 0 6961 0 6986 3 Vdd!
rlabel metal1 0 6999 0 7009 3 SDI
rlabel metal1 0 5224 0 5234 3 nReset
rlabel metal1 0 5247 0 5257 3 Test
rlabel metal1 0 5270 0 5280 3 Clock
rlabel metal1 0 5293 0 5318 3 GND!
rlabel metal1 0 5938 0 5963 3 Vdd!
rlabel metal1 0 5976 0 5986 3 SDI
rlabel metal1 0 4201 0 4211 3 nReset
rlabel metal1 0 4224 0 4234 3 Test
rlabel metal1 0 4247 0 4257 3 Clock
rlabel metal1 0 4270 0 4295 3 GND!
rlabel metal1 0 4915 0 4940 3 Vdd!
rlabel metal1 0 4953 0 4963 3 SDI
rlabel metal1 0 3178 0 3188 3 nReset
rlabel metal1 0 3201 0 3211 3 Test
rlabel metal1 0 3224 0 3234 3 Clock
rlabel metal1 0 3247 0 3272 3 GND!
rlabel metal1 0 3892 0 3917 3 Vdd!
rlabel metal1 0 3930 0 3940 3 SDI
rlabel metal1 0 2155 0 2165 3 nReset
rlabel metal1 0 2178 0 2188 3 Test
rlabel metal1 0 2201 0 2211 3 Clock
rlabel metal1 0 2224 0 2249 3 GND!
rlabel metal1 0 2869 0 2894 3 Vdd!
rlabel metal1 0 2907 0 2917 3 SDI
rlabel metal1 0 12385 0 12395 3 nReset
rlabel metal1 0 12408 0 12418 3 Test
rlabel metal1 0 12431 0 12441 3 Clock
rlabel metal1 0 12454 0 12479 3 GND!
rlabel metal1 0 13137 0 13147 3 SDI
rlabel metal1 0 13099 0 13124 3 Vdd!
rlabel metal1 0 1080 0 1090 3 Ir[1]
rlabel metal1 0 1100 0 1110 3 IrIn[1]
rlabel metal1 0 2103 0 2113 3 Ir[2]
rlabel metal1 0 2123 0 2133 3 IrIn[2]
rlabel metal1 0 3126 0 3136 3 Ir[3]
rlabel metal1 0 3146 0 3156 3 IrIn[3]
rlabel metal1 0 4149 0 4159 3 Ir[4]
rlabel metal1 0 4169 0 4179 3 IrIn[4]
rlabel metal1 0 5172 0 5182 3 Ir[5]
rlabel metal1 0 5192 0 5202 3 IrIn[5]
rlabel metal1 0 6195 0 6205 3 Ir[6]
rlabel metal1 0 6215 0 6225 3 IrIn[6]
rlabel metal1 0 7218 0 7228 3 Ir[7]
rlabel metal1 0 7238 0 7248 3 IrIn[7]
rlabel metal1 0 8241 0 8251 3 Ir[8]
rlabel metal1 0 8261 0 8271 3 IrIn[8]
rlabel metal1 0 9264 0 9274 3 Ir[9]
rlabel metal1 0 9284 0 9294 3 IrIn[9]
rlabel metal1 0 10287 0 10297 3 Ir[10]
rlabel metal1 0 10307 0 10317 3 IrIn[10]
rlabel metal1 0 11310 0 11320 3 Ir[11]
rlabel metal1 0 11330 0 11340 3 IrIn[11]
rlabel metal1 0 12333 0 12343 3 Ir[12]
rlabel metal1 0 12353 0 12363 3 IrIn[12]
rlabel metal1 0 13356 0 13366 3 Ir[13]
rlabel metal1 0 13376 0 13386 3 IrIn[13]
rlabel metal1 0 14379 0 14389 3 Ir[14]
rlabel metal1 0 14399 0 14409 3 IrIn[14]
rlabel metal1 0 15402 0 15412 3 Ir[15]
rlabel metal1 0 15422 0 15432 3 IrIn[15]
rlabel metal2 912 16419 924 16419 5 ImmSel
rlabel metal2 120 16419 132 16419 5 IrWe
rlabel metal1 1121 15402 1121 15412 7 Imm[15]
rlabel metal1 1121 14379 1121 14389 7 Imm[14]
rlabel metal1 1121 13356 1121 13366 7 Imm[13]
rlabel metal1 1121 12333 1121 12343 7 Imm[12]
rlabel metal1 1121 11310 1121 11320 7 Imm[11]
rlabel metal1 1121 10287 1121 10297 7 Imm[10]
rlabel metal1 1121 9264 1121 9274 7 Imm[9]
rlabel metal1 1121 8241 1121 8251 7 Imm[8]
rlabel metal1 1121 7218 1121 7228 7 Imm[7]
rlabel metal1 1121 6195 1121 6205 7 Imm[6]
rlabel metal1 1121 5172 1121 5182 7 Imm[5]
rlabel metal1 1121 4149 1121 4159 7 Imm[4]
rlabel metal1 1121 3126 1121 3136 7 Imm[3]
rlabel metal1 1121 2103 1121 2113 7 Imm[2]
rlabel metal1 1121 1080 1121 1090 7 Imm[1]
rlabel metal1 1121 57 1121 67 7 Imm[0]
<< end >>
