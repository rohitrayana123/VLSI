magic
tech c035u
timestamp 1396393625
<< metal1 >>
rect 901 898 2039 908
rect 2053 898 3191 908
rect 3205 898 4343 908
rect 4357 898 5495 908
rect 5509 898 6647 908
rect 6661 898 7799 908
rect 7813 898 8951 908
rect 8965 898 9216 908
rect 37 873 1175 883
rect 1189 873 2327 883
rect 2342 873 3479 883
rect 3493 873 4631 883
rect 4645 873 5783 883
rect 5797 873 6934 883
rect 6949 873 8087 883
rect 9181 876 9216 886
rect 614 850 743 860
rect 757 850 959 860
rect 1764 850 1895 860
rect 1909 850 2111 860
rect 2916 850 3047 860
rect 3061 850 3263 860
rect 4068 849 4199 859
rect 4213 849 4415 859
rect 5221 849 5351 859
rect 5365 849 5567 859
rect 6372 849 6503 859
rect 6517 849 6719 859
rect 7524 849 7655 859
rect 7669 849 7871 859
rect 8677 850 8807 860
rect 8821 850 9023 860
rect 1117 28 2255 38
rect 2269 28 3407 38
rect 3421 28 4559 38
rect 4573 28 5711 38
rect 5725 28 6863 38
rect 6877 28 8014 38
rect 8030 28 9167 38
<< m2contact >>
rect 887 896 901 910
rect 2039 896 2053 910
rect 3191 896 3205 910
rect 4343 896 4357 910
rect 5495 896 5509 910
rect 6647 896 6661 910
rect 7799 896 7813 910
rect 8951 896 8965 910
rect 23 871 37 885
rect 1175 872 1189 886
rect 2327 872 2342 886
rect 3479 872 3493 886
rect 4631 872 4645 886
rect 5783 872 5797 886
rect 6934 871 6949 885
rect 8087 871 8101 885
rect 9167 874 9181 888
rect 599 849 614 863
rect 743 848 757 862
rect 959 847 973 861
rect 1750 848 1764 862
rect 1895 847 1909 861
rect 2111 848 2125 862
rect 2902 848 2916 862
rect 3047 847 3061 861
rect 3263 848 3277 862
rect 4054 847 4068 861
rect 4199 847 4213 861
rect 4415 847 4429 861
rect 5207 847 5221 861
rect 5351 847 5365 861
rect 5567 847 5581 861
rect 6358 847 6372 861
rect 6503 847 6517 861
rect 6719 847 6733 861
rect 7510 847 7524 861
rect 7655 847 7669 861
rect 7871 847 7885 861
rect 8663 848 8677 862
rect 8807 847 8821 861
rect 9023 848 9037 862
rect 1103 26 1117 40
rect 2255 26 2269 40
rect 3407 26 3421 40
rect 4559 26 4573 40
rect 5711 26 5725 40
rect 6863 26 6877 40
rect 8014 26 8030 40
rect 9167 26 9181 40
<< metal2 >>
rect 24 885 36 915
rect 24 844 36 871
rect 72 844 84 915
rect 600 844 612 849
rect 744 844 756 848
rect 816 844 828 915
rect 888 844 900 896
rect 960 844 972 847
rect 1032 844 1044 915
rect 1176 844 1188 872
rect 1224 844 1236 915
rect 1752 844 1764 848
rect 1896 844 1908 847
rect 1968 844 1980 915
rect 2040 844 2052 896
rect 2112 844 2124 848
rect 2184 844 2196 915
rect 2328 844 2340 872
rect 2376 844 2388 915
rect 2904 844 2916 848
rect 3048 844 3060 847
rect 3120 844 3132 915
rect 3192 844 3204 896
rect 3264 844 3276 848
rect 3336 844 3348 915
rect 3480 844 3492 872
rect 3528 844 3540 915
rect 4056 844 4068 847
rect 4200 844 4212 847
rect 4272 844 4284 915
rect 4344 844 4356 896
rect 4416 844 4428 847
rect 4488 844 4500 915
rect 4632 844 4644 872
rect 4680 844 4692 915
rect 5208 844 5220 847
rect 5352 844 5364 847
rect 5424 844 5436 915
rect 5496 844 5508 896
rect 5568 844 5580 847
rect 5640 844 5652 915
rect 5784 844 5796 872
rect 5832 844 5844 915
rect 6360 844 6372 847
rect 6504 844 6516 847
rect 6576 844 6588 915
rect 6648 844 6660 896
rect 6720 844 6732 847
rect 6792 844 6804 915
rect 6936 844 6948 871
rect 6984 844 6996 915
rect 7512 844 7524 847
rect 7656 844 7668 847
rect 7728 844 7740 915
rect 7800 844 7812 896
rect 7872 844 7884 847
rect 7944 844 7956 915
rect 8088 844 8100 871
rect 8136 844 8148 915
rect 8664 844 8676 848
rect 8808 844 8820 847
rect 8880 844 8892 915
rect 8952 844 8964 896
rect 9024 844 9036 848
rect 9096 844 9108 915
rect 9168 844 9180 874
rect 72 21 84 45
rect 816 21 828 45
rect 1032 21 1044 45
rect 1104 40 1116 45
rect 1224 21 1236 45
rect 1968 21 1980 45
rect 2184 21 2196 45
rect 2256 40 2268 45
rect 2376 21 2388 45
rect 3120 21 3132 45
rect 3336 21 3348 45
rect 3408 40 3420 45
rect 3528 21 3540 45
rect 4272 21 4284 45
rect 4488 21 4500 45
rect 4560 40 4572 45
rect 4680 21 4692 45
rect 5424 21 5436 45
rect 5640 21 5652 45
rect 5712 40 5724 45
rect 5832 21 5844 45
rect 6576 21 6588 45
rect 6792 21 6804 45
rect 6864 40 6876 45
rect 6984 21 6996 45
rect 7728 21 7740 45
rect 7944 21 7956 45
rect 8016 40 8028 45
rect 8136 21 8148 45
rect 8880 21 8892 45
rect 9096 21 9108 45
rect 9168 40 9180 45
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 45
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 720 0 1 45
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 936 0 1 45
box 0 0 216 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 1152 0 1 45
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1872 0 1 45
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2088 0 1 45
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 2304 0 1 45
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3024 0 1 45
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3240 0 1 45
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 3456 0 1 45
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4176 0 1 45
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 4392 0 1 45
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 4608 0 1 45
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 5328 0 1 45
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 5544 0 1 45
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 5760 0 1 45
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 6480 0 1 45
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 6696 0 1 45
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 6912 0 1 45
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 7632 0 1 45
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 7848 0 1 45
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 8064 0 1 45
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 8784 0 1 45
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9000 0 1 45
box 0 0 216 799
<< labels >>
rlabel metal1 692 852 692 852 1 Reg0
rlabel metal1 1814 854 1814 854 1 Reg1
rlabel metal1 3107 855 3107 855 1 Reg2
rlabel metal1 4349 852 4349 852 1 Reg3
rlabel metal1 5402 853 5402 853 1 Reg4
rlabel metal1 6613 852 6613 852 1 Reg5
rlabel metal1 7783 854 7783 854 1 Reg6
rlabel metal1 8970 856 8970 856 1 Reg7Out
rlabel metal1 9216 876 9216 886 7 Rd2
rlabel metal1 9216 898 9216 908 7 Rd1
rlabel metal2 5424 915 5436 915 5 Rs1[4]
rlabel metal2 4680 915 4692 915 5 Rw[4]
rlabel metal2 4488 915 4500 915 5 Rs2[3]
rlabel metal2 4272 915 4284 915 5 Rs1[3]
rlabel metal2 3528 915 3540 915 5 Rw[3]
rlabel metal2 3336 915 3348 915 5 Rs2[2]
rlabel metal2 3120 915 3132 915 5 Rs1[2]
rlabel metal2 2376 915 2388 915 5 Rw[2]
rlabel metal2 2184 915 2196 915 5 Rs2[1]
rlabel metal2 1968 915 1980 915 5 Rs1[1]
rlabel metal2 1224 915 1236 915 5 Rw[1]
rlabel metal2 1032 915 1044 915 5 Rs2[0]
rlabel metal2 816 915 828 915 5 Rs1[0]
rlabel metal2 5640 915 5652 915 5 Rs2[4]
rlabel metal2 5832 915 5844 915 5 Rw[5]
rlabel metal2 6576 915 6588 915 5 Rs1[5]
rlabel metal2 6792 915 6804 915 5 Rs2[5]
rlabel metal2 6984 915 6996 915 5 Rw[6]
rlabel metal2 7728 915 7740 915 5 Rs1[6]
rlabel metal2 7944 915 7956 915 5 Rs2[6]
rlabel metal2 8880 915 8892 915 5 Rs1[7]
rlabel metal2 9096 915 9108 915 5 Rs2[7]
rlabel metal2 8136 915 8148 915 5 Rw[7]
rlabel metal2 72 915 84 915 5 Rw[0]
rlabel metal2 24 915 36 915 5 WData
rlabel metal2 816 21 828 21 1 Rs1[0]
rlabel metal2 2184 21 2196 21 1 Rs2[1]
rlabel metal2 5832 21 5844 21 5 Rw[5]
rlabel metal2 6576 21 6588 21 5 Rs1[5]
rlabel metal2 6792 21 6804 21 5 Rs2[5]
rlabel metal2 6984 21 6996 21 5 Rw[6]
rlabel metal2 7944 21 7956 21 5 Rs2[6]
rlabel metal2 8136 21 8148 21 5 Rw[7]
rlabel metal2 8880 21 8892 21 5 Rs1[7]
rlabel metal2 9096 21 9108 21 5 Rs2[7]
rlabel metal2 7728 21 7740 21 5 Rs1[6]
rlabel metal2 5640 21 5652 21 1 Rs2[4]
rlabel metal2 2376 21 2388 21 1 Rw[2]
rlabel metal2 5424 21 5436 21 5 Rs1[4]
rlabel metal2 4488 21 4500 21 5 Rs2[3]
rlabel metal2 4680 21 4692 21 5 Rw[4]
rlabel metal2 4272 21 4284 21 5 Rs1[3]
rlabel metal2 3336 21 3348 21 5 Rs2[2]
rlabel metal2 3528 21 3540 21 5 Rw[3]
rlabel metal2 3120 21 3132 21 5 Rs1[2]
rlabel metal2 1968 21 1980 21 5 Rs1[1]
rlabel metal2 1224 21 1236 21 5 Rw[1]
rlabel metal2 1032 21 1044 21 5 Rs2[0]
rlabel metal2 72 21 84 21 1 Rw[0]
<< end >>
