magic
tech c035u
timestamp 1393517329
<< metal1 >>
rect 614 1144 743 1154
rect 757 1144 2287 1154
rect 2301 1144 3439 1154
rect 3454 1144 4591 1154
rect 4605 1144 5743 1154
rect 5757 1144 6895 1154
rect 6909 1144 8046 1154
rect 8061 1144 9199 1154
rect 1332 1094 1855 1104
rect 1869 1094 2071 1104
rect 2876 1094 3007 1104
rect 3021 1094 3223 1104
rect 4028 1094 4159 1104
rect 4173 1094 4375 1104
rect 5180 1094 5311 1104
rect 5325 1094 5527 1104
rect 6332 1094 6463 1104
rect 6477 1094 6679 1104
rect 7484 1094 7615 1104
rect 7629 1094 7831 1104
rect 8636 1094 8767 1104
rect 8781 1094 8983 1104
rect 9788 1094 9919 1104
rect 9933 1094 10135 1104
rect 0 75 23 85
rect 37 75 10309 85
rect 0 40 1998 50
rect 2013 40 3150 50
rect 3165 40 4302 50
rect 4317 40 5455 50
rect 5470 40 6605 50
rect 6623 40 7757 50
rect 7775 40 8909 50
rect 8927 40 10063 50
rect 10077 40 10309 50
rect 0 5 2215 15
rect 2229 5 3367 15
rect 3381 5 4519 15
rect 4533 5 5671 15
rect 5686 5 6822 15
rect 6840 5 7974 15
rect 7992 5 9126 15
rect 9144 5 10279 15
rect 10293 5 10309 15
<< m2contact >>
rect 598 1139 614 1155
rect 743 1141 757 1155
rect 2287 1143 2301 1157
rect 3439 1143 3454 1157
rect 4591 1143 4605 1157
rect 5743 1143 5757 1157
rect 6895 1143 6909 1157
rect 8046 1142 8061 1156
rect 9199 1143 9214 1158
rect 1318 1092 1332 1106
rect 1855 1091 1869 1105
rect 2071 1091 2085 1105
rect 2862 1092 2876 1106
rect 3007 1091 3021 1105
rect 3223 1092 3237 1106
rect 4014 1092 4028 1106
rect 4159 1091 4173 1105
rect 4375 1092 4389 1106
rect 5166 1092 5180 1106
rect 5311 1091 5325 1105
rect 5527 1092 5541 1106
rect 6318 1092 6332 1106
rect 6463 1091 6477 1105
rect 6679 1092 6693 1106
rect 7470 1092 7484 1106
rect 7615 1091 7629 1105
rect 7831 1092 7845 1106
rect 8622 1092 8636 1106
rect 8767 1091 8781 1105
rect 8983 1092 8997 1106
rect 9774 1092 9788 1106
rect 9919 1091 9933 1105
rect 10135 1092 10149 1106
rect 23 74 37 88
rect 1998 38 2013 52
rect 3150 38 3165 52
rect 4302 38 4317 52
rect 5455 38 5470 53
rect 6605 38 6623 53
rect 7757 38 7775 53
rect 8909 38 8927 53
rect 10063 37 10077 52
rect 2215 4 2229 18
rect 3367 4 3381 18
rect 4519 4 4533 18
rect 5671 3 5686 18
rect 6822 0 6840 15
rect 7974 0 7992 15
rect 9126 0 9144 15
rect 10279 3 10293 18
<< metal2 >>
rect 24 1068 36 1194
rect 72 1068 84 1194
rect 600 1068 612 1139
rect 744 1068 756 1141
rect 792 1068 804 1194
rect 1320 1068 1332 1092
rect 1856 1068 1868 1091
rect 1928 1068 1940 1194
rect 2000 1068 2012 1194
rect 2072 1068 2084 1091
rect 2144 1068 2156 1194
rect 2216 1068 2228 1194
rect 2288 1068 2300 1143
rect 2336 1068 2348 1194
rect 2864 1068 2876 1092
rect 3008 1068 3020 1091
rect 3080 1068 3092 1194
rect 3152 1068 3164 1194
rect 3224 1068 3236 1092
rect 3296 1068 3308 1194
rect 3368 1068 3380 1194
rect 3440 1068 3452 1143
rect 3488 1068 3500 1194
rect 4016 1068 4028 1092
rect 4160 1068 4172 1091
rect 4232 1068 4244 1194
rect 4304 1068 4316 1194
rect 4376 1068 4388 1092
rect 4448 1068 4460 1194
rect 4520 1068 4532 1194
rect 4592 1068 4604 1143
rect 4640 1068 4652 1194
rect 5168 1068 5180 1092
rect 5312 1068 5324 1091
rect 5384 1068 5396 1194
rect 5456 1068 5468 1194
rect 5528 1068 5540 1092
rect 5600 1068 5612 1194
rect 5672 1068 5684 1194
rect 5744 1068 5756 1143
rect 5792 1068 5804 1194
rect 6320 1068 6332 1092
rect 6464 1068 6476 1091
rect 6536 1068 6548 1194
rect 6608 1068 6620 1194
rect 6680 1068 6692 1092
rect 6752 1068 6764 1194
rect 6824 1068 6836 1194
rect 6896 1068 6908 1143
rect 6944 1068 6956 1194
rect 7472 1068 7484 1092
rect 7616 1068 7628 1091
rect 7688 1068 7700 1194
rect 7760 1068 7772 1194
rect 7832 1068 7844 1092
rect 7904 1068 7916 1194
rect 7976 1068 7988 1194
rect 8048 1068 8060 1142
rect 8096 1068 8108 1194
rect 8624 1068 8636 1092
rect 8768 1068 8780 1091
rect 8840 1068 8852 1194
rect 8912 1068 8924 1194
rect 8984 1068 8996 1092
rect 9056 1068 9068 1194
rect 9128 1068 9140 1194
rect 9200 1068 9212 1143
rect 9248 1068 9260 1194
rect 9776 1068 9788 1092
rect 9920 1068 9932 1091
rect 9992 1068 10004 1194
rect 10064 1068 10076 1194
rect 10136 1068 10148 1092
rect 10208 1068 10220 1194
rect 10280 1068 10292 1194
rect 24 88 36 269
rect 2000 52 2012 269
rect 2216 18 2228 269
rect 3152 52 3164 269
rect 3368 18 3380 269
rect 4304 52 4316 269
rect 4520 18 4532 269
rect 5456 53 5468 269
rect 5672 18 5684 269
rect 6608 53 6620 269
rect 6824 15 6836 269
rect 7760 53 7772 269
rect 7976 15 7988 269
rect 8912 53 8924 269
rect 9128 15 9140 269
rect 10064 52 10076 269
rect 10280 18 10292 269
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 269
box 0 0 720 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 720 0 1 269
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 1832 0 1 269
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 2048 0 1 269
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 2264 0 1 269
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 2984 0 1 269
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 3200 0 1 269
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 3416 0 1 269
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 4136 0 1 269
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 4352 0 1 269
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 4568 0 1 269
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 5288 0 1 269
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 5504 0 1 269
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 5720 0 1 269
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 6440 0 1 269
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 6656 0 1 269
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 6872 0 1 269
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 7592 0 1 269
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 7808 0 1 269
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 8024 0 1 269
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 8744 0 1 269
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 8960 0 1 269
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 9176 0 1 269
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 9896 0 1 269
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 10112 0 1 269
box 0 0 216 799
<< labels >>
rlabel metal2 72 1194 84 1194 5 IRWc
rlabel metal2 792 1194 804 1194 5 WData[0]
rlabel metal2 9248 1194 9260 1194 5 WData[7]
rlabel metal2 8096 1194 8108 1194 5 WData[6]
rlabel metal2 6944 1194 6956 1194 5 WData[5]
rlabel metal2 5792 1194 5804 1194 5 WData[4]
rlabel metal2 4640 1194 4652 1194 5 WData[3]
rlabel metal2 3488 1194 3500 1194 5 WData[2]
rlabel metal2 2336 1194 2348 1194 5 WData[1]
<< end >>
