magic
tech c035u
timestamp 1394146861
<< error_s >>
rect 4103 2045 4117 2050
use ALUDecoder ALUDecoder_0
timestamp 1394146776
transform 1 0 0 0 1 2040
box 0 0 7450 1481
use LLIcell_U LLIcell_U_0
timestamp 1393855556
transform 1 0 6816 0 1 998
box 0 0 192 1042
use ALUSlice ALUSlice_1
timestamp 1394146137
transform 1 0 0 0 1 998
box 0 0 7224 1042
use LLIcell_L LLIcell_L_0
timestamp 1393855517
transform 1 0 6816 0 1 -44
box 0 0 192 1042
use ALUSlice ALUSlice_0
timestamp 1394146137
transform 1 0 0 0 1 -44
box 0 0 7224 1042
<< end >>
