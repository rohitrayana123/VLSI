magic
tech c035u
timestamp 1394295027
<< metal1 >>
rect 37 888 1175 898
rect 1189 888 2327 898
rect 2342 888 3479 898
rect 3493 888 4631 898
rect 4645 888 5783 898
rect 5797 888 6934 898
rect 6949 888 8087 898
rect 614 865 743 875
rect 757 865 959 875
rect 1764 865 1895 875
rect 1909 865 2111 875
rect 2916 865 3047 875
rect 3061 865 3263 875
rect 4068 864 4199 874
rect 4213 864 4415 874
rect 5221 864 5351 874
rect 5365 864 5567 874
rect 6372 864 6503 874
rect 6517 864 6719 874
rect 7524 864 7655 874
rect 7669 864 7871 874
rect 8677 865 8807 875
rect 8821 865 9023 875
rect 901 44 2038 54
rect 2053 44 3190 54
rect 3205 44 4343 54
rect 4358 44 5493 54
rect 5511 44 6645 54
rect 6663 44 7797 54
rect 7815 44 8951 54
rect 1117 21 2255 31
rect 2269 21 3407 31
rect 3421 21 4559 31
rect 4574 21 5710 31
rect 5728 21 6862 31
rect 6880 21 8014 31
rect 8032 21 9167 31
<< m2contact >>
rect 23 886 37 900
rect 1175 887 1189 901
rect 2327 887 2342 901
rect 3479 887 3493 901
rect 4631 887 4645 901
rect 5783 887 5797 901
rect 6934 886 6949 900
rect 8087 887 8102 902
rect 599 864 614 878
rect 743 863 757 877
rect 959 862 973 876
rect 1750 863 1764 877
rect 1895 862 1909 876
rect 2111 863 2125 877
rect 2902 863 2916 877
rect 3047 862 3061 876
rect 3263 863 3277 877
rect 4054 862 4068 876
rect 4199 862 4213 876
rect 4415 862 4429 876
rect 5207 862 5221 876
rect 5351 862 5365 876
rect 5567 862 5581 876
rect 6358 862 6372 876
rect 6503 862 6517 876
rect 6719 862 6733 876
rect 7510 862 7524 876
rect 7655 862 7669 876
rect 7871 862 7885 876
rect 8663 863 8677 877
rect 8807 862 8821 876
rect 9023 863 9037 877
rect 886 42 901 56
rect 2038 42 2053 56
rect 3190 42 3205 56
rect 4343 42 4358 57
rect 5493 42 5511 57
rect 6645 42 6663 57
rect 7797 42 7815 57
rect 8951 41 8965 56
rect 1103 20 1117 34
rect 2255 20 2269 34
rect 3407 20 3421 34
rect 4559 19 4574 34
rect 5710 16 5728 31
rect 6862 16 6880 31
rect 8014 16 8032 31
rect 9167 19 9181 34
<< metal2 >>
rect 24 900 36 939
rect 24 859 36 886
rect 72 859 84 939
rect 600 859 612 864
rect 744 859 756 863
rect 816 859 828 939
rect 960 859 972 862
rect 1032 859 1044 939
rect 1176 859 1188 887
rect 1224 859 1236 939
rect 1752 859 1764 863
rect 1896 859 1908 862
rect 1968 859 1980 939
rect 2112 859 2124 863
rect 2184 859 2196 939
rect 2328 859 2340 887
rect 2376 859 2388 939
rect 2904 859 2916 863
rect 3048 859 3060 862
rect 3120 859 3132 939
rect 3264 859 3276 863
rect 3336 859 3348 939
rect 3480 859 3492 887
rect 3528 859 3540 939
rect 4056 859 4068 862
rect 4200 859 4212 862
rect 4272 859 4284 939
rect 4416 859 4428 862
rect 4488 859 4500 939
rect 4632 859 4644 887
rect 4680 859 4692 939
rect 5208 859 5220 862
rect 5352 859 5364 862
rect 5424 859 5436 939
rect 5568 859 5580 862
rect 5640 859 5652 939
rect 5784 859 5796 887
rect 5832 859 5844 939
rect 6360 859 6372 862
rect 6504 859 6516 862
rect 6576 859 6588 939
rect 6720 859 6732 862
rect 6792 859 6804 939
rect 6936 859 6948 886
rect 6984 859 6996 939
rect 7512 859 7524 862
rect 7656 859 7668 862
rect 7728 859 7740 939
rect 7872 859 7884 862
rect 7944 859 7956 939
rect 8088 859 8100 887
rect 8136 859 8148 939
rect 8664 859 8676 863
rect 8808 859 8820 862
rect 8880 859 8892 939
rect 9024 859 9036 863
rect 9096 859 9108 939
rect 72 0 84 60
rect 816 0 828 60
rect 888 56 900 60
rect 1032 0 1044 60
rect 1104 34 1116 60
rect 1224 0 1236 60
rect 1968 0 1980 60
rect 2040 56 2052 60
rect 2184 0 2196 60
rect 2256 34 2268 60
rect 2376 0 2388 60
rect 3120 0 3132 60
rect 3192 56 3204 60
rect 3336 0 3348 60
rect 3408 34 3420 60
rect 3528 0 3540 60
rect 4272 0 4284 60
rect 4344 57 4356 60
rect 4488 0 4500 60
rect 4560 34 4572 60
rect 4680 0 4692 60
rect 5424 0 5436 60
rect 5496 57 5508 60
rect 5640 0 5652 60
rect 5712 31 5724 60
rect 5832 0 5844 60
rect 6576 0 6588 60
rect 6648 57 6660 60
rect 6792 0 6804 60
rect 6864 31 6876 60
rect 6984 0 6996 60
rect 7728 0 7740 60
rect 7800 57 7812 60
rect 7944 0 7956 60
rect 8016 31 8028 60
rect 8136 0 8148 60
rect 8880 0 8892 60
rect 8952 56 8964 60
rect 8952 0 8964 41
rect 9096 0 9108 60
rect 9168 34 9180 60
rect 9168 0 9180 19
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 0 0 1 60
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 720 0 1 60
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 936 0 1 60
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 1152 0 1 60
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1872 0 1 60
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2088 0 1 60
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 2304 0 1 60
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3024 0 1 60
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3240 0 1 60
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 3456 0 1 60
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4176 0 1 60
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 4392 0 1 60
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 4608 0 1 60
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 5328 0 1 60
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 5544 0 1 60
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 5760 0 1 60
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 6480 0 1 60
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 6696 0 1 60
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 6912 0 1 60
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 7632 0 1 60
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 7848 0 1 60
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 8064 0 1 60
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 8784 0 1 60
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9000 0 1 60
box 0 0 216 799
<< labels >>
rlabel metal2 5424 939 5436 939 5 Rs1[4]
rlabel metal2 4680 939 4692 939 5 Rw[4]
rlabel metal2 4488 939 4500 939 5 Rs2[3]
rlabel metal2 4272 939 4284 939 5 Rs1[3]
rlabel metal2 3528 939 3540 939 5 Rw[3]
rlabel metal2 3336 939 3348 939 5 Rs2[2]
rlabel metal2 3120 939 3132 939 5 Rs1[2]
rlabel metal2 2376 939 2388 939 5 Rw[2]
rlabel metal2 2184 939 2196 939 5 Rs2[1]
rlabel metal2 1968 939 1980 939 5 Rs1[1]
rlabel metal2 1224 939 1236 939 5 Rw[1]
rlabel metal2 1032 939 1044 939 5 Rs2[0]
rlabel metal2 816 939 828 939 5 Rs1[0]
rlabel metal2 5640 939 5652 939 5 Rs2[4]
rlabel metal2 5832 939 5844 939 5 Rw[5]
rlabel metal2 6576 939 6588 939 5 Rs1[5]
rlabel metal2 6792 939 6804 939 5 Rs2[5]
rlabel metal2 6984 939 6996 939 5 Rw[6]
rlabel metal2 7728 939 7740 939 5 Rs1[6]
rlabel metal2 7944 939 7956 939 5 Rs2[6]
rlabel metal2 8880 939 8892 939 5 Rs1[7]
rlabel metal2 9096 939 9108 939 5 Rs2[7]
rlabel metal2 8136 939 8148 939 5 Rw[7]
rlabel metal2 72 939 84 939 5 Rw[0]
rlabel metal2 72 0 84 0 1 Rw[0]
rlabel metal2 1032 0 1044 0 5 Rs2[0]
rlabel metal2 1224 0 1236 0 5 Rw[1]
rlabel metal2 1968 0 1980 0 5 Rs1[1]
rlabel metal2 3120 0 3132 0 5 Rs1[2]
rlabel metal2 3528 0 3540 0 5 Rw[3]
rlabel metal2 3336 0 3348 0 5 Rs2[2]
rlabel metal2 4272 0 4284 0 5 Rs1[3]
rlabel metal2 4680 0 4692 0 5 Rw[4]
rlabel metal2 4488 0 4500 0 5 Rs2[3]
rlabel metal2 5424 0 5436 0 5 Rs1[4]
rlabel metal2 2376 0 2388 0 1 Rw[2]
rlabel metal2 5640 0 5652 0 1 Rs2[4]
rlabel metal2 7728 0 7740 0 5 Rs1[6]
rlabel metal2 9096 0 9108 0 5 Rs2[7]
rlabel metal2 8880 0 8892 0 5 Rs1[7]
rlabel metal2 8136 0 8148 0 5 Rw[7]
rlabel metal2 7944 0 7956 0 5 Rs2[6]
rlabel metal2 6984 0 6996 0 5 Rw[6]
rlabel metal2 6792 0 6804 0 5 Rs2[5]
rlabel metal2 6576 0 6588 0 5 Rs1[5]
rlabel metal2 5832 0 5844 0 5 Rw[5]
rlabel metal2 2184 0 2196 0 1 Rs2[1]
rlabel metal2 816 0 828 0 1 Rs1[0]
rlabel metal2 8952 0 8964 0 1 Rd1
rlabel metal2 9168 0 9180 0 1 Rd2
rlabel metal2 24 939 36 939 5 WData
<< end >>
