magic
tech c035u
timestamp 1394217247
<< metal1 >>
rect 0 1021 23 1031
rect 38 1021 1175 1031
rect 1189 1021 2327 1031
rect 2342 1021 3479 1031
rect 3493 1021 4631 1031
rect 4645 1021 5783 1031
rect 5797 1021 6934 1031
rect 6949 1021 8087 1031
rect 614 984 743 994
rect 757 984 959 994
rect 1764 971 1895 981
rect 1909 971 2111 981
rect 2916 971 3047 981
rect 3061 971 3263 981
rect 4068 971 4199 981
rect 4213 971 4415 981
rect 5220 971 5351 981
rect 5365 971 5567 981
rect 6372 971 6503 981
rect 6517 971 6719 981
rect 7524 971 7655 981
rect 7669 971 7871 981
rect 8676 971 8807 981
rect 8821 971 9023 981
rect 0 60 886 70
rect 901 60 2038 70
rect 2053 60 3190 70
rect 3205 60 4343 70
rect 4358 60 5493 70
rect 5511 60 6645 70
rect 6663 60 7797 70
rect 7815 60 8951 70
rect 8965 60 9216 70
rect 0 25 1103 35
rect 1117 25 2255 35
rect 2269 25 3407 35
rect 3421 25 4559 35
rect 4574 25 5710 35
rect 5728 25 6862 35
rect 6880 25 8014 35
rect 8032 25 9167 35
rect 9181 25 9216 35
<< m2contact >>
rect 23 1018 38 1034
rect 1175 1020 1189 1034
rect 2327 1020 2342 1034
rect 3479 1020 3493 1034
rect 4631 1020 4645 1034
rect 5783 1020 5797 1034
rect 6934 1019 6949 1033
rect 8087 1020 8102 1035
rect 599 983 614 997
rect 743 982 757 996
rect 959 981 973 995
rect 1750 969 1764 983
rect 1895 968 1909 982
rect 2111 969 2125 983
rect 2902 969 2916 983
rect 3047 968 3061 982
rect 3263 969 3277 983
rect 4054 969 4068 983
rect 4199 968 4213 982
rect 4415 969 4429 983
rect 5206 969 5220 983
rect 5351 968 5365 982
rect 5567 969 5581 983
rect 6358 969 6372 983
rect 6503 968 6517 982
rect 6719 969 6733 983
rect 7510 969 7524 983
rect 7655 968 7669 982
rect 7871 969 7885 983
rect 8662 969 8676 983
rect 8807 968 8821 982
rect 9023 969 9037 983
rect 886 58 901 72
rect 2038 58 2053 72
rect 3190 58 3205 72
rect 4343 58 4358 73
rect 5493 58 5511 73
rect 6645 58 6663 73
rect 7797 58 7815 73
rect 8951 57 8965 72
rect 1103 24 1117 38
rect 2255 24 2269 38
rect 3407 24 3421 38
rect 4559 23 4574 38
rect 5710 20 5728 35
rect 6862 20 6880 35
rect 8014 20 8032 35
rect 9167 23 9181 38
<< metal2 >>
rect 24 945 36 1018
rect 72 945 84 1075
rect 600 945 612 983
rect 744 945 756 982
rect 816 945 828 1075
rect 960 945 972 981
rect 1032 945 1044 1075
rect 1176 945 1188 1020
rect 1224 945 1236 1075
rect 1752 945 1764 969
rect 1896 945 1908 968
rect 1968 945 1980 1075
rect 2112 945 2124 969
rect 2184 945 2196 1075
rect 2328 945 2340 1020
rect 2376 945 2388 1075
rect 2904 945 2916 969
rect 3048 945 3060 968
rect 3120 945 3132 1075
rect 3264 945 3276 969
rect 3336 945 3348 1075
rect 3480 945 3492 1020
rect 3528 945 3540 1075
rect 4056 945 4068 969
rect 4200 945 4212 968
rect 4272 945 4284 1075
rect 4416 945 4428 969
rect 4488 945 4500 1075
rect 4632 945 4644 1020
rect 4680 945 4692 1075
rect 5208 945 5220 969
rect 5352 945 5364 968
rect 5424 945 5436 1075
rect 5568 945 5580 969
rect 5640 945 5652 1075
rect 5784 945 5796 1020
rect 5832 945 5844 1075
rect 6360 945 6372 969
rect 6504 945 6516 968
rect 6576 945 6588 1075
rect 6720 945 6732 969
rect 6792 945 6804 1075
rect 6936 945 6948 1019
rect 6984 945 6996 1075
rect 7512 945 7524 969
rect 7656 945 7668 968
rect 7728 945 7740 1075
rect 7872 945 7884 969
rect 7944 945 7956 1075
rect 8088 945 8100 1020
rect 8136 945 8148 1075
rect 8664 945 8676 969
rect 8808 945 8820 968
rect 8880 945 8892 1075
rect 9024 945 9036 969
rect 9096 945 9108 1075
rect 72 0 84 146
rect 816 0 828 146
rect 888 72 900 146
rect 1032 0 1044 146
rect 1104 38 1116 146
rect 1224 0 1236 146
rect 1968 0 1980 146
rect 2040 72 2052 146
rect 2184 0 2196 146
rect 2256 38 2268 146
rect 2376 0 2388 146
rect 3120 0 3132 146
rect 3192 72 3204 146
rect 3336 0 3348 146
rect 3408 38 3420 146
rect 3528 0 3540 146
rect 4272 0 4284 146
rect 4344 73 4356 146
rect 4488 0 4500 146
rect 4560 38 4572 146
rect 4680 0 4692 146
rect 5424 0 5436 146
rect 5496 73 5508 146
rect 5640 0 5652 146
rect 5712 35 5724 146
rect 5832 0 5844 146
rect 6576 0 6588 146
rect 6648 73 6660 146
rect 6792 0 6804 146
rect 6864 35 6876 146
rect 6984 0 6996 146
rect 7728 0 7740 146
rect 7800 73 7812 146
rect 7944 0 7956 146
rect 8016 35 8028 146
rect 8136 0 8148 146
rect 8880 0 8892 146
rect 8952 72 8964 146
rect 9096 0 9108 146
rect 9168 38 9180 146
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 0 0 1 146
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 720 0 1 146
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 936 0 1 146
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 1152 0 1 146
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1872 0 1 146
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2088 0 1 146
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 2304 0 1 146
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3024 0 1 146
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3240 0 1 146
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 3456 0 1 146
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4176 0 1 146
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 4392 0 1 146
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 4608 0 1 146
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 5328 0 1 146
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 5544 0 1 146
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 5760 0 1 146
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 6480 0 1 146
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 6696 0 1 146
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 6912 0 1 146
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 7632 0 1 146
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 7848 0 1 146
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 8064 0 1 146
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 8784 0 1 146
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9000 0 1 146
box 0 0 216 799
<< labels >>
rlabel metal2 5424 1075 5436 1075 5 Rs1[4]
rlabel metal2 4680 1075 4692 1075 5 Rw[4]
rlabel metal2 4488 1075 4500 1075 5 Rs2[3]
rlabel metal2 4272 1075 4284 1075 5 Rs1[3]
rlabel metal2 3528 1075 3540 1075 5 Rw[3]
rlabel metal2 3336 1075 3348 1075 5 Rs2[2]
rlabel metal2 3120 1075 3132 1075 5 Rs1[2]
rlabel metal2 2376 1075 2388 1075 5 Rw[2]
rlabel metal2 2184 1075 2196 1075 5 Rs2[1]
rlabel metal2 1968 1075 1980 1075 5 Rs1[1]
rlabel metal2 1224 1075 1236 1075 5 Rw[1]
rlabel metal2 1032 1075 1044 1075 5 Rs2[0]
rlabel metal2 816 1075 828 1075 5 Rs1[0]
rlabel metal2 72 0 84 0 1 Rw[0]
rlabel metal2 1032 0 1044 0 5 Rs2[0]
rlabel metal2 1224 0 1236 0 5 Rw[1]
rlabel metal2 1968 0 1980 0 5 Rs1[1]
rlabel metal2 3120 0 3132 0 5 Rs1[2]
rlabel metal2 3528 0 3540 0 5 Rw[3]
rlabel metal2 3336 0 3348 0 5 Rs2[2]
rlabel metal2 4272 0 4284 0 5 Rs1[3]
rlabel metal2 4680 0 4692 0 5 Rw[4]
rlabel metal2 4488 0 4500 0 5 Rs2[3]
rlabel metal2 5424 0 5436 0 5 Rs1[4]
rlabel metal2 2376 0 2388 0 1 Rw[2]
rlabel metal2 5640 0 5652 0 1 Rs2[4]
rlabel metal2 7728 0 7740 0 5 Rs1[6]
rlabel metal2 9096 0 9108 0 5 Rs2[7]
rlabel metal2 8880 0 8892 0 5 Rs1[7]
rlabel metal2 8136 0 8148 0 5 Rw[7]
rlabel metal2 7944 0 7956 0 5 Rs2[6]
rlabel metal2 6984 0 6996 0 5 Rw[6]
rlabel metal2 6792 0 6804 0 5 Rs2[5]
rlabel metal2 6576 0 6588 0 5 Rs1[5]
rlabel metal2 5832 0 5844 0 5 Rw[5]
rlabel metal2 5640 1075 5652 1075 5 Rs2[4]
rlabel metal2 5832 1075 5844 1075 5 Rw[5]
rlabel metal2 6576 1075 6588 1075 5 Rs1[5]
rlabel metal2 6792 1075 6804 1075 5 Rs2[5]
rlabel metal2 6984 1075 6996 1075 5 Rw[6]
rlabel metal2 7728 1075 7740 1075 5 Rs1[6]
rlabel metal2 7944 1075 7956 1075 5 Rs2[6]
rlabel metal2 8880 1075 8892 1075 5 Rs1[7]
rlabel metal2 9096 1075 9108 1075 5 Rs2[7]
rlabel metal2 8136 1075 8148 1075 5 Rw[7]
rlabel metal2 2184 0 2196 0 1 Rs2[1]
rlabel metal2 72 1075 84 1075 5 Rw[0]
rlabel metal2 816 0 828 0 1 Rs1[0]
rlabel metal1 0 60 0 70 3 Rd1
rlabel metal1 0 25 0 35 3 Rd2
rlabel metal1 0 1021 0 1031 1 WData
rlabel metal1 9216 25 9216 35 7 Rd2
rlabel metal1 9216 60 9216 70 7 Rd1
<< end >>
