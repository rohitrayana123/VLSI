magic
tech c035u
timestamp 1394620980
<< error_s >>
rect 2026 16111 2058 16113
rect 2242 16111 2274 16113
rect 58 15913 68 15919
rect 58 15903 68 15906
rect 58 15890 68 15896
rect 58 15880 68 15883
rect 77 15842 78 15848
rect 58 15197 68 15200
rect 58 15184 68 15190
rect 58 15174 68 15177
rect 58 15161 68 15167
rect 58 15151 68 15154
rect 58 15138 68 15144
rect 58 14913 68 14919
rect 58 14903 68 14906
rect 58 14890 68 14896
rect 58 14880 68 14883
rect 77 14842 78 14848
rect 58 14197 68 14200
rect 58 14184 68 14190
rect 58 14174 68 14177
rect 58 14161 68 14167
rect 58 14151 68 14154
rect 58 14138 68 14144
rect 58 13913 68 13919
rect 58 13903 68 13906
rect 58 13890 68 13896
rect 58 13880 68 13883
rect 77 13842 78 13848
rect 58 13197 68 13200
rect 58 13184 68 13190
rect 58 13174 68 13177
rect 58 13161 68 13167
rect 58 13151 68 13154
rect 58 13138 68 13144
rect 58 12913 68 12919
rect 58 12903 68 12906
rect 58 12890 68 12896
rect 58 12880 68 12883
rect 77 12842 78 12848
rect 58 12197 68 12200
rect 58 12184 68 12190
rect 58 12174 68 12177
rect 58 12161 68 12167
rect 58 12151 68 12154
rect 58 12138 68 12144
rect 58 11913 68 11919
rect 58 11903 68 11906
rect 58 11890 68 11896
rect 58 11880 68 11883
rect 77 11842 78 11848
rect 58 11197 68 11200
rect 58 11184 68 11190
rect 58 11174 68 11177
rect 58 11161 68 11167
rect 58 11151 68 11154
rect 58 11138 68 11144
rect 58 10913 68 10919
rect 58 10903 68 10906
rect 58 10890 68 10896
rect 58 10880 68 10883
rect 77 10842 78 10848
rect 58 10197 68 10200
rect 58 10184 68 10190
rect 58 10174 68 10177
rect 58 10161 68 10167
rect 58 10151 68 10154
rect 58 10138 68 10144
rect 58 9913 68 9919
rect 58 9903 68 9906
rect 58 9890 68 9896
rect 58 9880 68 9883
rect 77 9842 78 9848
rect 58 9197 68 9200
rect 58 9184 68 9190
rect 58 9174 68 9177
rect 58 9161 68 9167
rect 58 9151 68 9154
rect 58 9138 68 9144
rect 58 8913 68 8919
rect 58 8903 68 8906
rect 58 8890 68 8896
rect 58 8880 68 8883
rect 77 8842 78 8848
rect 58 8197 68 8200
rect 58 8184 68 8190
rect 58 8174 68 8177
rect 58 8161 68 8167
rect 58 8151 68 8154
rect 58 8138 68 8144
rect 58 7913 68 7919
rect 58 7903 68 7906
rect 58 7890 68 7896
rect 58 7880 68 7883
rect 77 7842 78 7848
rect 58 7197 68 7200
rect 58 7184 68 7190
rect 58 7174 68 7177
rect 58 7161 68 7167
rect 58 7151 68 7154
rect 58 7138 68 7144
rect 58 6913 68 6919
rect 58 6903 68 6906
rect 58 6890 68 6896
rect 58 6880 68 6883
rect 77 6842 78 6848
rect 58 6197 68 6200
rect 58 6184 68 6190
rect 58 6174 68 6177
rect 58 6161 68 6167
rect 58 6151 68 6154
rect 58 6138 68 6144
rect 58 5913 68 5919
rect 58 5903 68 5906
rect 58 5890 68 5896
rect 58 5880 68 5883
rect 77 5842 78 5848
rect 58 5197 68 5200
rect 58 5184 68 5190
rect 58 5174 68 5177
rect 58 5161 68 5167
rect 58 5151 68 5154
rect 58 5138 68 5144
rect 58 4913 68 4919
rect 58 4903 68 4906
rect 58 4890 68 4896
rect 58 4880 68 4883
rect 77 4842 78 4848
rect 58 4197 68 4200
rect 58 4184 68 4190
rect 58 4174 68 4177
rect 58 4161 68 4167
rect 58 4151 68 4154
rect 58 4138 68 4144
rect 58 3913 68 3919
rect 58 3903 68 3906
rect 58 3890 68 3896
rect 58 3880 68 3883
rect 77 3842 78 3848
rect 58 3197 68 3200
rect 58 3184 68 3190
rect 58 3174 68 3177
rect 58 3161 68 3167
rect 58 3151 68 3154
rect 58 3138 68 3144
rect 58 2913 68 2919
rect 58 2903 68 2906
rect 58 2890 68 2896
rect 58 2880 68 2883
rect 77 2842 78 2848
rect 58 2197 68 2200
rect 58 2184 68 2190
rect 58 2174 68 2177
rect 58 2161 68 2167
rect 58 2151 68 2154
rect 58 2138 68 2144
rect 58 1913 68 1919
rect 58 1903 68 1906
rect 58 1890 68 1896
rect 58 1880 68 1883
rect 77 1842 78 1848
rect 58 1197 68 1200
rect 58 1184 68 1190
rect 58 1174 68 1177
rect 58 1161 68 1167
rect 58 1151 68 1154
rect 58 1138 68 1144
rect 58 913 68 919
rect 58 903 68 906
rect 58 890 68 896
rect 58 880 68 883
rect 77 842 78 848
rect 58 197 68 200
rect 58 184 68 190
rect 58 174 68 177
rect 58 161 68 167
rect 58 151 68 154
rect 58 138 68 144
<< metal1 >>
rect 0 16010 91 16020
rect 0 15903 68 15913
rect 0 15880 68 15890
rect 0 15842 68 15867
rect 0 15197 68 15222
rect 0 15174 68 15184
rect 0 15151 68 15161
rect 0 15128 68 15138
rect 9249 15045 9313 15055
rect 0 15010 91 15020
rect 9033 15023 9313 15033
rect 0 14903 68 14913
rect 0 14880 68 14890
rect 0 14842 68 14867
rect 0 14197 68 14222
rect 0 14174 68 14184
rect 0 14151 68 14161
rect 0 14128 68 14138
rect 9249 14045 9313 14055
rect 0 14010 91 14020
rect 9033 14023 9313 14033
rect 0 13903 68 13913
rect 0 13880 68 13890
rect 0 13842 68 13867
rect 0 13197 68 13222
rect 0 13174 68 13184
rect 0 13151 68 13161
rect 0 13128 68 13138
rect 9249 13045 9313 13055
rect 0 13010 91 13020
rect 9033 13023 9313 13033
rect 0 12903 68 12913
rect 0 12880 68 12890
rect 0 12842 68 12867
rect 0 12197 68 12222
rect 0 12174 68 12184
rect 0 12151 68 12161
rect 0 12128 68 12138
rect 9249 12045 9313 12055
rect 0 12010 91 12020
rect 9033 12023 9313 12033
rect 0 11903 68 11913
rect 0 11880 68 11890
rect 0 11842 68 11867
rect 0 11197 68 11222
rect 0 11174 68 11184
rect 0 11151 68 11161
rect 0 11128 68 11138
rect 9249 11045 9313 11055
rect 0 11010 91 11020
rect 9033 11023 9313 11033
rect 0 10903 68 10913
rect 0 10880 68 10890
rect 0 10842 68 10867
rect 0 10197 68 10222
rect 0 10174 68 10184
rect 0 10151 68 10161
rect 0 10128 68 10138
rect 9249 10045 9313 10055
rect 0 10010 91 10020
rect 9033 10023 9313 10033
rect 0 9903 68 9913
rect 0 9880 68 9890
rect 0 9842 68 9867
rect 0 9197 68 9222
rect 0 9174 68 9184
rect 0 9151 68 9161
rect 0 9128 68 9138
rect 9249 9045 9313 9055
rect 0 9010 91 9020
rect 9033 9023 9313 9033
rect 0 8903 68 8913
rect 0 8880 68 8890
rect 0 8842 68 8867
rect 0 8197 68 8222
rect 0 8174 68 8184
rect 0 8151 68 8161
rect 0 8128 68 8138
rect 9249 8045 9313 8055
rect 0 8010 91 8020
rect 9033 8023 9313 8033
rect 0 7903 68 7913
rect 0 7880 68 7890
rect 0 7842 68 7867
rect 0 7197 68 7222
rect 0 7174 68 7184
rect 0 7151 68 7161
rect 0 7128 68 7138
rect 9249 7045 9313 7055
rect 0 7010 91 7020
rect 9033 7023 9313 7033
rect 0 6903 68 6913
rect 0 6880 68 6890
rect 0 6842 68 6867
rect 0 6197 68 6222
rect 0 6174 68 6184
rect 0 6151 68 6161
rect 0 6128 68 6138
rect 9249 6045 9313 6055
rect 0 6010 91 6020
rect 9033 6023 9313 6033
rect 0 5903 68 5913
rect 0 5880 68 5890
rect 0 5842 68 5867
rect 0 5197 68 5222
rect 0 5174 68 5184
rect 0 5151 68 5161
rect 0 5128 68 5138
rect 9249 5045 9313 5055
rect 0 5010 91 5020
rect 9033 5023 9313 5033
rect 0 4903 68 4913
rect 0 4880 68 4890
rect 0 4842 68 4867
rect 0 4197 68 4222
rect 0 4174 68 4184
rect 0 4151 68 4161
rect 0 4128 68 4138
rect 9249 4045 9313 4055
rect 0 4010 91 4020
rect 9033 4023 9313 4033
rect 0 3903 68 3913
rect 0 3880 68 3890
rect 0 3842 68 3867
rect 0 3197 68 3222
rect 0 3174 68 3184
rect 0 3151 68 3161
rect 0 3128 68 3138
rect 9249 3045 9313 3055
rect 0 3010 91 3020
rect 9033 3023 9313 3033
rect 0 2903 68 2913
rect 0 2880 68 2890
rect 0 2842 68 2867
rect 0 2197 68 2222
rect 0 2174 68 2184
rect 0 2151 68 2161
rect 0 2128 68 2138
rect 9249 2045 9313 2055
rect 0 2010 91 2020
rect 9033 2023 9313 2033
rect 0 1903 68 1913
rect 0 1880 68 1890
rect 0 1842 68 1867
rect 0 1197 68 1222
rect 0 1174 68 1184
rect 0 1151 68 1161
rect 0 1128 68 1138
rect 9249 1045 9313 1055
rect 0 1010 91 1020
rect 9033 1023 9313 1033
rect 0 903 68 913
rect 0 880 68 890
rect 0 842 68 867
rect 0 197 68 222
rect 0 174 68 184
rect 0 151 68 161
rect 0 128 68 138
rect 9249 45 9313 55
rect 9033 23 9313 33
<< m2contact >>
rect 91 16008 105 16022
rect 9235 15043 9249 15057
rect 91 15008 105 15022
rect 9019 15021 9033 15035
rect 9235 14043 9249 14057
rect 91 14008 105 14022
rect 9019 14021 9033 14035
rect 9235 13043 9249 13057
rect 91 13008 105 13022
rect 9019 13021 9033 13035
rect 9235 12043 9249 12057
rect 91 12008 105 12022
rect 9019 12021 9033 12035
rect 9235 11043 9249 11057
rect 91 11008 105 11022
rect 9019 11021 9033 11035
rect 9235 10043 9249 10057
rect 91 10008 105 10022
rect 9019 10021 9033 10035
rect 9235 9043 9249 9057
rect 91 9008 105 9022
rect 9019 9021 9033 9035
rect 9235 8043 9249 8057
rect 91 8008 105 8022
rect 9019 8021 9033 8035
rect 9235 7043 9249 7057
rect 91 7008 105 7022
rect 9019 7021 9033 7035
rect 9235 6043 9249 6057
rect 91 6008 105 6022
rect 9019 6021 9033 6035
rect 9235 5043 9249 5057
rect 91 5008 105 5022
rect 9019 5021 9033 5035
rect 9235 4043 9249 4057
rect 91 4008 105 4022
rect 9019 4021 9033 4035
rect 9235 3043 9249 3057
rect 91 3008 105 3022
rect 9019 3021 9033 3035
rect 9235 2043 9249 2057
rect 91 2008 105 2022
rect 9019 2021 9033 2035
rect 9235 1043 9249 1057
rect 91 1008 105 1022
rect 9019 1021 9033 1035
rect 9235 43 9249 57
rect 9019 21 9033 35
<< metal2 >>
rect 92 17649 104 17662
rect 116 17649 128 17662
rect 140 17649 152 17662
rect 190 17649 202 17662
rect 356 17649 368 17662
rect 380 17649 392 17662
rect 404 17649 416 17662
rect 500 17649 512 17662
rect 524 17649 536 17662
rect 548 17649 560 17662
rect 92 16000 104 16008
rect 140 16000 152 16031
rect 884 16000 896 16031
rect 1100 16000 1112 16031
rect 1292 16000 1304 16031
rect 2036 16000 2048 16031
rect 2252 16000 2264 16031
rect 2444 16000 2456 16031
rect 3188 16000 3200 16031
rect 3404 16000 3416 16031
rect 3596 16000 3608 16031
rect 4340 16000 4352 16031
rect 4556 16000 4568 16031
rect 4748 16000 4760 16031
rect 5492 16000 5504 16031
rect 5708 16000 5720 16031
rect 5900 16000 5912 16031
rect 6644 16000 6656 16031
rect 6860 16000 6872 16031
rect 7052 16000 7064 16031
rect 7796 16000 7808 16031
rect 8012 16000 8024 16031
rect 8204 16000 8216 16031
rect 8948 16000 8960 16031
rect 9164 16000 9176 16031
rect 92 15000 104 15008
rect 140 15000 152 15061
rect 884 15000 896 15061
rect 1100 15000 1112 15061
rect 1292 15000 1304 15061
rect 2036 15000 2048 15061
rect 2252 15000 2264 15061
rect 2444 15000 2456 15061
rect 3188 15000 3200 15061
rect 3404 15000 3416 15061
rect 3596 15000 3608 15061
rect 4340 15000 4352 15061
rect 4556 15000 4568 15061
rect 4748 15000 4760 15061
rect 5492 15000 5504 15061
rect 5708 15000 5720 15061
rect 5900 15000 5912 15061
rect 6644 15000 6656 15061
rect 6860 15000 6872 15061
rect 7052 15000 7064 15061
rect 7796 15000 7808 15061
rect 8012 15000 8024 15061
rect 8204 15000 8216 15061
rect 8948 15000 8960 15061
rect 9020 15035 9032 15061
rect 9164 15000 9176 15061
rect 9236 15057 9248 15061
rect 92 14000 104 14008
rect 140 14000 152 14061
rect 884 14000 896 14061
rect 1100 14000 1112 14061
rect 1292 14000 1304 14061
rect 2036 14000 2048 14061
rect 2252 14000 2264 14061
rect 2444 14000 2456 14061
rect 3188 14000 3200 14061
rect 3404 14000 3416 14061
rect 3596 14000 3608 14061
rect 4340 14000 4352 14061
rect 4556 14000 4568 14061
rect 4748 14000 4760 14061
rect 5492 14000 5504 14061
rect 5708 14000 5720 14061
rect 5900 14000 5912 14061
rect 6644 14000 6656 14061
rect 6860 14000 6872 14061
rect 7052 14000 7064 14061
rect 7796 14000 7808 14061
rect 8012 14000 8024 14061
rect 8204 14000 8216 14061
rect 8948 14000 8960 14061
rect 9020 14035 9032 14061
rect 9164 14000 9176 14061
rect 9236 14057 9248 14061
rect 92 13000 104 13008
rect 140 13000 152 13061
rect 884 13000 896 13061
rect 1100 13000 1112 13061
rect 1292 13000 1304 13061
rect 2036 13000 2048 13061
rect 2252 13000 2264 13061
rect 2444 13000 2456 13061
rect 3188 13000 3200 13061
rect 3404 13000 3416 13061
rect 3596 13000 3608 13061
rect 4340 13000 4352 13061
rect 4556 13000 4568 13061
rect 4748 13000 4760 13061
rect 5492 13000 5504 13061
rect 5708 13000 5720 13061
rect 5900 13000 5912 13061
rect 6644 13000 6656 13061
rect 6860 13000 6872 13061
rect 7052 13000 7064 13061
rect 7796 13000 7808 13061
rect 8012 13000 8024 13061
rect 8204 13000 8216 13061
rect 8948 13000 8960 13061
rect 9020 13035 9032 13061
rect 9164 13000 9176 13061
rect 9236 13057 9248 13061
rect 92 12000 104 12008
rect 140 12000 152 12061
rect 884 12000 896 12061
rect 1100 12000 1112 12061
rect 1292 12000 1304 12061
rect 2036 12000 2048 12061
rect 2252 12000 2264 12061
rect 2444 12000 2456 12061
rect 3188 12000 3200 12061
rect 3404 12000 3416 12061
rect 3596 12000 3608 12061
rect 4340 12000 4352 12061
rect 4556 12000 4568 12061
rect 4748 12000 4760 12061
rect 5492 12000 5504 12061
rect 5708 12000 5720 12061
rect 5900 12000 5912 12061
rect 6644 12000 6656 12061
rect 6860 12000 6872 12061
rect 7052 12000 7064 12061
rect 7796 12000 7808 12061
rect 8012 12000 8024 12061
rect 8204 12000 8216 12061
rect 8948 12000 8960 12061
rect 9020 12035 9032 12061
rect 9164 12000 9176 12061
rect 9236 12057 9248 12061
rect 92 11000 104 11008
rect 140 11000 152 11061
rect 884 11000 896 11061
rect 1100 11000 1112 11061
rect 1292 11000 1304 11061
rect 2036 11000 2048 11061
rect 2252 11000 2264 11061
rect 2444 11000 2456 11061
rect 3188 11000 3200 11061
rect 3404 11000 3416 11061
rect 3596 11000 3608 11061
rect 4340 11000 4352 11061
rect 4556 11000 4568 11061
rect 4748 11000 4760 11061
rect 5492 11000 5504 11061
rect 5708 11000 5720 11061
rect 5900 11000 5912 11061
rect 6644 11000 6656 11061
rect 6860 11000 6872 11061
rect 7052 11000 7064 11061
rect 7796 11000 7808 11061
rect 8012 11000 8024 11061
rect 8204 11000 8216 11061
rect 8948 11000 8960 11061
rect 9020 11035 9032 11061
rect 9164 11000 9176 11061
rect 9236 11057 9248 11061
rect 92 10000 104 10008
rect 140 10000 152 10061
rect 884 10000 896 10061
rect 1100 10000 1112 10061
rect 1292 10000 1304 10061
rect 2036 10000 2048 10061
rect 2252 10000 2264 10061
rect 2444 10000 2456 10061
rect 3188 10000 3200 10061
rect 3404 10000 3416 10061
rect 3596 10000 3608 10061
rect 4340 10000 4352 10061
rect 4556 10000 4568 10061
rect 4748 10000 4760 10061
rect 5492 10000 5504 10061
rect 5708 10000 5720 10061
rect 5900 10000 5912 10061
rect 6644 10000 6656 10061
rect 6860 10000 6872 10061
rect 7052 10000 7064 10061
rect 7796 10000 7808 10061
rect 8012 10000 8024 10061
rect 8204 10000 8216 10061
rect 8948 10000 8960 10061
rect 9020 10035 9032 10061
rect 9164 10000 9176 10061
rect 9236 10057 9248 10061
rect 92 9000 104 9008
rect 140 9000 152 9061
rect 884 9000 896 9061
rect 1100 9000 1112 9061
rect 1292 9000 1304 9061
rect 2036 9000 2048 9061
rect 2252 9000 2264 9061
rect 2444 9000 2456 9061
rect 3188 9000 3200 9061
rect 3404 9000 3416 9061
rect 3596 9000 3608 9061
rect 4340 9000 4352 9061
rect 4556 9000 4568 9061
rect 4748 9000 4760 9061
rect 5492 9000 5504 9061
rect 5708 9000 5720 9061
rect 5900 9000 5912 9061
rect 6644 9000 6656 9061
rect 6860 9000 6872 9061
rect 7052 9000 7064 9061
rect 7796 9000 7808 9061
rect 8012 9000 8024 9061
rect 8204 9000 8216 9061
rect 8948 9000 8960 9061
rect 9020 9035 9032 9061
rect 9164 9000 9176 9061
rect 9236 9057 9248 9061
rect 92 8000 104 8008
rect 140 8000 152 8061
rect 884 8000 896 8061
rect 1100 8000 1112 8061
rect 1292 8000 1304 8061
rect 2036 8000 2048 8061
rect 2252 8000 2264 8061
rect 2444 8000 2456 8061
rect 3188 8000 3200 8061
rect 3404 8000 3416 8061
rect 3596 8000 3608 8061
rect 4340 8000 4352 8061
rect 4556 8000 4568 8061
rect 4748 8000 4760 8061
rect 5492 8000 5504 8061
rect 5708 8000 5720 8061
rect 5900 8000 5912 8061
rect 6644 8000 6656 8061
rect 6860 8000 6872 8061
rect 7052 8000 7064 8061
rect 7796 8000 7808 8061
rect 8012 8000 8024 8061
rect 8204 8000 8216 8061
rect 8948 8000 8960 8061
rect 9020 8035 9032 8061
rect 9164 8000 9176 8061
rect 9236 8057 9248 8061
rect 92 7000 104 7008
rect 140 7000 152 7061
rect 884 7000 896 7061
rect 1100 7000 1112 7061
rect 1292 7000 1304 7061
rect 2036 7000 2048 7061
rect 2252 7000 2264 7061
rect 2444 7000 2456 7061
rect 3188 7000 3200 7061
rect 3404 7000 3416 7061
rect 3596 7000 3608 7061
rect 4340 7000 4352 7061
rect 4556 7000 4568 7061
rect 4748 7000 4760 7061
rect 5492 7000 5504 7061
rect 5708 7000 5720 7061
rect 5900 7000 5912 7061
rect 6644 7000 6656 7061
rect 6860 7000 6872 7061
rect 7052 7000 7064 7061
rect 7796 7000 7808 7061
rect 8012 7000 8024 7061
rect 8204 7000 8216 7061
rect 8948 7000 8960 7061
rect 9020 7035 9032 7061
rect 9164 7000 9176 7061
rect 9236 7057 9248 7061
rect 92 6000 104 6008
rect 140 6000 152 6061
rect 884 6000 896 6061
rect 1100 6000 1112 6061
rect 1292 6000 1304 6061
rect 2036 6000 2048 6061
rect 2252 6000 2264 6061
rect 2444 6000 2456 6061
rect 3188 6000 3200 6061
rect 3404 6000 3416 6061
rect 3596 6000 3608 6061
rect 4340 6000 4352 6061
rect 4556 6000 4568 6061
rect 4748 6000 4760 6061
rect 5492 6000 5504 6061
rect 5708 6000 5720 6061
rect 5900 6000 5912 6061
rect 6644 6000 6656 6061
rect 6860 6000 6872 6061
rect 7052 6000 7064 6061
rect 7796 6000 7808 6061
rect 8012 6000 8024 6061
rect 8204 6000 8216 6061
rect 8948 6000 8960 6061
rect 9020 6035 9032 6061
rect 9164 6000 9176 6061
rect 9236 6057 9248 6061
rect 92 5000 104 5008
rect 140 5000 152 5061
rect 884 5000 896 5061
rect 1100 5000 1112 5061
rect 1292 5000 1304 5061
rect 2036 5000 2048 5061
rect 2252 5000 2264 5061
rect 2444 5000 2456 5061
rect 3188 5000 3200 5061
rect 3404 5000 3416 5061
rect 3596 5000 3608 5061
rect 4340 5000 4352 5061
rect 4556 5000 4568 5061
rect 4748 5000 4760 5061
rect 5492 5000 5504 5061
rect 5708 5000 5720 5061
rect 5900 5000 5912 5061
rect 6644 5000 6656 5061
rect 6860 5000 6872 5061
rect 7052 5000 7064 5061
rect 7796 5000 7808 5061
rect 8012 5000 8024 5061
rect 8204 5000 8216 5061
rect 8948 5000 8960 5061
rect 9020 5035 9032 5061
rect 9164 5000 9176 5061
rect 9236 5057 9248 5061
rect 92 4000 104 4008
rect 140 4000 152 4061
rect 884 4000 896 4061
rect 1100 4000 1112 4061
rect 1292 4000 1304 4061
rect 2036 4000 2048 4061
rect 2252 4000 2264 4061
rect 2444 4000 2456 4061
rect 3188 4000 3200 4061
rect 3404 4000 3416 4061
rect 3596 4000 3608 4061
rect 4340 4000 4352 4061
rect 4556 4000 4568 4061
rect 4748 4000 4760 4061
rect 5492 4000 5504 4061
rect 5708 4000 5720 4061
rect 5900 4000 5912 4061
rect 6644 4000 6656 4061
rect 6860 4000 6872 4061
rect 7052 4000 7064 4061
rect 7796 4000 7808 4061
rect 8012 4000 8024 4061
rect 8204 4000 8216 4061
rect 8948 4000 8960 4061
rect 9020 4035 9032 4061
rect 9164 4000 9176 4061
rect 9236 4057 9248 4061
rect 92 3000 104 3008
rect 140 3000 152 3061
rect 884 3000 896 3061
rect 1100 3000 1112 3061
rect 1292 3000 1304 3061
rect 2036 3000 2048 3061
rect 2252 3000 2264 3061
rect 2444 3000 2456 3061
rect 3188 3000 3200 3061
rect 3404 3000 3416 3061
rect 3596 3000 3608 3061
rect 4340 3000 4352 3061
rect 4556 3000 4568 3061
rect 4748 3000 4760 3061
rect 5492 3000 5504 3061
rect 5708 3000 5720 3061
rect 5900 3000 5912 3061
rect 6644 3000 6656 3061
rect 6860 3000 6872 3061
rect 7052 3000 7064 3061
rect 7796 3000 7808 3061
rect 8012 3000 8024 3061
rect 8204 3000 8216 3061
rect 8948 3000 8960 3061
rect 9020 3035 9032 3061
rect 9164 3000 9176 3061
rect 9236 3057 9248 3061
rect 92 2000 104 2008
rect 140 2000 152 2061
rect 884 2000 896 2061
rect 1100 2000 1112 2061
rect 1292 2000 1304 2061
rect 2036 2000 2048 2061
rect 2252 2000 2264 2061
rect 2444 2000 2456 2061
rect 3188 2000 3200 2061
rect 3404 2000 3416 2061
rect 3596 2000 3608 2061
rect 4340 2000 4352 2061
rect 4556 2000 4568 2061
rect 4748 2000 4760 2061
rect 5492 2000 5504 2061
rect 5708 2000 5720 2061
rect 5900 2000 5912 2061
rect 6644 2000 6656 2061
rect 6860 2000 6872 2061
rect 7052 2000 7064 2061
rect 7796 2000 7808 2061
rect 8012 2000 8024 2061
rect 8204 2000 8216 2061
rect 8948 2000 8960 2061
rect 9020 2035 9032 2061
rect 9164 2000 9176 2061
rect 9236 2057 9248 2061
rect 92 1000 104 1008
rect 140 1000 152 1061
rect 884 1000 896 1061
rect 1100 1000 1112 1061
rect 1292 1000 1304 1061
rect 2036 1000 2048 1061
rect 2252 1000 2264 1061
rect 2444 1000 2456 1061
rect 3188 1000 3200 1061
rect 3404 1000 3416 1061
rect 3596 1000 3608 1061
rect 4340 1000 4352 1061
rect 4556 1000 4568 1061
rect 4748 1000 4760 1061
rect 5492 1000 5504 1061
rect 5708 1000 5720 1061
rect 5900 1000 5912 1061
rect 6644 1000 6656 1061
rect 6860 1000 6872 1061
rect 7052 1000 7064 1061
rect 7796 1000 7808 1061
rect 8012 1000 8024 1061
rect 8204 1000 8216 1061
rect 8948 1000 8960 1061
rect 9020 1035 9032 1061
rect 9164 1000 9176 1061
rect 9236 1057 9248 1061
rect 140 0 152 61
rect 884 0 896 61
rect 1100 0 1112 61
rect 1292 0 1304 61
rect 2036 0 2048 61
rect 2252 0 2264 61
rect 2444 0 2456 61
rect 3188 0 3200 61
rect 3404 0 3416 61
rect 3596 0 3608 61
rect 4340 0 4352 61
rect 4556 0 4568 61
rect 4748 0 4760 61
rect 5492 0 5504 61
rect 5708 0 5720 61
rect 5900 0 5912 61
rect 6644 0 6656 61
rect 6860 0 6872 61
rect 7052 0 7064 61
rect 7796 0 7808 61
rect 8012 0 8024 61
rect 8204 0 8216 61
rect 8948 0 8960 61
rect 9020 35 9032 61
rect 9164 0 9176 61
rect 9236 57 9248 61
use regBlock_decoder regBlock_decoder_0
timestamp 1394493274
transform 1 0 68 0 1 16031
box 0 0 9216 1618
use regBlock_slice regBlock_slice_0
array 0 0 9313 0 15 1000
timestamp 1394620980
transform 1 0 68 0 1 61
box 0 0 9216 1042
<< labels >>
rlabel metal1 9313 45 9313 55 7 Rd2[0]
rlabel metal1 9313 1045 9313 1055 7 Rd2[1]
rlabel metal1 9313 2045 9313 2055 7 Rd2[2]
rlabel metal1 9313 3045 9313 3055 7 Rd2[3]
rlabel metal1 9313 4045 9313 4055 7 Rd2[4]
rlabel metal1 9313 5045 9313 5055 7 Rd2[5]
rlabel metal1 9313 6045 9313 6055 7 Rd2[6]
rlabel metal1 9313 7045 9313 7055 7 Rd2[7]
rlabel metal1 9313 8045 9313 8055 7 Rd2[8]
rlabel metal1 9313 9045 9313 9055 7 Rd2[9]
rlabel metal1 9313 10045 9313 10055 7 Rd2[10]
rlabel metal1 9313 11045 9313 11055 7 Rd2[11]
rlabel metal1 9313 12045 9313 12055 7 Rd2[12]
rlabel metal1 9313 13045 9313 13055 7 Rd2[13]
rlabel metal1 9313 14045 9313 14055 7 Rd2[14]
rlabel metal1 9313 15045 9313 15055 7 Rd2[15]
rlabel metal1 9313 23 9313 33 7 Rd1[0]
rlabel metal1 9313 1023 9313 1033 7 Rd1[1]
rlabel metal1 9313 2023 9313 2033 7 Rd1[2]
rlabel metal1 9313 3023 9313 3033 7 Rd1[3]
rlabel metal1 9313 4023 9313 4033 7 Rd1[4]
rlabel metal1 9313 5023 9313 5033 7 Rd1[5]
rlabel metal1 9313 6023 9313 6033 7 Rd1[6]
rlabel metal1 9313 7023 9313 7033 7 Rd1[7]
rlabel metal1 9313 8023 9313 8033 7 Rd1[8]
rlabel metal1 9313 9023 9313 9033 7 Rd1[9]
rlabel metal1 9313 10023 9313 10033 7 Rd1[10]
rlabel metal1 9313 11023 9313 11033 7 Rd1[11]
rlabel metal1 9313 12023 9313 12033 7 Rd1[12]
rlabel metal1 9313 13023 9313 13033 7 Rd1[13]
rlabel metal1 9313 14023 9313 14033 7 Rd1[14]
rlabel metal1 9313 15023 9313 15033 7 Rd1[15]
rlabel metal1 0 128 0 138 3 nReset
rlabel metal1 0 1128 0 1138 3 nReset
rlabel metal1 0 2128 0 2138 3 nReset
rlabel metal1 0 3128 0 3138 3 nReset
rlabel metal1 0 4128 0 4138 3 nReset
rlabel metal1 0 5128 0 5138 3 nReset
rlabel metal1 0 6128 0 6138 3 nReset
rlabel metal1 0 7128 0 7138 3 nReset
rlabel metal1 0 8128 0 8138 3 nReset
rlabel metal1 0 9128 0 9138 3 nReset
rlabel metal1 0 10128 0 10138 3 nReset
rlabel metal1 0 11128 0 11138 3 nReset
rlabel metal1 0 12128 0 12138 3 nReset
rlabel metal1 0 13128 0 13138 3 nReset
rlabel metal1 0 14128 0 14138 3 nReset
rlabel metal1 0 15128 0 15138 3 nReset
rlabel metal1 0 151 0 161 3 Test
rlabel metal1 0 1151 0 1161 3 Test
rlabel metal1 0 2151 0 2161 3 Test
rlabel metal1 0 3151 0 3161 3 Test
rlabel metal1 0 4151 0 4161 3 Test
rlabel metal1 0 5151 0 5161 3 Test
rlabel metal1 0 6151 0 6161 3 Test
rlabel metal1 0 7151 0 7161 3 Test
rlabel metal1 0 8151 0 8161 3 Test
rlabel metal1 0 9151 0 9161 3 Test
rlabel metal1 0 10151 0 10161 3 Test
rlabel metal1 0 11151 0 11161 3 Test
rlabel metal1 0 12151 0 12161 3 Test
rlabel metal1 0 13151 0 13161 3 Test
rlabel metal1 0 14151 0 14161 3 Test
rlabel metal1 0 15151 0 15161 3 Test
rlabel metal1 0 174 0 184 3 Clock
rlabel metal1 0 1174 0 1184 3 Clock
rlabel metal1 0 2174 0 2184 3 Clock
rlabel metal1 0 3174 0 3184 3 Clock
rlabel metal1 0 4174 0 4184 3 Clock
rlabel metal1 0 5174 0 5184 3 Clock
rlabel metal1 0 6174 0 6184 3 Clock
rlabel metal1 0 7174 0 7184 3 Clock
rlabel metal1 0 8174 0 8184 3 Clock
rlabel metal1 0 9174 0 9184 3 Clock
rlabel metal1 0 10174 0 10184 3 Clock
rlabel metal1 0 11174 0 11184 3 Clock
rlabel metal1 0 12174 0 12184 3 Clock
rlabel metal1 0 13174 0 13184 3 Clock
rlabel metal1 0 14174 0 14184 3 Clock
rlabel metal1 0 15174 0 15184 3 Clock
rlabel metal1 0 197 0 222 3 GND!
rlabel metal1 0 1197 0 1222 3 GND!
rlabel metal1 0 2197 0 2222 3 GND!
rlabel metal1 0 3197 0 3222 3 GND!
rlabel metal1 0 4197 0 4222 3 GND!
rlabel metal1 0 5197 0 5222 3 GND!
rlabel metal1 0 6197 0 6222 3 GND!
rlabel metal1 0 7197 0 7222 3 GND!
rlabel metal1 0 8197 0 8222 3 GND!
rlabel metal1 0 9197 0 9222 3 GND!
rlabel metal1 0 10197 0 10222 3 GND!
rlabel metal1 0 11197 0 11222 3 GND!
rlabel metal1 0 12197 0 12222 3 GND!
rlabel metal1 0 13197 0 13222 3 GND!
rlabel metal1 0 14197 0 14222 3 GND!
rlabel metal1 0 15197 0 15222 3 GND!
rlabel metal1 0 842 0 867 3 Vdd!
rlabel metal1 0 1842 0 1867 3 Vdd!
rlabel metal1 0 2842 0 2867 3 Vdd!
rlabel metal1 0 3842 0 3867 3 Vdd!
rlabel metal1 0 4842 0 4867 3 Vdd!
rlabel metal1 0 5842 0 5867 3 Vdd!
rlabel metal1 0 6842 0 6867 3 Vdd!
rlabel metal1 0 7842 0 7867 3 Vdd!
rlabel metal1 0 8842 0 8867 3 Vdd!
rlabel metal1 0 9842 0 9867 3 Vdd!
rlabel metal1 0 10842 0 10867 3 Vdd!
rlabel metal1 0 11842 0 11867 3 Vdd!
rlabel metal1 0 12842 0 12867 3 Vdd!
rlabel metal1 0 13842 0 13867 3 Vdd!
rlabel metal1 0 14842 0 14867 3 Vdd!
rlabel metal1 0 15842 0 15867 3 Vdd!
rlabel metal1 0 880 0 890 3 SDI
rlabel metal1 0 1880 0 1890 3 SDI
rlabel metal1 0 2880 0 2890 3 SDI
rlabel metal1 0 3880 0 3890 3 SDI
rlabel metal1 0 4880 0 4890 3 SDI
rlabel metal1 0 5880 0 5890 3 SDI
rlabel metal1 0 6880 0 6890 3 SDI
rlabel metal1 0 7880 0 7890 3 SDI
rlabel metal1 0 8880 0 8890 3 SDI
rlabel metal1 0 9880 0 9890 3 SDI
rlabel metal1 0 10880 0 10890 3 SDI
rlabel metal1 0 11880 0 11890 3 SDI
rlabel metal1 0 12880 0 12890 3 SDI
rlabel metal1 0 13880 0 13890 3 SDI
rlabel metal1 0 14880 0 14890 3 SDI
rlabel metal1 0 15880 0 15890 3 SDI
rlabel metal1 0 903 0 913 3 ScanReturn
rlabel metal1 0 1903 0 1913 3 ScanReturn
rlabel metal1 0 2903 0 2913 3 ScanReturn
rlabel metal1 0 3903 0 3913 3 ScanReturn
rlabel metal1 0 4903 0 4913 3 ScanReturn
rlabel metal1 0 5903 0 5913 3 ScanReturn
rlabel metal1 0 6903 0 6913 3 ScanReturn
rlabel metal1 0 7903 0 7913 3 ScanReturn
rlabel metal1 0 8903 0 8913 3 ScanReturn
rlabel metal1 0 9903 0 9913 3 ScanReturn
rlabel metal1 0 10903 0 10913 3 ScanReturn
rlabel metal1 0 11903 0 11913 3 ScanReturn
rlabel metal1 0 12903 0 12913 3 ScanReturn
rlabel metal1 0 13903 0 13913 3 ScanReturn
rlabel metal1 0 14903 0 14913 3 ScanReturn
rlabel metal1 0 15903 0 15913 3 ScanReturn
rlabel metal1 0 1010 0 1020 3 WData[0]
rlabel metal1 0 2010 0 2020 3 WData[1]
rlabel metal1 0 3010 0 3020 3 WData[2]
rlabel metal1 0 4010 0 4020 3 WData[3]
rlabel metal1 0 5010 0 5020 3 WData[4]
rlabel metal1 0 6010 0 6020 3 WData[5]
rlabel metal1 0 7010 0 7020 3 WData[6]
rlabel metal1 0 8010 0 8020 3 WData[7]
rlabel metal1 0 9010 0 9020 3 WData[8]
rlabel metal1 0 10010 0 10020 3 WData[9]
rlabel metal1 0 11010 0 11020 3 WData[10]
rlabel metal1 0 12010 0 12020 3 WData[11]
rlabel metal1 0 13010 0 13020 3 WData[12]
rlabel metal1 0 14010 0 14020 3 WData[13]
rlabel metal1 0 15010 0 15020 3 WData[14]
rlabel metal1 0 16010 0 16020 3 WData[15]
rlabel metal2 356 17662 368 17662 5 Rs1[0]
rlabel metal2 380 17662 392 17662 5 Rs1[1]
rlabel metal2 404 17662 416 17662 5 Rs1[2]
rlabel metal2 500 17662 512 17662 5 Rs2[0]
rlabel metal2 524 17662 536 17662 5 Rs2[1]
rlabel metal2 548 17662 560 17662 5 Rs2[2]
rlabel metal2 92 17662 104 17662 5 Rw[0]
rlabel metal2 116 17662 128 17662 5 Rw[1]
rlabel metal2 140 17662 152 17662 5 Rw[2]
rlabel metal2 190 17662 202 17662 5 We
<< end >>
