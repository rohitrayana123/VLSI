../behavioural/monitor.sv