magic
tech c035u
timestamp 1396906397
<< nwell >>
rect 26811 1155 27123 1553
<< pwell >>
rect 26811 754 27123 1155
<< pohmic >>
rect 26811 830 27123 840
<< nohmic >>
rect 26811 1490 27123 1500
<< metal1 >>
rect 5416 7966 5858 7976
rect 7456 7966 27170 7976
rect 2392 7942 2450 7952
rect 3952 7942 21926 7952
rect 84 7918 1706 7928
rect 2008 7918 14366 7928
rect 84 7894 1754 7904
rect 2200 7894 3302 7904
rect 3664 7894 11822 7904
rect 13504 7894 16898 7904
rect 2428 7870 9986 7880
rect 10096 7870 14570 7880
rect 16036 7870 16442 7880
rect 16696 7868 16714 7882
rect 17632 7868 17650 7882
rect 18556 7870 18770 7880
rect 19264 7868 19282 7882
rect 24436 7870 26354 7880
rect 4408 7846 27122 7856
rect 4984 7822 9650 7832
rect 10948 7822 14906 7832
rect 15568 7822 22766 7832
rect 23584 7822 26126 7832
rect 27112 7822 27493 7832
rect 5836 7798 10898 7808
rect 11800 7798 17834 7808
rect 18736 7798 20246 7808
rect 21088 7796 21106 7810
rect 22672 7798 25286 7808
rect 27160 7798 27493 7808
rect 7540 7774 7994 7784
rect 8392 7774 11786 7784
rect 13624 7774 24446 7784
rect 24808 7774 27146 7784
rect 27184 7774 27493 7784
rect 9244 7750 19706 7760
rect 19768 7748 19786 7762
rect 25048 7750 27493 7760
rect 14356 7726 23210 7736
rect 27136 7726 27493 7736
rect 14176 6893 14690 6903
rect 14008 6869 15458 6879
rect 17440 6869 20306 6879
rect 24400 6869 24674 6879
rect 25888 6869 25898 6879
rect 12712 6845 24386 6855
rect 24400 6845 25874 6855
rect 12448 6821 14306 6831
rect 14656 6821 17426 6831
rect 12232 6797 12698 6807
rect 13864 6797 17858 6807
rect 12184 6773 27493 6783
rect 11512 6749 14162 6759
rect 14416 6749 15050 6759
rect 10816 6725 17642 6735
rect 10408 6701 14138 6711
rect 14224 6701 14882 6711
rect 17968 6701 17978 6711
rect 19192 6701 26738 6711
rect 9832 6677 10490 6687
rect 10744 6677 11810 6687
rect 11824 6677 12866 6687
rect 12880 6677 13586 6687
rect 13600 6677 23474 6687
rect 9808 6653 15074 6663
rect 15088 6653 23858 6663
rect 9616 6629 10610 6639
rect 10720 6629 10874 6639
rect 11320 6629 17018 6639
rect 17032 6629 22130 6639
rect 22144 6629 23762 6639
rect 9352 6605 13538 6615
rect 13552 6605 18074 6615
rect 18088 6605 22226 6615
rect 22240 6605 25082 6615
rect 9328 6581 13178 6591
rect 13192 6581 21290 6591
rect 21784 6581 22154 6591
rect 9208 6557 10466 6567
rect 10480 6557 19178 6567
rect 19192 6557 21770 6567
rect 21784 6557 24170 6567
rect 24184 6557 26042 6567
rect 9160 6533 26570 6543
rect 9112 6509 9182 6519
rect 9280 6509 17954 6519
rect 9088 6485 14006 6495
rect 14020 6485 17306 6495
rect 9040 6461 16874 6471
rect 8848 6437 10802 6447
rect 10816 6437 25730 6447
rect 8728 6413 14042 6423
rect 14056 6413 17786 6423
rect 8680 6389 12914 6399
rect 13576 6389 18578 6399
rect 18592 6389 26570 6399
rect 26584 6389 26690 6399
rect 8536 6365 21746 6375
rect 8488 6341 13754 6351
rect 13840 6341 18986 6351
rect 19000 6341 26858 6351
rect 8416 6317 11162 6327
rect 11224 6317 21362 6327
rect 8224 6293 17402 6303
rect 8176 6269 21530 6279
rect 21544 6269 25298 6279
rect 25312 6269 26234 6279
rect 8152 6245 8210 6255
rect 8392 6245 12626 6255
rect 12640 6245 20690 6255
rect 8104 6221 20978 6231
rect 7960 6197 15890 6207
rect 20008 6197 21194 6207
rect 7936 6173 25130 6183
rect 7912 6149 10850 6159
rect 10912 6149 10922 6159
rect 11152 6149 19730 6159
rect 19744 6149 20714 6159
rect 7888 6125 23018 6135
rect 7864 6101 12266 6111
rect 12280 6101 15434 6111
rect 19528 6101 19670 6111
rect 19864 6101 20318 6111
rect 7792 6077 10298 6087
rect 10312 6077 11378 6087
rect 11392 6077 14834 6087
rect 14848 6077 19514 6087
rect 19528 6077 20642 6087
rect 20656 6077 20666 6087
rect 20680 6077 23234 6087
rect 7720 6053 23882 6063
rect 7624 6029 22610 6039
rect 7552 6005 11426 6015
rect 11440 6005 12338 6015
rect 12352 6005 15914 6015
rect 17176 6005 22202 6015
rect 7528 5981 12842 5991
rect 12856 5981 15626 5991
rect 15640 5981 21074 5991
rect 7288 5957 8114 5967
rect 8128 5957 11402 5967
rect 11416 5957 11762 5967
rect 11776 5957 14426 5967
rect 14440 5957 23282 5967
rect 23296 5957 23834 5967
rect 7216 5933 26882 5943
rect 7048 5909 12242 5919
rect 12256 5909 13802 5919
rect 13816 5909 16298 5919
rect 16312 5909 17798 5919
rect 17812 5909 20018 5919
rect 20032 5909 24290 5919
rect 24304 5909 25106 5919
rect 6832 5885 8258 5895
rect 8272 5885 8402 5895
rect 8464 5885 14786 5895
rect 17152 5885 18242 5895
rect 19816 5885 20210 5895
rect 20512 5885 21302 5895
rect 6664 5861 20858 5871
rect 20872 5861 22178 5871
rect 6616 5837 10622 5847
rect 10636 5837 17354 5847
rect 17368 5837 18194 5847
rect 18208 5837 24098 5847
rect 24112 5837 25802 5847
rect 6568 5813 7010 5823
rect 7024 5813 7826 5823
rect 7840 5813 13130 5823
rect 13144 5813 20498 5823
rect 21064 5813 21506 5823
rect 6472 5789 7082 5799
rect 7192 5789 12434 5799
rect 13528 5789 14690 5799
rect 14704 5789 19610 5799
rect 19624 5789 24122 5799
rect 6328 5765 8594 5775
rect 8608 5765 9050 5775
rect 9064 5765 10778 5775
rect 10792 5765 11690 5775
rect 11704 5765 13946 5775
rect 13960 5765 16610 5775
rect 16624 5765 18866 5775
rect 18880 5765 19994 5775
rect 20008 5765 23978 5775
rect 6304 5741 6314 5751
rect 6448 5741 16730 5751
rect 17056 5741 26090 5751
rect 6256 5717 11042 5727
rect 11104 5717 22250 5727
rect 6232 5693 7094 5703
rect 7108 5693 22658 5703
rect 6208 5669 12866 5679
rect 12880 5669 21050 5679
rect 21064 5669 23930 5679
rect 23944 5669 26666 5679
rect 6184 5645 26498 5655
rect 5800 5621 14474 5631
rect 14584 5621 14690 5631
rect 15160 5621 18362 5631
rect 19504 5621 19970 5631
rect 5776 5597 6146 5607
rect 6160 5597 10826 5607
rect 10840 5597 17594 5607
rect 19336 5597 19946 5607
rect 20488 5597 21206 5607
rect 5752 5573 11522 5583
rect 11608 5573 14762 5583
rect 15040 5573 17522 5583
rect 19312 5573 19466 5583
rect 19600 5573 21794 5583
rect 5656 5549 11474 5559
rect 11488 5549 15170 5559
rect 15520 5549 26378 5559
rect 5560 5525 11018 5535
rect 11080 5525 11906 5535
rect 12040 5525 21914 5535
rect 5512 5501 13634 5511
rect 13648 5501 17210 5511
rect 17224 5501 19154 5511
rect 19168 5501 24194 5511
rect 24208 5501 25826 5511
rect 5464 5477 11858 5487
rect 11872 5477 14618 5487
rect 14632 5477 24914 5487
rect 24928 5477 25610 5487
rect 5416 5453 7634 5463
rect 7648 5453 10406 5463
rect 10420 5453 11354 5463
rect 11368 5453 15722 5463
rect 15736 5453 22946 5463
rect 5320 5429 6722 5439
rect 6736 5429 21098 5439
rect 21112 5429 21938 5439
rect 5032 5405 17186 5415
rect 17488 5405 17738 5415
rect 19216 5405 24578 5415
rect 5008 5381 24746 5391
rect 4984 5357 4994 5367
rect 5128 5357 5954 5367
rect 6088 5357 12026 5367
rect 12088 5357 15506 5367
rect 15520 5357 18146 5367
rect 18160 5357 20474 5367
rect 4912 5333 5126 5343
rect 5272 5333 6674 5343
rect 6688 5333 17762 5343
rect 18184 5333 24650 5343
rect 4864 5309 21386 5319
rect 21400 5309 23690 5319
rect 4816 5285 24842 5295
rect 4792 5261 10346 5271
rect 10360 5261 12218 5271
rect 12232 5261 16490 5271
rect 16504 5261 19130 5271
rect 19144 5261 21146 5271
rect 21160 5261 22874 5271
rect 4744 5237 22010 5247
rect 4720 5213 26162 5223
rect 4552 5189 6026 5199
rect 6040 5189 11666 5199
rect 11896 5189 12170 5199
rect 12688 5189 12722 5199
rect 12808 5189 12926 5199
rect 13072 5189 19850 5199
rect 4528 5165 24434 5175
rect 4432 5141 23306 5151
rect 4384 5117 8306 5127
rect 8320 5117 10442 5127
rect 10576 5117 19802 5127
rect 20248 5117 20426 5127
rect 4336 5093 14858 5103
rect 14920 5093 14930 5103
rect 15016 5093 23642 5103
rect 4288 5069 26018 5079
rect 4144 5045 6626 5055
rect 6640 5045 20882 5055
rect 4120 5021 12482 5031
rect 12664 5021 15554 5031
rect 15568 5021 23954 5031
rect 4096 4997 7298 5007
rect 7312 4997 19778 5007
rect 19792 4997 26906 5007
rect 3976 4973 10034 4983
rect 10240 4973 15770 4983
rect 16552 4973 18938 4983
rect 18952 4973 19670 4983
rect 19768 4973 20042 4983
rect 20200 4973 21506 4983
rect 3856 4949 9314 4959
rect 9328 4949 9698 4959
rect 9712 4949 10490 4959
rect 10504 4949 21338 4959
rect 3808 4925 3938 4935
rect 4000 4925 23306 4935
rect 3784 4901 14450 4911
rect 14512 4901 18458 4911
rect 19120 4901 19922 4911
rect 19936 4901 22082 4911
rect 3736 4877 5210 4887
rect 5224 4877 20234 4887
rect 3520 4853 6386 4863
rect 6400 4853 14810 4863
rect 14824 4853 20618 4863
rect 21256 4853 21866 4863
rect 3472 4829 7514 4839
rect 7528 4829 19898 4839
rect 19912 4829 20834 4839
rect 21040 4829 21626 4839
rect 3448 4805 5690 4815
rect 5704 4805 7154 4815
rect 7168 4805 12146 4815
rect 12160 4805 12674 4815
rect 12688 4805 14210 4815
rect 14224 4805 17546 4815
rect 17560 4805 20522 4815
rect 20536 4805 25538 4815
rect 25552 4805 26426 4815
rect 26440 4805 26474 4815
rect 3376 4781 13346 4791
rect 13408 4781 22154 4791
rect 22168 4781 25466 4791
rect 3352 4757 6818 4767
rect 6832 4757 10058 4767
rect 10072 4757 23618 4767
rect 23632 4757 25202 4767
rect 3328 4733 4250 4743
rect 4264 4733 23066 4743
rect 23512 4733 23546 4743
rect 25576 4733 25586 4743
rect 3160 4709 5186 4719
rect 5200 4709 7850 4719
rect 7864 4709 9026 4719
rect 9040 4709 9698 4719
rect 9712 4709 13274 4719
rect 13288 4709 25562 4719
rect 3064 4685 4298 4695
rect 4312 4685 4850 4695
rect 4864 4685 6530 4695
rect 6544 4685 6890 4695
rect 6904 4685 7994 4695
rect 8008 4685 8690 4695
rect 8704 4685 13442 4695
rect 13456 4685 23498 4695
rect 3040 4661 22994 4671
rect 2920 4637 9626 4647
rect 9640 4637 13154 4647
rect 13216 4637 21674 4647
rect 21688 4637 23330 4647
rect 2872 4613 21698 4623
rect 2824 4589 11570 4599
rect 11584 4589 13058 4599
rect 13072 4589 23426 4599
rect 2776 4565 17450 4575
rect 17848 4565 24074 4575
rect 2752 4541 4226 4551
rect 4240 4541 7442 4551
rect 7456 4541 10250 4551
rect 10264 4541 10946 4551
rect 10960 4541 20162 4551
rect 20776 4541 21506 4551
rect 24256 4541 24362 4551
rect 2728 4517 4562 4527
rect 4576 4517 6938 4527
rect 6952 4517 7946 4527
rect 7960 4517 8330 4527
rect 8344 4517 11978 4527
rect 11992 4517 13106 4527
rect 13120 4517 20954 4527
rect 20968 4517 21458 4527
rect 21472 4517 21890 4527
rect 24232 4517 26834 4527
rect 2704 4493 4010 4503
rect 4024 4493 5066 4503
rect 5080 4493 6914 4503
rect 6928 4493 8066 4503
rect 8080 4493 9278 4503
rect 9292 4493 11954 4503
rect 11968 4493 13202 4503
rect 13216 4493 17666 4503
rect 17680 4493 20114 4503
rect 20128 4493 20738 4503
rect 20944 4493 22514 4503
rect 24160 4493 24254 4503
rect 26632 4493 26642 4503
rect 2680 4469 6962 4479
rect 6976 4469 8138 4479
rect 8152 4469 12314 4479
rect 12328 4469 12602 4479
rect 12616 4469 20018 4479
rect 20080 4469 26618 4479
rect 2656 4445 6866 4455
rect 6928 4445 7094 4455
rect 7144 4445 8618 4455
rect 8632 4445 17210 4455
rect 17344 4445 22034 4455
rect 23920 4445 24674 4455
rect 2632 4421 9146 4431
rect 9160 4421 13082 4431
rect 13096 4421 24410 4431
rect 24904 4421 26762 4431
rect 2608 4397 12530 4407
rect 12544 4397 15242 4407
rect 15256 4397 21026 4407
rect 21040 4397 23210 4407
rect 23224 4397 26978 4407
rect 2584 4373 22058 4383
rect 22072 4373 25970 4383
rect 2536 4349 16586 4359
rect 16696 4349 20186 4359
rect 20272 4349 21410 4359
rect 23752 4349 26642 4359
rect 2512 4325 24338 4335
rect 24640 4325 25658 4335
rect 2440 4301 4466 4311
rect 4480 4301 7034 4311
rect 7048 4301 9554 4311
rect 9568 4301 18002 4311
rect 18016 4301 19490 4311
rect 19504 4301 20906 4311
rect 20920 4301 25922 4311
rect 2392 4277 4970 4287
rect 4984 4277 6074 4287
rect 6088 4277 6578 4287
rect 6592 4277 6650 4287
rect 6664 4277 7610 4287
rect 7624 4277 9938 4287
rect 9952 4277 11258 4287
rect 11272 4277 12458 4287
rect 12472 4277 12530 4287
rect 12544 4277 12554 4287
rect 12568 4277 15698 4287
rect 15712 4277 22586 4287
rect 23464 4277 25034 4287
rect 2368 4253 9242 4263
rect 9256 4253 15962 4263
rect 15976 4253 16514 4263
rect 16528 4253 21338 4263
rect 21352 4253 23186 4263
rect 23200 4253 25754 4263
rect 25864 4253 27122 4263
rect 2296 4229 12362 4239
rect 12616 4229 12626 4239
rect 12976 4229 22850 4239
rect 22936 4229 24458 4239
rect 24616 4229 26714 4239
rect 2272 4205 8930 4215
rect 8944 4205 9458 4215
rect 9472 4205 10706 4215
rect 10768 4205 21434 4215
rect 22024 4205 22226 4215
rect 22552 4205 24314 4215
rect 24328 4205 24746 4215
rect 25768 4205 25802 4215
rect 2200 4181 2402 4191
rect 2416 4181 8450 4191
rect 8464 4181 10514 4191
rect 10528 4181 10826 4191
rect 10840 4181 11282 4191
rect 11296 4181 12794 4191
rect 12808 4181 15722 4191
rect 15736 4181 24866 4191
rect 2176 4157 14306 4167
rect 14320 4157 24554 4167
rect 2128 4133 7250 4143
rect 7264 4133 7586 4143
rect 7672 4133 10658 4143
rect 10768 4133 13682 4143
rect 13696 4133 17762 4143
rect 18304 4133 25898 4143
rect 2080 4109 4322 4119
rect 4336 4109 4826 4119
rect 4840 4109 6938 4119
rect 6952 4109 7562 4119
rect 7576 4109 11786 4119
rect 11800 4109 24434 4119
rect 2056 4085 8042 4095
rect 8056 4085 14258 4095
rect 14512 4085 23546 4095
rect 23560 4085 25346 4095
rect 1984 4061 5306 4071
rect 5320 4061 9458 4071
rect 9472 4061 20162 4071
rect 20176 4061 23162 4071
rect 23632 4061 23690 4071
rect 24208 4061 24938 4071
rect 1960 4037 6770 4047
rect 6784 4037 16850 4047
rect 17056 4037 23378 4047
rect 24352 4037 24794 4047
rect 1888 4013 7130 4023
rect 7144 4013 13922 4023
rect 13936 4013 14354 4023
rect 14560 4013 20210 4023
rect 21472 4013 21938 4023
rect 22264 4013 23810 4023
rect 24424 4013 25850 4023
rect 25864 4013 26402 4023
rect 1840 3989 3530 3999
rect 3544 3989 4898 3999
rect 4912 3989 5090 3999
rect 5104 3989 8906 3999
rect 8920 3989 20714 3999
rect 20728 3989 21242 3999
rect 23008 3989 23018 3999
rect 23176 3989 23234 3999
rect 1816 3965 6410 3975
rect 6424 3965 8354 3975
rect 8368 3965 14090 3975
rect 14104 3965 16922 3975
rect 16936 3965 25322 3975
rect 1744 3941 9914 3951
rect 10048 3941 10406 3951
rect 10552 3941 13370 3951
rect 13840 3941 19346 3951
rect 19888 3941 23114 3951
rect 1696 3917 9890 3927
rect 10144 3917 21650 3927
rect 1672 3893 16778 3903
rect 17248 3893 19538 3903
rect 19912 3893 20318 3903
rect 21664 3893 22082 3903
rect 1648 3869 4178 3879
rect 4192 3869 5714 3879
rect 5728 3869 7706 3879
rect 7720 3869 7754 3879
rect 7768 3869 8906 3879
rect 8920 3869 10394 3879
rect 10408 3869 11282 3879
rect 11296 3869 25610 3879
rect 1624 3845 24050 3855
rect 84 3821 8186 3831
rect 8200 3821 12002 3831
rect 12016 3821 17282 3831
rect 17296 3821 17690 3831
rect 19288 3821 19634 3831
rect 20104 3821 24530 3831
rect 84 3797 19946 3807
rect 24064 3797 25250 3807
rect 1624 3773 3170 3783
rect 3184 3773 3266 3783
rect 3280 3773 3314 3783
rect 3328 3773 7730 3783
rect 7744 3773 13298 3783
rect 13312 3773 14234 3783
rect 14248 3773 15314 3783
rect 15328 3773 17906 3783
rect 17920 3773 19082 3783
rect 19096 3773 19754 3783
rect 19768 3773 21122 3783
rect 21136 3773 23090 3783
rect 23104 3773 23402 3783
rect 23416 3773 26138 3783
rect 1648 3749 3290 3759
rect 3304 3749 4946 3759
rect 4960 3749 5594 3759
rect 5608 3749 6506 3759
rect 6520 3749 6554 3759
rect 6568 3749 7586 3759
rect 7600 3749 8258 3759
rect 8272 3749 9098 3759
rect 9112 3749 9674 3759
rect 9688 3749 10082 3759
rect 10096 3749 12986 3759
rect 13000 3749 15122 3759
rect 15136 3749 16250 3759
rect 16264 3749 21266 3759
rect 21280 3749 21482 3759
rect 21496 3749 21554 3759
rect 21568 3749 23042 3759
rect 23056 3749 23378 3759
rect 23392 3749 23594 3759
rect 1672 3725 2306 3735
rect 2320 3725 12458 3735
rect 13120 3725 13322 3735
rect 13864 3725 17618 3735
rect 17680 3725 17798 3735
rect 19336 3725 20042 3735
rect 21136 3725 21674 3735
rect 1720 3701 4538 3711
rect 4624 3701 5378 3711
rect 5392 3701 14402 3711
rect 14608 3701 17714 3711
rect 1768 3677 17906 3687
rect 1936 3653 14450 3663
rect 14728 3653 15098 3663
rect 15160 3653 21962 3663
rect 2224 3629 14858 3639
rect 15544 3629 27146 3639
rect 2224 3605 4202 3615
rect 4216 3605 5618 3615
rect 5632 3605 6842 3615
rect 6856 3605 7922 3615
rect 7936 3605 10202 3615
rect 10216 3605 12650 3615
rect 12664 3605 12986 3615
rect 13000 3605 13706 3615
rect 13720 3605 14114 3615
rect 14128 3605 24026 3615
rect 2272 3581 6482 3591
rect 6496 3581 7058 3591
rect 7072 3581 10586 3591
rect 10600 3581 21866 3591
rect 21880 3581 21986 3591
rect 22000 3581 25514 3591
rect 2464 3557 6698 3567
rect 6712 3557 7490 3567
rect 7504 3557 10370 3567
rect 10384 3557 11186 3567
rect 11200 3557 12242 3567
rect 12256 3557 13898 3567
rect 13912 3557 14330 3567
rect 14344 3557 16970 3567
rect 16984 3557 21818 3567
rect 24040 3557 24074 3567
rect 2488 3533 17618 3543
rect 17728 3533 24002 3543
rect 2536 3509 2834 3519
rect 2848 3509 4682 3519
rect 4696 3509 8882 3519
rect 8896 3509 16082 3519
rect 16096 3509 16874 3519
rect 17512 3509 20402 3519
rect 2560 3485 2786 3495
rect 2800 3485 2954 3495
rect 2968 3485 4994 3495
rect 5008 3485 6290 3495
rect 6304 3485 8762 3495
rect 8776 3485 9218 3495
rect 9232 3485 13898 3495
rect 13912 3485 14714 3495
rect 14728 3485 16898 3495
rect 16912 3485 20546 3495
rect 20560 3485 21794 3495
rect 21808 3485 24146 3495
rect 24160 3485 24482 3495
rect 2584 3461 3818 3471
rect 3832 3461 13250 3471
rect 13264 3461 25706 3471
rect 2608 3437 19394 3447
rect 20416 3437 24722 3447
rect 2680 3413 11618 3423
rect 12136 3413 20810 3423
rect 2752 3389 5834 3399
rect 5992 3389 14738 3399
rect 14752 3389 16034 3399
rect 16048 3389 18050 3399
rect 18064 3389 23522 3399
rect 2824 3365 6266 3375
rect 6280 3365 13034 3375
rect 13048 3365 22730 3375
rect 22744 3365 27026 3375
rect 2968 3341 14522 3351
rect 15712 3341 21890 3351
rect 21904 3341 24254 3351
rect 3112 3317 7346 3327
rect 7408 3317 16946 3327
rect 16960 3317 24290 3327
rect 3232 3293 18098 3303
rect 3376 3269 3410 3279
rect 3424 3269 3746 3279
rect 3760 3269 10106 3279
rect 10120 3269 12746 3279
rect 12760 3269 17258 3279
rect 17272 3269 18410 3279
rect 18424 3269 25394 3279
rect 3544 3245 3866 3255
rect 3880 3245 6674 3255
rect 6688 3245 8786 3255
rect 8800 3245 18026 3255
rect 18040 3245 19658 3255
rect 3568 3221 4586 3231
rect 4672 3221 6746 3231
rect 6760 3221 7322 3231
rect 7432 3221 7874 3231
rect 7888 3221 16754 3231
rect 16768 3221 19298 3231
rect 19312 3221 19418 3231
rect 19432 3221 24314 3231
rect 24328 3221 25010 3231
rect 3568 3197 26786 3207
rect 3616 3173 24098 3183
rect 26800 3173 26834 3183
rect 3616 3149 5162 3159
rect 5176 3149 8282 3159
rect 8296 3149 8570 3159
rect 8584 3149 9746 3159
rect 9760 3149 15026 3159
rect 15040 3149 17114 3159
rect 17128 3149 17786 3159
rect 18040 3149 18722 3159
rect 19432 3149 19706 3159
rect 3640 3125 8954 3135
rect 8968 3125 20354 3135
rect 20368 3125 22706 3135
rect 22720 3125 23354 3135
rect 3664 3101 19826 3111
rect 19840 3101 20570 3111
rect 20584 3101 22106 3111
rect 22120 3101 23810 3111
rect 3736 3077 3842 3087
rect 3856 3077 4346 3087
rect 4360 3077 16802 3087
rect 16816 3077 21626 3087
rect 3784 3053 4658 3063
rect 4672 3053 14834 3063
rect 14848 3053 21002 3063
rect 3880 3029 5882 3039
rect 6040 3029 6722 3039
rect 6736 3029 9650 3039
rect 9664 3029 13922 3039
rect 13936 3029 14186 3039
rect 14200 3029 15578 3039
rect 15592 3029 17930 3039
rect 20368 3029 20858 3039
rect 3904 3005 20114 3015
rect 3904 2981 7370 2991
rect 7384 2981 12818 2991
rect 12832 2981 24242 2991
rect 3928 2957 27493 2967
rect 4000 2933 10274 2943
rect 10336 2933 14882 2943
rect 15784 2933 20426 2943
rect 4048 2909 11186 2919
rect 11272 2909 26930 2919
rect 4048 2885 12098 2895
rect 12112 2885 14978 2895
rect 17272 2885 17642 2895
rect 4096 2861 10154 2871
rect 10168 2861 19970 2871
rect 19984 2861 24722 2871
rect 4216 2837 19562 2847
rect 19576 2837 20378 2847
rect 20392 2837 26258 2847
rect 4456 2813 20786 2823
rect 4504 2789 10898 2799
rect 11032 2789 21302 2799
rect 4768 2765 15866 2775
rect 20392 2765 21074 2775
rect 5008 2741 9962 2751
rect 10168 2741 16634 2751
rect 5080 2717 5126 2727
rect 5176 2717 9002 2727
rect 9016 2717 20762 2727
rect 20776 2717 23666 2727
rect 5152 2693 6986 2703
rect 7000 2693 25178 2703
rect 5224 2669 18770 2679
rect 5272 2645 6314 2655
rect 6328 2645 12770 2655
rect 12784 2645 20282 2655
rect 20296 2645 24818 2655
rect 24832 2645 26450 2655
rect 5536 2621 5978 2631
rect 6112 2621 16634 2631
rect 5800 2597 12722 2607
rect 12832 2597 21206 2607
rect 5848 2573 12890 2583
rect 12904 2573 26354 2583
rect 6112 2549 20450 2559
rect 6160 2525 25778 2535
rect 6328 2501 8162 2511
rect 8176 2501 8474 2511
rect 8488 2501 8666 2511
rect 8680 2501 10010 2511
rect 10024 2501 10922 2511
rect 10936 2501 12554 2511
rect 12568 2501 13490 2511
rect 13504 2501 14378 2511
rect 14392 2501 15842 2511
rect 15856 2501 21362 2511
rect 21376 2501 25946 2511
rect 6352 2477 16802 2487
rect 20464 2477 26186 2487
rect 6496 2453 21506 2463
rect 25792 2453 26810 2463
rect 6616 2429 14954 2439
rect 6808 2405 8978 2415
rect 8992 2405 26306 2415
rect 6856 2381 21722 2391
rect 6976 2357 10682 2367
rect 10864 2357 17378 2367
rect 7192 2333 7274 2343
rect 7288 2333 9338 2343
rect 9352 2333 9986 2343
rect 10000 2333 11042 2343
rect 11056 2333 13394 2343
rect 13408 2333 13466 2343
rect 13480 2333 13970 2343
rect 13984 2333 14282 2343
rect 14296 2333 16994 2343
rect 17008 2333 17882 2343
rect 17896 2333 20594 2343
rect 20608 2333 22850 2343
rect 7264 2309 7442 2319
rect 7504 2309 7514 2319
rect 7768 2309 21602 2319
rect 7432 2285 10874 2295
rect 11128 2285 25634 2295
rect 7480 2261 9746 2271
rect 9760 2261 10586 2271
rect 10600 2261 19466 2271
rect 19480 2261 24626 2271
rect 24640 2261 25418 2271
rect 7528 2237 9842 2247
rect 10192 2237 25586 2247
rect 7816 2213 17474 2223
rect 7984 2189 8210 2199
rect 8224 2189 14738 2199
rect 14752 2189 22418 2199
rect 8200 2165 9434 2175
rect 9448 2165 15098 2175
rect 15112 2165 22370 2175
rect 8248 2141 8882 2151
rect 8896 2141 9122 2151
rect 9136 2141 9770 2151
rect 9784 2141 12314 2151
rect 12328 2141 13010 2151
rect 13024 2141 21698 2151
rect 8368 2117 9482 2127
rect 9544 2117 15050 2127
rect 17008 2117 17066 2127
rect 8728 2093 9182 2103
rect 9232 2093 17090 2103
rect 17104 2093 20138 2103
rect 20152 2093 22778 2103
rect 8776 2069 13418 2079
rect 13960 2069 14006 2079
rect 14056 2069 14666 2079
rect 14992 2069 15170 2079
rect 8800 2045 19250 2055
rect 19264 2045 21170 2055
rect 9016 2021 9050 2031
rect 9184 2021 9866 2031
rect 10288 2021 10622 2031
rect 11176 2021 11714 2031
rect 12280 2021 24506 2031
rect 9064 1997 10106 2007
rect 10120 1997 14618 2007
rect 14632 1997 22802 2007
rect 22816 1997 23258 2007
rect 9256 1973 9278 1983
rect 9400 1973 17882 1983
rect 17896 1973 21578 1983
rect 9400 1949 26546 1959
rect 9496 1925 16442 1935
rect 9544 1901 17978 1911
rect 9592 1877 15218 1887
rect 9592 1853 17570 1863
rect 9808 1829 17738 1839
rect 9880 1805 24986 1815
rect 10336 1781 24506 1791
rect 24520 1781 24962 1791
rect 10384 1757 10778 1767
rect 11224 1757 19370 1767
rect 19384 1757 27098 1767
rect 10432 1733 10682 1743
rect 10696 1733 21842 1743
rect 10624 1709 12926 1719
rect 12940 1709 18434 1719
rect 18448 1709 19058 1719
rect 19072 1709 24842 1719
rect 24856 1709 25442 1719
rect 25456 1709 26378 1719
rect 11368 1685 11426 1695
rect 11512 1685 19442 1695
rect 21856 1685 22202 1695
rect 11416 1661 24698 1671
rect 12760 1637 12842 1647
rect 13168 1637 13178 1647
rect 13360 1637 13538 1647
rect 14008 1637 24362 1647
rect 13432 1613 13586 1623
rect 14272 1613 18818 1623
rect 18832 1613 24650 1623
rect 14536 1589 15074 1599
rect 17584 1589 17858 1599
rect 27160 1589 27493 1599
rect 14680 1565 14690 1575
rect 27136 1565 27493 1575
rect 26811 1536 27123 1546
rect 26811 1513 27123 1523
rect 26811 1475 27123 1500
rect 26811 830 27123 855
rect 26811 807 27123 817
rect 26811 784 27123 794
rect 26811 761 27123 771
rect 17176 732 22274 742
rect 13024 708 22922 718
rect 12928 684 14018 694
rect 15400 684 26642 694
rect 12496 660 13754 670
rect 15280 660 17690 670
rect 18016 660 25802 670
rect 11464 636 20546 646
rect 20992 636 23738 646
rect 10984 612 21002 622
rect 21232 612 25898 622
rect 10216 588 26018 598
rect 9640 564 25010 574
rect 9568 540 13586 550
rect 13696 540 13802 550
rect 14896 540 22322 550
rect 9448 516 21482 526
rect 8056 492 17522 502
rect 17824 492 24266 502
rect 8008 468 14906 478
rect 15112 468 22082 478
rect 7384 444 21290 454
rect 7096 420 23690 430
rect 26800 420 27493 430
rect 6760 396 15194 406
rect 15208 396 22490 406
rect 22960 396 24770 406
rect 24976 396 24986 406
rect 26752 396 27493 406
rect 6232 372 13778 382
rect 14368 372 17978 382
rect 18328 372 23978 382
rect 24952 370 24970 384
rect 26584 372 26786 382
rect 6064 348 8570 358
rect 8584 348 9914 358
rect 9976 348 18218 358
rect 18352 348 24986 358
rect 5440 324 14066 334
rect 15496 324 25082 334
rect 5296 300 7682 310
rect 7696 300 7802 310
rect 7816 300 20882 310
rect 20896 300 21530 310
rect 5104 276 15338 286
rect 16240 276 18986 286
rect 19936 276 24674 286
rect 4768 252 8282 262
rect 8656 252 23546 262
rect 4504 228 24866 238
rect 4144 204 6386 214
rect 6448 204 26690 214
rect 3520 180 12770 190
rect 12784 180 15818 190
rect 15832 180 22634 190
rect 22648 180 22826 190
rect 2848 156 4610 166
rect 4720 156 10634 166
rect 10936 156 11066 166
rect 11128 154 11146 168
rect 11320 156 17858 166
rect 18592 156 23090 166
rect 2728 132 3674 142
rect 3760 132 8834 142
rect 9280 132 19250 142
rect 20056 132 23282 142
rect 2704 108 6338 118
rect 6424 108 7634 118
rect 7960 108 12170 118
rect 12400 108 13538 118
rect 16840 108 25202 118
rect 84 84 1730 94
rect 1864 84 4778 94
rect 5056 84 13466 94
rect 13528 84 21602 94
rect 84 60 23042 70
rect 5992 36 27493 46
rect 17440 10 17458 24
rect 20152 12 21962 22
rect 26800 12 27493 22
<< m2contact >>
rect 5402 7964 5416 7978
rect 5858 7964 5872 7978
rect 7442 7964 7456 7978
rect 27170 7964 27184 7978
rect 2378 7940 2392 7954
rect 2450 7940 2464 7954
rect 3938 7940 3952 7954
rect 21926 7940 21940 7954
rect 70 7916 84 7930
rect 1706 7916 1720 7930
rect 1994 7916 2008 7930
rect 14366 7916 14380 7930
rect 70 7892 84 7906
rect 1754 7892 1768 7906
rect 2186 7892 2200 7906
rect 3302 7892 3316 7906
rect 3650 7892 3664 7906
rect 11822 7892 11836 7906
rect 13490 7892 13504 7906
rect 16898 7892 16912 7906
rect 2414 7868 2428 7882
rect 9986 7868 10000 7882
rect 10082 7868 10096 7882
rect 14570 7868 14584 7882
rect 16022 7868 16036 7882
rect 16442 7868 16456 7882
rect 16682 7868 16696 7882
rect 17618 7868 17632 7882
rect 18542 7868 18556 7882
rect 18770 7868 18784 7882
rect 19250 7868 19264 7882
rect 24422 7868 24436 7882
rect 26354 7868 26368 7882
rect 4394 7844 4408 7858
rect 27122 7844 27136 7858
rect 4970 7820 4984 7834
rect 9650 7820 9664 7834
rect 10934 7820 10948 7834
rect 14906 7820 14920 7834
rect 15554 7820 15568 7834
rect 22766 7820 22780 7834
rect 23570 7820 23584 7834
rect 26126 7820 26140 7834
rect 27098 7820 27112 7834
rect 27493 7820 27507 7834
rect 5822 7796 5836 7810
rect 10898 7796 10912 7810
rect 11786 7796 11800 7810
rect 17834 7796 17848 7810
rect 18722 7796 18736 7810
rect 20246 7796 20260 7810
rect 21074 7796 21088 7810
rect 22658 7796 22672 7810
rect 25286 7796 25300 7810
rect 27146 7796 27160 7810
rect 27493 7796 27507 7810
rect 7526 7772 7540 7786
rect 7994 7772 8008 7786
rect 8378 7772 8392 7786
rect 11786 7772 11800 7786
rect 13610 7772 13624 7786
rect 24446 7772 24460 7786
rect 24794 7772 24808 7786
rect 27146 7772 27160 7786
rect 27170 7772 27184 7786
rect 27493 7772 27507 7786
rect 9230 7748 9244 7762
rect 19706 7748 19720 7762
rect 19754 7748 19768 7762
rect 25034 7748 25048 7762
rect 27493 7748 27507 7762
rect 14342 7724 14356 7738
rect 23210 7724 23224 7738
rect 27122 7724 27136 7738
rect 27493 7724 27507 7738
rect 14162 6891 14176 6905
rect 14690 6891 14704 6905
rect 13994 6867 14008 6881
rect 15458 6867 15472 6881
rect 17426 6867 17440 6881
rect 20306 6867 20320 6881
rect 24386 6867 24400 6881
rect 24674 6867 24688 6881
rect 25874 6867 25888 6881
rect 25898 6867 25912 6881
rect 12698 6843 12712 6857
rect 24386 6843 24400 6857
rect 25874 6843 25888 6857
rect 12434 6819 12448 6833
rect 14306 6819 14320 6833
rect 14642 6819 14656 6833
rect 17426 6819 17440 6833
rect 12218 6795 12232 6809
rect 12698 6795 12712 6809
rect 13850 6795 13864 6809
rect 17858 6795 17872 6809
rect 12170 6771 12184 6785
rect 27493 6771 27507 6785
rect 11498 6747 11512 6761
rect 14162 6747 14176 6761
rect 14402 6747 14416 6761
rect 15050 6747 15064 6761
rect 10802 6723 10816 6737
rect 17642 6723 17656 6737
rect 10394 6699 10408 6713
rect 14138 6699 14152 6713
rect 14210 6699 14224 6713
rect 14882 6699 14896 6713
rect 17954 6699 17968 6713
rect 17978 6699 17992 6713
rect 19178 6699 19192 6713
rect 26738 6699 26752 6713
rect 9818 6675 9832 6689
rect 10490 6675 10504 6689
rect 10730 6675 10744 6689
rect 11810 6675 11824 6689
rect 12866 6675 12880 6689
rect 13586 6675 13600 6689
rect 23474 6675 23488 6689
rect 9794 6651 9808 6665
rect 15074 6651 15088 6665
rect 23858 6651 23872 6665
rect 9602 6627 9616 6641
rect 10610 6627 10624 6641
rect 10706 6627 10720 6641
rect 10874 6627 10888 6641
rect 11306 6627 11320 6641
rect 17018 6627 17032 6641
rect 22130 6627 22144 6641
rect 23762 6627 23776 6641
rect 9338 6603 9352 6617
rect 13538 6603 13552 6617
rect 18074 6603 18088 6617
rect 22226 6603 22240 6617
rect 25082 6603 25096 6617
rect 9314 6579 9328 6593
rect 13178 6579 13192 6593
rect 21290 6579 21304 6593
rect 21770 6579 21784 6593
rect 22154 6579 22168 6593
rect 9194 6555 9208 6569
rect 10466 6555 10480 6569
rect 19178 6555 19192 6569
rect 21770 6555 21784 6569
rect 24170 6555 24184 6569
rect 26042 6555 26056 6569
rect 9146 6531 9160 6545
rect 26570 6531 26584 6545
rect 9098 6507 9112 6521
rect 9182 6507 9196 6521
rect 9266 6507 9280 6521
rect 17954 6507 17968 6521
rect 9074 6483 9088 6497
rect 14006 6483 14020 6497
rect 17306 6483 17320 6497
rect 9026 6459 9040 6473
rect 16874 6459 16888 6473
rect 8834 6435 8848 6449
rect 10802 6435 10816 6449
rect 25730 6435 25744 6449
rect 8714 6411 8728 6425
rect 14042 6411 14056 6425
rect 17786 6411 17800 6425
rect 8666 6387 8680 6401
rect 12914 6387 12928 6401
rect 13562 6387 13576 6401
rect 18578 6387 18592 6401
rect 26570 6387 26584 6401
rect 26690 6387 26704 6401
rect 8522 6363 8536 6377
rect 21746 6363 21760 6377
rect 8474 6339 8488 6353
rect 13754 6339 13768 6353
rect 13826 6339 13840 6353
rect 18986 6339 19000 6353
rect 26858 6339 26872 6353
rect 8402 6315 8416 6329
rect 11162 6315 11176 6329
rect 11210 6315 11224 6329
rect 21362 6315 21376 6329
rect 8210 6291 8224 6305
rect 17402 6291 17416 6305
rect 8162 6267 8176 6281
rect 21530 6267 21544 6281
rect 25298 6267 25312 6281
rect 26234 6267 26248 6281
rect 8138 6243 8152 6257
rect 8210 6243 8224 6257
rect 8378 6243 8392 6257
rect 12626 6243 12640 6257
rect 20690 6243 20704 6257
rect 8090 6219 8104 6233
rect 20978 6219 20992 6233
rect 7946 6195 7960 6209
rect 15890 6195 15904 6209
rect 19994 6195 20008 6209
rect 21194 6195 21208 6209
rect 7922 6171 7936 6185
rect 25130 6171 25144 6185
rect 7898 6147 7912 6161
rect 10850 6147 10864 6161
rect 10898 6147 10912 6161
rect 10922 6147 10936 6161
rect 11138 6147 11152 6161
rect 19730 6147 19744 6161
rect 20714 6147 20728 6161
rect 7874 6123 7888 6137
rect 23018 6123 23032 6137
rect 7850 6099 7864 6113
rect 12266 6099 12280 6113
rect 15434 6099 15448 6113
rect 19514 6099 19528 6113
rect 19670 6099 19684 6113
rect 19850 6099 19864 6113
rect 20318 6099 20332 6113
rect 7778 6075 7792 6089
rect 10298 6075 10312 6089
rect 11378 6075 11392 6089
rect 14834 6075 14848 6089
rect 19514 6075 19528 6089
rect 20642 6075 20656 6089
rect 20666 6075 20680 6089
rect 23234 6075 23248 6089
rect 7706 6051 7720 6065
rect 23882 6051 23896 6065
rect 7610 6027 7624 6041
rect 22610 6027 22624 6041
rect 7538 6003 7552 6017
rect 11426 6003 11440 6017
rect 12338 6003 12352 6017
rect 15914 6003 15928 6017
rect 17162 6003 17176 6017
rect 22202 6003 22216 6017
rect 7514 5979 7528 5993
rect 12842 5979 12856 5993
rect 15626 5979 15640 5993
rect 21074 5979 21088 5993
rect 7274 5955 7288 5969
rect 8114 5955 8128 5969
rect 11402 5955 11416 5969
rect 11762 5955 11776 5969
rect 14426 5955 14440 5969
rect 23282 5955 23296 5969
rect 23834 5955 23848 5969
rect 7202 5931 7216 5945
rect 26882 5931 26896 5945
rect 7034 5907 7048 5921
rect 12242 5907 12256 5921
rect 13802 5907 13816 5921
rect 16298 5907 16312 5921
rect 17798 5907 17812 5921
rect 20018 5907 20032 5921
rect 24290 5907 24304 5921
rect 25106 5907 25120 5921
rect 6818 5883 6832 5897
rect 8258 5883 8272 5897
rect 8402 5883 8416 5897
rect 8450 5883 8464 5897
rect 14786 5883 14800 5897
rect 17138 5883 17152 5897
rect 18242 5883 18256 5897
rect 19802 5883 19816 5897
rect 20210 5883 20224 5897
rect 20498 5883 20512 5897
rect 21302 5883 21316 5897
rect 6650 5859 6664 5873
rect 20858 5859 20872 5873
rect 22178 5859 22192 5873
rect 6602 5835 6616 5849
rect 10622 5835 10636 5849
rect 17354 5835 17368 5849
rect 18194 5835 18208 5849
rect 24098 5835 24112 5849
rect 25802 5835 25816 5849
rect 6554 5811 6568 5825
rect 7010 5811 7024 5825
rect 7826 5811 7840 5825
rect 13130 5811 13144 5825
rect 20498 5811 20512 5825
rect 21050 5811 21064 5825
rect 21506 5811 21520 5825
rect 6458 5787 6472 5801
rect 7082 5787 7096 5801
rect 7178 5787 7192 5801
rect 12434 5787 12448 5801
rect 13514 5787 13528 5801
rect 14690 5787 14704 5801
rect 19610 5787 19624 5801
rect 24122 5787 24136 5801
rect 6314 5763 6328 5777
rect 8594 5763 8608 5777
rect 9050 5763 9064 5777
rect 10778 5763 10792 5777
rect 11690 5763 11704 5777
rect 13946 5763 13960 5777
rect 16610 5763 16624 5777
rect 18866 5763 18880 5777
rect 19994 5763 20008 5777
rect 23978 5763 23992 5777
rect 6290 5739 6304 5753
rect 6314 5739 6328 5753
rect 6434 5739 6448 5753
rect 16730 5739 16744 5753
rect 17042 5739 17056 5753
rect 26090 5739 26104 5753
rect 6242 5715 6256 5729
rect 11042 5715 11056 5729
rect 11090 5715 11104 5729
rect 22250 5715 22264 5729
rect 6218 5691 6232 5705
rect 7094 5691 7108 5705
rect 22658 5691 22672 5705
rect 6194 5667 6208 5681
rect 12866 5667 12880 5681
rect 21050 5667 21064 5681
rect 23930 5667 23944 5681
rect 26666 5667 26680 5681
rect 6170 5643 6184 5657
rect 26498 5643 26512 5657
rect 5786 5619 5800 5633
rect 14474 5619 14488 5633
rect 14570 5619 14584 5633
rect 14690 5619 14704 5633
rect 15146 5619 15160 5633
rect 18362 5619 18376 5633
rect 19490 5619 19504 5633
rect 19970 5619 19984 5633
rect 5762 5595 5776 5609
rect 6146 5595 6160 5609
rect 10826 5595 10840 5609
rect 17594 5595 17608 5609
rect 19322 5595 19336 5609
rect 19946 5595 19960 5609
rect 20474 5595 20488 5609
rect 21206 5595 21220 5609
rect 5738 5571 5752 5585
rect 11522 5571 11536 5585
rect 11594 5571 11608 5585
rect 14762 5571 14776 5585
rect 15026 5571 15040 5585
rect 17522 5571 17536 5585
rect 19298 5571 19312 5585
rect 19466 5571 19480 5585
rect 19586 5571 19600 5585
rect 21794 5571 21808 5585
rect 5642 5547 5656 5561
rect 11474 5547 11488 5561
rect 15170 5547 15184 5561
rect 15506 5547 15520 5561
rect 26378 5547 26392 5561
rect 5546 5523 5560 5537
rect 11018 5523 11032 5537
rect 11066 5523 11080 5537
rect 11906 5523 11920 5537
rect 12026 5523 12040 5537
rect 21914 5523 21928 5537
rect 5498 5499 5512 5513
rect 13634 5499 13648 5513
rect 17210 5499 17224 5513
rect 19154 5499 19168 5513
rect 24194 5499 24208 5513
rect 25826 5499 25840 5513
rect 5450 5475 5464 5489
rect 11858 5475 11872 5489
rect 14618 5475 14632 5489
rect 24914 5475 24928 5489
rect 25610 5475 25624 5489
rect 5402 5451 5416 5465
rect 7634 5451 7648 5465
rect 10406 5451 10420 5465
rect 11354 5451 11368 5465
rect 15722 5451 15736 5465
rect 22946 5451 22960 5465
rect 5306 5427 5320 5441
rect 6722 5427 6736 5441
rect 21098 5427 21112 5441
rect 21938 5427 21952 5441
rect 5018 5403 5032 5417
rect 17186 5403 17200 5417
rect 17474 5403 17488 5417
rect 17738 5403 17752 5417
rect 19202 5403 19216 5417
rect 24578 5403 24592 5417
rect 4994 5379 5008 5393
rect 24746 5379 24760 5393
rect 4970 5355 4984 5369
rect 4994 5355 5008 5369
rect 5114 5355 5128 5369
rect 5954 5355 5968 5369
rect 6074 5355 6088 5369
rect 12026 5355 12040 5369
rect 12074 5355 12088 5369
rect 15506 5355 15520 5369
rect 18146 5355 18160 5369
rect 20474 5355 20488 5369
rect 4898 5331 4912 5345
rect 5126 5331 5140 5345
rect 5258 5331 5272 5345
rect 6674 5331 6688 5345
rect 17762 5331 17776 5345
rect 18170 5331 18184 5345
rect 24650 5331 24664 5345
rect 4850 5307 4864 5321
rect 21386 5307 21400 5321
rect 23690 5307 23704 5321
rect 4802 5283 4816 5297
rect 24842 5283 24856 5297
rect 4778 5259 4792 5273
rect 10346 5259 10360 5273
rect 12218 5259 12232 5273
rect 16490 5259 16504 5273
rect 19130 5259 19144 5273
rect 21146 5259 21160 5273
rect 22874 5259 22888 5273
rect 4730 5235 4744 5249
rect 22010 5235 22024 5249
rect 4706 5211 4720 5225
rect 26162 5211 26176 5225
rect 4538 5187 4552 5201
rect 6026 5187 6040 5201
rect 11666 5187 11680 5201
rect 11882 5187 11896 5201
rect 12170 5187 12184 5201
rect 12674 5187 12688 5201
rect 12722 5187 12736 5201
rect 12794 5187 12808 5201
rect 12926 5187 12940 5201
rect 13058 5187 13072 5201
rect 19850 5187 19864 5201
rect 4514 5163 4528 5177
rect 24434 5163 24448 5177
rect 4418 5139 4432 5153
rect 23306 5139 23320 5153
rect 4370 5115 4384 5129
rect 8306 5115 8320 5129
rect 10442 5115 10456 5129
rect 10562 5115 10576 5129
rect 19802 5115 19816 5129
rect 20234 5115 20248 5129
rect 20426 5115 20440 5129
rect 4322 5091 4336 5105
rect 14858 5091 14872 5105
rect 14906 5091 14920 5105
rect 14930 5091 14944 5105
rect 15002 5091 15016 5105
rect 23642 5091 23656 5105
rect 4274 5067 4288 5081
rect 26018 5067 26032 5081
rect 4130 5043 4144 5057
rect 6626 5043 6640 5057
rect 20882 5043 20896 5057
rect 4106 5019 4120 5033
rect 12482 5019 12496 5033
rect 12650 5019 12664 5033
rect 15554 5019 15568 5033
rect 23954 5019 23968 5033
rect 4082 4995 4096 5009
rect 7298 4995 7312 5009
rect 19778 4995 19792 5009
rect 26906 4995 26920 5009
rect 3962 4971 3976 4985
rect 10034 4971 10048 4985
rect 10226 4971 10240 4985
rect 15770 4971 15784 4985
rect 16538 4971 16552 4985
rect 18938 4971 18952 4985
rect 19670 4971 19684 4985
rect 19754 4971 19768 4985
rect 20042 4971 20056 4985
rect 20186 4971 20200 4985
rect 21506 4971 21520 4985
rect 3842 4947 3856 4961
rect 9314 4947 9328 4961
rect 9698 4947 9712 4961
rect 10490 4947 10504 4961
rect 21338 4947 21352 4961
rect 3794 4923 3808 4937
rect 3938 4923 3952 4937
rect 3986 4923 4000 4937
rect 23306 4923 23320 4937
rect 3770 4899 3784 4913
rect 14450 4899 14464 4913
rect 14498 4899 14512 4913
rect 18458 4899 18472 4913
rect 19106 4899 19120 4913
rect 19922 4899 19936 4913
rect 22082 4899 22096 4913
rect 3722 4875 3736 4889
rect 5210 4875 5224 4889
rect 20234 4875 20248 4889
rect 3506 4851 3520 4865
rect 6386 4851 6400 4865
rect 14810 4851 14824 4865
rect 20618 4851 20632 4865
rect 21242 4851 21256 4865
rect 21866 4851 21880 4865
rect 3458 4827 3472 4841
rect 7514 4827 7528 4841
rect 19898 4827 19912 4841
rect 20834 4827 20848 4841
rect 21026 4827 21040 4841
rect 21626 4827 21640 4841
rect 3434 4803 3448 4817
rect 5690 4803 5704 4817
rect 7154 4803 7168 4817
rect 12146 4803 12160 4817
rect 12674 4803 12688 4817
rect 14210 4803 14224 4817
rect 17546 4803 17560 4817
rect 20522 4803 20536 4817
rect 25538 4803 25552 4817
rect 26426 4803 26440 4817
rect 26474 4803 26488 4817
rect 3362 4779 3376 4793
rect 13346 4779 13360 4793
rect 13394 4779 13408 4793
rect 22154 4779 22168 4793
rect 25466 4779 25480 4793
rect 3338 4755 3352 4769
rect 6818 4755 6832 4769
rect 10058 4755 10072 4769
rect 23618 4755 23632 4769
rect 25202 4755 25216 4769
rect 3314 4731 3328 4745
rect 4250 4731 4264 4745
rect 23066 4731 23080 4745
rect 23498 4731 23512 4745
rect 23546 4731 23560 4745
rect 25562 4731 25576 4745
rect 25586 4731 25600 4745
rect 3146 4707 3160 4721
rect 5186 4707 5200 4721
rect 7850 4707 7864 4721
rect 9026 4707 9040 4721
rect 9698 4707 9712 4721
rect 13274 4707 13288 4721
rect 25562 4707 25576 4721
rect 3050 4683 3064 4697
rect 4298 4683 4312 4697
rect 4850 4683 4864 4697
rect 6530 4683 6544 4697
rect 6890 4683 6904 4697
rect 7994 4683 8008 4697
rect 8690 4683 8704 4697
rect 13442 4683 13456 4697
rect 23498 4683 23512 4697
rect 3026 4659 3040 4673
rect 22994 4659 23008 4673
rect 2906 4635 2920 4649
rect 9626 4635 9640 4649
rect 13154 4635 13168 4649
rect 13202 4635 13216 4649
rect 21674 4635 21688 4649
rect 23330 4635 23344 4649
rect 2858 4611 2872 4625
rect 21698 4611 21712 4625
rect 2810 4587 2824 4601
rect 11570 4587 11584 4601
rect 13058 4587 13072 4601
rect 23426 4587 23440 4601
rect 2762 4563 2776 4577
rect 17450 4563 17464 4577
rect 17834 4563 17848 4577
rect 24074 4563 24088 4577
rect 2738 4539 2752 4553
rect 4226 4539 4240 4553
rect 7442 4539 7456 4553
rect 10250 4539 10264 4553
rect 10946 4539 10960 4553
rect 20162 4539 20176 4553
rect 20762 4539 20776 4553
rect 21506 4539 21520 4553
rect 24242 4539 24256 4553
rect 24362 4539 24376 4553
rect 2714 4515 2728 4529
rect 4562 4515 4576 4529
rect 6938 4515 6952 4529
rect 7946 4515 7960 4529
rect 8330 4515 8344 4529
rect 11978 4515 11992 4529
rect 13106 4515 13120 4529
rect 20954 4515 20968 4529
rect 21458 4515 21472 4529
rect 21890 4515 21904 4529
rect 24218 4515 24232 4529
rect 26834 4515 26848 4529
rect 2690 4491 2704 4505
rect 4010 4491 4024 4505
rect 5066 4491 5080 4505
rect 6914 4491 6928 4505
rect 8066 4491 8080 4505
rect 9278 4491 9292 4505
rect 11954 4491 11968 4505
rect 13202 4491 13216 4505
rect 17666 4491 17680 4505
rect 20114 4491 20128 4505
rect 20738 4491 20752 4505
rect 20930 4491 20944 4505
rect 22514 4491 22528 4505
rect 24146 4491 24160 4505
rect 24254 4491 24268 4505
rect 26618 4491 26632 4505
rect 26642 4491 26656 4505
rect 2666 4467 2680 4481
rect 6962 4467 6976 4481
rect 8138 4467 8152 4481
rect 12314 4467 12328 4481
rect 12602 4467 12616 4481
rect 20018 4467 20032 4481
rect 20066 4467 20080 4481
rect 26618 4467 26632 4481
rect 2642 4443 2656 4457
rect 6866 4443 6880 4457
rect 6914 4443 6928 4457
rect 7094 4443 7108 4457
rect 7130 4443 7144 4457
rect 8618 4443 8632 4457
rect 17210 4443 17224 4457
rect 17330 4443 17344 4457
rect 22034 4443 22048 4457
rect 23906 4443 23920 4457
rect 24674 4443 24688 4457
rect 2618 4419 2632 4433
rect 9146 4419 9160 4433
rect 13082 4419 13096 4433
rect 24410 4419 24424 4433
rect 24890 4419 24904 4433
rect 26762 4419 26776 4433
rect 2594 4395 2608 4409
rect 12530 4395 12544 4409
rect 15242 4395 15256 4409
rect 21026 4395 21040 4409
rect 23210 4395 23224 4409
rect 26978 4395 26992 4409
rect 2570 4371 2584 4385
rect 22058 4371 22072 4385
rect 25970 4371 25984 4385
rect 2522 4347 2536 4361
rect 16586 4347 16600 4361
rect 16682 4347 16696 4361
rect 20186 4347 20200 4361
rect 20258 4347 20272 4361
rect 21410 4347 21424 4361
rect 23738 4347 23752 4361
rect 26642 4347 26656 4361
rect 2498 4323 2512 4337
rect 24338 4323 24352 4337
rect 24626 4323 24640 4337
rect 25658 4323 25672 4337
rect 2426 4299 2440 4313
rect 4466 4299 4480 4313
rect 7034 4299 7048 4313
rect 9554 4299 9568 4313
rect 18002 4299 18016 4313
rect 19490 4299 19504 4313
rect 20906 4299 20920 4313
rect 25922 4299 25936 4313
rect 2378 4275 2392 4289
rect 4970 4275 4984 4289
rect 6074 4275 6088 4289
rect 6578 4275 6592 4289
rect 6650 4275 6664 4289
rect 7610 4275 7624 4289
rect 9938 4275 9952 4289
rect 11258 4275 11272 4289
rect 12458 4275 12472 4289
rect 12530 4275 12544 4289
rect 12554 4275 12568 4289
rect 15698 4275 15712 4289
rect 22586 4275 22600 4289
rect 23450 4275 23464 4289
rect 25034 4275 25048 4289
rect 2354 4251 2368 4265
rect 9242 4251 9256 4265
rect 15962 4251 15976 4265
rect 16514 4251 16528 4265
rect 21338 4251 21352 4265
rect 23186 4251 23200 4265
rect 25754 4251 25768 4265
rect 25850 4251 25864 4265
rect 27122 4251 27136 4265
rect 2282 4227 2296 4241
rect 12362 4227 12376 4241
rect 12602 4227 12616 4241
rect 12626 4227 12640 4241
rect 12962 4227 12976 4241
rect 22850 4227 22864 4241
rect 22922 4227 22936 4241
rect 24458 4227 24472 4241
rect 24602 4227 24616 4241
rect 26714 4227 26728 4241
rect 2258 4203 2272 4217
rect 8930 4203 8944 4217
rect 9458 4203 9472 4217
rect 10706 4203 10720 4217
rect 10754 4203 10768 4217
rect 21434 4203 21448 4217
rect 22010 4203 22024 4217
rect 22226 4203 22240 4217
rect 22538 4203 22552 4217
rect 24314 4203 24328 4217
rect 24746 4203 24760 4217
rect 25754 4203 25768 4217
rect 25802 4203 25816 4217
rect 2186 4179 2200 4193
rect 2402 4179 2416 4193
rect 8450 4179 8464 4193
rect 10514 4179 10528 4193
rect 10826 4179 10840 4193
rect 11282 4179 11296 4193
rect 12794 4179 12808 4193
rect 15722 4179 15736 4193
rect 24866 4179 24880 4193
rect 2162 4155 2176 4169
rect 14306 4155 14320 4169
rect 24554 4155 24568 4169
rect 2114 4131 2128 4145
rect 7250 4131 7264 4145
rect 7586 4131 7600 4145
rect 7658 4131 7672 4145
rect 10658 4131 10672 4145
rect 10754 4131 10768 4145
rect 13682 4131 13696 4145
rect 17762 4131 17776 4145
rect 18290 4131 18304 4145
rect 25898 4131 25912 4145
rect 2066 4107 2080 4121
rect 4322 4107 4336 4121
rect 4826 4107 4840 4121
rect 6938 4107 6952 4121
rect 7562 4107 7576 4121
rect 11786 4107 11800 4121
rect 24434 4107 24448 4121
rect 2042 4083 2056 4097
rect 8042 4083 8056 4097
rect 14258 4083 14272 4097
rect 14498 4083 14512 4097
rect 23546 4083 23560 4097
rect 25346 4083 25360 4097
rect 1970 4059 1984 4073
rect 5306 4059 5320 4073
rect 9458 4059 9472 4073
rect 20162 4059 20176 4073
rect 23162 4059 23176 4073
rect 23618 4059 23632 4073
rect 23690 4059 23704 4073
rect 24194 4059 24208 4073
rect 24938 4059 24952 4073
rect 1946 4035 1960 4049
rect 6770 4035 6784 4049
rect 16850 4035 16864 4049
rect 17042 4035 17056 4049
rect 23378 4035 23392 4049
rect 24338 4035 24352 4049
rect 24794 4035 24808 4049
rect 1874 4011 1888 4025
rect 7130 4011 7144 4025
rect 13922 4011 13936 4025
rect 14354 4011 14368 4025
rect 14546 4011 14560 4025
rect 20210 4011 20224 4025
rect 21458 4011 21472 4025
rect 21938 4011 21952 4025
rect 22250 4011 22264 4025
rect 23810 4011 23824 4025
rect 24410 4011 24424 4025
rect 25850 4011 25864 4025
rect 26402 4011 26416 4025
rect 1826 3987 1840 4001
rect 3530 3987 3544 4001
rect 4898 3987 4912 4001
rect 5090 3987 5104 4001
rect 8906 3987 8920 4001
rect 20714 3987 20728 4001
rect 21242 3987 21256 4001
rect 22994 3987 23008 4001
rect 23018 3987 23032 4001
rect 23162 3987 23176 4001
rect 23234 3987 23248 4001
rect 1802 3963 1816 3977
rect 6410 3963 6424 3977
rect 8354 3963 8368 3977
rect 14090 3963 14104 3977
rect 16922 3963 16936 3977
rect 25322 3963 25336 3977
rect 1730 3939 1744 3953
rect 9914 3939 9928 3953
rect 10034 3939 10048 3953
rect 10406 3939 10420 3953
rect 10538 3939 10552 3953
rect 13370 3939 13384 3953
rect 13826 3939 13840 3953
rect 19346 3939 19360 3953
rect 19874 3939 19888 3953
rect 23114 3939 23128 3953
rect 1682 3915 1696 3929
rect 9890 3915 9904 3929
rect 10130 3915 10144 3929
rect 21650 3915 21664 3929
rect 1658 3891 1672 3905
rect 16778 3891 16792 3905
rect 17234 3891 17248 3905
rect 19538 3891 19552 3905
rect 19898 3891 19912 3905
rect 20318 3891 20332 3905
rect 21650 3891 21664 3905
rect 22082 3891 22096 3905
rect 1634 3867 1648 3881
rect 4178 3867 4192 3881
rect 5714 3867 5728 3881
rect 7706 3867 7720 3881
rect 7754 3867 7768 3881
rect 8906 3867 8920 3881
rect 10394 3867 10408 3881
rect 11282 3867 11296 3881
rect 25610 3867 25624 3881
rect 1610 3843 1624 3857
rect 24050 3843 24064 3857
rect 70 3819 84 3833
rect 8186 3819 8200 3833
rect 12002 3819 12016 3833
rect 17282 3819 17296 3833
rect 17690 3819 17704 3833
rect 19274 3819 19288 3833
rect 19634 3819 19648 3833
rect 20090 3819 20104 3833
rect 24530 3819 24544 3833
rect 70 3795 84 3809
rect 19946 3795 19960 3809
rect 24050 3795 24064 3809
rect 25250 3795 25264 3809
rect 1610 3771 1624 3785
rect 3170 3771 3184 3785
rect 3266 3771 3280 3785
rect 3314 3771 3328 3785
rect 7730 3771 7744 3785
rect 13298 3771 13312 3785
rect 14234 3771 14248 3785
rect 15314 3771 15328 3785
rect 17906 3771 17920 3785
rect 19082 3771 19096 3785
rect 19754 3771 19768 3785
rect 21122 3771 21136 3785
rect 23090 3771 23104 3785
rect 23402 3771 23416 3785
rect 26138 3771 26152 3785
rect 1634 3747 1648 3761
rect 3290 3747 3304 3761
rect 4946 3747 4960 3761
rect 5594 3747 5608 3761
rect 6506 3747 6520 3761
rect 6554 3747 6568 3761
rect 7586 3747 7600 3761
rect 8258 3747 8272 3761
rect 9098 3747 9112 3761
rect 9674 3747 9688 3761
rect 10082 3747 10096 3761
rect 12986 3747 13000 3761
rect 15122 3747 15136 3761
rect 16250 3747 16264 3761
rect 21266 3747 21280 3761
rect 21482 3747 21496 3761
rect 21554 3747 21568 3761
rect 23042 3747 23056 3761
rect 23378 3747 23392 3761
rect 23594 3747 23608 3761
rect 1658 3723 1672 3737
rect 2306 3723 2320 3737
rect 12458 3723 12472 3737
rect 13106 3723 13120 3737
rect 13322 3723 13336 3737
rect 13850 3723 13864 3737
rect 17618 3723 17632 3737
rect 17666 3723 17680 3737
rect 17798 3723 17812 3737
rect 19322 3723 19336 3737
rect 20042 3723 20056 3737
rect 21122 3723 21136 3737
rect 21674 3723 21688 3737
rect 1706 3699 1720 3713
rect 4538 3699 4552 3713
rect 4610 3699 4624 3713
rect 5378 3699 5392 3713
rect 14402 3699 14416 3713
rect 14594 3699 14608 3713
rect 17714 3699 17728 3713
rect 1754 3675 1768 3689
rect 17906 3675 17920 3689
rect 1922 3651 1936 3665
rect 14450 3651 14464 3665
rect 14714 3651 14728 3665
rect 15098 3651 15112 3665
rect 15146 3651 15160 3665
rect 21962 3651 21976 3665
rect 2210 3627 2224 3641
rect 14858 3627 14872 3641
rect 15530 3627 15544 3641
rect 27146 3627 27160 3641
rect 2210 3603 2224 3617
rect 4202 3603 4216 3617
rect 5618 3603 5632 3617
rect 6842 3603 6856 3617
rect 7922 3603 7936 3617
rect 10202 3603 10216 3617
rect 12650 3603 12664 3617
rect 12986 3603 13000 3617
rect 13706 3603 13720 3617
rect 14114 3603 14128 3617
rect 24026 3603 24040 3617
rect 2258 3579 2272 3593
rect 6482 3579 6496 3593
rect 7058 3579 7072 3593
rect 10586 3579 10600 3593
rect 21866 3579 21880 3593
rect 21986 3579 22000 3593
rect 25514 3579 25528 3593
rect 2450 3555 2464 3569
rect 6698 3555 6712 3569
rect 7490 3555 7504 3569
rect 10370 3555 10384 3569
rect 11186 3555 11200 3569
rect 12242 3555 12256 3569
rect 13898 3555 13912 3569
rect 14330 3555 14344 3569
rect 16970 3555 16984 3569
rect 21818 3555 21832 3569
rect 24026 3555 24040 3569
rect 24074 3555 24088 3569
rect 2474 3531 2488 3545
rect 17618 3531 17632 3545
rect 17714 3531 17728 3545
rect 24002 3531 24016 3545
rect 2522 3507 2536 3521
rect 2834 3507 2848 3521
rect 4682 3507 4696 3521
rect 8882 3507 8896 3521
rect 16082 3507 16096 3521
rect 16874 3507 16888 3521
rect 17498 3507 17512 3521
rect 20402 3507 20416 3521
rect 2546 3483 2560 3497
rect 2786 3483 2800 3497
rect 2954 3483 2968 3497
rect 4994 3483 5008 3497
rect 6290 3483 6304 3497
rect 8762 3483 8776 3497
rect 9218 3483 9232 3497
rect 13898 3483 13912 3497
rect 14714 3483 14728 3497
rect 16898 3483 16912 3497
rect 20546 3483 20560 3497
rect 21794 3483 21808 3497
rect 24146 3483 24160 3497
rect 24482 3483 24496 3497
rect 2570 3459 2584 3473
rect 3818 3459 3832 3473
rect 13250 3459 13264 3473
rect 25706 3459 25720 3473
rect 2594 3435 2608 3449
rect 19394 3435 19408 3449
rect 20402 3435 20416 3449
rect 24722 3435 24736 3449
rect 2666 3411 2680 3425
rect 11618 3411 11632 3425
rect 12122 3411 12136 3425
rect 20810 3411 20824 3425
rect 2738 3387 2752 3401
rect 5834 3387 5848 3401
rect 5978 3387 5992 3401
rect 14738 3387 14752 3401
rect 16034 3387 16048 3401
rect 18050 3387 18064 3401
rect 23522 3387 23536 3401
rect 2810 3363 2824 3377
rect 6266 3363 6280 3377
rect 13034 3363 13048 3377
rect 22730 3363 22744 3377
rect 27026 3363 27040 3377
rect 2954 3339 2968 3353
rect 14522 3339 14536 3353
rect 15698 3339 15712 3353
rect 21890 3339 21904 3353
rect 24254 3339 24268 3353
rect 3098 3315 3112 3329
rect 7346 3315 7360 3329
rect 7394 3315 7408 3329
rect 16946 3315 16960 3329
rect 24290 3315 24304 3329
rect 3218 3291 3232 3305
rect 18098 3291 18112 3305
rect 3362 3267 3376 3281
rect 3410 3267 3424 3281
rect 3746 3267 3760 3281
rect 10106 3267 10120 3281
rect 12746 3267 12760 3281
rect 17258 3267 17272 3281
rect 18410 3267 18424 3281
rect 25394 3267 25408 3281
rect 3530 3243 3544 3257
rect 3866 3243 3880 3257
rect 6674 3243 6688 3257
rect 8786 3243 8800 3257
rect 18026 3243 18040 3257
rect 19658 3243 19672 3257
rect 3554 3219 3568 3233
rect 4586 3219 4600 3233
rect 4658 3219 4672 3233
rect 6746 3219 6760 3233
rect 7322 3219 7336 3233
rect 7418 3219 7432 3233
rect 7874 3219 7888 3233
rect 16754 3219 16768 3233
rect 19298 3219 19312 3233
rect 19418 3219 19432 3233
rect 24314 3219 24328 3233
rect 25010 3219 25024 3233
rect 3554 3195 3568 3209
rect 26786 3195 26800 3209
rect 3602 3171 3616 3185
rect 24098 3171 24112 3185
rect 26786 3171 26800 3185
rect 26834 3171 26848 3185
rect 3602 3147 3616 3161
rect 5162 3147 5176 3161
rect 8282 3147 8296 3161
rect 8570 3147 8584 3161
rect 9746 3147 9760 3161
rect 15026 3147 15040 3161
rect 17114 3147 17128 3161
rect 17786 3147 17800 3161
rect 18026 3147 18040 3161
rect 18722 3147 18736 3161
rect 19418 3147 19432 3161
rect 19706 3147 19720 3161
rect 3626 3123 3640 3137
rect 8954 3123 8968 3137
rect 20354 3123 20368 3137
rect 22706 3123 22720 3137
rect 23354 3123 23368 3137
rect 3650 3099 3664 3113
rect 19826 3099 19840 3113
rect 20570 3099 20584 3113
rect 22106 3099 22120 3113
rect 23810 3099 23824 3113
rect 3722 3075 3736 3089
rect 3842 3075 3856 3089
rect 4346 3075 4360 3089
rect 16802 3075 16816 3089
rect 21626 3075 21640 3089
rect 3770 3051 3784 3065
rect 4658 3051 4672 3065
rect 14834 3051 14848 3065
rect 21002 3051 21016 3065
rect 3866 3027 3880 3041
rect 5882 3027 5896 3041
rect 6026 3027 6040 3041
rect 6722 3027 6736 3041
rect 9650 3027 9664 3041
rect 13922 3027 13936 3041
rect 14186 3027 14200 3041
rect 15578 3027 15592 3041
rect 17930 3027 17944 3041
rect 20354 3027 20368 3041
rect 20858 3027 20872 3041
rect 3890 3003 3904 3017
rect 20114 3003 20128 3017
rect 3890 2979 3904 2993
rect 7370 2979 7384 2993
rect 12818 2979 12832 2993
rect 24242 2979 24256 2993
rect 3914 2955 3928 2969
rect 27493 2955 27507 2969
rect 3986 2931 4000 2945
rect 10274 2931 10288 2945
rect 10322 2931 10336 2945
rect 14882 2931 14896 2945
rect 15770 2931 15784 2945
rect 20426 2931 20440 2945
rect 4034 2907 4048 2921
rect 11186 2907 11200 2921
rect 11258 2907 11272 2921
rect 26930 2907 26944 2921
rect 4034 2883 4048 2897
rect 12098 2883 12112 2897
rect 14978 2883 14992 2897
rect 17258 2883 17272 2897
rect 17642 2883 17656 2897
rect 4082 2859 4096 2873
rect 10154 2859 10168 2873
rect 19970 2859 19984 2873
rect 24722 2859 24736 2873
rect 4202 2835 4216 2849
rect 19562 2835 19576 2849
rect 20378 2835 20392 2849
rect 26258 2835 26272 2849
rect 4442 2811 4456 2825
rect 20786 2811 20800 2825
rect 4490 2787 4504 2801
rect 10898 2787 10912 2801
rect 11018 2787 11032 2801
rect 21302 2787 21316 2801
rect 4754 2763 4768 2777
rect 15866 2763 15880 2777
rect 20378 2763 20392 2777
rect 21074 2763 21088 2777
rect 4994 2739 5008 2753
rect 9962 2739 9976 2753
rect 10154 2739 10168 2753
rect 16634 2739 16648 2753
rect 5066 2715 5080 2729
rect 5126 2715 5140 2729
rect 5162 2715 5176 2729
rect 9002 2715 9016 2729
rect 20762 2715 20776 2729
rect 23666 2715 23680 2729
rect 5138 2691 5152 2705
rect 6986 2691 7000 2705
rect 25178 2691 25192 2705
rect 5210 2667 5224 2681
rect 18770 2667 18784 2681
rect 5258 2643 5272 2657
rect 6314 2643 6328 2657
rect 12770 2643 12784 2657
rect 20282 2643 20296 2657
rect 24818 2643 24832 2657
rect 26450 2643 26464 2657
rect 5522 2619 5536 2633
rect 5978 2619 5992 2633
rect 6098 2619 6112 2633
rect 16634 2619 16648 2633
rect 5786 2595 5800 2609
rect 12722 2595 12736 2609
rect 12818 2595 12832 2609
rect 21206 2595 21220 2609
rect 5834 2571 5848 2585
rect 12890 2571 12904 2585
rect 26354 2571 26368 2585
rect 6098 2547 6112 2561
rect 20450 2547 20464 2561
rect 6146 2523 6160 2537
rect 25778 2523 25792 2537
rect 6314 2499 6328 2513
rect 8162 2499 8176 2513
rect 8474 2499 8488 2513
rect 8666 2499 8680 2513
rect 10010 2499 10024 2513
rect 10922 2499 10936 2513
rect 12554 2499 12568 2513
rect 13490 2499 13504 2513
rect 14378 2499 14392 2513
rect 15842 2499 15856 2513
rect 21362 2499 21376 2513
rect 25946 2499 25960 2513
rect 6338 2475 6352 2489
rect 16802 2475 16816 2489
rect 20450 2475 20464 2489
rect 26186 2475 26200 2489
rect 6482 2451 6496 2465
rect 21506 2451 21520 2465
rect 25778 2451 25792 2465
rect 26810 2451 26824 2465
rect 6602 2427 6616 2441
rect 14954 2427 14968 2441
rect 6794 2403 6808 2417
rect 8978 2403 8992 2417
rect 26306 2403 26320 2417
rect 6842 2379 6856 2393
rect 21722 2379 21736 2393
rect 6962 2355 6976 2369
rect 10682 2355 10696 2369
rect 10850 2355 10864 2369
rect 17378 2355 17392 2369
rect 7178 2331 7192 2345
rect 7274 2331 7288 2345
rect 9338 2331 9352 2345
rect 9986 2331 10000 2345
rect 11042 2331 11056 2345
rect 13394 2331 13408 2345
rect 13466 2331 13480 2345
rect 13970 2331 13984 2345
rect 14282 2331 14296 2345
rect 16994 2331 17008 2345
rect 17882 2331 17896 2345
rect 20594 2331 20608 2345
rect 22850 2331 22864 2345
rect 7250 2307 7264 2321
rect 7442 2307 7456 2321
rect 7490 2307 7504 2321
rect 7514 2307 7528 2321
rect 7754 2307 7768 2321
rect 21602 2307 21616 2321
rect 7418 2283 7432 2297
rect 10874 2283 10888 2297
rect 11114 2283 11128 2297
rect 25634 2283 25648 2297
rect 7466 2259 7480 2273
rect 9746 2259 9760 2273
rect 10586 2259 10600 2273
rect 19466 2259 19480 2273
rect 24626 2259 24640 2273
rect 25418 2259 25432 2273
rect 7514 2235 7528 2249
rect 9842 2235 9856 2249
rect 10178 2235 10192 2249
rect 25586 2235 25600 2249
rect 7802 2211 7816 2225
rect 17474 2211 17488 2225
rect 7970 2187 7984 2201
rect 8210 2187 8224 2201
rect 14738 2187 14752 2201
rect 22418 2187 22432 2201
rect 8186 2163 8200 2177
rect 9434 2163 9448 2177
rect 15098 2163 15112 2177
rect 22370 2163 22384 2177
rect 8234 2139 8248 2153
rect 8882 2139 8896 2153
rect 9122 2139 9136 2153
rect 9770 2139 9784 2153
rect 12314 2139 12328 2153
rect 13010 2139 13024 2153
rect 21698 2139 21712 2153
rect 8354 2115 8368 2129
rect 9482 2115 9496 2129
rect 9530 2115 9544 2129
rect 15050 2115 15064 2129
rect 16994 2115 17008 2129
rect 17066 2115 17080 2129
rect 8714 2091 8728 2105
rect 9182 2091 9196 2105
rect 9218 2091 9232 2105
rect 17090 2091 17104 2105
rect 20138 2091 20152 2105
rect 22778 2091 22792 2105
rect 8762 2067 8776 2081
rect 13418 2067 13432 2081
rect 13946 2067 13960 2081
rect 14006 2067 14020 2081
rect 14042 2067 14056 2081
rect 14666 2067 14680 2081
rect 14978 2067 14992 2081
rect 15170 2067 15184 2081
rect 8786 2043 8800 2057
rect 19250 2043 19264 2057
rect 21170 2043 21184 2057
rect 9002 2019 9016 2033
rect 9050 2019 9064 2033
rect 9170 2019 9184 2033
rect 9866 2019 9880 2033
rect 10274 2019 10288 2033
rect 10622 2019 10636 2033
rect 11162 2019 11176 2033
rect 11714 2019 11728 2033
rect 12266 2019 12280 2033
rect 24506 2019 24520 2033
rect 9050 1995 9064 2009
rect 10106 1995 10120 2009
rect 14618 1995 14632 2009
rect 22802 1995 22816 2009
rect 23258 1995 23272 2009
rect 9242 1971 9256 1985
rect 9278 1971 9292 1985
rect 9386 1971 9400 1985
rect 17882 1971 17896 1985
rect 21578 1971 21592 1985
rect 9386 1947 9400 1961
rect 26546 1947 26560 1961
rect 9482 1923 9496 1937
rect 16442 1923 16456 1937
rect 9530 1899 9544 1913
rect 17978 1899 17992 1913
rect 9578 1875 9592 1889
rect 15218 1875 15232 1889
rect 9578 1851 9592 1865
rect 17570 1851 17584 1865
rect 9794 1827 9808 1841
rect 17738 1827 17752 1841
rect 9866 1803 9880 1817
rect 24986 1803 25000 1817
rect 10322 1779 10336 1793
rect 24506 1779 24520 1793
rect 24962 1779 24976 1793
rect 10370 1755 10384 1769
rect 10778 1755 10792 1769
rect 11210 1755 11224 1769
rect 19370 1755 19384 1769
rect 27098 1755 27112 1769
rect 10418 1731 10432 1745
rect 10682 1731 10696 1745
rect 21842 1731 21856 1745
rect 10610 1707 10624 1721
rect 12926 1707 12940 1721
rect 18434 1707 18448 1721
rect 19058 1707 19072 1721
rect 24842 1707 24856 1721
rect 25442 1707 25456 1721
rect 26378 1707 26392 1721
rect 11354 1683 11368 1697
rect 11426 1683 11440 1697
rect 11498 1683 11512 1697
rect 19442 1683 19456 1697
rect 21842 1683 21856 1697
rect 22202 1683 22216 1697
rect 11402 1659 11416 1673
rect 24698 1659 24712 1673
rect 12746 1635 12760 1649
rect 12842 1635 12856 1649
rect 13154 1635 13168 1649
rect 13178 1635 13192 1649
rect 13346 1635 13360 1649
rect 13538 1635 13552 1649
rect 13994 1635 14008 1649
rect 24362 1635 24376 1649
rect 13418 1611 13432 1625
rect 13586 1611 13600 1625
rect 14258 1611 14272 1625
rect 18818 1611 18832 1625
rect 24650 1611 24664 1625
rect 14522 1587 14536 1601
rect 15074 1587 15088 1601
rect 17570 1587 17584 1601
rect 17858 1587 17872 1601
rect 27146 1587 27160 1601
rect 27493 1587 27507 1601
rect 14666 1563 14680 1577
rect 14690 1563 14704 1577
rect 27122 1563 27136 1577
rect 27493 1563 27507 1577
rect 17162 730 17176 744
rect 22274 730 22288 744
rect 13010 706 13024 720
rect 22922 706 22936 720
rect 12914 682 12928 696
rect 14018 682 14032 696
rect 15386 682 15400 696
rect 26642 682 26656 696
rect 12482 658 12496 672
rect 13754 658 13768 672
rect 15266 658 15280 672
rect 17690 658 17704 672
rect 18002 658 18016 672
rect 25802 658 25816 672
rect 11450 634 11464 648
rect 20546 634 20560 648
rect 20978 634 20992 648
rect 23738 634 23752 648
rect 10970 610 10984 624
rect 21002 610 21016 624
rect 21218 610 21232 624
rect 25898 610 25912 624
rect 10202 586 10216 600
rect 26018 586 26032 600
rect 9626 562 9640 576
rect 25010 562 25024 576
rect 9554 538 9568 552
rect 13586 538 13600 552
rect 13682 538 13696 552
rect 13802 538 13816 552
rect 14882 538 14896 552
rect 22322 538 22336 552
rect 9434 514 9448 528
rect 21482 514 21496 528
rect 8042 490 8056 504
rect 17522 490 17536 504
rect 17810 490 17824 504
rect 24266 490 24280 504
rect 7994 466 8008 480
rect 14906 466 14920 480
rect 15098 466 15112 480
rect 22082 466 22096 480
rect 7370 442 7384 456
rect 21290 442 21304 456
rect 7082 418 7096 432
rect 23690 418 23704 432
rect 26786 418 26800 432
rect 27493 418 27507 432
rect 6746 394 6760 408
rect 15194 394 15208 408
rect 22490 394 22504 408
rect 22946 394 22960 408
rect 24770 394 24784 408
rect 24962 394 24976 408
rect 24986 394 25000 408
rect 26738 394 26752 408
rect 27493 394 27507 408
rect 6218 370 6232 384
rect 13778 370 13792 384
rect 14354 370 14368 384
rect 17978 370 17992 384
rect 18314 370 18328 384
rect 23978 370 23992 384
rect 24938 370 24952 384
rect 26570 370 26584 384
rect 26786 370 26800 384
rect 6050 346 6064 360
rect 8570 346 8584 360
rect 9914 346 9928 360
rect 9962 346 9976 360
rect 18218 346 18232 360
rect 18338 346 18352 360
rect 24986 346 25000 360
rect 5426 322 5440 336
rect 14066 322 14080 336
rect 15482 322 15496 336
rect 25082 322 25096 336
rect 5282 298 5296 312
rect 7682 298 7696 312
rect 7802 298 7816 312
rect 20882 298 20896 312
rect 21530 298 21544 312
rect 5090 274 5104 288
rect 15338 274 15352 288
rect 16226 274 16240 288
rect 18986 274 19000 288
rect 19922 274 19936 288
rect 24674 274 24688 288
rect 4754 250 4768 264
rect 8282 250 8296 264
rect 8642 250 8656 264
rect 23546 250 23560 264
rect 4490 226 4504 240
rect 24866 226 24880 240
rect 4130 202 4144 216
rect 6386 202 6400 216
rect 6434 202 6448 216
rect 26690 202 26704 216
rect 3506 178 3520 192
rect 12770 178 12784 192
rect 15818 178 15832 192
rect 22634 178 22648 192
rect 22826 178 22840 192
rect 2834 154 2848 168
rect 4610 154 4624 168
rect 4706 154 4720 168
rect 10634 154 10648 168
rect 10922 154 10936 168
rect 11066 154 11080 168
rect 11114 154 11128 168
rect 11306 154 11320 168
rect 17858 154 17872 168
rect 18578 154 18592 168
rect 23090 154 23104 168
rect 2714 130 2728 144
rect 3674 130 3688 144
rect 3746 130 3760 144
rect 8834 130 8848 144
rect 9266 130 9280 144
rect 19250 130 19264 144
rect 20042 130 20056 144
rect 23282 130 23296 144
rect 2690 106 2704 120
rect 6338 106 6352 120
rect 6410 106 6424 120
rect 7634 106 7648 120
rect 7946 106 7960 120
rect 12170 106 12184 120
rect 12386 106 12400 120
rect 13538 106 13552 120
rect 16826 106 16840 120
rect 25202 106 25216 120
rect 70 82 84 96
rect 1730 82 1744 96
rect 1850 82 1864 96
rect 4778 82 4792 96
rect 5042 82 5056 96
rect 13466 82 13480 96
rect 13514 82 13528 96
rect 21602 82 21616 96
rect 70 58 84 72
rect 23042 58 23056 72
rect 5978 34 5992 48
rect 27493 34 27507 48
rect 17426 10 17440 24
rect 20138 10 20152 24
rect 21962 10 21976 24
rect 26786 10 26800 24
rect 27493 10 27507 24
<< metal2 >>
rect 0 7917 70 7929
rect 0 7893 70 7905
rect 123 7714 323 7988
rect 339 7714 351 7988
rect 363 7714 375 7988
rect 387 7714 399 7988
rect 411 7714 423 7988
rect 1707 7714 1719 7916
rect 1755 7714 1767 7892
rect 1995 7714 2007 7916
rect 2187 7714 2199 7892
rect 2379 7714 2391 7940
rect 2415 7882 2427 7988
rect 2451 7954 2463 7988
rect 3303 7906 3315 7988
rect 3651 7714 3663 7892
rect 3939 7714 3951 7940
rect 4395 7714 4407 7844
rect 4971 7834 4983 7988
rect 5403 7714 5415 7964
rect 5823 7810 5835 7988
rect 5859 7978 5871 7988
rect 7443 7714 7455 7964
rect 7527 7786 7539 7988
rect 8379 7786 8391 7988
rect 7995 7714 8007 7772
rect 9231 7762 9243 7988
rect 10083 7882 10095 7988
rect 9651 7714 9663 7820
rect 9987 7714 9999 7868
rect 10935 7834 10947 7988
rect 11787 7810 11799 7988
rect 11823 7906 11835 7988
rect 13491 7906 13503 7988
rect 10899 7714 10911 7796
rect 11787 7714 11799 7772
rect 13611 7714 13623 7772
rect 14343 7738 14355 7988
rect 14367 7930 14379 7988
rect 16023 7882 16035 7988
rect 16695 7882 16707 7988
rect 16696 7868 16714 7882
rect 14571 7714 14583 7868
rect 14907 7714 14919 7820
rect 15555 7714 15567 7820
rect 16443 7714 16455 7868
rect 16683 7714 16695 7868
rect 16899 7714 16911 7892
rect 17631 7882 17643 7988
rect 18543 7882 18555 7988
rect 19263 7882 19275 7988
rect 17632 7868 17650 7882
rect 19264 7868 19282 7882
rect 17619 7714 17631 7868
rect 17835 7714 17847 7796
rect 18723 7714 18735 7796
rect 18771 7714 18783 7868
rect 19251 7714 19263 7868
rect 19767 7762 19779 7988
rect 20247 7810 20259 7988
rect 21087 7810 21099 7988
rect 21927 7954 21939 7988
rect 22767 7834 22779 7988
rect 24423 7882 24435 7988
rect 21088 7796 21106 7810
rect 19768 7748 19786 7762
rect 19707 7714 19719 7748
rect 19755 7714 19767 7748
rect 21075 7714 21087 7796
rect 22659 7714 22671 7796
rect 23211 7714 23223 7724
rect 23571 7714 23583 7820
rect 24447 7786 24459 7988
rect 25287 7810 25299 7988
rect 26127 7834 26139 7988
rect 24795 7714 24807 7772
rect 25035 7714 25047 7748
rect 26355 7714 26367 7868
rect 27099 7714 27111 7820
rect 27123 7738 27135 7844
rect 27147 7786 27159 7796
rect 27171 7786 27183 7964
rect 27243 7714 27443 7988
rect 27507 7821 27577 7833
rect 27507 7797 27577 7809
rect 27507 7773 27577 7785
rect 27507 7749 27577 7761
rect 27507 7725 27577 7737
rect 0 3820 70 3832
rect 0 3796 70 3808
rect 123 1553 323 6915
rect 339 1553 351 6915
rect 363 1553 375 6915
rect 387 1553 399 6915
rect 411 1553 423 6915
rect 1611 3857 1623 6915
rect 1635 3881 1647 6915
rect 1659 3905 1671 6915
rect 1611 1553 1623 3771
rect 1635 1553 1647 3747
rect 1659 1553 1671 3723
rect 1683 1553 1695 3915
rect 1707 3713 1719 6915
rect 1731 1553 1743 3939
rect 1755 3689 1767 6915
rect 1803 3977 1815 6915
rect 1827 4001 1839 6915
rect 1875 4025 1887 6915
rect 1923 3665 1935 6915
rect 1947 4049 1959 6915
rect 1971 4073 1983 6915
rect 2043 4097 2055 6915
rect 2067 4121 2079 6915
rect 2115 4145 2127 6915
rect 2163 4169 2175 6915
rect 2187 4193 2199 6915
rect 2211 3641 2223 6915
rect 2259 4217 2271 6915
rect 2283 4241 2295 6915
rect 2307 3737 2319 6915
rect 2355 4265 2367 6915
rect 2379 4289 2391 6915
rect 2427 4313 2439 6915
rect 2211 1553 2223 3603
rect 2259 1553 2271 3579
rect 2403 1553 2415 4179
rect 2451 1553 2463 3555
rect 2475 3545 2487 6915
rect 2499 4337 2511 6915
rect 2523 4361 2535 6915
rect 2571 4385 2583 6915
rect 2595 4409 2607 6915
rect 2619 4433 2631 6915
rect 2667 4481 2679 6915
rect 2691 4505 2703 6915
rect 2715 4529 2727 6915
rect 2739 4553 2751 6915
rect 2763 4577 2775 6915
rect 2811 4601 2823 6915
rect 2523 1553 2535 3507
rect 2547 1553 2559 3483
rect 2571 1553 2583 3459
rect 2595 1553 2607 3435
rect 2643 1553 2655 4443
rect 2835 3521 2847 6915
rect 2859 4625 2871 6915
rect 2907 4649 2919 6915
rect 2955 3497 2967 6915
rect 3027 4673 3039 6915
rect 3051 4697 3063 6915
rect 2667 1553 2679 3411
rect 2739 1553 2751 3387
rect 2787 1553 2799 3483
rect 2811 1553 2823 3363
rect 2955 1553 2967 3339
rect 3099 3329 3111 6915
rect 3147 4721 3159 6915
rect 3171 3785 3183 6915
rect 3219 3305 3231 6915
rect 3267 3785 3279 6915
rect 3291 3761 3303 6915
rect 3315 4745 3327 6915
rect 3339 4769 3351 6915
rect 3363 4793 3375 6915
rect 3315 1553 3327 3771
rect 3411 3281 3423 6915
rect 3435 4817 3447 6915
rect 3459 4841 3471 6915
rect 3507 4865 3519 6915
rect 3531 4001 3543 6915
rect 3363 1553 3375 3267
rect 3531 1553 3543 3243
rect 3555 3233 3567 6915
rect 3555 1553 3567 3195
rect 3603 3185 3615 6915
rect 3723 4889 3735 6915
rect 3747 3281 3759 6915
rect 3771 4913 3783 6915
rect 3603 1553 3615 3147
rect 3627 1553 3639 3123
rect 3651 1553 3663 3099
rect 3723 1553 3735 3075
rect 3771 1553 3783 3051
rect 3795 1553 3807 4923
rect 3819 3473 3831 6915
rect 3843 4961 3855 6915
rect 3867 3257 3879 6915
rect 3843 1553 3855 3075
rect 3867 1553 3879 3027
rect 3891 3017 3903 6915
rect 3939 4937 3951 6915
rect 3891 1553 3903 2979
rect 3915 1553 3927 2955
rect 3963 1553 3975 4971
rect 3987 4937 3999 6915
rect 4011 4505 4023 6915
rect 3987 1553 3999 2931
rect 4035 2921 4047 6915
rect 4083 5009 4095 6915
rect 4131 5057 4143 6915
rect 4035 1553 4047 2883
rect 4083 1553 4095 2859
rect 4107 1553 4119 5019
rect 4179 1553 4191 3867
rect 4203 3617 4215 6915
rect 4227 4553 4239 6915
rect 4275 5081 4287 6915
rect 4323 5105 4335 6915
rect 4203 1553 4215 2835
rect 4251 1553 4263 4731
rect 4299 1553 4311 4683
rect 4323 1553 4335 4107
rect 4347 3089 4359 6915
rect 4371 5129 4383 6915
rect 4419 1553 4431 5139
rect 4443 2825 4455 6915
rect 4467 4313 4479 6915
rect 4491 2801 4503 6915
rect 4539 5201 4551 6915
rect 4515 1553 4527 5163
rect 4563 4529 4575 6915
rect 4611 3713 4623 6915
rect 4539 1553 4551 3699
rect 4659 3233 4671 6915
rect 4683 3521 4695 6915
rect 4707 5225 4719 6915
rect 4587 1553 4599 3219
rect 4659 1553 4671 3051
rect 4731 1553 4743 5235
rect 4755 2777 4767 6915
rect 4779 5273 4791 6915
rect 4803 5297 4815 6915
rect 4851 5321 4863 6915
rect 4899 5345 4911 6915
rect 4971 5369 4983 6915
rect 4995 5393 5007 6915
rect 5019 5417 5031 6915
rect 4827 1553 4839 4107
rect 4851 1553 4863 4683
rect 4899 1553 4911 3987
rect 4947 1553 4959 3747
rect 4971 1553 4983 4275
rect 4995 3497 5007 5355
rect 5067 4505 5079 6915
rect 5091 4001 5103 6915
rect 5115 5369 5127 6915
rect 4995 1553 5007 2739
rect 5127 2729 5139 5331
rect 5163 3161 5175 6915
rect 5187 4721 5199 6915
rect 5211 4889 5223 6915
rect 5259 5345 5271 6915
rect 5307 5441 5319 6915
rect 5067 1553 5079 2715
rect 5139 1553 5151 2691
rect 5163 1553 5175 2715
rect 5211 1553 5223 2667
rect 5259 1553 5271 2643
rect 5307 1553 5319 4059
rect 5379 3713 5391 6915
rect 5403 5465 5415 6915
rect 5451 5489 5463 6915
rect 5499 5513 5511 6915
rect 5523 2633 5535 6915
rect 5547 5537 5559 6915
rect 5595 3761 5607 6915
rect 5619 3617 5631 6915
rect 5643 5561 5655 6915
rect 5691 4817 5703 6915
rect 5715 3881 5727 6915
rect 5739 5585 5751 6915
rect 5763 5609 5775 6915
rect 5787 5633 5799 6915
rect 5835 3401 5847 6915
rect 5883 3041 5895 6915
rect 5955 5369 5967 6915
rect 5979 3401 5991 6915
rect 6027 5201 6039 6915
rect 6075 5369 6087 6915
rect 5787 1553 5799 2595
rect 5835 1553 5847 2571
rect 5979 1553 5991 2619
rect 6027 1553 6039 3027
rect 6075 1553 6087 4275
rect 6099 2633 6111 6915
rect 6147 5609 6159 6915
rect 6195 5681 6207 6915
rect 6219 5705 6231 6915
rect 6243 5729 6255 6915
rect 6291 5753 6303 6915
rect 6315 5777 6327 6915
rect 6099 1553 6111 2547
rect 6147 1553 6159 2523
rect 6171 1553 6183 5643
rect 6267 1553 6279 3363
rect 6291 1553 6303 3483
rect 6315 2657 6327 5739
rect 6315 1553 6327 2499
rect 6339 2489 6351 6915
rect 6387 4865 6399 6915
rect 6411 3977 6423 6915
rect 6435 5753 6447 6915
rect 6459 1553 6471 5787
rect 6483 3593 6495 6915
rect 6507 3761 6519 6915
rect 6555 5825 6567 6915
rect 6603 5849 6615 6915
rect 6627 5057 6639 6915
rect 6651 5873 6663 6915
rect 6675 5345 6687 6915
rect 6723 5441 6735 6915
rect 6483 1553 6495 2451
rect 6531 1553 6543 4683
rect 6555 1553 6567 3747
rect 6579 1553 6591 4275
rect 6603 1553 6615 2427
rect 6651 1553 6663 4275
rect 6675 1553 6687 3243
rect 6699 1553 6711 3555
rect 6747 3233 6759 6915
rect 6771 4049 6783 6915
rect 6819 5897 6831 6915
rect 6723 1553 6735 3027
rect 6795 1553 6807 2403
rect 6819 1553 6831 4755
rect 6843 3617 6855 6915
rect 6867 4457 6879 6915
rect 6843 1553 6855 2379
rect 6891 1553 6903 4683
rect 6915 4505 6927 6915
rect 6939 4529 6951 6915
rect 6963 4481 6975 6915
rect 6915 1553 6927 4443
rect 6939 1553 6951 4107
rect 6987 2705 6999 6915
rect 7035 5921 7047 6915
rect 6963 1553 6975 2355
rect 7011 1553 7023 5811
rect 7035 1553 7047 4299
rect 7059 3593 7071 6915
rect 7083 5801 7095 6915
rect 7095 4457 7107 5691
rect 7131 4457 7143 6915
rect 7179 5801 7191 6915
rect 7131 1553 7143 4011
rect 7155 1553 7167 4803
rect 7179 1553 7191 2331
rect 7203 1553 7215 5931
rect 7251 4145 7263 6915
rect 7275 5969 7287 6915
rect 7251 1553 7263 2307
rect 7275 1553 7287 2331
rect 7299 1553 7311 4995
rect 7323 3233 7335 6915
rect 7347 1553 7359 3315
rect 7371 2993 7383 6915
rect 7395 3329 7407 6915
rect 7419 3233 7431 6915
rect 7443 2321 7455 4539
rect 7491 3569 7503 6915
rect 7515 5993 7527 6915
rect 7539 6017 7551 6915
rect 7515 2321 7527 4827
rect 7587 4145 7599 6915
rect 7611 6041 7623 6915
rect 7635 5465 7647 6915
rect 7419 1553 7431 2283
rect 7467 1553 7479 2259
rect 7491 1553 7503 2307
rect 7515 1553 7527 2235
rect 7563 1553 7575 4107
rect 7587 1553 7599 3747
rect 7611 1553 7623 4275
rect 7659 4145 7671 6915
rect 7707 6065 7719 6915
rect 7707 1553 7719 3867
rect 7731 3785 7743 6915
rect 7755 3881 7767 6915
rect 7779 6089 7791 6915
rect 7755 1553 7767 2307
rect 7803 2225 7815 6915
rect 7851 6113 7863 6915
rect 7875 6137 7887 6915
rect 7899 6161 7911 6915
rect 7923 6185 7935 6915
rect 7947 6209 7959 6915
rect 7827 1553 7839 5811
rect 7851 1553 7863 4707
rect 7995 4697 8007 6915
rect 7875 1553 7887 3219
rect 7923 1553 7935 3603
rect 7947 1553 7959 4515
rect 8043 4097 8055 6915
rect 7971 1553 7983 2187
rect 8067 1553 8079 4491
rect 8091 1553 8103 6219
rect 8115 5969 8127 6915
rect 8139 6257 8151 6915
rect 8163 6281 8175 6915
rect 8139 1553 8151 4467
rect 8187 3833 8199 6915
rect 8211 6305 8223 6915
rect 8163 1553 8175 2499
rect 8211 2201 8223 6243
rect 8259 5897 8271 6915
rect 8187 1553 8199 2163
rect 8235 1553 8247 2139
rect 8259 1553 8271 3747
rect 8283 3161 8295 6915
rect 8307 5129 8319 6915
rect 8331 1553 8343 4515
rect 8355 3977 8367 6915
rect 8379 6257 8391 6915
rect 8403 6329 8415 6915
rect 8451 5897 8463 6915
rect 8475 6353 8487 6915
rect 8523 6377 8535 6915
rect 8355 1553 8367 2115
rect 8403 1553 8415 5883
rect 8451 1553 8463 4179
rect 8571 3161 8583 6915
rect 8595 5777 8607 6915
rect 8619 4457 8631 6915
rect 8667 6401 8679 6915
rect 8691 4697 8703 6915
rect 8715 6425 8727 6915
rect 8763 3497 8775 6915
rect 8787 3257 8799 6915
rect 8835 6449 8847 6915
rect 8883 3521 8895 6915
rect 8907 4001 8919 6915
rect 8931 4217 8943 6915
rect 8475 1553 8487 2499
rect 8667 1553 8679 2499
rect 8715 1553 8727 2091
rect 8763 1553 8775 2067
rect 8787 1553 8799 2043
rect 8883 1553 8895 2139
rect 8907 1553 8919 3867
rect 8955 1553 8967 3123
rect 8979 2417 8991 6915
rect 9003 2729 9015 6915
rect 9027 6473 9039 6915
rect 9075 6497 9087 6915
rect 9099 6521 9111 6915
rect 9147 6545 9159 6915
rect 9195 6569 9207 6915
rect 9003 1553 9015 2019
rect 9027 1553 9039 4707
rect 9051 2033 9063 5763
rect 9051 1553 9063 1995
rect 9099 1553 9111 3747
rect 9123 1553 9135 2139
rect 9147 1553 9159 4419
rect 9183 2105 9195 6507
rect 9219 3497 9231 6915
rect 9243 4265 9255 6915
rect 9267 6521 9279 6915
rect 9315 6593 9327 6915
rect 9339 6617 9351 6915
rect 9171 1553 9183 2019
rect 9219 1553 9231 2091
rect 9279 1985 9291 4491
rect 9243 1553 9255 1971
rect 9315 1553 9327 4947
rect 9339 1553 9351 2331
rect 9387 1985 9399 6915
rect 9435 2177 9447 6915
rect 9459 4217 9471 6915
rect 9387 1553 9399 1947
rect 9459 1553 9471 4059
rect 9483 2129 9495 6915
rect 9531 2129 9543 6915
rect 9555 4313 9567 6915
rect 9483 1553 9495 1923
rect 9531 1553 9543 1899
rect 9579 1889 9591 6915
rect 9579 1553 9591 1851
rect 9603 1553 9615 6627
rect 9627 4649 9639 6915
rect 9651 3041 9663 6915
rect 9699 4961 9711 6915
rect 9675 1553 9687 3747
rect 9699 1553 9711 4707
rect 9747 3161 9759 6915
rect 9747 1553 9759 2259
rect 9771 2153 9783 6915
rect 9795 6665 9807 6915
rect 9795 1553 9807 1827
rect 9819 1553 9831 6675
rect 9843 2249 9855 6915
rect 9867 2033 9879 6915
rect 9891 3929 9903 6915
rect 9915 3953 9927 6915
rect 9867 1553 9879 1803
rect 9939 1553 9951 4275
rect 9963 2753 9975 6915
rect 9987 2345 9999 6915
rect 10035 4985 10047 6915
rect 10011 1553 10023 2499
rect 10035 1553 10047 3939
rect 10059 1553 10071 4755
rect 10083 3761 10095 6915
rect 10107 3281 10119 6915
rect 10107 1553 10119 1995
rect 10131 1553 10143 3915
rect 10155 2873 10167 6915
rect 10203 3617 10215 6915
rect 10227 4985 10239 6915
rect 10155 1553 10167 2739
rect 10179 1553 10191 2235
rect 10251 1553 10263 4539
rect 10275 2945 10287 6915
rect 10275 1553 10287 2019
rect 10299 1553 10311 6075
rect 10323 2945 10335 6915
rect 10347 5273 10359 6915
rect 10371 3569 10383 6915
rect 10395 6713 10407 6915
rect 10407 3953 10419 5451
rect 10443 5129 10455 6915
rect 10491 6689 10503 6915
rect 10323 1553 10335 1779
rect 10371 1553 10383 1755
rect 10395 1553 10407 3867
rect 10419 1553 10431 1731
rect 10467 1553 10479 6555
rect 10563 5129 10575 6915
rect 10491 1553 10503 4947
rect 10515 1553 10527 4179
rect 10539 1553 10551 3939
rect 10587 3593 10599 6915
rect 10611 6641 10623 6915
rect 10587 1553 10599 2259
rect 10623 2033 10635 5835
rect 10659 4145 10671 6915
rect 10683 2369 10695 6915
rect 10707 6641 10719 6915
rect 10731 6689 10743 6915
rect 10755 4217 10767 6915
rect 10803 6737 10815 6915
rect 10611 1553 10623 1707
rect 10683 1553 10695 1731
rect 10707 1553 10719 4203
rect 10755 1553 10767 4131
rect 10779 1769 10791 5763
rect 10803 1553 10815 6435
rect 10827 5609 10839 6915
rect 10851 6161 10863 6915
rect 10827 1553 10839 4179
rect 10851 1553 10863 2355
rect 10875 2297 10887 6627
rect 10899 6161 10911 6915
rect 10899 1553 10911 2787
rect 10923 2513 10935 6147
rect 10947 4553 10959 6915
rect 11019 5537 11031 6915
rect 11043 5729 11055 6915
rect 11067 5537 11079 6915
rect 11091 5729 11103 6915
rect 11139 6161 11151 6915
rect 11163 6329 11175 6915
rect 11187 3569 11199 6915
rect 11211 6329 11223 6915
rect 11259 4289 11271 6915
rect 11283 4193 11295 6915
rect 11307 6641 11319 6915
rect 11355 5465 11367 6915
rect 11019 1553 11031 2787
rect 11043 1553 11055 2331
rect 11115 1553 11127 2283
rect 11163 1553 11175 2019
rect 11187 1553 11199 2907
rect 11211 1553 11223 1755
rect 11259 1553 11271 2907
rect 11283 1553 11295 3867
rect 11355 1553 11367 1683
rect 11379 1553 11391 6075
rect 11403 5969 11415 6915
rect 11427 1697 11439 6003
rect 11475 5561 11487 6915
rect 11499 6761 11511 6915
rect 11523 5585 11535 6915
rect 11571 4601 11583 6915
rect 11595 5585 11607 6915
rect 11619 3425 11631 6915
rect 11667 5201 11679 6915
rect 11691 5777 11703 6915
rect 11715 2033 11727 6915
rect 11763 5969 11775 6915
rect 11787 4121 11799 6915
rect 11811 6689 11823 6915
rect 11859 5489 11871 6915
rect 11883 5201 11895 6915
rect 11907 5537 11919 6915
rect 11955 4505 11967 6915
rect 11979 4529 11991 6915
rect 12003 3833 12015 6915
rect 12027 5537 12039 6915
rect 12075 5369 12087 6915
rect 11403 1553 11415 1659
rect 11499 1553 11511 1683
rect 12027 1553 12039 5355
rect 12099 2897 12111 6915
rect 12123 3425 12135 6915
rect 12147 4817 12159 6915
rect 12171 6785 12183 6915
rect 12219 6809 12231 6915
rect 12243 5921 12255 6915
rect 12267 6113 12279 6915
rect 12171 1553 12183 5187
rect 12219 1553 12231 5259
rect 12315 4481 12327 6915
rect 12243 1553 12255 3555
rect 12267 1553 12279 2019
rect 12315 1553 12327 2139
rect 12339 1553 12351 6003
rect 12363 4241 12375 6915
rect 12435 6833 12447 6915
rect 12435 1553 12447 5787
rect 12459 4289 12471 6915
rect 12483 5033 12495 6915
rect 12531 4409 12543 6915
rect 12555 4289 12567 6915
rect 12603 4481 12615 6915
rect 12459 1553 12471 3723
rect 12531 1553 12543 4275
rect 12627 4241 12639 6243
rect 12651 5033 12663 6915
rect 12675 5201 12687 6915
rect 12699 6857 12711 6915
rect 12555 1553 12567 2499
rect 12603 1553 12615 4227
rect 12651 1553 12663 3603
rect 12675 1553 12687 4803
rect 12699 1553 12711 6795
rect 12723 2609 12735 5187
rect 12747 3281 12759 6915
rect 12771 2657 12783 6915
rect 12795 5201 12807 6915
rect 12747 1553 12759 1635
rect 12795 1553 12807 4179
rect 12819 2993 12831 6915
rect 12867 6689 12879 6915
rect 12915 6401 12927 6915
rect 12819 1553 12831 2595
rect 12843 1649 12855 5979
rect 12867 1553 12879 5667
rect 12891 1553 12903 2571
rect 12927 1721 12939 5187
rect 12963 1553 12975 4227
rect 12987 3761 12999 6915
rect 12987 1553 12999 3603
rect 13011 2153 13023 6915
rect 13035 3377 13047 6915
rect 13059 5201 13071 6915
rect 13059 1553 13071 4587
rect 13107 4529 13119 6915
rect 13131 5825 13143 6915
rect 13155 4649 13167 6915
rect 13083 1553 13095 4419
rect 13107 1553 13119 3723
rect 13179 1649 13191 6579
rect 13203 4649 13215 6915
rect 13155 1553 13167 1635
rect 13203 1553 13215 4491
rect 13251 3473 13263 6915
rect 13275 1553 13287 4707
rect 13299 1553 13311 3771
rect 13323 3737 13335 6915
rect 13347 4793 13359 6915
rect 13371 3953 13383 6915
rect 13395 4793 13407 6915
rect 13347 1553 13359 1635
rect 13395 1553 13407 2331
rect 13419 2081 13431 6915
rect 13419 1553 13431 1611
rect 13443 1553 13455 4683
rect 13467 2345 13479 6915
rect 13491 2513 13503 6915
rect 13515 5801 13527 6915
rect 13539 1649 13551 6603
rect 13563 6401 13575 6915
rect 13587 1625 13599 6675
rect 13635 1553 13647 5499
rect 13683 4145 13695 6915
rect 13707 3617 13719 6915
rect 13755 6353 13767 6915
rect 13803 5921 13815 6915
rect 13827 6353 13839 6915
rect 13851 6809 13863 6915
rect 13827 1553 13839 3939
rect 13851 1553 13863 3723
rect 13899 3569 13911 6915
rect 13923 4025 13935 6915
rect 13947 5777 13959 6915
rect 13899 1553 13911 3483
rect 13923 1553 13935 3027
rect 13971 2345 13983 6915
rect 13995 6881 14007 6915
rect 14007 2081 14019 6483
rect 14043 6425 14055 6915
rect 14091 3977 14103 6915
rect 14163 6905 14175 6915
rect 13947 1553 13959 2067
rect 13995 1553 14007 1635
rect 14043 1553 14055 2067
rect 14115 1553 14127 3603
rect 14139 1553 14151 6699
rect 14163 1553 14175 6747
rect 14187 3041 14199 6915
rect 14211 6713 14223 6915
rect 14211 1553 14223 4803
rect 14259 4097 14271 6915
rect 14235 1553 14247 3771
rect 14283 2345 14295 6915
rect 14307 6833 14319 6915
rect 14259 1553 14271 1611
rect 14307 1553 14319 4155
rect 14355 4025 14367 6915
rect 14331 1553 14343 3555
rect 14379 2513 14391 6915
rect 14403 6761 14415 6915
rect 14403 1553 14415 3699
rect 14427 1553 14439 5955
rect 14451 4913 14463 6915
rect 14475 5633 14487 6915
rect 14499 4913 14511 6915
rect 14451 1553 14463 3651
rect 14499 1553 14511 4083
rect 14523 3353 14535 6915
rect 14571 5633 14583 6915
rect 14619 5489 14631 6915
rect 14643 6833 14655 6915
rect 14523 1553 14535 1587
rect 14547 1553 14559 4011
rect 14595 1553 14607 3699
rect 14667 2081 14679 6915
rect 14691 5801 14703 6891
rect 14619 1553 14631 1995
rect 14691 1577 14703 5619
rect 14715 3665 14727 6915
rect 14667 1553 14679 1563
rect 14715 1553 14727 3483
rect 14739 3401 14751 6915
rect 14763 5585 14775 6915
rect 14739 1553 14751 2187
rect 14787 1553 14799 5883
rect 14811 4865 14823 6915
rect 14835 6089 14847 6915
rect 14859 5105 14871 6915
rect 14835 1553 14847 3051
rect 14859 1553 14871 3627
rect 14883 2945 14895 6699
rect 14907 5105 14919 6915
rect 14931 1553 14943 5091
rect 14955 2441 14967 6915
rect 14979 2897 14991 6915
rect 15003 5105 15015 6915
rect 15027 5585 15039 6915
rect 14979 1553 14991 2067
rect 15027 1553 15039 3147
rect 15051 2129 15063 6747
rect 15075 1601 15087 6651
rect 15147 5633 15159 6915
rect 15099 2177 15111 3651
rect 15123 1553 15135 3747
rect 15147 1553 15159 3651
rect 15171 2081 15183 5547
rect 15219 1553 15231 1875
rect 15243 1553 15255 4395
rect 15315 1553 15327 3771
rect 15435 1553 15447 6099
rect 15459 1553 15471 6867
rect 15507 5561 15519 6915
rect 15507 1553 15519 5355
rect 15555 5033 15567 6915
rect 15531 1553 15543 3627
rect 15579 1553 15591 3027
rect 15627 1553 15639 5979
rect 15699 4289 15711 6915
rect 15723 5465 15735 6915
rect 15771 4985 15783 6915
rect 15891 6209 15903 6915
rect 15699 1553 15711 3339
rect 15723 1553 15735 4179
rect 15771 1553 15783 2931
rect 15843 1553 15855 2499
rect 15867 1553 15879 2763
rect 15915 1553 15927 6003
rect 15963 1553 15975 4251
rect 16251 3761 16263 6915
rect 16299 5921 16311 6915
rect 16035 1553 16047 3387
rect 16083 1553 16095 3507
rect 16443 1937 16455 6915
rect 16491 5273 16503 6915
rect 16515 4265 16527 6915
rect 16539 4985 16551 6915
rect 16587 4361 16599 6915
rect 16611 5777 16623 6915
rect 16635 2753 16647 6915
rect 16683 4361 16695 6915
rect 16731 5753 16743 6915
rect 16755 3233 16767 6915
rect 16635 1553 16647 2619
rect 16779 1553 16791 3891
rect 16803 3089 16815 6915
rect 16851 4049 16863 6915
rect 16875 6473 16887 6915
rect 16803 1553 16815 2475
rect 16875 1553 16887 3507
rect 16899 1553 16911 3483
rect 16923 1553 16935 3963
rect 16971 3569 16983 6915
rect 16947 1553 16959 3315
rect 16995 2345 17007 6915
rect 16995 1553 17007 2115
rect 17019 1553 17031 6627
rect 17043 5753 17055 6915
rect 17043 1553 17055 4035
rect 17067 2129 17079 6915
rect 17139 5897 17151 6915
rect 17163 6017 17175 6915
rect 17187 5417 17199 6915
rect 17211 5513 17223 6915
rect 17091 1553 17103 2091
rect 17115 1553 17127 3147
rect 17211 1553 17223 4443
rect 17235 1553 17247 3891
rect 17259 3281 17271 6915
rect 17283 3833 17295 6915
rect 17259 1553 17271 2883
rect 17307 1553 17319 6483
rect 17331 4457 17343 6915
rect 17355 1553 17367 5835
rect 17379 2369 17391 6915
rect 17403 6305 17415 6915
rect 17427 6881 17439 6915
rect 17427 1553 17439 6819
rect 17451 4577 17463 6915
rect 17475 5417 17487 6915
rect 17523 5585 17535 6915
rect 17547 4817 17559 6915
rect 17475 1553 17487 2211
rect 17499 1553 17511 3507
rect 17571 1865 17583 6915
rect 17571 1553 17583 1587
rect 17595 1553 17607 5595
rect 17619 3737 17631 6915
rect 17619 1553 17631 3531
rect 17643 2897 17655 6723
rect 17667 4505 17679 6915
rect 17691 3833 17703 6915
rect 17667 1553 17679 3723
rect 17715 3713 17727 6915
rect 17715 1553 17727 3531
rect 17739 1841 17751 5403
rect 17763 5345 17775 6915
rect 17787 6425 17799 6915
rect 17763 1553 17775 4131
rect 17799 3737 17811 5907
rect 17835 4577 17847 6915
rect 17787 1553 17799 3147
rect 17859 1601 17871 6795
rect 17883 2345 17895 6915
rect 17907 3785 17919 6915
rect 17883 1553 17895 1971
rect 17907 1553 17919 3675
rect 17931 3041 17943 6915
rect 17955 6713 17967 6915
rect 17955 1553 17967 6507
rect 17979 1913 17991 6699
rect 18003 4313 18015 6915
rect 18027 3257 18039 6915
rect 18051 3401 18063 6915
rect 18027 1553 18039 3147
rect 18075 1553 18087 6603
rect 18099 1553 18111 3291
rect 18147 1553 18159 5355
rect 18171 5345 18183 6915
rect 18579 6401 18591 6915
rect 18195 1553 18207 5835
rect 18243 1553 18255 5883
rect 18291 1553 18303 4131
rect 18363 1553 18375 5619
rect 18411 1553 18423 3267
rect 18435 1553 18447 1707
rect 18459 1553 18471 4899
rect 18723 3161 18735 6915
rect 18771 2681 18783 6915
rect 18819 1625 18831 6915
rect 18867 5777 18879 6915
rect 18939 4985 18951 6915
rect 18987 6353 18999 6915
rect 19059 1721 19071 6915
rect 19083 3785 19095 6915
rect 19107 4913 19119 6915
rect 19155 5513 19167 6915
rect 19179 6713 19191 6915
rect 19131 1553 19143 5259
rect 19179 1553 19191 6555
rect 19203 5417 19215 6915
rect 19251 2057 19263 6915
rect 19299 5585 19311 6915
rect 19323 5609 19335 6915
rect 19347 3953 19359 6915
rect 19275 1553 19287 3819
rect 19299 1553 19311 3219
rect 19323 1553 19335 3723
rect 19395 3449 19407 6915
rect 19419 3233 19431 6915
rect 19371 1553 19383 1755
rect 19419 1553 19431 3147
rect 19443 1697 19455 6915
rect 19491 5633 19503 6915
rect 19515 6113 19527 6915
rect 19467 2273 19479 5571
rect 19491 1553 19503 4299
rect 19515 1553 19527 6075
rect 19539 3905 19551 6915
rect 19587 5585 19599 6915
rect 19563 1553 19575 2835
rect 19611 1553 19623 5787
rect 19635 3833 19647 6915
rect 19671 4985 19683 6099
rect 19659 1553 19671 3243
rect 19707 3161 19719 6915
rect 19731 1553 19743 6147
rect 19755 4985 19767 6915
rect 19803 5897 19815 6915
rect 19755 1553 19767 3771
rect 19779 1553 19791 4995
rect 19803 1553 19815 5115
rect 19827 3113 19839 6915
rect 19851 6113 19863 6915
rect 19851 1553 19863 5187
rect 19899 4841 19911 6915
rect 19923 4913 19935 6915
rect 19947 5609 19959 6915
rect 19995 6209 20007 6915
rect 20019 5921 20031 6915
rect 19875 1553 19887 3939
rect 19899 1553 19911 3891
rect 19947 1553 19959 3795
rect 19971 2873 19983 5619
rect 19995 1553 20007 5763
rect 20019 1553 20031 4467
rect 20043 3737 20055 4971
rect 20067 4481 20079 6915
rect 20115 4505 20127 6915
rect 20091 1553 20103 3819
rect 20115 1553 20127 3003
rect 20139 2105 20151 6915
rect 20163 4553 20175 6915
rect 20187 4985 20199 6915
rect 20163 1553 20175 4059
rect 20187 1553 20199 4347
rect 20211 4025 20223 5883
rect 20235 5129 20247 6915
rect 20235 1553 20247 4875
rect 20259 4361 20271 6915
rect 20307 6881 20319 6915
rect 20319 3905 20331 6099
rect 20355 3137 20367 6915
rect 20283 1553 20295 2643
rect 20355 1553 20367 3027
rect 20379 2849 20391 6915
rect 20403 3521 20415 6915
rect 20379 1553 20391 2763
rect 20403 1553 20415 3435
rect 20427 2945 20439 5115
rect 20451 2561 20463 6915
rect 20475 5609 20487 6915
rect 20499 5897 20511 6915
rect 20451 1553 20463 2475
rect 20475 1553 20487 5355
rect 20499 1553 20511 5811
rect 20523 1553 20535 4803
rect 20547 3497 20559 6915
rect 20571 3113 20583 6915
rect 20619 4865 20631 6915
rect 20667 6089 20679 6915
rect 20691 6257 20703 6915
rect 20715 6161 20727 6915
rect 20595 1553 20607 2331
rect 20643 1553 20655 6075
rect 20763 4553 20775 6915
rect 20715 1553 20727 3987
rect 20739 1553 20751 4491
rect 20811 3425 20823 6915
rect 20763 1553 20775 2715
rect 20787 1553 20799 2811
rect 20835 1553 20847 4827
rect 20859 3041 20871 5859
rect 20883 5057 20895 6915
rect 20907 4313 20919 6915
rect 20931 4505 20943 6915
rect 20979 6233 20991 6915
rect 20955 1553 20967 4515
rect 21003 3065 21015 6915
rect 21027 4841 21039 6915
rect 21051 5825 21063 6915
rect 21027 1553 21039 4395
rect 21051 1553 21063 5667
rect 21075 2777 21087 5979
rect 21099 1553 21111 5427
rect 21123 3785 21135 6915
rect 21147 5273 21159 6915
rect 21195 6209 21207 6915
rect 21123 1553 21135 3723
rect 21207 2609 21219 5595
rect 21243 4865 21255 6915
rect 21171 1553 21183 2043
rect 21243 1553 21255 3987
rect 21267 3761 21279 6915
rect 21291 6593 21303 6915
rect 21303 2801 21315 5883
rect 21339 4961 21351 6915
rect 21363 6329 21375 6915
rect 21339 1553 21351 4251
rect 21363 1553 21375 2499
rect 21387 1553 21399 5307
rect 21411 4361 21423 6915
rect 21459 4529 21471 6915
rect 21435 1553 21447 4203
rect 21459 1553 21471 4011
rect 21483 3761 21495 6915
rect 21531 6281 21543 6915
rect 21507 4985 21519 5811
rect 21507 2465 21519 4539
rect 21555 1553 21567 3747
rect 21579 1985 21591 6915
rect 21603 2321 21615 6915
rect 21627 3089 21639 4827
rect 21651 3929 21663 6915
rect 21651 1553 21663 3891
rect 21675 3737 21687 4635
rect 21699 4625 21711 6915
rect 21723 2393 21735 6915
rect 21747 6377 21759 6915
rect 21771 6593 21783 6915
rect 21699 1553 21711 2139
rect 21771 1553 21783 6555
rect 21795 5585 21807 6915
rect 21795 1553 21807 3483
rect 21819 1553 21831 3555
rect 21843 1745 21855 6915
rect 21867 3593 21879 4851
rect 21891 4529 21903 6915
rect 21843 1553 21855 1683
rect 21891 1553 21903 3339
rect 21915 1553 21927 5523
rect 21939 4025 21951 5427
rect 21963 3665 21975 6915
rect 21987 3593 21999 6915
rect 22011 5249 22023 6915
rect 22011 1553 22023 4203
rect 22035 1553 22047 4443
rect 22059 4385 22071 6915
rect 22083 3905 22095 4899
rect 22107 3113 22119 6915
rect 22131 1553 22143 6627
rect 22155 4793 22167 6579
rect 22179 1553 22191 5859
rect 22203 1697 22215 6003
rect 22227 4217 22239 6603
rect 22251 5729 22263 6915
rect 22611 6041 22623 6915
rect 22659 5705 22671 6915
rect 22251 1553 22263 4011
rect 22371 1553 22383 2163
rect 22419 1553 22431 2187
rect 22515 1553 22527 4491
rect 22539 1553 22551 4203
rect 22587 1553 22599 4275
rect 22707 1553 22719 3123
rect 22731 1553 22743 3363
rect 22779 1553 22791 2091
rect 22803 2009 22815 6915
rect 22851 4241 22863 6915
rect 22851 1553 22863 2331
rect 22875 1553 22887 5259
rect 22923 4241 22935 6915
rect 22947 5465 22959 6915
rect 22995 4673 23007 6915
rect 23019 4001 23031 6123
rect 22995 1553 23007 3987
rect 23043 3761 23055 6915
rect 23067 4745 23079 6915
rect 23091 3785 23103 6915
rect 23115 3953 23127 6915
rect 23163 4073 23175 6915
rect 23163 1553 23175 3987
rect 23187 1553 23199 4251
rect 23211 1553 23223 4395
rect 23235 4001 23247 6075
rect 23283 5969 23295 6915
rect 23307 5153 23319 6915
rect 23259 1553 23271 1995
rect 23307 1553 23319 4923
rect 23331 4649 23343 6915
rect 23379 4049 23391 6915
rect 23403 3785 23415 6915
rect 23355 1553 23367 3123
rect 23379 1553 23391 3747
rect 23427 1553 23439 4587
rect 23451 4289 23463 6915
rect 23475 1553 23487 6675
rect 23499 4745 23511 6915
rect 23499 1553 23511 4683
rect 23523 3401 23535 6915
rect 23619 4769 23631 6915
rect 23547 4097 23559 4731
rect 23595 1553 23607 3747
rect 23619 1553 23631 4059
rect 23643 1553 23655 5091
rect 23667 2729 23679 6915
rect 23691 4073 23703 5307
rect 23739 4361 23751 6915
rect 23763 6641 23775 6915
rect 23811 4025 23823 6915
rect 23859 6665 23871 6915
rect 23811 1553 23823 3099
rect 23835 1553 23847 5955
rect 23883 1553 23895 6051
rect 23907 4457 23919 6915
rect 23979 5777 23991 6915
rect 23931 1553 23943 5667
rect 23955 1553 23967 5019
rect 24003 3545 24015 6915
rect 24027 3617 24039 6915
rect 24051 3857 24063 6915
rect 24099 5849 24111 6915
rect 24123 5801 24135 6915
rect 24027 1553 24039 3555
rect 24051 1553 24063 3795
rect 24075 3569 24087 4563
rect 24147 4505 24159 6915
rect 24099 1553 24111 3171
rect 24147 1553 24159 3483
rect 24171 1553 24183 6555
rect 24195 5513 24207 6915
rect 24219 4529 24231 6915
rect 24243 4553 24255 6915
rect 24291 5921 24303 6915
rect 24195 1553 24207 4059
rect 24255 3353 24267 4491
rect 24315 4217 24327 6915
rect 24339 4337 24351 6915
rect 24387 6881 24399 6915
rect 24243 1553 24255 2979
rect 24291 1553 24303 3315
rect 24315 1553 24327 3219
rect 24339 1553 24351 4035
rect 24363 1649 24375 4539
rect 24387 1553 24399 6843
rect 24411 4433 24423 6915
rect 24435 5177 24447 6915
rect 24411 1553 24423 4011
rect 24435 1553 24447 4107
rect 24459 1553 24471 4227
rect 24483 3497 24495 6915
rect 24507 2033 24519 6915
rect 24531 3833 24543 6915
rect 24579 5417 24591 6915
rect 24603 4241 24615 6915
rect 24627 4337 24639 6915
rect 24651 5345 24663 6915
rect 24675 4457 24687 6867
rect 24507 1553 24519 1779
rect 24555 1553 24567 4155
rect 24627 1553 24639 2259
rect 24699 1673 24711 6915
rect 24723 3449 24735 6915
rect 24747 5393 24759 6915
rect 24651 1553 24663 1611
rect 24723 1553 24735 2859
rect 24747 1553 24759 4203
rect 24795 4049 24807 6915
rect 24843 5297 24855 6915
rect 24867 4193 24879 6915
rect 24891 4433 24903 6915
rect 24819 1553 24831 2643
rect 24843 1553 24855 1707
rect 24915 1553 24927 5475
rect 24939 4073 24951 6915
rect 24963 1793 24975 6915
rect 24987 1817 24999 6915
rect 25011 3233 25023 6915
rect 25083 6617 25095 6915
rect 25107 5921 25119 6915
rect 25131 6185 25143 6915
rect 25035 1553 25047 4275
rect 25179 2705 25191 6915
rect 25203 4769 25215 6915
rect 25251 3809 25263 6915
rect 25299 6281 25311 6915
rect 25323 3977 25335 6915
rect 25347 4097 25359 6915
rect 25395 3281 25407 6915
rect 25419 2273 25431 6915
rect 25443 1721 25455 6915
rect 25467 4793 25479 6915
rect 25515 3593 25527 6915
rect 25539 4817 25551 6915
rect 25563 4745 25575 6915
rect 25611 5489 25623 6915
rect 25563 1553 25575 4707
rect 25587 2249 25599 4731
rect 25611 1553 25623 3867
rect 25635 2297 25647 6915
rect 25659 4337 25671 6915
rect 25707 3473 25719 6915
rect 25731 6449 25743 6915
rect 25755 4265 25767 6915
rect 25755 1553 25767 4203
rect 25779 2537 25791 6915
rect 25803 4217 25815 5835
rect 25827 5513 25839 6915
rect 25851 4265 25863 6915
rect 25875 6881 25887 6915
rect 25779 1553 25791 2451
rect 25851 1553 25863 4011
rect 25875 1553 25887 6843
rect 25899 4145 25911 6867
rect 25923 4313 25935 6915
rect 25947 2513 25959 6915
rect 25971 4385 25983 6915
rect 26019 5081 26031 6915
rect 26043 6569 26055 6915
rect 26091 5753 26103 6915
rect 26139 3785 26151 6915
rect 26163 5225 26175 6915
rect 26187 2489 26199 6915
rect 26235 6281 26247 6915
rect 26259 2849 26271 6915
rect 26307 2417 26319 6915
rect 26355 2585 26367 6915
rect 26379 5561 26391 6915
rect 26403 4025 26415 6915
rect 26379 1553 26391 1707
rect 26427 1553 26439 4803
rect 26451 2657 26463 6915
rect 26475 4817 26487 6915
rect 26499 5657 26511 6915
rect 26547 1961 26559 6915
rect 26571 6545 26583 6915
rect 26571 1553 26583 6387
rect 26619 4505 26631 6915
rect 26667 5681 26679 6915
rect 26691 6401 26703 6915
rect 26619 1553 26631 4467
rect 26643 4361 26655 4491
rect 26715 4241 26727 6915
rect 26739 1553 26751 6699
rect 26763 4433 26775 6915
rect 26787 3209 26799 6915
rect 26787 1553 26799 3171
rect 26811 2465 26823 6915
rect 26859 6353 26871 6915
rect 26883 5945 26895 6915
rect 26907 5009 26919 6915
rect 26835 3185 26847 4515
rect 26931 2921 26943 6915
rect 26979 4409 26991 6915
rect 27027 3377 27039 6915
rect 27099 1769 27111 6915
rect 27123 1577 27135 4251
rect 27147 1601 27159 3627
rect 27243 1553 27443 6915
rect 27507 6772 27577 6784
rect 27507 2956 27577 2968
rect 27507 1588 27577 1600
rect 27507 1564 27577 1576
rect 0 83 70 95
rect 0 59 70 71
rect 123 0 323 754
rect 339 0 351 754
rect 363 0 375 754
rect 387 0 399 754
rect 411 0 423 754
rect 1731 96 1743 754
rect 1851 96 1863 754
rect 2691 120 2703 754
rect 2715 144 2727 754
rect 2835 168 2847 754
rect 3507 192 3519 754
rect 3675 144 3687 754
rect 3747 144 3759 754
rect 4131 216 4143 754
rect 4491 240 4503 754
rect 4611 168 4623 754
rect 4707 168 4719 754
rect 4755 264 4767 754
rect 4779 96 4791 754
rect 5043 96 5055 754
rect 5091 288 5103 754
rect 5283 312 5295 754
rect 5427 336 5439 754
rect 5979 48 5991 754
rect 6051 360 6063 754
rect 6219 384 6231 754
rect 6339 120 6351 754
rect 6387 216 6399 754
rect 6411 120 6423 754
rect 6435 216 6447 754
rect 6747 408 6759 754
rect 7083 432 7095 754
rect 7371 456 7383 754
rect 7635 120 7647 754
rect 7683 312 7695 754
rect 7803 312 7815 754
rect 7995 480 8007 754
rect 8043 504 8055 754
rect 8283 264 8295 754
rect 8571 360 8583 754
rect 8643 264 8655 754
rect 8835 144 8847 754
rect 9267 144 9279 754
rect 9435 528 9447 754
rect 9555 552 9567 754
rect 9627 576 9639 754
rect 9915 360 9927 754
rect 9963 360 9975 754
rect 10203 600 10215 754
rect 10635 168 10647 754
rect 10923 168 10935 754
rect 10971 624 10983 754
rect 11067 168 11079 754
rect 11115 168 11127 754
rect 11307 168 11319 754
rect 11451 648 11463 754
rect 11128 154 11146 168
rect 7947 0 7959 106
rect 11127 0 11139 154
rect 12171 120 12183 754
rect 12387 120 12399 754
rect 12483 672 12495 754
rect 12771 192 12783 754
rect 12915 696 12927 754
rect 13011 720 13023 754
rect 13467 96 13479 754
rect 13515 96 13527 754
rect 13539 120 13551 754
rect 13587 552 13599 754
rect 13683 552 13695 754
rect 13755 672 13767 754
rect 13779 384 13791 754
rect 13803 552 13815 754
rect 14019 696 14031 754
rect 14067 336 14079 754
rect 14355 384 14367 754
rect 14883 552 14895 754
rect 14907 480 14919 754
rect 15099 480 15111 754
rect 15195 408 15207 754
rect 15267 672 15279 754
rect 15339 288 15351 754
rect 15387 696 15399 754
rect 15483 336 15495 754
rect 15819 192 15831 754
rect 16227 288 16239 754
rect 16827 120 16839 754
rect 17163 744 17175 754
rect 17427 24 17439 754
rect 17523 504 17535 754
rect 17691 672 17703 754
rect 17811 504 17823 754
rect 17859 168 17871 754
rect 17979 384 17991 754
rect 18003 672 18015 754
rect 18219 360 18231 754
rect 18315 384 18327 754
rect 18339 360 18351 754
rect 18579 168 18591 754
rect 18987 288 18999 754
rect 19251 144 19263 754
rect 19923 288 19935 754
rect 20043 144 20055 754
rect 20139 24 20151 754
rect 20547 648 20559 754
rect 20883 312 20895 754
rect 20979 648 20991 754
rect 21003 624 21015 754
rect 21219 624 21231 754
rect 21291 456 21303 754
rect 21483 528 21495 754
rect 21531 312 21543 754
rect 21603 96 21615 754
rect 21963 24 21975 754
rect 22083 480 22095 754
rect 22275 744 22287 754
rect 22323 552 22335 754
rect 22491 408 22503 754
rect 22635 192 22647 754
rect 22827 192 22839 754
rect 22923 720 22935 754
rect 22947 408 22959 754
rect 23043 72 23055 754
rect 23091 168 23103 754
rect 23283 144 23295 754
rect 23547 264 23559 754
rect 23691 432 23703 754
rect 23739 648 23751 754
rect 23979 384 23991 754
rect 24267 504 24279 754
rect 24675 288 24687 754
rect 24771 408 24783 754
rect 24867 240 24879 754
rect 24939 384 24951 754
rect 24963 408 24975 754
rect 25011 576 25023 754
rect 24952 370 24970 384
rect 17440 10 17458 24
rect 17439 0 17451 10
rect 24951 0 24963 370
rect 24987 360 24999 394
rect 25083 336 25095 754
rect 25203 120 25215 754
rect 25803 672 25815 754
rect 25899 624 25911 754
rect 26019 600 26031 754
rect 26571 384 26583 754
rect 26643 696 26655 754
rect 26691 216 26703 754
rect 26739 408 26751 754
rect 26787 432 26799 754
rect 26787 24 26799 370
rect 27243 0 27443 754
rect 27507 419 27577 431
rect 27507 395 27577 407
rect 27507 35 27577 47
rect 27507 11 27577 23
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 6915
box 0 0 1464 799
use nand2 g8197
timestamp 1386234792
transform 1 0 1587 0 1 6915
box 0 0 96 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 1683 0 1 6915
box 0 0 48 799
use rowcrosser PcEn
timestamp 1386086759
transform 1 0 1731 0 1 6915
box 0 0 48 799
use nor2 g8032
timestamp 1386235306
transform 1 0 1779 0 1 6915
box 0 0 120 799
use nand3 g8316
timestamp 1386234893
transform 1 0 1899 0 1 6915
box 0 0 120 799
use nor2 g8043
timestamp 1386235306
transform 1 0 2019 0 1 6915
box 0 0 120 799
use nand2 g8112
timestamp 1386234792
transform 1 0 2139 0 1 6915
box 0 0 96 799
use nand2 g8291
timestamp 1386234792
transform 1 0 2235 0 1 6915
box 0 0 96 799
use and2 g8060
timestamp 1386234845
transform 1 0 2331 0 1 6915
box 0 0 120 799
use nand2 g8182
timestamp 1386234792
transform 1 0 2451 0 1 6915
box 0 0 96 799
use nand2 g8066
timestamp 1386234792
transform 1 0 2547 0 1 6915
box 0 0 96 799
use nand4 g8169
timestamp 1386234936
transform 1 0 2643 0 1 6915
box 0 0 144 799
use nand2 g8229
timestamp 1386234792
transform 1 0 2787 0 1 6915
box 0 0 96 799
use inv g8107
timestamp 1386238110
transform 1 0 2883 0 1 6915
box 0 0 120 799
use nor2 g8313
timestamp 1386235306
transform 1 0 3003 0 1 6915
box 0 0 120 799
use and2 g8039
timestamp 1386234845
transform 1 0 3123 0 1 6915
box 0 0 120 799
use nand4 g8344
timestamp 1386234936
transform 1 0 3243 0 1 6915
box 0 0 144 799
use nand2 g8123
timestamp 1386234792
transform 1 0 3387 0 1 6915
box 0 0 96 799
use nand2 g8046
timestamp 1386234792
transform 1 0 3483 0 1 6915
box 0 0 96 799
use inv g8222
timestamp 1386238110
transform 1 0 3579 0 1 6915
box 0 0 120 799
use nand2 g8102
timestamp 1386234792
transform 1 0 3699 0 1 6915
box 0 0 96 799
use nand3 g8098
timestamp 1386234893
transform 1 0 3795 0 1 6915
box 0 0 120 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 3915 0 1 6915
box 0 0 48 799
use nand2 g8327
timestamp 1386234792
transform 1 0 3963 0 1 6915
box 0 0 96 799
use inv g8314
timestamp 1386238110
transform 1 0 4059 0 1 6915
box 0 0 120 799
use and2 g8012
timestamp 1386234845
transform 1 0 4179 0 1 6915
box 0 0 120 799
use nand3 g8187
timestamp 1386234893
transform 1 0 4299 0 1 6915
box 0 0 120 799
use nand2 g8135
timestamp 1386234792
transform 1 0 4419 0 1 6915
box 0 0 96 799
use and2 g8171
timestamp 1386234845
transform 1 0 4515 0 1 6915
box 0 0 120 799
use nand2 g8295
timestamp 1386234792
transform 1 0 4635 0 1 6915
box 0 0 96 799
use nand2 g8287
timestamp 1386234792
transform 1 0 4731 0 1 6915
box 0 0 96 799
use inv g8154
timestamp 1386238110
transform 1 0 4827 0 1 6915
box 0 0 120 799
use nand2 g8276
timestamp 1386234792
transform 1 0 4947 0 1 6915
box 0 0 96 799
use nand2 g8261
timestamp 1386234792
transform 1 0 5043 0 1 6915
box 0 0 96 799
use nand2 g8130
timestamp 1386234792
transform 1 0 5139 0 1 6915
box 0 0 96 799
use inv g8082
timestamp 1386238110
transform 1 0 5235 0 1 6915
box 0 0 120 799
use and2 g8027
timestamp 1386234845
transform 1 0 5355 0 1 6915
box 0 0 120 799
use nand2 g8318
timestamp 1386234792
transform 1 0 5475 0 1 6915
box 0 0 96 799
use nand2 g8035
timestamp 1386234792
transform 1 0 5571 0 1 6915
box 0 0 96 799
use nand4 g8019
timestamp 1386234936
transform 1 0 5667 0 1 6915
box 0 0 144 799
use inv g8168
timestamp 1386238110
transform 1 0 5811 0 1 6915
box 0 0 120 799
use nor2 g8238
timestamp 1386235306
transform 1 0 5931 0 1 6915
box 0 0 120 799
use and2 g7989
timestamp 1386234845
transform 1 0 6051 0 1 6915
box 0 0 120 799
use nand2 g8225
timestamp 1386234792
transform 1 0 6171 0 1 6915
box 0 0 96 799
use nand2 g8143
timestamp 1386234792
transform 1 0 6267 0 1 6915
box 0 0 96 799
use nand2 g8333
timestamp 1386234792
transform 1 0 6363 0 1 6915
box 0 0 96 799
use nor2 g2
timestamp 1386235306
transform 1 0 6459 0 1 6915
box 0 0 120 799
use nand3 g8069
timestamp 1386234893
transform 1 0 6579 0 1 6915
box 0 0 120 799
use nand2 g8042
timestamp 1386234792
transform 1 0 6699 0 1 6915
box 0 0 96 799
use nand2 g8149
timestamp 1386234792
transform 1 0 6795 0 1 6915
box 0 0 96 799
use nand3 g8338
timestamp 1386234893
transform 1 0 6891 0 1 6915
box 0 0 120 799
use nand2 g8280
timestamp 1386234792
transform 1 0 7011 0 1 6915
box 0 0 96 799
use inv g8249
timestamp 1386238110
transform 1 0 7107 0 1 6915
box 0 0 120 799
use and2 g8064
timestamp 1386234845
transform 1 0 7227 0 1 6915
box 0 0 120 799
use nand3 g8310
timestamp 1386234893
transform 1 0 7347 0 1 6915
box 0 0 120 799
use nand2 g8235
timestamp 1386234792
transform 1 0 7467 0 1 6915
box 0 0 96 799
use nand3 g8058
timestamp 1386234893
transform 1 0 7563 0 1 6915
box 0 0 120 799
use nand4 g8009
timestamp 1386234936
transform 1 0 7683 0 1 6915
box 0 0 144 799
use nand4 g8362
timestamp 1386234936
transform 1 0 7827 0 1 6915
box 0 0 144 799
use inv g8088
timestamp 1386238110
transform 1 0 7971 0 1 6915
box 0 0 120 799
use nand4 g8055
timestamp 1386234936
transform 1 0 8091 0 1 6915
box 0 0 144 799
use nand2 g8214
timestamp 1386234792
transform 1 0 8235 0 1 6915
box 0 0 96 799
use nand2 g8056
timestamp 1386234792
transform 1 0 8331 0 1 6915
box 0 0 96 799
use nor2 g8281
timestamp 1386235306
transform 1 0 8427 0 1 6915
box 0 0 120 799
use nand2 g8269
timestamp 1386234792
transform 1 0 8547 0 1 6915
box 0 0 96 799
use nand2 g8183
timestamp 1386234792
transform 1 0 8643 0 1 6915
box 0 0 96 799
use and2 g8170
timestamp 1386234845
transform 1 0 8739 0 1 6915
box 0 0 120 799
use nand2 g8124
timestamp 1386234792
transform 1 0 8859 0 1 6915
box 0 0 96 799
use nand2 g8106
timestamp 1386234792
transform 1 0 8955 0 1 6915
box 0 0 96 799
use nor2 g8119
timestamp 1386235306
transform 1 0 9051 0 1 6915
box 0 0 120 799
use nand3 g8275
timestamp 1386234893
transform 1 0 9171 0 1 6915
box 0 0 120 799
use nor2 g8146
timestamp 1386235306
transform 1 0 9291 0 1 6915
box 0 0 120 799
use nand2 g8127
timestamp 1386234792
transform 1 0 9411 0 1 6915
box 0 0 96 799
use nand2 g8155
timestamp 1386234792
transform 1 0 9507 0 1 6915
box 0 0 96 799
use nor2 g8290
timestamp 1386235306
transform 1 0 9603 0 1 6915
box 0 0 120 799
use nand2 g8033
timestamp 1386234792
transform 1 0 9723 0 1 6915
box 0 0 96 799
use nand3 g8252
timestamp 1386234893
transform 1 0 9819 0 1 6915
box 0 0 120 799
use nor2 g8334
timestamp 1386235306
transform 1 0 9939 0 1 6915
box 0 0 120 799
use nor2 g8244
timestamp 1386235306
transform 1 0 10059 0 1 6915
box 0 0 120 799
use nor2 g8240
timestamp 1386235306
transform 1 0 10179 0 1 6915
box 0 0 120 799
use nand3 g8054
timestamp 1386234893
transform 1 0 10299 0 1 6915
box 0 0 120 799
use inv g8139
timestamp 1386238110
transform 1 0 10419 0 1 6915
box 0 0 120 799
use nand2 g8023
timestamp 1386234792
transform 1 0 10539 0 1 6915
box 0 0 96 799
use nand4 g8118
timestamp 1386234936
transform 1 0 10635 0 1 6915
box 0 0 144 799
use nand2 g8363
timestamp 1386234792
transform 1 0 10779 0 1 6915
box 0 0 96 799
use inv g7981
timestamp 1386238110
transform 1 0 10875 0 1 6915
box 0 0 120 799
use nand3 g8111
timestamp 1386234893
transform 1 0 10995 0 1 6915
box 0 0 120 799
use nand3 g8347
timestamp 1386234893
transform 1 0 11115 0 1 6915
box 0 0 120 799
use nand2 g8357
timestamp 1386234792
transform 1 0 11235 0 1 6915
box 0 0 96 799
use inv g8120
timestamp 1386238110
transform 1 0 11331 0 1 6915
box 0 0 120 799
use nand2 g8091
timestamp 1386234792
transform 1 0 11451 0 1 6915
box 0 0 96 799
use nand2 g8134
timestamp 1386234792
transform 1 0 11547 0 1 6915
box 0 0 96 799
use nand2 g8320
timestamp 1386234792
transform 1 0 11643 0 1 6915
box 0 0 96 799
use nand2 g8050
timestamp 1386234792
transform 1 0 11739 0 1 6915
box 0 0 96 799
use nand2 g8218
timestamp 1386234792
transform 1 0 11835 0 1 6915
box 0 0 96 799
use nand3 g7995
timestamp 1386234893
transform 1 0 11931 0 1 6915
box 0 0 120 799
use nand4 g8284
timestamp 1386234936
transform 1 0 12051 0 1 6915
box 0 0 144 799
use nand2 g8198
timestamp 1386234792
transform 1 0 12195 0 1 6915
box 0 0 96 799
use inv g8272
timestamp 1386238110
transform 1 0 12291 0 1 6915
box 0 0 120 799
use nand2 g8199
timestamp 1386234792
transform 1 0 12411 0 1 6915
box 0 0 96 799
use nor2 g8306
timestamp 1386235306
transform 1 0 12507 0 1 6915
box 0 0 120 799
use nand2 g8221
timestamp 1386234792
transform 1 0 12627 0 1 6915
box 0 0 96 799
use nand3 g8319
timestamp 1386234893
transform 1 0 12723 0 1 6915
box 0 0 120 799
use inv g8220
timestamp 1386238110
transform 1 0 12843 0 1 6915
box 0 0 120 799
use nand3 g8230
timestamp 1386234893
transform 1 0 12963 0 1 6915
box 0 0 120 799
use nand2 g8194
timestamp 1386234792
transform 1 0 13083 0 1 6915
box 0 0 96 799
use inv g8004
timestamp 1386238110
transform 1 0 13179 0 1 6915
box 0 0 120 799
use nand4 g8340
timestamp 1386234936
transform 1 0 13299 0 1 6915
box 0 0 144 799
use nand2 rm_assigns_buf_StatusReg_1
timestamp 1386234792
transform 1 0 13443 0 1 6915
box 0 0 96 799
use buffer g8074
timestamp 1386236986
transform 1 0 13539 0 1 6915
box 0 0 120 799
use and2 g8209
timestamp 1386234845
transform 1 0 13659 0 1 6915
box 0 0 120 799
use nand2 g8103
timestamp 1386234792
transform 1 0 13779 0 1 6915
box 0 0 96 799
use nand4 g8268
timestamp 1386234936
transform 1 0 13875 0 1 6915
box 0 0 144 799
use inv g8283
timestamp 1386238110
transform 1 0 14019 0 1 6915
box 0 0 120 799
use nand2 g8321
timestamp 1386234792
transform 1 0 14139 0 1 6915
box 0 0 96 799
use nand2 g8180
timestamp 1386234792
transform 1 0 14235 0 1 6915
box 0 0 96 799
use nand2 g8005
timestamp 1386234792
transform 1 0 14331 0 1 6915
box 0 0 96 799
use nand3 g8052
timestamp 1386234893
transform 1 0 14427 0 1 6915
box 0 0 120 799
use rowcrosser PcWe
timestamp 1386086759
transform 1 0 14547 0 1 6915
box 0 0 48 799
use nand2 g8136
timestamp 1386234792
transform 1 0 14595 0 1 6915
box 0 0 96 799
use nand2 g8110
timestamp 1386234792
transform 1 0 14691 0 1 6915
box 0 0 96 799
use nand2 g8153
timestamp 1386234792
transform 1 0 14787 0 1 6915
box 0 0 96 799
use rowcrosser ALE
timestamp 1386086759
transform 1 0 14883 0 1 6915
box 0 0 48 799
use nand3 StatusReg_reg_91_3_93_
timestamp 1386234893
transform 1 0 14931 0 1 6915
box 0 0 120 799
use scandtype g8308
timestamp 1386241841
transform 1 0 15051 0 1 6915
box 0 0 624 799
use nor2 stateSub_reg_91_2_93_
timestamp 1386235306
transform 1 0 15675 0 1 6915
box 0 0 120 799
use scandtype g8294
timestamp 1386241841
transform 1 0 15795 0 1 6915
box 0 0 624 799
use rowcrosser Op2Sel_91_1_93_
timestamp 1386086759
transform 1 0 16419 0 1 6915
box 0 0 48 799
use nand2 g8024
timestamp 1386234792
transform 1 0 16467 0 1 6915
box 0 0 96 799
use nand2 g8099
timestamp 1386234792
transform 1 0 16563 0 1 6915
box 0 0 96 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 16659 0 1 6915
box 0 0 48 799
use and2 g8057
timestamp 1386234845
transform 1 0 16707 0 1 6915
box 0 0 120 799
use nand2 g8190
timestamp 1386234792
transform 1 0 16827 0 1 6915
box 0 0 96 799
use mux2 g8045
timestamp 1386235218
transform 1 0 16923 0 1 6915
box 0 0 192 799
use nand3 g8304
timestamp 1386234893
transform 1 0 17115 0 1 6915
box 0 0 120 799
use nor2 g8018
timestamp 1386235306
transform 1 0 17235 0 1 6915
box 0 0 120 799
use nand4 g8092
timestamp 1386234936
transform 1 0 17355 0 1 6915
box 0 0 144 799
use nand2 g8277
timestamp 1386234792
transform 1 0 17499 0 1 6915
box 0 0 96 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 17595 0 1 6915
box 0 0 48 799
use nand2 g8081
timestamp 1386234792
transform 1 0 17643 0 1 6915
box 0 0 96 799
use nor2 g8296
timestamp 1386235306
transform 1 0 17739 0 1 6915
box 0 0 120 799
use nand3 g8234
timestamp 1386234893
transform 1 0 17859 0 1 6915
box 0 0 120 799
use nand2 StatusReg_reg_91_1_93_
timestamp 1386234792
transform 1 0 17979 0 1 6915
box 0 0 96 799
use scandtype g8324
timestamp 1386241841
transform 1 0 18075 0 1 6915
box 0 0 624 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 18699 0 1 6915
box 0 0 48 799
use rowcrosser Op1Sel
timestamp 1386086759
transform 1 0 18747 0 1 6915
box 0 0 48 799
use inv g8293
timestamp 1386238110
transform 1 0 18795 0 1 6915
box 0 0 120 799
use inv g8312
timestamp 1386238110
transform 1 0 18915 0 1 6915
box 0 0 120 799
use nand2 g8028
timestamp 1386234792
transform 1 0 19035 0 1 6915
box 0 0 96 799
use nand2 g8213
timestamp 1386234792
transform 1 0 19131 0 1 6915
box 0 0 96 799
use rowcrosser MemEn
timestamp 1386086759
transform 1 0 19227 0 1 6915
box 0 0 48 799
use nand2 g8096
timestamp 1386234792
transform 1 0 19275 0 1 6915
box 0 0 96 799
use nand2 g8212
timestamp 1386234792
transform 1 0 19371 0 1 6915
box 0 0 96 799
use nand2 g8015
timestamp 1386234792
transform 1 0 19467 0 1 6915
box 0 0 96 799
use inv g8084
timestamp 1386238110
transform 1 0 19563 0 1 6915
box 0 0 120 799
use rowcrosser AluEn
timestamp 1386086759
transform 1 0 19683 0 1 6915
box 0 0 48 799
use rowcrosser g8048
timestamp 1386086759
transform 1 0 19731 0 1 6915
box 0 0 48 799
use nand2 g8265
timestamp 1386234792
transform 1 0 19779 0 1 6915
box 0 0 96 799
use nand2 g8200
timestamp 1386234792
transform 1 0 19875 0 1 6915
box 0 0 96 799
use nor2 g8108
timestamp 1386235306
transform 1 0 19971 0 1 6915
box 0 0 120 799
use nand3 g8049
timestamp 1386234893
transform 1 0 20091 0 1 6915
box 0 0 120 799
use nor2 g8159
timestamp 1386235306
transform 1 0 20211 0 1 6915
box 0 0 120 799
use nand2 g8144
timestamp 1386234792
transform 1 0 20331 0 1 6915
box 0 0 96 799
use nand2 g8177
timestamp 1386234792
transform 1 0 20427 0 1 6915
box 0 0 96 799
use and2 g8251
timestamp 1386234845
transform 1 0 20523 0 1 6915
box 0 0 120 799
use nand2 g8036
timestamp 1386234792
transform 1 0 20643 0 1 6915
box 0 0 96 799
use inv g8226
timestamp 1386238110
transform 1 0 20739 0 1 6915
box 0 0 120 799
use nand2 g7979
timestamp 1386234792
transform 1 0 20859 0 1 6915
box 0 0 96 799
use nand4 g8264
timestamp 1386234936
transform 1 0 20955 0 1 6915
box 0 0 144 799
use and2 g8332
timestamp 1386234845
transform 1 0 21099 0 1 6915
box 0 0 120 799
use nand2 g8089
timestamp 1386234792
transform 1 0 21219 0 1 6915
box 0 0 96 799
use and2 g8206
timestamp 1386234845
transform 1 0 21315 0 1 6915
box 0 0 120 799
use and2 g8237
timestamp 1386234845
transform 1 0 21435 0 1 6915
box 0 0 120 799
use nor2 g8016
timestamp 1386235306
transform 1 0 21555 0 1 6915
box 0 0 120 799
use nand4 g8278
timestamp 1386234936
transform 1 0 21675 0 1 6915
box 0 0 144 799
use inv g8181
timestamp 1386238110
transform 1 0 21819 0 1 6915
box 0 0 120 799
use nand2 g8216
timestamp 1386234792
transform 1 0 21939 0 1 6915
box 0 0 96 799
use inv StatusReg_reg_91_0_93_
timestamp 1386238110
transform 1 0 22035 0 1 6915
box 0 0 120 799
use scandtype g8253
timestamp 1386241841
transform 1 0 22155 0 1 6915
box 0 0 624 799
use inv g8186
timestamp 1386238110
transform 1 0 22779 0 1 6915
box 0 0 120 799
use and2 g8090
timestamp 1386234845
transform 1 0 22899 0 1 6915
box 0 0 120 799
use nand3 g8223
timestamp 1386234893
transform 1 0 23019 0 1 6915
box 0 0 120 799
use inv g8195
timestamp 1386238110
transform 1 0 23139 0 1 6915
box 0 0 120 799
use nand2 g8077
timestamp 1386234792
transform 1 0 23259 0 1 6915
box 0 0 96 799
use and2 g8133
timestamp 1386234845
transform 1 0 23355 0 1 6915
box 0 0 120 799
use nor2 g8341
timestamp 1386235306
transform 1 0 23475 0 1 6915
box 0 0 120 799
use inv g8041
timestamp 1386238110
transform 1 0 23595 0 1 6915
box 0 0 120 799
use nor2 g8289
timestamp 1386235306
transform 1 0 23715 0 1 6915
box 0 0 120 799
use inv g8002
timestamp 1386238110
transform 1 0 23835 0 1 6915
box 0 0 120 799
use nand3 g8128
timestamp 1386234893
transform 1 0 23955 0 1 6915
box 0 0 120 799
use nand2 g8029
timestamp 1386234792
transform 1 0 24075 0 1 6915
box 0 0 96 799
use nand2 g8100
timestamp 1386234792
transform 1 0 24171 0 1 6915
box 0 0 96 799
use nand2 g8117
timestamp 1386234792
transform 1 0 24267 0 1 6915
box 0 0 96 799
use nand2 g8167
timestamp 1386234792
transform 1 0 24363 0 1 6915
box 0 0 96 799
use nand2 g7982
timestamp 1386234792
transform 1 0 24459 0 1 6915
box 0 0 96 799
use nand3 g8191
timestamp 1386234893
transform 1 0 24555 0 1 6915
box 0 0 120 799
use nand2 g8227
timestamp 1386234792
transform 1 0 24675 0 1 6915
box 0 0 96 799
use rowcrosser Op2Sel_91_0_93_
timestamp 1386086759
transform 1 0 24771 0 1 6915
box 0 0 48 799
use nand2 g7975
timestamp 1386234792
transform 1 0 24819 0 1 6915
box 0 0 96 799
use nand4 g8270
timestamp 1386234936
transform 1 0 24915 0 1 6915
box 0 0 144 799
use nand2 g8073
timestamp 1386234792
transform 1 0 25059 0 1 6915
box 0 0 96 799
use nor2 g8163
timestamp 1386235306
transform 1 0 25155 0 1 6915
box 0 0 120 799
use nand2 g8273
timestamp 1386234792
transform 1 0 25275 0 1 6915
box 0 0 96 799
use nand3 g8337
timestamp 1386234893
transform 1 0 25371 0 1 6915
box 0 0 120 799
use nand2 g8051
timestamp 1386234792
transform 1 0 25491 0 1 6915
box 0 0 96 799
use nand2 g8147
timestamp 1386234792
transform 1 0 25587 0 1 6915
box 0 0 96 799
use nand3 g8030
timestamp 1386234893
transform 1 0 25683 0 1 6915
box 0 0 120 799
use nand2 g8217
timestamp 1386234792
transform 1 0 25803 0 1 6915
box 0 0 96 799
use nand2 g8248
timestamp 1386234792
transform 1 0 25899 0 1 6915
box 0 0 96 799
use nor2 g8114
timestamp 1386235306
transform 1 0 25995 0 1 6915
box 0 0 120 799
use nand2 g8174
timestamp 1386234792
transform 1 0 26115 0 1 6915
box 0 0 96 799
use and2 g8305
timestamp 1386234845
transform 1 0 26211 0 1 6915
box 0 0 120 799
use nand2 g8241
timestamp 1386234792
transform 1 0 26331 0 1 6915
box 0 0 96 799
use nand2 g8067
timestamp 1386234792
transform 1 0 26427 0 1 6915
box 0 0 96 799
use nor2 g7990
timestamp 1386235306
transform 1 0 26523 0 1 6915
box 0 0 120 799
use nand2 g8158
timestamp 1386234792
transform 1 0 26643 0 1 6915
box 0 0 96 799
use nand2 g8063
timestamp 1386234792
transform 1 0 26739 0 1 6915
box 0 0 96 799
use nand3 g8257
timestamp 1386234893
transform 1 0 26835 0 1 6915
box 0 0 120 799
use inv ENB
timestamp 1386238110
transform 1 0 26955 0 1 6915
box 0 0 120 799
use rowcrosser AluOR_91_1_93_
timestamp 1386086759
transform 1 0 27075 0 1 6915
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27123 0 1 6915
box 0 0 320 799
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 754
box 0 0 1464 799
use nand3 stateSub_reg_91_0_93_
timestamp 1386234893
transform 1 0 1587 0 1 754
box 0 0 120 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 1707 0 1 754
box 0 0 48 799
use scandtype g8352
timestamp 1386241841
transform 1 0 1755 0 1 754
box 0 0 624 799
use inv g8150
timestamp 1386238110
transform 1 0 2379 0 1 754
box 0 0 120 799
use nand3 g8020
timestamp 1386234893
transform 1 0 2499 0 1 754
box 0 0 120 799
use nand4 g8178
timestamp 1386234936
transform 1 0 2619 0 1 754
box 0 0 144 799
use nand2 state_reg_91_1_93_
timestamp 1386234792
transform 1 0 2763 0 1 754
box 0 0 96 799
use scandtype g8250
timestamp 1386241841
transform 1 0 2859 0 1 754
box 0 0 624 799
use nand2 g8148
timestamp 1386234792
transform 1 0 3483 0 1 754
box 0 0 96 799
use nand3 g7976
timestamp 1386234893
transform 1 0 3579 0 1 754
box 0 0 120 799
use nand3 g7993
timestamp 1386234893
transform 1 0 3699 0 1 754
box 0 0 120 799
use nand3 g8196
timestamp 1386234893
transform 1 0 3819 0 1 754
box 0 0 120 799
use nor2 g8211
timestamp 1386235306
transform 1 0 3939 0 1 754
box 0 0 120 799
use nand2 g8175
timestamp 1386234792
transform 1 0 4059 0 1 754
box 0 0 96 799
use and2 g8300
timestamp 1386234845
transform 1 0 4155 0 1 754
box 0 0 120 799
use xor2 g8078
timestamp 1386237344
transform 1 0 4275 0 1 754
box 0 0 192 799
use nand2 g8093
timestamp 1386234792
transform 1 0 4467 0 1 754
box 0 0 96 799
use and2 g8104
timestamp 1386234845
transform 1 0 4563 0 1 754
box 0 0 120 799
use nand3 g8307
timestamp 1386234893
transform 1 0 4683 0 1 754
box 0 0 120 799
use nor2 g8335
timestamp 1386235306
transform 1 0 4803 0 1 754
box 0 0 120 799
use nand2 g8160
timestamp 1386234792
transform 1 0 4923 0 1 754
box 0 0 96 799
use nand2 g8076
timestamp 1386234792
transform 1 0 5019 0 1 754
box 0 0 96 799
use nor2 g8224
timestamp 1386235306
transform 1 0 5115 0 1 754
box 0 0 120 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 5235 0 1 754
box 0 0 96 799
use scandtype g8161
timestamp 1386241841
transform 1 0 5331 0 1 754
box 0 0 624 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 5955 0 1 754
box 0 0 48 799
use nand3 g8094
timestamp 1386234893
transform 1 0 6003 0 1 754
box 0 0 120 799
use and2 g8121
timestamp 1386234845
transform 1 0 6123 0 1 754
box 0 0 120 799
use nand3 g8037
timestamp 1386234893
transform 1 0 6243 0 1 754
box 0 0 120 799
use nand4 g8266
timestamp 1386234936
transform 1 0 6363 0 1 754
box 0 0 144 799
use nand3 g8189
timestamp 1386234893
transform 1 0 6507 0 1 754
box 0 0 120 799
use nand4 g8125
timestamp 1386234936
transform 1 0 6627 0 1 754
box 0 0 144 799
use nand2 g8297
timestamp 1386234792
transform 1 0 6771 0 1 754
box 0 0 96 799
use nand3 g8232
timestamp 1386234893
transform 1 0 6867 0 1 754
box 0 0 120 799
use nor2 g8152
timestamp 1386235306
transform 1 0 6987 0 1 754
box 0 0 120 799
use nand3 g8328
timestamp 1386234893
transform 1 0 7107 0 1 754
box 0 0 120 799
use nand2 g8080
timestamp 1386234792
transform 1 0 7227 0 1 754
box 0 0 96 799
use nor2 g8282
timestamp 1386235306
transform 1 0 7323 0 1 754
box 0 0 120 799
use nand2 g8267
timestamp 1386234792
transform 1 0 7443 0 1 754
box 0 0 96 799
use nand3 g8274
timestamp 1386234893
transform 1 0 7539 0 1 754
box 0 0 120 799
use and2 g8236
timestamp 1386234845
transform 1 0 7659 0 1 754
box 0 0 120 799
use nand3 g8101
timestamp 1386234893
transform 1 0 7779 0 1 754
box 0 0 120 799
use nand3 g8011
timestamp 1386234893
transform 1 0 7899 0 1 754
box 0 0 120 799
use nand2 g8185
timestamp 1386234792
transform 1 0 8019 0 1 754
box 0 0 96 799
use nand2 g8255
timestamp 1386234792
transform 1 0 8115 0 1 754
box 0 0 96 799
use nand2 g8086
timestamp 1386234792
transform 1 0 8211 0 1 754
box 0 0 96 799
use and2 g8301
timestamp 1386234845
transform 1 0 8307 0 1 754
box 0 0 120 799
use xor2 g8192
timestamp 1386237344
transform 1 0 8427 0 1 754
box 0 0 192 799
use nor2 g7988
timestamp 1386235306
transform 1 0 8619 0 1 754
box 0 0 120 799
use nor2 g8292
timestamp 1386235306
transform 1 0 8739 0 1 754
box 0 0 120 799
use and2 g8254
timestamp 1386234845
transform 1 0 8859 0 1 754
box 0 0 120 799
use nand2 g8116
timestamp 1386234792
transform 1 0 8979 0 1 754
box 0 0 96 799
use nand3 g8166
timestamp 1386234893
transform 1 0 9075 0 1 754
box 0 0 120 799
use nand2 g8145
timestamp 1386234792
transform 1 0 9195 0 1 754
box 0 0 96 799
use and2 g8001
timestamp 1386234845
transform 1 0 9291 0 1 754
box 0 0 120 799
use nand2 g8014
timestamp 1386234792
transform 1 0 9411 0 1 754
box 0 0 96 799
use nand4 g8315
timestamp 1386234936
transform 1 0 9507 0 1 754
box 0 0 144 799
use and2 g7998
timestamp 1386234845
transform 1 0 9651 0 1 754
box 0 0 120 799
use nor2 g8228
timestamp 1386235306
transform 1 0 9771 0 1 754
box 0 0 120 799
use nand2 g8342
timestamp 1386234792
transform 1 0 9891 0 1 754
box 0 0 96 799
use nand2 g7987
timestamp 1386234792
transform 1 0 9987 0 1 754
box 0 0 96 799
use nand4 g8072
timestamp 1386234936
transform 1 0 10083 0 1 754
box 0 0 144 799
use nand3 g8279
timestamp 1386234893
transform 1 0 10227 0 1 754
box 0 0 120 799
use nand2 g8105
timestamp 1386234792
transform 1 0 10347 0 1 754
box 0 0 96 799
use nand3 g8259
timestamp 1386234893
transform 1 0 10443 0 1 754
box 0 0 120 799
use nand2 g8129
timestamp 1386234792
transform 1 0 10563 0 1 754
box 0 0 96 799
use nor2 g8122
timestamp 1386235306
transform 1 0 10659 0 1 754
box 0 0 120 799
use nand2 g8059
timestamp 1386234792
transform 1 0 10779 0 1 754
box 0 0 96 799
use and2 g8097
timestamp 1386234845
transform 1 0 10875 0 1 754
box 0 0 120 799
use nand2 g8062
timestamp 1386234792
transform 1 0 10995 0 1 754
box 0 0 96 799
use rowcrosser SysBus_91_2_93_
timestamp 1386086759
transform 1 0 11091 0 1 754
box 0 0 48 799
use nand2 g8025
timestamp 1386234792
transform 1 0 11139 0 1 754
box 0 0 96 799
use nand2 g8247
timestamp 1386234792
transform 1 0 11235 0 1 754
box 0 0 96 799
use nand2 IntStatus_reg
timestamp 1386234792
transform 1 0 11331 0 1 754
box 0 0 96 799
use scanreg g8263
timestamp 1386241447
transform 1 0 11427 0 1 754
box 0 0 720 799
use rowcrosser Flags_91_0_93_
timestamp 1386086759
transform 1 0 12147 0 1 754
box 0 0 48 799
use nand2 g8256
timestamp 1386234792
transform 1 0 12195 0 1 754
box 0 0 96 799
use and2 g8087
timestamp 1386234845
transform 1 0 12291 0 1 754
box 0 0 120 799
use nand2 g8345
timestamp 1386234792
transform 1 0 12411 0 1 754
box 0 0 96 799
use and2 g8322
timestamp 1386234845
transform 1 0 12507 0 1 754
box 0 0 120 799
use nand2 g8286
timestamp 1386234792
transform 1 0 12627 0 1 754
box 0 0 96 799
use nand3 g7991
timestamp 1386234893
transform 1 0 12723 0 1 754
box 0 0 120 799
use nand2 g8201
timestamp 1386234792
transform 1 0 12843 0 1 754
box 0 0 96 799
use nand2 g8137
timestamp 1386234792
transform 1 0 12939 0 1 754
box 0 0 96 799
use nand2 g8331
timestamp 1386234792
transform 1 0 13035 0 1 754
box 0 0 96 799
use inv g8336
timestamp 1386238110
transform 1 0 13131 0 1 754
box 0 0 120 799
use nor2 g8242
timestamp 1386235306
transform 1 0 13251 0 1 754
box 0 0 120 799
use nand3 g8207
timestamp 1386234893
transform 1 0 13371 0 1 754
box 0 0 120 799
use nor2 g8044
timestamp 1386235306
transform 1 0 13491 0 1 754
box 0 0 120 799
use inv g8006
timestamp 1386238110
transform 1 0 13611 0 1 754
box 0 0 120 799
use nand4 g8173
timestamp 1386234936
transform 1 0 13731 0 1 754
box 0 0 144 799
use nand2 g7983
timestamp 1386234792
transform 1 0 13875 0 1 754
box 0 0 96 799
use nand3 g8157
timestamp 1386234893
transform 1 0 13971 0 1 754
box 0 0 120 799
use nand2 g8325
timestamp 1386234792
transform 1 0 14091 0 1 754
box 0 0 96 799
use nand2 g8040
timestamp 1386234792
transform 1 0 14187 0 1 754
box 0 0 96 799
use nand2 g8068
timestamp 1386234792
transform 1 0 14283 0 1 754
box 0 0 96 799
use nand2 g8140
timestamp 1386234792
transform 1 0 14379 0 1 754
box 0 0 96 799
use nand2 g8210
timestamp 1386234792
transform 1 0 14475 0 1 754
box 0 0 96 799
use nor2 g8141
timestamp 1386235306
transform 1 0 14571 0 1 754
box 0 0 120 799
use and2 g8003
timestamp 1386234845
transform 1 0 14691 0 1 754
box 0 0 120 799
use nand4 g8317
timestamp 1386234936
transform 1 0 14811 0 1 754
box 0 0 144 799
use inv g8203
timestamp 1386238110
transform 1 0 14955 0 1 754
box 0 0 120 799
use nand2 g8065
timestamp 1386234792
transform 1 0 15075 0 1 754
box 0 0 96 799
use nand3 g8113
timestamp 1386234893
transform 1 0 15171 0 1 754
box 0 0 120 799
use and2 g7977
timestamp 1386234845
transform 1 0 15291 0 1 754
box 0 0 120 799
use nand4 g8358
timestamp 1386234936
transform 1 0 15411 0 1 754
box 0 0 144 799
use inv g8070
timestamp 1386238110
transform 1 0 15555 0 1 754
box 0 0 120 799
use nor2 g8323
timestamp 1386235306
transform 1 0 15675 0 1 754
box 0 0 120 799
use nand2 g8309
timestamp 1386234792
transform 1 0 15795 0 1 754
box 0 0 96 799
use inv g8233
timestamp 1386238110
transform 1 0 15891 0 1 754
box 0 0 120 799
use inv IRQ2_reg
timestamp 1386238110
transform 1 0 16011 0 1 754
box 0 0 120 799
use scandtype g7980
timestamp 1386241841
transform 1 0 16131 0 1 754
box 0 0 624 799
use nand2 g8151
timestamp 1386234792
transform 1 0 16755 0 1 754
box 0 0 96 799
use nand3 g8138
timestamp 1386234893
transform 1 0 16851 0 1 754
box 0 0 120 799
use nand2 g8188
timestamp 1386234792
transform 1 0 16971 0 1 754
box 0 0 96 799
use and2 g8176
timestamp 1386234845
transform 1 0 17067 0 1 754
box 0 0 120 799
use nand2 g8172
timestamp 1386234792
transform 1 0 17187 0 1 754
box 0 0 96 799
use inv g8026
timestamp 1386238110
transform 1 0 17283 0 1 754
box 0 0 120 799
use rowcrosser SysBus_91_0_93_
timestamp 1386086759
transform 1 0 17403 0 1 754
box 0 0 48 799
use nand2 g8162
timestamp 1386234792
transform 1 0 17451 0 1 754
box 0 0 96 799
use nand2 g8031
timestamp 1386234792
transform 1 0 17547 0 1 754
box 0 0 96 799
use nand2 g8095
timestamp 1386234792
transform 1 0 17643 0 1 754
box 0 0 96 799
use nand2 g8008
timestamp 1386234792
transform 1 0 17739 0 1 754
box 0 0 96 799
use nand2 g8013
timestamp 1386234792
transform 1 0 17835 0 1 754
box 0 0 96 799
use nand3 g8299
timestamp 1386234893
transform 1 0 17931 0 1 754
box 0 0 120 799
use nor2 g8126
timestamp 1386235306
transform 1 0 18051 0 1 754
box 0 0 120 799
use nand2 g7984
timestamp 1386234792
transform 1 0 18171 0 1 754
box 0 0 96 799
use nand3 g8326
timestamp 1386234893
transform 1 0 18267 0 1 754
box 0 0 120 799
use nand2 IRQ1_reg
timestamp 1386234792
transform 1 0 18387 0 1 754
box 0 0 96 799
use scandtype g8329
timestamp 1386241841
transform 1 0 18483 0 1 754
box 0 0 624 799
use inv g7986
timestamp 1386238110
transform 1 0 19107 0 1 754
box 0 0 120 799
use nand3 rm_assigns_buf_MemEn
timestamp 1386234893
transform 1 0 19227 0 1 754
box 0 0 120 799
use buffer g8205
timestamp 1386236986
transform 1 0 19347 0 1 754
box 0 0 120 799
use and2 g8339
timestamp 1386234845
transform 1 0 19467 0 1 754
box 0 0 120 799
use inv g8164
timestamp 1386238110
transform 1 0 19587 0 1 754
box 0 0 120 799
use nand3 g8017
timestamp 1386234893
transform 1 0 19707 0 1 754
box 0 0 120 799
use nand4 g8165
timestamp 1386234936
transform 1 0 19827 0 1 754
box 0 0 144 799
use nand2 g8010
timestamp 1386234792
transform 1 0 19971 0 1 754
box 0 0 96 799
use nand4 g8260
timestamp 1386234936
transform 1 0 20067 0 1 754
box 0 0 144 799
use inv g8245
timestamp 1386238110
transform 1 0 20211 0 1 754
box 0 0 120 799
use nand2 g8034
timestamp 1386234792
transform 1 0 20331 0 1 754
box 0 0 96 799
use nand4 g8351
timestamp 1386234936
transform 1 0 20427 0 1 754
box 0 0 144 799
use inv g8215
timestamp 1386238110
transform 1 0 20571 0 1 754
box 0 0 120 799
use nand3 g8343
timestamp 1386234893
transform 1 0 20691 0 1 754
box 0 0 120 799
use inv g7999
timestamp 1386238110
transform 1 0 20811 0 1 754
box 0 0 120 799
use nand4 g8079
timestamp 1386234936
transform 1 0 20931 0 1 754
box 0 0 144 799
use and2 g8239
timestamp 1386234845
transform 1 0 21075 0 1 754
box 0 0 120 799
use and2 g8288
timestamp 1386234845
transform 1 0 21195 0 1 754
box 0 0 120 799
use nand2 g8007
timestamp 1386234792
transform 1 0 21315 0 1 754
box 0 0 96 799
use nand2 g8262
timestamp 1386234792
transform 1 0 21411 0 1 754
box 0 0 96 799
use and2 g8311
timestamp 1386234845
transform 1 0 21507 0 1 754
box 0 0 120 799
use inv g8109
timestamp 1386238110
transform 1 0 21627 0 1 754
box 0 0 120 799
use nand3 g8085
timestamp 1386234893
transform 1 0 21747 0 1 754
box 0 0 120 799
use and2 g8298
timestamp 1386234845
transform 1 0 21867 0 1 754
box 0 0 120 799
use nor2 g8346
timestamp 1386235306
transform 1 0 21987 0 1 754
box 0 0 120 799
use inv g8021
timestamp 1386238110
transform 1 0 22107 0 1 754
box 0 0 120 799
use nor2 g8184
timestamp 1386235306
transform 1 0 22227 0 1 754
box 0 0 120 799
use inv g8132
timestamp 1386238110
transform 1 0 22347 0 1 754
box 0 0 120 799
use nand2 g8355
timestamp 1386234792
transform 1 0 22467 0 1 754
box 0 0 96 799
use inv g8219
timestamp 1386238110
transform 1 0 22563 0 1 754
box 0 0 120 799
use and2 g8330
timestamp 1386234845
transform 1 0 22683 0 1 754
box 0 0 120 799
use nand2 g8061
timestamp 1386234792
transform 1 0 22803 0 1 754
box 0 0 96 799
use and2 g8360
timestamp 1386234845
transform 1 0 22899 0 1 754
box 0 0 120 799
use inv g8258
timestamp 1386238110
transform 1 0 23019 0 1 754
box 0 0 120 799
use nand2 g8115
timestamp 1386234792
transform 1 0 23139 0 1 754
box 0 0 96 799
use nand2 g8202
timestamp 1386234792
transform 1 0 23235 0 1 754
box 0 0 96 799
use and2 g8246
timestamp 1386234845
transform 1 0 23331 0 1 754
box 0 0 120 799
use nor2 g8208
timestamp 1386235306
transform 1 0 23451 0 1 754
box 0 0 120 799
use nand2 g8231
timestamp 1386234792
transform 1 0 23571 0 1 754
box 0 0 96 799
use inv g8156
timestamp 1386238110
transform 1 0 23667 0 1 754
box 0 0 120 799
use and2 g7992
timestamp 1386234845
transform 1 0 23787 0 1 754
box 0 0 120 799
use nand2 g8047
timestamp 1386234792
transform 1 0 23907 0 1 754
box 0 0 96 799
use nor2 g8179
timestamp 1386235306
transform 1 0 24003 0 1 754
box 0 0 120 799
use nand2 g8022
timestamp 1386234792
transform 1 0 24123 0 1 754
box 0 0 96 799
use nand4 g8193
timestamp 1386234936
transform 1 0 24219 0 1 754
box 0 0 144 799
use nand3 g8071
timestamp 1386234893
transform 1 0 24363 0 1 754
box 0 0 120 799
use inv g8285
timestamp 1386238110
transform 1 0 24483 0 1 754
box 0 0 120 799
use nand2 g8083
timestamp 1386234792
transform 1 0 24603 0 1 754
box 0 0 96 799
use nand2 g8204
timestamp 1386234792
transform 1 0 24699 0 1 754
box 0 0 96 799
use nand2 g8053
timestamp 1386234792
transform 1 0 24795 0 1 754
box 0 0 96 799
use nand2 g8000
timestamp 1386234792
transform 1 0 24891 0 1 754
box 0 0 96 799
use nor2 state_reg_91_0_93_
timestamp 1386235306
transform 1 0 24987 0 1 754
box 0 0 120 799
use scandtype g8142
timestamp 1386241841
transform 1 0 25107 0 1 754
box 0 0 624 799
use nand2 g8302
timestamp 1386234792
transform 1 0 25731 0 1 754
box 0 0 96 799
use nand2 stateSub_reg_91_1_93_
timestamp 1386234792
transform 1 0 25827 0 1 754
box 0 0 96 799
use scandtype g8075
timestamp 1386241841
transform 1 0 25923 0 1 754
box 0 0 624 799
use rowcrosser nWE
timestamp 1386086759
transform 1 0 26547 0 1 754
box 0 0 48 799
use nor2 SysBus_91_1_93_
timestamp 1386235306
transform 1 0 26595 0 1 754
box 0 0 120 799
use rowcrosser CFlag
timestamp 1386086759
transform 1 0 26715 0 1 754
box 0 0 48 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 26763 0 1 754
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27123 0 1 754
box 0 0 320 799
<< labels >>
rlabel m2contact 27177 7971 27177 7971 6 AluOR[0]
rlabel m2contact 27177 7779 27177 7779 6 AluOR[0]
rlabel m2contact 27153 7803 27153 7803 6 AluOR[1]
rlabel m2contact 27153 7779 27153 7779 6 AluOR[1]
rlabel m2contact 27129 7851 27129 7851 6 RwSel[1]
rlabel m2contact 27129 7731 27129 7731 6 RwSel[1]
rlabel m2contact 27105 7827 27105 7827 6 ENB
rlabel m2contact 26361 7875 26361 7875 6 StatusReg[2]
rlabel m2contact 26133 7827 26133 7827 6 StatusRegEn
rlabel m2contact 25293 7803 25293 7803 6 StatusReg[0]
rlabel m2contact 25041 7755 25041 7755 6 RegWe
rlabel m2contact 24801 7779 24801 7779 6 AluOR[1]
rlabel m2contact 24453 7779 24453 7779 6 StatusReg[1]
rlabel m2contact 24429 7875 24429 7875 6 StatusReg[2]
rlabel m2contact 23577 7827 23577 7827 6 StatusRegEn
rlabel m2contact 23217 7731 23217 7731 6 PcSel[2]
rlabel m2contact 22773 7827 22773 7827 6 StatusReg[3]
rlabel m2contact 22665 7803 22665 7803 6 StatusReg[0]
rlabel m2contact 21933 7947 21933 7947 6 AluEn
rlabel metal2 21099 7803 21099 7803 6 AluWe
rlabel m2contact 21081 7803 21081 7803 6 AluWe
rlabel m2contact 20253 7803 20253 7803 6 Op2Sel[0]
rlabel metal2 19779 7755 19779 7755 6 Op2Sel[1]
rlabel m2contact 19761 7755 19761 7755 6 Op2Sel[1]
rlabel m2contact 19713 7755 19713 7755 6 MemEn
rlabel metal2 19275 7875 19275 7875 6 Op1Sel
rlabel m2contact 19257 7875 19257 7875 6 Op1Sel
rlabel m2contact 18777 7875 18777 7875 6 WdSel
rlabel m2contact 18729 7803 18729 7803 6 Op2Sel[0]
rlabel m2contact 18549 7875 18549 7875 6 WdSel
rlabel m2contact 17841 7803 17841 7803 6 LrSel
rlabel metal2 17643 7875 17643 7875 6 PcEn
rlabel m2contact 17625 7875 17625 7875 6 PcEn
rlabel m2contact 16905 7899 16905 7899 6 LrEn
rlabel metal2 16707 7875 16707 7875 6 PcWe
rlabel m2contact 16689 7875 16689 7875 6 PcWe
rlabel m2contact 16449 7875 16449 7875 6 PcSel[0]
rlabel m2contact 16029 7875 16029 7875 6 PcSel[0]
rlabel m2contact 15561 7827 15561 7827 6 StatusReg[3]
rlabel m2contact 14913 7827 14913 7827 6 ImmSel
rlabel m2contact 14577 7875 14577 7875 6 IrWe
rlabel m2contact 14373 7923 14373 7923 6 PcSel[1]
rlabel m2contact 14349 7731 14349 7731 6 PcSel[2]
rlabel m2contact 13617 7779 13617 7779 4 StatusReg[1]
rlabel m2contact 13497 7899 13497 7899 4 LrEn
rlabel m2contact 11829 7899 11829 7899 4 LrWe
rlabel m2contact 11793 7779 11793 7779 4 OpcodeCondIn[0]
rlabel m2contact 11793 7803 11793 7803 4 LrSel
rlabel m2contact 10941 7827 10941 7827 4 ImmSel
rlabel m2contact 10905 7803 10905 7803 4 OpcodeCondIn[3]
rlabel m2contact 10089 7875 10089 7875 4 IrWe
rlabel m2contact 9993 7875 9993 7875 4 OpcodeCondIn[7]
rlabel m2contact 9657 7827 9657 7827 4 OpcodeCondIn[4]
rlabel m2contact 9237 7755 9237 7755 4 MemEn
rlabel m2contact 8385 7779 8385 7779 4 OpcodeCondIn[0]
rlabel m2contact 8001 7779 8001 7779 4 OpcodeCondIn[1]
rlabel m2contact 7533 7779 7533 7779 4 OpcodeCondIn[1]
rlabel m2contact 7449 7971 7449 7971 4 AluOR[0]
rlabel m2contact 5865 7971 5865 7971 4 OpcodeCondIn[2]
rlabel m2contact 5829 7803 5829 7803 4 OpcodeCondIn[3]
rlabel m2contact 5409 7971 5409 7971 4 OpcodeCondIn[2]
rlabel m2contact 4977 7827 4977 7827 4 OpcodeCondIn[4]
rlabel m2contact 4401 7851 4401 7851 4 RwSel[1]
rlabel m2contact 3945 7947 3945 7947 4 AluEn
rlabel m2contact 3657 7899 3657 7899 4 LrWe
rlabel m2contact 3309 7899 3309 7899 4 OpcodeCondIn[5]
rlabel m2contact 2457 7947 2457 7947 4 OpcodeCondIn[6]
rlabel m2contact 2421 7875 2421 7875 4 OpcodeCondIn[7]
rlabel m2contact 2385 7947 2385 7947 4 OpcodeCondIn[6]
rlabel m2contact 2193 7899 2193 7899 4 OpcodeCondIn[5]
rlabel m2contact 2001 7923 2001 7923 4 PcSel[1]
rlabel m2contact 1761 7899 1761 7899 4 nME
rlabel m2contact 1713 7923 1713 7923 4 ALE
rlabel m2contact 27153 3634 27153 3634 6 Rs1Sel[0]
rlabel m2contact 27153 1594 27153 1594 6 Rs1Sel[0]
rlabel m2contact 27129 4258 27129 4258 6 Flags[3]
rlabel m2contact 27129 1570 27129 1570 6 Flags[3]
rlabel m2contact 27105 1762 27105 1762 6 ENB
rlabel m2contact 27033 3370 27033 3370 6 n_179
rlabel m2contact 26985 4402 26985 4402 6 n_266
rlabel m2contact 26937 2914 26937 2914 6 n_254
rlabel m2contact 26913 5002 26913 5002 6 n_70
rlabel m2contact 26889 5938 26889 5938 6 n_163
rlabel m2contact 26865 6346 26865 6346 6 n_121
rlabel m2contact 26841 4522 26841 4522 6 Flags[2]
rlabel m2contact 26841 3178 26841 3178 6 Flags[2]
rlabel m2contact 26817 2458 26817 2458 6 n_132
rlabel m2contact 26793 3178 26793 3178 6 Flags[2]
rlabel m2contact 26793 3202 26793 3202 6 n_39
rlabel m2contact 26769 4426 26769 4426 6 n_86
rlabel m2contact 26745 6706 26745 6706 6 Flags[1]
rlabel m2contact 26721 4234 26721 4234 6 n_310
rlabel m2contact 26697 6394 26697 6394 6 CFlag
rlabel m2contact 26673 5674 26673 5674 6 n_309
rlabel m2contact 26649 4498 26649 4498 6 n_286
rlabel m2contact 26649 4354 26649 4354 6 n_286
rlabel m2contact 26625 4498 26625 4498 6 n_286
rlabel m2contact 26625 4474 26625 4474 6 n_91
rlabel m2contact 26577 6394 26577 6394 6 CFlag
rlabel m2contact 26577 6538 26577 6538 6 n_238
rlabel m2contact 26553 1954 26553 1954 6 n_221
rlabel m2contact 26505 5650 26505 5650 6 n_116
rlabel m2contact 26481 4810 26481 4810 6 stateSub[1]
rlabel m2contact 26457 2650 26457 2650 6 n_133
rlabel m2contact 26433 4810 26433 4810 6 stateSub[1]
rlabel m2contact 26409 4018 26409 4018 6 n_55
rlabel m2contact 26385 5554 26385 5554 6 n_398
rlabel m2contact 26385 1714 26385 1714 6 n_123
rlabel m2contact 26361 2578 26361 2578 6 StatusReg[2]
rlabel m2contact 26313 2410 26313 2410 6 n_226
rlabel m2contact 26265 2842 26265 2842 6 n_144
rlabel m2contact 26241 6274 26241 6274 6 n_157
rlabel m2contact 26193 2482 26193 2482 6 n_236
rlabel m2contact 26169 5218 26169 5218 6 n_152
rlabel m2contact 26145 3778 26145 3778 6 n_258
rlabel m2contact 26097 5746 26097 5746 6 n_64
rlabel m2contact 26049 6562 26049 6562 6 n_232
rlabel m2contact 26025 5074 26025 5074 6 n_13
rlabel m2contact 25977 4378 25977 4378 6 n_119
rlabel m2contact 25953 2506 25953 2506 6 OpcodeCondIn[3]
rlabel m2contact 25929 4306 25929 4306 6 n_128
rlabel m2contact 25905 6874 25905 6874 6 n_330
rlabel m2contact 25905 4138 25905 4138 6 n_330
rlabel m2contact 25881 6874 25881 6874 6 n_330
rlabel m2contact 25881 6850 25881 6850 6 n_54
rlabel m2contact 25857 4258 25857 4258 6 Flags[3]
rlabel m2contact 25857 4018 25857 4018 6 n_55
rlabel m2contact 25833 5506 25833 5506 6 n_332
rlabel m2contact 25809 5842 25809 5842 6 n_278
rlabel m2contact 25809 4210 25809 4210 6 n_278
rlabel m2contact 25785 2458 25785 2458 6 n_132
rlabel m2contact 25785 2530 25785 2530 6 n_276
rlabel m2contact 25761 4210 25761 4210 6 n_278
rlabel m2contact 25761 4258 25761 4258 6 n_231
rlabel m2contact 25737 6442 25737 6442 6 n_263
rlabel m2contact 25713 3466 25713 3466 6 n_241
rlabel m2contact 25665 4330 25665 4330 6 n_294
rlabel m2contact 25641 2290 25641 2290 6 SysBus[1]
rlabel m2contact 25617 5482 25617 5482 6 n_293
rlabel m2contact 25617 3874 25617 3874 6 state[0]
rlabel m2contact 25593 4738 25593 4738 6 n_7
rlabel m2contact 25593 2242 25593 2242 6 n_7
rlabel m2contact 25569 4738 25569 4738 6 n_7
rlabel m2contact 25569 4714 25569 4714 6 n_63
rlabel m2contact 25545 4810 25545 4810 6 stateSub[1]
rlabel m2contact 25521 3586 25521 3586 6 n_114
rlabel m2contact 25473 4786 25473 4786 6 n_299
rlabel m2contact 25449 1714 25449 1714 6 n_123
rlabel m2contact 25425 2266 25425 2266 6 n_78
rlabel m2contact 25401 3274 25401 3274 6 state[1]
rlabel m2contact 25353 4090 25353 4090 6 n_217
rlabel m2contact 25329 3970 25329 3970 6 n_219
rlabel m2contact 25305 6274 25305 6274 6 n_157
rlabel m2contact 25257 3802 25257 3802 6 n_213
rlabel m2contact 25209 4762 25209 4762 6 n_211
rlabel m2contact 25185 2698 25185 2698 6 n_212
rlabel m2contact 25137 6178 25137 6178 6 n_60
rlabel m2contact 25113 5914 25113 5914 6 stateSub[2]
rlabel m2contact 25089 6610 25089 6610 6 n_58
rlabel m2contact 25041 4282 25041 4282 6 n_209
rlabel m2contact 25017 3226 25017 3226 6 n_377
rlabel m2contact 24993 1810 24993 1810 6 n_375
rlabel m2contact 24969 1786 24969 1786 6 n_307
rlabel m2contact 24945 4066 24945 4066 6 n_178
rlabel m2contact 24921 5482 24921 5482 6 n_293
rlabel m2contact 24897 4426 24897 4426 6 n_86
rlabel m2contact 24873 4186 24873 4186 6 OpcodeCondIn[5]
rlabel m2contact 24849 1714 24849 1714 6 n_123
rlabel m2contact 24849 5290 24849 5290 6 n_53
rlabel m2contact 24825 2650 24825 2650 6 n_133
rlabel m2contact 24801 4042 24801 4042 6 AluOR[1]
rlabel m2contact 24753 4210 24753 4210 6 n_173
rlabel m2contact 24753 5386 24753 5386 6 n_93
rlabel m2contact 24729 3442 24729 3442 6 n_44
rlabel m2contact 24729 2866 24729 2866 6 n_106
rlabel m2contact 24705 1666 24705 1666 6 n_41
rlabel m2contact 24681 6874 24681 6874 6 n_98
rlabel m2contact 24681 4450 24681 4450 6 n_98
rlabel m2contact 24657 5338 24657 5338 6 n_360
rlabel m2contact 24657 1618 24657 1618 6 n_22
rlabel m2contact 24633 4330 24633 4330 6 n_294
rlabel m2contact 24633 2266 24633 2266 6 n_78
rlabel m2contact 24609 4234 24609 4234 6 n_310
rlabel m2contact 24585 5410 24585 5410 6 n_333
rlabel m2contact 24561 4162 24561 4162 6 n_340
rlabel m2contact 24537 3826 24537 3826 6 n_181
rlabel m2contact 24513 2026 24513 2026 6 n_36
rlabel m2contact 24513 1786 24513 1786 6 n_307
rlabel m2contact 24489 3490 24489 3490 6 n_229
rlabel m2contact 24465 4234 24465 4234 6 n_69
rlabel m2contact 24441 5170 24441 5170 6 n_196
rlabel m2contact 24441 4114 24441 4114 6 OpcodeCondIn[0]
rlabel m2contact 24417 4018 24417 4018 6 n_55
rlabel m2contact 24417 4426 24417 4426 6 n_195
rlabel m2contact 24393 6874 24393 6874 6 n_98
rlabel m2contact 24393 6850 24393 6850 6 n_54
rlabel m2contact 24369 4546 24369 4546 6 n_331
rlabel m2contact 24369 1642 24369 1642 6 n_331
rlabel m2contact 24345 4042 24345 4042 6 AluOR[1]
rlabel m2contact 24345 4330 24345 4330 6 n_174
rlabel m2contact 24321 4210 24321 4210 6 n_173
rlabel m2contact 24321 3226 24321 3226 6 n_377
rlabel m2contact 24297 3322 24297 3322 6 n_288
rlabel m2contact 24297 5914 24297 5914 6 stateSub[2]
rlabel m2contact 24261 4498 24261 4498 6 n_303
rlabel m2contact 24261 3346 24261 3346 6 n_303
rlabel m2contact 24249 4546 24249 4546 6 n_331
rlabel m2contact 24249 2986 24249 2986 6 n_322
rlabel m2contact 24225 4522 24225 4522 6 Flags[2]
rlabel m2contact 24201 4066 24201 4066 6 n_178
rlabel m2contact 24201 5506 24201 5506 6 n_332
rlabel m2contact 24177 6562 24177 6562 6 n_232
rlabel m2contact 24153 4498 24153 4498 6 n_303
rlabel m2contact 24153 3490 24153 3490 6 n_229
rlabel m2contact 24129 5794 24129 5794 6 n_29
rlabel m2contact 24105 5842 24105 5842 6 n_278
rlabel m2contact 24105 3178 24105 3178 6 n_339
rlabel m2contact 24081 4570 24081 4570 6 LrSel
rlabel m2contact 24081 3562 24081 3562 6 LrSel
rlabel m2contact 24057 3802 24057 3802 6 n_213
rlabel m2contact 24057 3850 24057 3850 6 n_357
rlabel m2contact 24033 3562 24033 3562 6 LrSel
rlabel m2contact 24033 3610 24033 3610 6 stateSub[0]
rlabel m2contact 24009 3538 24009 3538 6 n_318
rlabel m2contact 23985 5770 23985 5770 6 n_284
rlabel m2contact 23961 5026 23961 5026 6 StatusReg[3]
rlabel m2contact 23937 5674 23937 5674 6 n_309
rlabel m2contact 23913 4450 23913 4450 6 n_98
rlabel m2contact 23889 6058 23889 6058 6 n_161
rlabel m2contact 23865 6658 23865 6658 6 n_97
rlabel m2contact 23841 5962 23841 5962 6 n_249
rlabel m2contact 23817 4018 23817 4018 6 n_329
rlabel m2contact 23817 3106 23817 3106 6 n_184
rlabel m2contact 23769 6634 23769 6634 6 n_166
rlabel m2contact 23745 4354 23745 4354 6 n_286
rlabel m2contact 23697 5314 23697 5314 6 n_94
rlabel m2contact 23697 4066 23697 4066 6 n_94
rlabel m2contact 23673 2722 23673 2722 6 n_215
rlabel m2contact 23649 5098 23649 5098 6 n_108
rlabel m2contact 23625 4066 23625 4066 6 n_94
rlabel m2contact 23625 4762 23625 4762 6 n_211
rlabel m2contact 23601 3754 23601 3754 6 n_234
rlabel m2contact 23553 4738 23553 4738 6 n_217
rlabel m2contact 23553 4090 23553 4090 6 n_217
rlabel m2contact 23529 3394 23529 3394 6 n_188
rlabel m2contact 23505 4738 23505 4738 6 n_217
rlabel m2contact 23505 4690 23505 4690 6 OpcodeCondIn[1]
rlabel m2contact 23481 6682 23481 6682 6 n_75
rlabel m2contact 23457 4282 23457 4282 6 n_209
rlabel m2contact 23433 4594 23433 4594 6 n_186
rlabel m2contact 23409 3778 23409 3778 6 n_258
rlabel m2contact 23385 4042 23385 4042 6 n_167
rlabel m2contact 23385 3754 23385 3754 6 n_234
rlabel m2contact 23361 3130 23361 3130 6 n_145
rlabel m2contact 23337 4642 23337 4642 6 n_68
rlabel m2contact 23313 5146 23313 5146 6 n_17
rlabel m2contact 23313 4930 23313 4930 6 n_198
rlabel m2contact 23289 5962 23289 5962 6 n_249
rlabel m2contact 23265 2002 23265 2002 6 n_197
rlabel m2contact 23241 6082 23241 6082 6 n_257
rlabel m2contact 23241 3994 23241 3994 6 n_257
rlabel m2contact 23217 4402 23217 4402 6 n_266
rlabel m2contact 23193 4258 23193 4258 6 n_231
rlabel m2contact 23169 3994 23169 3994 6 n_257
rlabel m2contact 23169 4066 23169 4066 6 n_349
rlabel m2contact 23121 3946 23121 3946 6 n_208
rlabel m2contact 23097 3778 23097 3778 6 n_258
rlabel m2contact 23073 4738 23073 4738 6 n_200
rlabel m2contact 23049 3754 23049 3754 6 n_234
rlabel m2contact 23025 6130 23025 6130 6 n_255
rlabel m2contact 23025 3994 23025 3994 6 n_255
rlabel m2contact 23001 3994 23001 3994 6 n_255
rlabel m2contact 23001 4666 23001 4666 6 n_110
rlabel m2contact 22953 5458 22953 5458 6 OpcodeCondIn[2]
rlabel m2contact 22929 4234 22929 4234 6 n_69
rlabel m2contact 22881 5266 22881 5266 6 n_65
rlabel m2contact 22857 4234 22857 4234 6 n_82
rlabel m2contact 22857 2338 22857 2338 6 OpcodeCondIn[7]
rlabel m2contact 22809 2002 22809 2002 6 n_197
rlabel m2contact 22785 2098 22785 2098 6 n_155
rlabel m2contact 22737 3370 22737 3370 6 n_179
rlabel m2contact 22713 3130 22713 3130 6 n_145
rlabel m2contact 22665 5698 22665 5698 6 StatusReg[0]
rlabel m2contact 22617 6034 22617 6034 6 n_399
rlabel m2contact 22593 4282 22593 4282 6 OpcodeCondIn[6]
rlabel m2contact 22545 4210 22545 4210 6 n_173
rlabel m2contact 22521 4498 22521 4498 6 n_103
rlabel m2contact 22425 2194 22425 2194 6 n_243
rlabel m2contact 22377 2170 22377 2170 6 n_189
rlabel m2contact 22257 4018 22257 4018 6 n_329
rlabel m2contact 22257 5722 22257 5722 6 n_367
rlabel m2contact 22233 6610 22233 6610 6 n_58
rlabel m2contact 22233 4210 22233 4210 6 n_58
rlabel m2contact 22209 6010 22209 6010 6 n_203
rlabel m2contact 22209 1690 22209 1690 6 n_203
rlabel m2contact 22185 5866 22185 5866 6 n_43
rlabel m2contact 22161 6586 22161 6586 6 n_299
rlabel m2contact 22161 4786 22161 4786 6 n_299
rlabel m2contact 22137 6634 22137 6634 6 n_166
rlabel m2contact 22113 3106 22113 3106 6 n_184
rlabel m2contact 22089 4906 22089 4906 6 n_23
rlabel m2contact 22089 3898 22089 3898 6 n_23
rlabel m2contact 22065 4378 22065 4378 6 n_119
rlabel m2contact 22041 4450 22041 4450 6 n_5
rlabel m2contact 22017 4210 22017 4210 6 n_58
rlabel m2contact 22017 5242 22017 5242 6 n_130
rlabel m2contact 21993 3586 21993 3586 6 n_114
rlabel m2contact 21969 3658 21969 3658 6 n_90
rlabel m2contact 21945 5434 21945 5434 6 n_319
rlabel m2contact 21945 4018 21945 4018 6 n_319
rlabel m2contact 21921 5530 21921 5530 6 n_141
rlabel m2contact 21897 3346 21897 3346 6 n_303
rlabel m2contact 21897 4522 21897 4522 6 n_267
rlabel m2contact 21873 4858 21873 4858 6 n_114
rlabel m2contact 21873 3586 21873 3586 6 n_114
rlabel m2contact 21849 1690 21849 1690 6 n_203
rlabel m2contact 21849 1738 21849 1738 6 n_101
rlabel m2contact 21825 3562 21825 3562 6 n_202
rlabel m2contact 21801 5578 21801 5578 6 n_351
rlabel m2contact 21801 3490 21801 3490 6 n_229
rlabel m2contact 21777 6586 21777 6586 6 n_299
rlabel m2contact 21777 6562 21777 6562 6 n_232
rlabel m2contact 21753 6370 21753 6370 6 n_312
rlabel m2contact 21729 2386 21729 2386 6 n_227
rlabel m2contact 21705 2146 21705 2146 6 n_139
rlabel m2contact 21705 4618 21705 4618 6 n_154
rlabel m2contact 21681 4642 21681 4642 6 n_68
rlabel m2contact 21681 3730 21681 3730 6 n_68
rlabel m2contact 21657 3898 21657 3898 6 n_23
rlabel m2contact 21657 3922 21657 3922 6 n_85
rlabel m2contact 21633 4834 21633 4834 6 n_373
rlabel m2contact 21633 3082 21633 3082 6 n_373
rlabel m2contact 21609 2314 21609 2314 6 n_59
rlabel m2contact 21585 1978 21585 1978 6 n_84
rlabel m2contact 21561 3754 21561 3754 6 n_234
rlabel m2contact 21537 6274 21537 6274 6 n_157
rlabel m2contact 21513 5818 21513 5818 6 n_170
rlabel m2contact 21513 4978 21513 4978 6 n_170
rlabel m2contact 21513 4546 21513 4546 6 n_280
rlabel m2contact 21513 2458 21513 2458 6 n_280
rlabel m2contact 21489 3754 21489 3754 6 n_234
rlabel m2contact 21465 4018 21465 4018 6 n_319
rlabel m2contact 21465 4522 21465 4522 6 n_267
rlabel m2contact 21441 4210 21441 4210 6 n_273
rlabel m2contact 21417 4354 21417 4354 6 n_248
rlabel m2contact 21393 5314 21393 5314 6 n_94
rlabel m2contact 21369 6322 21369 6322 6 n_199
rlabel m2contact 21369 2506 21369 2506 6 OpcodeCondIn[3]
rlabel m2contact 21345 4954 21345 4954 6 n_240
rlabel m2contact 21345 4258 21345 4258 6 n_231
rlabel m2contact 21309 5890 21309 5890 6 n_113
rlabel m2contact 21309 2794 21309 2794 6 n_113
rlabel m2contact 21297 6586 21297 6586 6 n_21
rlabel m2contact 21273 3754 21273 3754 6 n_234
rlabel m2contact 21249 4858 21249 4858 6 n_114
rlabel m2contact 21249 3994 21249 3994 6 n_153
rlabel m2contact 21213 5602 21213 5602 6 n_26
rlabel m2contact 21213 2602 21213 2602 6 n_26
rlabel m2contact 21201 6202 21201 6202 6 n_35
rlabel m2contact 21177 2050 21177 2050 6 Op1Sel
rlabel m2contact 21153 5266 21153 5266 6 n_65
rlabel m2contact 21129 3730 21129 3730 6 n_68
rlabel m2contact 21129 3778 21129 3778 6 n_258
rlabel m2contact 21105 5434 21105 5434 6 n_319
rlabel m2contact 21081 5986 21081 5986 6 n_25
rlabel m2contact 21081 2770 21081 2770 6 n_25
rlabel m2contact 21057 5818 21057 5818 6 n_170
rlabel m2contact 21057 5674 21057 5674 6 n_309
rlabel m2contact 21033 4834 21033 4834 6 n_373
rlabel m2contact 21033 4402 21033 4402 6 n_266
rlabel m2contact 21009 3058 21009 3058 6 n_371
rlabel m2contact 20985 6226 20985 6226 6 n_324
rlabel m2contact 20961 4522 20961 4522 6 n_267
rlabel m2contact 20937 4498 20937 4498 6 n_103
rlabel m2contact 20913 4306 20913 4306 6 n_128
rlabel m2contact 20889 5050 20889 5050 6 n_79
rlabel m2contact 20865 5866 20865 5866 6 n_43
rlabel m2contact 20865 3034 20865 3034 6 n_43
rlabel m2contact 20841 4834 20841 4834 6 n_33
rlabel m2contact 20817 3418 20817 3418 6 n_301
rlabel m2contact 20793 2818 20793 2818 6 n_87
rlabel m2contact 20769 4546 20769 4546 6 n_280
rlabel m2contact 20769 2722 20769 2722 6 n_215
rlabel m2contact 20745 4498 20745 4498 6 n_245
rlabel m2contact 20721 6154 20721 6154 6 n_71
rlabel m2contact 20721 3994 20721 3994 6 n_153
rlabel m2contact 20697 6250 20697 6250 6 n_19
rlabel m2contact 20673 6082 20673 6082 6 n_257
rlabel m2contact 20649 6082 20649 6082 6 n_257
rlabel m2contact 20625 4858 20625 4858 6 n_260
rlabel m2contact 20601 2338 20601 2338 6 OpcodeCondIn[7]
rlabel m2contact 20577 3106 20577 3106 6 n_184
rlabel m2contact 20553 3490 20553 3490 6 n_229
rlabel m2contact 20529 4810 20529 4810 6 stateSub[1]
rlabel m2contact 20505 5890 20505 5890 6 n_113
rlabel m2contact 20505 5818 20505 5818 6 n_118
rlabel m2contact 20481 5602 20481 5602 6 n_26
rlabel m2contact 20481 5362 20481 5362 6 n_346
rlabel m2contact 20457 2482 20457 2482 6 n_236
rlabel m2contact 20457 2554 20457 2554 6 n_73
rlabel m2contact 20433 5122 20433 5122 6 n_308
rlabel m2contact 20433 2938 20433 2938 6 n_308
rlabel m2contact 20409 3442 20409 3442 6 n_44
rlabel m2contact 20409 3514 20409 3514 6 n_146
rlabel m2contact 20385 2770 20385 2770 6 n_25
rlabel m2contact 20385 2842 20385 2842 6 n_144
rlabel m2contact 20361 3034 20361 3034 6 n_43
rlabel m2contact 20361 3130 20361 3130 6 n_145
rlabel m2contact 20325 6106 20325 6106 6 n_274
rlabel m2contact 20325 3898 20325 3898 6 n_274
rlabel m2contact 20313 6874 20313 6874 6 n_336
rlabel m2contact 20289 2650 20289 2650 6 n_133
rlabel m2contact 20265 4354 20265 4354 6 n_248
rlabel m2contact 20241 5122 20241 5122 6 n_308
rlabel m2contact 20241 4882 20241 4882 6 n_81
rlabel m2contact 20217 5890 20217 5890 6 n_223
rlabel m2contact 20217 4018 20217 4018 6 n_223
rlabel m2contact 20193 4978 20193 4978 6 n_170
rlabel m2contact 20193 4354 20193 4354 6 PcWe
rlabel m2contact 20169 4546 20169 4546 6 n_169
rlabel m2contact 20169 4066 20169 4066 6 n_349
rlabel m2contact 20145 2098 20145 2098 6 n_155
rlabel m2contact 20121 3010 20121 3010 6 n_242
rlabel m2contact 20121 4498 20121 4498 6 n_245
rlabel m2contact 20097 3826 20097 3826 6 n_181
rlabel m2contact 20073 4474 20073 4474 6 n_91
rlabel m2contact 20049 4978 20049 4978 6 Op2Sel[1]
rlabel m2contact 20049 3730 20049 3730 6 Op2Sel[1]
rlabel m2contact 20025 5914 20025 5914 6 stateSub[2]
rlabel m2contact 20025 4474 20025 4474 6 n_159
rlabel m2contact 20001 6202 20001 6202 6 n_35
rlabel m2contact 20001 5770 20001 5770 6 n_284
rlabel m2contact 19977 5626 19977 5626 6 n_106
rlabel m2contact 19977 2866 19977 2866 6 n_106
rlabel m2contact 19953 5602 19953 5602 6 n_34
rlabel m2contact 19953 3802 19953 3802 6 nOE
rlabel m2contact 19929 4906 19929 4906 6 n_23
rlabel m2contact 19905 3898 19905 3898 6 n_274
rlabel m2contact 19905 4834 19905 4834 6 n_33
rlabel m2contact 19881 3946 19881 3946 6 n_208
rlabel m2contact 19857 6106 19857 6106 6 n_274
rlabel m2contact 19857 5194 19857 5194 6 n_140
rlabel m2contact 19833 3106 19833 3106 6 n_184
rlabel m2contact 19809 5890 19809 5890 6 n_223
rlabel m2contact 19809 5122 19809 5122 6 n_72
rlabel m2contact 19785 5002 19785 5002 6 n_70
rlabel m2contact 19761 4978 19761 4978 6 Op2Sel[1]
rlabel m2contact 19761 3778 19761 3778 6 n_258
rlabel m2contact 19737 6154 19737 6154 6 n_71
rlabel m2contact 19713 3154 19713 3154 6 MemEn
rlabel m2contact 19677 6106 19677 6106 6 n_96
rlabel m2contact 19677 4978 19677 4978 6 n_96
rlabel m2contact 19665 3250 19665 3250 6 n_177
rlabel m2contact 19641 3826 19641 3826 6 n_365
rlabel m2contact 19617 5794 19617 5794 6 n_29
rlabel m2contact 19593 5578 19593 5578 6 n_351
rlabel m2contact 19569 2842 19569 2842 6 n_144
rlabel m2contact 19545 3898 19545 3898 6 n_107
rlabel m2contact 19521 6106 19521 6106 6 n_96
rlabel m2contact 19521 6082 19521 6082 6 n_257
rlabel m2contact 19497 5626 19497 5626 6 n_106
rlabel m2contact 19497 4306 19497 4306 6 n_128
rlabel m2contact 19473 5578 19473 5578 6 n_78
rlabel m2contact 19473 2266 19473 2266 6 n_78
rlabel m2contact 19449 1690 19449 1690 6 n_265
rlabel m2contact 19425 3154 19425 3154 6 MemEn
rlabel m2contact 19425 3226 19425 3226 6 n_377
rlabel m2contact 19401 3442 19401 3442 6 n_205
rlabel m2contact 19377 1762 19377 1762 6 ENB
rlabel m2contact 19353 3946 19353 3946 6 n_88
rlabel m2contact 19329 3730 19329 3730 6 Op2Sel[1]
rlabel m2contact 19329 5602 19329 5602 6 n_34
rlabel m2contact 19305 5578 19305 5578 6 n_78
rlabel m2contact 19305 3226 19305 3226 6 n_377
rlabel m2contact 19281 3826 19281 3826 6 n_365
rlabel m2contact 19257 2050 19257 2050 6 Op1Sel
rlabel m2contact 19209 5410 19209 5410 6 n_333
rlabel m2contact 19185 6706 19185 6706 6 Flags[1]
rlabel m2contact 19185 6562 19185 6562 6 n_232
rlabel m2contact 19161 5506 19161 5506 6 n_332
rlabel m2contact 19137 5266 19137 5266 6 n_65
rlabel m2contact 19113 4906 19113 4906 6 n_23
rlabel m2contact 19089 3778 19089 3778 6 n_258
rlabel m2contact 19065 1714 19065 1714 6 n_123
rlabel m2contact 18993 6346 18993 6346 6 n_121
rlabel m2contact 18945 4978 18945 4978 6 n_96
rlabel m2contact 18873 5770 18873 5770 6 n_284
rlabel m2contact 18825 1618 18825 1618 6 n_22
rlabel m2contact 18777 2674 18777 2674 6 WdSel
rlabel m2contact 18729 3154 18729 3154 6 Op2Sel[0]
rlabel m2contact 18585 6394 18585 6394 6 CFlag
rlabel m2contact 18465 4906 18465 4906 6 n_11
rlabel m2contact 18441 1714 18441 1714 6 n_123
rlabel m2contact 18417 3274 18417 3274 6 state[1]
rlabel m2contact 18369 5626 18369 5626 6 n_358
rlabel m2contact 18297 4138 18297 4138 6 n_330
rlabel m2contact 18249 5890 18249 5890 6 n_279
rlabel m2contact 18201 5842 18201 5842 6 n_278
rlabel m2contact 18177 5338 18177 5338 6 n_360
rlabel m2contact 18153 5362 18153 5362 6 n_346
rlabel m2contact 18105 3298 18105 3298 6 n_16
rlabel m2contact 18081 6610 18081 6610 6 n_58
rlabel m2contact 18057 3394 18057 3394 6 n_188
rlabel m2contact 18033 3154 18033 3154 6 Op2Sel[0]
rlabel m2contact 18033 3250 18033 3250 6 n_177
rlabel m2contact 18009 4306 18009 4306 6 n_128
rlabel m2contact 17985 6706 17985 6706 6 n_31
rlabel m2contact 17985 1906 17985 1906 6 n_31
rlabel m2contact 17961 6706 17961 6706 6 n_31
rlabel m2contact 17961 6514 17961 6514 6 n_233
rlabel m2contact 17937 3034 17937 3034 6 OpcodeCondIn[4]
rlabel m2contact 17913 3682 17913 3682 6 nME
rlabel m2contact 17913 3778 17913 3778 6 n_258
rlabel m2contact 17889 1978 17889 1978 6 n_84
rlabel m2contact 17889 2338 17889 2338 6 OpcodeCondIn[7]
rlabel m2contact 17865 6802 17865 6802 6 n_122
rlabel m2contact 17865 1594 17865 1594 6 n_122
rlabel m2contact 17841 4570 17841 4570 6 LrSel
rlabel m2contact 17805 5914 17805 5914 6 stateSub[2]
rlabel m2contact 17805 3730 17805 3730 6 stateSub[2]
rlabel m2contact 17793 6418 17793 6418 6 n_102
rlabel m2contact 17793 3154 17793 3154 6 n_268
rlabel m2contact 17769 4138 17769 4138 6 n_269
rlabel m2contact 17769 5338 17769 5338 6 n_400
rlabel m2contact 17745 5410 17745 5410 6 n_368
rlabel m2contact 17745 1834 17745 1834 6 n_368
rlabel m2contact 17721 3538 17721 3538 6 n_318
rlabel m2contact 17721 3706 17721 3706 6 n_77
rlabel m2contact 17697 3826 17697 3826 6 nWait
rlabel m2contact 17673 3730 17673 3730 6 stateSub[2]
rlabel m2contact 17673 4498 17673 4498 6 n_245
rlabel m2contact 17649 6730 17649 6730 6 n_142
rlabel m2contact 17649 2890 17649 2890 6 n_142
rlabel m2contact 17625 3730 17625 3730 6 PcEn
rlabel m2contact 17625 3538 17625 3538 6 n_158
rlabel m2contact 17601 5602 17601 5602 6 n_193
rlabel m2contact 17577 1594 17577 1594 6 n_122
rlabel m2contact 17577 1858 17577 1858 6 n_207
rlabel m2contact 17553 4810 17553 4810 6 stateSub[1]
rlabel m2contact 17529 5578 17529 5578 6 n_165
rlabel m2contact 17505 3514 17505 3514 6 n_146
rlabel m2contact 17481 5410 17481 5410 6 n_368
rlabel m2contact 17481 2218 17481 2218 6 n_259
rlabel m2contact 17457 4570 17457 4570 6 n_160
rlabel m2contact 17433 6874 17433 6874 6 n_336
rlabel m2contact 17433 6826 17433 6826 6 SysBus[2]
rlabel m2contact 17409 6298 17409 6298 6 n_250
rlabel m2contact 17385 2362 17385 2362 6 n_264
rlabel m2contact 17361 5842 17361 5842 6 n_278
rlabel m2contact 17337 4450 17337 4450 6 n_5
rlabel m2contact 17313 6490 17313 6490 6 n_214
rlabel m2contact 17289 3826 17289 3826 6 nWait
rlabel m2contact 17265 2890 17265 2890 6 n_142
rlabel m2contact 17265 3274 17265 3274 6 state[1]
rlabel m2contact 17241 3898 17241 3898 6 n_107
rlabel m2contact 17217 4450 17217 4450 6 n_99
rlabel m2contact 17217 5506 17217 5506 6 n_332
rlabel m2contact 17193 5410 17193 5410 6 n_182
rlabel m2contact 17169 6010 17169 6010 6 n_203
rlabel m2contact 17145 5890 17145 5890 6 n_279
rlabel m2contact 17121 3154 17121 3154 6 n_268
rlabel m2contact 17097 2098 17097 2098 6 n_155
rlabel m2contact 17073 2122 17073 2122 6 n_127
rlabel m2contact 17049 4042 17049 4042 6 n_167
rlabel m2contact 17049 5746 17049 5746 6 n_64
rlabel m2contact 17025 6634 17025 6634 6 n_166
rlabel m2contact 17001 2122 17001 2122 6 n_127
rlabel m2contact 17001 2338 17001 2338 6 OpcodeCondIn[7]
rlabel m2contact 16977 3562 16977 3562 6 n_202
rlabel m2contact 16953 3322 16953 3322 6 n_288
rlabel m2contact 16929 3970 16929 3970 6 n_219
rlabel m2contact 16905 3490 16905 3490 6 n_229
rlabel m2contact 16881 6466 16881 6466 6 n_228
rlabel m2contact 16881 3514 16881 3514 6 n_204
rlabel m2contact 16857 4042 16857 4042 6 n_354
rlabel m2contact 16809 2482 16809 2482 6 n_134
rlabel m2contact 16809 3082 16809 3082 6 n_373
rlabel m2contact 16785 3898 16785 3898 6 n_370
rlabel m2contact 16761 3226 16761 3226 6 n_377
rlabel m2contact 16737 5746 16737 5746 6 n_261
rlabel m2contact 16689 4354 16689 4354 6 PcWe
rlabel m2contact 16641 2746 16641 2746 6 n_285
rlabel m2contact 16641 2626 16641 2626 6 IRQ2
rlabel m2contact 16617 5770 16617 5770 6 n_284
rlabel m2contact 16593 4354 16593 4354 6 n_256
rlabel m2contact 16545 4978 16545 4978 6 n_96
rlabel m2contact 16521 4258 16521 4258 6 n_231
rlabel m2contact 16497 5266 16497 5266 6 n_65
rlabel m2contact 16449 1930 16449 1930 6 PcSel[0]
rlabel m2contact 16305 5914 16305 5914 6 stateSub[2]
rlabel m2contact 16257 3754 16257 3754 6 n_234
rlabel m2contact 16089 3514 16089 3514 6 n_204
rlabel m2contact 16041 3394 16041 3394 6 n_188
rlabel m2contact 15969 4258 15969 4258 6 n_231
rlabel m2contact 15921 6010 15921 6010 6 n_40
rlabel m2contact 15897 6202 15897 6202 6 n_315
rlabel m2contact 15873 2770 15873 2770 6 n_10
rlabel m2contact 15849 2506 15849 2506 6 OpcodeCondIn[3]
rlabel m2contact 15777 2938 15777 2938 6 n_308
rlabel m2contact 15777 4978 15777 4978 6 n_6
rlabel m2contact 15729 5458 15729 5458 6 OpcodeCondIn[2]
rlabel m2contact 15729 4186 15729 4186 6 OpcodeCondIn[5]
rlabel m2contact 15705 3346 15705 3346 6 n_303
rlabel m2contact 15705 4282 15705 4282 6 OpcodeCondIn[6]
rlabel m2contact 15633 5986 15633 5986 6 n_25
rlabel m2contact 15585 3034 15585 3034 6 OpcodeCondIn[4]
rlabel m2contact 15561 5026 15561 5026 6 StatusReg[3]
rlabel m2contact 15537 3634 15537 3634 6 Rs1Sel[0]
rlabel m2contact 15513 5554 15513 5554 6 n_398
rlabel m2contact 15513 5362 15513 5362 6 n_346
rlabel m2contact 15465 6874 15465 6874 6 n_172
rlabel m2contact 15441 6106 15441 6106 6 n_314
rlabel m2contact 15321 3778 15321 3778 6 n_258
rlabel m2contact 15249 4402 15249 4402 6 n_266
rlabel m2contact 15225 1882 15225 1882 6 n_225
rlabel m2contact 15177 5554 15177 5554 6 n_28
rlabel m2contact 15177 2074 15177 2074 6 n_28
rlabel m2contact 15153 3658 15153 3658 6 n_90
rlabel m2contact 15153 5626 15153 5626 6 n_358
rlabel m2contact 15129 3754 15129 3754 6 n_234
rlabel m2contact 15105 3658 15105 3658 6 n_189
rlabel m2contact 15105 2170 15105 2170 6 n_189
rlabel m2contact 15081 6658 15081 6658 6 n_97
rlabel m2contact 15081 1594 15081 1594 6 n_97
rlabel m2contact 15057 6754 15057 6754 6 n_150
rlabel m2contact 15057 2122 15057 2122 6 n_150
rlabel m2contact 15033 5578 15033 5578 6 n_165
rlabel m2contact 15033 3154 15033 3154 6 n_268
rlabel m2contact 15009 5098 15009 5098 6 n_108
rlabel m2contact 14985 2074 14985 2074 6 n_28
rlabel m2contact 14985 2890 14985 2890 6 n_164
rlabel m2contact 14961 2434 14961 2434 6 n_20
rlabel m2contact 14937 5098 14937 5098 6 ImmSel
rlabel m2contact 14913 5098 14913 5098 6 ImmSel
rlabel m2contact 14889 6706 14889 6706 6 n_30
rlabel m2contact 14889 2938 14889 2938 6 n_30
rlabel m2contact 14865 5098 14865 5098 6 n_237
rlabel m2contact 14865 3634 14865 3634 6 n_341
rlabel m2contact 14841 6082 14841 6082 6 n_257
rlabel m2contact 14841 3058 14841 3058 6 n_371
rlabel m2contact 14817 4858 14817 4858 6 n_260
rlabel m2contact 14793 5890 14793 5890 6 n_222
rlabel m2contact 14769 5578 14769 5578 6 n_190
rlabel m2contact 14745 2194 14745 2194 6 n_243
rlabel m2contact 14745 3394 14745 3394 6 n_188
rlabel m2contact 14721 3658 14721 3658 6 n_189
rlabel m2contact 14721 3490 14721 3490 6 n_229
rlabel m2contact 14697 5626 14697 5626 6 IrWe
rlabel m2contact 14697 1570 14697 1570 6 IrWe
rlabel m2contact 14697 6898 14697 6898 6 n_29
rlabel m2contact 14697 5794 14697 5794 6 n_29
rlabel m2contact 14673 1570 14673 1570 6 IrWe
rlabel m2contact 14673 2074 14673 2074 6 n_292
rlabel m2contact 14649 6826 14649 6826 6 SysBus[2]
rlabel m2contact 14625 2002 14625 2002 6 n_197
rlabel m2contact 14625 5482 14625 5482 6 n_293
rlabel m2contact 14601 3706 14601 3706 6 n_77
rlabel m2contact 14577 5626 14577 5626 6 IrWe
rlabel m2contact 14553 4018 14553 4018 6 n_223
rlabel m2contact 14529 1594 14529 1594 6 n_97
rlabel m2contact 14529 3346 14529 3346 6 n_298
rlabel m2contact 14505 4906 14505 4906 6 n_11
rlabel m2contact 14505 4090 14505 4090 6 n_217
rlabel m2contact 14481 5626 14481 5626 6 n_206
rlabel m2contact 14457 4906 14457 4906 6 n_105
rlabel m2contact 14457 3658 14457 3658 6 n_252
rlabel m2contact 14433 5962 14433 5962 6 n_249
rlabel m2contact 14409 6754 14409 6754 6 n_150
rlabel m2contact 14409 3706 14409 3706 6 n_251
rlabel m2contact 14385 2506 14385 2506 6 OpcodeCondIn[3]
rlabel m2contact 14361 4018 14361 4018 6 n_162
rlabel m2contact 14337 3562 14337 3562 6 n_202
rlabel m2contact 14313 6826 14313 6826 6 n_15
rlabel m2contact 14313 4162 14313 4162 6 n_340
rlabel m2contact 14289 2338 14289 2338 6 OpcodeCondIn[7]
rlabel m2contact 14265 1618 14265 1618 6 n_22
rlabel m2contact 14265 4090 14265 4090 6 n_14
rlabel m2contact 14241 3778 14241 3778 6 n_258
rlabel m2contact 14217 6706 14217 6706 6 n_30
rlabel m2contact 14217 4810 14217 4810 6 stateSub[1]
rlabel m2contact 14193 3034 14193 3034 6 OpcodeCondIn[4]
rlabel m2contact 14169 6898 14169 6898 6 n_29
rlabel m2contact 14169 6754 14169 6754 6 n_111
rlabel m2contact 14145 6706 14145 6706 6 n_66
rlabel m2contact 14121 3610 14121 3610 6 stateSub[0]
rlabel m2contact 14097 3970 14097 3970 6 n_219
rlabel m2contact 14049 2074 14049 2074 6 n_292
rlabel m2contact 14049 6418 14049 6418 6 n_102
rlabel m2contact 14013 6490 14013 6490 6 n_214
rlabel m2contact 14013 2074 14013 2074 6 n_214
rlabel m2contact 14001 6874 14001 6874 6 n_172
rlabel m2contact 14001 1642 14001 1642 6 n_331
rlabel m2contact 13977 2338 13977 2338 4 OpcodeCondIn[7]
rlabel m2contact 13953 2074 13953 2074 4 n_214
rlabel m2contact 13953 5770 13953 5770 4 n_284
rlabel m2contact 13929 3034 13929 3034 4 OpcodeCondIn[4]
rlabel m2contact 13929 4018 13929 4018 4 n_162
rlabel m2contact 13905 3490 13905 3490 4 n_229
rlabel m2contact 13905 3562 13905 3562 4 n_202
rlabel m2contact 13857 6802 13857 6802 4 n_122
rlabel m2contact 13857 3730 13857 3730 4 PcEn
rlabel m2contact 13833 6346 13833 6346 4 n_121
rlabel m2contact 13833 3946 13833 3946 4 n_88
rlabel m2contact 13809 5914 13809 5914 4 stateSub[2]
rlabel m2contact 13761 6346 13761 6346 4 n_275
rlabel m2contact 13713 3610 13713 3610 4 stateSub[0]
rlabel m2contact 13689 4138 13689 4138 4 n_269
rlabel m2contact 13641 5506 13641 5506 4 n_332
rlabel m2contact 13593 6682 13593 6682 4 n_75
rlabel m2contact 13593 1618 13593 1618 4 n_75
rlabel m2contact 13569 6394 13569 6394 4 CFlag
rlabel m2contact 13545 6610 13545 6610 4 n_58
rlabel m2contact 13545 1642 13545 1642 4 n_58
rlabel m2contact 13521 5794 13521 5794 4 n_29
rlabel m2contact 13497 2506 13497 2506 4 OpcodeCondIn[3]
rlabel m2contact 13473 2338 13473 2338 4 OpcodeCondIn[7]
rlabel m2contact 13449 4690 13449 4690 4 OpcodeCondIn[1]
rlabel m2contact 13425 1618 13425 1618 4 n_75
rlabel m2contact 13425 2074 13425 2074 4 n_300
rlabel m2contact 13401 4786 13401 4786 4 n_299
rlabel m2contact 13401 2338 13401 2338 4 OpcodeCondIn[7]
rlabel m2contact 13377 3946 13377 3946 4 n_239
rlabel m2contact 13353 1642 13353 1642 4 n_58
rlabel m2contact 13353 4786 13353 4786 4 n_201
rlabel m2contact 13329 3730 13329 3730 4 n_187
rlabel m2contact 13305 3778 13305 3778 4 n_258
rlabel m2contact 13281 4714 13281 4714 4 n_63
rlabel m2contact 13257 3466 13257 3466 4 n_241
rlabel m2contact 13209 4642 13209 4642 4 n_68
rlabel m2contact 13209 4498 13209 4498 4 n_245
rlabel m2contact 13185 6586 13185 6586 4 n_21
rlabel m2contact 13185 1642 13185 1642 4 n_21
rlabel m2contact 13161 1642 13161 1642 4 n_21
rlabel m2contact 13161 4642 13161 4642 4 n_136
rlabel m2contact 13137 5818 13137 5818 4 n_118
rlabel m2contact 13113 3730 13113 3730 4 n_187
rlabel m2contact 13113 4522 13113 4522 4 n_267
rlabel m2contact 13089 4426 13089 4426 4 n_195
rlabel m2contact 13065 5194 13065 5194 4 n_140
rlabel m2contact 13065 4594 13065 4594 4 n_186
rlabel m2contact 13041 3370 13041 3370 4 n_179
rlabel m2contact 13017 2146 13017 2146 4 n_139
rlabel m2contact 12993 3610 12993 3610 4 stateSub[0]
rlabel m2contact 12993 3754 12993 3754 4 n_234
rlabel m2contact 12969 4234 12969 4234 4 n_82
rlabel m2contact 12933 5194 12933 5194 4 n_123
rlabel m2contact 12933 1714 12933 1714 4 n_123
rlabel m2contact 12921 6394 12921 6394 4 n_27
rlabel m2contact 12897 2578 12897 2578 4 StatusReg[2]
rlabel m2contact 12873 6682 12873 6682 4 n_75
rlabel m2contact 12873 5674 12873 5674 4 n_309
rlabel m2contact 12849 5986 12849 5986 4 n_25
rlabel m2contact 12849 1642 12849 1642 4 n_25
rlabel m2contact 12825 2602 12825 2602 4 n_26
rlabel m2contact 12825 2986 12825 2986 4 n_322
rlabel m2contact 12801 5194 12801 5194 4 n_123
rlabel m2contact 12801 4186 12801 4186 4 OpcodeCondIn[5]
rlabel m2contact 12777 2650 12777 2650 4 n_133
rlabel m2contact 12753 1642 12753 1642 4 n_25
rlabel m2contact 12753 3274 12753 3274 4 state[1]
rlabel m2contact 12729 5194 12729 5194 4 n_397
rlabel m2contact 12729 2602 12729 2602 4 n_397
rlabel m2contact 12705 6850 12705 6850 4 n_54
rlabel m2contact 12705 6802 12705 6802 4 n_4
rlabel m2contact 12681 5194 12681 5194 4 n_397
rlabel m2contact 12681 4810 12681 4810 4 stateSub[1]
rlabel m2contact 12657 5026 12657 5026 4 StatusReg[3]
rlabel m2contact 12657 3610 12657 3610 4 stateSub[0]
rlabel m2contact 12633 6250 12633 6250 4 n_19
rlabel m2contact 12633 4234 12633 4234 4 n_19
rlabel m2contact 12609 4234 12609 4234 4 n_19
rlabel m2contact 12609 4474 12609 4474 4 n_159
rlabel m2contact 12561 2506 12561 2506 4 OpcodeCondIn[3]
rlabel m2contact 12561 4282 12561 4282 4 OpcodeCondIn[6]
rlabel m2contact 12537 4402 12537 4402 4 n_266
rlabel m2contact 12537 4282 12537 4282 4 OpcodeCondIn[6]
rlabel m2contact 12489 5026 12489 5026 4 n_49
rlabel m2contact 12465 4282 12465 4282 4 OpcodeCondIn[6]
rlabel m2contact 12465 3730 12465 3730 4 n_271
rlabel m2contact 12441 6826 12441 6826 4 n_15
rlabel m2contact 12441 5794 12441 5794 4 n_100
rlabel m2contact 12369 4234 12369 4234 4 n_126
rlabel m2contact 12345 6010 12345 6010 4 n_40
rlabel m2contact 12321 2146 12321 2146 4 n_139
rlabel m2contact 12321 4474 12321 4474 4 n_159
rlabel m2contact 12273 2026 12273 2026 4 n_36
rlabel m2contact 12273 6106 12273 6106 4 n_314
rlabel m2contact 12249 5914 12249 5914 4 stateSub[2]
rlabel m2contact 12249 3562 12249 3562 4 n_202
rlabel m2contact 12225 6802 12225 6802 4 n_4
rlabel m2contact 12225 5266 12225 5266 4 n_65
rlabel m2contact 12177 6778 12177 6778 4 RwSel[0]
rlabel m2contact 12177 5194 12177 5194 4 SysBus[0]
rlabel m2contact 12153 4810 12153 4810 4 stateSub[1]
rlabel m2contact 12129 3418 12129 3418 4 n_301
rlabel m2contact 12105 2890 12105 2890 4 n_164
rlabel m2contact 12081 5362 12081 5362 4 n_346
rlabel m2contact 12033 5530 12033 5530 4 n_141
rlabel m2contact 12033 5362 12033 5362 4 IntStatus
rlabel m2contact 12009 3826 12009 3826 4 nWait
rlabel m2contact 11985 4522 11985 4522 4 n_267
rlabel m2contact 11961 4498 11961 4498 4 n_245
rlabel m2contact 11913 5530 11913 5530 4 n_295
rlabel m2contact 11889 5194 11889 5194 4 SysBus[0]
rlabel m2contact 11865 5482 11865 5482 4 n_293
rlabel m2contact 11817 6682 11817 6682 4 n_75
rlabel m2contact 11793 4114 11793 4114 4 OpcodeCondIn[0]
rlabel m2contact 11769 5962 11769 5962 4 n_249
rlabel m2contact 11721 2026 11721 2026 4 n_192
rlabel m2contact 11697 5770 11697 5770 4 n_284
rlabel m2contact 11673 5194 11673 5194 4 n_191
rlabel m2contact 11625 3418 11625 3418 4 n_247
rlabel m2contact 11601 5578 11601 5578 4 n_190
rlabel m2contact 11577 4594 11577 4594 4 n_186
rlabel m2contact 11529 5578 11529 5578 4 n_148
rlabel m2contact 11505 6754 11505 6754 4 n_111
rlabel m2contact 11505 1690 11505 1690 4 n_265
rlabel m2contact 11481 5554 11481 5554 4 n_28
rlabel m2contact 11433 6010 11433 6010 4 n_40
rlabel m2contact 11433 1690 11433 1690 4 n_40
rlabel m2contact 11409 1666 11409 1666 4 n_41
rlabel m2contact 11409 5962 11409 5962 4 n_249
rlabel m2contact 11385 6082 11385 6082 4 n_257
rlabel m2contact 11361 1690 11361 1690 4 n_40
rlabel m2contact 11361 5458 11361 5458 4 OpcodeCondIn[2]
rlabel m2contact 11313 6634 11313 6634 4 n_166
rlabel m2contact 11289 4186 11289 4186 4 OpcodeCondIn[5]
rlabel m2contact 11289 3874 11289 3874 4 state[0]
rlabel m2contact 11265 2914 11265 2914 4 n_254
rlabel m2contact 11265 4282 11265 4282 4 OpcodeCondIn[6]
rlabel m2contact 11217 1762 11217 1762 4 ENB
rlabel m2contact 11217 6322 11217 6322 4 n_199
rlabel m2contact 11193 2914 11193 2914 4 n_246
rlabel m2contact 11193 3562 11193 3562 4 n_202
rlabel m2contact 11169 2026 11169 2026 4 n_192
rlabel m2contact 11169 6322 11169 6322 4 n_120
rlabel m2contact 11145 6154 11145 6154 4 n_71
rlabel m2contact 11121 2290 11121 2290 4 SysBus[1]
rlabel m2contact 11097 5722 11097 5722 4 n_367
rlabel m2contact 11073 5530 11073 5530 4 n_295
rlabel m2contact 11049 2338 11049 2338 4 OpcodeCondIn[7]
rlabel m2contact 11049 5722 11049 5722 4 n_311
rlabel m2contact 11025 2794 11025 2794 4 n_113
rlabel m2contact 11025 5530 11025 5530 4 n_334
rlabel m2contact 10953 4546 10953 4546 4 n_169
rlabel m2contact 10929 6154 10929 6154 4 OpcodeCondIn[3]
rlabel m2contact 10929 2506 10929 2506 4 OpcodeCondIn[3]
rlabel m2contact 10905 6154 10905 6154 4 OpcodeCondIn[3]
rlabel m2contact 10905 2794 10905 2794 4 n_129
rlabel m2contact 10881 6634 10881 6634 4 n_176
rlabel m2contact 10881 2290 10881 2290 4 n_176
rlabel m2contact 10857 2362 10857 2362 4 n_264
rlabel m2contact 10857 6154 10857 6154 4 n_194
rlabel m2contact 10833 5602 10833 5602 4 n_193
rlabel m2contact 10833 4186 10833 4186 4 OpcodeCondIn[5]
rlabel m2contact 10809 6730 10809 6730 4 n_142
rlabel m2contact 10809 6442 10809 6442 4 n_263
rlabel m2contact 10785 5770 10785 5770 4 n_284
rlabel m2contact 10785 1762 10785 1762 4 n_284
rlabel m2contact 10761 4138 10761 4138 4 n_269
rlabel m2contact 10761 4210 10761 4210 4 n_273
rlabel m2contact 10737 6682 10737 6682 4 n_75
rlabel m2contact 10713 6634 10713 6634 4 n_176
rlabel m2contact 10713 4210 10713 4210 4 n_224
rlabel m2contact 10689 1738 10689 1738 4 n_101
rlabel m2contact 10689 2362 10689 2362 4 n_8
rlabel m2contact 10665 4138 10665 4138 4 n_46
rlabel m2contact 10629 5842 10629 5842 4 n_278
rlabel m2contact 10629 2026 10629 2026 4 n_278
rlabel m2contact 10617 1714 10617 1714 4 n_123
rlabel m2contact 10617 6634 10617 6634 4 n_115
rlabel m2contact 10593 2266 10593 2266 4 n_78
rlabel m2contact 10593 3586 10593 3586 4 n_114
rlabel m2contact 10569 5122 10569 5122 4 n_72
rlabel m2contact 10545 3946 10545 3946 4 n_239
rlabel m2contact 10521 4186 10521 4186 4 OpcodeCondIn[5]
rlabel m2contact 10497 6682 10497 6682 4 n_326
rlabel m2contact 10497 4954 10497 4954 4 n_240
rlabel m2contact 10473 6562 10473 6562 4 n_232
rlabel m2contact 10449 5122 10449 5122 4 n_325
rlabel m2contact 10425 1738 10425 1738 4 n_101
rlabel m2contact 10413 5458 10413 5458 4 OpcodeCondIn[2]
rlabel m2contact 10413 3946 10413 3946 4 OpcodeCondIn[2]
rlabel m2contact 10401 6706 10401 6706 4 n_66
rlabel m2contact 10401 3874 10401 3874 4 state[0]
rlabel m2contact 10377 1762 10377 1762 4 n_284
rlabel m2contact 10377 3562 10377 3562 4 n_202
rlabel m2contact 10353 5266 10353 5266 4 n_65
rlabel m2contact 10329 1786 10329 1786 4 n_307
rlabel m2contact 10329 2938 10329 2938 4 n_30
rlabel m2contact 10305 6082 10305 6082 4 n_257
rlabel m2contact 10281 2026 10281 2026 4 n_278
rlabel m2contact 10281 2938 10281 2938 4 n_32
rlabel m2contact 10257 4546 10257 4546 4 n_169
rlabel m2contact 10233 4978 10233 4978 4 n_6
rlabel m2contact 10209 3610 10209 3610 4 stateSub[0]
rlabel m2contact 10185 2242 10185 2242 4 n_7
rlabel m2contact 10161 2746 10161 2746 4 n_285
rlabel m2contact 10161 2866 10161 2866 4 n_106
rlabel m2contact 10137 3922 10137 3922 4 n_85
rlabel m2contact 10113 2002 10113 2002 4 n_197
rlabel m2contact 10113 3274 10113 3274 4 state[1]
rlabel m2contact 10089 3754 10089 3754 4 n_234
rlabel m2contact 10065 4762 10065 4762 4 n_211
rlabel m2contact 10041 3946 10041 3946 4 OpcodeCondIn[2]
rlabel m2contact 10041 4978 10041 4978 4 n_38
rlabel m2contact 10017 2506 10017 2506 4 OpcodeCondIn[3]
rlabel m2contact 9993 2338 9993 2338 4 OpcodeCondIn[7]
rlabel m2contact 9969 2746 9969 2746 4 n_9
rlabel m2contact 9945 4282 9945 4282 4 OpcodeCondIn[6]
rlabel m2contact 9921 3946 9921 3946 4 nWE
rlabel m2contact 9897 3922 9897 3922 4 n_297
rlabel m2contact 9873 1810 9873 1810 4 n_375
rlabel m2contact 9873 2026 9873 2026 4 n_235
rlabel m2contact 9849 2242 9849 2242 4 n_51
rlabel m2contact 9825 6682 9825 6682 4 n_326
rlabel m2contact 9801 1834 9801 1834 4 n_368
rlabel m2contact 9801 6658 9801 6658 4 n_97
rlabel m2contact 9777 2146 9777 2146 4 n_139
rlabel m2contact 9753 2266 9753 2266 4 n_78
rlabel m2contact 9753 3154 9753 3154 4 n_268
rlabel m2contact 9705 4954 9705 4954 4 n_240
rlabel m2contact 9705 4714 9705 4714 4 n_63
rlabel m2contact 9681 3754 9681 3754 4 n_234
rlabel m2contact 9657 3034 9657 3034 4 OpcodeCondIn[4]
rlabel m2contact 9633 4642 9633 4642 4 n_136
rlabel m2contact 9609 6634 9609 6634 4 n_115
rlabel m2contact 9585 1858 9585 1858 4 n_207
rlabel m2contact 9585 1882 9585 1882 4 n_225
rlabel m2contact 9561 4306 9561 4306 4 n_128
rlabel m2contact 9537 1906 9537 1906 4 n_31
rlabel m2contact 9537 2122 9537 2122 4 n_150
rlabel m2contact 9489 1930 9489 1930 4 PcSel[0]
rlabel m2contact 9489 2122 9489 2122 4 n_220
rlabel m2contact 9465 4210 9465 4210 4 n_224
rlabel m2contact 9465 4066 9465 4066 4 n_349
rlabel m2contact 9441 2170 9441 2170 4 n_189
rlabel m2contact 9393 1954 9393 1954 4 n_221
rlabel m2contact 9393 1978 9393 1978 4 n_84
rlabel m2contact 9345 6610 9345 6610 4 n_58
rlabel m2contact 9345 2338 9345 2338 4 OpcodeCondIn[7]
rlabel m2contact 9321 6586 9321 6586 4 n_21
rlabel m2contact 9321 4954 9321 4954 4 n_240
rlabel m2contact 9285 4498 9285 4498 4 n_245
rlabel m2contact 9285 1978 9285 1978 4 n_245
rlabel m2contact 9273 6514 9273 6514 4 n_233
rlabel m2contact 9249 1978 9249 1978 4 n_245
rlabel m2contact 9249 4258 9249 4258 4 n_231
rlabel m2contact 9225 2098 9225 2098 4 n_155
rlabel m2contact 9225 3490 9225 3490 4 n_229
rlabel m2contact 9201 6562 9201 6562 4 n_232
rlabel m2contact 9189 6514 9189 6514 4 n_92
rlabel m2contact 9189 2098 9189 2098 4 n_92
rlabel m2contact 9177 2026 9177 2026 4 n_235
rlabel m2contact 9153 6538 9153 6538 4 n_238
rlabel m2contact 9153 4426 9153 4426 4 n_195
rlabel m2contact 9129 2146 9129 2146 4 n_139
rlabel m2contact 9105 6514 9105 6514 4 n_92
rlabel m2contact 9105 3754 9105 3754 4 n_234
rlabel m2contact 9081 6490 9081 6490 4 n_214
rlabel m2contact 9057 2002 9057 2002 4 n_197
rlabel m2contact 9057 5770 9057 5770 4 n_284
rlabel m2contact 9057 2026 9057 2026 4 n_284
rlabel m2contact 9033 6466 9033 6466 4 n_228
rlabel m2contact 9033 4714 9033 4714 4 n_63
rlabel m2contact 9009 2026 9009 2026 4 n_284
rlabel m2contact 9009 2722 9009 2722 4 n_215
rlabel m2contact 8985 2410 8985 2410 4 n_226
rlabel m2contact 8961 3130 8961 3130 4 n_145
rlabel m2contact 8937 4210 8937 4210 4 n_224
rlabel m2contact 8913 3994 8913 3994 4 n_153
rlabel m2contact 8913 3874 8913 3874 4 state[0]
rlabel m2contact 8889 2146 8889 2146 4 n_139
rlabel m2contact 8889 3514 8889 3514 4 n_204
rlabel m2contact 8841 6442 8841 6442 4 n_263
rlabel m2contact 8793 2050 8793 2050 4 Op1Sel
rlabel m2contact 8793 3250 8793 3250 4 n_177
rlabel m2contact 8769 2074 8769 2074 4 n_300
rlabel m2contact 8769 3490 8769 3490 4 n_229
rlabel m2contact 8721 2098 8721 2098 4 n_92
rlabel m2contact 8721 6418 8721 6418 4 n_102
rlabel m2contact 8697 4690 8697 4690 4 OpcodeCondIn[1]
rlabel m2contact 8673 6394 8673 6394 4 n_27
rlabel m2contact 8673 2506 8673 2506 4 OpcodeCondIn[3]
rlabel m2contact 8625 4450 8625 4450 4 n_99
rlabel m2contact 8601 5770 8601 5770 4 n_284
rlabel m2contact 8577 3154 8577 3154 4 n_268
rlabel m2contact 8529 6370 8529 6370 4 n_312
rlabel m2contact 8481 6346 8481 6346 4 n_275
rlabel m2contact 8481 2506 8481 2506 4 OpcodeCondIn[3]
rlabel m2contact 8457 5890 8457 5890 4 n_222
rlabel m2contact 8457 4186 8457 4186 4 OpcodeCondIn[5]
rlabel m2contact 8409 6322 8409 6322 4 n_120
rlabel m2contact 8409 5890 8409 5890 4 n_313
rlabel m2contact 8385 6250 8385 6250 4 n_19
rlabel m2contact 8361 2122 8361 2122 4 n_220
rlabel m2contact 8361 3970 8361 3970 4 n_219
rlabel m2contact 8337 4522 8337 4522 4 n_267
rlabel m2contact 8313 5122 8313 5122 4 n_325
rlabel m2contact 8289 3154 8289 3154 4 n_268
rlabel m2contact 8265 5890 8265 5890 4 n_313
rlabel m2contact 8265 3754 8265 3754 4 n_234
rlabel m2contact 8241 2146 8241 2146 4 n_139
rlabel m2contact 8217 6298 8217 6298 4 n_250
rlabel m2contact 8217 6250 8217 6250 4 n_243
rlabel m2contact 8217 2194 8217 2194 4 n_243
rlabel m2contact 8193 2170 8193 2170 4 n_189
rlabel m2contact 8193 3826 8193 3826 4 nWait
rlabel m2contact 8169 6274 8169 6274 4 n_157
rlabel m2contact 8169 2506 8169 2506 4 OpcodeCondIn[3]
rlabel m2contact 8145 6250 8145 6250 4 n_243
rlabel m2contact 8145 4474 8145 4474 4 n_159
rlabel m2contact 8121 5962 8121 5962 4 n_249
rlabel m2contact 8097 6226 8097 6226 4 n_324
rlabel m2contact 8073 4498 8073 4498 4 n_245
rlabel m2contact 8049 4090 8049 4090 4 n_14
rlabel m2contact 8001 4690 8001 4690 4 OpcodeCondIn[1]
rlabel m2contact 7977 2194 7977 2194 4 n_243
rlabel m2contact 7953 6202 7953 6202 4 n_315
rlabel m2contact 7953 4522 7953 4522 4 n_267
rlabel m2contact 7929 6178 7929 6178 4 n_60
rlabel m2contact 7929 3610 7929 3610 4 stateSub[0]
rlabel m2contact 7905 6154 7905 6154 4 n_194
rlabel m2contact 7881 6130 7881 6130 4 n_255
rlabel m2contact 7881 3226 7881 3226 4 n_377
rlabel m2contact 7857 6106 7857 6106 4 n_314
rlabel m2contact 7857 4714 7857 4714 4 n_63
rlabel m2contact 7833 5818 7833 5818 4 n_118
rlabel m2contact 7809 2218 7809 2218 4 n_259
rlabel m2contact 7785 6082 7785 6082 4 n_257
rlabel m2contact 7761 2314 7761 2314 4 n_59
rlabel m2contact 7761 3874 7761 3874 4 state[0]
rlabel m2contact 7737 3778 7737 3778 4 n_258
rlabel m2contact 7713 6058 7713 6058 4 n_161
rlabel m2contact 7713 3874 7713 3874 4 state[0]
rlabel m2contact 7665 4138 7665 4138 4 n_46
rlabel m2contact 7641 5458 7641 5458 4 OpcodeCondIn[2]
rlabel m2contact 7617 6034 7617 6034 4 n_399
rlabel m2contact 7617 4282 7617 4282 4 OpcodeCondIn[6]
rlabel m2contact 7593 4138 7593 4138 4 n_45
rlabel m2contact 7593 3754 7593 3754 4 n_234
rlabel m2contact 7569 4114 7569 4114 4 OpcodeCondIn[0]
rlabel m2contact 7545 6010 7545 6010 4 n_40
rlabel m2contact 7521 2242 7521 2242 4 n_51
rlabel m2contact 7521 5986 7521 5986 4 n_25
rlabel m2contact 7521 4834 7521 4834 4 n_33
rlabel m2contact 7521 2314 7521 2314 4 n_33
rlabel m2contact 7497 2314 7497 2314 4 n_33
rlabel m2contact 7497 3562 7497 3562 4 n_202
rlabel m2contact 7473 2266 7473 2266 4 n_78
rlabel m2contact 7449 4546 7449 4546 4 n_169
rlabel m2contact 7449 2314 7449 2314 4 n_169
rlabel m2contact 7425 2290 7425 2290 4 n_176
rlabel m2contact 7425 3226 7425 3226 4 n_377
rlabel m2contact 7401 3322 7401 3322 4 n_288
rlabel m2contact 7377 2986 7377 2986 4 n_322
rlabel m2contact 7353 3322 7353 3322 4 n_135
rlabel m2contact 7329 3226 7329 3226 4 n_151
rlabel m2contact 7305 5002 7305 5002 4 n_70
rlabel m2contact 7281 5962 7281 5962 4 n_249
rlabel m2contact 7281 2338 7281 2338 4 OpcodeCondIn[7]
rlabel m2contact 7257 2314 7257 2314 4 n_169
rlabel m2contact 7257 4138 7257 4138 4 n_45
rlabel m2contact 7209 5938 7209 5938 4 n_163
rlabel m2contact 7185 2338 7185 2338 4 OpcodeCondIn[7]
rlabel m2contact 7185 5794 7185 5794 4 n_100
rlabel m2contact 7161 4810 7161 4810 4 stateSub[1]
rlabel m2contact 7137 4450 7137 4450 4 n_99
rlabel m2contact 7137 4018 7137 4018 4 n_162
rlabel m2contact 7101 5698 7101 5698 4 StatusReg[0]
rlabel m2contact 7101 4450 7101 4450 4 StatusReg[0]
rlabel m2contact 7089 5794 7089 5794 4 n_12
rlabel m2contact 7065 3586 7065 3586 4 n_114
rlabel m2contact 7041 5914 7041 5914 4 stateSub[2]
rlabel m2contact 7041 4306 7041 4306 4 n_128
rlabel m2contact 7017 5818 7017 5818 4 n_118
rlabel m2contact 6993 2698 6993 2698 4 n_212
rlabel m2contact 6969 2362 6969 2362 4 n_8
rlabel m2contact 6969 4474 6969 4474 4 n_159
rlabel m2contact 6945 4522 6945 4522 4 n_267
rlabel m2contact 6945 4114 6945 4114 4 OpcodeCondIn[0]
rlabel m2contact 6921 4450 6921 4450 4 StatusReg[0]
rlabel m2contact 6921 4498 6921 4498 4 n_245
rlabel m2contact 6897 4690 6897 4690 4 OpcodeCondIn[1]
rlabel m2contact 6873 4450 6873 4450 4 n_316
rlabel m2contact 6849 2386 6849 2386 4 n_227
rlabel m2contact 6849 3610 6849 3610 4 stateSub[0]
rlabel m2contact 6825 5890 6825 5890 4 n_313
rlabel m2contact 6825 4762 6825 4762 4 n_211
rlabel m2contact 6801 2410 6801 2410 4 n_226
rlabel m2contact 6777 4042 6777 4042 4 n_354
rlabel m2contact 6753 3226 6753 3226 4 n_151
rlabel m2contact 6729 3034 6729 3034 4 OpcodeCondIn[4]
rlabel m2contact 6729 5434 6729 5434 4 n_319
rlabel m2contact 6705 3562 6705 3562 4 n_202
rlabel m2contact 6681 5338 6681 5338 4 n_400
rlabel m2contact 6681 3250 6681 3250 4 n_177
rlabel m2contact 6657 5866 6657 5866 4 n_43
rlabel m2contact 6657 4282 6657 4282 4 OpcodeCondIn[6]
rlabel m2contact 6633 5050 6633 5050 4 n_79
rlabel m2contact 6609 2434 6609 2434 4 n_20
rlabel m2contact 6609 5842 6609 5842 4 n_278
rlabel m2contact 6585 4282 6585 4282 4 OpcodeCondIn[6]
rlabel m2contact 6561 5818 6561 5818 4 n_118
rlabel m2contact 6561 3754 6561 3754 4 n_234
rlabel m2contact 6537 4690 6537 4690 4 OpcodeCondIn[1]
rlabel m2contact 6513 3754 6513 3754 4 n_234
rlabel m2contact 6489 2458 6489 2458 4 n_280
rlabel m2contact 6489 3586 6489 3586 4 n_114
rlabel m2contact 6465 5794 6465 5794 4 n_12
rlabel m2contact 6441 5746 6441 5746 4 n_261
rlabel m2contact 6417 3970 6417 3970 4 n_219
rlabel m2contact 6393 4858 6393 4858 4 n_260
rlabel m2contact 6345 2482 6345 2482 4 n_134
rlabel m2contact 6321 2506 6321 2506 4 OpcodeCondIn[3]
rlabel m2contact 6321 5770 6321 5770 4 n_284
rlabel m2contact 6321 5746 6321 5746 4 n_133
rlabel m2contact 6321 2650 6321 2650 4 n_133
rlabel m2contact 6297 5746 6297 5746 4 n_133
rlabel m2contact 6297 3490 6297 3490 4 n_229
rlabel m2contact 6273 3370 6273 3370 4 n_179
rlabel m2contact 6249 5722 6249 5722 4 n_311
rlabel m2contact 6225 5698 6225 5698 4 StatusReg[0]
rlabel m2contact 6201 5674 6201 5674 4 n_309
rlabel m2contact 6177 5650 6177 5650 4 n_116
rlabel m2contact 6153 2530 6153 2530 4 n_276
rlabel m2contact 6153 5602 6153 5602 4 n_193
rlabel m2contact 6105 2554 6105 2554 4 n_73
rlabel m2contact 6105 2626 6105 2626 4 IRQ2
rlabel m2contact 6081 5362 6081 5362 4 IntStatus
rlabel m2contact 6081 4282 6081 4282 4 OpcodeCondIn[6]
rlabel m2contact 6033 3034 6033 3034 4 OpcodeCondIn[4]
rlabel m2contact 6033 5194 6033 5194 4 n_191
rlabel m2contact 5985 3394 5985 3394 4 n_188
rlabel m2contact 5985 2626 5985 2626 4 Flags[0]
rlabel m2contact 5961 5362 5961 5362 4 n_74
rlabel m2contact 5889 3034 5889 3034 4 n_361
rlabel m2contact 5841 2578 5841 2578 4 StatusReg[2]
rlabel m2contact 5841 3394 5841 3394 4 n_345
rlabel m2contact 5793 2602 5793 2602 4 n_397
rlabel m2contact 5793 5626 5793 5626 4 n_206
rlabel m2contact 5769 5602 5769 5602 4 n_193
rlabel m2contact 5745 5578 5745 5578 4 n_148
rlabel m2contact 5721 3874 5721 3874 4 state[0]
rlabel m2contact 5697 4810 5697 4810 4 stateSub[1]
rlabel m2contact 5649 5554 5649 5554 4 n_28
rlabel m2contact 5625 3610 5625 3610 4 stateSub[0]
rlabel m2contact 5601 3754 5601 3754 4 n_234
rlabel m2contact 5553 5530 5553 5530 4 n_334
rlabel m2contact 5529 2626 5529 2626 4 Flags[0]
rlabel m2contact 5505 5506 5505 5506 4 n_332
rlabel m2contact 5457 5482 5457 5482 4 n_293
rlabel m2contact 5409 5458 5409 5458 4 OpcodeCondIn[2]
rlabel m2contact 5385 3706 5385 3706 4 n_251
rlabel m2contact 5313 5434 5313 5434 4 n_319
rlabel m2contact 5313 4066 5313 4066 4 n_349
rlabel m2contact 5265 2650 5265 2650 4 n_133
rlabel m2contact 5265 5338 5265 5338 4 n_400
rlabel m2contact 5217 2674 5217 2674 4 WdSel
rlabel m2contact 5217 4882 5217 4882 4 n_81
rlabel m2contact 5193 4714 5193 4714 4 n_63
rlabel m2contact 5169 2722 5169 2722 4 n_215
rlabel m2contact 5169 3154 5169 3154 4 n_268
rlabel m2contact 5145 2698 5145 2698 4 n_212
rlabel m2contact 5133 5338 5133 5338 4 n_95
rlabel m2contact 5133 2722 5133 2722 4 n_95
rlabel m2contact 5121 5362 5121 5362 4 n_74
rlabel m2contact 5097 3994 5097 3994 4 n_153
rlabel m2contact 5073 2722 5073 2722 4 n_95
rlabel m2contact 5073 4498 5073 4498 4 n_245
rlabel m2contact 5025 5410 5025 5410 4 n_182
rlabel m2contact 5001 2746 5001 2746 4 n_9
rlabel m2contact 5001 5386 5001 5386 4 n_93
rlabel m2contact 5001 5362 5001 5362 4 n_229
rlabel m2contact 5001 3490 5001 3490 4 n_229
rlabel m2contact 4977 5362 4977 5362 4 n_229
rlabel m2contact 4977 4282 4977 4282 4 OpcodeCondIn[6]
rlabel m2contact 4953 3754 4953 3754 4 n_234
rlabel m2contact 4905 5338 4905 5338 4 n_95
rlabel m2contact 4905 3994 4905 3994 4 n_153
rlabel m2contact 4857 5314 4857 5314 4 n_94
rlabel m2contact 4857 4690 4857 4690 4 OpcodeCondIn[1]
rlabel m2contact 4833 4114 4833 4114 4 OpcodeCondIn[0]
rlabel m2contact 4809 5290 4809 5290 4 n_53
rlabel m2contact 4785 5266 4785 5266 4 n_65
rlabel m2contact 4761 2770 4761 2770 4 n_10
rlabel m2contact 4737 5242 4737 5242 4 n_130
rlabel m2contact 4713 5218 4713 5218 4 n_152
rlabel m2contact 4689 3514 4689 3514 4 n_204
rlabel m2contact 4665 3226 4665 3226 4 n_151
rlabel m2contact 4665 3058 4665 3058 4 n_371
rlabel m2contact 4617 3706 4617 3706 4 n_251
rlabel m2contact 4593 3226 4593 3226 4 n_262
rlabel m2contact 4569 4522 4569 4522 4 n_267
rlabel m2contact 4545 5194 4545 5194 4 n_191
rlabel m2contact 4545 3706 4545 3706 4 ALE
rlabel m2contact 4521 5170 4521 5170 4 n_196
rlabel m2contact 4497 2794 4497 2794 4 n_129
rlabel m2contact 4473 4306 4473 4306 4 n_128
rlabel m2contact 4449 2818 4449 2818 4 n_87
rlabel m2contact 4425 5146 4425 5146 4 n_17
rlabel m2contact 4377 5122 4377 5122 4 n_325
rlabel m2contact 4353 3082 4353 3082 4 n_373
rlabel m2contact 4329 5098 4329 5098 4 n_237
rlabel m2contact 4329 4114 4329 4114 4 OpcodeCondIn[0]
rlabel m2contact 4305 4690 4305 4690 4 OpcodeCondIn[1]
rlabel m2contact 4281 5074 4281 5074 4 n_13
rlabel m2contact 4257 4738 4257 4738 4 n_200
rlabel m2contact 4233 4546 4233 4546 4 n_169
rlabel m2contact 4209 2842 4209 2842 4 n_144
rlabel m2contact 4209 3610 4209 3610 4 stateSub[0]
rlabel m2contact 4185 3874 4185 3874 4 state[0]
rlabel m2contact 4137 5050 4137 5050 4 n_79
rlabel m2contact 4113 5026 4113 5026 4 n_49
rlabel m2contact 4089 2866 4089 2866 4 n_106
rlabel m2contact 4089 5002 4089 5002 4 n_70
rlabel m2contact 4041 2890 4041 2890 4 n_164
rlabel m2contact 4041 2914 4041 2914 4 n_246
rlabel m2contact 4017 4498 4017 4498 4 n_245
rlabel m2contact 3993 2938 3993 2938 4 n_32
rlabel m2contact 3993 4930 3993 4930 4 n_198
rlabel m2contact 3969 4978 3969 4978 4 n_38
rlabel m2contact 3945 4930 3945 4930 4 AluEn
rlabel m2contact 3921 2962 3921 2962 4 Rs1Sel[1]
rlabel m2contact 3897 2986 3897 2986 4 n_322
rlabel m2contact 3897 3010 3897 3010 4 n_242
rlabel m2contact 3873 3034 3873 3034 4 n_361
rlabel m2contact 3873 3250 3873 3250 4 n_177
rlabel m2contact 3849 4954 3849 4954 4 n_240
rlabel m2contact 3849 3082 3849 3082 4 n_373
rlabel m2contact 3825 3466 3825 3466 4 n_241
rlabel m2contact 3801 4930 3801 4930 4 AluEn
rlabel m2contact 3777 3058 3777 3058 4 n_371
rlabel m2contact 3777 4906 3777 4906 4 n_105
rlabel m2contact 3753 3274 3753 3274 4 state[1]
rlabel m2contact 3729 3082 3729 3082 4 n_373
rlabel m2contact 3729 4882 3729 4882 4 n_81
rlabel m2contact 3657 3106 3657 3106 4 n_184
rlabel m2contact 3633 3130 3633 3130 4 n_145
rlabel m2contact 3609 3154 3609 3154 4 n_268
rlabel m2contact 3609 3178 3609 3178 4 n_339
rlabel m2contact 3561 3202 3561 3202 4 n_39
rlabel m2contact 3561 3226 3561 3226 4 n_262
rlabel m2contact 3537 3250 3537 3250 4 n_177
rlabel m2contact 3537 3994 3537 3994 4 n_153
rlabel m2contact 3513 4858 3513 4858 4 n_260
rlabel m2contact 3465 4834 3465 4834 4 n_33
rlabel m2contact 3441 4810 3441 4810 4 stateSub[1]
rlabel m2contact 3417 3274 3417 3274 4 state[1]
rlabel m2contact 3369 3274 3369 3274 4 state[1]
rlabel m2contact 3369 4786 3369 4786 4 n_201
rlabel m2contact 3345 4762 3345 4762 4 n_211
rlabel m2contact 3321 4738 3321 4738 4 n_200
rlabel m2contact 3321 3778 3321 3778 4 n_258
rlabel m2contact 3297 3754 3297 3754 4 n_234
rlabel m2contact 3273 3778 3273 3778 4 n_258
rlabel m2contact 3225 3298 3225 3298 4 n_16
rlabel m2contact 3177 3778 3177 3778 4 n_258
rlabel m2contact 3153 4714 3153 4714 4 n_63
rlabel m2contact 3105 3322 3105 3322 4 n_135
rlabel m2contact 3057 4690 3057 4690 4 OpcodeCondIn[1]
rlabel m2contact 3033 4666 3033 4666 4 n_110
rlabel m2contact 2961 3346 2961 3346 4 n_298
rlabel m2contact 2961 3490 2961 3490 4 n_229
rlabel m2contact 2913 4642 2913 4642 4 n_136
rlabel m2contact 2865 4618 2865 4618 4 n_154
rlabel m2contact 2841 3514 2841 3514 4 n_204
rlabel m2contact 2817 3370 2817 3370 4 n_179
rlabel m2contact 2817 4594 2817 4594 4 n_186
rlabel m2contact 2793 3490 2793 3490 4 n_229
rlabel m2contact 2769 4570 2769 4570 4 n_160
rlabel m2contact 2745 3394 2745 3394 4 n_345
rlabel m2contact 2745 4546 2745 4546 4 n_169
rlabel m2contact 2721 4522 2721 4522 4 n_267
rlabel m2contact 2697 4498 2697 4498 4 n_245
rlabel m2contact 2673 3418 2673 3418 4 n_247
rlabel m2contact 2673 4474 2673 4474 4 n_159
rlabel m2contact 2649 4450 2649 4450 4 n_316
rlabel m2contact 2625 4426 2625 4426 4 n_195
rlabel m2contact 2601 3442 2601 3442 4 n_205
rlabel m2contact 2601 4402 2601 4402 4 n_266
rlabel m2contact 2577 3466 2577 3466 4 n_241
rlabel m2contact 2577 4378 2577 4378 4 n_119
rlabel m2contact 2553 3490 2553 3490 4 n_229
rlabel m2contact 2529 3514 2529 3514 4 n_204
rlabel m2contact 2529 4354 2529 4354 4 n_256
rlabel m2contact 2505 4330 2505 4330 4 n_174
rlabel m2contact 2481 3538 2481 3538 4 n_158
rlabel m2contact 2457 3562 2457 3562 4 n_202
rlabel m2contact 2433 4306 2433 4306 4 n_128
rlabel m2contact 2409 4186 2409 4186 4 OpcodeCondIn[5]
rlabel m2contact 2385 4282 2385 4282 4 OpcodeCondIn[6]
rlabel m2contact 2361 4258 2361 4258 4 n_231
rlabel m2contact 2313 3730 2313 3730 4 n_271
rlabel m2contact 2289 4234 2289 4234 4 n_126
rlabel m2contact 2265 3586 2265 3586 4 n_114
rlabel m2contact 2265 4210 2265 4210 4 n_224
rlabel m2contact 2217 3610 2217 3610 4 stateSub[0]
rlabel m2contact 2217 3634 2217 3634 4 n_341
rlabel m2contact 2193 4186 2193 4186 4 OpcodeCondIn[5]
rlabel m2contact 2169 4162 2169 4162 4 n_340
rlabel m2contact 2121 4138 2121 4138 4 n_45
rlabel m2contact 2073 4114 2073 4114 4 OpcodeCondIn[0]
rlabel m2contact 2049 4090 2049 4090 4 n_14
rlabel m2contact 1977 4066 1977 4066 4 n_349
rlabel m2contact 1953 4042 1953 4042 4 n_354
rlabel m2contact 1929 3658 1929 3658 4 n_252
rlabel m2contact 1881 4018 1881 4018 4 n_162
rlabel m2contact 1833 3994 1833 3994 4 n_153
rlabel m2contact 1809 3970 1809 3970 4 n_219
rlabel m2contact 1761 3682 1761 3682 4 nME
rlabel m2contact 1737 3946 1737 3946 4 nWE
rlabel m2contact 1713 3706 1713 3706 4 ALE
rlabel m2contact 1689 3922 1689 3922 4 n_297
rlabel m2contact 1665 3898 1665 3898 4 n_370
rlabel m2contact 1665 3730 1665 3730 4 n_271
rlabel m2contact 1641 3754 1641 3754 4 n_234
rlabel m2contact 1641 3874 1641 3874 4 state[0]
rlabel m2contact 1617 3778 1617 3778 4 n_258
rlabel m2contact 1617 3850 1617 3850 4 n_357
rlabel m2contact 26793 377 26793 377 8 CFlag
rlabel m2contact 26793 17 26793 17 8 CFlag
rlabel m2contact 26793 425 26793 425 8 Flags[2]
rlabel m2contact 26745 401 26745 401 8 Flags[1]
rlabel m2contact 26697 209 26697 209 8 n_210
rlabel m2contact 26649 689 26649 689 8 n_168
rlabel m2contact 26577 377 26577 377 8 CFlag
rlabel m2contact 26025 593 26025 593 8 n_337
rlabel m2contact 25905 617 25905 617 8 n_56
rlabel m2contact 25809 665 25809 665 8 n_277
rlabel m2contact 25209 113 25209 113 8 n_379
rlabel m2contact 25089 329 25089 329 8 n_317
rlabel m2contact 25017 569 25017 569 8 n_290
rlabel m2contact 24993 401 24993 401 8 n_291
rlabel m2contact 24993 353 24993 353 8 n_291
rlabel m2contact 24969 401 24969 401 8 n_291
rlabel metal2 24963 377 24963 377 8 SysBus[3]
rlabel m2contact 24945 377 24945 377 8 SysBus[3]
rlabel m2contact 24873 233 24873 233 8 n_124
rlabel m2contact 24777 401 24777 401 8 n_175
rlabel m2contact 24681 281 24681 281 8 n_50
rlabel m2contact 24273 497 24273 497 8 n_270
rlabel m2contact 23985 377 23985 377 8 n_305
rlabel m2contact 23745 641 23745 641 8 n_117
rlabel m2contact 23697 425 23697 425 8 n_104
rlabel m2contact 23553 257 23553 257 8 n_42
rlabel m2contact 23289 137 23289 137 8 n_143
rlabel m2contact 23097 161 23097 161 8 n_1
rlabel m2contact 23049 65 23049 65 8 nIRQ
rlabel m2contact 22953 401 22953 401 8 n_175
rlabel m2contact 22929 713 22929 713 8 n_125
rlabel m2contact 22833 185 22833 185 8 n_24
rlabel m2contact 22641 185 22641 185 8 n_24
rlabel m2contact 22497 401 22497 401 8 n_147
rlabel m2contact 22329 545 22329 545 8 n_344
rlabel m2contact 22281 737 22281 737 8 n_149
rlabel m2contact 22089 473 22089 473 8 n_52
rlabel m2contact 21969 17 21969 17 8 n_304
rlabel m2contact 21609 89 21609 89 8 n_57
rlabel m2contact 21537 305 21537 305 8 n_67
rlabel m2contact 21489 521 21489 521 8 n_328
rlabel m2contact 21297 449 21297 449 8 n_83
rlabel m2contact 21225 617 21225 617 8 n_56
rlabel m2contact 21009 617 21009 617 8 n_183
rlabel m2contact 20985 641 20985 641 8 n_117
rlabel m2contact 20889 305 20889 305 8 n_67
rlabel m2contact 20553 641 20553 641 8 n_281
rlabel m2contact 20145 17 20145 17 8 n_304
rlabel m2contact 20049 137 20049 137 8 n_143
rlabel m2contact 19929 281 19929 281 8 n_50
rlabel m2contact 19257 137 19257 137 8 n_156
rlabel m2contact 18993 281 18993 281 8 IRQ1
rlabel m2contact 18585 161 18585 161 8 n_1
rlabel m2contact 18345 353 18345 353 8 n_291
rlabel m2contact 18321 377 18321 377 8 n_305
rlabel m2contact 18225 353 18225 353 8 n_48
rlabel m2contact 18009 665 18009 665 8 n_277
rlabel m2contact 17985 377 17985 377 8 n_342
rlabel m2contact 17865 161 17865 161 8 n_283
rlabel m2contact 17817 497 17817 497 8 n_270
rlabel m2contact 17697 665 17697 665 8 n_287
rlabel m2contact 17529 497 17529 497 8 n_282
rlabel metal2 17451 17 17451 17 8 SysBus[2]
rlabel m2contact 17433 17 17433 17 8 SysBus[2]
rlabel m2contact 17169 737 17169 737 8 n_149
rlabel m2contact 16833 113 16833 113 8 n_379
rlabel m2contact 16233 281 16233 281 8 IRQ1
rlabel m2contact 15825 185 15825 185 8 n_24
rlabel m2contact 15489 329 15489 329 8 n_317
rlabel m2contact 15393 689 15393 689 8 n_168
rlabel m2contact 15345 281 15345 281 8 n_131
rlabel m2contact 15273 665 15273 665 8 n_287
rlabel m2contact 15201 401 15201 401 8 n_147
rlabel m2contact 15105 473 15105 473 8 n_52
rlabel m2contact 14913 473 14913 473 8 n_244
rlabel m2contact 14889 545 14889 545 8 n_344
rlabel m2contact 14361 377 14361 377 8 n_342
rlabel m2contact 14073 329 14073 329 8 n_359
rlabel m2contact 14025 689 14025 689 8 n_306
rlabel m2contact 13809 545 13809 545 2 n_327
rlabel m2contact 13785 377 13785 377 2 n_302
rlabel m2contact 13761 665 13761 665 2 n_272
rlabel m2contact 13689 545 13689 545 2 n_327
rlabel m2contact 13593 545 13593 545 2 n_109
rlabel m2contact 13545 113 13545 113 2 n_61
rlabel m2contact 13521 89 13521 89 2 n_57
rlabel m2contact 13473 89 13473 89 2 n_76
rlabel m2contact 13017 713 13017 713 2 n_125
rlabel m2contact 12921 689 12921 689 2 n_306
rlabel m2contact 12777 185 12777 185 2 n_24
rlabel m2contact 12489 665 12489 665 2 n_272
rlabel m2contact 12393 113 12393 113 2 n_61
rlabel m2contact 12177 113 12177 113 2 SysBus[0]
rlabel m2contact 11457 641 11457 641 2 n_281
rlabel m2contact 11313 161 11313 161 2 n_283
rlabel metal2 11139 161 11139 161 2 SysBus[1]
rlabel m2contact 11121 161 11121 161 2 SysBus[1]
rlabel m2contact 11073 161 11073 161 2 n_137
rlabel m2contact 10977 617 10977 617 2 n_183
rlabel m2contact 10929 161 10929 161 2 n_137
rlabel m2contact 10641 161 10641 161 2 n_37
rlabel m2contact 10209 593 10209 593 2 n_337
rlabel m2contact 9969 353 9969 353 2 n_48
rlabel m2contact 9921 353 9921 353 2 n_47
rlabel m2contact 9633 569 9633 569 2 n_290
rlabel m2contact 9561 545 9561 545 2 n_109
rlabel m2contact 9441 521 9441 521 2 n_328
rlabel m2contact 9273 137 9273 137 2 n_156
rlabel m2contact 8841 137 8841 137 2 n_353
rlabel m2contact 8649 257 8649 257 2 n_42
rlabel m2contact 8577 353 8577 353 2 n_47
rlabel m2contact 8289 257 8289 257 2 n_62
rlabel m2contact 8049 497 8049 497 2 n_282
rlabel m2contact 8001 473 8001 473 2 n_244
rlabel m2contact 7953 113 7953 113 2 SysBus[0]
rlabel m2contact 7809 305 7809 305 2 n_67
rlabel m2contact 7689 305 7689 305 2 n_67
rlabel m2contact 7641 113 7641 113 2 n_18
rlabel m2contact 7377 449 7377 449 2 n_83
rlabel m2contact 7089 425 7089 425 2 n_104
rlabel m2contact 6753 401 6753 401 2 n_147
rlabel m2contact 6441 209 6441 209 2 n_210
rlabel m2contact 6417 113 6417 113 2 n_18
rlabel m2contact 6393 209 6393 209 2 n_89
rlabel m2contact 6345 113 6345 113 2 n_230
rlabel m2contact 6225 377 6225 377 2 n_302
rlabel m2contact 6057 353 6057 353 2 n_47
rlabel m2contact 5985 41 5985 41 2 Flags[0]
rlabel m2contact 5433 329 5433 329 2 n_359
rlabel m2contact 5289 305 5289 305 2 n_67
rlabel m2contact 5097 281 5097 281 2 n_131
rlabel m2contact 5049 89 5049 89 2 n_76
rlabel m2contact 4785 89 4785 89 2 n_171
rlabel m2contact 4761 257 4761 257 2 n_62
rlabel m2contact 4713 161 4713 161 2 n_37
rlabel m2contact 4617 161 4617 161 2 n_180
rlabel m2contact 4497 233 4497 233 2 n_124
rlabel m2contact 4137 209 4137 209 2 n_89
rlabel m2contact 3753 137 3753 137 2 n_353
rlabel m2contact 3681 137 3681 137 2 n_185
rlabel m2contact 3513 185 3513 185 2 n_24
rlabel m2contact 2841 161 2841 161 2 n_180
rlabel m2contact 2721 137 2721 137 2 n_185
rlabel m2contact 2697 113 2697 113 2 n_230
rlabel m2contact 1857 89 1857 89 2 n_171
rlabel m2contact 1737 89 1737 89 2 nWE
rlabel metal2 26127 7988 26139 7988 6 StatusRegEn
rlabel metal2 25287 7988 25299 7988 6 StatusReg[0]
rlabel metal2 24447 7988 24459 7988 6 StatusReg[1]
rlabel metal2 24423 7988 24435 7988 6 StatusReg[2]
rlabel metal2 22767 7988 22779 7988 6 StatusReg[3]
rlabel metal2 21927 7988 21939 7988 6 AluEn
rlabel metal2 21087 7988 21099 7988 6 AluWe
rlabel metal2 20247 7988 20259 7988 6 Op2Sel[0]
rlabel metal2 19767 7988 19779 7988 6 Op2Sel[1]
rlabel metal2 19263 7988 19275 7988 6 Op1Sel
rlabel metal2 18543 7988 18555 7988 6 WdSel
rlabel metal2 17631 7988 17643 7988 6 PcEn
rlabel metal2 16695 7988 16707 7988 6 PcWe
rlabel metal2 16023 7988 16035 7988 6 PcSel[0]
rlabel metal2 14367 7988 14379 7988 6 PcSel[1]
rlabel metal2 14343 7988 14355 7988 6 PcSel[2]
rlabel metal2 13491 7988 13503 7988 4 LrEn
rlabel metal2 11823 7988 11835 7988 4 LrWe
rlabel metal2 11787 7988 11799 7988 4 LrSel
rlabel metal2 10935 7988 10947 7988 4 ImmSel
rlabel metal2 10083 7988 10095 7988 4 IrWe
rlabel metal2 9231 7988 9243 7988 4 MemEn
rlabel metal2 8379 7988 8391 7988 4 OpcodeCondIn[0]
rlabel metal2 7527 7988 7539 7988 4 OpcodeCondIn[1]
rlabel metal2 5859 7988 5871 7988 4 OpcodeCondIn[2]
rlabel metal2 5823 7988 5835 7988 4 OpcodeCondIn[3]
rlabel metal2 4971 7988 4983 7988 4 OpcodeCondIn[4]
rlabel metal2 3303 7988 3315 7988 4 OpcodeCondIn[5]
rlabel metal2 2451 7988 2463 7988 4 OpcodeCondIn[6]
rlabel metal2 2415 7988 2427 7988 4 OpcodeCondIn[7]
rlabel metal2 24951 0 24963 0 8 SysBus[3]
rlabel metal2 17439 0 17451 0 8 SysBus[2]
rlabel metal2 11127 0 11139 0 2 SysBus[1]
rlabel metal2 7947 0 7959 0 2 SysBus[0]
rlabel metal2 27577 419 27577 431 8 Flags[2]
rlabel metal2 27577 395 27577 407 8 Flags[1]
rlabel metal2 27577 35 27577 47 8 Flags[0]
rlabel metal2 27577 11 27577 23 8 CFlag
rlabel metal2 27577 6772 27577 6784 6 RwSel[0]
rlabel metal2 27577 2956 27577 2968 6 Rs1Sel[1]
rlabel metal2 27577 1588 27577 1600 6 Rs1Sel[0]
rlabel metal2 27577 1564 27577 1576 6 Flags[3]
rlabel metal2 27577 7821 27577 7833 6 ENB
rlabel metal2 27577 7797 27577 7809 6 AluOR[1]
rlabel metal2 27577 7773 27577 7785 6 AluOR[0]
rlabel metal2 27577 7749 27577 7761 6 RegWe
rlabel metal2 27577 7725 27577 7737 6 RwSel[1]
rlabel metal2 27243 0 27443 0 1 GND!
rlabel metal2 27243 7988 27443 7988 5 GND!
rlabel metal2 0 83 0 95 2 nWE
rlabel metal2 0 59 0 71 2 nIRQ
rlabel metal2 0 3820 0 3832 4 nWait
rlabel metal2 0 3796 0 3808 4 nOE
rlabel metal2 0 7917 0 7929 4 ALE
rlabel metal2 0 7893 0 7905 4 nME
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 339 7988 351 7988 5 SDO
rlabel metal2 387 7988 399 7988 5 Clock
rlabel metal2 363 7988 375 7988 5 Test
rlabel metal2 411 7988 423 7988 5 nReset
rlabel metal2 123 7988 323 7988 5 Vdd!
<< end >>
