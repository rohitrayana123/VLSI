magic
tech c035u
timestamp 1394626552
<< metal1 >>
rect 481 22062 16460 22072
rect 16474 22062 23764 22072
rect 504 22038 16580 22048
rect 16594 22038 23764 22048
rect 527 22014 16700 22024
rect 16714 22014 23764 22024
rect 550 21990 16820 22000
rect 16834 21990 23764 22000
rect 573 21966 16940 21976
rect 16954 21966 23764 21976
rect 596 21942 4148 21952
rect 4162 21942 23764 21952
rect 619 21918 4580 21928
rect 4594 21918 23764 21928
rect 642 21894 5012 21904
rect 5026 21894 23764 21904
rect 665 21870 4196 21880
rect 4210 21870 23764 21880
rect 688 21846 4628 21856
rect 4642 21846 23764 21856
rect 711 21822 5060 21832
rect 5074 21822 23764 21832
rect 734 21798 7148 21808
rect 7162 21798 23764 21808
rect 757 21774 7124 21784
rect 7138 21774 22364 21784
rect 22378 21774 23764 21784
rect 780 21750 7100 21760
rect 7114 21750 22556 21760
rect 22570 21750 23764 21760
rect 803 21726 22676 21736
rect 22690 21726 23764 21736
rect 826 21702 22796 21712
rect 22810 21702 23764 21712
rect 23565 18891 23757 18901
rect 0 17893 467 17903
rect 481 17893 832 17903
rect 0 17861 832 17871
rect 0 17827 832 17837
rect 23565 17827 23757 17837
rect 23565 17715 23757 17725
rect 0 16717 490 16727
rect 504 16717 832 16727
rect 0 16685 832 16695
rect 0 16651 832 16661
rect 23565 16651 23757 16661
rect 23565 16539 23757 16549
rect 0 15541 513 15551
rect 527 15541 832 15551
rect 0 15509 832 15519
rect 0 15475 832 15485
rect 23565 15475 23757 15485
rect 23565 15363 23757 15373
rect 0 14365 536 14375
rect 550 14365 832 14375
rect 0 14333 832 14343
rect 0 14299 832 14309
rect 23565 14299 23757 14309
rect 23565 14187 23757 14197
rect 0 13189 559 13199
rect 573 13189 832 13199
rect 0 13157 832 13167
rect 0 13123 832 13133
rect 23565 13123 23757 13133
rect 23565 13011 23757 13021
rect 0 12013 582 12023
rect 596 12013 832 12023
rect 0 11981 832 11991
rect 0 11947 832 11957
rect 23565 11947 23757 11957
rect 23565 11835 23757 11845
rect 0 10837 605 10847
rect 619 10837 832 10847
rect 0 10805 832 10815
rect 0 10771 832 10781
rect 23565 10771 23757 10781
rect 23565 10659 23757 10669
rect 0 9661 628 9671
rect 642 9661 832 9671
rect 0 9629 832 9639
rect 0 9595 832 9605
rect 23565 9595 23757 9605
rect 23565 9483 23757 9493
rect 0 8485 651 8495
rect 665 8485 832 8495
rect 0 8453 832 8463
rect 0 8419 832 8429
rect 23565 8419 23757 8429
rect 23565 8307 23757 8317
rect 0 7309 674 7319
rect 688 7309 832 7319
rect 0 7277 832 7287
rect 0 7243 832 7253
rect 23565 7243 23757 7253
rect 23565 7131 23757 7141
rect 0 6133 697 6143
rect 711 6133 832 6143
rect 0 6101 832 6111
rect 0 6067 832 6077
rect 23565 6067 23757 6077
rect 23565 5955 23757 5965
rect 0 4957 720 4967
rect 734 4957 832 4967
rect 0 4925 832 4935
rect 0 4891 832 4901
rect 23565 4891 23757 4901
rect 23565 4779 23757 4789
rect 0 3781 743 3791
rect 757 3781 832 3791
rect 0 3749 832 3759
rect 0 3715 832 3725
rect 23565 3715 23757 3725
rect 23565 3603 23757 3613
rect 0 2605 766 2615
rect 780 2605 832 2615
rect 0 2573 832 2583
rect 0 2539 832 2549
rect 23565 2539 23757 2549
rect 23565 2427 23757 2437
rect 0 1429 789 1439
rect 803 1429 832 1439
rect 0 1397 832 1407
rect 0 1363 832 1373
rect 23565 1363 23757 1373
rect 23565 1251 23757 1261
rect 0 253 812 263
rect 826 253 832 263
rect 0 221 832 231
rect 0 187 832 197
rect 23565 187 23757 197
rect 2522 72 17252 82
rect 17266 72 19916 82
rect 19930 72 19963 82
rect 19977 72 20012 82
rect 20026 72 20060 82
rect 20074 72 20108 82
rect 20122 72 20156 82
rect 20170 72 20204 82
rect 20218 72 20252 82
rect 20266 72 20564 82
rect 20578 72 20612 82
rect 20626 72 20659 82
rect 20673 72 20708 82
rect 20722 72 21020 82
rect 21034 72 21068 82
rect 21082 72 21452 82
rect 21466 72 24813 82
rect 1037 51 3740 61
<< m2contact >>
rect 467 22060 481 22074
rect 16460 22061 16474 22075
rect 490 22036 504 22050
rect 16580 22036 16594 22050
rect 513 22012 527 22026
rect 16700 22012 16714 22026
rect 536 21988 550 22002
rect 16820 21988 16834 22002
rect 559 21964 573 21978
rect 16940 21964 16954 21978
rect 582 21940 596 21954
rect 4148 21940 4162 21954
rect 605 21916 619 21930
rect 4580 21916 4594 21930
rect 628 21892 642 21906
rect 5012 21892 5026 21906
rect 651 21868 665 21882
rect 4196 21868 4210 21882
rect 674 21844 688 21858
rect 4628 21844 4642 21858
rect 697 21820 711 21834
rect 5060 21820 5074 21834
rect 720 21796 734 21810
rect 7148 21796 7162 21810
rect 743 21772 757 21786
rect 7124 21772 7138 21786
rect 22364 21772 22378 21786
rect 766 21748 780 21762
rect 7100 21748 7114 21762
rect 22556 21747 22570 21761
rect 789 21724 803 21738
rect 22676 21724 22690 21738
rect 812 21700 826 21714
rect 22796 21700 22810 21714
rect 467 17891 481 17905
rect 490 16715 504 16729
rect 513 15539 527 15553
rect 536 14363 550 14377
rect 559 13187 573 13201
rect 582 12011 596 12025
rect 605 10835 619 10849
rect 628 9659 642 9673
rect 651 8483 665 8497
rect 674 7307 688 7321
rect 697 6131 711 6145
rect 720 4955 734 4969
rect 743 3779 757 3793
rect 766 2603 780 2617
rect 789 1427 803 1441
rect 812 251 826 265
rect 17252 70 17266 84
rect 19916 70 19930 84
rect 19963 70 19977 84
rect 20012 70 20026 84
rect 20060 70 20074 84
rect 20108 70 20122 84
rect 20156 70 20170 84
rect 20204 70 20218 84
rect 20252 70 20266 84
rect 20564 70 20578 84
rect 20612 70 20626 84
rect 20659 70 20673 84
rect 20708 70 20722 84
rect 21020 70 21034 84
rect 21068 70 21082 84
rect 21452 70 21466 84
rect 24813 70 24827 84
rect 1023 49 1037 63
rect 3740 48 3754 62
<< metal2 >>
rect 468 17905 480 22060
rect 491 16729 503 22036
rect 514 15553 526 22012
rect 537 14377 549 21988
rect 560 13201 572 21964
rect 583 12025 595 21940
rect 606 10849 618 21916
rect 629 9673 641 21892
rect 652 8497 664 21868
rect 675 7321 687 21844
rect 698 6145 710 21820
rect 721 4969 733 21796
rect 744 3793 756 21772
rect 767 2617 779 21748
rect 790 1441 802 21724
rect 813 265 825 21700
rect 837 21691 1037 22218
rect 1053 21691 1065 22218
rect 1077 21691 1089 22218
rect 1101 21691 1113 22218
rect 1125 21691 1137 22218
rect 4125 21691 4137 22218
rect 4149 21691 4161 21940
rect 4197 21691 4209 21868
rect 4365 21691 4377 22218
rect 4581 21691 4593 21916
rect 4629 21691 4641 21844
rect 5013 21691 5025 21892
rect 5061 21691 5073 21820
rect 5421 21691 5433 22218
rect 5661 21691 5673 22218
rect 6791 21691 6803 22218
rect 7101 21691 7113 21748
rect 7125 21691 7137 21772
rect 7149 21691 7161 21796
rect 16461 21691 16473 22061
rect 16581 21691 16593 22036
rect 16701 21691 16713 22012
rect 16821 21691 16833 21988
rect 16941 21691 16953 21964
rect 18045 21691 18057 22218
rect 18477 21691 18489 22218
rect 18669 21691 18681 22218
rect 18741 21691 18753 22218
rect 18837 21691 18849 22218
rect 22365 21691 22377 21772
rect 22557 21691 22569 21747
rect 22677 21691 22689 21724
rect 22797 21691 22809 21700
rect 24813 21691 25013 22218
rect 23613 18885 23625 18908
rect 23613 17709 23625 17843
rect 23613 16533 23625 16667
rect 23613 15357 23625 15491
rect 23613 14181 23625 14315
rect 23613 13005 23625 13139
rect 23613 11829 23625 11963
rect 23613 10653 23625 10787
rect 23613 9477 23625 9611
rect 23613 8301 23625 8435
rect 23613 7125 23625 7259
rect 23613 5949 23625 6083
rect 23613 4773 23625 4907
rect 23613 3597 23625 3731
rect 23613 2421 23625 2555
rect 23613 1245 23625 1379
rect 23613 92 23625 203
rect 837 63 1037 92
rect 837 49 1023 63
rect 837 0 1037 49
rect 1053 0 1065 92
rect 1077 0 1089 92
rect 1101 0 1113 92
rect 1125 0 1137 92
rect 2397 0 2409 92
rect 2589 0 2601 92
rect 3381 0 3393 92
rect 3741 62 3753 92
rect 3885 0 3897 92
rect 4101 0 4113 92
rect 4845 0 4857 92
rect 5013 0 5025 92
rect 5397 0 5409 92
rect 5613 0 5625 92
rect 6357 0 6369 92
rect 6525 0 6537 92
rect 15933 0 15945 92
rect 16125 0 16137 92
rect 16773 83 16785 92
rect 16965 83 16977 92
rect 17253 84 17265 92
rect 19917 84 19929 92
rect 19965 84 19977 92
rect 20013 84 20025 92
rect 20061 84 20073 92
rect 20109 84 20121 92
rect 20157 84 20169 92
rect 20205 84 20217 92
rect 20253 84 20265 92
rect 20565 84 20577 92
rect 20613 84 20625 92
rect 20661 84 20673 92
rect 20709 84 20721 92
rect 21021 84 21033 92
rect 21069 84 21081 92
rect 21453 84 21465 92
rect 16773 71 16977 83
rect 23829 0 23841 92
rect 24573 0 24585 92
rect 24813 84 25013 92
rect 24827 70 25013 84
rect 24813 0 25013 70
use slice17 slice17_0
timestamp 1394626552
transform 1 0 837 0 1 18908
box 0 0 24176 2783
use leftbuf_slice leftbuf_slice_0
array 0 0 1685 0 15 1176
timestamp 1394551156
transform 1 0 832 0 1 98
box 0 -6 1685 1170
use IrAA IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 2517 0 1 9611
box 0 -111 1008 1065
use IrBA IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 2517 0 1 6083
box 0 -111 1008 1065
use IrBB IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 2517 0 1 204
box 0 -112 1008 1064
use Datapath_slice Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394620980
transform 1 0 3525 0 1 92
box 0 0 20040 1176
use LLIcell_U LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1394560148
transform 1 0 23565 0 1 9611
box 0 0 192 1042
use LLIcell_L LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 23565 0 1 203
box 0 0 192 1042
use Datapath_end Datapath_end_0
array 0 0 1256 0 15 1176
timestamp 1394624888
transform 1 0 23757 0 1 92
box 0 0 1256 1176
<< labels >>
rlabel metal1 0 187 0 197 3 SysBus[0]
rlabel metal1 0 1363 0 1373 3 SysBus[1]
rlabel metal1 0 2539 0 2549 3 SysBus[2]
rlabel metal1 0 3715 0 3725 3 SysBus[3]
rlabel metal1 0 4891 0 4901 3 SysBus[4]
rlabel metal1 0 6067 0 6077 3 SysBus[5]
rlabel metal1 0 7243 0 7253 3 SysBus[6]
rlabel metal1 0 8419 0 8429 3 SysBus[7]
rlabel metal1 0 9595 0 9605 3 SysBus[8]
rlabel metal1 0 10771 0 10781 3 SysBus[9]
rlabel metal1 0 11947 0 11957 3 SysBus[10]
rlabel metal1 0 13123 0 13133 3 SysBus[11]
rlabel metal1 0 14299 0 14309 3 SysBus[12]
rlabel metal1 0 15475 0 15485 3 SysBus[13]
rlabel metal1 0 16651 0 16661 3 SysBus[14]
rlabel metal1 0 17827 0 17837 3 SysBus[15]
rlabel metal1 0 253 0 263 3 Ir[0]
rlabel metal1 0 1429 0 1439 3 Ir[1]
rlabel metal1 0 2605 0 2615 3 Ir[2]
rlabel metal1 0 3781 0 3791 3 Ir[3]
rlabel metal1 0 4957 0 4967 3 Ir[4]
rlabel metal1 0 6133 0 6143 3 Ir[5]
rlabel metal1 0 7309 0 7319 3 Ir[6]
rlabel metal1 0 8485 0 8495 3 Ir[7]
rlabel metal1 0 9661 0 9671 3 Ir[8]
rlabel metal1 0 10837 0 10847 3 Ir[9]
rlabel metal1 0 12013 0 12023 3 Ir[10]
rlabel metal1 0 13189 0 13199 3 Ir[11]
rlabel metal1 0 14365 0 14375 3 Ir[12]
rlabel metal1 0 15541 0 15551 3 Ir[13]
rlabel metal1 0 16717 0 16727 3 Ir[14]
rlabel metal1 0 17893 0 17903 3 Ir[15]
rlabel metal2 837 0 1037 0 1 Vdd!
rlabel metal2 1053 0 1065 0 1 SDI
rlabel metal2 1077 0 1089 0 1 Test
rlabel metal2 1101 0 1113 0 1 Clock
rlabel metal2 1125 0 1137 0 1 nReset
rlabel metal2 3885 0 3897 0 1 LrSel
rlabel metal2 4101 0 4113 0 1 LrWe
rlabel metal2 4845 0 4857 0 1 LrEn
rlabel metal2 5013 0 5025 0 1 PcSel[0]
rlabel metal2 5397 0 5409 0 1 PcSel[1]
rlabel metal2 5613 0 5625 0 1 PcWe
rlabel metal2 6357 0 6369 0 1 PcEn
rlabel metal2 6525 0 6537 0 1 WdSel
rlabel metal2 16125 0 16137 0 1 Op2Sel
rlabel metal2 15933 0 15945 0 1 Op1Sel
rlabel metal2 3381 0 3393 0 1 ImmSel
rlabel metal2 2589 0 2601 0 1 IrWe
rlabel metal1 0 221 0 231 3 DataIn[0]
rlabel metal1 0 17861 0 17871 3 DataIn[15]
rlabel metal1 0 16685 0 16695 3 DataIn[14]
rlabel metal1 0 15509 0 15519 3 DataIn[13]
rlabel metal1 0 14333 0 14343 3 DataIn[12]
rlabel metal1 0 13157 0 13167 3 DataIn[11]
rlabel metal1 0 11981 0 11991 3 DataIn[10]
rlabel metal1 0 10805 0 10815 3 DataIn[9]
rlabel metal1 0 9629 0 9639 3 DataIn[8]
rlabel metal1 0 8453 0 8463 3 DataIn[7]
rlabel metal1 0 7277 0 7287 3 DataIn[6]
rlabel metal1 0 6101 0 6111 3 DataIn[5]
rlabel metal1 0 4925 0 4935 3 DataIn[4]
rlabel metal1 0 3749 0 3759 3 DataIn[3]
rlabel metal1 0 2573 0 2583 3 DataIn[2]
rlabel metal1 0 1397 0 1407 3 DataIn[1]
rlabel metal2 2397 0 2409 0 1 MemEn
rlabel metal2 24813 0 25013 0 1 GND!
rlabel metal2 24573 0 24585 0 1 AluEn
rlabel metal2 23829 0 23841 0 1 AluWe
rlabel metal2 750 21769 750 21769 1 Ir[3]
rlabel metal2 727 21770 727 21770 1 Ir[4]
rlabel metal2 704 21769 704 21769 1 Ir[5]
rlabel metal2 681 21768 681 21768 1 Ir[6]
rlabel metal2 658 21767 658 21767 1 Ir[7]
rlabel metal2 635 21765 635 21765 1 Ir[8]
rlabel metal2 612 21765 612 21765 1 Ir[9]
rlabel metal2 589 21764 589 21764 1 Ir[10]
rlabel metal2 566 21765 566 21765 1 Ir[11]
rlabel metal2 543 21765 543 21765 1 Ir[12]
rlabel metal2 520 21764 520 21764 1 Ir[13]
rlabel metal2 497 21764 497 21764 1 Ir[14]
rlabel metal2 473 21765 473 21765 1 Ir[15]
rlabel metal2 1077 22218 1089 22218 1 Test
rlabel metal2 1101 22218 1113 22218 1 Clock
rlabel metal2 1125 22218 1137 22218 1 nReset
rlabel metal2 837 22218 1037 22218 5 Vdd!
rlabel metal2 6791 22218 6803 22218 5 RegWe
rlabel metal2 7105 21740 7105 21740 1 Ir[2]
rlabel metal2 7131 21764 7131 21764 1 Ir[3]
rlabel metal2 7154 21788 7154 21788 1 Ir[4]
rlabel metal2 4125 22218 4137 22218 5 Rs1Sel[0]
rlabel metal2 4365 22218 4377 22218 5 Rs1Sel[1]
rlabel metal1 4606 21947 4606 21947 1 Ir[10]
rlabel metal2 5421 22218 5433 22218 5 RwSel[0]
rlabel metal2 5661 22218 5673 22218 5 RwSel[1]
rlabel metal2 4154 21933 4154 21933 1 Ir[10]
rlabel metal2 4203 21860 4203 21860 1 Ir[7]
rlabel metal2 4586 21908 4586 21908 1 Ir[9]
rlabel metal2 4635 21837 4635 21837 1 Ir[6]
rlabel metal2 5018 21885 5018 21885 1 Ir[8]
rlabel metal2 5068 21814 5068 21814 1 Ir[5]
rlabel metal2 24813 22218 25013 22218 1 GND!
rlabel metal2 1053 22218 1065 22218 5 SDO
rlabel metal2 16466 22054 16466 22054 1 Ir[15]
rlabel metal2 16585 22029 16585 22029 1 Ir[14]
rlabel metal2 16706 22006 16706 22006 1 Ir[13]
rlabel metal2 16827 21982 16827 21982 1 Ir[12]
rlabel metal2 16947 21957 16947 21957 1 Ir[11]
rlabel metal2 18045 22218 18057 22218 5 CFlag
rlabel metal2 18477 22218 18489 22218 5 Flags[2]
rlabel metal2 18669 22218 18681 22218 5 Flags[1]
rlabel metal2 18741 22218 18753 22218 5 Flags[3]
rlabel metal2 18837 22218 18849 22218 5 Flags[0]
rlabel metal2 22371 21767 22371 21767 1 Ir[3]
rlabel metal2 22562 21742 22562 21742 1 Ir[2]
rlabel metal2 22682 21717 22682 21717 1 Ir[1]
rlabel metal2 22803 21695 22803 21695 1 Ir[0]
<< end >>
