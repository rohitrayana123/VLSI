magic
tech c035u
timestamp 1394047590
<< metal1 >>
rect 13455 1865 16752 1875
rect 12303 1837 16367 1847
rect 3133 1785 6670 1795
rect 9998 1781 14330 1791
rect 11150 1717 14246 1727
rect 2416 1680 14400 1690
rect 2416 1495 2426 1680
rect 3091 1655 13248 1665
rect 2933 1635 12096 1645
rect 2825 1615 10944 1625
rect 2703 1590 9792 1600
rect 2546 1557 8639 1569
rect 8847 1567 15699 1577
rect 2639 1533 7487 1543
rect 2483 1506 6335 1517
rect 2270 1485 2426 1495
rect 5990 1485 14184 1495
rect 2030 1455 3078 1465
rect 5750 1455 13031 1465
rect 16357 1465 16367 1837
rect 16356 1455 16512 1465
rect 1791 1430 2920 1440
rect 5511 1430 11880 1440
rect 14261 1430 16272 1440
rect 1551 1407 2809 1417
rect 5271 1407 10728 1417
rect 14344 1407 16031 1417
rect 63 1383 1366 1393
rect 1385 1383 1608 1393
rect 1622 1383 1848 1393
rect 1862 1383 2088 1393
rect 3784 1383 5086 1393
rect 5105 1383 5328 1393
rect 5342 1383 5568 1393
rect 5582 1383 5808 1393
rect 14559 1383 15862 1393
rect 15881 1383 16104 1393
rect 16118 1383 16344 1393
rect 16358 1383 16584 1393
rect 350 1358 455 1368
rect 470 1358 936 1368
rect 950 1358 1416 1368
rect 1430 1358 1896 1368
rect 4070 1358 4175 1368
rect 4190 1358 4656 1368
rect 4670 1358 5136 1368
rect 5150 1358 5616 1368
rect 14846 1358 14951 1368
rect 14966 1358 15432 1368
rect 15446 1358 15912 1368
rect 15926 1358 16392 1368
rect 184 1332 912 1342
rect 926 1332 1152 1342
rect 1166 1332 1872 1342
rect 1886 1332 2112 1342
rect 3904 1332 4632 1342
rect 4646 1332 4872 1342
rect 4886 1332 5592 1342
rect 5606 1332 5832 1342
rect 7695 1340 13937 1350
rect 14680 1332 15408 1342
rect 15422 1332 15648 1342
rect 15662 1332 16368 1342
rect 16382 1332 16608 1342
rect 111 1297 408 1307
rect 422 1297 648 1307
rect 662 1297 888 1307
rect 902 1297 1124 1307
rect 1311 1295 2689 1305
rect 3831 1297 4128 1307
rect 4142 1297 4368 1307
rect 4382 1297 4608 1307
rect 4622 1297 4844 1307
rect 5031 1295 9574 1305
rect 14607 1297 14904 1307
rect 14918 1297 15144 1307
rect 15158 1297 15384 1307
rect 15398 1297 15620 1307
rect 15713 1295 15790 1305
rect 303 1275 695 1285
rect 1072 1273 2531 1283
rect 4023 1275 4415 1285
rect 4792 1273 8424 1283
rect 14799 1275 15191 1285
rect 15520 1275 15551 1285
rect 230 1246 431 1257
rect 447 1246 672 1257
rect 686 1246 1392 1257
rect 1406 1246 1632 1257
rect 3950 1246 4151 1257
rect 4167 1246 4392 1257
rect 4406 1246 5112 1257
rect 5126 1246 5352 1257
rect 6543 1250 7428 1260
rect 831 1221 2623 1231
rect 4551 1221 7272 1231
rect 7418 1231 7428 1250
rect 14726 1246 14927 1257
rect 14943 1246 15168 1257
rect 15182 1246 15888 1257
rect 15902 1246 16128 1257
rect 7418 1221 15311 1231
rect 754 1198 1176 1208
rect 1191 1198 1656 1208
rect 1670 1198 2136 1208
rect 4472 1198 4896 1208
rect 4911 1198 5376 1208
rect 5390 1198 5856 1208
rect 15244 1198 15672 1208
rect 15687 1198 16152 1208
rect 16166 1198 16632 1208
rect 590 1176 2469 1187
rect 4310 1176 6120 1187
rect 6690 1180 15072 1190
rect 15124 1165 15503 1175
rect 2919 1144 3048 1154
rect 3062 1144 6480 1154
rect 6494 1144 7632 1154
rect 7647 1144 8784 1154
rect 8798 1144 9936 1154
rect 9950 1144 11088 1154
rect 11102 1144 12239 1154
rect 12254 1144 13392 1154
rect 15124 1161 15134 1165
rect 13951 1151 15134 1161
rect 3638 1107 6048 1117
rect 6062 1107 6264 1117
rect 494 1074 528 1084
rect 734 1075 768 1085
rect 974 1075 1008 1085
rect 1215 1080 1248 1090
rect 1454 1080 1488 1090
rect 1694 1080 1728 1090
rect 1934 1080 1968 1090
rect 2175 1080 2207 1090
rect 4214 1074 4248 1084
rect 4454 1075 4488 1085
rect 4694 1075 4728 1085
rect 4935 1080 4968 1090
rect 5174 1080 5208 1090
rect 5414 1080 5448 1090
rect 7069 1094 7200 1104
rect 5654 1080 5688 1090
rect 5895 1080 5927 1090
rect 7214 1094 7416 1104
rect 8221 1094 8352 1104
rect 8366 1094 8568 1104
rect 9373 1094 9504 1104
rect 9518 1094 9720 1104
rect 10525 1094 10656 1104
rect 10670 1094 10872 1104
rect 11677 1094 11808 1104
rect 11822 1094 12024 1104
rect 12829 1094 12960 1104
rect 12974 1094 13176 1104
rect 13981 1094 14112 1104
rect 14126 1094 14328 1104
rect 14990 1074 15024 1084
rect 15230 1075 15264 1085
rect 15470 1075 15504 1085
rect 15711 1080 15744 1090
rect 15950 1080 15984 1090
rect 16190 1080 16224 1090
rect 16430 1080 16464 1090
rect 16671 1080 16703 1090
rect 0 990 25 1015
rect 16801 990 16815 1015
rect 0 345 25 370
rect 16801 345 16815 370
rect 0 322 25 332
rect 16801 322 16815 332
rect 0 276 25 286
rect 16801 276 16815 286
rect 0 75 2328 85
rect 2342 75 16815 85
rect 0 40 6191 50
rect 6206 40 7343 50
rect 7358 40 8495 50
rect 8510 40 9648 50
rect 9663 40 10798 50
rect 10816 40 11950 50
rect 11968 40 13102 50
rect 13120 40 14256 50
rect 14270 40 16815 50
rect 0 5 6408 15
rect 6422 5 7560 15
rect 7574 5 8712 15
rect 8726 5 9864 15
rect 9879 5 11015 15
rect 11033 5 12167 15
rect 12185 5 13319 15
rect 13337 5 14472 15
rect 14486 5 16815 15
<< m2contact >>
rect 13440 1863 13455 1877
rect 16752 1863 16766 1877
rect 12288 1835 12303 1849
rect 3118 1784 3133 1798
rect 6670 1776 6691 1799
rect 9982 1779 9998 1793
rect 14330 1779 14345 1793
rect 11136 1716 11150 1730
rect 14246 1716 14260 1730
rect 2256 1484 2270 1498
rect 14400 1679 14414 1693
rect 3075 1655 3091 1669
rect 13248 1654 13262 1668
rect 2918 1635 2933 1649
rect 12096 1631 12110 1645
rect 2808 1613 2825 1627
rect 10944 1611 10958 1625
rect 2688 1587 2703 1602
rect 9792 1589 9806 1603
rect 2530 1554 2546 1570
rect 8639 1555 8657 1570
rect 8829 1564 8847 1580
rect 15699 1566 15713 1580
rect 2625 1532 2639 1546
rect 7487 1531 7502 1545
rect 2469 1505 2483 1519
rect 6335 1505 6350 1519
rect 5976 1482 5990 1496
rect 14184 1484 14198 1498
rect 2016 1453 2030 1467
rect 3078 1454 3092 1468
rect 5736 1453 5750 1467
rect 13031 1453 13047 1467
rect 16512 1453 16526 1467
rect 1776 1428 1791 1442
rect 2920 1429 2934 1443
rect 5496 1428 5511 1442
rect 11880 1429 11894 1443
rect 14247 1428 14261 1442
rect 16272 1428 16287 1442
rect 1535 1404 1551 1419
rect 2809 1405 2823 1419
rect 5255 1404 5271 1419
rect 10728 1405 10742 1419
rect 14330 1405 14344 1419
rect 16031 1404 16047 1419
rect 49 1382 63 1396
rect 1366 1381 1385 1397
rect 1608 1380 1622 1394
rect 1848 1382 1862 1396
rect 2088 1382 2103 1396
rect 3769 1382 3784 1396
rect 5086 1381 5105 1397
rect 5328 1380 5342 1394
rect 5568 1382 5582 1396
rect 5808 1382 5823 1396
rect 14545 1382 14559 1396
rect 15862 1381 15881 1397
rect 16104 1380 16118 1394
rect 16344 1382 16358 1396
rect 16584 1382 16599 1396
rect 336 1357 350 1371
rect 455 1357 470 1371
rect 936 1357 950 1371
rect 1416 1357 1430 1371
rect 1896 1356 1911 1370
rect 4056 1357 4070 1371
rect 4175 1357 4190 1371
rect 4656 1357 4670 1371
rect 5136 1357 5150 1371
rect 5616 1356 5631 1370
rect 14832 1357 14846 1371
rect 14951 1357 14966 1371
rect 15432 1357 15446 1371
rect 15912 1357 15926 1371
rect 16392 1356 16407 1370
rect 167 1330 184 1344
rect 912 1332 926 1346
rect 1152 1331 1166 1345
rect 1872 1331 1886 1345
rect 2112 1330 2127 1344
rect 3887 1330 3904 1344
rect 4632 1332 4646 1346
rect 4872 1331 4886 1345
rect 5592 1331 5606 1345
rect 5832 1330 5847 1344
rect 7681 1339 7695 1353
rect 13937 1338 13952 1352
rect 14663 1330 14680 1344
rect 15408 1332 15422 1346
rect 15648 1331 15662 1345
rect 16368 1331 16382 1345
rect 16608 1330 16623 1344
rect 96 1295 111 1309
rect 408 1295 422 1309
rect 648 1296 662 1310
rect 888 1296 902 1310
rect 1124 1295 1141 1312
rect 1294 1293 1311 1307
rect 2689 1294 2703 1308
rect 3816 1295 3831 1309
rect 4128 1295 4142 1309
rect 4368 1296 4382 1310
rect 4608 1296 4622 1310
rect 4844 1295 4861 1312
rect 5014 1293 5031 1307
rect 9574 1293 9593 1310
rect 14592 1295 14607 1309
rect 14904 1295 14918 1309
rect 15144 1296 15158 1310
rect 15384 1296 15398 1310
rect 15620 1295 15637 1312
rect 15699 1293 15713 1307
rect 15790 1293 15807 1307
rect 288 1273 303 1287
rect 695 1269 711 1287
rect 1055 1270 1072 1285
rect 2531 1271 2545 1285
rect 4008 1273 4023 1287
rect 4415 1269 4431 1287
rect 4775 1270 4792 1285
rect 8424 1271 8438 1285
rect 14784 1273 14799 1287
rect 15191 1269 15207 1287
rect 15503 1271 15520 1286
rect 15551 1270 15568 1285
rect 216 1245 230 1259
rect 431 1244 447 1258
rect 672 1245 686 1259
rect 1392 1245 1406 1259
rect 1632 1245 1646 1259
rect 3936 1245 3950 1259
rect 4151 1244 4167 1258
rect 4392 1245 4406 1259
rect 5112 1245 5126 1259
rect 5352 1245 5366 1259
rect 6528 1248 6543 1262
rect 815 1219 831 1233
rect 2623 1220 2637 1234
rect 4535 1219 4551 1233
rect 7272 1220 7287 1234
rect 14712 1245 14726 1259
rect 14927 1244 14943 1258
rect 15168 1245 15182 1259
rect 15888 1245 15902 1259
rect 16128 1245 16142 1259
rect 15311 1219 15327 1233
rect 740 1197 754 1211
rect 1176 1197 1191 1211
rect 1656 1197 1670 1211
rect 2136 1197 2150 1211
rect 4458 1197 4472 1211
rect 4896 1197 4911 1211
rect 5376 1197 5390 1211
rect 5856 1197 5870 1211
rect 15230 1197 15244 1211
rect 15672 1197 15687 1211
rect 16152 1197 16166 1211
rect 16632 1197 16646 1211
rect 576 1176 590 1190
rect 2469 1175 2483 1189
rect 4296 1176 4310 1190
rect 6120 1175 6134 1189
rect 6674 1177 6690 1193
rect 15072 1176 15086 1190
rect 2903 1139 2919 1155
rect 3048 1141 3062 1155
rect 6480 1143 6494 1157
rect 7632 1143 7647 1157
rect 8784 1143 8798 1157
rect 9936 1143 9950 1157
rect 11088 1143 11102 1157
rect 12239 1142 12254 1156
rect 13392 1143 13407 1158
rect 13937 1150 13951 1164
rect 15503 1161 15520 1176
rect 3624 1105 3638 1119
rect 6048 1105 6062 1119
rect 6264 1104 6278 1118
rect 480 1071 494 1085
rect 528 1071 542 1085
rect 720 1074 734 1088
rect 768 1073 782 1087
rect 960 1074 974 1088
rect 1008 1074 1022 1088
rect 1200 1078 1215 1092
rect 1248 1078 1263 1092
rect 1439 1078 1454 1092
rect 1488 1078 1503 1092
rect 1680 1079 1694 1093
rect 1728 1078 1742 1092
rect 1920 1079 1934 1093
rect 1968 1078 1982 1092
rect 2160 1078 2175 1092
rect 2207 1078 2222 1092
rect 4200 1071 4214 1085
rect 4248 1071 4262 1085
rect 4440 1074 4454 1088
rect 4488 1073 4502 1087
rect 4680 1074 4694 1088
rect 4728 1074 4742 1088
rect 4920 1078 4935 1092
rect 4968 1078 4983 1092
rect 5159 1078 5174 1092
rect 5208 1078 5223 1092
rect 5400 1079 5414 1093
rect 5448 1078 5462 1092
rect 5640 1079 5654 1093
rect 7055 1092 7069 1106
rect 5688 1078 5702 1092
rect 5880 1078 5895 1092
rect 5927 1078 5942 1092
rect 7200 1091 7214 1105
rect 7416 1092 7430 1106
rect 8207 1092 8221 1106
rect 8352 1091 8366 1105
rect 8568 1092 8582 1106
rect 9359 1092 9373 1106
rect 9504 1091 9518 1105
rect 9720 1092 9734 1106
rect 10511 1092 10525 1106
rect 10656 1091 10670 1105
rect 10872 1092 10886 1106
rect 11663 1092 11677 1106
rect 11808 1091 11822 1105
rect 12024 1092 12038 1106
rect 12815 1092 12829 1106
rect 12960 1091 12974 1105
rect 13176 1092 13190 1106
rect 13967 1092 13981 1106
rect 14112 1091 14126 1105
rect 14328 1092 14342 1106
rect 14976 1071 14990 1085
rect 15024 1071 15038 1085
rect 15216 1074 15230 1088
rect 15264 1073 15278 1087
rect 15456 1074 15470 1088
rect 15504 1074 15518 1088
rect 15696 1078 15711 1092
rect 15744 1078 15759 1092
rect 15935 1078 15950 1092
rect 15984 1078 15999 1092
rect 16176 1079 16190 1093
rect 16224 1078 16238 1092
rect 16416 1079 16430 1093
rect 16464 1078 16478 1092
rect 16656 1078 16671 1092
rect 16703 1078 16717 1092
rect 2328 74 2342 88
rect 6191 38 6206 52
rect 7343 38 7358 52
rect 8495 38 8510 52
rect 9648 38 9663 53
rect 10798 38 10816 53
rect 11950 38 11968 53
rect 13102 38 13120 53
rect 14256 37 14270 52
rect 6408 4 6422 18
rect 7560 4 7574 18
rect 8712 4 8726 18
rect 9864 3 9879 18
rect 11015 0 11033 15
rect 12167 0 12185 15
rect 13319 0 13337 15
rect 14472 3 14486 18
<< metal2 >>
rect 49 1396 61 1895
rect 49 1068 61 1382
rect 169 1344 181 1895
rect 97 1068 109 1295
rect 169 1068 181 1330
rect 289 1287 301 1895
rect 217 1068 229 1245
rect 289 1068 301 1273
rect 337 1068 349 1357
rect 409 1068 421 1295
rect 433 1068 445 1244
rect 457 1068 469 1357
rect 481 1068 493 1071
rect 529 1068 541 1071
rect 577 1068 589 1176
rect 649 1068 661 1296
rect 711 1273 752 1285
rect 673 1068 685 1245
rect 697 1068 709 1269
rect 740 1211 752 1273
rect 721 1068 733 1074
rect 769 1068 781 1073
rect 817 1068 829 1219
rect 889 1068 901 1296
rect 913 1068 925 1332
rect 937 1068 949 1357
rect 961 1068 973 1074
rect 1009 1068 1021 1074
rect 1057 1068 1069 1270
rect 1129 1068 1141 1295
rect 1153 1068 1165 1331
rect 1177 1068 1189 1197
rect 1201 1068 1213 1078
rect 1249 1068 1261 1078
rect 1297 1068 1309 1293
rect 1369 1068 1381 1381
rect 1393 1068 1405 1245
rect 1417 1068 1429 1357
rect 1441 1068 1453 1078
rect 1489 1068 1501 1078
rect 1537 1068 1549 1404
rect 1609 1068 1621 1380
rect 1633 1068 1645 1245
rect 1657 1068 1669 1197
rect 1681 1068 1693 1079
rect 1729 1068 1741 1078
rect 1777 1068 1789 1428
rect 1849 1068 1861 1382
rect 1873 1068 1885 1331
rect 1897 1068 1909 1356
rect 1921 1068 1933 1079
rect 1969 1068 1981 1078
rect 2017 1068 2029 1453
rect 2089 1068 2101 1382
rect 2113 1068 2125 1330
rect 2137 1068 2149 1197
rect 2161 1068 2173 1078
rect 2209 1068 2221 1078
rect 2257 1068 2269 1484
rect 2377 1068 2389 1895
rect 3119 1798 3131 1895
rect 2470 1189 2482 1505
rect 2532 1285 2544 1554
rect 2625 1234 2637 1532
rect 2690 1308 2702 1587
rect 2810 1419 2822 1613
rect 2920 1443 2932 1635
rect 3079 1468 3091 1655
rect 3119 1223 3131 1784
rect 3097 1211 3131 1223
rect 3769 1396 3781 1895
rect 2905 1068 2917 1139
rect 3049 1068 3061 1141
rect 3097 1068 3109 1211
rect 3625 1068 3637 1105
rect 3769 1068 3781 1382
rect 3889 1344 3901 1895
rect 3817 1068 3829 1295
rect 3889 1068 3901 1330
rect 4009 1287 4021 1895
rect 3937 1068 3949 1245
rect 4009 1068 4021 1273
rect 4057 1068 4069 1357
rect 4129 1068 4141 1295
rect 4153 1068 4165 1244
rect 4177 1068 4189 1357
rect 4201 1068 4213 1071
rect 4249 1068 4261 1071
rect 4297 1068 4309 1176
rect 4369 1068 4381 1296
rect 4431 1273 4471 1285
rect 4393 1068 4405 1245
rect 4417 1068 4429 1269
rect 4459 1211 4471 1273
rect 4441 1068 4453 1074
rect 4489 1068 4501 1073
rect 4537 1068 4549 1219
rect 4609 1068 4621 1296
rect 4633 1068 4645 1332
rect 4657 1068 4669 1357
rect 4681 1068 4693 1074
rect 4729 1068 4741 1074
rect 4777 1068 4789 1270
rect 4849 1068 4861 1295
rect 4873 1068 4885 1331
rect 4897 1068 4909 1197
rect 4921 1068 4933 1078
rect 4969 1068 4981 1078
rect 5017 1068 5029 1293
rect 5089 1068 5101 1381
rect 5113 1068 5125 1245
rect 5137 1068 5149 1357
rect 5161 1068 5173 1078
rect 5209 1068 5221 1078
rect 5257 1068 5269 1404
rect 5329 1068 5341 1380
rect 5353 1068 5365 1245
rect 5377 1068 5389 1197
rect 5401 1068 5413 1079
rect 5449 1068 5461 1078
rect 5497 1068 5509 1428
rect 5569 1068 5581 1382
rect 5593 1068 5605 1331
rect 5617 1068 5629 1356
rect 5641 1068 5653 1079
rect 5689 1068 5701 1078
rect 5737 1068 5749 1453
rect 5809 1068 5821 1382
rect 5833 1068 5845 1330
rect 5857 1068 5869 1197
rect 5881 1068 5893 1078
rect 5929 1068 5941 1078
rect 5977 1068 5989 1482
rect 6049 1068 6061 1105
rect 6121 1068 6133 1175
rect 6265 1068 6277 1104
rect 6337 1068 6349 1505
rect 6481 1068 6493 1143
rect 6529 1068 6541 1248
rect 6675 1193 6687 1776
rect 7057 1068 7069 1092
rect 7201 1068 7213 1091
rect 7273 1068 7285 1220
rect 7417 1068 7429 1092
rect 7489 1068 7501 1531
rect 7633 1068 7645 1143
rect 7681 1068 7693 1339
rect 8209 1068 8221 1092
rect 8353 1068 8365 1091
rect 8425 1068 8437 1271
rect 8569 1068 8581 1092
rect 8641 1068 8653 1555
rect 8785 1068 8797 1143
rect 8833 1068 8845 1564
rect 9361 1068 9373 1092
rect 9505 1068 9517 1091
rect 9577 1068 9589 1293
rect 9721 1068 9733 1092
rect 9793 1068 9805 1589
rect 9937 1068 9949 1143
rect 9985 1068 9997 1779
rect 10513 1068 10525 1092
rect 10657 1068 10669 1091
rect 10729 1068 10741 1405
rect 10873 1068 10885 1092
rect 10945 1068 10957 1611
rect 11089 1068 11101 1143
rect 11137 1068 11149 1716
rect 11665 1068 11677 1092
rect 11809 1068 11821 1091
rect 11881 1068 11893 1429
rect 12025 1068 12037 1092
rect 12097 1068 12109 1631
rect 12241 1068 12253 1142
rect 12289 1068 12301 1835
rect 12817 1068 12829 1092
rect 12961 1068 12973 1091
rect 13033 1068 13045 1453
rect 13177 1068 13189 1092
rect 13249 1068 13261 1654
rect 13393 1068 13405 1143
rect 13441 1068 13453 1863
rect 13938 1164 13950 1338
rect 13969 1068 13981 1092
rect 14113 1068 14125 1091
rect 14185 1068 14197 1484
rect 14247 1442 14259 1716
rect 14331 1419 14343 1779
rect 14329 1068 14341 1092
rect 14401 1068 14413 1679
rect 14545 1396 14557 1895
rect 14545 1068 14557 1382
rect 14665 1344 14677 1895
rect 14593 1068 14605 1295
rect 14665 1068 14677 1330
rect 14785 1287 14797 1895
rect 14713 1068 14725 1245
rect 14785 1068 14797 1273
rect 14833 1068 14845 1357
rect 14905 1068 14917 1295
rect 14929 1068 14941 1244
rect 14953 1068 14965 1357
rect 14977 1068 14989 1071
rect 15025 1068 15037 1071
rect 15073 1068 15085 1176
rect 15145 1068 15157 1296
rect 15207 1274 15242 1286
rect 15169 1068 15181 1245
rect 15193 1068 15205 1269
rect 15230 1211 15242 1274
rect 15217 1068 15229 1074
rect 15265 1068 15277 1073
rect 15313 1068 15325 1219
rect 15385 1068 15397 1296
rect 15409 1068 15421 1332
rect 15433 1068 15445 1357
rect 15505 1176 15517 1271
rect 15457 1068 15469 1074
rect 15505 1068 15517 1074
rect 15553 1068 15565 1270
rect 15625 1068 15637 1295
rect 15649 1068 15661 1331
rect 15700 1307 15712 1566
rect 15673 1068 15685 1197
rect 15697 1068 15709 1078
rect 15745 1068 15757 1078
rect 15793 1068 15805 1293
rect 15865 1068 15877 1381
rect 15889 1068 15901 1245
rect 15913 1068 15925 1357
rect 15937 1068 15949 1078
rect 15985 1068 15997 1078
rect 16033 1068 16045 1404
rect 16105 1068 16117 1380
rect 16129 1068 16141 1245
rect 16153 1068 16165 1197
rect 16177 1068 16189 1079
rect 16225 1068 16237 1078
rect 16273 1068 16285 1428
rect 16345 1068 16357 1382
rect 16369 1068 16381 1331
rect 16393 1068 16405 1356
rect 16417 1068 16429 1079
rect 16465 1068 16477 1078
rect 16513 1068 16525 1453
rect 16585 1068 16597 1382
rect 16609 1068 16621 1330
rect 16633 1068 16645 1197
rect 16657 1068 16669 1078
rect 16705 1068 16717 1078
rect 16753 1068 16765 1863
rect 2329 88 2341 269
rect 6193 52 6205 269
rect 6409 18 6421 269
rect 7345 52 7357 269
rect 7561 18 7573 269
rect 8497 52 8509 269
rect 8713 18 8725 269
rect 9649 53 9661 269
rect 9865 18 9877 269
rect 10801 53 10813 269
rect 11017 15 11029 269
rect 11953 53 11965 269
rect 12169 15 12181 269
rect 13105 53 13117 269
rect 13321 15 13333 269
rect 14257 52 14269 269
rect 14473 18 14485 269
use inv inv_11
timestamp 1386238110
transform 1 0 25 0 1 269
box 0 0 120 799
use inv inv_12
timestamp 1386238110
transform 1 0 145 0 1 269
box 0 0 120 799
use inv inv_13
timestamp 1386238110
transform 1 0 265 0 1 269
box 0 0 120 799
use nand3 nand3_8
timestamp 1386234893
transform 1 0 385 0 1 269
box 0 0 120 799
use inv inv_14
timestamp 1386238110
transform 1 0 505 0 1 269
box 0 0 120 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 625 0 1 269
box 0 0 120 799
use inv inv_15
timestamp 1386238110
transform 1 0 745 0 1 269
box 0 0 120 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 865 0 1 269
box 0 0 120 799
use inv inv_16
timestamp 1386238110
transform 1 0 985 0 1 269
box 0 0 120 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 1105 0 1 269
box 0 0 120 799
use inv inv_17
timestamp 1386238110
transform 1 0 1225 0 1 269
box 0 0 120 799
use nand3 nand3_12
timestamp 1386234893
transform 1 0 1345 0 1 269
box 0 0 120 799
use inv inv_18
timestamp 1386238110
transform 1 0 1465 0 1 269
box 0 0 120 799
use nand3 nand3_13
timestamp 1386234893
transform 1 0 1585 0 1 269
box 0 0 120 799
use inv inv_19
timestamp 1386238110
transform 1 0 1705 0 1 269
box 0 0 120 799
use nand3 nand3_14
timestamp 1386234893
transform 1 0 1825 0 1 269
box 0 0 120 799
use inv inv_20
timestamp 1386238110
transform 1 0 1945 0 1 269
box 0 0 120 799
use nand3 nand3_15
timestamp 1386234893
transform 1 0 2065 0 1 269
box 0 0 120 799
use inv inv_21
timestamp 1386238110
transform 1 0 2185 0 1 269
box 0 0 120 799
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 2305 0 1 269
box 0 0 720 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 3025 0 1 269
box 0 0 720 799
use inv inv_0
timestamp 1386238110
transform 1 0 3745 0 1 269
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 3865 0 1 269
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 3985 0 1 269
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 4105 0 1 269
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 4225 0 1 269
box 0 0 120 799
use nand3 nand3_1
timestamp 1386234893
transform 1 0 4345 0 1 269
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 4465 0 1 269
box 0 0 120 799
use nand3 nand3_2
timestamp 1386234893
transform 1 0 4585 0 1 269
box 0 0 120 799
use inv inv_5
timestamp 1386238110
transform 1 0 4705 0 1 269
box 0 0 120 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 4825 0 1 269
box 0 0 120 799
use inv inv_6
timestamp 1386238110
transform 1 0 4945 0 1 269
box 0 0 120 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 5065 0 1 269
box 0 0 120 799
use inv inv_7
timestamp 1386238110
transform 1 0 5185 0 1 269
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 5305 0 1 269
box 0 0 120 799
use inv inv_8
timestamp 1386238110
transform 1 0 5425 0 1 269
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 5545 0 1 269
box 0 0 120 799
use inv inv_9
timestamp 1386238110
transform 1 0 5665 0 1 269
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 5785 0 1 269
box 0 0 120 799
use inv inv_10
timestamp 1386238110
transform 1 0 5905 0 1 269
box 0 0 120 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 6025 0 1 269
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 6241 0 1 269
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 6457 0 1 269
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 7177 0 1 269
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 7393 0 1 269
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 7609 0 1 269
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 8329 0 1 269
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 8545 0 1 269
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 8761 0 1 269
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 9481 0 1 269
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 9697 0 1 269
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 9913 0 1 269
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 10633 0 1 269
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 10849 0 1 269
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 11065 0 1 269
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 11785 0 1 269
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 12001 0 1 269
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 12217 0 1 269
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 12937 0 1 269
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 13153 0 1 269
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 13369 0 1 269
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 14089 0 1 269
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 14305 0 1 269
box 0 0 216 799
use inv inv_22
timestamp 1386238110
transform 1 0 14521 0 1 269
box 0 0 120 799
use inv inv_23
timestamp 1386238110
transform 1 0 14641 0 1 269
box 0 0 120 799
use inv inv_24
timestamp 1386238110
transform 1 0 14761 0 1 269
box 0 0 120 799
use nand3 nand3_16
timestamp 1386234893
transform 1 0 14881 0 1 269
box 0 0 120 799
use inv inv_25
timestamp 1386238110
transform 1 0 15001 0 1 269
box 0 0 120 799
use nand3 nand3_17
timestamp 1386234893
transform 1 0 15121 0 1 269
box 0 0 120 799
use inv inv_26
timestamp 1386238110
transform 1 0 15241 0 1 269
box 0 0 120 799
use nand3 nand3_18
timestamp 1386234893
transform 1 0 15361 0 1 269
box 0 0 120 799
use inv inv_27
timestamp 1386238110
transform 1 0 15481 0 1 269
box 0 0 120 799
use nand3 nand3_19
timestamp 1386234893
transform 1 0 15601 0 1 269
box 0 0 120 799
use inv inv_28
timestamp 1386238110
transform 1 0 15721 0 1 269
box 0 0 120 799
use nand3 nand3_20
timestamp 1386234893
transform 1 0 15841 0 1 269
box 0 0 120 799
use inv inv_29
timestamp 1386238110
transform 1 0 15961 0 1 269
box 0 0 120 799
use nand3 nand3_21
timestamp 1386234893
transform 1 0 16081 0 1 269
box 0 0 120 799
use inv inv_30
timestamp 1386238110
transform 1 0 16201 0 1 269
box 0 0 120 799
use nand3 nand3_22
timestamp 1386234893
transform 1 0 16321 0 1 269
box 0 0 120 799
use inv inv_31
timestamp 1386238110
transform 1 0 16441 0 1 269
box 0 0 120 799
use nand3 nand3_23
timestamp 1386234893
transform 1 0 16561 0 1 269
box 0 0 120 799
use inv inv_32
timestamp 1386238110
transform 1 0 16681 0 1 269
box 0 0 120 799
<< labels >>
rlabel metal2 49 1895 61 1895 5 Rs2[0]
rlabel metal2 169 1895 181 1895 5 Rs2[1]
rlabel metal2 289 1895 301 1895 5 Rs2[2]
rlabel metal2 3769 1895 3781 1895 5 Rs1[0]
rlabel metal2 3889 1895 3901 1895 5 Rs1[1]
rlabel metal2 4009 1895 4021 1895 5 Rs1[2]
rlabel metal2 3119 1895 3131 1895 5 WData[0]
rlabel metal1 0 75 0 85 3 Databus
rlabel metal1 0 40 0 50 3 Rd1[0]
rlabel metal1 0 5 0 15 3 Rd2[0]
rlabel metal1 0 990 0 1015 3 Vdd!
rlabel metal1 0 345 0 370 3 GND!
rlabel metal1 0 322 0 332 3 Clock
rlabel metal1 0 276 0 286 3 nReset
rlabel metal1 16815 345 16815 370 7 GND!
rlabel metal1 16815 322 16815 332 7 Clock
rlabel metal1 16815 276 16815 286 7 nReset
rlabel metal1 16815 75 16815 85 7 Databus
rlabel metal1 16815 40 16815 50 7 Rd1[0]
rlabel metal1 16815 5 16815 15 7 Rd2[0]
rlabel metal1 16815 990 16815 1015 7 Vdd!
rlabel metal2 14545 1895 14557 1895 5 Rw[0]
rlabel metal2 14665 1895 14677 1895 5 Rw[1]
rlabel metal2 14785 1895 14797 1895 5 Rw[2]
rlabel metal2 2377 1895 2389 1895 5 We
<< end >>
