../../../Design/Implementation/verilog/behavioural/decoder.sv