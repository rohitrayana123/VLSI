magic
tech c035u
timestamp 1394310524
<< pwell >>
rect 1332 16954 1386 16979
rect 1332 15875 1386 15900
rect 1332 14796 1386 14821
rect 1332 13717 1386 13742
rect 1332 12638 1386 12663
rect 1332 11559 1386 11584
rect 1332 10480 1386 10505
rect 1332 9401 1386 9426
rect 1332 8322 1386 8347
rect 1332 7243 1386 7268
rect 1332 6164 1386 6189
rect 1332 5085 1386 5110
rect 1332 4006 1386 4031
rect 1332 2927 1386 2952
rect 1332 1848 1386 1873
rect 1332 769 1386 794
<< metal1 >>
rect 1332 17660 1386 17670
rect 1332 17637 1386 17647
rect 1332 17599 1386 17624
rect 1332 16954 1386 16979
rect 1332 16931 1386 16941
rect 1332 16908 1386 16918
rect 1332 16885 1386 16895
rect 1332 16862 1386 16872
rect 1332 16802 1386 16812
rect 2394 16780 2423 16790
rect 1332 16581 1386 16591
rect 1332 16558 1386 16568
rect 1332 16520 1386 16545
rect 1332 15875 1386 15900
rect 1332 15852 1386 15862
rect 1332 15829 1386 15839
rect 1332 15806 1386 15816
rect 1332 15783 1386 15793
rect 1332 15723 1386 15733
rect 2394 15701 2423 15711
rect 1332 15502 1386 15512
rect 1332 15479 1386 15489
rect 1332 15441 1386 15466
rect 1332 14796 1386 14821
rect 1332 14773 1386 14783
rect 1332 14750 1386 14760
rect 1332 14727 1386 14737
rect 1332 14704 1386 14714
rect 1332 14644 1386 14654
rect 2394 14622 2423 14632
rect 1332 14423 1386 14433
rect 1332 14400 1386 14410
rect 1332 14362 1386 14387
rect 1332 13717 1386 13742
rect 1332 13694 1386 13704
rect 1332 13671 1386 13681
rect 1332 13648 1386 13658
rect 1332 13625 1386 13635
rect 1332 13565 1386 13575
rect 2394 13543 2423 13553
rect 1332 13344 1386 13354
rect 1332 13321 1386 13331
rect 1332 13283 1386 13308
rect 1332 12638 1386 12663
rect 1332 12615 1386 12625
rect 1332 12592 1386 12602
rect 1332 12569 1386 12579
rect 1332 12546 1386 12556
rect 1332 12486 1386 12496
rect 2394 12464 2423 12474
rect 1332 12265 1386 12275
rect 1332 12242 1386 12252
rect 1332 12204 1386 12229
rect 1332 11559 1386 11584
rect 1332 11536 1386 11546
rect 1332 11513 1386 11523
rect 1332 11490 1386 11500
rect 1332 11467 1386 11477
rect 1332 11407 1386 11417
rect 2394 11385 2423 11395
rect 1332 11186 1386 11196
rect 1332 11163 1386 11173
rect 1332 11125 1386 11150
rect 1332 10480 1386 10505
rect 1332 10457 1386 10467
rect 1332 10434 1386 10444
rect 1332 10411 1386 10421
rect 1332 10388 1386 10398
rect 1332 10328 1386 10338
rect 2394 10306 2423 10316
rect 1332 10107 1386 10117
rect 1332 10084 1386 10094
rect 1332 10046 1386 10071
rect 1332 9401 1386 9426
rect 1332 9378 1386 9388
rect 1332 9355 1386 9365
rect 1332 9332 1386 9342
rect 1332 9309 1386 9319
rect 1332 9249 1386 9259
rect 2394 9227 2423 9237
rect 1332 9028 1386 9038
rect 1332 9005 1386 9015
rect 1332 8967 1386 8992
rect 1332 8322 1386 8347
rect 1332 8299 1386 8309
rect 1332 8276 1386 8286
rect 1332 8253 1386 8263
rect 1332 8230 1386 8240
rect 1332 8170 1386 8180
rect 2394 8148 2423 8158
rect 1332 7949 1386 7959
rect 1332 7926 1386 7936
rect 1332 7888 1386 7913
rect 1332 7243 1386 7268
rect 1332 7220 1386 7230
rect 1332 7197 1386 7207
rect 1332 7174 1386 7184
rect 1332 7151 1386 7161
rect 1332 7091 1386 7101
rect 2394 7069 2423 7079
rect 1332 6870 1386 6880
rect 1332 6847 1386 6857
rect 1332 6809 1386 6834
rect 1332 6164 1386 6189
rect 1332 6141 1386 6151
rect 1332 6118 1386 6128
rect 1332 6095 1386 6105
rect 1332 6072 1386 6082
rect 1332 6012 1386 6022
rect 2394 5990 2423 6000
rect 1332 5791 1386 5801
rect 1332 5768 1386 5778
rect 1332 5730 1386 5755
rect 1332 5085 1386 5110
rect 1332 5062 1386 5072
rect 1332 5039 1386 5049
rect 1332 5016 1386 5026
rect 1332 4993 1386 5003
rect 1332 4933 1386 4943
rect 2394 4911 2423 4921
rect 1332 4712 1386 4722
rect 1332 4689 1386 4699
rect 1332 4651 1386 4676
rect 1332 4006 1386 4031
rect 1332 3983 1386 3993
rect 1332 3960 1386 3970
rect 1332 3937 1386 3947
rect 1332 3914 1386 3924
rect 1332 3854 1386 3864
rect 2394 3832 2423 3842
rect 1332 3633 1386 3643
rect 1332 3610 1386 3620
rect 1332 3572 1386 3597
rect 1332 2927 1386 2952
rect 1332 2904 1386 2914
rect 1332 2881 1386 2891
rect 1332 2858 1386 2868
rect 1332 2835 1386 2845
rect 1332 2775 1386 2785
rect 2394 2753 2423 2763
rect 1332 2554 1386 2564
rect 1332 2531 1386 2541
rect 1332 2493 1386 2518
rect 1332 1848 1386 1873
rect 1332 1825 1386 1835
rect 1332 1802 1386 1812
rect 1332 1779 1386 1789
rect 1332 1756 1386 1766
rect 1332 1696 1386 1706
rect 2394 1674 2423 1684
rect 1332 1475 1386 1485
rect 1332 1452 1386 1462
rect 1332 1414 1386 1439
rect 1332 769 1386 794
rect 1332 746 1386 756
rect 1332 723 1386 733
rect 1332 700 1386 710
rect 1332 677 1386 687
rect 1332 617 1386 627
rect 2394 595 2423 605
use IrAA  IrAA_0
array 0 0 1008 0 7 1079
timestamp 1394309515
transform 1 0 1386 0 1 9154
box 0 0 1008 1079
use IrBA  IrBA_0
array 0 0 1008 0 2 1079
timestamp 1394309607
transform 1 0 1386 0 1 5917
box 0 0 1008 1079
use IrBB  IrBB_0
array 0 0 1008 0 4 1079
timestamp 1394309685
transform 1 0 1386 0 1 633
box 0 -111 1008 968
<< labels >>
rlabel metal1 1332 617 1332 627 3 SysBus[0]
rlabel metal1 1332 1696 1332 1706 3 SysBus[1]
rlabel metal1 1332 2775 1332 2785 3 SysBus[2]
rlabel metal1 1332 3854 1332 3864 3 SysBus[3]
rlabel metal1 1332 4933 1332 4943 3 SysBus[4]
rlabel metal1 1332 6012 1332 6022 3 SysBus[5]
rlabel metal1 1332 7091 1332 7101 3 SysBus[6]
rlabel metal1 1332 8170 1332 8180 3 SysBus[7]
rlabel metal1 1332 9249 1332 9259 3 SysBus[8]
rlabel metal1 1332 10328 1332 10338 3 SysBus[9]
rlabel metal1 1332 11407 1332 11417 3 SysBus[10]
rlabel metal1 1332 12486 1332 12496 3 SysBus[11]
rlabel metal1 1332 13565 1332 13575 3 SysBus[12]
rlabel metal1 1332 14644 1332 14654 3 SysBus[13]
rlabel metal1 1332 15723 1332 15733 3 SysBus[14]
rlabel metal1 1332 16802 1332 16812 3 SysBus[15]
rlabel metal1 1332 677 1332 687 3 Ir[0]
rlabel metal1 1332 1756 1332 1766 3 Ir[1]
rlabel metal1 1332 2835 1332 2845 3 Ir[2]
rlabel metal1 1332 3914 1332 3924 3 Ir[3]
rlabel metal1 1332 4993 1332 5003 3 Ir[4]
rlabel metal1 1332 6072 1332 6082 3 Ir[5]
rlabel metal1 1332 7151 1332 7161 3 Ir[6]
rlabel metal1 1332 8230 1332 8240 3 Ir[7]
rlabel metal1 1332 9309 1332 9319 3 Ir[8]
rlabel metal1 1332 10388 1332 10398 3 Ir[9]
rlabel metal1 1332 11467 1332 11477 3 Ir[10]
rlabel metal1 1332 12546 1332 12556 3 Ir[11]
rlabel metal1 1332 13625 1332 13635 3 Ir[12]
rlabel metal1 1332 14704 1332 14714 3 Ir[13]
rlabel metal1 1332 15783 1332 15793 3 Ir[14]
rlabel metal1 1332 16862 1332 16872 3 Ir[15]
rlabel metal1 1332 700 1332 710 3 nReset
rlabel metal1 1332 1779 1332 1789 3 nReset
rlabel metal1 1332 2858 1332 2868 3 nReset
rlabel metal1 1332 3937 1332 3947 3 nReset
rlabel metal1 1332 5016 1332 5026 3 nReset
rlabel metal1 1332 6095 1332 6105 3 nReset
rlabel metal1 1332 7174 1332 7184 3 nReset
rlabel metal1 1332 8253 1332 8263 3 nReset
rlabel metal1 1332 9332 1332 9342 3 nReset
rlabel metal1 1332 10411 1332 10421 3 nReset
rlabel metal1 1332 11490 1332 11500 3 nReset
rlabel metal1 1332 12569 1332 12579 3 nReset
rlabel metal1 1332 13648 1332 13658 3 nReset
rlabel metal1 1332 14727 1332 14737 3 nReset
rlabel metal1 1332 15806 1332 15816 3 nReset
rlabel metal1 1332 16885 1332 16895 3 nReset
rlabel metal1 1332 723 1332 733 3 Test
rlabel metal1 1332 1802 1332 1812 3 Test
rlabel metal1 1332 2881 1332 2891 3 Test
rlabel metal1 1332 3960 1332 3970 3 Test
rlabel metal1 1332 5039 1332 5049 3 Test
rlabel metal1 1332 6118 1332 6128 3 Test
rlabel metal1 1332 7197 1332 7207 3 Test
rlabel metal1 1332 8276 1332 8286 3 Test
rlabel metal1 1332 9355 1332 9365 3 Test
rlabel metal1 1332 10434 1332 10444 3 Test
rlabel metal1 1332 11513 1332 11523 3 Test
rlabel metal1 1332 12592 1332 12602 3 Test
rlabel metal1 1332 13671 1332 13681 3 Test
rlabel metal1 1332 14750 1332 14760 3 Test
rlabel metal1 1332 15829 1332 15839 3 Test
rlabel metal1 1332 16908 1332 16918 3 Test
rlabel metal1 1332 746 1332 756 3 Clock
rlabel metal1 1332 1825 1332 1835 3 Clock
rlabel metal1 1332 2904 1332 2914 3 Clock
rlabel metal1 1332 3983 1332 3993 3 Clock
rlabel metal1 1332 5062 1332 5072 3 Clock
rlabel metal1 1332 6141 1332 6151 3 Clock
rlabel metal1 1332 7220 1332 7230 3 Clock
rlabel metal1 1332 8299 1332 8309 3 Clock
rlabel metal1 1332 9378 1332 9388 3 Clock
rlabel metal1 1332 10457 1332 10467 3 Clock
rlabel metal1 1332 11536 1332 11546 3 Clock
rlabel metal1 1332 12615 1332 12625 3 Clock
rlabel metal1 1332 13694 1332 13704 3 Clock
rlabel metal1 1332 14773 1332 14783 3 Clock
rlabel metal1 1332 15852 1332 15862 3 Clock
rlabel metal1 1332 16931 1332 16941 3 Clock
rlabel metal1 1332 769 1332 794 3 GND
rlabel metal1 1332 1848 1332 1873 3 GND
rlabel metal1 1332 2927 1332 2952 3 GND
rlabel metal1 1332 4006 1332 4031 3 GND
rlabel metal1 1332 5085 1332 5110 3 GND
rlabel metal1 1332 6164 1332 6189 3 GND
rlabel metal1 1332 7243 1332 7268 3 GND
rlabel metal1 1332 8322 1332 8347 3 GND
rlabel metal1 1332 9401 1332 9426 3 GND
rlabel metal1 1332 10480 1332 10505 3 GND
rlabel metal1 1332 11559 1332 11584 3 GND
rlabel metal1 1332 12638 1332 12663 3 GND
rlabel metal1 1332 13717 1332 13742 3 GND
rlabel metal1 1332 14796 1332 14821 3 GND
rlabel metal1 1332 15875 1332 15900 3 GND
rlabel metal1 1332 16954 1332 16979 3 GND
rlabel metal1 1332 1414 1332 1439 3 Vdd!
rlabel metal1 1332 2493 1332 2518 3 Vdd!
rlabel metal1 1332 3572 1332 3597 3 Vdd!
rlabel metal1 1332 4651 1332 4676 3 Vdd!
rlabel metal1 1332 5730 1332 5755 3 Vdd!
rlabel metal1 1332 6809 1332 6834 3 Vdd!
rlabel metal1 1332 7888 1332 7913 3 Vdd!
rlabel metal1 1332 8967 1332 8992 3 Vdd!
rlabel metal1 1332 10046 1332 10071 3 Vdd!
rlabel metal1 1332 11125 1332 11150 3 Vdd!
rlabel metal1 1332 12204 1332 12229 3 Vdd!
rlabel metal1 1332 13283 1332 13308 3 Vdd!
rlabel metal1 1332 14362 1332 14387 3 Vdd!
rlabel metal1 1332 15441 1332 15466 3 Vdd!
rlabel metal1 1332 16520 1332 16545 3 Vdd!
rlabel metal1 1332 17599 1332 17624 3 Vdd!
rlabel metal1 1332 1452 1332 1462 3 SDI
rlabel metal1 1332 2531 1332 2541 3 SDI
rlabel metal1 1332 3610 1332 3620 3 SDI
rlabel metal1 1332 4689 1332 4699 3 SDI
rlabel metal1 1332 5768 1332 5778 3 SDI
rlabel metal1 1332 6847 1332 6857 3 SDI
rlabel metal1 1332 7926 1332 7936 3 SDI
rlabel metal1 1332 9005 1332 9015 3 SDI
rlabel metal1 1332 10084 1332 10094 3 SDI
rlabel metal1 1332 11163 1332 11173 3 SDI
rlabel metal1 1332 12242 1332 12252 3 SDI
rlabel metal1 1332 13321 1332 13331 3 SDI
rlabel metal1 1332 14400 1332 14410 3 SDI
rlabel metal1 1332 15479 1332 15489 3 SDI
rlabel metal1 1332 16558 1332 16568 3 SDI
rlabel metal1 1332 17637 1332 17647 3 SDI
rlabel metal1 1332 1475 1332 1485 3 ScanReturn
rlabel metal1 1332 2554 1332 2564 3 ScanReturn
rlabel metal1 1332 3633 1332 3643 3 ScanReturn
rlabel metal1 1332 4712 1332 4722 3 ScanReturn
rlabel metal1 1332 5791 1332 5801 3 ScanReturn
rlabel metal1 1332 6870 1332 6880 3 ScanReturn
rlabel metal1 1332 7949 1332 7959 3 ScanReturn
rlabel metal1 1332 9028 1332 9038 3 ScanReturn
rlabel metal1 1332 10107 1332 10117 3 ScanReturn
rlabel metal1 1332 11186 1332 11196 3 ScanReturn
rlabel metal1 1332 12265 1332 12275 3 ScanReturn
rlabel metal1 1332 13344 1332 13354 3 ScanReturn
rlabel metal1 1332 14423 1332 14433 3 ScanReturn
rlabel metal1 1332 15502 1332 15512 3 ScanReturn
rlabel metal1 1332 16581 1332 16591 3 ScanReturn
rlabel metal1 1332 17660 1332 17670 3 ScanReturn
rlabel metal1 2423 595 2423 605 7 Imm[0]
rlabel metal1 2423 1674 2423 1684 7 Imm[1]
rlabel metal1 2423 2753 2423 2763 7 Imm[2]
rlabel metal1 2423 3832 2423 3842 7 Imm[3]
rlabel metal1 2423 4911 2423 4921 7 Imm[4]
rlabel metal1 2423 5990 2423 6000 7 Imm[5]
rlabel metal1 2423 7069 2423 7079 7 Imm[6]
rlabel metal1 2423 8148 2423 8158 7 Imm[7]
rlabel metal1 2423 9227 2423 9237 7 Imm[8]
rlabel metal1 2423 10306 2423 10316 7 Imm[9]
rlabel metal1 2423 11385 2423 11395 7 Imm[10]
rlabel metal1 2423 12464 2423 12474 7 Imm[11]
rlabel metal1 2423 13543 2423 13553 7 Imm[12]
rlabel metal1 2423 14622 2423 14632 7 Imm[13]
rlabel metal1 2423 15701 2423 15711 7 Imm[14]
rlabel metal1 2423 16780 2423 16790 7 Imm[15]
<< end >>
