magic
tech c035u
timestamp 1394107240
<< metal1 >>
rect 0 1001 73 1011
rect 88 1001 1225 1011
rect 1239 1001 2377 1011
rect 2392 1001 3529 1011
rect 3543 1001 4681 1011
rect 4695 1001 5833 1011
rect 5847 1001 6984 1011
rect 6999 1001 8137 1011
rect 664 964 793 974
rect 807 964 1009 974
rect 1814 951 1945 961
rect 1959 951 2161 961
rect 2966 951 3097 961
rect 3111 951 3313 961
rect 4118 951 4249 961
rect 4263 951 4465 961
rect 5270 951 5401 961
rect 5415 951 5617 961
rect 6422 951 6553 961
rect 6567 951 6769 961
rect 7574 951 7705 961
rect 7719 951 7921 961
rect 8726 951 8857 961
rect 8871 951 9073 961
rect 0 908 50 918
rect 9266 908 9385 918
rect 0 885 50 895
rect 9266 885 9385 895
rect 9266 847 9385 872
rect 0 202 50 227
rect 9266 202 9385 227
rect 0 179 50 189
rect 9266 179 9385 189
rect 0 156 50 166
rect 9266 156 9385 166
rect 0 133 50 143
rect 9266 133 9385 143
rect 0 40 936 50
rect 951 40 2088 50
rect 2103 40 3240 50
rect 3255 40 4393 50
rect 4408 40 5543 50
rect 5561 40 6695 50
rect 6713 40 7847 50
rect 7865 40 9001 50
rect 9015 40 9385 50
rect 0 5 1153 15
rect 1167 5 2305 15
rect 2319 5 3457 15
rect 3471 5 4609 15
rect 4624 5 5760 15
rect 5778 5 6912 15
rect 6930 5 8064 15
rect 8082 5 9217 15
rect 9231 5 9385 15
<< m2contact >>
rect 73 998 88 1014
rect 1225 1000 1239 1014
rect 2377 1000 2392 1014
rect 3529 1000 3543 1014
rect 4681 1000 4695 1014
rect 5833 1000 5847 1014
rect 6984 999 6999 1013
rect 8137 1000 8152 1015
rect 649 963 664 977
rect 793 962 807 976
rect 1009 961 1023 975
rect 1800 949 1814 963
rect 1945 948 1959 962
rect 2161 949 2175 963
rect 2952 949 2966 963
rect 3097 948 3111 962
rect 3313 949 3327 963
rect 4104 949 4118 963
rect 4249 948 4263 962
rect 4465 949 4479 963
rect 5256 949 5270 963
rect 5401 948 5415 962
rect 5617 949 5631 963
rect 6408 949 6422 963
rect 6553 948 6567 962
rect 6769 949 6783 963
rect 7560 949 7574 963
rect 7705 948 7719 962
rect 7921 949 7935 963
rect 8712 949 8726 963
rect 8857 948 8871 962
rect 9073 949 9087 963
rect 936 38 951 52
rect 2088 38 2103 52
rect 3240 38 3255 52
rect 4393 38 4408 53
rect 5543 38 5561 53
rect 6695 38 6713 53
rect 7847 38 7865 53
rect 9001 37 9015 52
rect 1153 4 1167 18
rect 2305 4 2319 18
rect 3457 4 3471 18
rect 4609 3 4624 18
rect 5760 0 5778 15
rect 6912 0 6930 15
rect 8064 0 8082 15
rect 9217 3 9231 18
<< metal2 >>
rect 74 925 86 998
rect 122 925 134 1177
rect 650 925 662 963
rect 794 925 806 962
rect 866 925 878 1177
rect 1010 925 1022 961
rect 1082 925 1094 1177
rect 1226 925 1238 1000
rect 1274 925 1286 1177
rect 1802 925 1814 949
rect 1946 925 1958 948
rect 2018 925 2030 1177
rect 2162 925 2174 949
rect 2234 925 2246 1177
rect 2378 925 2390 1000
rect 2426 925 2438 1177
rect 2954 925 2966 949
rect 3098 925 3110 948
rect 3170 925 3182 1177
rect 3314 925 3326 949
rect 3386 925 3398 1177
rect 3530 925 3542 1000
rect 3578 925 3590 1177
rect 4106 925 4118 949
rect 4250 925 4262 948
rect 4322 925 4334 1177
rect 4466 925 4478 949
rect 4538 925 4550 1177
rect 4682 925 4694 1000
rect 4730 925 4742 1177
rect 5258 925 5270 949
rect 5402 925 5414 948
rect 5474 925 5486 1177
rect 5618 925 5630 949
rect 5690 925 5702 1177
rect 5834 925 5846 1000
rect 5882 925 5894 1177
rect 6410 925 6422 949
rect 6554 925 6566 948
rect 6626 925 6638 1177
rect 6770 925 6782 949
rect 6842 925 6854 1177
rect 6986 925 6998 999
rect 7034 925 7046 1177
rect 7562 925 7574 949
rect 7706 925 7718 948
rect 7778 925 7790 1177
rect 7922 925 7934 949
rect 7994 925 8006 1177
rect 8138 925 8150 1000
rect 8186 925 8198 1177
rect 8714 925 8726 949
rect 8858 925 8870 948
rect 8930 925 8942 1177
rect 9074 925 9086 949
rect 9146 925 9158 1177
rect 938 52 950 126
rect 1154 18 1166 126
rect 2090 52 2102 126
rect 2306 18 2318 126
rect 3242 52 3254 126
rect 3458 18 3470 126
rect 4394 53 4406 126
rect 4610 18 4622 126
rect 5546 53 5558 126
rect 5762 15 5774 126
rect 6698 53 6710 126
rect 6914 15 6926 126
rect 7850 53 7862 126
rect 8066 15 8078 126
rect 9002 52 9014 126
rect 9218 18 9230 126
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 50 0 1 126
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 770 0 1 126
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 986 0 1 126
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 1202 0 1 126
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1922 0 1 126
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2138 0 1 126
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 2354 0 1 126
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3074 0 1 126
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3290 0 1 126
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 3506 0 1 126
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4226 0 1 126
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 4442 0 1 126
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 4658 0 1 126
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 5378 0 1 126
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 5594 0 1 126
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 5810 0 1 126
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 6530 0 1 126
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 6746 0 1 126
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 6962 0 1 126
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 7682 0 1 126
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 7898 0 1 126
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 8114 0 1 126
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 8834 0 1 126
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9050 0 1 126
box 0 0 216 799
<< labels >>
rlabel metal2 122 1177 134 1177 5 Rw[0]
rlabel metal2 866 1177 878 1177 5 Rs1[0]
rlabel metal2 1082 1177 1094 1177 5 Rs2[0]
rlabel metal2 1274 1177 1286 1177 5 Rw[1]
rlabel metal2 2018 1177 2030 1177 5 Rs1[1]
rlabel metal2 2234 1177 2246 1177 5 Rs2[1]
rlabel metal2 2426 1177 2438 1177 5 Rw[2]
rlabel metal2 3170 1177 3182 1177 5 Rs1[2]
rlabel metal2 3386 1177 3398 1177 5 Rs2[2]
rlabel metal2 3578 1177 3590 1177 5 Rw[3]
rlabel metal2 4322 1177 4334 1177 5 Rs1[3]
rlabel metal2 4538 1177 4550 1177 5 Rs2[3]
rlabel metal2 4730 1177 4742 1177 5 Rw[4]
rlabel metal2 5474 1177 5486 1177 5 Rs1[4]
rlabel metal2 5690 1177 5702 1177 5 Rs2[4]
rlabel metal2 5882 1177 5894 1177 5 Rw[5]
rlabel metal2 6626 1177 6638 1177 5 Rs1[5]
rlabel metal2 6842 1177 6854 1177 5 Rs2[5]
rlabel metal2 7034 1177 7046 1177 5 Rw[6]
rlabel metal2 7778 1177 7790 1177 5 Rs1[6]
rlabel metal2 7994 1177 8006 1177 5 Rs2[6]
rlabel metal2 8186 1177 8198 1177 5 Rsw[7]
rlabel metal2 8930 1177 8942 1177 5 Rs1[7]
rlabel metal2 9146 1177 9158 1177 5 Rs2[7]
rlabel metal1 0 1001 0 1011 1 WData
rlabel metal1 0 40 0 50 3 Rd1
rlabel metal1 0 5 0 15 3 Rd2
rlabel metal1 9385 203 9385 227 7 GND!
rlabel metal1 9385 179 9385 189 7 Clock
rlabel metal1 9385 156 9385 166 7 Test
rlabel metal1 9385 133 9385 143 7 nReset
rlabel metal1 9385 847 9385 872 7 Vdd!
rlabel metal1 9385 908 9385 918 7 ScanReturn
rlabel metal1 9385 885 9385 895 7 Scan
rlabel metal1 9385 40 9385 50 7 Rd1
rlabel metal1 9385 5 9385 15 7 Rd2
rlabel metal1 0 908 0 918 3 ScanReturn
rlabel metal1 0 885 0 895 3 SDI
rlabel metal1 0 133 0 143 3 nReset
rlabel metal1 0 156 0 166 3 Test
rlabel metal1 0 179 0 189 3 Clock
rlabel metal1 0 202 0 227 3 GND!
<< end >>
