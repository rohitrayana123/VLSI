magic
tech c035u
timestamp 1395690245
<< metal1 >>
rect 1573 1159 3215 1169
rect 3229 1159 20472 1169
rect 12552 1030 12623 1040
rect 12552 1008 12863 1018
rect 12901 1009 13055 1019
rect 13141 1003 13176 1013
rect 12709 981 13176 991
rect 12973 149 13103 159
rect 0 95 3095 105
rect 3109 95 3263 105
rect 3277 95 20472 105
rect 0 73 12815 83
rect 2821 51 12671 61
rect 0 29 20472 39
<< m2contact >>
rect 1559 1157 1573 1171
rect 3215 1157 3229 1171
rect 12623 1028 12637 1042
rect 12863 1006 12877 1020
rect 12887 1005 12901 1019
rect 13055 1007 13069 1021
rect 13127 1001 13141 1015
rect 12695 979 12709 993
rect 12959 145 12973 159
rect 13103 147 13117 161
rect 3095 93 3109 107
rect 3263 93 3277 107
rect 12815 71 12829 85
rect 2807 49 2821 63
rect 12671 49 12685 63
<< metal2 >>
rect 216 1153 228 1176
rect 360 1153 372 1176
rect 576 1153 588 1176
rect 1320 1153 1332 1176
rect 1488 1153 1500 1176
rect 1560 1153 1572 1157
rect 1872 1153 1884 1176
rect 2064 1153 2076 1176
rect 2280 1153 2292 1176
rect 3024 1153 3036 1176
rect 3192 976 3204 1176
rect 3216 976 3228 1157
rect 3288 1153 3372 1165
rect 3408 1153 3420 1176
rect 4152 1153 4164 1176
rect 4368 1153 4380 1176
rect 4560 1153 4572 1176
rect 5304 1153 5316 1176
rect 5520 1153 5532 1176
rect 5712 1153 5724 1176
rect 6456 1153 6468 1176
rect 6672 1153 6684 1176
rect 6864 1153 6876 1176
rect 7608 1153 7620 1176
rect 7824 1153 7836 1176
rect 8016 1153 8028 1176
rect 8760 1153 8772 1176
rect 8976 1153 8988 1176
rect 9168 1153 9180 1176
rect 9912 1153 9924 1176
rect 10128 1153 10140 1176
rect 10320 1153 10332 1176
rect 11064 1153 11076 1176
rect 11280 1153 11292 1176
rect 11472 1153 11484 1176
rect 12216 1153 12228 1176
rect 12432 1153 12444 1176
rect 3288 976 3300 1153
rect 12600 976 12612 1176
rect 12624 976 12636 1028
rect 12696 976 12708 979
rect 12792 976 12804 1176
rect 12864 976 12876 1006
rect 12888 976 12900 1005
rect 13032 976 13044 1176
rect 13248 1153 13260 1176
rect 13512 1153 13524 1176
rect 13680 1153 13692 1176
rect 13848 1153 13860 1176
rect 13872 1153 13884 1176
rect 13944 1153 13956 1176
rect 14160 1153 14172 1176
rect 14304 1153 14316 1176
rect 14640 1153 14652 1176
rect 15000 1153 15012 1176
rect 15408 1153 15420 1176
rect 15744 1153 15756 1176
rect 16056 1153 16068 1176
rect 16392 1153 16404 1176
rect 16512 1153 16524 1176
rect 16560 1153 16572 1176
rect 16728 1153 16740 1176
rect 16824 1153 16836 1176
rect 16872 1153 16884 1176
rect 16920 1153 16932 1176
rect 16968 1153 16980 1176
rect 17016 1153 17028 1176
rect 17064 1153 17076 1176
rect 17112 1153 17124 1176
rect 17160 1153 17172 1176
rect 17472 1153 17484 1176
rect 17520 1153 17532 1176
rect 17568 1153 17580 1176
rect 17616 1153 17628 1176
rect 17928 1153 17940 1176
rect 17976 1153 17988 1176
rect 18360 1153 18372 1176
rect 18528 1153 18540 1176
rect 18553 1153 18565 1176
rect 18600 1153 18612 1176
rect 18648 1153 18660 1176
rect 18696 1153 18708 1176
rect 18744 1153 18756 1176
rect 18792 1153 18804 1176
rect 18840 1153 18852 1176
rect 18888 1153 18900 1176
rect 18936 1153 18948 1176
rect 19176 1153 19188 1176
rect 19248 1153 19260 1176
rect 19296 1153 19308 1176
rect 19344 1153 19356 1176
rect 19392 1153 19404 1176
rect 19632 1153 19644 1176
rect 19704 1153 19716 1176
rect 19752 1153 19764 1176
rect 19992 1153 20004 1176
rect 20064 1153 20076 1176
rect 20352 1153 20364 1176
rect 13056 976 13068 1007
rect 13128 976 13140 1001
rect 216 0 228 111
rect 360 0 372 111
rect 576 0 588 111
rect 1320 0 1332 111
rect 1488 0 1500 111
rect 1872 0 1884 111
rect 2064 0 2076 111
rect 2280 0 2292 111
rect 2808 63 2820 111
rect 3024 0 3036 111
rect 3096 107 3108 111
rect 3192 0 3204 177
rect 3264 107 3276 177
rect 3408 0 3420 111
rect 4152 0 4164 111
rect 4368 0 4380 111
rect 4560 0 4572 111
rect 5304 0 5316 111
rect 5520 0 5532 111
rect 5712 0 5724 111
rect 6456 0 6468 111
rect 6672 0 6684 111
rect 6864 0 6876 111
rect 7608 0 7620 111
rect 7824 0 7836 111
rect 8016 0 8028 111
rect 8760 0 8772 111
rect 8976 0 8988 111
rect 9168 0 9180 111
rect 9912 0 9924 111
rect 10128 0 10140 111
rect 10320 0 10332 111
rect 11064 0 11076 111
rect 11280 0 11292 111
rect 11472 0 11484 111
rect 12216 0 12228 111
rect 12432 0 12444 111
rect 12600 0 12612 177
rect 12672 63 12684 177
rect 12792 0 12804 177
rect 12816 85 12828 177
rect 12960 159 12972 177
rect 13032 0 13044 177
rect 13104 161 13116 177
rect 13248 0 13260 111
rect 13512 0 13524 111
rect 13680 0 13692 111
rect 13872 0 13884 111
rect 14160 0 14172 111
rect 14304 0 14316 111
rect 14640 0 14652 111
rect 15000 0 15012 111
rect 15408 0 15420 111
rect 15744 0 15756 111
rect 16056 0 16068 111
rect 16392 0 16404 111
rect 16560 0 16572 111
rect 16728 0 16740 111
rect 16824 0 16836 111
rect 16872 0 16884 111
rect 16920 0 16932 111
rect 16968 0 16980 111
rect 17016 0 17028 111
rect 17064 0 17076 111
rect 17112 0 17124 111
rect 17160 0 17172 111
rect 17472 0 17484 111
rect 17520 0 17532 111
rect 17568 0 17580 111
rect 17616 0 17628 111
rect 17928 0 17940 111
rect 17976 0 17988 111
rect 18360 0 18372 111
rect 18528 0 18540 111
rect 18553 0 18565 111
rect 18600 0 18612 111
rect 18648 0 18660 111
rect 18696 0 18708 111
rect 18744 0 18756 111
rect 18792 0 18804 111
rect 18840 0 18852 111
rect 18888 0 18900 111
rect 18936 0 18948 111
rect 19176 0 19188 111
rect 19248 0 19260 111
rect 19296 0 19308 111
rect 19344 0 19356 111
rect 19392 0 19404 111
rect 19632 0 19644 111
rect 19704 0 19716 111
rect 19752 0 19764 111
rect 19992 0 20004 111
rect 20064 0 20076 111
rect 20352 0 20364 111
use Pc_slice Pc_slice_0
timestamp 1394724028
transform 1 0 0 0 1 111
box 0 0 3144 1042
use mux2 mux2_0
timestamp 1386235218
transform 1 0 3144 0 1 177
box 0 0 192 799
use regBlock_slice regBlock_slice_0
timestamp 1395689161
transform 1 0 3336 0 1 111
box 0 0 9216 1042
use mux2 mux2_1
timestamp 1386235218
transform 1 0 12552 0 1 177
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 12744 0 1 177
box 0 0 192 799
use tielow tielow_0
timestamp 1386086605
transform 1 0 12936 0 1 177
box 0 0 48 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 12984 0 1 177
box 0 0 192 799
use ALUSlice ALUSlice_0
timestamp 1394559926
transform 1 0 13176 0 1 111
box 0 0 7296 1042
<< labels >>
rlabel metal2 12792 1176 12804 1176 5 Op2Sel[0]
rlabel metal2 13032 1176 13044 1176 5 Op2Sel[1]
rlabel metal1 13163 1007 13163 1007 1 B
rlabel metal2 13032 0 13044 0 1 Op2Sel[1]
rlabel metal2 20064 1176 20076 1176 5 Sh1_R_in
rlabel metal2 16824 1176 16836 1176 5 Sh8Z_L
rlabel metal2 17160 1176 17172 1176 5 Sh8G_L
rlabel metal2 17064 1176 17076 1176 5 Sh8E_L
rlabel metal2 17112 1176 17124 1176 5 Sh8F_L
rlabel metal2 16920 1176 16932 1176 5 Sh8B_L
rlabel metal2 17016 1176 17028 1176 5 Sh8D_L
rlabel metal2 16968 1176 16980 1176 5 Sh8C_L
rlabel metal2 16872 1176 16884 1176 5 Sh8A_L
rlabel metal1 20472 95 20472 105 7 SysBus
rlabel metal1 20472 1159 20472 1169 7 AluOut
rlabel metal2 16512 1176 16524 1176 5 A
rlabel metal2 18360 1176 18372 1176 5 Sh1_L_Out
rlabel metal2 18528 1176 18540 1176 5 Sh8
rlabel metal2 18696 1176 18708 1176 5 Sh8C_R
rlabel metal2 18648 1176 18660 1176 5 Sh8B_R
rlabel metal2 18600 1176 18612 1176 5 Sh8A_R
rlabel metal2 17616 1176 17628 1176 5 Sh4C_L
rlabel metal2 17568 1176 17580 1176 5 Sh4B_L
rlabel metal2 17976 1176 17988 1176 5 Sh2B_L
rlabel metal2 17928 1176 17940 1176 5 Sh2A_L
rlabel metal2 18553 1176 18565 1176 5 ShR
rlabel metal2 17520 1176 17532 1176 5 Sh4A_L
rlabel metal2 17472 1176 17484 1176 5 Sh4Z_L
rlabel metal2 19248 1176 19260 1176 5 Sh4Z_R
rlabel metal2 19992 1176 20004 1176 5 Sh1
rlabel metal2 19632 1176 19644 1176 5 Sh2
rlabel metal2 20352 1176 20364 1176 5 ShOut
rlabel metal2 19752 1176 19764 1176 5 Sh2B_R
rlabel metal2 19704 1176 19716 1176 5 Sh2A_R
rlabel metal2 19392 1176 19404 1176 5 Sh4C_R
rlabel metal2 19344 1176 19356 1176 5 Sh4B_R
rlabel metal2 19296 1176 19308 1176 5 Sh4A_R
rlabel metal2 19176 1176 19188 1176 5 Sh4
rlabel metal2 18744 1176 18756 1176 5 Sh8D_R
rlabel metal2 18792 1176 18804 1176 5 Sh8E_R
rlabel metal2 18840 1176 18852 1176 5 Sh8F_R
rlabel metal2 18888 1176 18900 1176 5 Sh8G_R
rlabel metal2 18936 1176 18948 1176 5 Sh8H_R
rlabel metal2 13248 1176 13260 1176 5 ZeroA
rlabel metal2 13680 1176 13692 1176 5 CIn
rlabel metal2 13944 1176 13956 1176 5 Sum
rlabel metal2 13872 1176 13884 1176 5 COut
rlabel metal2 16560 1176 16572 1176 5 ShB
rlabel metal2 16392 1176 16404 1176 5 NOR
rlabel metal2 16056 1176 16068 1176 5 NAND
rlabel metal2 15744 1176 15756 1176 5 NOT
rlabel metal2 15408 1176 15420 1176 5 XOR
rlabel metal2 15000 1176 15012 1176 5 OR
rlabel metal2 14640 1176 14652 1176 5 AND
rlabel metal2 13512 1176 13524 1176 5 SUB
rlabel metal2 14160 1176 14172 1176 5 nZ
rlabel metal2 14304 1176 14316 1176 5 FAOut
rlabel metal2 16728 1176 16740 1176 5 ShL
rlabel metal2 13848 1176 13860 1176 5 CIn_Slice
rlabel metal2 17112 0 17124 0 1 Sh8G_L
rlabel metal2 17064 0 17076 0 1 Sh8F_L
rlabel metal2 17016 0 17028 0 1 Sh8E_L
rlabel metal2 16968 0 16980 0 1 Sh8D_L
rlabel metal2 18360 0 18372 0 1 Sh1_L_In
rlabel metal2 18600 0 18612 0 1 Sh8Z_R
rlabel metal2 18648 0 18660 0 1 Sh8A_R
rlabel metal2 18696 0 18708 0 1 Sh8B_R
rlabel metal2 17616 0 17628 0 1 Sh4D_L
rlabel metal2 17568 0 17580 0 1 Sh4C_L
rlabel metal2 17520 0 17532 0 1 Sh4B_L
rlabel metal2 17976 0 17988 0 1 Sh2C_L
rlabel metal2 17928 0 17940 0 1 Sh2B_L
rlabel metal2 18553 0 18565 0 1 ShR
rlabel metal2 18528 0 18540 0 1 Sh8
rlabel metal2 17472 0 17484 0 1 Sh4A_L
rlabel metal2 17160 0 17172 0 1 Sh8H_L
rlabel metal2 19248 0 19260 0 1 Sh4Y_L
rlabel metal2 20064 0 20076 0 1 Sh1_R_Out
rlabel metal2 19752 0 19764 0 1 Sh2A_R
rlabel metal2 19704 0 19716 0 1 Sh2Z_R
rlabel metal2 19296 0 19308 0 1 Sh4Z_R
rlabel metal2 19344 0 19356 0 1 Sh4A_R
rlabel metal2 19392 0 19404 0 1 Sh4B_R
rlabel metal2 20352 0 20364 0 1 ShOut
rlabel metal2 19632 0 19644 0 1 Sh2
rlabel metal2 19992 0 20004 0 1 Sh1
rlabel metal2 19176 0 19188 0 1 Sh4
rlabel metal2 18744 0 18756 0 1 Sh8C_R
rlabel metal2 18792 0 18804 0 1 Sh8D_R
rlabel metal2 18840 0 18852 0 1 Sh8E_R
rlabel metal2 18888 0 18900 0 1 Sh8F_R
rlabel metal2 18936 0 18948 0 1 Sh8G_R
rlabel metal2 16824 0 16836 0 1 Sh8A_L
rlabel metal2 16920 0 16932 0 1 Sh8C_L
rlabel metal2 16872 0 16884 0 1 Sh8B_L
rlabel metal2 13248 0 13260 0 1 ZeroA
rlabel metal2 14304 0 14316 0 1 FAOut
rlabel metal2 13680 0 13692 0 1 CIn
rlabel metal2 14640 0 14652 0 1 AND
rlabel metal2 15000 0 15012 0 1 OR
rlabel metal2 15408 0 15420 0 1 XOR
rlabel metal2 15744 0 15756 0 1 NOT
rlabel metal2 16056 0 16068 0 1 NAND
rlabel metal2 16392 0 16404 0 1 NOR
rlabel metal2 16728 0 16740 0 1 ShL
rlabel metal2 16560 0 16572 0 1 ShB
rlabel metal2 13512 0 13524 0 1 SUB
rlabel metal2 14160 0 14172 0 1 nZ_prev
rlabel metal2 13872 0 13884 0 1 CIn_Slice
rlabel metal2 12792 0 12804 0 1 Op2Sel[0]
rlabel metal1 12815 987 12815 987 1 A
rlabel metal1 12942 1164 12942 1164 6 AluOut
rlabel metal2 12600 1176 12612 1176 5 Op1Sel
rlabel metal1 12925 99 12925 99 1 SysBus
rlabel metal2 12600 0 12612 0 1 Op1Sel
rlabel metal2 3192 1176 3204 1176 5 WdSel
rlabel metal2 3408 1176 3420 1176 5 Rw[0]
rlabel metal2 4152 1176 4164 1176 5 Rs1[0]
rlabel metal2 4368 1176 4380 1176 5 Rs2[0]
rlabel metal2 4560 1176 4572 1176 5 Rw[1]
rlabel metal2 5304 1176 5316 1176 5 Rs1[1]
rlabel metal2 5520 1176 5532 1176 5 Rs2[1]
rlabel metal2 5712 1176 5724 1176 5 Rw[2]
rlabel metal2 6456 1176 6468 1176 5 Rs1[2]
rlabel metal2 6672 1176 6684 1176 5 Rs2[2]
rlabel metal2 6864 1176 6876 1176 5 Rw[3]
rlabel metal2 7608 1176 7620 1176 5 Rs1[3]
rlabel metal2 7824 1176 7836 1176 5 Rs2[3]
rlabel metal2 8016 1176 8028 1176 5 Rw[4]
rlabel metal2 8760 1176 8772 1176 5 Rs1[4]
rlabel metal2 8976 1176 8988 1176 5 Rs2[4]
rlabel metal2 9168 1176 9180 1176 5 Rw[5]
rlabel metal2 10128 1176 10140 1176 5 Rs2[5]
rlabel metal2 9912 1176 9924 1176 5 Rs1[5]
rlabel metal2 10320 1176 10332 1176 5 Rw[6]
rlabel metal2 11064 1176 11076 1176 5 Rs1[6]
rlabel metal2 11280 1176 11292 1176 5 Rs2[6]
rlabel metal2 11472 1176 11484 1176 5 Rw[7]
rlabel metal2 12216 1176 12228 1176 5 Rs1[7]
rlabel metal2 12432 1176 12444 1176 5 Rs2[7]
rlabel metal2 4368 0 4380 0 1 Rs2[0]
rlabel metal2 3408 0 3420 0 1 Rw[0]
rlabel metal1 12546 56 12546 56 1 Pc
rlabel metal1 12545 78 12545 78 1 Imm
rlabel metal1 12544 100 12544 100 1 SysBus
rlabel metal2 12432 0 12444 0 1 Rs2[7]
rlabel metal2 12216 0 12228 0 1 Rs1[7]
rlabel metal2 11472 0 11484 0 1 Rw[7]
rlabel metal2 11280 0 11292 0 1 Rs2[6]
rlabel metal2 11064 0 11076 0 1 Rs1[6]
rlabel metal2 10320 0 10332 0 1 Rw[6]
rlabel metal2 10128 0 10140 0 1 Rs2[5]
rlabel metal2 9912 0 9924 0 1 Rs1[5]
rlabel metal2 9168 0 9180 0 1 Rw[5]
rlabel metal2 8976 0 8988 0 1 Rs2[4]
rlabel metal2 8760 0 8772 0 1 Rs1[4]
rlabel metal2 8016 0 8028 0 1 Rw[4]
rlabel metal2 7824 0 7836 0 1 Rs2[3]
rlabel metal2 7608 0 7620 0 1 Rs1[3]
rlabel metal2 6864 0 6876 0 1 Rw[3]
rlabel metal2 6672 0 6684 0 1 Rs2[2]
rlabel metal2 6456 0 6468 0 1 Rs1[2]
rlabel metal2 5712 0 5724 0 1 Rw[2]
rlabel metal2 5520 0 5532 0 1 Rs2[1]
rlabel metal2 5304 0 5316 0 1 Rs1[1]
rlabel metal2 4560 0 4572 0 1 Rw[1]
rlabel metal2 4152 0 4164 0 1 Rs1[0]
rlabel metal2 3192 0 3204 0 1 WdSel
rlabel metal1 3288 100 3288 100 1 SysBus
rlabel metal2 3024 1176 3036 1176 5 PcEn
rlabel metal2 3024 0 3036 0 1 PcEn
rlabel metal2 2280 0 2292 0 1 PcWe
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 1872 1176 1884 1176 5 PcSel[1]
rlabel metal2 1488 1176 1500 1176 5 PcSel[0]
rlabel metal2 1320 1176 1332 1176 5 LrEn
rlabel metal2 576 1176 588 1176 5 LrWe
rlabel metal2 360 1176 372 1176 5 LrSel
rlabel metal2 216 1176 228 1176 5 PcIncCout
rlabel metal2 2280 1176 2292 1176 5 PcWe
rlabel metal1 0 95 0 105 1 SysBus
rlabel metal1 0 73 0 83 1 Imm
rlabel metal2 2064 0 2076 0 1 PcSel[2]
rlabel metal2 2064 1176 2076 1176 5 PcSel[2]
rlabel metal1 0 29 0 39 3 DataIn
rlabel metal1 20472 29 20472 39 7 DataIn
rlabel metal1 12577 1035 12577 1035 1 Rd1
rlabel metal1 12579 1013 12579 1013 1 Rd2
<< end >>
