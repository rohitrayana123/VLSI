magic
tech c035u
timestamp 1394109793
<< metal1 >>
rect -10 875 71 885
rect 85 875 311 885
rect 325 875 431 885
rect 445 875 671 885
rect 685 875 887 885
rect 901 875 1127 885
rect 1141 875 1343 885
rect 1357 875 1679 885
rect -10 853 47 863
rect 61 853 191 863
rect 205 853 551 863
rect 565 853 647 863
rect 661 853 863 863
rect 877 853 1223 863
rect 1237 853 1319 863
rect 1333 853 1559 863
rect 1573 853 1693 863
rect -10 830 23 840
rect 37 830 167 840
rect 181 830 407 840
rect 421 830 767 840
rect 781 830 1007 840
rect 1021 830 1103 840
rect 1117 830 1439 840
rect 1453 830 1535 840
rect 1549 830 1693 840
rect -10 782 0 792
rect -10 759 0 769
rect -10 721 0 746
rect -10 53 0 63
rect -10 30 0 40
rect -10 7 0 17
<< m2contact >>
rect 71 873 85 887
rect 311 873 325 887
rect 431 873 445 887
rect 671 873 685 887
rect 887 873 901 887
rect 1127 873 1141 887
rect 1343 873 1357 887
rect 1679 873 1693 887
rect 47 851 61 865
rect 191 851 205 865
rect 551 851 565 865
rect 647 851 661 865
rect 863 851 877 865
rect 1223 851 1237 865
rect 1319 851 1333 865
rect 1559 851 1573 865
rect 23 828 37 842
rect 167 828 181 842
rect 407 828 421 842
rect 767 828 781 842
rect 1007 828 1021 842
rect 1103 828 1117 842
rect 1439 828 1453 842
rect 1535 828 1549 842
<< metal2 >>
rect 24 799 36 828
rect 48 799 60 851
rect 72 799 84 873
rect 168 799 180 828
rect 192 799 204 851
rect 312 799 324 873
rect 408 799 420 828
rect 432 799 444 873
rect 552 799 564 851
rect 648 799 660 851
rect 672 799 684 873
rect 768 799 780 828
rect 864 799 876 851
rect 888 799 900 873
rect 1008 799 1020 828
rect 1104 799 1116 828
rect 1128 799 1140 873
rect 1224 799 1236 851
rect 1320 799 1332 851
rect 1344 799 1356 873
rect 1440 799 1452 828
rect 1536 799 1548 828
rect 1560 799 1572 851
rect 1680 799 1692 873
rect 120 -45 132 0
rect 240 -12 300 0
rect 360 -45 372 0
rect 480 -12 540 0
rect 600 -45 612 0
rect 696 -12 756 0
rect 816 -45 828 0
rect 936 -12 996 0
rect 1056 -45 1068 0
rect 1152 -12 1212 0
rect 1272 -45 1284 0
rect 1368 -12 1428 0
rect 1488 -45 1500 0
rect 1608 -12 1668 0
rect 1728 -45 1740 0
use nor3 nor3_0
timestamp 1386235396
transform 1 0 0 0 1 0
box 0 0 144 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 144 0 1 0
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 264 0 1 0
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 384 0 1 0
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 504 0 1 0
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 624 0 1 0
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 720 0 1 0
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 840 0 1 0
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 960 0 1 0
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1080 0 1 0
box 0 0 96 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 1176 0 1 0
box 0 0 120 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 1296 0 1 0
box 0 0 96 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 1392 0 1 0
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 1512 0 1 0
box 0 0 120 799
use and2 and2_4
timestamp 1386234845
transform 1 0 1632 0 1 0
box 0 0 120 799
<< labels >>
rlabel metal2 120 -45 132 -45 1 Out[0]
rlabel metal2 360 -45 372 -45 1 Out[1]
rlabel metal2 600 -45 612 -45 1 Out[2]
rlabel metal2 816 -45 828 -45 1 Out[3]
rlabel metal2 1056 -45 1068 -45 1 Out[4]
rlabel metal2 1272 -45 1284 -45 1 Out[5]
rlabel metal2 1488 -45 1500 -45 1 Out[6]
rlabel metal2 1728 -45 1740 -45 1 Out[7]
rlabel metal1 -10 830 -10 840 3 In[0]
rlabel metal1 -10 853 -10 863 3 In[1]
rlabel metal1 -10 875 -10 885 4 In[2]
rlabel metal1 -10 782 -10 792 3 ScanReturn
rlabel metal1 -10 759 -10 769 3 Scan
rlabel metal1 -10 721 -10 746 3 Vdd!
rlabel metal1 -10 7 -10 17 3 nReset
rlabel metal1 -10 30 -10 40 3 Test
rlabel metal1 -10 53 -10 63 3 Clock
<< end >>
