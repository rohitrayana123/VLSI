magic
tech c035u
timestamp 1394708291
<< metal1 >>
rect 37 894 1175 904
rect 1189 894 2327 904
rect 2342 894 3479 904
rect 3493 894 4631 904
rect 4645 894 5783 904
rect 5797 894 6934 904
rect 6949 894 8087 904
rect 614 871 743 881
rect 757 871 959 881
rect 1764 871 1895 881
rect 1909 871 2111 881
rect 2916 871 3047 881
rect 3061 871 3263 881
rect 4068 870 4199 880
rect 4213 870 4415 880
rect 5221 870 5351 880
rect 5365 870 5567 880
rect 6372 870 6503 880
rect 6517 870 6719 880
rect 7524 870 7655 880
rect 7669 870 7871 880
rect 8677 871 8807 881
rect 8821 871 9023 881
rect 901 50 2038 60
rect 2053 50 3190 60
rect 3205 50 4343 60
rect 4358 50 5493 60
rect 5511 50 6645 60
rect 6663 50 7797 60
rect 7815 50 8951 60
rect 1117 27 2255 37
rect 2269 27 3407 37
rect 3421 27 4559 37
rect 4574 27 5710 37
rect 5728 27 6862 37
rect 6880 27 8014 37
rect 8032 27 9167 37
<< m2contact >>
rect 23 892 37 906
rect 1175 893 1189 907
rect 2327 893 2342 907
rect 3479 893 3493 907
rect 4631 893 4645 907
rect 5783 893 5797 907
rect 6934 892 6949 906
rect 8087 892 8101 906
rect 599 870 614 884
rect 743 869 757 883
rect 959 868 973 882
rect 1750 869 1764 883
rect 1895 868 1909 882
rect 2111 869 2125 883
rect 2902 869 2916 883
rect 3047 868 3061 882
rect 3263 869 3277 883
rect 4054 868 4068 882
rect 4199 868 4213 882
rect 4415 868 4429 882
rect 5207 868 5221 882
rect 5351 868 5365 882
rect 5567 868 5581 882
rect 6358 868 6372 882
rect 6503 868 6517 882
rect 6719 868 6733 882
rect 7510 868 7524 882
rect 7655 868 7669 882
rect 7871 868 7885 882
rect 8663 869 8677 883
rect 8807 868 8821 882
rect 9023 869 9037 883
rect 886 48 901 62
rect 2038 48 2053 62
rect 3190 48 3205 62
rect 4343 48 4358 63
rect 5493 48 5511 63
rect 6645 48 6663 63
rect 7797 48 7815 63
rect 8951 47 8965 62
rect 1103 26 1117 40
rect 2255 26 2269 40
rect 3407 26 3421 40
rect 4559 25 4574 40
rect 5710 22 5728 37
rect 6862 22 6880 37
rect 8014 22 8032 37
rect 9167 25 9181 40
<< metal2 >>
rect 24 906 36 1042
rect 24 865 36 892
rect 72 865 84 1042
rect 600 865 612 870
rect 744 865 756 869
rect 816 865 828 1042
rect 960 865 972 868
rect 1032 865 1044 1042
rect 1176 865 1188 893
rect 1224 865 1236 1042
rect 1752 865 1764 869
rect 1896 865 1908 868
rect 1968 865 1980 1042
rect 2112 865 2124 869
rect 2184 865 2196 1042
rect 2328 865 2340 893
rect 2376 865 2388 1042
rect 2904 865 2916 869
rect 3048 865 3060 868
rect 3120 865 3132 1042
rect 3264 865 3276 869
rect 3336 865 3348 1042
rect 3480 865 3492 893
rect 3528 865 3540 1042
rect 4056 865 4068 868
rect 4200 865 4212 868
rect 4272 865 4284 1042
rect 4416 865 4428 868
rect 4488 865 4500 1042
rect 4632 865 4644 893
rect 4680 865 4692 1042
rect 5208 865 5220 868
rect 5352 865 5364 868
rect 5424 865 5436 1042
rect 5568 865 5580 868
rect 5640 865 5652 1042
rect 5784 865 5796 893
rect 5832 865 5844 1042
rect 6360 865 6372 868
rect 6504 865 6516 868
rect 6576 865 6588 1042
rect 6720 865 6732 868
rect 6792 865 6804 1042
rect 6936 865 6948 892
rect 6984 865 6996 1042
rect 7512 865 7524 868
rect 7656 865 7668 868
rect 7728 865 7740 1042
rect 7872 865 7884 868
rect 7944 865 7956 1042
rect 8088 865 8100 892
rect 8136 865 8148 1042
rect 8664 865 8676 869
rect 8808 865 8820 868
rect 8880 865 8892 1042
rect 9024 865 9036 869
rect 9096 865 9108 1042
rect 72 0 84 66
rect 816 0 828 66
rect 888 62 900 66
rect 1032 0 1044 66
rect 1104 40 1116 66
rect 1224 0 1236 66
rect 1968 0 1980 66
rect 2040 62 2052 66
rect 2184 0 2196 66
rect 2256 40 2268 66
rect 2376 0 2388 66
rect 3120 0 3132 66
rect 3192 62 3204 66
rect 3336 0 3348 66
rect 3408 40 3420 66
rect 3528 0 3540 66
rect 4272 0 4284 66
rect 4344 63 4356 66
rect 4488 0 4500 66
rect 4560 40 4572 66
rect 4680 0 4692 66
rect 5424 0 5436 66
rect 5496 63 5508 66
rect 5640 0 5652 66
rect 5712 37 5724 66
rect 5832 0 5844 66
rect 6576 0 6588 66
rect 6648 63 6660 66
rect 6792 0 6804 66
rect 6864 37 6876 66
rect 6984 0 6996 66
rect 7728 0 7740 66
rect 7800 63 7812 66
rect 7944 0 7956 66
rect 8016 37 8028 66
rect 8136 0 8148 66
rect 8880 0 8892 66
rect 8952 62 8964 66
rect 8952 0 8964 47
rect 9096 0 9108 66
rect 9168 40 9180 66
rect 9168 0 9180 25
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 66
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 720 0 1 66
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 936 0 1 66
box 0 0 216 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 1152 0 1 66
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1872 0 1 66
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2088 0 1 66
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 2304 0 1 66
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3024 0 1 66
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3240 0 1 66
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 3456 0 1 66
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4176 0 1 66
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 4392 0 1 66
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 4608 0 1 66
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 5328 0 1 66
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 5544 0 1 66
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 5760 0 1 66
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 6480 0 1 66
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 6696 0 1 66
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 6912 0 1 66
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 7632 0 1 66
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 7848 0 1 66
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 8064 0 1 66
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 8784 0 1 66
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9000 0 1 66
box 0 0 216 799
<< labels >>
rlabel metal2 72 0 84 0 1 Rw[0]
rlabel metal2 1032 0 1044 0 5 Rs2[0]
rlabel metal2 1224 0 1236 0 5 Rw[1]
rlabel metal2 1968 0 1980 0 5 Rs1[1]
rlabel metal2 3120 0 3132 0 5 Rs1[2]
rlabel metal2 3528 0 3540 0 5 Rw[3]
rlabel metal2 3336 0 3348 0 5 Rs2[2]
rlabel metal2 4272 0 4284 0 5 Rs1[3]
rlabel metal2 4680 0 4692 0 5 Rw[4]
rlabel metal2 4488 0 4500 0 5 Rs2[3]
rlabel metal2 5424 0 5436 0 5 Rs1[4]
rlabel metal2 2376 0 2388 0 1 Rw[2]
rlabel metal2 5640 0 5652 0 1 Rs2[4]
rlabel metal2 7728 0 7740 0 5 Rs1[6]
rlabel metal2 9096 0 9108 0 5 Rs2[7]
rlabel metal2 8880 0 8892 0 5 Rs1[7]
rlabel metal2 8136 0 8148 0 5 Rw[7]
rlabel metal2 7944 0 7956 0 5 Rs2[6]
rlabel metal2 6984 0 6996 0 5 Rw[6]
rlabel metal2 6792 0 6804 0 5 Rs2[5]
rlabel metal2 6576 0 6588 0 5 Rs1[5]
rlabel metal2 5832 0 5844 0 5 Rw[5]
rlabel metal2 2184 0 2196 0 1 Rs2[1]
rlabel metal2 816 0 828 0 1 Rs1[0]
rlabel metal2 8952 0 8964 0 1 Rd1
rlabel metal2 9168 0 9180 0 1 Rd2
rlabel metal2 5424 1042 5436 1042 5 Rs1[4]
rlabel metal2 4680 1042 4692 1042 5 Rw[4]
rlabel metal2 4488 1042 4500 1042 5 Rs2[3]
rlabel metal2 4272 1042 4284 1042 5 Rs1[3]
rlabel metal2 3528 1042 3540 1042 5 Rw[3]
rlabel metal2 3336 1042 3348 1042 5 Rs2[2]
rlabel metal2 3120 1042 3132 1042 5 Rs1[2]
rlabel metal2 2376 1042 2388 1042 5 Rw[2]
rlabel metal2 2184 1042 2196 1042 5 Rs2[1]
rlabel metal2 1968 1042 1980 1042 5 Rs1[1]
rlabel metal2 1224 1042 1236 1042 5 Rw[1]
rlabel metal2 1032 1042 1044 1042 5 Rs2[0]
rlabel metal2 816 1042 828 1042 5 Rs1[0]
rlabel metal2 5640 1042 5652 1042 5 Rs2[4]
rlabel metal2 5832 1042 5844 1042 5 Rw[5]
rlabel metal2 6576 1042 6588 1042 5 Rs1[5]
rlabel metal2 6792 1042 6804 1042 5 Rs2[5]
rlabel metal2 6984 1042 6996 1042 5 Rw[6]
rlabel metal2 7728 1042 7740 1042 5 Rs1[6]
rlabel metal2 7944 1042 7956 1042 5 Rs2[6]
rlabel metal2 8880 1042 8892 1042 5 Rs1[7]
rlabel metal2 9096 1042 9108 1042 5 Rs2[7]
rlabel metal2 8136 1042 8148 1042 5 Rw[7]
rlabel metal2 72 1042 84 1042 5 Rw[0]
rlabel metal2 24 1042 36 1042 5 WData
rlabel metal1 692 873 692 873 1 Reg0
rlabel metal1 1814 875 1814 875 1 Reg1
rlabel metal1 3107 876 3107 876 1 Reg2
rlabel metal1 4349 873 4349 873 1 Reg3
rlabel metal1 5402 874 5402 874 1 Reg4
rlabel metal1 6613 873 6613 873 1 Reg5
rlabel metal1 7783 875 7783 875 1 Reg6
rlabel metal1 8970 877 8970 877 1 Reg7Out
<< end >>
