magic
tech c035u
timestamp 1395432264
<< metal1 >>
rect 7440 41410 7450 41452
rect 7488 41410 7498 41452
rect 7440 41400 7498 41410
rect 6450 40416 6514 40426
rect 6504 40405 6514 40416
rect 7440 40405 7450 41400
rect 7536 40405 7546 41452
rect 11472 41266 11482 41452
rect 11520 41293 11530 41452
rect 15600 41437 15610 41452
rect 15648 41437 15658 41452
rect 19728 41437 19738 41452
rect 19776 41437 19786 41452
rect 19920 41437 19930 41452
rect 27984 41437 27994 41452
rect 28032 41437 28042 41452
rect 28176 41410 28186 41452
rect 32112 41437 32122 41452
rect 32160 41437 32170 41452
rect 11629 41400 28186 41410
rect 32304 41410 32314 41452
rect 36240 41437 36250 41452
rect 36288 41413 36298 41452
rect 36432 41437 36442 41452
rect 28213 41400 32314 41410
rect 32341 41400 36263 41410
rect 36312 41400 36778 41410
rect 11592 41376 28031 41386
rect 11592 41338 11602 41376
rect 28069 41376 32111 41386
rect 32125 41376 36239 41386
rect 36312 41386 36322 41400
rect 36253 41376 36322 41386
rect 36336 41376 36431 41386
rect 11640 41352 15647 41362
rect 11640 41341 11650 41352
rect 15685 41352 36287 41362
rect 36336 41362 36346 41376
rect 36768 41386 36778 41400
rect 36768 41376 36802 41386
rect 36312 41352 36346 41362
rect 36624 41352 36778 41362
rect 11568 41328 11602 41338
rect 11568 41293 11578 41328
rect 11677 41328 32159 41338
rect 32184 41328 32327 41338
rect 32184 41314 32194 41328
rect 36312 41338 36322 41352
rect 36277 41328 36322 41338
rect 11592 41304 32194 41314
rect 11592 41293 11602 41304
rect 11701 41280 19775 41290
rect 19813 41280 28199 41290
rect 11472 41256 15599 41266
rect 11520 40405 11530 41231
rect 11544 40378 11554 41256
rect 15637 41256 19727 41266
rect 19741 41256 27983 41266
rect 27997 41256 28055 41266
rect 11712 41232 19919 41242
rect 6450 40368 11554 40378
rect 6504 35722 6514 40343
rect 6528 35749 6538 40368
rect 7440 39082 7450 40343
rect 7536 39109 7546 40343
rect 11520 39301 11530 40343
rect 11568 39274 11578 41231
rect 11592 39277 11602 41231
rect 11616 39277 11626 41231
rect 11640 39277 11650 41231
rect 11664 39277 11674 41231
rect 11688 39277 11698 41231
rect 11712 39277 11722 41232
rect 11736 41208 19799 41218
rect 11736 39277 11746 41208
rect 11760 41184 15671 41194
rect 11760 39277 11770 41184
rect 11784 41160 15623 41170
rect 11784 39277 11794 41160
rect 11485 39264 11578 39274
rect 11437 39240 11818 39250
rect 11389 39216 11591 39226
rect 11808 39226 11818 39240
rect 11808 39216 11866 39226
rect 11365 39192 11831 39202
rect 11856 39202 11866 39216
rect 11856 39192 11890 39202
rect 11304 39168 11866 39178
rect 11304 39157 11314 39168
rect 11341 39144 11818 39154
rect 11280 39120 11471 39130
rect 11280 39109 11290 39120
rect 11509 39120 11783 39130
rect 11808 39109 11818 39144
rect 11413 39096 11783 39106
rect 11832 39106 11842 39143
rect 11856 39133 11866 39168
rect 11880 39154 11890 39192
rect 15600 39181 15610 41135
rect 27253 39240 29122 39250
rect 26533 39216 29087 39226
rect 29112 39226 29122 39240
rect 29112 39216 29290 39226
rect 26269 39192 29255 39202
rect 29280 39202 29290 39216
rect 29280 39192 29399 39202
rect 36624 39181 36634 41352
rect 18277 39168 29471 39178
rect 36768 39178 36778 41352
rect 36792 40642 36802 41376
rect 36792 40632 41538 40642
rect 41472 40621 41482 40632
rect 41448 40584 41538 40594
rect 41448 40477 41458 40584
rect 41472 40477 41482 40559
rect 41424 40440 41538 40450
rect 36768 39168 36802 39178
rect 36792 39157 36802 39168
rect 11880 39144 36778 39154
rect 17245 39120 29351 39130
rect 29389 39120 29423 39130
rect 29461 39120 36647 39130
rect 36768 39130 36778 39144
rect 36768 39120 36874 39130
rect 36864 39109 36874 39120
rect 11832 39096 11879 39106
rect 17053 39096 29063 39106
rect 29101 39096 36839 39106
rect 7440 39072 11831 39082
rect 11869 39072 36887 39082
rect 11448 39048 11855 39058
rect 6504 35712 6562 35722
rect 6450 35688 6514 35698
rect 6504 35677 6514 35688
rect 6528 35650 6538 35687
rect 6450 35640 6538 35650
rect 6504 30997 6514 35615
rect 6528 30994 6538 35640
rect 6552 31021 6562 35712
rect 6528 30984 6586 30994
rect 6450 30960 6538 30970
rect 6528 30949 6538 30960
rect 6576 30922 6586 30984
rect 6450 30912 6586 30922
rect 6504 26317 6514 30887
rect 6528 26317 6538 30887
rect 6552 26314 6562 30887
rect 6552 26304 6586 26314
rect 6450 26280 6562 26290
rect 6504 21685 6514 26255
rect 6528 21685 6538 26255
rect 6552 21685 6562 26280
rect 6576 21685 6586 26304
rect 6450 21648 6610 21658
rect 6504 16957 6514 21623
rect 6528 16957 6538 21623
rect 6552 16954 6562 21623
rect 6576 16981 6586 21623
rect 6600 18034 6610 21648
rect 7536 18061 7546 39047
rect 11304 39010 11314 39047
rect 11328 39013 11338 39047
rect 11352 39013 11362 39047
rect 11376 39013 11386 39047
rect 11400 39013 11410 39047
rect 11424 39013 11434 39047
rect 11448 39013 11458 39048
rect 11893 39048 11914 39058
rect 11472 39024 11879 39034
rect 11472 39013 11482 39024
rect 11904 39034 11914 39048
rect 16093 39048 29375 39058
rect 29413 39048 36767 39058
rect 36805 39048 36946 39058
rect 11904 39024 36911 39034
rect 36936 39034 36946 39048
rect 36936 39024 36959 39034
rect 11269 39000 11314 39010
rect 41424 39010 41434 40440
rect 11557 39000 41434 39010
rect 11232 38976 11279 38986
rect 11232 38941 11242 38976
rect 11317 38976 12191 38986
rect 15853 38976 29447 38986
rect 29485 38976 36815 38986
rect 36877 38976 36983 38986
rect 11280 38952 11759 38962
rect 11280 38914 11290 38952
rect 11893 38952 12311 38962
rect 15600 38962 15610 38975
rect 15600 38952 29338 38962
rect 11568 38928 11735 38938
rect 11568 38917 11578 38928
rect 11221 38904 11290 38914
rect 11605 38904 11711 38914
rect 11784 38893 11794 38951
rect 11197 38880 11687 38890
rect 11808 38890 11818 38951
rect 11832 38914 11842 38951
rect 11856 38938 11866 38951
rect 11856 38928 29303 38938
rect 29328 38938 29338 38952
rect 29365 38952 36863 38962
rect 36901 38952 37007 38962
rect 29328 38928 36623 38938
rect 36661 38928 36887 38938
rect 36925 38928 37042 38938
rect 37032 38917 37042 38928
rect 11832 38904 12167 38914
rect 12205 38904 29399 38914
rect 29437 38904 36946 38914
rect 36936 38893 36946 38904
rect 11808 38880 29039 38890
rect 29077 38880 36911 38890
rect 37008 38890 37018 38903
rect 37008 38880 37066 38890
rect 37056 38869 37066 38880
rect 11173 38856 11231 38866
rect 11293 38856 37007 38866
rect 11136 38832 11183 38842
rect 11136 36109 11146 38832
rect 41448 38842 41458 40415
rect 11245 38832 41458 38842
rect 11184 38808 11663 38818
rect 11160 36109 11170 38807
rect 11184 36109 11194 38808
rect 11797 38808 12298 38818
rect 12288 38797 12298 38808
rect 12325 38808 29242 38818
rect 29232 38797 29242 38808
rect 29269 38808 36802 38818
rect 11208 36109 11218 38783
rect 11232 36109 11242 38783
rect 11256 36109 11266 38783
rect 11280 36109 11290 38783
rect 11304 36109 11314 38783
rect 11328 36109 11338 38783
rect 11352 36109 11362 38783
rect 11376 36109 11386 38783
rect 11400 36109 11410 38783
rect 11424 36109 11434 38783
rect 11448 36109 11458 38783
rect 11472 36109 11482 38783
rect 11496 36109 11506 38783
rect 11520 36109 11530 38783
rect 11544 36109 11554 38783
rect 11568 36109 11578 38783
rect 11592 36082 11602 38783
rect 11616 36085 11626 38783
rect 11640 36085 11650 38783
rect 11112 36072 11602 36082
rect 11112 36034 11122 36072
rect 11664 36058 11698 36061
rect 11605 36051 11698 36058
rect 11605 36048 11674 36051
rect 11112 36029 11674 36034
rect 11112 36024 11698 36029
rect 11664 36019 11698 36024
rect 11136 35986 11146 35999
rect 11664 35986 11698 35995
rect 11136 35985 11698 35986
rect 11136 35976 11674 35985
rect 11160 34933 11170 35951
rect 11184 34933 11194 35951
rect 11208 34933 11218 35951
rect 11232 34933 11242 35951
rect 11256 34933 11266 35951
rect 11280 34933 11290 35951
rect 11304 34933 11314 35951
rect 11328 34933 11338 35951
rect 11352 34933 11362 35951
rect 11376 34933 11386 35951
rect 11400 34933 11410 35951
rect 11424 34933 11434 35951
rect 11448 34933 11458 35951
rect 11472 34933 11482 35951
rect 11496 34933 11506 35951
rect 11520 34933 11530 35951
rect 11544 34933 11554 35951
rect 11568 34933 11578 35951
rect 11592 34933 11602 35951
rect 11616 34906 11626 35951
rect 11640 34909 11650 35951
rect 11136 34896 11626 34906
rect 11136 34858 11146 34896
rect 11664 34882 11698 34885
rect 11629 34875 11698 34882
rect 11629 34872 11674 34875
rect 11136 34853 11674 34858
rect 11136 34848 11698 34853
rect 11664 34843 11698 34848
rect 11160 34810 11170 34823
rect 11664 34810 11698 34819
rect 11160 34809 11698 34810
rect 11160 34800 11674 34809
rect 11184 33757 11194 34775
rect 11208 33757 11218 34775
rect 11232 33757 11242 34775
rect 11256 33757 11266 34775
rect 11280 33757 11290 34775
rect 11304 33757 11314 34775
rect 11328 33757 11338 34775
rect 11352 33757 11362 34775
rect 11376 33757 11386 34775
rect 11400 33757 11410 34775
rect 11424 33757 11434 34775
rect 11448 33757 11458 34775
rect 11472 33757 11482 34775
rect 11496 33757 11506 34775
rect 11520 33757 11530 34775
rect 11544 33757 11554 34775
rect 11568 33730 11578 34775
rect 11592 33733 11602 34775
rect 11616 33733 11626 34775
rect 11640 33733 11650 34775
rect 11160 33720 11578 33730
rect 11160 33682 11170 33720
rect 11664 33706 11698 33709
rect 11581 33699 11698 33706
rect 11581 33696 11674 33699
rect 11160 33677 11674 33682
rect 11160 33672 11698 33677
rect 11664 33667 11698 33672
rect 11184 33634 11194 33647
rect 11664 33634 11698 33643
rect 11184 33633 11698 33634
rect 11184 33624 11674 33633
rect 11208 32581 11218 33599
rect 11232 32581 11242 33599
rect 11256 32581 11266 33599
rect 11280 32581 11290 33599
rect 11304 32581 11314 33599
rect 11328 32581 11338 33599
rect 11352 32581 11362 33599
rect 11376 32554 11386 33599
rect 11400 32557 11410 33599
rect 11424 32557 11434 33599
rect 11448 32557 11458 33599
rect 11472 32557 11482 33599
rect 11496 32557 11506 33599
rect 11520 32557 11530 33599
rect 11544 32557 11554 33599
rect 11568 32557 11578 33599
rect 11592 32557 11602 33599
rect 11616 32557 11626 33599
rect 11640 32557 11650 33599
rect 11184 32544 11386 32554
rect 11184 32506 11194 32544
rect 11664 32530 11698 32533
rect 11389 32523 11698 32530
rect 11389 32520 11674 32523
rect 11184 32501 11674 32506
rect 11184 32496 11698 32501
rect 11664 32491 11698 32496
rect 11208 32458 11218 32471
rect 11664 32458 11698 32467
rect 11208 32457 11698 32458
rect 11208 32448 11674 32457
rect 11232 31405 11242 32423
rect 11256 31405 11266 32423
rect 11280 31405 11290 32423
rect 11304 31405 11314 32423
rect 11328 31405 11338 32423
rect 11352 31405 11362 32423
rect 11376 31405 11386 32423
rect 11400 31405 11410 32423
rect 11424 31405 11434 32423
rect 11448 31405 11458 32423
rect 11472 31405 11482 32423
rect 11496 31405 11506 32423
rect 11520 31405 11530 32423
rect 11544 31378 11554 32423
rect 11568 31381 11578 32423
rect 11592 31381 11602 32423
rect 11616 31381 11626 32423
rect 11640 31381 11650 32423
rect 11208 31368 11554 31378
rect 11208 31330 11218 31368
rect 11664 31354 11698 31357
rect 11557 31347 11698 31354
rect 11557 31344 11674 31347
rect 11208 31325 11674 31330
rect 11208 31320 11698 31325
rect 11664 31315 11698 31320
rect 11232 31282 11242 31295
rect 11664 31282 11698 31291
rect 11232 31281 11698 31282
rect 11232 31272 11674 31281
rect 11256 30229 11266 31247
rect 11280 30229 11290 31247
rect 11304 30229 11314 31247
rect 11328 30229 11338 31247
rect 11352 30202 11362 31247
rect 11376 30205 11386 31247
rect 11400 30205 11410 31247
rect 11424 30205 11434 31247
rect 11448 30205 11458 31247
rect 11472 30205 11482 31247
rect 11496 30205 11506 31247
rect 11520 30205 11530 31247
rect 11544 30205 11554 31247
rect 11568 30205 11578 31247
rect 11592 30205 11602 31247
rect 11616 30205 11626 31247
rect 11640 30205 11650 31247
rect 11232 30192 11362 30202
rect 11232 30154 11242 30192
rect 11664 30178 11698 30181
rect 11365 30171 11698 30178
rect 11365 30168 11674 30171
rect 11232 30149 11674 30154
rect 11232 30144 11698 30149
rect 11664 30139 11698 30144
rect 11256 30106 11266 30119
rect 11664 30106 11698 30115
rect 11256 30105 11698 30106
rect 11256 30096 11674 30105
rect 11280 29053 11290 30071
rect 11304 29053 11314 30071
rect 11328 29053 11338 30071
rect 11352 29053 11362 30071
rect 11376 29053 11386 30071
rect 11400 29053 11410 30071
rect 11424 29026 11434 30071
rect 11448 29029 11458 30071
rect 11472 29029 11482 30071
rect 11496 29029 11506 30071
rect 11520 29029 11530 30071
rect 11544 29029 11554 30071
rect 11568 29029 11578 30071
rect 11592 29029 11602 30071
rect 11616 29029 11626 30071
rect 11640 29029 11650 30071
rect 11256 29016 11434 29026
rect 11256 28978 11266 29016
rect 11664 29002 11698 29005
rect 11437 28995 11698 29002
rect 11437 28992 11674 28995
rect 11256 28973 11674 28978
rect 11256 28968 11698 28973
rect 11664 28963 11698 28968
rect 11280 28930 11290 28943
rect 11664 28930 11698 28939
rect 11280 28929 11698 28930
rect 11280 28920 11674 28929
rect 11304 27877 11314 28895
rect 11328 27877 11338 28895
rect 11352 27877 11362 28895
rect 11376 27877 11386 28895
rect 11400 27877 11410 28895
rect 11424 27877 11434 28895
rect 11448 27877 11458 28895
rect 11472 27877 11482 28895
rect 11496 27877 11506 28895
rect 11520 27877 11530 28895
rect 11544 27877 11554 28895
rect 11568 27877 11578 28895
rect 11592 27877 11602 28895
rect 11616 27877 11626 28895
rect 11640 27850 11650 28895
rect 11293 27840 11650 27850
rect 11256 27816 11471 27826
rect 11256 27805 11266 27816
rect 11664 27826 11698 27829
rect 11653 27819 11698 27826
rect 11653 27816 11674 27819
rect 11472 27797 11674 27802
rect 11472 27792 11698 27797
rect 11448 27778 11458 27791
rect 11472 27781 11482 27792
rect 11664 27787 11698 27792
rect 11232 27768 11458 27778
rect 11232 26650 11242 27768
rect 11664 27754 11698 27763
rect 11448 27753 11698 27754
rect 11448 27744 11674 27753
rect 11256 26653 11266 27743
rect 11280 26653 11290 27743
rect 11304 26653 11314 27743
rect 11328 26653 11338 27743
rect 11352 26653 11362 27743
rect 11376 26653 11386 27743
rect 11400 26653 11410 27743
rect 11424 26653 11434 27743
rect 11448 26653 11458 27744
rect 11472 26653 11482 27719
rect 11496 26653 11506 27719
rect 11520 26653 11530 27719
rect 11544 26653 11554 27719
rect 11568 26653 11578 27719
rect 11592 26653 11602 27719
rect 11616 26653 11626 27719
rect 11640 26653 11650 27719
rect 11208 26640 11242 26650
rect 11208 26629 11218 26640
rect 11245 26621 11674 26626
rect 11245 26616 11698 26621
rect 11664 26611 11698 26616
rect 11184 26592 11303 26602
rect 11184 25501 11194 26592
rect 11664 26578 11698 26587
rect 11304 26577 11698 26578
rect 11304 26568 11674 26577
rect 11208 25501 11218 26567
rect 11232 25501 11242 26567
rect 11256 25501 11266 26567
rect 11280 25501 11290 26567
rect 11304 25501 11314 26568
rect 11328 25501 11338 26543
rect 11352 25501 11362 26543
rect 11376 25501 11386 26543
rect 11400 25501 11410 26543
rect 11424 25501 11434 26543
rect 11448 25474 11458 26543
rect 11472 25477 11482 26543
rect 11496 25477 11506 26543
rect 11520 25477 11530 26543
rect 11544 25477 11554 26543
rect 11568 25477 11578 26543
rect 11592 25477 11602 26543
rect 11616 25477 11626 26543
rect 11640 25477 11650 26543
rect 11160 25464 11458 25474
rect 11160 25453 11170 25464
rect 11448 25445 11674 25450
rect 11448 25440 11698 25445
rect 11400 25426 11410 25439
rect 11448 25429 11458 25440
rect 11664 25435 11698 25440
rect 11136 25416 11410 25426
rect 11136 24325 11146 25416
rect 11664 25402 11698 25411
rect 11400 25401 11698 25402
rect 11400 25392 11674 25401
rect 11160 24325 11170 25391
rect 11184 24325 11194 25391
rect 11208 24325 11218 25391
rect 11232 24325 11242 25391
rect 11256 24325 11266 25391
rect 11280 24325 11290 25391
rect 11304 24325 11314 25391
rect 11328 24325 11338 25391
rect 11352 24325 11362 25391
rect 11376 24325 11386 25391
rect 11400 24325 11410 25392
rect 11424 24325 11434 25367
rect 11448 24325 11458 25367
rect 11472 24298 11482 25367
rect 11496 24301 11506 25367
rect 11520 24301 11530 25367
rect 11544 24301 11554 25367
rect 11568 24301 11578 25367
rect 11592 24301 11602 25367
rect 11616 24301 11626 25367
rect 11640 24301 11650 25367
rect 11112 24288 11482 24298
rect 11112 24277 11122 24288
rect 11472 24269 11674 24274
rect 11472 24264 11698 24269
rect 11208 24250 11218 24263
rect 11472 24253 11482 24264
rect 11664 24259 11698 24264
rect 11088 24240 11218 24250
rect 11088 23149 11098 24240
rect 11664 24226 11698 24235
rect 11208 24225 11698 24226
rect 11208 24216 11674 24225
rect 11112 23149 11122 24215
rect 11136 23149 11146 24215
rect 11160 23149 11170 24215
rect 11184 23149 11194 24215
rect 11208 23149 11218 24216
rect 11232 23149 11242 24191
rect 11256 23149 11266 24191
rect 11280 23149 11290 24191
rect 11304 23149 11314 24191
rect 11328 23149 11338 24191
rect 11352 23149 11362 24191
rect 11376 23149 11386 24191
rect 11400 23149 11410 24191
rect 11424 23149 11434 24191
rect 11448 23149 11458 24191
rect 11472 23149 11482 24191
rect 11496 23149 11506 24191
rect 11520 23149 11530 24191
rect 11544 23149 11554 24191
rect 11568 23122 11578 24191
rect 11592 23125 11602 24191
rect 11616 23125 11626 24191
rect 11640 23125 11650 24191
rect 11064 23112 11578 23122
rect 11064 23101 11074 23112
rect 11568 23093 11674 23098
rect 11568 23088 11698 23093
rect 11352 23074 11362 23087
rect 11568 23077 11578 23088
rect 11664 23083 11698 23088
rect 11040 23064 11362 23074
rect 11040 21973 11050 23064
rect 11664 23050 11698 23059
rect 11352 23049 11698 23050
rect 11352 23040 11674 23049
rect 11064 21973 11074 23039
rect 11088 21973 11098 23039
rect 11112 21973 11122 23039
rect 11136 21973 11146 23039
rect 11160 21973 11170 23039
rect 11184 21973 11194 23039
rect 11208 21973 11218 23039
rect 11232 21973 11242 23039
rect 11256 21973 11266 23039
rect 11280 21973 11290 23039
rect 11304 21973 11314 23039
rect 11328 21973 11338 23039
rect 11352 21973 11362 23040
rect 11376 21973 11386 23015
rect 11400 21973 11410 23015
rect 11424 21973 11434 23015
rect 11448 21973 11458 23015
rect 11472 21973 11482 23015
rect 11496 21973 11506 23015
rect 11520 21973 11530 23015
rect 11544 21973 11554 23015
rect 11568 21946 11578 23015
rect 11592 21949 11602 23015
rect 11616 21949 11626 23015
rect 11640 21949 11650 23015
rect 11016 21936 11578 21946
rect 11016 21925 11026 21936
rect 11568 21917 11674 21922
rect 11568 21912 11698 21917
rect 11448 21898 11458 21911
rect 11568 21901 11578 21912
rect 11664 21907 11698 21912
rect 10992 21888 11458 21898
rect 10992 20797 11002 21888
rect 11664 21874 11698 21883
rect 11448 21873 11698 21874
rect 11448 21864 11674 21873
rect 11016 20797 11026 21863
rect 11040 20770 11050 21863
rect 11064 20773 11074 21863
rect 11088 20773 11098 21863
rect 11112 20773 11122 21863
rect 11136 20773 11146 21863
rect 11160 20773 11170 21863
rect 11184 20773 11194 21863
rect 11208 20773 11218 21863
rect 11232 20773 11242 21863
rect 11256 20773 11266 21863
rect 11280 20773 11290 21863
rect 11304 20773 11314 21863
rect 11328 20773 11338 21863
rect 11352 20773 11362 21863
rect 11376 20773 11386 21863
rect 11400 20773 11410 21863
rect 11424 20773 11434 21863
rect 11448 20773 11458 21864
rect 11472 20773 11482 21839
rect 11496 20773 11506 21839
rect 11520 20773 11530 21839
rect 11544 20773 11554 21839
rect 11568 20773 11578 21839
rect 11592 20773 11602 21839
rect 11616 20773 11626 21839
rect 11640 20773 11650 21839
rect 10968 20760 11050 20770
rect 10968 20749 10978 20760
rect 11053 20741 11674 20746
rect 11053 20736 11698 20741
rect 11664 20731 11698 20736
rect 10944 20712 11063 20722
rect 10944 19669 10954 20712
rect 11664 20698 11698 20707
rect 11064 20697 11698 20698
rect 11064 20688 11674 20697
rect 10968 19669 10978 20687
rect 10992 19642 11002 20687
rect 11016 19645 11026 20687
rect 11040 19645 11050 20687
rect 11064 19645 11074 20688
rect 11088 19645 11098 20663
rect 11112 19645 11122 20663
rect 11136 19645 11146 20663
rect 11160 19645 11170 20663
rect 11184 19645 11194 20663
rect 11208 19645 11218 20663
rect 11232 19645 11242 20663
rect 11256 19645 11266 20663
rect 11280 19645 11290 20663
rect 11304 19645 11314 20663
rect 11328 19645 11338 20663
rect 11352 19645 11362 20663
rect 11376 19645 11386 20663
rect 11400 19645 11410 20663
rect 11424 19645 11434 20663
rect 11448 19645 11458 20663
rect 11472 19645 11482 20663
rect 11496 19645 11506 20663
rect 10920 19632 11002 19642
rect 10920 19621 10930 19632
rect 11520 19618 11530 20663
rect 11005 19608 11530 19618
rect 11544 19594 11554 20663
rect 11568 19597 11578 20663
rect 11592 19597 11602 20663
rect 11616 19597 11626 20663
rect 11640 19597 11650 20663
rect 10896 19584 11554 19594
rect 10896 19570 10906 19584
rect 10896 19560 11530 19570
rect 11520 19549 11530 19560
rect 11544 19565 11674 19570
rect 11544 19560 11698 19565
rect 11544 19549 11554 19560
rect 11664 19555 11698 19560
rect 10896 19536 11111 19546
rect 10896 18445 10906 19536
rect 11664 19522 11698 19531
rect 11112 19521 11698 19522
rect 11112 19512 11674 19521
rect 10920 18445 10930 19511
rect 10944 18445 10954 19511
rect 10968 18445 10978 19511
rect 10992 18445 11002 19511
rect 11016 18445 11026 19511
rect 11040 18445 11050 19511
rect 11064 18445 11074 19511
rect 11088 18445 11098 19511
rect 11112 18445 11122 19512
rect 11136 18445 11146 19487
rect 11160 18445 11170 19487
rect 11184 18445 11194 19487
rect 11208 18418 11218 19487
rect 11232 18421 11242 19487
rect 11256 18421 11266 19487
rect 11280 18421 11290 19487
rect 11304 18421 11314 19487
rect 11328 18421 11338 19487
rect 11352 18421 11362 19487
rect 11376 18421 11386 19487
rect 11400 18421 11410 19487
rect 11424 18421 11434 19487
rect 11448 18421 11458 19487
rect 11472 18421 11482 19487
rect 11496 18421 11506 19487
rect 11520 18421 11530 19487
rect 11544 18421 11554 19487
rect 11568 18421 11578 19487
rect 11592 18421 11602 19487
rect 11616 18421 11626 19487
rect 11640 18421 11650 19487
rect 10872 18408 11218 18418
rect 10872 18397 10882 18408
rect 11221 18389 11674 18394
rect 11221 18384 11698 18389
rect 11664 18379 11698 18384
rect 10848 18360 11399 18370
rect 10848 18154 10858 18360
rect 11664 18346 11698 18355
rect 11400 18345 11698 18346
rect 11400 18336 11674 18345
rect 10872 18181 10882 18335
rect 10896 18181 10906 18335
rect 10920 18181 10930 18335
rect 10944 18181 10954 18335
rect 10968 18181 10978 18335
rect 10992 18181 11002 18335
rect 11016 18181 11026 18335
rect 11040 18181 11050 18335
rect 11064 18181 11074 18335
rect 11088 18181 11098 18335
rect 11112 18181 11122 18335
rect 11136 18181 11146 18335
rect 11160 18181 11170 18335
rect 11184 18181 11194 18335
rect 11208 18181 11218 18335
rect 11232 18181 11242 18335
rect 11256 18181 11266 18335
rect 11280 18181 11290 18335
rect 11304 18181 11314 18335
rect 11328 18181 11338 18335
rect 11352 18181 11362 18335
rect 11376 18181 11386 18335
rect 11400 18181 11410 18336
rect 11424 18181 11434 18311
rect 11448 18181 11458 18311
rect 11472 18181 11482 18311
rect 11496 18181 11506 18311
rect 11520 18181 11530 18311
rect 11544 18181 11554 18311
rect 11568 18181 11578 18311
rect 11592 18181 11602 18311
rect 11616 18181 11626 18311
rect 11640 18181 11650 18311
rect 36768 18181 36778 38783
rect 36792 18178 36802 38808
rect 36816 18205 36826 38807
rect 36840 18205 36850 38807
rect 36864 18205 36874 38807
rect 36888 18205 36898 38807
rect 36912 18205 36922 38807
rect 36936 18202 36946 38807
rect 36960 26314 36970 38807
rect 36984 30994 36994 38807
rect 37008 31138 37018 38807
rect 37032 35722 37042 38807
rect 37056 35866 37066 38807
rect 41472 35914 41482 40415
rect 41472 35904 41538 35914
rect 41472 35893 41482 35904
rect 37056 35856 41538 35866
rect 41472 35749 41482 35831
rect 37032 35712 41538 35722
rect 41472 31186 41482 35687
rect 41472 31176 41538 31186
rect 41472 31165 41482 31176
rect 37008 31128 41538 31138
rect 41472 31021 41482 31103
rect 36984 30984 41538 30994
rect 41472 26341 41482 30959
rect 36960 26304 41495 26314
rect 36936 18192 36959 18202
rect 36792 18168 36994 18178
rect 10848 18144 36935 18154
rect 36984 18154 36994 18168
rect 36984 18144 37018 18154
rect 37008 18133 37018 18144
rect 10885 18120 36983 18130
rect 10909 18096 36791 18106
rect 36949 18096 37042 18106
rect 10933 18072 36935 18082
rect 37032 18082 37042 18096
rect 37032 18072 37066 18082
rect 10957 18048 37042 18058
rect 37032 18037 37042 18048
rect 6600 18024 12287 18034
rect 13045 18024 36287 18034
rect 37056 18034 37066 18072
rect 37056 18024 37090 18034
rect 10981 18000 37066 18010
rect 6552 16944 6610 16954
rect 6450 16920 6562 16930
rect 6504 12586 6514 16895
rect 6528 16594 6538 16895
rect 6552 16618 6562 16920
rect 6576 16642 6586 16919
rect 6600 16690 6610 16944
rect 7536 16717 7546 17999
rect 37056 17989 37066 18000
rect 37080 17989 37090 18024
rect 11677 17976 12311 17986
rect 14544 17976 35543 17986
rect 12360 17962 12370 17975
rect 10968 17952 12370 17962
rect 10968 17098 10978 17952
rect 11688 17928 12335 17938
rect 10383 17088 10978 17098
rect 10992 17074 11002 17927
rect 9888 17064 11002 17074
rect 9888 17050 9898 17064
rect 9864 17040 9898 17050
rect 9864 17026 9874 17040
rect 11016 17050 11026 17927
rect 9925 17040 11026 17050
rect 9840 17016 9874 17026
rect 9840 17002 9850 17016
rect 11040 17026 11050 17927
rect 9901 17016 11050 17026
rect 9816 16992 9850 17002
rect 9816 16978 9826 16992
rect 11064 17002 11074 17927
rect 9877 16992 11074 17002
rect 9792 16968 9826 16978
rect 9792 16954 9802 16968
rect 11088 16978 11098 17927
rect 9853 16968 11098 16978
rect 9768 16944 9802 16954
rect 9768 16930 9778 16944
rect 11112 16954 11122 17927
rect 9829 16944 11122 16954
rect 9696 16920 9778 16930
rect 9696 16906 9706 16920
rect 11136 16930 11146 17927
rect 9805 16920 11146 16930
rect 11160 16930 11170 17927
rect 11184 16957 11194 17927
rect 11208 16957 11218 17927
rect 11232 16957 11242 17927
rect 11256 16957 11266 17927
rect 11280 16957 11290 17927
rect 11304 16957 11314 17927
rect 11328 16957 11338 17927
rect 11352 16957 11362 17927
rect 11376 16957 11386 17927
rect 11400 16957 11410 17927
rect 11424 16957 11434 17927
rect 11448 16957 11458 17927
rect 11472 16957 11482 17927
rect 11496 16957 11506 17927
rect 11520 16957 11530 17927
rect 11544 16957 11554 17927
rect 11568 16957 11578 17927
rect 11592 16957 11602 17927
rect 11616 16957 11626 17927
rect 11640 16957 11650 17927
rect 11664 16957 11674 17927
rect 11688 16957 11698 17928
rect 11712 17904 12167 17914
rect 11712 16957 11722 17904
rect 13032 16957 13042 17975
rect 13632 16957 13642 17975
rect 13824 16957 13834 17975
rect 14544 16957 14554 17976
rect 14592 17952 27839 17962
rect 14592 16957 14602 17952
rect 36624 17962 36634 17975
rect 36624 17952 37114 17962
rect 16896 17928 27599 17938
rect 14616 16957 14626 17927
rect 15168 16957 15178 17927
rect 15384 16957 15394 17927
rect 16128 16957 16138 17927
rect 16296 16954 16306 17927
rect 16680 16978 16690 17927
rect 16872 17026 16882 17927
rect 16896 17053 16906 17928
rect 20592 17904 27407 17914
rect 17088 17026 17098 17903
rect 17832 17050 17842 17903
rect 18000 17074 18010 17903
rect 20592 17077 20602 17904
rect 18000 17064 19103 17074
rect 17832 17040 22138 17050
rect 16872 17016 16930 17026
rect 17088 17016 22103 17026
rect 16885 16992 16895 17002
rect 16920 17002 16930 17016
rect 22128 17026 22138 17040
rect 22128 17016 22151 17026
rect 16920 16992 24431 17002
rect 16680 16968 25151 16978
rect 36768 16957 36778 17927
rect 36792 16957 36802 17927
rect 36816 16957 36826 17927
rect 36840 16957 36850 17927
rect 36864 16957 36874 17927
rect 36888 16957 36898 17927
rect 16296 16944 28130 16954
rect 36912 16954 36922 17927
rect 36936 16978 36946 17927
rect 36960 17002 36970 17927
rect 36984 17026 36994 17927
rect 37008 17050 37018 17927
rect 37032 17074 37042 17927
rect 37056 17098 37066 17927
rect 37080 17122 37090 17927
rect 37104 17146 37114 17952
rect 37104 17136 37295 17146
rect 37080 17112 37655 17122
rect 37056 17088 37679 17098
rect 37032 17064 37703 17074
rect 37008 17040 37727 17050
rect 36984 17016 37751 17026
rect 36960 16992 37775 17002
rect 36936 16968 37799 16978
rect 41472 16978 41482 26279
rect 41472 16968 41538 16978
rect 41472 16957 41482 16968
rect 36912 16944 37823 16954
rect 11160 16920 41538 16930
rect 9672 16896 9706 16906
rect 9672 16882 9682 16896
rect 9733 16896 11183 16906
rect 16141 16896 28154 16906
rect 36901 16896 37871 16906
rect 9648 16872 9682 16882
rect 9648 16858 9658 16872
rect 11208 16882 11218 16895
rect 9709 16872 11218 16882
rect 11232 16882 11242 16895
rect 11232 16872 11746 16882
rect 11736 16861 11746 16872
rect 9624 16848 9658 16858
rect 9624 16834 9634 16848
rect 9685 16848 11255 16858
rect 9600 16824 9634 16834
rect 9600 16810 9610 16824
rect 11280 16834 11290 16847
rect 9661 16824 11290 16834
rect 11304 16834 11314 16847
rect 11304 16824 11770 16834
rect 11760 16813 11770 16824
rect 13032 16813 13042 16895
rect 13632 16813 13642 16895
rect 9576 16800 9610 16810
rect 9576 16789 9586 16800
rect 9637 16800 11327 16810
rect 13824 16810 13834 16895
rect 14544 16837 14554 16895
rect 14592 16837 14602 16895
rect 14616 16834 14626 16895
rect 15168 16858 15178 16895
rect 15384 16882 15394 16895
rect 15384 16872 30551 16882
rect 15168 16848 32218 16858
rect 14616 16824 19079 16834
rect 19117 16824 30527 16834
rect 30565 16824 32183 16834
rect 32208 16834 32218 16848
rect 32208 16824 32663 16834
rect 13824 16800 34151 16810
rect 36768 16810 36778 16895
rect 36792 16837 36802 16895
rect 36816 16834 36826 16895
rect 36840 16858 36850 16895
rect 36864 16882 36874 16895
rect 36864 16872 37895 16882
rect 36840 16848 37991 16858
rect 36816 16824 38015 16834
rect 41472 16813 41482 16895
rect 36768 16800 38039 16810
rect 11352 16786 11362 16799
rect 9613 16776 11362 16786
rect 11376 16786 11386 16799
rect 11376 16776 36778 16786
rect 9565 16752 11399 16762
rect 11437 16752 11807 16762
rect 13645 16752 35663 16762
rect 36768 16762 36778 16776
rect 36805 16776 41538 16786
rect 36768 16752 38098 16762
rect 38088 16741 38098 16752
rect 9541 16728 11447 16738
rect 11485 16728 38063 16738
rect 9493 16704 11495 16714
rect 11533 16704 11783 16714
rect 11821 16704 37967 16714
rect 38005 16704 38146 16714
rect 38136 16693 38146 16704
rect 6600 16680 10175 16690
rect 10189 16680 11711 16690
rect 11749 16680 38122 16690
rect 9445 16656 11567 16666
rect 11629 16656 11722 16666
rect 6576 16632 9743 16642
rect 9781 16632 11543 16642
rect 11581 16632 11687 16642
rect 6552 16608 11615 16618
rect 11629 16608 11663 16618
rect 11712 16618 11722 16656
rect 11797 16656 37991 16666
rect 38112 16666 38122 16680
rect 38112 16656 38170 16666
rect 11760 16642 11770 16655
rect 11760 16632 38122 16642
rect 11712 16608 37954 16618
rect 6528 16584 10210 16594
rect 7464 16560 10175 16570
rect 7464 12613 7474 16560
rect 10200 16570 10210 16584
rect 10360 16584 11567 16594
rect 11605 16584 37930 16594
rect 10200 16560 10306 16570
rect 10176 16549 10186 16559
rect 10296 16549 10306 16560
rect 10324 16560 11615 16570
rect 10324 16549 10334 16560
rect 11653 16560 37858 16570
rect 7536 16323 7546 16535
rect 9432 16357 9442 16535
rect 9480 16357 9490 16535
rect 9528 16357 9538 16535
rect 9552 16357 9562 16535
rect 9576 16347 9586 16535
rect 9600 16381 9610 16535
rect 9624 16381 9634 16535
rect 9648 16371 9658 16535
rect 9672 16398 9682 16535
rect 9696 16398 9706 16535
rect 9720 16398 9730 16535
rect 9744 16398 9754 16535
rect 9768 16398 9778 16535
rect 9792 16398 9802 16535
rect 9816 16398 9826 16535
rect 9840 16398 9850 16535
rect 9864 16398 9874 16535
rect 9888 16398 9898 16535
rect 9912 16398 9922 16535
rect 37656 16399 37666 16535
rect 37680 16399 37690 16535
rect 37704 16399 37714 16535
rect 37728 16399 37738 16535
rect 37752 16399 37762 16535
rect 37776 16399 37786 16535
rect 37800 16399 37810 16535
rect 37824 16399 37834 16535
rect 37848 16399 37858 16560
rect 37872 16399 37882 16559
rect 37896 16399 37906 16559
rect 37920 16399 37930 16584
rect 37944 16399 37954 16608
rect 37968 16399 37978 16607
rect 37992 16399 38002 16607
rect 38016 16399 38026 16607
rect 9648 16361 9935 16371
rect 38040 16372 38050 16607
rect 37645 16362 38050 16372
rect 9576 16337 9935 16347
rect 37645 16338 38015 16348
rect 7536 16313 9935 16323
rect 37645 16314 37823 16324
rect 9432 12613 9442 16282
rect 37645 16290 37775 16300
rect 9480 12613 9490 16281
rect 9528 12613 9538 16281
rect 9552 12613 9562 16281
rect 9600 12613 9610 16281
rect 9624 12613 9634 16281
rect 9672 12730 9682 16288
rect 9696 12733 9706 16288
rect 9720 12733 9730 16288
rect 9744 12733 9754 16288
rect 9768 12733 9778 16288
rect 9792 12733 9802 16288
rect 9816 12733 9826 16288
rect 9648 12720 9682 12730
rect 9648 12613 9658 12720
rect 9840 12706 9850 16288
rect 9864 12709 9874 16288
rect 9672 12696 9850 12706
rect 9672 12613 9682 12696
rect 9888 12682 9898 16288
rect 9840 12672 9898 12682
rect 9696 12613 9706 12671
rect 9720 12613 9730 12671
rect 9744 12634 9754 12671
rect 9840 12661 9850 12672
rect 9912 12658 9922 16288
rect 37896 16276 37906 16313
rect 37645 16266 37906 16276
rect 37920 16255 37930 16313
rect 37944 16255 37954 16313
rect 37968 16255 37978 16313
rect 37992 16255 38002 16313
rect 38064 16255 38074 16607
rect 38088 16255 38098 16607
rect 38112 16570 38122 16632
rect 38136 16597 38146 16631
rect 38160 16594 38170 16656
rect 38160 16584 41375 16594
rect 41472 16594 41482 16751
rect 41437 16584 41482 16594
rect 38112 16560 41482 16570
rect 37645 16242 37871 16252
rect 38136 16228 38146 16535
rect 37645 16218 38146 16228
rect 9901 12648 9922 12658
rect 9744 12624 9922 12634
rect 9757 12600 9887 12610
rect 9912 12610 9922 12624
rect 9912 12600 9935 12610
rect 6504 12576 9935 12586
rect 9901 12552 9935 12562
rect 6450 12192 6514 12202
rect 6504 8098 6514 12192
rect 7464 8125 7474 12551
rect 9432 8125 9442 12551
rect 9480 12538 9490 12551
rect 9480 12528 9935 12538
rect 9528 8125 9538 12503
rect 9552 8125 9562 12503
rect 9600 8125 9610 12503
rect 9624 8417 9634 12503
rect 9648 8465 9658 12503
rect 9672 8492 9682 12503
rect 9696 8492 9706 12503
rect 9720 8492 9730 12503
rect 9744 8492 9754 12503
rect 9768 8492 9778 12503
rect 9792 8492 9802 12503
rect 9816 8492 9826 12503
rect 9840 8492 9850 12503
rect 9864 8492 9874 12503
rect 9888 8492 9898 12503
rect 9912 8492 9922 12528
rect 37656 10333 37666 16193
rect 37680 10333 37690 16193
rect 37704 10333 37714 16193
rect 37728 10306 37738 16193
rect 37645 10296 37738 10306
rect 37656 10213 37666 10271
rect 37680 10213 37690 10271
rect 37704 10213 37714 10271
rect 37752 10213 37762 16193
rect 37800 10213 37810 16193
rect 37848 10213 37858 16193
rect 37920 10213 37930 16193
rect 37944 10213 37954 16193
rect 37968 10213 37978 16193
rect 37992 10186 38002 16193
rect 37645 10176 38002 10186
rect 37645 10152 37967 10162
rect 37656 8515 37666 10127
rect 37680 8515 37690 10127
rect 37704 8515 37714 10127
rect 37752 8515 37762 10127
rect 37800 8515 37810 10127
rect 37848 8488 37858 10127
rect 37645 8478 37858 8488
rect 9648 8455 9935 8465
rect 9685 8431 9935 8441
rect 37680 8441 37690 8454
rect 37645 8431 37690 8441
rect 9624 8407 9935 8417
rect 37920 8417 37930 10127
rect 37645 8407 37930 8417
rect 9733 8383 9935 8393
rect 37944 8393 37954 10127
rect 38064 8396 38074 16193
rect 37645 8383 37954 8393
rect 9696 8125 9706 8382
rect 38088 8369 38098 16193
rect 41376 12058 41386 16535
rect 41424 12250 41434 16535
rect 41472 12274 41482 16560
rect 41461 12264 41482 12274
rect 41424 12240 41538 12250
rect 41472 12229 41482 12240
rect 41448 12202 41458 12215
rect 41448 12192 41538 12202
rect 41472 12085 41482 12167
rect 41376 12048 41538 12058
rect 37645 8359 38098 8369
rect 9744 8290 9754 8358
rect 9768 8317 9778 8358
rect 9792 8317 9802 8358
rect 9816 8317 9826 8358
rect 9840 8317 9850 8358
rect 9864 8317 9874 8358
rect 9888 8317 9898 8358
rect 9912 8317 9922 8358
rect 37645 8335 37703 8345
rect 9744 8280 9935 8290
rect 10296 8290 10306 8303
rect 10008 8280 10306 8290
rect 9853 8256 9959 8266
rect 9768 8146 9778 8255
rect 9792 8218 9802 8255
rect 9877 8232 9983 8242
rect 10008 8218 10018 8280
rect 10372 8266 10382 8303
rect 37752 8290 37762 8334
rect 9792 8208 10018 8218
rect 10032 8256 10382 8266
rect 36456 8280 37762 8290
rect 9829 8184 10007 8194
rect 10032 8170 10042 8256
rect 9877 8160 10042 8170
rect 10056 8232 10346 8242
rect 9768 8136 10042 8146
rect 10032 8125 10042 8136
rect 10056 8098 10066 8232
rect 6504 8088 10066 8098
rect 7464 7501 7474 8063
rect 9432 7501 9442 8063
rect 9528 7501 9538 8063
rect 9552 7501 9562 8063
rect 9600 7501 9610 8063
rect 9696 7501 9706 8063
rect 9864 7474 9874 8063
rect 6450 7464 9874 7474
rect 7464 6565 7474 7439
rect 9432 6586 9442 7439
rect 9528 6613 9538 7439
rect 9552 6658 9562 7439
rect 9600 6685 9610 7439
rect 9696 6685 9706 7439
rect 9888 6685 9898 8063
rect 9912 6685 9922 8063
rect 9936 6685 9946 8063
rect 9960 6682 9970 8063
rect 9984 6706 9994 8063
rect 10008 6730 10018 8063
rect 10032 6754 10042 8063
rect 10032 6744 11567 6754
rect 10008 6720 11711 6730
rect 9984 6696 15695 6706
rect 9960 6672 15850 6682
rect 9552 6648 11687 6658
rect 11725 6648 15815 6658
rect 15840 6658 15850 6672
rect 15840 6648 19799 6658
rect 9949 6624 19967 6634
rect 9600 6610 9610 6623
rect 9600 6600 28090 6610
rect 9432 6576 28055 6586
rect 28080 6586 28090 6600
rect 28080 6576 28234 6586
rect 9541 6552 28199 6562
rect 28224 6562 28234 6576
rect 36456 6565 36466 8280
rect 37656 7474 37666 8255
rect 37800 7501 37810 8334
rect 38064 7501 38074 8334
rect 41472 7522 41482 12023
rect 41472 7512 41538 7522
rect 37656 7464 41538 7474
rect 37800 7330 37810 7439
rect 38064 7357 38074 7439
rect 37800 7320 41538 7330
rect 28224 6552 32207 6562
rect 7440 6528 9887 6538
rect 7440 6514 7450 6528
rect 9925 6528 11735 6538
rect 11749 6528 15863 6538
rect 15877 6528 19991 6538
rect 20005 6528 28247 6538
rect 28261 6528 32362 6538
rect 7416 6504 7450 6514
rect 7416 6450 7426 6504
rect 7477 6504 7522 6514
rect 7464 6450 7474 6503
rect 7512 6450 7522 6504
rect 9709 6504 11554 6514
rect 11544 6450 11554 6504
rect 11581 6504 15682 6514
rect 11688 6450 11698 6479
rect 11736 6450 11746 6479
rect 15672 6450 15682 6504
rect 15709 6504 19954 6514
rect 15816 6450 15826 6479
rect 15864 6450 15874 6479
rect 19800 6450 19810 6479
rect 19944 6450 19954 6504
rect 19981 6504 32194 6514
rect 19992 6450 20002 6479
rect 28056 6450 28066 6479
rect 28200 6450 28210 6479
rect 28248 6450 28258 6479
rect 32184 6450 32194 6504
rect 32352 6514 32362 6528
rect 36325 6528 36538 6538
rect 36528 6514 36538 6528
rect 38064 6514 38074 7295
rect 32221 6504 32338 6514
rect 32352 6504 36514 6514
rect 36528 6504 38074 6514
rect 32328 6450 32338 6504
rect 32376 6450 32386 6504
rect 36312 6450 36322 6479
rect 36456 6450 36466 6479
rect 36504 6450 36514 6504
<< m2contact >>
rect 15599 41423 15613 41437
rect 15647 41423 15661 41437
rect 19727 41423 19741 41437
rect 19775 41423 19789 41437
rect 19919 41423 19933 41437
rect 27983 41423 27997 41437
rect 28031 41423 28045 41437
rect 11615 41399 11629 41413
rect 32111 41423 32125 41437
rect 32159 41423 32173 41437
rect 28199 41399 28213 41413
rect 36239 41423 36253 41437
rect 36431 41423 36445 41437
rect 32327 41399 32341 41413
rect 36263 41399 36277 41413
rect 36287 41399 36301 41413
rect 28031 41375 28045 41389
rect 28055 41375 28069 41389
rect 32111 41375 32125 41389
rect 36239 41375 36253 41389
rect 15647 41351 15661 41365
rect 15671 41351 15685 41365
rect 36287 41351 36301 41365
rect 36431 41375 36445 41389
rect 11639 41327 11653 41341
rect 11663 41327 11677 41341
rect 32159 41327 32173 41341
rect 32327 41327 32341 41341
rect 36263 41327 36277 41341
rect 11519 41279 11533 41293
rect 11567 41279 11581 41293
rect 11591 41279 11605 41293
rect 11687 41279 11701 41293
rect 19775 41279 19789 41293
rect 19799 41279 19813 41293
rect 28199 41279 28213 41293
rect 11519 41231 11533 41245
rect 6503 40391 6517 40405
rect 7439 40391 7453 40405
rect 7535 40391 7549 40405
rect 11519 40391 11533 40405
rect 15599 41255 15613 41269
rect 15623 41255 15637 41269
rect 19727 41255 19741 41269
rect 27983 41255 27997 41269
rect 28055 41255 28069 41269
rect 11567 41231 11581 41245
rect 11591 41231 11605 41245
rect 11615 41231 11629 41245
rect 11639 41231 11653 41245
rect 11663 41231 11677 41245
rect 11687 41231 11701 41245
rect 6503 40343 6517 40357
rect 7439 40343 7453 40357
rect 7535 40343 7549 40357
rect 11519 40343 11533 40357
rect 11519 39287 11533 39301
rect 11471 39263 11485 39277
rect 19919 41231 19933 41245
rect 19799 41207 19813 41221
rect 15671 41183 15685 41197
rect 15623 41159 15637 41173
rect 15599 41135 15613 41149
rect 11591 39263 11605 39277
rect 11615 39263 11629 39277
rect 11639 39263 11653 39277
rect 11663 39263 11677 39277
rect 11687 39263 11701 39277
rect 11711 39263 11725 39277
rect 11735 39263 11749 39277
rect 11759 39263 11773 39277
rect 11783 39263 11797 39277
rect 11423 39239 11437 39253
rect 11375 39215 11389 39229
rect 11591 39215 11605 39229
rect 11351 39191 11365 39205
rect 11831 39191 11845 39205
rect 11303 39143 11317 39157
rect 11327 39143 11341 39157
rect 11471 39119 11485 39133
rect 11495 39119 11509 39133
rect 11783 39119 11797 39133
rect 11831 39143 11845 39157
rect 7535 39095 7549 39109
rect 11279 39095 11293 39109
rect 11399 39095 11413 39109
rect 11783 39095 11797 39109
rect 11807 39095 11821 39109
rect 27239 39239 27253 39253
rect 26519 39215 26533 39229
rect 29087 39215 29101 39229
rect 26255 39191 26269 39205
rect 29255 39191 29269 39205
rect 29399 39191 29413 39205
rect 15599 39167 15613 39181
rect 18263 39167 18277 39181
rect 29471 39167 29485 39181
rect 36623 39167 36637 39181
rect 41471 40607 41485 40621
rect 41471 40559 41485 40573
rect 41447 40463 41461 40477
rect 41471 40463 41485 40477
rect 11855 39119 11869 39133
rect 17231 39119 17245 39133
rect 29351 39119 29365 39133
rect 29375 39119 29389 39133
rect 29423 39119 29437 39133
rect 29447 39119 29461 39133
rect 36647 39119 36661 39133
rect 36791 39143 36805 39157
rect 11879 39095 11893 39109
rect 17039 39095 17053 39109
rect 29063 39095 29077 39109
rect 29087 39095 29101 39109
rect 36839 39095 36853 39109
rect 36863 39095 36877 39109
rect 11831 39071 11845 39085
rect 11855 39071 11869 39085
rect 36887 39071 36901 39085
rect 7535 39047 7549 39061
rect 11303 39047 11317 39061
rect 11327 39047 11341 39061
rect 11351 39047 11365 39061
rect 11375 39047 11389 39061
rect 11399 39047 11413 39061
rect 11423 39047 11437 39061
rect 6527 35735 6541 35749
rect 6527 35687 6541 35701
rect 6503 35663 6517 35677
rect 6503 35615 6517 35629
rect 6503 30983 6517 30997
rect 6551 31007 6565 31021
rect 6527 30935 6541 30949
rect 6503 30887 6517 30901
rect 6527 30887 6541 30901
rect 6551 30887 6565 30901
rect 6503 26303 6517 26317
rect 6527 26303 6541 26317
rect 6503 26255 6517 26269
rect 6527 26255 6541 26269
rect 6503 21671 6517 21685
rect 6527 21671 6541 21685
rect 6551 21671 6565 21685
rect 6575 21671 6589 21685
rect 6503 21623 6517 21637
rect 6527 21623 6541 21637
rect 6551 21623 6565 21637
rect 6575 21623 6589 21637
rect 6503 16943 6517 16957
rect 6527 16943 6541 16957
rect 11255 38999 11269 39013
rect 11855 39047 11869 39061
rect 11879 39047 11893 39061
rect 11879 39023 11893 39037
rect 16079 39047 16093 39061
rect 29375 39047 29389 39061
rect 29399 39047 29413 39061
rect 36767 39047 36781 39061
rect 36791 39047 36805 39061
rect 36911 39023 36925 39037
rect 36959 39023 36973 39037
rect 11327 38999 11341 39013
rect 11351 38999 11365 39013
rect 11375 38999 11389 39013
rect 11399 38999 11413 39013
rect 11423 38999 11437 39013
rect 11447 38999 11461 39013
rect 11471 38999 11485 39013
rect 11543 38999 11557 39013
rect 41447 40415 41461 40429
rect 41471 40415 41485 40429
rect 11279 38975 11293 38989
rect 11303 38975 11317 38989
rect 12191 38975 12205 38989
rect 15599 38975 15613 38989
rect 15839 38975 15853 38989
rect 29447 38975 29461 38989
rect 29471 38975 29485 38989
rect 36815 38975 36829 38989
rect 36863 38975 36877 38989
rect 36983 38975 36997 38989
rect 11231 38927 11245 38941
rect 11207 38903 11221 38917
rect 11759 38951 11773 38965
rect 11783 38951 11797 38965
rect 11807 38951 11821 38965
rect 11831 38951 11845 38965
rect 11855 38951 11869 38965
rect 11879 38951 11893 38965
rect 12311 38951 12325 38965
rect 11735 38927 11749 38941
rect 11567 38903 11581 38917
rect 11591 38903 11605 38917
rect 11711 38903 11725 38917
rect 11183 38879 11197 38893
rect 11687 38879 11701 38893
rect 11783 38879 11797 38893
rect 29303 38927 29317 38941
rect 29351 38951 29365 38965
rect 36863 38951 36877 38965
rect 36887 38951 36901 38965
rect 37007 38951 37021 38965
rect 36623 38927 36637 38941
rect 36647 38927 36661 38941
rect 36887 38927 36901 38941
rect 36911 38927 36925 38941
rect 12167 38903 12181 38917
rect 12191 38903 12205 38917
rect 29399 38903 29413 38917
rect 29423 38903 29437 38917
rect 37007 38903 37021 38917
rect 37031 38903 37045 38917
rect 29039 38879 29053 38893
rect 29063 38879 29077 38893
rect 36911 38879 36925 38893
rect 36935 38879 36949 38893
rect 11159 38855 11173 38869
rect 11231 38855 11245 38869
rect 11279 38855 11293 38869
rect 37007 38855 37021 38869
rect 37055 38855 37069 38869
rect 11183 38831 11197 38845
rect 11231 38831 11245 38845
rect 11159 38807 11173 38821
rect 11663 38807 11677 38821
rect 11783 38807 11797 38821
rect 12311 38807 12325 38821
rect 29255 38807 29269 38821
rect 11207 38783 11221 38797
rect 11231 38783 11245 38797
rect 11255 38783 11269 38797
rect 11279 38783 11293 38797
rect 11303 38783 11317 38797
rect 11327 38783 11341 38797
rect 11351 38783 11365 38797
rect 11375 38783 11389 38797
rect 11399 38783 11413 38797
rect 11423 38783 11437 38797
rect 11447 38783 11461 38797
rect 11471 38783 11485 38797
rect 11495 38783 11509 38797
rect 11519 38783 11533 38797
rect 11543 38783 11557 38797
rect 11567 38783 11581 38797
rect 11591 38783 11605 38797
rect 11615 38783 11629 38797
rect 11639 38783 11653 38797
rect 12287 38783 12301 38797
rect 29231 38783 29245 38797
rect 36767 38783 36781 38797
rect 11135 36095 11149 36109
rect 11159 36095 11173 36109
rect 11183 36095 11197 36109
rect 11207 36095 11221 36109
rect 11231 36095 11245 36109
rect 11255 36095 11269 36109
rect 11279 36095 11293 36109
rect 11303 36095 11317 36109
rect 11327 36095 11341 36109
rect 11351 36095 11365 36109
rect 11375 36095 11389 36109
rect 11399 36095 11413 36109
rect 11423 36095 11437 36109
rect 11447 36095 11461 36109
rect 11471 36095 11485 36109
rect 11495 36095 11509 36109
rect 11519 36095 11533 36109
rect 11543 36095 11557 36109
rect 11567 36095 11581 36109
rect 11615 36071 11629 36085
rect 11639 36071 11653 36085
rect 11591 36047 11605 36061
rect 11135 35999 11149 36013
rect 11159 35951 11173 35965
rect 11183 35951 11197 35965
rect 11207 35951 11221 35965
rect 11231 35951 11245 35965
rect 11255 35951 11269 35965
rect 11279 35951 11293 35965
rect 11303 35951 11317 35965
rect 11327 35951 11341 35965
rect 11351 35951 11365 35965
rect 11375 35951 11389 35965
rect 11399 35951 11413 35965
rect 11423 35951 11437 35965
rect 11447 35951 11461 35965
rect 11471 35951 11485 35965
rect 11495 35951 11509 35965
rect 11519 35951 11533 35965
rect 11543 35951 11557 35965
rect 11567 35951 11581 35965
rect 11591 35951 11605 35965
rect 11615 35951 11629 35965
rect 11639 35951 11653 35965
rect 11159 34919 11173 34933
rect 11183 34919 11197 34933
rect 11207 34919 11221 34933
rect 11231 34919 11245 34933
rect 11255 34919 11269 34933
rect 11279 34919 11293 34933
rect 11303 34919 11317 34933
rect 11327 34919 11341 34933
rect 11351 34919 11365 34933
rect 11375 34919 11389 34933
rect 11399 34919 11413 34933
rect 11423 34919 11437 34933
rect 11447 34919 11461 34933
rect 11471 34919 11485 34933
rect 11495 34919 11509 34933
rect 11519 34919 11533 34933
rect 11543 34919 11557 34933
rect 11567 34919 11581 34933
rect 11591 34919 11605 34933
rect 11639 34895 11653 34909
rect 11615 34871 11629 34885
rect 11159 34823 11173 34837
rect 11183 34775 11197 34789
rect 11207 34775 11221 34789
rect 11231 34775 11245 34789
rect 11255 34775 11269 34789
rect 11279 34775 11293 34789
rect 11303 34775 11317 34789
rect 11327 34775 11341 34789
rect 11351 34775 11365 34789
rect 11375 34775 11389 34789
rect 11399 34775 11413 34789
rect 11423 34775 11437 34789
rect 11447 34775 11461 34789
rect 11471 34775 11485 34789
rect 11495 34775 11509 34789
rect 11519 34775 11533 34789
rect 11543 34775 11557 34789
rect 11567 34775 11581 34789
rect 11591 34775 11605 34789
rect 11615 34775 11629 34789
rect 11639 34775 11653 34789
rect 11183 33743 11197 33757
rect 11207 33743 11221 33757
rect 11231 33743 11245 33757
rect 11255 33743 11269 33757
rect 11279 33743 11293 33757
rect 11303 33743 11317 33757
rect 11327 33743 11341 33757
rect 11351 33743 11365 33757
rect 11375 33743 11389 33757
rect 11399 33743 11413 33757
rect 11423 33743 11437 33757
rect 11447 33743 11461 33757
rect 11471 33743 11485 33757
rect 11495 33743 11509 33757
rect 11519 33743 11533 33757
rect 11543 33743 11557 33757
rect 11591 33719 11605 33733
rect 11615 33719 11629 33733
rect 11639 33719 11653 33733
rect 11567 33695 11581 33709
rect 11183 33647 11197 33661
rect 11207 33599 11221 33613
rect 11231 33599 11245 33613
rect 11255 33599 11269 33613
rect 11279 33599 11293 33613
rect 11303 33599 11317 33613
rect 11327 33599 11341 33613
rect 11351 33599 11365 33613
rect 11375 33599 11389 33613
rect 11399 33599 11413 33613
rect 11423 33599 11437 33613
rect 11447 33599 11461 33613
rect 11471 33599 11485 33613
rect 11495 33599 11509 33613
rect 11519 33599 11533 33613
rect 11543 33599 11557 33613
rect 11567 33599 11581 33613
rect 11591 33599 11605 33613
rect 11615 33599 11629 33613
rect 11639 33599 11653 33613
rect 11207 32567 11221 32581
rect 11231 32567 11245 32581
rect 11255 32567 11269 32581
rect 11279 32567 11293 32581
rect 11303 32567 11317 32581
rect 11327 32567 11341 32581
rect 11351 32567 11365 32581
rect 11399 32543 11413 32557
rect 11423 32543 11437 32557
rect 11447 32543 11461 32557
rect 11471 32543 11485 32557
rect 11495 32543 11509 32557
rect 11519 32543 11533 32557
rect 11543 32543 11557 32557
rect 11567 32543 11581 32557
rect 11591 32543 11605 32557
rect 11615 32543 11629 32557
rect 11639 32543 11653 32557
rect 11375 32519 11389 32533
rect 11207 32471 11221 32485
rect 11231 32423 11245 32437
rect 11255 32423 11269 32437
rect 11279 32423 11293 32437
rect 11303 32423 11317 32437
rect 11327 32423 11341 32437
rect 11351 32423 11365 32437
rect 11375 32423 11389 32437
rect 11399 32423 11413 32437
rect 11423 32423 11437 32437
rect 11447 32423 11461 32437
rect 11471 32423 11485 32437
rect 11495 32423 11509 32437
rect 11519 32423 11533 32437
rect 11543 32423 11557 32437
rect 11567 32423 11581 32437
rect 11591 32423 11605 32437
rect 11615 32423 11629 32437
rect 11639 32423 11653 32437
rect 11231 31391 11245 31405
rect 11255 31391 11269 31405
rect 11279 31391 11293 31405
rect 11303 31391 11317 31405
rect 11327 31391 11341 31405
rect 11351 31391 11365 31405
rect 11375 31391 11389 31405
rect 11399 31391 11413 31405
rect 11423 31391 11437 31405
rect 11447 31391 11461 31405
rect 11471 31391 11485 31405
rect 11495 31391 11509 31405
rect 11519 31391 11533 31405
rect 11567 31367 11581 31381
rect 11591 31367 11605 31381
rect 11615 31367 11629 31381
rect 11639 31367 11653 31381
rect 11543 31343 11557 31357
rect 11231 31295 11245 31309
rect 11255 31247 11269 31261
rect 11279 31247 11293 31261
rect 11303 31247 11317 31261
rect 11327 31247 11341 31261
rect 11351 31247 11365 31261
rect 11375 31247 11389 31261
rect 11399 31247 11413 31261
rect 11423 31247 11437 31261
rect 11447 31247 11461 31261
rect 11471 31247 11485 31261
rect 11495 31247 11509 31261
rect 11519 31247 11533 31261
rect 11543 31247 11557 31261
rect 11567 31247 11581 31261
rect 11591 31247 11605 31261
rect 11615 31247 11629 31261
rect 11639 31247 11653 31261
rect 11255 30215 11269 30229
rect 11279 30215 11293 30229
rect 11303 30215 11317 30229
rect 11327 30215 11341 30229
rect 11375 30191 11389 30205
rect 11399 30191 11413 30205
rect 11423 30191 11437 30205
rect 11447 30191 11461 30205
rect 11471 30191 11485 30205
rect 11495 30191 11509 30205
rect 11519 30191 11533 30205
rect 11543 30191 11557 30205
rect 11567 30191 11581 30205
rect 11591 30191 11605 30205
rect 11615 30191 11629 30205
rect 11639 30191 11653 30205
rect 11351 30167 11365 30181
rect 11255 30119 11269 30133
rect 11279 30071 11293 30085
rect 11303 30071 11317 30085
rect 11327 30071 11341 30085
rect 11351 30071 11365 30085
rect 11375 30071 11389 30085
rect 11399 30071 11413 30085
rect 11423 30071 11437 30085
rect 11447 30071 11461 30085
rect 11471 30071 11485 30085
rect 11495 30071 11509 30085
rect 11519 30071 11533 30085
rect 11543 30071 11557 30085
rect 11567 30071 11581 30085
rect 11591 30071 11605 30085
rect 11615 30071 11629 30085
rect 11639 30071 11653 30085
rect 11279 29039 11293 29053
rect 11303 29039 11317 29053
rect 11327 29039 11341 29053
rect 11351 29039 11365 29053
rect 11375 29039 11389 29053
rect 11399 29039 11413 29053
rect 11447 29015 11461 29029
rect 11471 29015 11485 29029
rect 11495 29015 11509 29029
rect 11519 29015 11533 29029
rect 11543 29015 11557 29029
rect 11567 29015 11581 29029
rect 11591 29015 11605 29029
rect 11615 29015 11629 29029
rect 11639 29015 11653 29029
rect 11423 28991 11437 29005
rect 11279 28943 11293 28957
rect 11303 28895 11317 28909
rect 11327 28895 11341 28909
rect 11351 28895 11365 28909
rect 11375 28895 11389 28909
rect 11399 28895 11413 28909
rect 11423 28895 11437 28909
rect 11447 28895 11461 28909
rect 11471 28895 11485 28909
rect 11495 28895 11509 28909
rect 11519 28895 11533 28909
rect 11543 28895 11557 28909
rect 11567 28895 11581 28909
rect 11591 28895 11605 28909
rect 11615 28895 11629 28909
rect 11639 28895 11653 28909
rect 11303 27863 11317 27877
rect 11327 27863 11341 27877
rect 11351 27863 11365 27877
rect 11375 27863 11389 27877
rect 11399 27863 11413 27877
rect 11423 27863 11437 27877
rect 11447 27863 11461 27877
rect 11471 27863 11485 27877
rect 11495 27863 11509 27877
rect 11519 27863 11533 27877
rect 11543 27863 11557 27877
rect 11567 27863 11581 27877
rect 11591 27863 11605 27877
rect 11615 27863 11629 27877
rect 11279 27839 11293 27853
rect 11471 27815 11485 27829
rect 11639 27815 11653 27829
rect 11255 27791 11269 27805
rect 11447 27791 11461 27805
rect 11471 27767 11485 27781
rect 11255 27743 11269 27757
rect 11279 27743 11293 27757
rect 11303 27743 11317 27757
rect 11327 27743 11341 27757
rect 11351 27743 11365 27757
rect 11375 27743 11389 27757
rect 11399 27743 11413 27757
rect 11423 27743 11437 27757
rect 11471 27719 11485 27733
rect 11495 27719 11509 27733
rect 11519 27719 11533 27733
rect 11543 27719 11557 27733
rect 11567 27719 11581 27733
rect 11591 27719 11605 27733
rect 11615 27719 11629 27733
rect 11639 27719 11653 27733
rect 11255 26639 11269 26653
rect 11279 26639 11293 26653
rect 11303 26639 11317 26653
rect 11327 26639 11341 26653
rect 11351 26639 11365 26653
rect 11375 26639 11389 26653
rect 11399 26639 11413 26653
rect 11423 26639 11437 26653
rect 11447 26639 11461 26653
rect 11471 26639 11485 26653
rect 11495 26639 11509 26653
rect 11519 26639 11533 26653
rect 11543 26639 11557 26653
rect 11567 26639 11581 26653
rect 11591 26639 11605 26653
rect 11615 26639 11629 26653
rect 11639 26639 11653 26653
rect 11207 26615 11221 26629
rect 11231 26615 11245 26629
rect 11303 26591 11317 26605
rect 11207 26567 11221 26581
rect 11231 26567 11245 26581
rect 11255 26567 11269 26581
rect 11279 26567 11293 26581
rect 11327 26543 11341 26557
rect 11351 26543 11365 26557
rect 11375 26543 11389 26557
rect 11399 26543 11413 26557
rect 11423 26543 11437 26557
rect 11447 26543 11461 26557
rect 11471 26543 11485 26557
rect 11495 26543 11509 26557
rect 11519 26543 11533 26557
rect 11543 26543 11557 26557
rect 11567 26543 11581 26557
rect 11591 26543 11605 26557
rect 11615 26543 11629 26557
rect 11639 26543 11653 26557
rect 11183 25487 11197 25501
rect 11207 25487 11221 25501
rect 11231 25487 11245 25501
rect 11255 25487 11269 25501
rect 11279 25487 11293 25501
rect 11303 25487 11317 25501
rect 11327 25487 11341 25501
rect 11351 25487 11365 25501
rect 11375 25487 11389 25501
rect 11399 25487 11413 25501
rect 11423 25487 11437 25501
rect 11471 25463 11485 25477
rect 11495 25463 11509 25477
rect 11519 25463 11533 25477
rect 11543 25463 11557 25477
rect 11567 25463 11581 25477
rect 11591 25463 11605 25477
rect 11615 25463 11629 25477
rect 11639 25463 11653 25477
rect 11159 25439 11173 25453
rect 11399 25439 11413 25453
rect 11447 25415 11461 25429
rect 11159 25391 11173 25405
rect 11183 25391 11197 25405
rect 11207 25391 11221 25405
rect 11231 25391 11245 25405
rect 11255 25391 11269 25405
rect 11279 25391 11293 25405
rect 11303 25391 11317 25405
rect 11327 25391 11341 25405
rect 11351 25391 11365 25405
rect 11375 25391 11389 25405
rect 11423 25367 11437 25381
rect 11447 25367 11461 25381
rect 11471 25367 11485 25381
rect 11495 25367 11509 25381
rect 11519 25367 11533 25381
rect 11543 25367 11557 25381
rect 11567 25367 11581 25381
rect 11591 25367 11605 25381
rect 11615 25367 11629 25381
rect 11639 25367 11653 25381
rect 11135 24311 11149 24325
rect 11159 24311 11173 24325
rect 11183 24311 11197 24325
rect 11207 24311 11221 24325
rect 11231 24311 11245 24325
rect 11255 24311 11269 24325
rect 11279 24311 11293 24325
rect 11303 24311 11317 24325
rect 11327 24311 11341 24325
rect 11351 24311 11365 24325
rect 11375 24311 11389 24325
rect 11399 24311 11413 24325
rect 11423 24311 11437 24325
rect 11447 24311 11461 24325
rect 11495 24287 11509 24301
rect 11519 24287 11533 24301
rect 11543 24287 11557 24301
rect 11567 24287 11581 24301
rect 11591 24287 11605 24301
rect 11615 24287 11629 24301
rect 11639 24287 11653 24301
rect 11111 24263 11125 24277
rect 11207 24263 11221 24277
rect 11471 24239 11485 24253
rect 11111 24215 11125 24229
rect 11135 24215 11149 24229
rect 11159 24215 11173 24229
rect 11183 24215 11197 24229
rect 11231 24191 11245 24205
rect 11255 24191 11269 24205
rect 11279 24191 11293 24205
rect 11303 24191 11317 24205
rect 11327 24191 11341 24205
rect 11351 24191 11365 24205
rect 11375 24191 11389 24205
rect 11399 24191 11413 24205
rect 11423 24191 11437 24205
rect 11447 24191 11461 24205
rect 11471 24191 11485 24205
rect 11495 24191 11509 24205
rect 11519 24191 11533 24205
rect 11543 24191 11557 24205
rect 11567 24191 11581 24205
rect 11591 24191 11605 24205
rect 11615 24191 11629 24205
rect 11639 24191 11653 24205
rect 11087 23135 11101 23149
rect 11111 23135 11125 23149
rect 11135 23135 11149 23149
rect 11159 23135 11173 23149
rect 11183 23135 11197 23149
rect 11207 23135 11221 23149
rect 11231 23135 11245 23149
rect 11255 23135 11269 23149
rect 11279 23135 11293 23149
rect 11303 23135 11317 23149
rect 11327 23135 11341 23149
rect 11351 23135 11365 23149
rect 11375 23135 11389 23149
rect 11399 23135 11413 23149
rect 11423 23135 11437 23149
rect 11447 23135 11461 23149
rect 11471 23135 11485 23149
rect 11495 23135 11509 23149
rect 11519 23135 11533 23149
rect 11543 23135 11557 23149
rect 11591 23111 11605 23125
rect 11615 23111 11629 23125
rect 11639 23111 11653 23125
rect 11063 23087 11077 23101
rect 11351 23087 11365 23101
rect 11567 23063 11581 23077
rect 11063 23039 11077 23053
rect 11087 23039 11101 23053
rect 11111 23039 11125 23053
rect 11135 23039 11149 23053
rect 11159 23039 11173 23053
rect 11183 23039 11197 23053
rect 11207 23039 11221 23053
rect 11231 23039 11245 23053
rect 11255 23039 11269 23053
rect 11279 23039 11293 23053
rect 11303 23039 11317 23053
rect 11327 23039 11341 23053
rect 11375 23015 11389 23029
rect 11399 23015 11413 23029
rect 11423 23015 11437 23029
rect 11447 23015 11461 23029
rect 11471 23015 11485 23029
rect 11495 23015 11509 23029
rect 11519 23015 11533 23029
rect 11543 23015 11557 23029
rect 11567 23015 11581 23029
rect 11591 23015 11605 23029
rect 11615 23015 11629 23029
rect 11639 23015 11653 23029
rect 11039 21959 11053 21973
rect 11063 21959 11077 21973
rect 11087 21959 11101 21973
rect 11111 21959 11125 21973
rect 11135 21959 11149 21973
rect 11159 21959 11173 21973
rect 11183 21959 11197 21973
rect 11207 21959 11221 21973
rect 11231 21959 11245 21973
rect 11255 21959 11269 21973
rect 11279 21959 11293 21973
rect 11303 21959 11317 21973
rect 11327 21959 11341 21973
rect 11351 21959 11365 21973
rect 11375 21959 11389 21973
rect 11399 21959 11413 21973
rect 11423 21959 11437 21973
rect 11447 21959 11461 21973
rect 11471 21959 11485 21973
rect 11495 21959 11509 21973
rect 11519 21959 11533 21973
rect 11543 21959 11557 21973
rect 11591 21935 11605 21949
rect 11615 21935 11629 21949
rect 11639 21935 11653 21949
rect 11015 21911 11029 21925
rect 11447 21911 11461 21925
rect 11567 21887 11581 21901
rect 11015 21863 11029 21877
rect 11039 21863 11053 21877
rect 11063 21863 11077 21877
rect 11087 21863 11101 21877
rect 11111 21863 11125 21877
rect 11135 21863 11149 21877
rect 11159 21863 11173 21877
rect 11183 21863 11197 21877
rect 11207 21863 11221 21877
rect 11231 21863 11245 21877
rect 11255 21863 11269 21877
rect 11279 21863 11293 21877
rect 11303 21863 11317 21877
rect 11327 21863 11341 21877
rect 11351 21863 11365 21877
rect 11375 21863 11389 21877
rect 11399 21863 11413 21877
rect 11423 21863 11437 21877
rect 10991 20783 11005 20797
rect 11015 20783 11029 20797
rect 11471 21839 11485 21853
rect 11495 21839 11509 21853
rect 11519 21839 11533 21853
rect 11543 21839 11557 21853
rect 11567 21839 11581 21853
rect 11591 21839 11605 21853
rect 11615 21839 11629 21853
rect 11639 21839 11653 21853
rect 11063 20759 11077 20773
rect 11087 20759 11101 20773
rect 11111 20759 11125 20773
rect 11135 20759 11149 20773
rect 11159 20759 11173 20773
rect 11183 20759 11197 20773
rect 11207 20759 11221 20773
rect 11231 20759 11245 20773
rect 11255 20759 11269 20773
rect 11279 20759 11293 20773
rect 11303 20759 11317 20773
rect 11327 20759 11341 20773
rect 11351 20759 11365 20773
rect 11375 20759 11389 20773
rect 11399 20759 11413 20773
rect 11423 20759 11437 20773
rect 11447 20759 11461 20773
rect 11471 20759 11485 20773
rect 11495 20759 11509 20773
rect 11519 20759 11533 20773
rect 11543 20759 11557 20773
rect 11567 20759 11581 20773
rect 11591 20759 11605 20773
rect 11615 20759 11629 20773
rect 11639 20759 11653 20773
rect 10967 20735 10981 20749
rect 11039 20735 11053 20749
rect 11063 20711 11077 20725
rect 10967 20687 10981 20701
rect 10991 20687 11005 20701
rect 11015 20687 11029 20701
rect 11039 20687 11053 20701
rect 10943 19655 10957 19669
rect 10967 19655 10981 19669
rect 11087 20663 11101 20677
rect 11111 20663 11125 20677
rect 11135 20663 11149 20677
rect 11159 20663 11173 20677
rect 11183 20663 11197 20677
rect 11207 20663 11221 20677
rect 11231 20663 11245 20677
rect 11255 20663 11269 20677
rect 11279 20663 11293 20677
rect 11303 20663 11317 20677
rect 11327 20663 11341 20677
rect 11351 20663 11365 20677
rect 11375 20663 11389 20677
rect 11399 20663 11413 20677
rect 11423 20663 11437 20677
rect 11447 20663 11461 20677
rect 11471 20663 11485 20677
rect 11495 20663 11509 20677
rect 11519 20663 11533 20677
rect 11543 20663 11557 20677
rect 11567 20663 11581 20677
rect 11591 20663 11605 20677
rect 11615 20663 11629 20677
rect 11639 20663 11653 20677
rect 11015 19631 11029 19645
rect 11039 19631 11053 19645
rect 11063 19631 11077 19645
rect 11087 19631 11101 19645
rect 11111 19631 11125 19645
rect 11135 19631 11149 19645
rect 11159 19631 11173 19645
rect 11183 19631 11197 19645
rect 11207 19631 11221 19645
rect 11231 19631 11245 19645
rect 11255 19631 11269 19645
rect 11279 19631 11293 19645
rect 11303 19631 11317 19645
rect 11327 19631 11341 19645
rect 11351 19631 11365 19645
rect 11375 19631 11389 19645
rect 11399 19631 11413 19645
rect 11423 19631 11437 19645
rect 11447 19631 11461 19645
rect 11471 19631 11485 19645
rect 11495 19631 11509 19645
rect 10919 19607 10933 19621
rect 10991 19607 11005 19621
rect 11567 19583 11581 19597
rect 11591 19583 11605 19597
rect 11615 19583 11629 19597
rect 11639 19583 11653 19597
rect 11111 19535 11125 19549
rect 11519 19535 11533 19549
rect 11543 19535 11557 19549
rect 10919 19511 10933 19525
rect 10943 19511 10957 19525
rect 10967 19511 10981 19525
rect 10991 19511 11005 19525
rect 11015 19511 11029 19525
rect 11039 19511 11053 19525
rect 11063 19511 11077 19525
rect 11087 19511 11101 19525
rect 11135 19487 11149 19501
rect 11159 19487 11173 19501
rect 11183 19487 11197 19501
rect 11207 19487 11221 19501
rect 11231 19487 11245 19501
rect 11255 19487 11269 19501
rect 11279 19487 11293 19501
rect 11303 19487 11317 19501
rect 11327 19487 11341 19501
rect 11351 19487 11365 19501
rect 11375 19487 11389 19501
rect 11399 19487 11413 19501
rect 11423 19487 11437 19501
rect 11447 19487 11461 19501
rect 11471 19487 11485 19501
rect 11495 19487 11509 19501
rect 11519 19487 11533 19501
rect 11543 19487 11557 19501
rect 11567 19487 11581 19501
rect 11591 19487 11605 19501
rect 11615 19487 11629 19501
rect 11639 19487 11653 19501
rect 10895 18431 10909 18445
rect 10919 18431 10933 18445
rect 10943 18431 10957 18445
rect 10967 18431 10981 18445
rect 10991 18431 11005 18445
rect 11015 18431 11029 18445
rect 11039 18431 11053 18445
rect 11063 18431 11077 18445
rect 11087 18431 11101 18445
rect 11111 18431 11125 18445
rect 11135 18431 11149 18445
rect 11159 18431 11173 18445
rect 11183 18431 11197 18445
rect 11231 18407 11245 18421
rect 11255 18407 11269 18421
rect 11279 18407 11293 18421
rect 11303 18407 11317 18421
rect 11327 18407 11341 18421
rect 11351 18407 11365 18421
rect 11375 18407 11389 18421
rect 11399 18407 11413 18421
rect 11423 18407 11437 18421
rect 11447 18407 11461 18421
rect 11471 18407 11485 18421
rect 11495 18407 11509 18421
rect 11519 18407 11533 18421
rect 11543 18407 11557 18421
rect 11567 18407 11581 18421
rect 11591 18407 11605 18421
rect 11615 18407 11629 18421
rect 11639 18407 11653 18421
rect 10871 18383 10885 18397
rect 11207 18383 11221 18397
rect 11399 18359 11413 18373
rect 10871 18335 10885 18349
rect 10895 18335 10909 18349
rect 10919 18335 10933 18349
rect 10943 18335 10957 18349
rect 10967 18335 10981 18349
rect 10991 18335 11005 18349
rect 11015 18335 11029 18349
rect 11039 18335 11053 18349
rect 11063 18335 11077 18349
rect 11087 18335 11101 18349
rect 11111 18335 11125 18349
rect 11135 18335 11149 18349
rect 11159 18335 11173 18349
rect 11183 18335 11197 18349
rect 11207 18335 11221 18349
rect 11231 18335 11245 18349
rect 11255 18335 11269 18349
rect 11279 18335 11293 18349
rect 11303 18335 11317 18349
rect 11327 18335 11341 18349
rect 11351 18335 11365 18349
rect 11375 18335 11389 18349
rect 11423 18311 11437 18325
rect 11447 18311 11461 18325
rect 11471 18311 11485 18325
rect 11495 18311 11509 18325
rect 11519 18311 11533 18325
rect 11543 18311 11557 18325
rect 11567 18311 11581 18325
rect 11591 18311 11605 18325
rect 11615 18311 11629 18325
rect 11639 18311 11653 18325
rect 10871 18167 10885 18181
rect 10895 18167 10909 18181
rect 10919 18167 10933 18181
rect 10943 18167 10957 18181
rect 10967 18167 10981 18181
rect 10991 18167 11005 18181
rect 11015 18167 11029 18181
rect 11039 18167 11053 18181
rect 11063 18167 11077 18181
rect 11087 18167 11101 18181
rect 11111 18167 11125 18181
rect 11135 18167 11149 18181
rect 11159 18167 11173 18181
rect 11183 18167 11197 18181
rect 11207 18167 11221 18181
rect 11231 18167 11245 18181
rect 11255 18167 11269 18181
rect 11279 18167 11293 18181
rect 11303 18167 11317 18181
rect 11327 18167 11341 18181
rect 11351 18167 11365 18181
rect 11375 18167 11389 18181
rect 11399 18167 11413 18181
rect 11423 18167 11437 18181
rect 11447 18167 11461 18181
rect 11471 18167 11485 18181
rect 11495 18167 11509 18181
rect 11519 18167 11533 18181
rect 11543 18167 11557 18181
rect 11567 18167 11581 18181
rect 11591 18167 11605 18181
rect 11615 18167 11629 18181
rect 11639 18167 11653 18181
rect 36767 18167 36781 18181
rect 36815 38807 36829 38821
rect 36839 38807 36853 38821
rect 36863 38807 36877 38821
rect 36887 38807 36901 38821
rect 36911 38807 36925 38821
rect 36935 38807 36949 38821
rect 36959 38807 36973 38821
rect 36983 38807 36997 38821
rect 37007 38807 37021 38821
rect 37031 38807 37045 38821
rect 37055 38807 37069 38821
rect 36815 18191 36829 18205
rect 36839 18191 36853 18205
rect 36863 18191 36877 18205
rect 36887 18191 36901 18205
rect 36911 18191 36925 18205
rect 41471 35879 41485 35893
rect 41471 35831 41485 35845
rect 41471 35735 41485 35749
rect 41471 35687 41485 35701
rect 41471 31151 41485 31165
rect 41471 31103 41485 31117
rect 41471 31007 41485 31021
rect 41471 30959 41485 30973
rect 41471 26327 41485 26341
rect 41495 26303 41509 26317
rect 41471 26279 41485 26293
rect 36959 18191 36973 18205
rect 36935 18143 36949 18157
rect 10871 18119 10885 18133
rect 36983 18119 36997 18133
rect 37007 18119 37021 18133
rect 10895 18095 10909 18109
rect 36791 18095 36805 18109
rect 36935 18095 36949 18109
rect 10919 18071 10933 18085
rect 36935 18071 36949 18085
rect 7535 18047 7549 18061
rect 10943 18047 10957 18061
rect 12287 18023 12301 18037
rect 13031 18023 13045 18037
rect 36287 18023 36301 18037
rect 37031 18023 37045 18037
rect 7535 17999 7549 18013
rect 10967 17999 10981 18013
rect 6575 16967 6589 16981
rect 6503 16895 6517 16909
rect 6527 16895 6541 16909
rect 6575 16919 6589 16933
rect 11663 17975 11677 17989
rect 12311 17975 12325 17989
rect 12359 17975 12373 17989
rect 13031 17975 13045 17989
rect 13631 17975 13645 17989
rect 13823 17975 13837 17989
rect 10369 17087 10383 17101
rect 10991 17927 11005 17941
rect 11015 17927 11029 17941
rect 11039 17927 11053 17941
rect 11063 17927 11077 17941
rect 11087 17927 11101 17941
rect 11111 17927 11125 17941
rect 11135 17927 11149 17941
rect 11159 17927 11173 17941
rect 11183 17927 11197 17941
rect 11207 17927 11221 17941
rect 11231 17927 11245 17941
rect 11255 17927 11269 17941
rect 11279 17927 11293 17941
rect 11303 17927 11317 17941
rect 11327 17927 11341 17941
rect 11351 17927 11365 17941
rect 11375 17927 11389 17941
rect 11399 17927 11413 17941
rect 11423 17927 11437 17941
rect 11447 17927 11461 17941
rect 11471 17927 11485 17941
rect 11495 17927 11509 17941
rect 11519 17927 11533 17941
rect 11543 17927 11557 17941
rect 11567 17927 11581 17941
rect 11591 17927 11605 17941
rect 11615 17927 11629 17941
rect 11639 17927 11653 17941
rect 11663 17927 11677 17941
rect 9911 17039 9925 17053
rect 9887 17015 9901 17029
rect 9863 16991 9877 17005
rect 9839 16967 9853 16981
rect 9815 16943 9829 16957
rect 9791 16919 9805 16933
rect 12335 17927 12349 17941
rect 12167 17903 12181 17917
rect 35543 17975 35557 17989
rect 36623 17975 36637 17989
rect 37055 17975 37069 17989
rect 37079 17975 37093 17989
rect 27839 17951 27853 17965
rect 14615 17927 14629 17941
rect 15167 17927 15181 17941
rect 15383 17927 15397 17941
rect 16127 17927 16141 17941
rect 16295 17927 16309 17941
rect 16679 17927 16693 17941
rect 16871 17927 16885 17941
rect 11183 16943 11197 16957
rect 11207 16943 11221 16957
rect 11231 16943 11245 16957
rect 11255 16943 11269 16957
rect 11279 16943 11293 16957
rect 11303 16943 11317 16957
rect 11327 16943 11341 16957
rect 11351 16943 11365 16957
rect 11375 16943 11389 16957
rect 11399 16943 11413 16957
rect 11423 16943 11437 16957
rect 11447 16943 11461 16957
rect 11471 16943 11485 16957
rect 11495 16943 11509 16957
rect 11519 16943 11533 16957
rect 11543 16943 11557 16957
rect 11567 16943 11581 16957
rect 11591 16943 11605 16957
rect 11615 16943 11629 16957
rect 11639 16943 11653 16957
rect 11663 16943 11677 16957
rect 11687 16943 11701 16957
rect 11711 16943 11725 16957
rect 13031 16943 13045 16957
rect 13631 16943 13645 16957
rect 13823 16943 13837 16957
rect 14543 16943 14557 16957
rect 14591 16943 14605 16957
rect 14615 16943 14629 16957
rect 15167 16943 15181 16957
rect 15383 16943 15397 16957
rect 16127 16943 16141 16957
rect 27599 17927 27613 17941
rect 36767 17927 36781 17941
rect 36791 17927 36805 17941
rect 36815 17927 36829 17941
rect 36839 17927 36853 17941
rect 36863 17927 36877 17941
rect 36887 17927 36901 17941
rect 36911 17927 36925 17941
rect 36935 17927 36949 17941
rect 36959 17927 36973 17941
rect 36983 17927 36997 17941
rect 37007 17927 37021 17941
rect 37031 17927 37045 17941
rect 37055 17927 37069 17941
rect 37079 17927 37093 17941
rect 17087 17903 17101 17917
rect 17831 17903 17845 17917
rect 17999 17903 18013 17917
rect 16895 17039 16909 17053
rect 27407 17903 27421 17917
rect 19103 17063 19117 17077
rect 20591 17063 20605 17077
rect 16871 16991 16885 17005
rect 16895 16991 16909 17005
rect 22103 17015 22117 17029
rect 22151 17015 22165 17029
rect 24431 16991 24445 17005
rect 25151 16967 25165 16981
rect 28130 16943 28144 16957
rect 36767 16943 36781 16957
rect 36791 16943 36805 16957
rect 36815 16943 36829 16957
rect 36839 16943 36853 16957
rect 36863 16943 36877 16957
rect 36887 16943 36901 16957
rect 37295 17135 37309 17149
rect 37655 17111 37669 17125
rect 37679 17087 37693 17101
rect 37703 17063 37717 17077
rect 37727 17039 37741 17053
rect 37751 17015 37765 17029
rect 37775 16991 37789 17005
rect 37799 16967 37813 16981
rect 37823 16943 37837 16957
rect 41471 16943 41485 16957
rect 9719 16895 9733 16909
rect 11183 16895 11197 16909
rect 11207 16895 11221 16909
rect 11231 16895 11245 16909
rect 13031 16895 13045 16909
rect 13631 16895 13645 16909
rect 13823 16895 13837 16909
rect 14543 16895 14557 16909
rect 14591 16895 14605 16909
rect 14615 16895 14629 16909
rect 15167 16895 15181 16909
rect 15383 16895 15397 16909
rect 16127 16895 16141 16909
rect 28154 16895 28168 16909
rect 36767 16895 36781 16909
rect 36791 16895 36805 16909
rect 36815 16895 36829 16909
rect 36839 16895 36853 16909
rect 36863 16895 36877 16909
rect 36887 16895 36901 16909
rect 37871 16895 37885 16909
rect 41471 16895 41485 16909
rect 9695 16871 9709 16885
rect 9671 16847 9685 16861
rect 11255 16847 11269 16861
rect 11279 16847 11293 16861
rect 11303 16847 11317 16861
rect 11735 16847 11749 16861
rect 9647 16823 9661 16837
rect 9623 16799 9637 16813
rect 11327 16799 11341 16813
rect 11351 16799 11365 16813
rect 11375 16799 11389 16813
rect 11759 16799 11773 16813
rect 13031 16799 13045 16813
rect 13631 16799 13645 16813
rect 14543 16823 14557 16837
rect 14591 16823 14605 16837
rect 30551 16871 30565 16885
rect 19079 16823 19093 16837
rect 19103 16823 19117 16837
rect 30527 16823 30541 16837
rect 30551 16823 30565 16837
rect 32183 16823 32197 16837
rect 32663 16823 32677 16837
rect 34151 16799 34165 16813
rect 36791 16823 36805 16837
rect 37895 16871 37909 16885
rect 37991 16847 38005 16861
rect 38015 16823 38029 16837
rect 38039 16799 38053 16813
rect 41471 16799 41485 16813
rect 9575 16775 9589 16789
rect 9599 16775 9613 16789
rect 9551 16751 9565 16765
rect 11399 16751 11413 16765
rect 11423 16751 11437 16765
rect 11807 16751 11821 16765
rect 13631 16751 13645 16765
rect 35663 16751 35677 16765
rect 36791 16775 36805 16789
rect 41471 16751 41485 16765
rect 9527 16727 9541 16741
rect 11447 16727 11461 16741
rect 11471 16727 11485 16741
rect 38063 16727 38077 16741
rect 38087 16727 38101 16741
rect 7535 16703 7549 16717
rect 9479 16703 9493 16717
rect 11495 16703 11509 16717
rect 11519 16703 11533 16717
rect 11783 16703 11797 16717
rect 11807 16703 11821 16717
rect 37967 16703 37981 16717
rect 37991 16703 38005 16717
rect 10175 16679 10189 16693
rect 11711 16679 11725 16693
rect 11735 16679 11749 16693
rect 9431 16655 9445 16669
rect 11567 16655 11581 16669
rect 11615 16655 11629 16669
rect 9743 16631 9757 16645
rect 9767 16631 9781 16645
rect 11543 16631 11557 16645
rect 11567 16631 11581 16645
rect 11687 16631 11701 16645
rect 11615 16607 11629 16621
rect 11663 16607 11677 16621
rect 11759 16655 11773 16669
rect 11783 16655 11797 16669
rect 37991 16655 38005 16669
rect 38135 16679 38149 16693
rect 10175 16559 10189 16573
rect 10346 16583 10360 16597
rect 11567 16583 11581 16597
rect 11591 16583 11605 16597
rect 11615 16559 11629 16573
rect 11639 16559 11653 16573
rect 7535 16535 7549 16549
rect 9431 16535 9445 16549
rect 9479 16535 9493 16549
rect 9527 16535 9541 16549
rect 9551 16535 9565 16549
rect 9575 16535 9589 16549
rect 9599 16535 9613 16549
rect 9623 16535 9637 16549
rect 9647 16535 9661 16549
rect 9671 16535 9685 16549
rect 9695 16535 9709 16549
rect 9719 16535 9733 16549
rect 9743 16535 9757 16549
rect 9767 16535 9781 16549
rect 9791 16535 9805 16549
rect 9815 16535 9829 16549
rect 9839 16535 9853 16549
rect 9863 16535 9877 16549
rect 9887 16535 9901 16549
rect 9911 16535 9925 16549
rect 10175 16535 10189 16549
rect 10295 16535 10309 16549
rect 10322 16535 10336 16549
rect 37655 16535 37669 16549
rect 37679 16535 37693 16549
rect 37703 16535 37717 16549
rect 37727 16535 37741 16549
rect 37751 16535 37765 16549
rect 37775 16535 37789 16549
rect 37799 16535 37813 16549
rect 37823 16535 37837 16549
rect 9431 16343 9445 16357
rect 9479 16343 9493 16357
rect 9527 16343 9541 16357
rect 9551 16343 9565 16357
rect 9599 16367 9613 16381
rect 9623 16367 9637 16381
rect 37871 16559 37885 16573
rect 37895 16559 37909 16573
rect 37967 16607 37981 16621
rect 37991 16607 38005 16621
rect 38015 16607 38029 16621
rect 38039 16607 38053 16621
rect 38063 16607 38077 16621
rect 38087 16607 38101 16621
rect 9671 16384 9685 16398
rect 9695 16384 9709 16398
rect 9719 16384 9733 16398
rect 9743 16384 9757 16398
rect 9767 16384 9781 16398
rect 9791 16384 9805 16398
rect 9815 16384 9829 16398
rect 9839 16384 9853 16398
rect 9863 16384 9877 16398
rect 9887 16384 9901 16398
rect 9911 16384 9925 16398
rect 37655 16385 37669 16399
rect 37679 16385 37693 16399
rect 37703 16385 37717 16399
rect 37727 16385 37741 16399
rect 37751 16385 37765 16399
rect 37775 16385 37789 16399
rect 37799 16385 37813 16399
rect 37823 16385 37837 16399
rect 37847 16385 37861 16399
rect 37871 16385 37885 16399
rect 37895 16385 37909 16399
rect 37919 16385 37933 16399
rect 37943 16385 37957 16399
rect 37967 16385 37981 16399
rect 37991 16385 38005 16399
rect 38015 16385 38029 16399
rect 9935 16360 9949 16374
rect 37631 16361 37645 16375
rect 9935 16336 9949 16350
rect 37631 16337 37645 16351
rect 38015 16337 38029 16351
rect 9935 16312 9949 16326
rect 37631 16313 37645 16327
rect 37823 16313 37837 16327
rect 37895 16313 37909 16327
rect 37919 16313 37933 16327
rect 37943 16313 37957 16327
rect 37967 16313 37981 16327
rect 37991 16313 38005 16327
rect 9431 16282 9445 16296
rect 9479 16281 9493 16295
rect 9527 16281 9541 16295
rect 9551 16281 9565 16295
rect 9599 16281 9613 16295
rect 9623 16281 9637 16295
rect 9671 16288 9685 16302
rect 9695 16288 9709 16302
rect 9719 16288 9733 16302
rect 9743 16288 9757 16302
rect 9767 16288 9781 16302
rect 9791 16288 9805 16302
rect 9815 16288 9829 16302
rect 9839 16288 9853 16302
rect 9863 16288 9877 16302
rect 9887 16288 9901 16302
rect 9911 16288 9925 16302
rect 37631 16289 37645 16303
rect 37775 16289 37789 16303
rect 9695 12719 9709 12733
rect 9719 12719 9733 12733
rect 9743 12719 9757 12733
rect 9767 12719 9781 12733
rect 9791 12719 9805 12733
rect 9815 12719 9829 12733
rect 9863 12695 9877 12709
rect 9695 12671 9709 12685
rect 9719 12671 9733 12685
rect 9743 12671 9757 12685
rect 9839 12647 9853 12661
rect 9887 12647 9901 12661
rect 37631 16265 37645 16279
rect 38135 16631 38149 16645
rect 38135 16583 38149 16597
rect 41375 16583 41389 16597
rect 41423 16583 41437 16597
rect 38135 16535 38149 16549
rect 41375 16535 41389 16549
rect 41423 16535 41437 16549
rect 37631 16241 37645 16255
rect 37871 16241 37885 16255
rect 37919 16241 37933 16255
rect 37943 16241 37957 16255
rect 37967 16241 37981 16255
rect 37991 16241 38005 16255
rect 38063 16241 38077 16255
rect 38087 16241 38101 16255
rect 37631 16217 37645 16231
rect 37655 16193 37669 16207
rect 37679 16193 37693 16207
rect 37703 16193 37717 16207
rect 37727 16193 37741 16207
rect 37751 16193 37765 16207
rect 37799 16193 37813 16207
rect 37847 16193 37861 16207
rect 37919 16193 37933 16207
rect 37943 16193 37957 16207
rect 37967 16193 37981 16207
rect 37991 16193 38005 16207
rect 38063 16193 38077 16207
rect 38087 16193 38101 16207
rect 7463 12599 7477 12613
rect 9431 12599 9445 12613
rect 9479 12599 9493 12613
rect 9527 12599 9541 12613
rect 9551 12599 9565 12613
rect 9599 12599 9613 12613
rect 9623 12599 9637 12613
rect 9647 12599 9661 12613
rect 9671 12599 9685 12613
rect 9695 12599 9709 12613
rect 9719 12599 9733 12613
rect 9743 12599 9757 12613
rect 9887 12599 9901 12613
rect 9935 12599 9949 12613
rect 9935 12575 9949 12589
rect 7463 12551 7477 12565
rect 9431 12551 9445 12565
rect 9479 12551 9493 12565
rect 9887 12551 9901 12565
rect 9935 12551 9949 12565
rect 9527 12503 9541 12517
rect 9551 12503 9565 12517
rect 9599 12503 9613 12517
rect 9623 12503 9637 12517
rect 9647 12503 9661 12517
rect 9671 12503 9685 12517
rect 9695 12503 9709 12517
rect 9719 12503 9733 12517
rect 9743 12503 9757 12517
rect 9767 12503 9781 12517
rect 9791 12503 9805 12517
rect 9815 12503 9829 12517
rect 9839 12503 9853 12517
rect 9863 12503 9877 12517
rect 9887 12503 9901 12517
rect 9935 12527 9949 12541
rect 37655 10319 37669 10333
rect 37679 10319 37693 10333
rect 37703 10319 37717 10333
rect 37631 10295 37645 10309
rect 37655 10271 37669 10285
rect 37679 10271 37693 10285
rect 37703 10271 37717 10285
rect 37655 10199 37669 10213
rect 37679 10199 37693 10213
rect 37703 10199 37717 10213
rect 37751 10199 37765 10213
rect 37799 10199 37813 10213
rect 37847 10199 37861 10213
rect 37919 10199 37933 10213
rect 37943 10199 37957 10213
rect 37967 10199 37981 10213
rect 37631 10175 37645 10189
rect 37631 10151 37645 10165
rect 37967 10151 37981 10165
rect 37655 10127 37669 10141
rect 37679 10127 37693 10141
rect 37703 10127 37717 10141
rect 37751 10127 37765 10141
rect 37799 10127 37813 10141
rect 37847 10127 37861 10141
rect 37919 10127 37933 10141
rect 37943 10127 37957 10141
rect 37655 8501 37669 8515
rect 37679 8501 37693 8515
rect 37703 8501 37717 8515
rect 37751 8501 37765 8515
rect 37799 8501 37813 8515
rect 9671 8478 9685 8492
rect 9695 8478 9709 8492
rect 9719 8478 9733 8492
rect 9743 8478 9757 8492
rect 9767 8478 9781 8492
rect 9791 8478 9805 8492
rect 9815 8478 9829 8492
rect 9839 8478 9853 8492
rect 9863 8478 9877 8492
rect 9887 8478 9901 8492
rect 9911 8478 9925 8492
rect 37631 8477 37645 8491
rect 9935 8454 9949 8468
rect 37679 8454 37693 8468
rect 9671 8430 9685 8444
rect 9935 8430 9949 8444
rect 37631 8430 37645 8444
rect 9935 8406 9949 8420
rect 37631 8406 37645 8420
rect 9695 8382 9709 8396
rect 9719 8382 9733 8396
rect 9935 8382 9949 8396
rect 37631 8382 37645 8396
rect 38063 8382 38077 8396
rect 9743 8358 9757 8372
rect 9767 8358 9781 8372
rect 9791 8358 9805 8372
rect 9815 8358 9829 8372
rect 9839 8358 9853 8372
rect 9863 8358 9877 8372
rect 9887 8358 9901 8372
rect 9911 8358 9925 8372
rect 37631 8358 37645 8372
rect 41447 12263 41461 12277
rect 41447 12215 41461 12229
rect 41471 12215 41485 12229
rect 41471 12167 41485 12181
rect 41471 12071 41485 12085
rect 41471 12023 41485 12037
rect 37631 8334 37645 8348
rect 37703 8334 37717 8348
rect 37751 8334 37765 8348
rect 37799 8334 37813 8348
rect 38063 8334 38077 8348
rect 9767 8303 9781 8317
rect 9791 8303 9805 8317
rect 9815 8303 9829 8317
rect 9839 8303 9853 8317
rect 9863 8303 9877 8317
rect 9887 8303 9901 8317
rect 9911 8303 9925 8317
rect 10295 8303 10309 8317
rect 10370 8303 10384 8317
rect 9935 8279 9949 8293
rect 9767 8255 9781 8269
rect 9791 8255 9805 8269
rect 9839 8255 9853 8269
rect 9959 8255 9973 8269
rect 9863 8231 9877 8245
rect 9983 8231 9997 8245
rect 9815 8183 9829 8197
rect 10007 8183 10021 8197
rect 9863 8159 9877 8173
rect 7463 8111 7477 8125
rect 9431 8111 9445 8125
rect 9527 8111 9541 8125
rect 9551 8111 9565 8125
rect 9599 8111 9613 8125
rect 9695 8111 9709 8125
rect 10031 8111 10045 8125
rect 10346 8231 10360 8245
rect 7463 8063 7477 8077
rect 9431 8063 9445 8077
rect 9527 8063 9541 8077
rect 9551 8063 9565 8077
rect 9599 8063 9613 8077
rect 9695 8063 9709 8077
rect 9863 8063 9877 8077
rect 9887 8063 9901 8077
rect 9911 8063 9925 8077
rect 9935 8063 9949 8077
rect 9959 8063 9973 8077
rect 9983 8063 9997 8077
rect 10007 8063 10021 8077
rect 10031 8063 10045 8077
rect 7463 7487 7477 7501
rect 9431 7487 9445 7501
rect 9527 7487 9541 7501
rect 9551 7487 9565 7501
rect 9599 7487 9613 7501
rect 9695 7487 9709 7501
rect 7463 7439 7477 7453
rect 9431 7439 9445 7453
rect 9527 7439 9541 7453
rect 9551 7439 9565 7453
rect 9599 7439 9613 7453
rect 9695 7439 9709 7453
rect 9599 6671 9613 6685
rect 9695 6671 9709 6685
rect 9887 6671 9901 6685
rect 9911 6671 9925 6685
rect 9935 6671 9949 6685
rect 11567 6743 11581 6757
rect 11711 6719 11725 6733
rect 15695 6695 15709 6709
rect 11687 6647 11701 6661
rect 11711 6647 11725 6661
rect 15815 6647 15829 6661
rect 19799 6647 19813 6661
rect 9599 6623 9613 6637
rect 9935 6623 9949 6637
rect 19967 6623 19981 6637
rect 9527 6599 9541 6613
rect 28055 6575 28069 6589
rect 7463 6551 7477 6565
rect 9527 6551 9541 6565
rect 28199 6551 28213 6565
rect 37655 8255 37669 8269
rect 37799 7487 37813 7501
rect 38063 7487 38077 7501
rect 37799 7439 37813 7453
rect 38063 7439 38077 7453
rect 38063 7343 38077 7357
rect 38063 7295 38077 7309
rect 32207 6551 32221 6565
rect 36455 6551 36469 6565
rect 9887 6527 9901 6541
rect 9911 6527 9925 6541
rect 11735 6527 11749 6541
rect 15863 6527 15877 6541
rect 19991 6527 20005 6541
rect 28247 6527 28261 6541
rect 7463 6503 7477 6517
rect 9695 6503 9709 6517
rect 11567 6503 11581 6517
rect 11687 6479 11701 6493
rect 11735 6479 11749 6493
rect 15695 6503 15709 6517
rect 15815 6479 15829 6493
rect 15863 6479 15877 6493
rect 19799 6479 19813 6493
rect 19967 6503 19981 6517
rect 19991 6479 20005 6493
rect 28055 6479 28069 6493
rect 28199 6479 28213 6493
rect 28247 6479 28261 6493
rect 32207 6503 32221 6517
rect 36311 6527 36325 6541
rect 36311 6479 36325 6493
rect 36455 6479 36469 6493
<< metal2 >>
rect 11520 41245 11532 41279
rect 11568 41245 11580 41279
rect 11592 41245 11604 41279
rect 11616 41245 11628 41399
rect 11640 41245 11652 41327
rect 11664 41245 11676 41327
rect 11688 41245 11700 41279
rect 15600 41269 15612 41423
rect 15648 41365 15660 41423
rect 15600 41149 15612 41255
rect 15624 41173 15636 41255
rect 15672 41197 15684 41351
rect 19728 41269 19740 41423
rect 19776 41293 19788 41423
rect 19800 41221 19812 41279
rect 19920 41245 19932 41423
rect 27984 41269 27996 41423
rect 28032 41389 28044 41423
rect 28056 41269 28068 41375
rect 28200 41293 28212 41399
rect 32112 41389 32124 41423
rect 32160 41341 32172 41423
rect 32328 41341 32340 41399
rect 36240 41389 36252 41423
rect 36264 41341 36276 41399
rect 36288 41365 36300 41399
rect 36432 41389 36444 41423
rect 41472 40573 41484 40607
rect 41448 40429 41460 40463
rect 41472 40429 41484 40463
rect 6504 40357 6516 40391
rect 7440 40357 7452 40391
rect 7536 40357 7548 40391
rect 11520 40357 11532 40391
rect 7536 39061 7548 39095
rect 11160 38821 11172 38855
rect 11184 38845 11196 38879
rect 11208 38797 11220 38903
rect 11232 38869 11244 38927
rect 11232 38797 11244 38831
rect 11256 38797 11268 38999
rect 11280 38989 11292 39095
rect 11304 39061 11316 39143
rect 11328 39061 11340 39143
rect 11352 39061 11364 39191
rect 11376 39061 11388 39215
rect 11400 39061 11412 39095
rect 11424 39061 11436 39239
rect 11472 39133 11484 39263
rect 11280 38797 11292 38855
rect 11304 38797 11316 38975
rect 11328 38797 11340 38999
rect 11352 38797 11364 38999
rect 11376 38797 11388 38999
rect 11400 38797 11412 38999
rect 11424 38797 11436 38999
rect 11448 38797 11460 38999
rect 11472 38797 11484 38999
rect 11496 38797 11508 39119
rect 11520 38797 11532 39287
rect 11592 39229 11604 39263
rect 11544 38797 11556 38999
rect 11568 38797 11580 38903
rect 11592 38797 11604 38903
rect 11616 38797 11628 39263
rect 11640 38797 11652 39263
rect 11664 38821 11676 39263
rect 11688 38893 11700 39263
rect 11712 38917 11724 39263
rect 11736 38941 11748 39263
rect 11760 38965 11772 39263
rect 11784 39133 11796 39263
rect 11832 39157 11844 39191
rect 11784 38965 11796 39095
rect 11808 38965 11820 39095
rect 11856 39085 11868 39119
rect 11832 38965 11844 39071
rect 11880 39061 11892 39095
rect 11856 38965 11868 39047
rect 11880 38965 11892 39023
rect 15600 38989 15612 39167
rect 12192 38917 12204 38975
rect 11784 38821 11796 38879
rect 12168 38773 12180 38903
rect 12312 38821 12324 38951
rect 15840 38796 15852 38975
rect 16080 38796 16092 39047
rect 17040 38796 17052 39095
rect 17232 38796 17244 39119
rect 18264 38796 18276 39167
rect 26256 38796 26268 39191
rect 26520 38796 26532 39215
rect 27240 38796 27252 39239
rect 29088 39109 29100 39215
rect 29064 38893 29076 39095
rect 29040 38796 29052 38879
rect 29256 38821 29268 39191
rect 29352 38965 29364 39119
rect 29376 39061 29388 39119
rect 29400 39061 29412 39191
rect 15840 38784 15853 38796
rect 16080 38784 16093 38796
rect 17040 38784 17053 38796
rect 17232 38784 17245 38796
rect 18264 38784 18279 38796
rect 26256 38784 26270 38796
rect 26520 38784 26534 38796
rect 27240 38784 27254 38796
rect 29040 38784 29053 38796
rect 12289 38773 12301 38783
rect 15841 38773 15853 38784
rect 16081 38773 16093 38784
rect 17041 38773 17053 38784
rect 17233 38773 17245 38784
rect 18267 38773 18279 38784
rect 26258 38773 26270 38784
rect 26522 38773 26534 38784
rect 27242 38773 27254 38784
rect 29041 38773 29053 38784
rect 29304 38796 29316 38927
rect 29424 38917 29436 39119
rect 29448 38989 29460 39119
rect 29472 38989 29484 39167
rect 36624 38941 36636 39167
rect 36648 38941 36660 39119
rect 36792 39061 36804 39143
rect 29400 38796 29412 38903
rect 29304 38784 29317 38796
rect 29400 38784 29413 38796
rect 29233 38773 29245 38783
rect 29305 38773 29317 38784
rect 29401 38773 29413 38784
rect 36624 38773 36636 38927
rect 36768 38797 36780 39047
rect 36816 38821 36828 38975
rect 36840 38821 36852 39095
rect 36864 38989 36876 39095
rect 36888 38965 36900 39071
rect 36864 38821 36876 38951
rect 36912 38941 36924 39023
rect 36888 38821 36900 38927
rect 36912 38821 36924 38879
rect 36936 38821 36948 38879
rect 36960 38821 36972 39023
rect 36984 38821 36996 38975
rect 37008 38917 37020 38951
rect 37008 38821 37020 38855
rect 37032 38821 37044 38903
rect 37056 38821 37068 38855
rect 11136 36013 11148 36095
rect 11160 35965 11172 36095
rect 11184 35965 11196 36095
rect 11208 35965 11220 36095
rect 11232 35965 11244 36095
rect 11256 35965 11268 36095
rect 11280 35965 11292 36095
rect 11304 35965 11316 36095
rect 11328 35965 11340 36095
rect 11352 35965 11364 36095
rect 11376 35965 11388 36095
rect 11400 35965 11412 36095
rect 11424 35965 11436 36095
rect 11448 35965 11460 36095
rect 11472 35965 11484 36095
rect 11496 35965 11508 36095
rect 11520 35965 11532 36095
rect 11544 35965 11556 36095
rect 11568 35965 11580 36095
rect 11592 35965 11604 36047
rect 11616 35965 11628 36071
rect 11640 35965 11652 36071
rect 41472 35845 41484 35879
rect 6528 35701 6540 35735
rect 41472 35701 41484 35735
rect 6504 35629 6516 35663
rect 11160 34837 11172 34919
rect 11184 34789 11196 34919
rect 11208 34789 11220 34919
rect 11232 34789 11244 34919
rect 11256 34789 11268 34919
rect 11280 34789 11292 34919
rect 11304 34789 11316 34919
rect 11328 34789 11340 34919
rect 11352 34789 11364 34919
rect 11376 34789 11388 34919
rect 11400 34789 11412 34919
rect 11424 34789 11436 34919
rect 11448 34789 11460 34919
rect 11472 34789 11484 34919
rect 11496 34789 11508 34919
rect 11520 34789 11532 34919
rect 11544 34789 11556 34919
rect 11568 34789 11580 34919
rect 11592 34789 11604 34919
rect 11616 34789 11628 34871
rect 11640 34789 11652 34895
rect 11184 33661 11196 33743
rect 11208 33613 11220 33743
rect 11232 33613 11244 33743
rect 11256 33613 11268 33743
rect 11280 33613 11292 33743
rect 11304 33613 11316 33743
rect 11328 33613 11340 33743
rect 11352 33613 11364 33743
rect 11376 33613 11388 33743
rect 11400 33613 11412 33743
rect 11424 33613 11436 33743
rect 11448 33613 11460 33743
rect 11472 33613 11484 33743
rect 11496 33613 11508 33743
rect 11520 33613 11532 33743
rect 11544 33613 11556 33743
rect 11568 33613 11580 33695
rect 11592 33613 11604 33719
rect 11616 33613 11628 33719
rect 11640 33613 11652 33719
rect 11208 32485 11220 32567
rect 11232 32437 11244 32567
rect 11256 32437 11268 32567
rect 11280 32437 11292 32567
rect 11304 32437 11316 32567
rect 11328 32437 11340 32567
rect 11352 32437 11364 32567
rect 11376 32437 11388 32519
rect 11400 32437 11412 32543
rect 11424 32437 11436 32543
rect 11448 32437 11460 32543
rect 11472 32437 11484 32543
rect 11496 32437 11508 32543
rect 11520 32437 11532 32543
rect 11544 32437 11556 32543
rect 11568 32437 11580 32543
rect 11592 32437 11604 32543
rect 11616 32437 11628 32543
rect 11640 32437 11652 32543
rect 11232 31309 11244 31391
rect 11256 31261 11268 31391
rect 11280 31261 11292 31391
rect 11304 31261 11316 31391
rect 11328 31261 11340 31391
rect 11352 31261 11364 31391
rect 11376 31261 11388 31391
rect 11400 31261 11412 31391
rect 11424 31261 11436 31391
rect 11448 31261 11460 31391
rect 11472 31261 11484 31391
rect 11496 31261 11508 31391
rect 11520 31261 11532 31391
rect 11544 31261 11556 31343
rect 11568 31261 11580 31367
rect 11592 31261 11604 31367
rect 11616 31261 11628 31367
rect 11640 31261 11652 31367
rect 41472 31117 41484 31151
rect 6504 30901 6516 30983
rect 6528 30901 6540 30935
rect 6552 30901 6564 31007
rect 41472 30973 41484 31007
rect 11256 30133 11268 30215
rect 11280 30085 11292 30215
rect 11304 30085 11316 30215
rect 11328 30085 11340 30215
rect 11352 30085 11364 30167
rect 11376 30085 11388 30191
rect 11400 30085 11412 30191
rect 11424 30085 11436 30191
rect 11448 30085 11460 30191
rect 11472 30085 11484 30191
rect 11496 30085 11508 30191
rect 11520 30085 11532 30191
rect 11544 30085 11556 30191
rect 11568 30085 11580 30191
rect 11592 30085 11604 30191
rect 11616 30085 11628 30191
rect 11640 30085 11652 30191
rect 11280 28957 11292 29039
rect 11304 28909 11316 29039
rect 11328 28909 11340 29039
rect 11352 28909 11364 29039
rect 11376 28909 11388 29039
rect 11400 28909 11412 29039
rect 11424 28909 11436 28991
rect 11448 28909 11460 29015
rect 11472 28909 11484 29015
rect 11496 28909 11508 29015
rect 11520 28909 11532 29015
rect 11544 28909 11556 29015
rect 11568 28909 11580 29015
rect 11592 28909 11604 29015
rect 11616 28909 11628 29015
rect 11640 28909 11652 29015
rect 11256 27757 11268 27791
rect 11280 27757 11292 27839
rect 11304 27757 11316 27863
rect 11328 27757 11340 27863
rect 11352 27757 11364 27863
rect 11376 27757 11388 27863
rect 11400 27757 11412 27863
rect 11424 27757 11436 27863
rect 11448 27805 11460 27863
rect 11472 27829 11484 27863
rect 11472 27733 11484 27767
rect 11496 27733 11508 27863
rect 11520 27733 11532 27863
rect 11544 27733 11556 27863
rect 11568 27733 11580 27863
rect 11592 27733 11604 27863
rect 11616 27733 11628 27863
rect 11640 27733 11652 27815
rect 11208 26581 11220 26615
rect 11232 26581 11244 26615
rect 11256 26581 11268 26639
rect 11280 26581 11292 26639
rect 11304 26605 11316 26639
rect 11328 26557 11340 26639
rect 11352 26557 11364 26639
rect 11376 26557 11388 26639
rect 11400 26557 11412 26639
rect 11424 26557 11436 26639
rect 11448 26557 11460 26639
rect 11472 26557 11484 26639
rect 11496 26557 11508 26639
rect 11520 26557 11532 26639
rect 11544 26557 11556 26639
rect 11568 26557 11580 26639
rect 11592 26557 11604 26639
rect 11616 26557 11628 26639
rect 11640 26557 11652 26639
rect 6504 26269 6516 26303
rect 6528 26269 6540 26303
rect 41472 26293 41484 26327
rect 41509 26304 41538 26316
rect 11160 25405 11172 25439
rect 11184 25405 11196 25487
rect 11208 25405 11220 25487
rect 11232 25405 11244 25487
rect 11256 25405 11268 25487
rect 11280 25405 11292 25487
rect 11304 25405 11316 25487
rect 11328 25405 11340 25487
rect 11352 25405 11364 25487
rect 11376 25405 11388 25487
rect 11400 25453 11412 25487
rect 11424 25381 11436 25487
rect 11448 25381 11460 25415
rect 11472 25381 11484 25463
rect 11496 25381 11508 25463
rect 11520 25381 11532 25463
rect 11544 25381 11556 25463
rect 11568 25381 11580 25463
rect 11592 25381 11604 25463
rect 11616 25381 11628 25463
rect 11640 25381 11652 25463
rect 11112 24229 11124 24263
rect 11136 24229 11148 24311
rect 11160 24229 11172 24311
rect 11184 24229 11196 24311
rect 11208 24277 11220 24311
rect 11232 24205 11244 24311
rect 11256 24205 11268 24311
rect 11280 24205 11292 24311
rect 11304 24205 11316 24311
rect 11328 24205 11340 24311
rect 11352 24205 11364 24311
rect 11376 24205 11388 24311
rect 11400 24205 11412 24311
rect 11424 24205 11436 24311
rect 11448 24205 11460 24311
rect 11472 24205 11484 24239
rect 11496 24205 11508 24287
rect 11520 24205 11532 24287
rect 11544 24205 11556 24287
rect 11568 24205 11580 24287
rect 11592 24205 11604 24287
rect 11616 24205 11628 24287
rect 11640 24205 11652 24287
rect 11064 23053 11076 23087
rect 11088 23053 11100 23135
rect 11112 23053 11124 23135
rect 11136 23053 11148 23135
rect 11160 23053 11172 23135
rect 11184 23053 11196 23135
rect 11208 23053 11220 23135
rect 11232 23053 11244 23135
rect 11256 23053 11268 23135
rect 11280 23053 11292 23135
rect 11304 23053 11316 23135
rect 11328 23053 11340 23135
rect 11352 23101 11364 23135
rect 11376 23029 11388 23135
rect 11400 23029 11412 23135
rect 11424 23029 11436 23135
rect 11448 23029 11460 23135
rect 11472 23029 11484 23135
rect 11496 23029 11508 23135
rect 11520 23029 11532 23135
rect 11544 23029 11556 23135
rect 11568 23029 11580 23063
rect 11592 23029 11604 23111
rect 11616 23029 11628 23111
rect 11640 23029 11652 23111
rect 11016 21877 11028 21911
rect 11040 21877 11052 21959
rect 11064 21877 11076 21959
rect 11088 21877 11100 21959
rect 11112 21877 11124 21959
rect 11136 21877 11148 21959
rect 11160 21877 11172 21959
rect 11184 21877 11196 21959
rect 11208 21877 11220 21959
rect 11232 21877 11244 21959
rect 11256 21877 11268 21959
rect 11280 21877 11292 21959
rect 11304 21877 11316 21959
rect 11328 21877 11340 21959
rect 11352 21877 11364 21959
rect 11376 21877 11388 21959
rect 11400 21877 11412 21959
rect 11424 21877 11436 21959
rect 11448 21925 11460 21959
rect 11472 21853 11484 21959
rect 11496 21853 11508 21959
rect 11520 21853 11532 21959
rect 11544 21853 11556 21959
rect 11568 21853 11580 21887
rect 11592 21853 11604 21935
rect 11616 21853 11628 21935
rect 11640 21853 11652 21935
rect 6504 21637 6516 21671
rect 6528 21637 6540 21671
rect 6552 21637 6564 21671
rect 6576 21637 6588 21671
rect 10968 20701 10980 20735
rect 10992 20701 11004 20783
rect 11016 20701 11028 20783
rect 11040 20701 11052 20735
rect 11064 20725 11076 20759
rect 11088 20677 11100 20759
rect 11112 20677 11124 20759
rect 11136 20677 11148 20759
rect 11160 20677 11172 20759
rect 11184 20677 11196 20759
rect 11208 20677 11220 20759
rect 11232 20677 11244 20759
rect 11256 20677 11268 20759
rect 11280 20677 11292 20759
rect 11304 20677 11316 20759
rect 11328 20677 11340 20759
rect 11352 20677 11364 20759
rect 11376 20677 11388 20759
rect 11400 20677 11412 20759
rect 11424 20677 11436 20759
rect 11448 20677 11460 20759
rect 11472 20677 11484 20759
rect 11496 20677 11508 20759
rect 11520 20677 11532 20759
rect 11544 20677 11556 20759
rect 11568 20677 11580 20759
rect 11592 20677 11604 20759
rect 11616 20677 11628 20759
rect 11640 20677 11652 20759
rect 10920 19525 10932 19607
rect 10944 19525 10956 19655
rect 10968 19525 10980 19655
rect 10992 19525 11004 19607
rect 11016 19525 11028 19631
rect 11040 19525 11052 19631
rect 11064 19525 11076 19631
rect 11088 19525 11100 19631
rect 11112 19549 11124 19631
rect 11136 19501 11148 19631
rect 11160 19501 11172 19631
rect 11184 19501 11196 19631
rect 11208 19501 11220 19631
rect 11232 19501 11244 19631
rect 11256 19501 11268 19631
rect 11280 19501 11292 19631
rect 11304 19501 11316 19631
rect 11328 19501 11340 19631
rect 11352 19501 11364 19631
rect 11376 19501 11388 19631
rect 11400 19501 11412 19631
rect 11424 19501 11436 19631
rect 11448 19501 11460 19631
rect 11472 19501 11484 19631
rect 11496 19501 11508 19631
rect 11520 19501 11532 19535
rect 11544 19501 11556 19535
rect 11568 19501 11580 19583
rect 11592 19501 11604 19583
rect 11616 19501 11628 19583
rect 11640 19501 11652 19583
rect 10872 18349 10884 18383
rect 10896 18349 10908 18431
rect 10920 18349 10932 18431
rect 10944 18349 10956 18431
rect 10968 18349 10980 18431
rect 10992 18349 11004 18431
rect 11016 18349 11028 18431
rect 11040 18349 11052 18431
rect 11064 18349 11076 18431
rect 11088 18349 11100 18431
rect 11112 18349 11124 18431
rect 11136 18349 11148 18431
rect 11160 18349 11172 18431
rect 11184 18349 11196 18431
rect 11208 18349 11220 18383
rect 11232 18349 11244 18407
rect 11256 18349 11268 18407
rect 11280 18349 11292 18407
rect 11304 18349 11316 18407
rect 11328 18349 11340 18407
rect 11352 18349 11364 18407
rect 11376 18349 11388 18407
rect 11400 18373 11412 18407
rect 11424 18325 11436 18407
rect 11448 18325 11460 18407
rect 11472 18325 11484 18407
rect 11496 18325 11508 18407
rect 11520 18325 11532 18407
rect 11544 18325 11556 18407
rect 11568 18325 11580 18407
rect 11592 18325 11604 18407
rect 11616 18325 11628 18407
rect 11640 18325 11652 18407
rect 10872 18133 10884 18167
rect 10896 18109 10908 18167
rect 10920 18085 10932 18167
rect 10944 18061 10956 18167
rect 7536 18013 7548 18047
rect 10968 18013 10980 18167
rect 10992 17941 11004 18167
rect 11016 17941 11028 18167
rect 11040 17941 11052 18167
rect 11064 17941 11076 18167
rect 11088 17941 11100 18167
rect 11112 17941 11124 18167
rect 11136 17941 11148 18167
rect 11160 17941 11172 18167
rect 11184 17941 11196 18167
rect 11208 17941 11220 18167
rect 11232 17941 11244 18167
rect 11256 17941 11268 18167
rect 11280 17941 11292 18167
rect 11304 17941 11316 18167
rect 11328 17941 11340 18167
rect 11352 17941 11364 18167
rect 11376 17941 11388 18167
rect 11400 17941 11412 18167
rect 11424 17941 11436 18167
rect 11448 17941 11460 18167
rect 11472 17941 11484 18167
rect 11496 17941 11508 18167
rect 11520 17941 11532 18167
rect 11544 17941 11556 18167
rect 11568 17941 11580 18167
rect 11592 17941 11604 18167
rect 11616 17941 11628 18167
rect 11640 17941 11652 18167
rect 11664 17941 11676 17975
rect 12168 17917 12180 18201
rect 12289 18180 12301 18201
rect 12313 18180 12325 18201
rect 12337 18180 12349 18201
rect 12361 18180 12373 18201
rect 13633 18180 13645 18201
rect 13825 18180 13837 18201
rect 14617 18180 14629 18201
rect 15169 18180 15181 18201
rect 15385 18180 15397 18201
rect 16129 18180 16141 18201
rect 16297 18180 16309 18201
rect 16681 18180 16693 18201
rect 16873 18180 16885 18201
rect 17089 18180 17101 18201
rect 17833 18180 17845 18201
rect 18001 18180 18013 18201
rect 27409 18180 27421 18201
rect 27601 18180 27613 18201
rect 27841 18180 27853 18201
rect 35545 18180 35557 18201
rect 36289 18180 36301 18201
rect 12288 18168 12301 18180
rect 12312 18168 12325 18180
rect 12336 18168 12349 18180
rect 12360 18168 12373 18180
rect 13632 18168 13645 18180
rect 13824 18168 13837 18180
rect 14616 18168 14629 18180
rect 15168 18168 15181 18180
rect 15384 18168 15397 18180
rect 16128 18168 16141 18180
rect 16296 18168 16309 18180
rect 16680 18168 16693 18180
rect 16872 18168 16885 18180
rect 17088 18168 17101 18180
rect 17832 18168 17845 18180
rect 18000 18168 18013 18180
rect 27408 18168 27421 18180
rect 27600 18168 27613 18180
rect 27840 18168 27853 18180
rect 35544 18168 35557 18180
rect 36288 18168 36301 18180
rect 12288 18037 12300 18168
rect 12312 17989 12324 18168
rect 12336 17941 12348 18168
rect 12360 17989 12372 18168
rect 13032 17989 13044 18023
rect 13632 17989 13644 18168
rect 13824 17989 13836 18168
rect 14616 17941 14628 18168
rect 15168 17941 15180 18168
rect 15384 17941 15396 18168
rect 16128 17941 16140 18168
rect 16296 17941 16308 18168
rect 16680 17941 16692 18168
rect 16872 17941 16884 18168
rect 17088 17917 17100 18168
rect 17832 17917 17844 18168
rect 18000 17917 18012 18168
rect 27408 17917 27420 18168
rect 27600 17941 27612 18168
rect 27840 17965 27852 18168
rect 35544 17989 35556 18168
rect 36288 18037 36300 18168
rect 36624 17989 36636 18201
rect 36768 17941 36780 18167
rect 36792 17941 36804 18095
rect 36816 17941 36828 18191
rect 36840 17941 36852 18191
rect 36864 17941 36876 18191
rect 36888 17941 36900 18191
rect 36912 17941 36924 18191
rect 36936 18109 36948 18143
rect 36936 17941 36948 18071
rect 36960 17941 36972 18191
rect 36984 17941 36996 18119
rect 37008 17941 37020 18119
rect 37032 17941 37044 18023
rect 37056 17941 37068 17975
rect 37080 17941 37092 17975
rect 6504 16909 6516 16943
rect 6528 16909 6540 16943
rect 6576 16933 6588 16967
rect 7536 16549 7548 16703
rect 9432 16549 9444 16655
rect 9480 16549 9492 16703
rect 9528 16549 9540 16727
rect 9552 16549 9564 16751
rect 9576 16549 9588 16775
rect 9600 16549 9612 16775
rect 9624 16549 9636 16799
rect 9648 16549 9660 16823
rect 9672 16549 9684 16847
rect 9696 16549 9708 16871
rect 9720 16549 9732 16895
rect 9744 16549 9756 16631
rect 9768 16549 9780 16631
rect 9792 16549 9804 16919
rect 9816 16549 9828 16943
rect 9840 16549 9852 16967
rect 9864 16549 9876 16991
rect 9888 16549 9900 17015
rect 9912 16549 9924 17039
rect 10176 16573 10188 16679
rect 10309 16535 10311 16549
rect 10176 16504 10188 16535
rect 10299 16504 10311 16535
rect 10323 16504 10335 16535
rect 10347 16504 10359 16583
rect 10371 16504 10383 17087
rect 16896 17005 16908 17039
rect 11184 16909 11196 16943
rect 11208 16909 11220 16943
rect 11232 16909 11244 16943
rect 11256 16861 11268 16943
rect 11280 16861 11292 16943
rect 11304 16861 11316 16943
rect 11328 16813 11340 16943
rect 11352 16813 11364 16943
rect 11376 16813 11388 16943
rect 11400 16765 11412 16943
rect 11424 16765 11436 16943
rect 11448 16741 11460 16943
rect 11472 16741 11484 16943
rect 11496 16717 11508 16943
rect 11520 16717 11532 16943
rect 11544 16645 11556 16943
rect 11568 16669 11580 16943
rect 11568 16597 11580 16631
rect 11592 16597 11604 16943
rect 11616 16669 11628 16943
rect 11616 16573 11628 16607
rect 11640 16573 11652 16943
rect 11664 16621 11676 16943
rect 11688 16645 11700 16943
rect 11712 16693 11724 16943
rect 13032 16909 13044 16943
rect 13632 16909 13644 16943
rect 13824 16909 13836 16943
rect 14544 16909 14556 16943
rect 14592 16909 14604 16943
rect 14616 16909 14628 16943
rect 15168 16909 15180 16943
rect 15384 16909 15396 16943
rect 16128 16909 16140 16943
rect 11736 16693 11748 16847
rect 11760 16669 11772 16799
rect 11808 16717 11820 16751
rect 11784 16669 11796 16703
rect 13032 16548 13044 16799
rect 13632 16765 13644 16799
rect 14544 16548 14556 16823
rect 14592 16548 14604 16823
rect 16872 16548 16884 16991
rect 19104 16837 19116 17063
rect 13032 16536 13047 16548
rect 14544 16536 14559 16548
rect 13035 16504 13047 16536
rect 14547 16504 14559 16536
rect 14583 16536 14604 16548
rect 16863 16536 16884 16548
rect 19080 16548 19092 16823
rect 20592 16548 20604 17063
rect 22104 16548 22116 17015
rect 22152 16548 22164 17015
rect 24432 16548 24444 16991
rect 19080 16536 19095 16548
rect 20592 16536 20607 16548
rect 22104 16536 22119 16548
rect 14583 16504 14595 16536
rect 16863 16504 16875 16536
rect 19083 16504 19095 16536
rect 20595 16504 20607 16536
rect 22107 16504 22119 16536
rect 22143 16536 22164 16548
rect 24423 16536 24444 16548
rect 25152 16548 25164 16967
rect 25152 16536 25167 16548
rect 22143 16504 22155 16536
rect 24423 16504 24435 16536
rect 25155 16504 25167 16536
rect 28131 16504 28143 16943
rect 36768 16909 36780 16943
rect 36792 16909 36804 16943
rect 36816 16909 36828 16943
rect 36840 16909 36852 16943
rect 36864 16909 36876 16943
rect 36888 16909 36900 16943
rect 28155 16504 28167 16895
rect 30552 16837 30564 16871
rect 30528 16548 30540 16823
rect 32184 16548 32196 16823
rect 32664 16548 32676 16823
rect 30519 16536 30540 16548
rect 32175 16536 32196 16548
rect 32655 16536 32676 16548
rect 34152 16548 34164 16799
rect 36792 16789 36804 16823
rect 35664 16548 35676 16751
rect 34152 16536 34167 16548
rect 30519 16504 30531 16536
rect 32175 16504 32187 16536
rect 32655 16504 32667 16536
rect 34155 16504 34167 16536
rect 35655 16536 35676 16548
rect 35655 16504 35667 16536
rect 37296 16504 37308 17135
rect 37656 16549 37668 17111
rect 37680 16549 37692 17087
rect 37704 16549 37716 17063
rect 37728 16549 37740 17039
rect 37752 16549 37764 17015
rect 37776 16549 37788 16991
rect 37800 16549 37812 16967
rect 37824 16549 37836 16943
rect 41472 16909 41484 16943
rect 37872 16573 37884 16895
rect 37896 16573 37908 16871
rect 37992 16717 38004 16847
rect 37968 16621 37980 16703
rect 37992 16621 38004 16655
rect 38016 16621 38028 16823
rect 38040 16621 38052 16799
rect 41472 16765 41484 16799
rect 38064 16621 38076 16727
rect 38088 16621 38100 16727
rect 38136 16645 38148 16679
rect 38136 16549 38148 16583
rect 41376 16549 41388 16583
rect 41424 16549 41436 16583
rect 9432 16296 9444 16343
rect 9480 16295 9492 16343
rect 9528 16295 9540 16343
rect 9552 16295 9564 16343
rect 9600 16295 9612 16367
rect 9624 16295 9636 16367
rect 9672 16302 9684 16384
rect 9696 16302 9708 16384
rect 9720 16302 9732 16384
rect 9744 16302 9756 16384
rect 9768 16302 9780 16384
rect 9792 16302 9804 16384
rect 9816 16302 9828 16384
rect 9840 16302 9852 16384
rect 9864 16302 9876 16384
rect 9888 16302 9900 16384
rect 9912 16302 9924 16384
rect 9949 16361 9960 16373
rect 37609 16361 37631 16373
rect 9949 16337 9960 16349
rect 37609 16337 37631 16349
rect 9949 16313 9960 16325
rect 37609 16313 37631 16325
rect 37609 16289 37631 16301
rect 37609 16265 37631 16277
rect 37609 16241 37631 16253
rect 37609 16217 37631 16229
rect 37656 16207 37668 16385
rect 37680 16207 37692 16385
rect 37704 16207 37716 16385
rect 37728 16207 37740 16385
rect 37752 16207 37764 16385
rect 37776 16303 37788 16385
rect 37800 16207 37812 16385
rect 37824 16327 37836 16385
rect 37848 16207 37860 16385
rect 37872 16255 37884 16385
rect 37896 16327 37908 16385
rect 37920 16327 37932 16385
rect 37944 16327 37956 16385
rect 37968 16327 37980 16385
rect 37992 16327 38004 16385
rect 38016 16351 38028 16385
rect 37920 16207 37932 16241
rect 37944 16207 37956 16241
rect 37968 16207 37980 16241
rect 37992 16207 38004 16241
rect 38064 16207 38076 16241
rect 38088 16207 38100 16241
rect 9696 12685 9708 12719
rect 9720 12685 9732 12719
rect 9744 12685 9756 12719
rect 7464 12565 7476 12599
rect 9432 12565 9444 12599
rect 9480 12565 9492 12599
rect 9528 12517 9540 12599
rect 9552 12517 9564 12599
rect 9600 12517 9612 12599
rect 9624 12517 9636 12599
rect 9648 12517 9660 12599
rect 9672 12517 9684 12599
rect 9696 12517 9708 12599
rect 9720 12517 9732 12599
rect 9744 12517 9756 12599
rect 9768 12517 9780 12719
rect 9792 12517 9804 12719
rect 9816 12517 9828 12719
rect 9840 12517 9852 12647
rect 9864 12517 9876 12695
rect 9888 12613 9900 12647
rect 9949 12600 9960 12612
rect 9949 12576 9960 12588
rect 9949 12552 9960 12564
rect 9888 12517 9900 12551
rect 9949 12528 9960 12540
rect 41448 12229 41460 12263
rect 41472 12181 41484 12215
rect 41472 12037 41484 12071
rect 37609 10296 37631 10308
rect 37656 10285 37668 10319
rect 37680 10285 37692 10319
rect 37704 10285 37716 10319
rect 37609 10176 37631 10188
rect 37609 10152 37631 10164
rect 37656 10141 37668 10199
rect 37680 10141 37692 10199
rect 37704 10141 37716 10199
rect 37752 10141 37764 10199
rect 37800 10141 37812 10199
rect 37848 10141 37860 10199
rect 37920 10141 37932 10199
rect 37944 10141 37956 10199
rect 37968 10165 37980 10199
rect 37609 8479 37631 8491
rect 9672 8444 9684 8478
rect 9696 8396 9708 8478
rect 9720 8396 9732 8478
rect 9744 8372 9756 8478
rect 9768 8372 9780 8478
rect 9792 8372 9804 8478
rect 9816 8372 9828 8478
rect 9840 8372 9852 8478
rect 9864 8372 9876 8478
rect 9888 8372 9900 8478
rect 9912 8372 9924 8478
rect 9949 8455 9960 8467
rect 9949 8431 9960 8443
rect 37609 8431 37631 8443
rect 9949 8407 9960 8419
rect 37609 8407 37631 8419
rect 9949 8383 9960 8395
rect 37609 8383 37631 8395
rect 37609 8359 37631 8371
rect 37609 8335 37631 8347
rect 10299 8317 10311 8334
rect 10309 8303 10311 8317
rect 9768 8269 9780 8303
rect 9792 8269 9804 8303
rect 9816 8197 9828 8303
rect 9840 8269 9852 8303
rect 9864 8245 9876 8303
rect 7464 8077 7476 8111
rect 9432 8077 9444 8111
rect 9528 8077 9540 8111
rect 9552 8077 9564 8111
rect 9600 8077 9612 8111
rect 9696 8077 9708 8111
rect 9864 8077 9876 8159
rect 9888 8077 9900 8303
rect 9912 8077 9924 8303
rect 9936 8077 9948 8279
rect 9960 8077 9972 8255
rect 10347 8245 10359 8334
rect 10371 8317 10383 8334
rect 37656 8269 37668 8501
rect 37680 8468 37692 8501
rect 37704 8348 37716 8501
rect 37752 8348 37764 8501
rect 37800 8348 37812 8501
rect 38064 8348 38076 8382
rect 9984 8077 9996 8231
rect 10008 8077 10020 8183
rect 10032 8077 10044 8111
rect 7464 7453 7476 7487
rect 9432 7453 9444 7487
rect 9528 7453 9540 7487
rect 9552 7453 9564 7487
rect 9600 7453 9612 7487
rect 9696 7453 9708 7487
rect 37800 7453 37812 7487
rect 38064 7453 38076 7487
rect 38064 7309 38076 7343
rect 9600 6637 9612 6671
rect 9528 6565 9540 6599
rect 7464 6517 7476 6551
rect 9696 6517 9708 6671
rect 9888 6541 9900 6671
rect 9912 6541 9924 6671
rect 9936 6637 9948 6671
rect 11568 6517 11580 6743
rect 11712 6661 11724 6719
rect 11688 6493 11700 6647
rect 11736 6493 11748 6527
rect 15696 6517 15708 6695
rect 15816 6493 15828 6647
rect 15864 6493 15876 6527
rect 19800 6493 19812 6647
rect 19968 6517 19980 6623
rect 19992 6493 20004 6527
rect 28056 6493 28068 6575
rect 28200 6493 28212 6551
rect 28248 6493 28260 6527
rect 32208 6517 32220 6551
rect 36312 6493 36324 6527
rect 36456 6493 36468 6551
<< metal4 >>
rect 6702 46264 8262 47824
rect 10830 46264 12390 47824
rect 14958 46264 16518 47824
rect 19086 46264 20646 47824
rect 23214 46264 24774 47824
rect 27342 46264 28902 47824
rect 31470 46264 33030 47824
rect 35598 46264 37158 47824
rect 39726 46264 41286 47824
rect 78 39726 1638 41286
rect 46350 39726 47910 41286
rect 78 34996 1638 36556
rect 46350 34996 47910 36556
rect 78 30266 1638 31826
rect 46350 30266 47910 31826
rect 78 25536 1638 27096
rect 46350 25536 47910 27096
rect 78 20806 1638 22366
rect 46350 20806 47910 22366
rect 78 16076 1638 17636
rect 46350 16076 47910 17636
rect 78 11346 1638 12906
rect 46350 11346 47910 12906
rect 78 6616 1638 8176
rect 46350 6616 47910 8176
rect 6702 78 8262 1638
rect 10830 78 12390 1638
rect 14958 78 16518 1638
rect 19086 78 20646 1638
rect 23214 78 24774 1638
rect 27342 78 28902 1638
rect 31470 78 33030 1638
rect 35598 78 37158 1638
rect 39726 78 41286 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 0 -1 0 47902
box 0 0 6450 6450
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform 0 -1 6536 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform 0 -1 6622 1 0 41452
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 8342 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform 0 -1 8428 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform 0 -1 8514 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform 0 -1 8600 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform 0 -1 8686 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform 0 -1 8772 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform 0 -1 8858 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform 0 -1 8944 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform 0 -1 9030 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform 0 -1 9116 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform 0 -1 9202 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform 0 -1 9288 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform 0 -1 9374 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform 0 -1 9460 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform 0 -1 9546 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform 0 -1 9632 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform 0 -1 9718 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform 0 -1 9804 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform 0 -1 9890 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform 0 -1 9976 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform 0 -1 10062 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform 0 -1 10148 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform 0 -1 10234 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform 0 -1 10320 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform 0 -1 10406 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform 0 -1 10492 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform 0 -1 10578 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform 0 -1 10664 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform 0 -1 10750 1 0 41452
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 12470 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform 0 -1 12556 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform 0 -1 12642 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform 0 -1 12728 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform 0 -1 12814 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform 0 -1 12900 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform 0 -1 12986 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform 0 -1 13072 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform 0 -1 13158 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform 0 -1 13244 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform 0 -1 13330 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform 0 -1 13416 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform 0 -1 13502 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform 0 -1 13588 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform 0 -1 13674 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform 0 -1 13760 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform 0 -1 13846 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform 0 -1 13932 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform 0 -1 14018 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform 0 -1 14104 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform 0 -1 14190 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform 0 -1 14276 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform 0 -1 14362 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform 0 -1 14448 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform 0 -1 14534 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform 0 -1 14620 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform 0 -1 14706 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform 0 -1 14792 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform 0 -1 14878 1 0 41452
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 16598 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform 0 -1 16684 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform 0 -1 16770 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform 0 -1 16856 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform 0 -1 16942 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform 0 -1 17028 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform 0 -1 17114 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform 0 -1 17200 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform 0 -1 17286 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform 0 -1 17372 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform 0 -1 17458 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform 0 -1 17544 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform 0 -1 17630 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform 0 -1 17716 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform 0 -1 17802 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform 0 -1 17888 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform 0 -1 17974 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform 0 -1 18060 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform 0 -1 18146 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform 0 -1 18232 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform 0 -1 18318 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform 0 -1 18404 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform 0 -1 18490 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform 0 -1 18576 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform 0 -1 18662 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform 0 -1 18748 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform 0 -1 18834 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform 0 -1 18920 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform 0 -1 19006 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 20726 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform 0 -1 20812 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform 0 -1 20898 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform 0 -1 20984 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform 0 -1 21070 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform 0 -1 21156 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform 0 -1 21242 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform 0 -1 21328 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform 0 -1 21414 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform 0 -1 21500 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform 0 -1 21586 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform 0 -1 21672 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform 0 -1 21758 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform 0 -1 21844 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform 0 -1 21930 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform 0 -1 22016 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform 0 -1 22102 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform 0 -1 22188 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform 0 -1 22274 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform 0 -1 22360 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform 0 -1 22446 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform 0 -1 22532 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform 0 -1 22618 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform 0 -1 22704 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform 0 -1 22790 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform 0 -1 22876 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform 0 -1 22962 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform 0 -1 23048 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform 0 -1 23134 1 0 41452
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 24854 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform 0 -1 24940 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform 0 -1 25026 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform 0 -1 25112 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform 0 -1 25198 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform 0 -1 25284 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform 0 -1 25370 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform 0 -1 25456 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform 0 -1 25542 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform 0 -1 25628 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform 0 -1 25714 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform 0 -1 25800 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform 0 -1 25886 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform 0 -1 25972 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform 0 -1 26058 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform 0 -1 26144 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform 0 -1 26230 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform 0 -1 26316 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform 0 -1 26402 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform 0 -1 26488 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform 0 -1 26574 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform 0 -1 26660 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform 0 -1 26746 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform 0 -1 26832 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform 0 -1 26918 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform 0 -1 27004 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 27090 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 27176 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 27262 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 28982 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 29068 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 29154 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 29240 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 29326 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 29412 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 29498 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 29584 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 29670 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 29756 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 29842 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 29928 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 30014 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 30100 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 30186 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 30272 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 30358 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 30444 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 0 -1 30530 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 0 -1 30616 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 0 -1 30702 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 0 -1 30788 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 0 -1 30874 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 0 -1 30960 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 0 -1 31046 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 0 -1 31132 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 0 -1 31218 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 0 -1 31304 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 0 -1 31390 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 33110 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 0 -1 33196 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 0 -1 33282 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 0 -1 33368 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 0 -1 33454 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 33540 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 33626 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 33712 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 33798 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 33884 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 33970 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 34056 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 34142 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 34228 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 34314 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 34400 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 34486 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 34572 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 34658 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 34744 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 34830 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 34916 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 35002 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 35088 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 35174 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 35260 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 35346 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 35432 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 35518 1 0 41452
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 37238 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 37324 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 37410 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 37496 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 37582 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 37668 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 37754 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 37840 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 37926 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 38012 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 38098 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 38184 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 38270 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 38356 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 38442 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 38528 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 38614 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 38700 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 38786 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 38872 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 38958 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 39044 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 39130 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 39216 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 39302 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 39388 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 39474 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 39560 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 39646 1 0 41452
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 41366 1 0 41452
box 0 0 6450 1720
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 41452 1 0 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 41538 1 0 41452
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 47988 0 -1 47902
box 0 0 6450 6450
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 6450 0 -1 41452
box 0 0 6450 86
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 6450 0 -1 41366
box 0 0 6450 1720
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 6450 0 -1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 6450 0 -1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 6450 0 -1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 6450 0 -1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 6450 0 -1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 6450 0 -1 39216
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 6450 0 -1 39130
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 6450 0 -1 39044
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 6450 0 -1 38958
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 6450 0 -1 38872
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 6450 0 -1 38786
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 1 0 41538 0 1 41366
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 41538 0 1 39646
box 0 0 6450 1720
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 1 0 41538 0 1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 1 0 41538 0 1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 1 0 41538 0 1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 1 0 41538 0 1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 1 0 41538 0 1 39216
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 1 0 41538 0 1 39130
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 1 0 41538 0 1 39044
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 1 0 41538 0 1 38958
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 1 0 41538 0 1 38872
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 1 0 41538 0 1 38786
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 6450 0 -1 38700
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 6450 0 -1 38614
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 6450 0 -1 38528
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform -1 0 6450 0 -1 38442
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform -1 0 6450 0 -1 38356
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform -1 0 6450 0 -1 38270
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform -1 0 6450 0 -1 38184
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform -1 0 6450 0 -1 38098
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform -1 0 6450 0 -1 38012
box 0 0 6450 86
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform -1 0 6450 0 -1 37926
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform -1 0 6450 0 -1 37840
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform -1 0 6450 0 -1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform -1 0 6450 0 -1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform -1 0 6450 0 -1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform -1 0 6450 0 -1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform -1 0 6450 0 -1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform -1 0 6450 0 -1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform -1 0 6450 0 -1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform -1 0 6450 0 -1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform -1 0 6450 0 -1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform -1 0 6450 0 -1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform -1 0 6450 0 -1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform -1 0 6450 0 -1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform -1 0 6450 0 -1 36722
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 6450 0 -1 36636
box 0 0 6450 1720
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform -1 0 6450 0 -1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform -1 0 6450 0 -1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform -1 0 6450 0 -1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform -1 0 6450 0 -1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform -1 0 6450 0 -1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform -1 0 6450 0 -1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform -1 0 6450 0 -1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform -1 0 6450 0 -1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform -1 0 6450 0 -1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform -1 0 6450 0 -1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform -1 0 6450 0 -1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform -1 0 6450 0 -1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform -1 0 6450 0 -1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform -1 0 6450 0 -1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform -1 0 6450 0 -1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform -1 0 6450 0 -1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform -1 0 6450 0 -1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform -1 0 6450 0 -1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform -1 0 6450 0 -1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform -1 0 6450 0 -1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform -1 0 6450 0 -1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform -1 0 6450 0 -1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform -1 0 6450 0 -1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform -1 0 6450 0 -1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform -1 0 6450 0 -1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform -1 0 6450 0 -1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform -1 0 6450 0 -1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform -1 0 6450 0 -1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform -1 0 6450 0 -1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform -1 0 6450 0 -1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform -1 0 6450 0 -1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform -1 0 6450 0 -1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform -1 0 6450 0 -1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform -1 0 6450 0 -1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform -1 0 6450 0 -1 31992
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 6450 0 -1 31906
box 0 0 6450 1720
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform -1 0 6450 0 -1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform -1 0 6450 0 -1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform -1 0 6450 0 -1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform -1 0 6450 0 -1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform -1 0 6450 0 -1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform -1 0 6450 0 -1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform -1 0 6450 0 -1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform -1 0 6450 0 -1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform -1 0 6450 0 -1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform -1 0 6450 0 -1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform -1 0 6450 0 -1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform -1 0 6450 0 -1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform -1 0 6450 0 -1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform -1 0 6450 0 -1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_788
timestamp 1300117811
transform -1 0 6450 0 -1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_789
timestamp 1300117811
transform -1 0 6450 0 -1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_790
timestamp 1300117811
transform -1 0 6450 0 -1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_791
timestamp 1300117811
transform -1 0 6450 0 -1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_792
timestamp 1300117811
transform -1 0 6450 0 -1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_793
timestamp 1300117811
transform -1 0 6450 0 -1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_794
timestamp 1300117811
transform -1 0 6450 0 -1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_795
timestamp 1300117811
transform -1 0 6450 0 -1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_796
timestamp 1300117811
transform -1 0 6450 0 -1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_797
timestamp 1300117811
transform -1 0 6450 0 -1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_798
timestamp 1300117811
transform -1 0 6450 0 -1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_799
timestamp 1300117811
transform -1 0 6450 0 -1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_800
timestamp 1300117811
transform -1 0 6450 0 -1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_801
timestamp 1300117811
transform -1 0 6450 0 -1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_802
timestamp 1300117811
transform -1 0 6450 0 -1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_803
timestamp 1300117811
transform -1 0 6450 0 -1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_804
timestamp 1300117811
transform -1 0 6450 0 -1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_805
timestamp 1300117811
transform -1 0 6450 0 -1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_806
timestamp 1300117811
transform -1 0 6450 0 -1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_807
timestamp 1300117811
transform -1 0 6450 0 -1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_808
timestamp 1300117811
transform -1 0 6450 0 -1 27262
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 6450 0 -1 27176
box 0 0 6450 1720
use fillpp_mt fillpp_mt_809
timestamp 1300117811
transform -1 0 6450 0 -1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_810
timestamp 1300117811
transform -1 0 6450 0 -1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_811
timestamp 1300117811
transform -1 0 6450 0 -1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_812
timestamp 1300117811
transform -1 0 6450 0 -1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_813
timestamp 1300117811
transform -1 0 6450 0 -1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_814
timestamp 1300117811
transform -1 0 6450 0 -1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_815
timestamp 1300117811
transform -1 0 6450 0 -1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_816
timestamp 1300117811
transform -1 0 6450 0 -1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_817
timestamp 1300117811
transform -1 0 6450 0 -1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_818
timestamp 1300117811
transform -1 0 6450 0 -1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_819
timestamp 1300117811
transform -1 0 6450 0 -1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_820
timestamp 1300117811
transform -1 0 6450 0 -1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_821
timestamp 1300117811
transform -1 0 6450 0 -1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_822
timestamp 1300117811
transform -1 0 6450 0 -1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_823
timestamp 1300117811
transform -1 0 6450 0 -1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_824
timestamp 1300117811
transform -1 0 6450 0 -1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_825
timestamp 1300117811
transform -1 0 6450 0 -1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_826
timestamp 1300117811
transform -1 0 6450 0 -1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_827
timestamp 1300117811
transform -1 0 6450 0 -1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_828
timestamp 1300117811
transform -1 0 6450 0 -1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_829
timestamp 1300117811
transform -1 0 6450 0 -1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_830
timestamp 1300117811
transform -1 0 6450 0 -1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_831
timestamp 1300117811
transform -1 0 6450 0 -1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_832
timestamp 1300117811
transform -1 0 6450 0 -1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_833
timestamp 1300117811
transform -1 0 6450 0 -1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_834
timestamp 1300117811
transform -1 0 6450 0 -1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_835
timestamp 1300117811
transform -1 0 6450 0 -1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_836
timestamp 1300117811
transform -1 0 6450 0 -1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_837
timestamp 1300117811
transform -1 0 6450 0 -1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_838
timestamp 1300117811
transform -1 0 6450 0 -1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_839
timestamp 1300117811
transform -1 0 6450 0 -1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_840
timestamp 1300117811
transform -1 0 6450 0 -1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_841
timestamp 1300117811
transform -1 0 6450 0 -1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_842
timestamp 1300117811
transform -1 0 6450 0 -1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_843
timestamp 1300117811
transform -1 0 6450 0 -1 22532
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 6450 0 -1 22446
box 0 0 6450 1720
use fillpp_mt fillpp_mt_844
timestamp 1300117811
transform -1 0 6450 0 -1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_845
timestamp 1300117811
transform -1 0 6450 0 -1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_846
timestamp 1300117811
transform -1 0 6450 0 -1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_847
timestamp 1300117811
transform -1 0 6450 0 -1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_848
timestamp 1300117811
transform -1 0 6450 0 -1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_849
timestamp 1300117811
transform -1 0 6450 0 -1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_850
timestamp 1300117811
transform -1 0 6450 0 -1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_851
timestamp 1300117811
transform -1 0 6450 0 -1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_852
timestamp 1300117811
transform -1 0 6450 0 -1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_853
timestamp 1300117811
transform -1 0 6450 0 -1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_854
timestamp 1300117811
transform -1 0 6450 0 -1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_855
timestamp 1300117811
transform -1 0 6450 0 -1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_856
timestamp 1300117811
transform -1 0 6450 0 -1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_857
timestamp 1300117811
transform -1 0 6450 0 -1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_858
timestamp 1300117811
transform -1 0 6450 0 -1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_859
timestamp 1300117811
transform -1 0 6450 0 -1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_860
timestamp 1300117811
transform -1 0 6450 0 -1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_861
timestamp 1300117811
transform -1 0 6450 0 -1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_862
timestamp 1300117811
transform -1 0 6450 0 -1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_863
timestamp 1300117811
transform -1 0 6450 0 -1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_864
timestamp 1300117811
transform -1 0 6450 0 -1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_865
timestamp 1300117811
transform -1 0 6450 0 -1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_866
timestamp 1300117811
transform -1 0 6450 0 -1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_867
timestamp 1300117811
transform -1 0 6450 0 -1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_868
timestamp 1300117811
transform -1 0 6450 0 -1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_869
timestamp 1300117811
transform -1 0 6450 0 -1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_870
timestamp 1300117811
transform -1 0 6450 0 -1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_871
timestamp 1300117811
transform -1 0 6450 0 -1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_872
timestamp 1300117811
transform -1 0 6450 0 -1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_873
timestamp 1300117811
transform -1 0 6450 0 -1 18232
box 0 0 6450 86
use datapath datapath_0
timestamp 1395340701
transform 1 0 11284 0 1 18158
box 414 43 25445 20615
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 1 0 41538 0 1 38700
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 1 0 41538 0 1 38614
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 1 0 41538 0 1 38528
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 1 0 41538 0 1 38442
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 1 0 41538 0 1 38356
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 1 0 41538 0 1 38270
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 1 0 41538 0 1 38184
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 1 0 41538 0 1 38098
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 1 0 41538 0 1 38012
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 1 0 41538 0 1 37926
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 1 0 41538 0 1 37840
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 1 0 41538 0 1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 1 0 41538 0 1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 1 0 41538 0 1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 1 0 41538 0 1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 1 0 41538 0 1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 1 0 41538 0 1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 1 0 41538 0 1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 1 0 41538 0 1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 1 0 41538 0 1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 1 0 41538 0 1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 1 0 41538 0 1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 1 0 41538 0 1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 1 0 41538 0 1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 1 0 41538 0 1 36636
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 41538 0 1 34916
box 0 0 6450 1720
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 1 0 41538 0 1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 1 0 41538 0 1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 1 0 41538 0 1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 1 0 41538 0 1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 1 0 41538 0 1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 1 0 41538 0 1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 1 0 41538 0 1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 1 0 41538 0 1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 1 0 41538 0 1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 1 0 41538 0 1 34056
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 1 0 41538 0 1 33970
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 1 0 41538 0 1 33884
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 1 0 41538 0 1 33798
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 1 0 41538 0 1 33712
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 1 0 41538 0 1 33626
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 1 0 41538 0 1 33540
box 0 0 6450 86
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 1 0 41538 0 1 33454
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 1 0 41538 0 1 33368
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 1 0 41538 0 1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 1 0 41538 0 1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 1 0 41538 0 1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 1 0 41538 0 1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 1 0 41538 0 1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 1 0 41538 0 1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 1 0 41538 0 1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 1 0 41538 0 1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 1 0 41538 0 1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 1 0 41538 0 1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 1 0 41538 0 1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 1 0 41538 0 1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 1 0 41538 0 1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 1 0 41538 0 1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 1 0 41538 0 1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 1 0 41538 0 1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 1 0 41538 0 1 31906
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 41538 0 1 30186
box 0 0 6450 1720
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 1 0 41538 0 1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 1 0 41538 0 1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 1 0 41538 0 1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 1 0 41538 0 1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 1 0 41538 0 1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 1 0 41538 0 1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 1 0 41538 0 1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 1 0 41538 0 1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 1 0 41538 0 1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 1 0 41538 0 1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 41538 0 1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 41538 0 1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 41538 0 1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 41538 0 1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 41538 0 1 28896
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 41538 0 1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 41538 0 1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 41538 0 1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 41538 0 1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 41538 0 1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 41538 0 1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 41538 0 1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 41538 0 1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 41538 0 1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 41538 0 1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 41538 0 1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 41538 0 1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 41538 0 1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 41538 0 1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 41538 0 1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 41538 0 1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 41538 0 1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 41538 0 1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 41538 0 1 27262
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 41538 0 1 27176
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 41538 0 1 25456
box 0 0 6450 1720
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 41538 0 1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 41538 0 1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 41538 0 1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 41538 0 1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 41538 0 1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 41538 0 1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 41538 0 1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 41538 0 1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 41538 0 1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 41538 0 1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 41538 0 1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 41538 0 1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 41538 0 1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 41538 0 1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 41538 0 1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 41538 0 1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 41538 0 1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 41538 0 1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 41538 0 1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 41538 0 1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 41538 0 1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 41538 0 1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 41538 0 1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 41538 0 1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 41538 0 1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 41538 0 1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 41538 0 1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 41538 0 1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 41538 0 1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 41538 0 1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 41538 0 1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 41538 0 1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 41538 0 1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 41538 0 1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 41538 0 1 22446
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 41538 0 1 20726
box 0 0 6450 1720
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 41538 0 1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 41538 0 1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 41538 0 1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 41538 0 1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 41538 0 1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 41538 0 1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 41538 0 1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 41538 0 1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 41538 0 1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 41538 0 1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 41538 0 1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 41538 0 1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 41538 0 1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 41538 0 1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 41538 0 1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 41538 0 1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 41538 0 1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 41538 0 1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 41538 0 1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 41538 0 1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 41538 0 1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 41538 0 1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 41538 0 1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 41538 0 1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 41538 0 1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 41538 0 1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 41538 0 1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 41538 0 1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 41538 0 1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_874
timestamp 1300117811
transform -1 0 6450 0 -1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_875
timestamp 1300117811
transform -1 0 6450 0 -1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_876
timestamp 1300117811
transform -1 0 6450 0 -1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_877
timestamp 1300117811
transform -1 0 6450 0 -1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_878
timestamp 1300117811
transform -1 0 6450 0 -1 17802
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 6450 0 -1 17716
box 0 0 6450 1720
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 41538 0 1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 41538 0 1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 41538 0 1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 41538 0 1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 41538 0 1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 41538 0 1 17716
box 0 0 6450 86
use fillpp_mt fillpp_mt_879
timestamp 1300117811
transform -1 0 6450 0 -1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_880
timestamp 1300117811
transform -1 0 6450 0 -1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_881
timestamp 1300117811
transform -1 0 6450 0 -1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_882
timestamp 1300117811
transform -1 0 6450 0 -1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_883
timestamp 1300117811
transform -1 0 6450 0 -1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_884
timestamp 1300117811
transform -1 0 6450 0 -1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_885
timestamp 1300117811
transform -1 0 6450 0 -1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_886
timestamp 1300117811
transform -1 0 6450 0 -1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_887
timestamp 1300117811
transform -1 0 6450 0 -1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_888
timestamp 1300117811
transform -1 0 6450 0 -1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_889
timestamp 1300117811
transform -1 0 6450 0 -1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_890
timestamp 1300117811
transform -1 0 6450 0 -1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_891
timestamp 1300117811
transform -1 0 6450 0 -1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_892
timestamp 1300117811
transform -1 0 6450 0 -1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_893
timestamp 1300117811
transform -1 0 6450 0 -1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_894
timestamp 1300117811
transform -1 0 6450 0 -1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_895
timestamp 1300117811
transform -1 0 6450 0 -1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_896
timestamp 1300117811
transform -1 0 6450 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_897
timestamp 1300117811
transform -1 0 6450 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_898
timestamp 1300117811
transform -1 0 6450 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_899
timestamp 1300117811
transform -1 0 6450 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_900
timestamp 1300117811
transform -1 0 6450 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_901
timestamp 1300117811
transform -1 0 6450 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_902
timestamp 1300117811
transform -1 0 6450 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_903
timestamp 1300117811
transform -1 0 6450 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_904
timestamp 1300117811
transform -1 0 6450 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_905
timestamp 1300117811
transform -1 0 6450 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_906
timestamp 1300117811
transform -1 0 6450 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_907
timestamp 1300117811
transform -1 0 6450 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_908
timestamp 1300117811
transform -1 0 6450 0 -1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_909
timestamp 1300117811
transform -1 0 6450 0 -1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_910
timestamp 1300117811
transform -1 0 6450 0 -1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_911
timestamp 1300117811
transform -1 0 6450 0 -1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_912
timestamp 1300117811
transform -1 0 6450 0 -1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_913
timestamp 1300117811
transform -1 0 6450 0 -1 13072
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 6450 0 -1 12986
box 0 0 6450 1720
use fillpp_mt fillpp_mt_914
timestamp 1300117811
transform -1 0 6450 0 -1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_915
timestamp 1300117811
transform -1 0 6450 0 -1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_916
timestamp 1300117811
transform -1 0 6450 0 -1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_917
timestamp 1300117811
transform -1 0 6450 0 -1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_918
timestamp 1300117811
transform -1 0 6450 0 -1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_919
timestamp 1300117811
transform -1 0 6450 0 -1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_920
timestamp 1300117811
transform -1 0 6450 0 -1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_921
timestamp 1300117811
transform -1 0 6450 0 -1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_922
timestamp 1300117811
transform -1 0 6450 0 -1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_923
timestamp 1300117811
transform -1 0 6450 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_924
timestamp 1300117811
transform -1 0 6450 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_925
timestamp 1300117811
transform -1 0 6450 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_926
timestamp 1300117811
transform -1 0 6450 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_927
timestamp 1300117811
transform -1 0 6450 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_928
timestamp 1300117811
transform -1 0 6450 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_929
timestamp 1300117811
transform -1 0 6450 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_930
timestamp 1300117811
transform -1 0 6450 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_931
timestamp 1300117811
transform -1 0 6450 0 -1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_932
timestamp 1300117811
transform -1 0 6450 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_933
timestamp 1300117811
transform -1 0 6450 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_934
timestamp 1300117811
transform -1 0 6450 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_935
timestamp 1300117811
transform -1 0 6450 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_936
timestamp 1300117811
transform -1 0 6450 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_937
timestamp 1300117811
transform -1 0 6450 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_938
timestamp 1300117811
transform -1 0 6450 0 -1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_939
timestamp 1300117811
transform -1 0 6450 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_940
timestamp 1300117811
transform -1 0 6450 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_941
timestamp 1300117811
transform -1 0 6450 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_942
timestamp 1300117811
transform -1 0 6450 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_943
timestamp 1300117811
transform -1 0 6450 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_944
timestamp 1300117811
transform -1 0 6450 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_945
timestamp 1300117811
transform -1 0 6450 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_946
timestamp 1300117811
transform -1 0 6450 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_947
timestamp 1300117811
transform -1 0 6450 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_948
timestamp 1300117811
transform -1 0 6450 0 -1 8342
box 0 0 6450 86
use control control_0
timestamp 1395431750
transform 1 0 9960 0 1 8334
box 0 0 27649 8170
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 41538 0 1 15996
box 0 0 6450 1720
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 41538 0 1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 41538 0 1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 41538 0 1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 41538 0 1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 41538 0 1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 41538 0 1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 41538 0 1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 41538 0 1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 41538 0 1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 41538 0 1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 41538 0 1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 41538 0 1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 41538 0 1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 41538 0 1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 41538 0 1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 41538 0 1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 41538 0 1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 41538 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 41538 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 41538 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 41538 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 41538 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 41538 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 41538 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 41538 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 41538 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 41538 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 41538 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 41538 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 41538 0 1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 41538 0 1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 41538 0 1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 41538 0 1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 41538 0 1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 41538 0 1 12986
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 41538 0 1 11266
box 0 0 6450 1720
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 41538 0 1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 41538 0 1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 41538 0 1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 41538 0 1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 41538 0 1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 41538 0 1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 41538 0 1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 41538 0 1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 41538 0 1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 41538 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 41538 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 41538 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 41538 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 41538 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 41538 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 41538 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 41538 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 41538 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 41538 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 41538 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 41538 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 41538 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 41538 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 41538 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 41538 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 41538 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 41538 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 41538 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 41538 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 41538 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 41538 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 41538 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 41538 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 41538 0 1 8342
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 6450 0 -1 8256
box 0 0 6450 1720
use fillpp_mt fillpp_mt_949
timestamp 1300117811
transform -1 0 6450 0 -1 6536
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 41538 0 1 8256
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 41538 0 1 6536
box 0 0 6450 1720
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 41538 0 1 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 0 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 6450 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 6536 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6622 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 8342 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 8428 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 8514 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 8600 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8686 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8772 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8858 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8944 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 9030 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 9116 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 9202 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 9288 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 9374 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 9460 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 9546 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9632 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9718 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9804 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9890 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9976 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 10062 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 10148 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 10234 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 10320 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 10406 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 10492 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 10578 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 10664 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10750 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 12470 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 12556 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 12642 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 12728 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 12814 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12900 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12986 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 13072 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 13158 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 13244 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 13330 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 13416 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 13502 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 13588 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 13674 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 13760 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 13846 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 13932 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 14018 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 14104 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 14190 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 14276 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 14362 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 14448 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 14534 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 14620 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 14706 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 14792 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 14878 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 16598 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 16684 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 16770 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 16856 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 16942 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 17028 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 17114 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 17200 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 17286 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 17372 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 17458 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 17544 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 17630 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 17716 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 17802 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 17888 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 17974 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 18060 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 18146 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 18232 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 18318 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 18404 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 18490 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 18576 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 18662 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 18748 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 18834 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 18920 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 19006 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 20726 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 20812 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 20898 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 20984 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 21070 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 21156 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 21242 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 21328 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 21414 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 21500 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 21586 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 21672 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 21758 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 21844 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 21930 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 22016 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 22102 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 22188 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 22274 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 22360 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 22446 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 22532 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 22618 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 22704 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 22790 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 22876 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 22962 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 23048 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 23134 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 24854 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 24940 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 25026 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 25112 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 25198 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 25284 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 25370 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 25456 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 25542 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 25628 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 25714 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 25800 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 25886 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 25972 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 26058 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 26144 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 26230 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 26316 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 26402 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 26488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 26574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 26660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 26746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 26832 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 26918 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 27004 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 27090 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 27176 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 27262 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 28982 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 29068 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 29154 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 29240 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 29326 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 29412 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 29498 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 29584 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 29670 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 29756 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 29842 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 29928 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 30014 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 30100 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 30186 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 30272 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 30358 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 30444 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 30530 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 30616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 30702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 30788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 30874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 30960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 31046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 31132 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 31218 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 31304 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 31390 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 0 1 33110 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 0 1 33196 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 0 1 33282 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 0 1 33368 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 0 1 33454 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 0 1 33540 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 0 1 33626 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 0 1 33712 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 0 1 33798 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 0 1 33884 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 0 1 33970 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 0 1 34056 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 0 1 34142 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 0 1 34228 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 0 1 34314 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 0 1 34400 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 0 1 34486 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 0 1 34572 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 0 1 34658 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 0 1 34744 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 0 1 34830 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 0 1 34916 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 0 1 35002 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 0 1 35088 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 0 1 35174 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 0 1 35260 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 0 1 35346 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 0 1 35432 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 35518 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 0 1 37238 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 0 1 37324 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 0 1 37410 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 0 1 37496 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 0 1 37582 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 0 1 37668 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 0 1 37754 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 0 1 37840 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 0 1 37926 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 0 1 38012 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 0 1 38098 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 0 1 38184 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 0 1 38270 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 0 1 38356 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 0 1 38442 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 0 1 38528 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 0 1 38614 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 0 1 38700 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 0 1 38786 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 0 1 38872 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 0 1 38958 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 0 1 39044 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 0 1 39130 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 0 1 39216 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 0 1 39302 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 0 1 39388 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 0 1 39474 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 0 1 39560 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 39646 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 0 1 41366 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 0 1 41452 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 47988 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 6702 78 8262 1638 0 nIRQ
rlabel metal4 10830 78 12390 1638 0 Data[0]
rlabel metal4 14958 78 16518 1638 0 Data[1]
rlabel metal4 19086 78 20646 1638 0 Data[2]
rlabel metal4 23214 78 24774 1638 0 vdde!
rlabel metal4 27342 78 28902 1638 0 Data[3]
rlabel metal4 31470 78 33030 1638 0 Data[4]
rlabel metal4 35598 78 37158 1638 0 Data[5]
rlabel metal4 39726 78 41286 1638 0 gnde!
rlabel metal4 46350 6616 47910 8176 0 Data[6]
rlabel metal4 46350 11346 47910 12906 0 Data[7]
rlabel metal4 46350 16076 47910 17636 0 Data[8]
rlabel metal4 46350 20806 47910 22366 0 gnde!
rlabel metal4 46350 25536 47910 27096 0 GND!
rlabel metal4 46350 30266 47910 31826 0 Data[9]
rlabel metal4 46350 34996 47910 36556 0 Data[10]
rlabel metal4 46350 39726 47910 41286 0 Data[11]
rlabel metal4 39726 46264 41286 47824 0 vdde!
rlabel metal4 35598 46264 37158 47824 0 Data[12]
rlabel metal4 31470 46264 33030 47824 0 Data[13]
rlabel metal4 27342 46264 28902 47824 0 Data[14]
rlabel metal4 23214 46264 24774 47824 0 gnde!
rlabel metal4 19086 46264 20646 47824 0 Data[15]
rlabel metal4 14958 46264 16518 47824 0 ALE
rlabel metal4 10830 46264 12390 47824 0 nME
rlabel metal4 6702 46264 8262 47824 0 nWait
rlabel metal4 78 39726 1638 41286 0 nOE
rlabel metal4 78 34996 1638 36556 0 RnW
rlabel metal4 78 30266 1638 31826 0 SDO
rlabel metal4 78 25536 1638 27096 0 Vdd!
rlabel metal4 78 20806 1638 22366 0 SDI
rlabel metal4 78 16076 1638 17636 0 Test
rlabel metal4 78 11346 1638 12906 0 Clock
rlabel metal4 78 6616 1638 8176 0 nReset
<< end >>
