magic
tech c035u
timestamp 1395929462
<< metal1 >>
rect 21736 8036 21754 8050
rect 12760 8014 19454 8024
rect 21052 8014 24434 8024
rect 8488 7988 8506 8002
rect 9376 7988 9394 8002
rect 12184 7990 14786 8000
rect 17704 7988 17722 8002
rect 17896 7990 26066 8000
rect 3640 7966 4046 7976
rect 5248 7964 5266 7978
rect 7288 7966 9986 7976
rect 10264 7964 10282 7978
rect 11368 7966 24746 7976
rect 3496 7942 13022 7952
rect 13936 7942 24278 7952
rect 3280 7918 14630 7928
rect 15040 7918 16238 7928
rect 17296 7918 26114 7928
rect 84 7894 1682 7904
rect 2392 7894 5330 7904
rect 6304 7894 23474 7904
rect 26008 7894 26042 7904
rect 84 7870 2234 7880
rect 3016 7870 5678 7880
rect 7288 7870 15434 7880
rect 16360 7870 18650 7880
rect 20896 7870 21866 7880
rect 3208 7846 6794 7856
rect 8008 7844 8026 7858
rect 8440 7846 12206 7856
rect 12256 7846 22670 7856
rect 26104 7846 26437 7856
rect 4024 7822 11402 7832
rect 11632 7822 26018 7832
rect 26080 7822 26437 7832
rect 12208 7798 14090 7808
rect 14104 7798 17138 7808
rect 17152 7798 26090 7808
rect 26128 7798 26437 7808
rect 14620 7774 15146 7784
rect 15280 7774 25082 7784
rect 26056 7774 26437 7784
rect 18640 7750 23618 7760
rect 26032 7750 26437 7760
rect 12136 6917 12338 6927
rect 20488 6917 20498 6927
rect 12112 6893 25778 6903
rect 12064 6869 20474 6879
rect 11704 6845 15386 6855
rect 22288 6845 22298 6855
rect 11440 6821 11834 6831
rect 12040 6821 12254 6831
rect 12544 6821 22802 6831
rect 10816 6797 12914 6807
rect 12928 6797 22274 6807
rect 10576 6773 14450 6783
rect 14464 6773 21482 6783
rect 10408 6749 16034 6759
rect 16048 6749 16370 6759
rect 16384 6749 21938 6759
rect 21952 6749 23474 6759
rect 10360 6725 19298 6735
rect 10120 6701 11690 6711
rect 12016 6701 24650 6711
rect 9424 6677 9530 6687
rect 9688 6677 25490 6687
rect 9184 6653 21674 6663
rect 8968 6629 21530 6639
rect 8920 6605 8954 6615
rect 9160 6605 20402 6615
rect 8848 6581 16082 6591
rect 8824 6557 13946 6567
rect 8560 6533 11066 6543
rect 11080 6533 11234 6543
rect 11248 6533 16154 6543
rect 16168 6533 21026 6543
rect 21040 6533 22706 6543
rect 8560 6509 17906 6519
rect 8488 6485 15578 6495
rect 8488 6461 17690 6471
rect 8344 6437 11810 6447
rect 11920 6437 12170 6447
rect 12496 6437 16538 6447
rect 17416 6437 24746 6447
rect 8176 6413 8234 6423
rect 8320 6413 10058 6423
rect 10072 6413 22058 6423
rect 7936 6389 24074 6399
rect 7912 6365 10970 6375
rect 11296 6365 11330 6375
rect 11392 6365 20834 6375
rect 7888 6341 22490 6351
rect 7840 6317 25538 6327
rect 7456 6293 8618 6303
rect 8632 6293 8930 6303
rect 8944 6293 22586 6303
rect 7408 6269 21122 6279
rect 7288 6245 7970 6255
rect 8056 6245 19418 6255
rect 7240 6221 10778 6231
rect 10864 6221 11450 6231
rect 11656 6221 20066 6231
rect 7240 6197 19226 6207
rect 7192 6173 23930 6183
rect 7144 6149 11954 6159
rect 11968 6149 14834 6159
rect 14848 6149 25562 6159
rect 6880 6125 9482 6135
rect 9496 6125 12362 6135
rect 12376 6125 13826 6135
rect 16624 6125 16634 6135
rect 17344 6125 18938 6135
rect 22984 6125 23066 6135
rect 6832 6101 22970 6111
rect 6736 6077 22106 6087
rect 6712 6053 6722 6063
rect 6808 6053 6842 6063
rect 6904 6053 17738 6063
rect 17752 6053 25514 6063
rect 25624 6053 25826 6063
rect 6688 6029 8018 6039
rect 8080 6029 13322 6039
rect 16072 6029 16346 6039
rect 16576 6029 23282 6039
rect 23296 6029 25610 6039
rect 6472 6005 15218 6015
rect 15232 6005 21626 6015
rect 21640 6005 23306 6015
rect 6376 5981 7394 5991
rect 7408 5981 7682 5991
rect 7696 5981 8666 5991
rect 8680 5981 12002 5991
rect 12016 5981 24938 5991
rect 24952 5981 25802 5991
rect 6328 5957 6962 5967
rect 7024 5957 19778 5967
rect 6160 5933 14114 5943
rect 15208 5933 17882 5943
rect 6064 5909 7322 5919
rect 7336 5909 8858 5919
rect 8872 5909 10946 5919
rect 10960 5909 16202 5919
rect 16216 5909 18554 5919
rect 18568 5909 21074 5919
rect 6016 5885 16442 5895
rect 16504 5885 24938 5895
rect 5968 5861 9002 5871
rect 9064 5861 9170 5871
rect 9328 5861 25634 5871
rect 5968 5837 7034 5847
rect 7096 5837 10562 5847
rect 10576 5837 23402 5847
rect 25360 5837 25418 5847
rect 5800 5813 8594 5823
rect 8800 5813 19034 5823
rect 25312 5813 25322 5823
rect 25768 5813 25874 5823
rect 5800 5789 12578 5799
rect 12664 5789 13562 5799
rect 13576 5789 15986 5799
rect 16000 5789 21290 5799
rect 21304 5789 24026 5799
rect 24040 5789 24506 5799
rect 24520 5789 25730 5799
rect 5704 5765 15194 5775
rect 16024 5765 25754 5775
rect 5680 5741 5690 5751
rect 5776 5741 6530 5751
rect 6592 5741 7034 5751
rect 7048 5741 8066 5751
rect 8080 5741 11618 5751
rect 11632 5741 16178 5751
rect 16192 5741 18074 5751
rect 18088 5741 18854 5751
rect 18868 5741 19178 5751
rect 19192 5741 20690 5751
rect 20704 5741 25346 5751
rect 5656 5717 19046 5727
rect 19060 5717 25298 5727
rect 5656 5693 15482 5703
rect 15712 5693 25418 5703
rect 5608 5669 8282 5679
rect 8296 5669 10154 5679
rect 10216 5669 23978 5679
rect 5608 5645 6170 5655
rect 6232 5645 16730 5655
rect 17296 5645 17546 5655
rect 5584 5621 13874 5631
rect 15688 5621 24986 5631
rect 5584 5597 25994 5607
rect 5560 5573 6290 5583
rect 6304 5573 6362 5583
rect 6424 5573 10682 5583
rect 10768 5573 21950 5583
rect 5464 5549 16106 5559
rect 16480 5549 23378 5559
rect 5440 5525 6074 5535
rect 6088 5525 18122 5535
rect 5392 5501 11354 5511
rect 11368 5501 18410 5511
rect 18424 5501 25442 5511
rect 5320 5477 11522 5487
rect 11536 5477 18986 5487
rect 19000 5477 21986 5487
rect 5272 5453 16274 5463
rect 16336 5453 20066 5463
rect 5272 5429 9746 5439
rect 10120 5429 19682 5439
rect 5248 5405 7466 5415
rect 7480 5405 9074 5415
rect 9088 5405 10322 5415
rect 10336 5405 12074 5415
rect 12088 5405 14666 5415
rect 14680 5405 17402 5415
rect 17416 5405 20594 5415
rect 20608 5405 21842 5415
rect 21856 5405 25370 5415
rect 5152 5381 7754 5391
rect 7768 5381 21746 5391
rect 4984 5357 6866 5367
rect 6880 5357 10610 5367
rect 10624 5357 18290 5367
rect 4912 5333 12698 5343
rect 13288 5333 19994 5343
rect 4864 5309 11762 5319
rect 11872 5309 22826 5319
rect 4816 5285 7346 5295
rect 7360 5285 13370 5295
rect 13384 5285 20138 5295
rect 4792 5261 11882 5271
rect 11992 5261 20618 5271
rect 4672 5237 8330 5247
rect 8344 5237 11666 5247
rect 11752 5237 14618 5247
rect 15544 5237 23786 5247
rect 4624 5213 7826 5223
rect 7840 5213 18626 5223
rect 18640 5213 24554 5223
rect 4600 5189 9218 5199
rect 9232 5189 12674 5199
rect 13264 5189 13442 5199
rect 13528 5189 13586 5199
rect 14656 5189 14714 5199
rect 15328 5189 15506 5199
rect 15568 5189 15770 5199
rect 15928 5189 19274 5199
rect 4552 5165 25706 5175
rect 4360 5141 4658 5151
rect 4672 5141 9002 5151
rect 9016 5141 9674 5151
rect 9688 5141 11138 5151
rect 11152 5141 22106 5151
rect 22120 5141 23882 5151
rect 4336 5117 23738 5127
rect 4312 5093 13706 5103
rect 13936 5093 21458 5103
rect 21472 5093 21698 5103
rect 4264 5069 23018 5079
rect 4240 5045 9410 5055
rect 9640 5045 18266 5055
rect 18280 5045 22874 5055
rect 4144 5021 25850 5031
rect 4096 4997 13298 5007
rect 13408 4997 15410 5007
rect 15472 4997 20858 5007
rect 20872 4997 23474 5007
rect 4096 4973 17642 4983
rect 23368 4973 23438 4983
rect 4072 4949 13106 4959
rect 13216 4949 23570 4959
rect 4000 4925 7010 4935
rect 7024 4925 11186 4935
rect 11200 4925 12218 4935
rect 12232 4925 13226 4935
rect 13240 4925 14594 4935
rect 14608 4925 15434 4935
rect 15448 4925 18194 4935
rect 18208 4925 19922 4935
rect 19936 4925 23114 4935
rect 23128 4925 23234 4935
rect 23248 4925 23354 4935
rect 23368 4925 23834 4935
rect 3904 4901 18242 4911
rect 19984 4901 20306 4911
rect 3880 4877 7562 4887
rect 7576 4877 19970 4887
rect 3832 4853 17618 4863
rect 17632 4853 23762 4863
rect 3808 4829 7586 4839
rect 7600 4829 7706 4839
rect 7720 4829 9938 4839
rect 9952 4829 14282 4839
rect 14296 4829 18218 4839
rect 18232 4829 19538 4839
rect 19552 4829 23162 4839
rect 23176 4829 24146 4839
rect 3784 4805 7106 4815
rect 7120 4805 9242 4815
rect 9256 4805 9554 4815
rect 9568 4805 15890 4815
rect 15904 4805 17378 4815
rect 17392 4805 20570 4815
rect 3736 4781 4106 4791
rect 4168 4781 4466 4791
rect 4552 4781 16298 4791
rect 16432 4781 18746 4791
rect 22696 4781 22922 4791
rect 3712 4757 4226 4767
rect 4240 4757 6818 4767
rect 6832 4757 7970 4767
rect 7984 4757 7994 4767
rect 8008 4757 8090 4767
rect 8104 4757 9506 4767
rect 9520 4757 16130 4767
rect 16144 4757 19010 4767
rect 19024 4757 20258 4767
rect 20272 4757 22682 4767
rect 22696 4757 24098 4767
rect 3688 4733 4850 4743
rect 4864 4733 7514 4743
rect 7528 4733 7778 4743
rect 7792 4733 16106 4743
rect 16120 4733 23498 4743
rect 3664 4709 9698 4719
rect 9712 4709 12818 4719
rect 12832 4709 13850 4719
rect 13864 4709 22202 4719
rect 22216 4709 23042 4719
rect 3592 4685 22442 4695
rect 3544 4661 10922 4671
rect 10936 4661 14474 4671
rect 14488 4661 17354 4671
rect 17368 4661 18410 4671
rect 3544 4637 8210 4647
rect 8272 4637 10178 4647
rect 10192 4637 21506 4647
rect 3400 4613 14234 4623
rect 14392 4613 25082 4623
rect 3376 4589 12146 4599
rect 12448 4589 17810 4599
rect 20056 4589 25322 4599
rect 3352 4565 14498 4575
rect 14608 4565 14618 4575
rect 14896 4565 20042 4575
rect 22336 4565 22418 4575
rect 3232 4541 3458 4551
rect 3472 4541 7250 4551
rect 7264 4541 15122 4551
rect 15136 4541 18602 4551
rect 20248 4541 24338 4551
rect 3184 4517 5738 4527
rect 5752 4517 14042 4527
rect 14056 4517 19730 4527
rect 19744 4517 22322 4527
rect 23152 4517 23798 4527
rect 3136 4493 3266 4503
rect 3280 4493 8762 4503
rect 8776 4493 10082 4503
rect 10096 4493 13010 4503
rect 13024 4493 16418 4503
rect 16432 4493 21890 4503
rect 21904 4493 22658 4503
rect 22672 4493 25466 4503
rect 3112 4469 21578 4479
rect 21592 4469 21818 4479
rect 21832 4469 23138 4479
rect 3064 4445 12122 4455
rect 12328 4445 15938 4455
rect 15952 4445 17738 4455
rect 17800 4445 17822 4455
rect 20128 4445 20498 4455
rect 21208 4445 24482 4455
rect 3016 4421 5810 4431
rect 5824 4421 6578 4431
rect 6592 4421 8906 4431
rect 8920 4421 12026 4431
rect 12040 4421 17306 4431
rect 17320 4421 17786 4431
rect 18712 4421 18950 4431
rect 19096 4421 19154 4431
rect 19840 4421 19898 4431
rect 20104 4421 22370 4431
rect 2992 4397 6386 4407
rect 6400 4397 18722 4407
rect 18904 4397 22922 4407
rect 2968 4373 8402 4383
rect 8464 4373 8954 4383
rect 8968 4373 9842 4383
rect 10024 4373 17570 4383
rect 18184 4373 18302 4383
rect 18496 4373 22778 4383
rect 22912 4373 22922 4383
rect 2944 4349 21554 4359
rect 21808 4349 22178 4359
rect 22192 4349 22634 4359
rect 22648 4349 24266 4359
rect 24640 4349 24722 4359
rect 25720 4349 25874 4359
rect 2920 4325 4994 4335
rect 5008 4325 5186 4335
rect 5200 4325 8258 4335
rect 8272 4325 13034 4335
rect 13048 4325 15818 4335
rect 15832 4325 18506 4335
rect 18616 4325 25202 4335
rect 2896 4301 4418 4311
rect 4432 4301 5666 4311
rect 5680 4301 8282 4311
rect 8296 4301 20354 4311
rect 20368 4301 21770 4311
rect 21784 4301 22538 4311
rect 22624 4301 26437 4311
rect 2872 4277 7610 4287
rect 7624 4277 10202 4287
rect 10216 4277 11162 4287
rect 11176 4277 11282 4287
rect 11296 4277 18122 4287
rect 18136 4277 24650 4287
rect 2800 4253 4970 4263
rect 5032 4253 11714 4263
rect 11800 4253 12866 4263
rect 12880 4253 21146 4263
rect 21784 4253 21842 4263
rect 21904 4253 21950 4263
rect 22456 4253 22706 4263
rect 2728 4229 21866 4239
rect 2680 4205 7130 4215
rect 7144 4205 11090 4215
rect 11104 4205 16442 4215
rect 16456 4205 23330 4215
rect 2656 4181 8570 4191
rect 8656 4181 18338 4191
rect 18352 4181 22250 4191
rect 22264 4181 24362 4191
rect 2608 4157 11090 4167
rect 11320 4157 11426 4167
rect 11584 4157 13994 4167
rect 14008 4157 19370 4167
rect 20776 4157 23666 4167
rect 2536 4133 3962 4143
rect 3976 4133 6626 4143
rect 6640 4133 8162 4143
rect 8176 4133 10226 4143
rect 10240 4133 13154 4143
rect 13168 4133 15842 4143
rect 15856 4133 19826 4143
rect 19840 4133 21266 4143
rect 21280 4133 21602 4143
rect 2464 4109 7442 4119
rect 7456 4109 8882 4119
rect 8896 4109 13514 4119
rect 13528 4109 18530 4119
rect 18544 4109 23210 4119
rect 2416 4085 13106 4095
rect 13120 4085 20714 4095
rect 20824 4085 21722 4095
rect 2344 4061 5210 4071
rect 5224 4061 7946 4071
rect 7960 4061 9122 4071
rect 9136 4061 14858 4071
rect 14872 4061 17690 4071
rect 17704 4061 20450 4071
rect 21088 4061 23066 4071
rect 2296 4037 7202 4047
rect 7216 4037 12050 4047
rect 12064 4037 15650 4047
rect 16024 4037 23618 4047
rect 2200 4013 22154 4023
rect 2176 3989 18818 3999
rect 19024 3989 19046 3999
rect 21280 3989 21290 3999
rect 2104 3965 10418 3975
rect 10432 3965 12794 3975
rect 12808 3965 25154 3975
rect 2056 3941 6794 3951
rect 6808 3941 7730 3951
rect 7744 3941 10994 3951
rect 11368 3941 16466 3951
rect 16480 3941 21242 3951
rect 21256 3941 21386 3951
rect 1984 3917 2186 3927
rect 2200 3917 4370 3927
rect 4384 3917 8738 3927
rect 8752 3917 10826 3927
rect 10840 3917 11018 3927
rect 11032 3917 13178 3927
rect 13192 3917 17618 3927
rect 17632 3917 18362 3927
rect 18376 3917 19802 3927
rect 19816 3917 20666 3927
rect 1960 3893 9458 3903
rect 9472 3893 11546 3903
rect 11560 3893 12194 3903
rect 12208 3893 22586 3903
rect 22600 3893 23234 3903
rect 1912 3869 5066 3879
rect 5080 3869 12722 3879
rect 12736 3869 20786 3879
rect 1888 3845 3938 3855
rect 3952 3845 6554 3855
rect 6568 3845 9434 3855
rect 9448 3845 9866 3855
rect 9880 3845 11042 3855
rect 11056 3845 13538 3855
rect 13552 3845 18578 3855
rect 18592 3845 23714 3855
rect 1864 3821 2738 3831
rect 2752 3821 16226 3831
rect 16240 3821 22346 3831
rect 1816 3797 5858 3807
rect 5920 3797 22538 3807
rect 1768 3773 7802 3783
rect 7816 3773 9314 3783
rect 9376 3773 21206 3783
rect 1720 3749 20282 3759
rect 1648 3725 1730 3735
rect 1744 3725 2210 3735
rect 2224 3725 2234 3735
rect 2248 3725 3338 3735
rect 3352 3725 4754 3735
rect 4768 3725 5090 3735
rect 5104 3725 9050 3735
rect 9064 3725 14570 3735
rect 14584 3725 15218 3735
rect 15232 3725 16226 3735
rect 16240 3725 20162 3735
rect 20176 3725 23858 3735
rect 23872 3725 25922 3735
rect 1624 3701 21914 3711
rect 21928 3701 22394 3711
rect 84 3677 2378 3687
rect 2392 3677 7370 3687
rect 7384 3677 13082 3687
rect 13096 3677 23906 3687
rect 84 3653 13418 3663
rect 13672 3653 17474 3663
rect 18472 3653 19130 3663
rect 19144 3653 20210 3663
rect 23920 3653 24146 3663
rect 2008 3629 18698 3639
rect 2512 3605 4586 3615
rect 4600 3605 4730 3615
rect 4744 3605 5474 3615
rect 5488 3605 5978 3615
rect 5992 3605 15314 3615
rect 15328 3605 18338 3615
rect 18592 3605 18626 3615
rect 18736 3605 18854 3615
rect 2536 3581 9650 3591
rect 9664 3581 9962 3591
rect 9976 3581 14258 3591
rect 14272 3581 14642 3591
rect 14656 3581 18050 3591
rect 18064 3581 19850 3591
rect 19864 3581 24626 3591
rect 2560 3557 19082 3567
rect 2608 3533 4706 3543
rect 4720 3533 5330 3543
rect 5344 3533 6770 3543
rect 6784 3533 14738 3543
rect 14752 3533 22010 3543
rect 2632 3509 4298 3519
rect 4312 3509 4754 3519
rect 4768 3509 6842 3519
rect 6856 3509 11474 3519
rect 11488 3509 14762 3519
rect 14920 3509 25682 3519
rect 2704 3485 15434 3495
rect 15496 3485 15578 3495
rect 16096 3485 16370 3495
rect 16528 3485 24410 3495
rect 2800 3461 18170 3471
rect 18184 3461 18914 3471
rect 2824 3437 6506 3447
rect 6520 3437 24218 3447
rect 2848 3413 13346 3423
rect 13360 3413 16298 3423
rect 17440 3413 18674 3423
rect 18688 3413 19946 3423
rect 2896 3389 14978 3399
rect 14992 3389 22898 3399
rect 22912 3389 23690 3399
rect 23704 3389 24842 3399
rect 2920 3365 3362 3375
rect 3376 3365 11210 3375
rect 11224 3365 13058 3375
rect 13072 3365 15338 3375
rect 16264 3365 16394 3375
rect 2944 3341 4250 3351
rect 4264 3341 5114 3351
rect 5128 3341 5234 3351
rect 5248 3341 8810 3351
rect 8824 3341 9986 3351
rect 10000 3341 15362 3351
rect 15376 3341 15746 3351
rect 15760 3341 17954 3351
rect 17968 3341 20546 3351
rect 20560 3341 21410 3351
rect 21424 3341 24122 3351
rect 3016 3317 3626 3327
rect 3640 3317 5474 3327
rect 5488 3317 5690 3327
rect 5704 3317 7250 3327
rect 7264 3317 7922 3327
rect 7936 3317 11330 3327
rect 11344 3317 12938 3327
rect 12952 3317 16058 3327
rect 16072 3317 17978 3327
rect 17992 3317 18002 3327
rect 18016 3317 19106 3327
rect 19120 3317 24962 3327
rect 3040 3293 3218 3303
rect 3232 3293 11402 3303
rect 11416 3293 13250 3303
rect 13264 3293 18434 3303
rect 18448 3293 22154 3303
rect 22168 3293 22994 3303
rect 3064 3269 15506 3279
rect 15520 3269 23642 3279
rect 3112 3245 4514 3255
rect 4528 3245 6674 3255
rect 6688 3245 19874 3255
rect 3136 3221 6938 3231
rect 6952 3221 14882 3231
rect 14896 3221 19634 3231
rect 19648 3221 21818 3231
rect 3184 3197 9146 3207
rect 9160 3197 22730 3207
rect 3400 3173 10298 3183
rect 10312 3173 15794 3183
rect 15808 3173 18146 3183
rect 18160 3173 19154 3183
rect 19168 3173 20234 3183
rect 20248 3173 24674 3183
rect 3424 3149 14954 3159
rect 14968 3149 18218 3159
rect 3448 3125 9506 3135
rect 9736 3125 14402 3135
rect 14560 3125 15722 3135
rect 15736 3125 17654 3135
rect 17668 3125 20186 3135
rect 20200 3125 21314 3135
rect 3568 3101 18842 3111
rect 3904 3077 6698 3087
rect 6712 3077 9266 3087
rect 9280 3077 10730 3087
rect 10744 3077 10802 3087
rect 10816 3077 11906 3087
rect 11920 3077 12458 3087
rect 12472 3077 13634 3087
rect 13648 3077 17282 3087
rect 17296 3077 18098 3087
rect 18112 3077 19034 3087
rect 19048 3077 21362 3087
rect 3928 3053 8138 3063
rect 8200 3053 9890 3063
rect 9976 3053 17522 3063
rect 21376 3053 21746 3063
rect 4024 3029 5018 3039
rect 5152 3029 17498 3039
rect 4216 3005 15362 3015
rect 15760 3005 15818 3015
rect 17536 3005 17882 3015
rect 4288 2981 6746 2991
rect 6928 2981 8378 2991
rect 8392 2981 15098 2991
rect 15304 2981 19202 2991
rect 19216 2981 20906 2991
rect 20920 2981 22298 2991
rect 22312 2981 22658 2991
rect 4504 2957 25562 2967
rect 4624 2933 7418 2943
rect 7432 2933 9530 2943
rect 9544 2933 10538 2943
rect 10552 2933 10874 2943
rect 10888 2933 11306 2943
rect 11320 2933 15554 2943
rect 15568 2933 17762 2943
rect 17776 2933 21650 2943
rect 21664 2933 22130 2943
rect 22144 2933 22466 2943
rect 22480 2933 24482 2943
rect 4648 2909 21410 2919
rect 22144 2909 22178 2919
rect 4696 2885 26437 2895
rect 4744 2861 20882 2871
rect 20896 2861 25274 2871
rect 4840 2837 7562 2847
rect 7576 2837 10442 2847
rect 10456 2837 11810 2847
rect 11824 2837 22922 2847
rect 22936 2837 23522 2847
rect 4888 2813 6482 2823
rect 6496 2813 13202 2823
rect 13216 2813 14810 2823
rect 14824 2813 20378 2823
rect 20392 2813 22226 2823
rect 22240 2813 24002 2823
rect 24016 2813 25130 2823
rect 5008 2789 25946 2799
rect 5200 2765 14690 2775
rect 14704 2765 18650 2775
rect 18664 2765 20306 2775
rect 20320 2765 23438 2775
rect 23452 2765 25034 2775
rect 5320 2741 9098 2751
rect 9112 2741 17594 2751
rect 19216 2741 20330 2751
rect 20896 2741 20906 2751
rect 22240 2741 22250 2751
rect 5368 2717 9290 2727
rect 9304 2717 15650 2727
rect 17608 2717 17654 2727
rect 5416 2693 6722 2703
rect 6736 2693 9890 2703
rect 9904 2693 23954 2703
rect 5560 2669 9794 2679
rect 9808 2669 11594 2679
rect 11608 2669 16562 2679
rect 16576 2669 17858 2679
rect 17872 2669 21986 2679
rect 5752 2645 6266 2655
rect 6280 2645 14066 2655
rect 14080 2645 21674 2655
rect 21688 2645 25250 2655
rect 5848 2621 10154 2631
rect 10264 2621 11498 2631
rect 11656 2621 26437 2631
rect 6112 2597 13394 2607
rect 13888 2597 14138 2607
rect 14152 2597 24698 2607
rect 6208 2573 14090 2583
rect 14200 2573 14786 2583
rect 15112 2573 24890 2583
rect 6520 2549 6530 2559
rect 6640 2549 9170 2559
rect 9184 2549 17930 2559
rect 17944 2549 23426 2559
rect 6568 2525 11426 2535
rect 11440 2525 12254 2535
rect 12268 2525 22850 2535
rect 6976 2501 15866 2511
rect 15880 2501 19490 2511
rect 7000 2477 16610 2487
rect 7336 2453 7394 2463
rect 7528 2453 8234 2463
rect 8416 2453 23546 2463
rect 7360 2429 19322 2439
rect 7384 2405 9770 2415
rect 9880 2405 12098 2415
rect 12112 2405 12338 2415
rect 12352 2405 13130 2415
rect 13144 2405 13490 2415
rect 13504 2405 14714 2415
rect 14728 2405 15626 2415
rect 15640 2405 15770 2415
rect 15784 2405 16346 2415
rect 16360 2405 16586 2415
rect 16600 2405 18794 2415
rect 18808 2405 22562 2415
rect 7648 2381 17822 2391
rect 17836 2381 20330 2391
rect 20344 2381 23258 2391
rect 7720 2357 7754 2367
rect 7816 2357 10658 2367
rect 10720 2357 20114 2367
rect 20128 2357 22466 2367
rect 7768 2333 15962 2343
rect 15976 2333 23114 2343
rect 7864 2309 21626 2319
rect 21640 2309 25658 2319
rect 7888 2285 26437 2295
rect 8128 2261 21002 2271
rect 25672 2261 25778 2271
rect 8224 2237 15530 2247
rect 15544 2237 22418 2247
rect 8536 2213 24698 2223
rect 8584 2189 8594 2199
rect 8704 2189 18650 2199
rect 18664 2189 24386 2199
rect 8608 2165 13586 2175
rect 13936 2165 15602 2175
rect 15976 2165 16034 2175
rect 16600 2165 17546 2175
rect 8752 2141 23594 2151
rect 8896 2117 8930 2127
rect 8992 2117 15674 2127
rect 23608 2117 23798 2127
rect 8968 2093 13442 2103
rect 13456 2093 14354 2103
rect 14368 2093 20018 2103
rect 9088 2069 15074 2079
rect 9280 2045 10634 2055
rect 10648 2045 16490 2055
rect 16504 2045 18026 2055
rect 18040 2045 18302 2055
rect 18316 2045 21170 2055
rect 21184 2045 23090 2055
rect 23104 2045 25178 2055
rect 9400 2021 18950 2031
rect 18964 2021 19610 2031
rect 19624 2021 19898 2031
rect 19912 2021 20282 2031
rect 20296 2021 23882 2031
rect 23896 2021 25058 2031
rect 25072 2021 25586 2031
rect 9472 1997 12170 2007
rect 12256 1997 18770 2007
rect 18784 1997 25898 2007
rect 9784 1973 12962 1983
rect 13072 1973 13322 1983
rect 13384 1973 23186 1983
rect 10480 1949 21242 1959
rect 23104 1949 24026 1959
rect 10528 1925 15026 1935
rect 21184 1925 21206 1935
rect 10552 1901 10562 1911
rect 10624 1901 17714 1911
rect 17728 1901 22754 1911
rect 10576 1877 11258 1887
rect 11272 1877 14234 1887
rect 14248 1877 15338 1887
rect 15352 1877 24170 1887
rect 24184 1877 24722 1887
rect 10744 1853 10778 1863
rect 10912 1853 17450 1863
rect 17464 1853 22514 1863
rect 22768 1853 24050 1863
rect 10984 1829 25394 1839
rect 11488 1805 11666 1815
rect 11728 1805 11930 1815
rect 11944 1805 12074 1815
rect 12304 1805 16634 1815
rect 11752 1781 24602 1791
rect 13360 1757 21434 1767
rect 21448 1757 24818 1767
rect 25779 1728 26019 1738
rect 25779 1705 26019 1715
rect 25779 1667 26019 1692
rect 25779 1022 26019 1047
rect 11416 924 20498 934
rect 11224 900 13466 910
rect 13480 900 24434 910
rect 10456 876 15002 886
rect 15016 876 17138 886
rect 10312 852 20930 862
rect 10264 828 13322 838
rect 13768 828 22562 838
rect 10096 804 15890 814
rect 10024 780 11594 790
rect 12352 780 21290 790
rect 9928 756 14978 766
rect 17656 756 22250 766
rect 9832 732 21338 742
rect 9208 708 15074 718
rect 16744 708 19610 718
rect 20200 708 25778 718
rect 9040 684 18938 694
rect 19768 682 19786 696
rect 19888 684 20978 694
rect 8728 660 15578 670
rect 16360 660 22418 670
rect 8680 636 15146 646
rect 15472 636 22178 646
rect 8536 612 21722 622
rect 8440 588 22034 598
rect 8392 564 24818 574
rect 8320 540 19946 550
rect 19960 540 23810 550
rect 8104 516 21026 526
rect 25768 516 25802 526
rect 8008 492 25514 502
rect 25720 492 26437 502
rect 7696 468 11858 478
rect 11968 468 13034 478
rect 13168 468 21050 478
rect 23176 468 25754 478
rect 7684 444 22346 454
rect 7096 420 15818 430
rect 6736 396 6914 406
rect 6928 396 17834 406
rect 6328 372 21482 382
rect 5704 348 9626 358
rect 9736 348 17474 358
rect 17488 348 23546 358
rect 5512 324 13610 334
rect 13792 324 14066 334
rect 14176 324 22922 334
rect 5440 300 22706 310
rect 4960 276 7178 286
rect 7480 276 10490 286
rect 10672 276 16154 286
rect 4912 252 11426 262
rect 13024 252 15242 262
rect 4504 228 11018 238
rect 11152 228 24770 238
rect 4456 204 18818 214
rect 4432 180 10346 190
rect 10432 180 12146 190
rect 13288 180 17906 190
rect 2440 156 7154 166
rect 7504 156 12866 166
rect 12880 156 14954 166
rect 1672 132 9362 142
rect 9568 132 17954 142
rect 1648 108 17330 118
rect 1624 84 2546 94
rect 4144 84 4394 94
rect 4408 84 5714 94
rect 5848 84 9578 94
rect 9808 84 15770 94
rect 84 60 21938 70
rect 25816 60 26437 70
rect 84 36 1706 46
rect 1840 36 5042 46
rect 5344 36 14306 46
rect 25768 36 26437 46
rect 6520 12 19898 22
rect 25792 12 26437 22
<< m2contact >>
rect 21722 8036 21736 8050
rect 12746 8012 12760 8026
rect 19454 8012 19468 8026
rect 21038 8012 21052 8026
rect 24434 8012 24448 8026
rect 8474 7988 8488 8002
rect 9362 7988 9376 8002
rect 12170 7988 12184 8002
rect 14786 7988 14800 8002
rect 17690 7988 17704 8002
rect 17882 7988 17896 8002
rect 26066 7988 26080 8002
rect 3626 7964 3640 7978
rect 4046 7964 4060 7978
rect 5234 7964 5248 7978
rect 7274 7964 7288 7978
rect 9986 7964 10000 7978
rect 10250 7964 10264 7978
rect 11354 7964 11368 7978
rect 24746 7964 24760 7978
rect 3482 7940 3496 7954
rect 13022 7940 13036 7954
rect 13922 7940 13936 7954
rect 24278 7940 24292 7954
rect 3266 7916 3280 7930
rect 14630 7916 14644 7930
rect 15026 7916 15040 7930
rect 16238 7916 16252 7930
rect 17282 7916 17296 7930
rect 26114 7916 26128 7930
rect 70 7892 84 7906
rect 1682 7892 1696 7906
rect 2378 7892 2392 7906
rect 5330 7892 5344 7906
rect 6290 7892 6304 7906
rect 23474 7892 23488 7906
rect 25994 7892 26008 7906
rect 26042 7892 26056 7906
rect 70 7868 84 7882
rect 2234 7868 2248 7882
rect 3002 7868 3016 7882
rect 5678 7868 5692 7882
rect 7274 7868 7288 7882
rect 15434 7868 15448 7882
rect 16346 7868 16360 7882
rect 18650 7868 18664 7882
rect 20882 7868 20896 7882
rect 21866 7868 21880 7882
rect 3194 7844 3208 7858
rect 6794 7844 6808 7858
rect 7994 7844 8008 7858
rect 8426 7844 8440 7858
rect 12206 7844 12220 7858
rect 12242 7844 12256 7858
rect 22670 7844 22684 7858
rect 26090 7844 26104 7858
rect 26437 7844 26451 7858
rect 4010 7820 4024 7834
rect 11402 7820 11416 7834
rect 11618 7820 11632 7834
rect 26018 7820 26032 7834
rect 26066 7820 26080 7834
rect 26437 7820 26451 7834
rect 12194 7796 12208 7810
rect 14090 7796 14104 7810
rect 17138 7796 17152 7810
rect 26090 7796 26104 7810
rect 26114 7796 26128 7810
rect 26437 7796 26451 7810
rect 14606 7772 14620 7786
rect 15146 7772 15160 7786
rect 15266 7772 15280 7786
rect 25082 7772 25096 7786
rect 26042 7772 26056 7786
rect 26437 7772 26451 7786
rect 18626 7748 18640 7762
rect 23618 7748 23632 7762
rect 26018 7748 26032 7762
rect 26437 7748 26451 7762
rect 12122 6915 12136 6929
rect 12338 6915 12352 6929
rect 20474 6915 20488 6929
rect 20498 6915 20512 6929
rect 12098 6891 12112 6905
rect 25778 6891 25792 6905
rect 12050 6867 12064 6881
rect 20474 6867 20488 6881
rect 11690 6843 11704 6857
rect 15386 6843 15400 6857
rect 22274 6843 22288 6857
rect 22298 6843 22312 6857
rect 11426 6819 11440 6833
rect 11834 6819 11848 6833
rect 12026 6819 12040 6833
rect 12254 6819 12268 6833
rect 12530 6819 12544 6833
rect 22802 6819 22816 6833
rect 10802 6795 10816 6809
rect 12914 6795 12928 6809
rect 22274 6795 22288 6809
rect 10562 6771 10576 6785
rect 14450 6771 14464 6785
rect 21482 6771 21496 6785
rect 10394 6747 10408 6761
rect 16034 6747 16048 6761
rect 16370 6747 16384 6761
rect 21938 6747 21952 6761
rect 23474 6747 23488 6761
rect 10346 6723 10360 6737
rect 19298 6723 19312 6737
rect 10106 6699 10120 6713
rect 11690 6699 11704 6713
rect 12002 6699 12016 6713
rect 24650 6699 24664 6713
rect 9410 6675 9424 6689
rect 9530 6675 9544 6689
rect 9674 6675 9688 6689
rect 25490 6675 25504 6689
rect 9170 6651 9184 6665
rect 21674 6651 21688 6665
rect 8954 6627 8968 6641
rect 21530 6627 21544 6641
rect 8906 6603 8920 6617
rect 8954 6603 8968 6617
rect 9146 6603 9160 6617
rect 20402 6603 20416 6617
rect 8834 6579 8848 6593
rect 16082 6579 16096 6593
rect 8810 6555 8824 6569
rect 13946 6555 13960 6569
rect 8546 6531 8560 6545
rect 11066 6531 11080 6545
rect 11234 6531 11248 6545
rect 16154 6531 16168 6545
rect 21026 6531 21040 6545
rect 22706 6531 22720 6545
rect 8546 6507 8560 6521
rect 17906 6507 17920 6521
rect 8474 6483 8488 6497
rect 15578 6483 15592 6497
rect 8474 6459 8488 6473
rect 17690 6459 17704 6473
rect 8330 6435 8344 6449
rect 11810 6435 11824 6449
rect 11906 6435 11920 6449
rect 12170 6435 12184 6449
rect 12482 6435 12496 6449
rect 16538 6435 16552 6449
rect 17402 6435 17416 6449
rect 24746 6435 24760 6449
rect 8162 6411 8176 6425
rect 8234 6411 8248 6425
rect 8306 6411 8320 6425
rect 10058 6411 10072 6425
rect 22058 6411 22072 6425
rect 7922 6387 7936 6401
rect 24074 6387 24088 6401
rect 7898 6363 7912 6377
rect 10970 6363 10984 6377
rect 11282 6363 11296 6377
rect 11330 6363 11344 6377
rect 11378 6363 11392 6377
rect 20834 6363 20848 6377
rect 7874 6339 7888 6353
rect 22490 6339 22504 6353
rect 7826 6315 7840 6329
rect 25538 6315 25552 6329
rect 7442 6291 7456 6305
rect 8618 6291 8632 6305
rect 8930 6291 8944 6305
rect 22586 6291 22600 6305
rect 7394 6267 7408 6281
rect 21122 6267 21136 6281
rect 7274 6243 7288 6257
rect 7970 6243 7984 6257
rect 8042 6243 8056 6257
rect 19418 6243 19432 6257
rect 7226 6219 7240 6233
rect 10778 6219 10792 6233
rect 10850 6219 10864 6233
rect 11450 6219 11464 6233
rect 11642 6219 11656 6233
rect 20066 6219 20080 6233
rect 7226 6195 7240 6209
rect 19226 6195 19240 6209
rect 7178 6171 7192 6185
rect 23930 6171 23944 6185
rect 7130 6147 7144 6161
rect 11954 6147 11968 6161
rect 14834 6147 14848 6161
rect 25562 6147 25576 6161
rect 6866 6123 6880 6137
rect 9482 6123 9496 6137
rect 12362 6123 12376 6137
rect 13826 6123 13840 6137
rect 16610 6123 16624 6137
rect 16634 6123 16648 6137
rect 17330 6123 17344 6137
rect 18938 6123 18952 6137
rect 22970 6123 22984 6137
rect 23066 6123 23080 6137
rect 6818 6099 6832 6113
rect 22970 6099 22984 6113
rect 6722 6075 6736 6089
rect 22106 6075 22120 6089
rect 6698 6051 6712 6065
rect 6722 6051 6736 6065
rect 6794 6051 6808 6065
rect 6842 6051 6856 6065
rect 6890 6051 6904 6065
rect 17738 6051 17752 6065
rect 25514 6051 25528 6065
rect 25610 6051 25624 6065
rect 25826 6051 25840 6065
rect 6674 6027 6688 6041
rect 8018 6027 8032 6041
rect 8066 6027 8080 6041
rect 13322 6027 13336 6041
rect 16058 6027 16072 6041
rect 16346 6027 16360 6041
rect 16562 6027 16576 6041
rect 23282 6027 23296 6041
rect 25610 6027 25624 6041
rect 6458 6003 6472 6017
rect 15218 6003 15232 6017
rect 21626 6003 21640 6017
rect 23306 6003 23320 6017
rect 6362 5979 6376 5993
rect 7394 5979 7408 5993
rect 7682 5979 7696 5993
rect 8666 5979 8680 5993
rect 12002 5979 12016 5993
rect 24938 5979 24952 5993
rect 25802 5979 25816 5993
rect 6314 5955 6328 5969
rect 6962 5955 6976 5969
rect 7010 5955 7024 5969
rect 19778 5955 19792 5969
rect 6146 5931 6160 5945
rect 14114 5931 14128 5945
rect 15194 5931 15208 5945
rect 17882 5931 17896 5945
rect 6050 5907 6064 5921
rect 7322 5907 7336 5921
rect 8858 5907 8872 5921
rect 10946 5907 10960 5921
rect 16202 5907 16216 5921
rect 18554 5907 18568 5921
rect 21074 5907 21088 5921
rect 6002 5883 6016 5897
rect 16442 5883 16456 5897
rect 16490 5883 16504 5897
rect 24938 5883 24952 5897
rect 5954 5859 5968 5873
rect 9002 5859 9016 5873
rect 9050 5859 9064 5873
rect 9170 5859 9184 5873
rect 9314 5859 9328 5873
rect 25634 5859 25648 5873
rect 5954 5835 5968 5849
rect 7034 5835 7048 5849
rect 7082 5835 7096 5849
rect 10562 5835 10576 5849
rect 23402 5835 23416 5849
rect 25346 5835 25360 5849
rect 25418 5835 25432 5849
rect 5786 5811 5800 5825
rect 8594 5811 8608 5825
rect 8786 5811 8800 5825
rect 19034 5811 19048 5825
rect 25298 5811 25312 5825
rect 25322 5811 25336 5825
rect 25754 5811 25768 5825
rect 25874 5811 25888 5825
rect 5786 5787 5800 5801
rect 12578 5787 12592 5801
rect 12650 5787 12664 5801
rect 13562 5787 13576 5801
rect 15986 5787 16000 5801
rect 21290 5787 21304 5801
rect 24026 5787 24040 5801
rect 24506 5787 24520 5801
rect 25730 5787 25744 5801
rect 5690 5763 5704 5777
rect 15194 5763 15208 5777
rect 16010 5763 16024 5777
rect 25754 5763 25768 5777
rect 5666 5739 5680 5753
rect 5690 5739 5704 5753
rect 5762 5739 5776 5753
rect 6530 5739 6544 5753
rect 6578 5739 6592 5753
rect 7034 5739 7048 5753
rect 8066 5739 8080 5753
rect 11618 5739 11632 5753
rect 16178 5739 16192 5753
rect 18074 5739 18088 5753
rect 18854 5739 18868 5753
rect 19178 5739 19192 5753
rect 20690 5739 20704 5753
rect 25346 5739 25360 5753
rect 5642 5715 5656 5729
rect 19046 5715 19060 5729
rect 25298 5715 25312 5729
rect 5642 5691 5656 5705
rect 15482 5691 15496 5705
rect 15698 5691 15712 5705
rect 25418 5691 25432 5705
rect 5594 5667 5608 5681
rect 8282 5667 8296 5681
rect 10154 5667 10168 5681
rect 10202 5667 10216 5681
rect 23978 5667 23992 5681
rect 5594 5643 5608 5657
rect 6170 5643 6184 5657
rect 6218 5643 6232 5657
rect 16730 5643 16744 5657
rect 17282 5643 17296 5657
rect 17546 5643 17560 5657
rect 5570 5619 5584 5633
rect 13874 5619 13888 5633
rect 15674 5619 15688 5633
rect 24986 5619 25000 5633
rect 5570 5595 5584 5609
rect 25994 5595 26008 5609
rect 5546 5571 5560 5585
rect 6290 5571 6304 5585
rect 6362 5571 6376 5585
rect 6410 5571 6424 5585
rect 10682 5571 10696 5585
rect 10754 5571 10768 5585
rect 21950 5571 21964 5585
rect 5450 5547 5464 5561
rect 16106 5547 16120 5561
rect 16466 5547 16480 5561
rect 23378 5547 23392 5561
rect 5426 5523 5440 5537
rect 6074 5523 6088 5537
rect 18122 5523 18136 5537
rect 5378 5499 5392 5513
rect 11354 5499 11368 5513
rect 18410 5499 18424 5513
rect 25442 5499 25456 5513
rect 5306 5475 5320 5489
rect 11522 5475 11536 5489
rect 18986 5475 19000 5489
rect 21986 5475 22000 5489
rect 5258 5451 5272 5465
rect 16274 5451 16288 5465
rect 16322 5451 16336 5465
rect 20066 5451 20080 5465
rect 5258 5427 5272 5441
rect 9746 5427 9760 5441
rect 10106 5427 10120 5441
rect 19682 5427 19696 5441
rect 5234 5403 5248 5417
rect 7466 5403 7480 5417
rect 9074 5403 9088 5417
rect 10322 5403 10336 5417
rect 12074 5403 12088 5417
rect 14666 5403 14680 5417
rect 17402 5403 17416 5417
rect 20594 5403 20608 5417
rect 21842 5403 21856 5417
rect 25370 5403 25384 5417
rect 5138 5379 5152 5393
rect 7754 5379 7768 5393
rect 21746 5379 21760 5393
rect 4970 5355 4984 5369
rect 6866 5355 6880 5369
rect 10610 5355 10624 5369
rect 18290 5355 18304 5369
rect 4898 5331 4912 5345
rect 12698 5331 12712 5345
rect 13274 5331 13288 5345
rect 19994 5331 20008 5345
rect 4850 5307 4864 5321
rect 11762 5307 11776 5321
rect 11858 5307 11872 5321
rect 22826 5307 22840 5321
rect 4802 5283 4816 5297
rect 7346 5283 7360 5297
rect 13370 5283 13384 5297
rect 20138 5283 20152 5297
rect 4778 5259 4792 5273
rect 11882 5259 11896 5273
rect 11978 5259 11992 5273
rect 20618 5259 20632 5273
rect 4658 5235 4672 5249
rect 8330 5235 8344 5249
rect 11666 5235 11680 5249
rect 11738 5235 11752 5249
rect 14618 5235 14632 5249
rect 15530 5235 15544 5249
rect 23786 5235 23800 5249
rect 4610 5211 4624 5225
rect 7826 5211 7840 5225
rect 18626 5211 18640 5225
rect 24554 5211 24568 5225
rect 4586 5187 4600 5201
rect 9218 5187 9232 5201
rect 12674 5187 12688 5201
rect 13250 5187 13264 5201
rect 13442 5187 13456 5201
rect 13514 5187 13528 5201
rect 13586 5187 13600 5201
rect 14642 5187 14656 5201
rect 14714 5187 14728 5201
rect 15314 5187 15328 5201
rect 15506 5187 15520 5201
rect 15554 5187 15568 5201
rect 15770 5187 15784 5201
rect 15914 5187 15928 5201
rect 19274 5187 19288 5201
rect 4538 5163 4552 5177
rect 25706 5163 25720 5177
rect 4346 5139 4360 5153
rect 4658 5139 4672 5153
rect 9002 5139 9016 5153
rect 9674 5139 9688 5153
rect 11138 5139 11152 5153
rect 22106 5139 22120 5153
rect 23882 5139 23896 5153
rect 4322 5115 4336 5129
rect 23738 5115 23752 5129
rect 4298 5091 4312 5105
rect 13706 5091 13720 5105
rect 13922 5091 13936 5105
rect 21458 5091 21472 5105
rect 21698 5091 21712 5105
rect 4250 5067 4264 5081
rect 23018 5067 23032 5081
rect 4226 5043 4240 5057
rect 9410 5043 9424 5057
rect 9626 5043 9640 5057
rect 18266 5043 18280 5057
rect 22874 5043 22888 5057
rect 4130 5019 4144 5033
rect 25850 5019 25864 5033
rect 4082 4995 4096 5009
rect 13298 4995 13312 5009
rect 13394 4995 13408 5009
rect 15410 4995 15424 5009
rect 15458 4995 15472 5009
rect 20858 4995 20872 5009
rect 23474 4995 23488 5009
rect 4082 4971 4096 4985
rect 17642 4971 17656 4985
rect 23354 4971 23368 4985
rect 23438 4971 23452 4985
rect 4058 4947 4072 4961
rect 13106 4947 13120 4961
rect 13202 4947 13216 4961
rect 23570 4947 23584 4961
rect 3986 4923 4000 4937
rect 7010 4923 7024 4937
rect 11186 4923 11200 4937
rect 12218 4923 12232 4937
rect 13226 4923 13240 4937
rect 14594 4923 14608 4937
rect 15434 4923 15448 4937
rect 18194 4923 18208 4937
rect 19922 4923 19936 4937
rect 23114 4923 23128 4937
rect 23234 4923 23248 4937
rect 23354 4923 23368 4937
rect 23834 4923 23848 4937
rect 3890 4899 3904 4913
rect 18242 4899 18256 4913
rect 19970 4899 19984 4913
rect 20306 4899 20320 4913
rect 3866 4875 3880 4889
rect 7562 4875 7576 4889
rect 19970 4875 19984 4889
rect 3818 4851 3832 4865
rect 17618 4851 17632 4865
rect 23762 4851 23776 4865
rect 3794 4827 3808 4841
rect 7586 4827 7600 4841
rect 7706 4827 7720 4841
rect 9938 4827 9952 4841
rect 14282 4827 14296 4841
rect 18218 4827 18232 4841
rect 19538 4827 19552 4841
rect 23162 4827 23176 4841
rect 24146 4827 24160 4841
rect 3770 4803 3784 4817
rect 7106 4803 7120 4817
rect 9242 4803 9256 4817
rect 9554 4803 9568 4817
rect 15890 4803 15904 4817
rect 17378 4803 17392 4817
rect 20570 4803 20584 4817
rect 3722 4779 3736 4793
rect 4106 4779 4120 4793
rect 4154 4779 4168 4793
rect 4466 4779 4480 4793
rect 4538 4779 4552 4793
rect 16298 4779 16312 4793
rect 16418 4779 16432 4793
rect 18746 4779 18760 4793
rect 22682 4779 22696 4793
rect 22922 4779 22936 4793
rect 3698 4755 3712 4769
rect 4226 4755 4240 4769
rect 6818 4755 6832 4769
rect 7970 4755 7984 4769
rect 7994 4755 8008 4769
rect 8090 4755 8104 4769
rect 9506 4755 9520 4769
rect 16130 4755 16144 4769
rect 19010 4755 19024 4769
rect 20258 4755 20272 4769
rect 22682 4755 22696 4769
rect 24098 4755 24112 4769
rect 3674 4731 3688 4745
rect 4850 4731 4864 4745
rect 7514 4731 7528 4745
rect 7778 4731 7792 4745
rect 16106 4731 16120 4745
rect 23498 4731 23512 4745
rect 3650 4707 3664 4721
rect 9698 4707 9712 4721
rect 12818 4707 12832 4721
rect 13850 4707 13864 4721
rect 22202 4707 22216 4721
rect 23042 4707 23056 4721
rect 3578 4683 3592 4697
rect 22442 4683 22456 4697
rect 3530 4659 3544 4673
rect 10922 4659 10936 4673
rect 14474 4659 14488 4673
rect 17354 4659 17368 4673
rect 18410 4659 18424 4673
rect 3530 4635 3544 4649
rect 8210 4635 8224 4649
rect 8258 4635 8272 4649
rect 10178 4635 10192 4649
rect 21506 4635 21520 4649
rect 3386 4611 3400 4625
rect 14234 4611 14248 4625
rect 14378 4611 14392 4625
rect 25082 4611 25096 4625
rect 3362 4587 3376 4601
rect 12146 4587 12160 4601
rect 12434 4587 12448 4601
rect 17810 4587 17824 4601
rect 20042 4587 20056 4601
rect 25322 4587 25336 4601
rect 3338 4563 3352 4577
rect 14498 4563 14512 4577
rect 14594 4563 14608 4577
rect 14618 4563 14632 4577
rect 14882 4563 14896 4577
rect 20042 4563 20056 4577
rect 22322 4563 22336 4577
rect 22418 4563 22432 4577
rect 3218 4539 3232 4553
rect 3458 4539 3472 4553
rect 7250 4539 7264 4553
rect 15122 4539 15136 4553
rect 18602 4539 18616 4553
rect 20234 4539 20248 4553
rect 24338 4539 24352 4553
rect 3170 4515 3184 4529
rect 5738 4515 5752 4529
rect 14042 4515 14056 4529
rect 19730 4515 19744 4529
rect 22322 4515 22336 4529
rect 23138 4515 23152 4529
rect 23798 4515 23812 4529
rect 3122 4491 3136 4505
rect 3266 4491 3280 4505
rect 8762 4491 8776 4505
rect 10082 4491 10096 4505
rect 13010 4491 13024 4505
rect 16418 4491 16432 4505
rect 21890 4491 21904 4505
rect 22658 4491 22672 4505
rect 25466 4491 25480 4505
rect 3098 4467 3112 4481
rect 21578 4467 21592 4481
rect 21818 4467 21832 4481
rect 23138 4467 23152 4481
rect 3050 4443 3064 4457
rect 12122 4443 12136 4457
rect 12314 4443 12328 4457
rect 15938 4443 15952 4457
rect 17738 4443 17752 4457
rect 17786 4443 17800 4457
rect 17822 4443 17836 4457
rect 20114 4443 20128 4457
rect 20498 4443 20512 4457
rect 21194 4443 21208 4457
rect 24482 4443 24496 4457
rect 3002 4419 3016 4433
rect 5810 4419 5824 4433
rect 6578 4419 6592 4433
rect 8906 4419 8920 4433
rect 12026 4419 12040 4433
rect 17306 4419 17320 4433
rect 17786 4419 17800 4433
rect 18698 4419 18712 4433
rect 18950 4419 18964 4433
rect 19082 4419 19096 4433
rect 19154 4419 19168 4433
rect 19826 4419 19840 4433
rect 19898 4419 19912 4433
rect 20090 4419 20104 4433
rect 22370 4419 22384 4433
rect 2978 4395 2992 4409
rect 6386 4395 6400 4409
rect 18722 4395 18736 4409
rect 18890 4395 18904 4409
rect 22922 4395 22936 4409
rect 2954 4371 2968 4385
rect 8402 4371 8416 4385
rect 8450 4371 8464 4385
rect 8954 4371 8968 4385
rect 9842 4371 9856 4385
rect 10010 4371 10024 4385
rect 17570 4371 17584 4385
rect 18170 4371 18184 4385
rect 18302 4371 18316 4385
rect 18482 4371 18496 4385
rect 22778 4371 22792 4385
rect 22898 4371 22912 4385
rect 22922 4371 22936 4385
rect 2930 4347 2944 4361
rect 21554 4347 21568 4361
rect 21794 4347 21808 4361
rect 22178 4347 22192 4361
rect 22634 4347 22648 4361
rect 24266 4347 24280 4361
rect 24626 4347 24640 4361
rect 24722 4347 24736 4361
rect 25706 4347 25720 4361
rect 25874 4347 25888 4361
rect 2906 4323 2920 4337
rect 4994 4323 5008 4337
rect 5186 4323 5200 4337
rect 8258 4323 8272 4337
rect 13034 4323 13048 4337
rect 15818 4323 15832 4337
rect 18506 4323 18520 4337
rect 18602 4323 18616 4337
rect 25202 4323 25216 4337
rect 2882 4299 2896 4313
rect 4418 4299 4432 4313
rect 5666 4299 5680 4313
rect 8282 4299 8296 4313
rect 20354 4299 20368 4313
rect 21770 4299 21784 4313
rect 22538 4299 22552 4313
rect 22610 4299 22624 4313
rect 26437 4299 26451 4313
rect 2858 4275 2872 4289
rect 7610 4275 7624 4289
rect 10202 4275 10216 4289
rect 11162 4275 11176 4289
rect 11282 4275 11296 4289
rect 18122 4275 18136 4289
rect 24650 4275 24664 4289
rect 2786 4251 2800 4265
rect 4970 4251 4984 4265
rect 5018 4251 5032 4265
rect 11714 4251 11728 4265
rect 11786 4251 11800 4265
rect 12866 4251 12880 4265
rect 21146 4251 21160 4265
rect 21770 4251 21784 4265
rect 21842 4251 21856 4265
rect 21890 4251 21904 4265
rect 21950 4251 21964 4265
rect 22442 4251 22456 4265
rect 22706 4251 22720 4265
rect 2714 4227 2728 4241
rect 21866 4227 21880 4241
rect 2666 4203 2680 4217
rect 7130 4203 7144 4217
rect 11090 4203 11104 4217
rect 16442 4203 16456 4217
rect 23330 4203 23344 4217
rect 2642 4179 2656 4193
rect 8570 4179 8584 4193
rect 8642 4179 8656 4193
rect 18338 4179 18352 4193
rect 22250 4179 22264 4193
rect 24362 4179 24376 4193
rect 2594 4155 2608 4169
rect 11090 4155 11104 4169
rect 11306 4155 11320 4169
rect 11426 4155 11440 4169
rect 11570 4155 11584 4169
rect 13994 4155 14008 4169
rect 19370 4155 19384 4169
rect 20762 4155 20776 4169
rect 23666 4155 23680 4169
rect 2522 4131 2536 4145
rect 3962 4131 3976 4145
rect 6626 4131 6640 4145
rect 8162 4131 8176 4145
rect 10226 4131 10240 4145
rect 13154 4131 13168 4145
rect 15842 4131 15856 4145
rect 19826 4131 19840 4145
rect 21266 4131 21280 4145
rect 21602 4131 21616 4145
rect 2450 4107 2464 4121
rect 7442 4107 7456 4121
rect 8882 4107 8896 4121
rect 13514 4107 13528 4121
rect 18530 4107 18544 4121
rect 23210 4107 23224 4121
rect 2402 4083 2416 4097
rect 13106 4083 13120 4097
rect 20714 4083 20728 4097
rect 20810 4083 20824 4097
rect 21722 4083 21736 4097
rect 2330 4059 2344 4073
rect 5210 4059 5224 4073
rect 7946 4059 7960 4073
rect 9122 4059 9136 4073
rect 14858 4059 14872 4073
rect 17690 4059 17704 4073
rect 20450 4059 20464 4073
rect 21074 4059 21088 4073
rect 23066 4059 23080 4073
rect 2282 4035 2296 4049
rect 7202 4035 7216 4049
rect 12050 4035 12064 4049
rect 15650 4035 15664 4049
rect 16010 4035 16024 4049
rect 23618 4035 23632 4049
rect 2186 4011 2200 4025
rect 22154 4011 22168 4025
rect 2162 3987 2176 4001
rect 18818 3987 18832 4001
rect 19010 3987 19024 4001
rect 19046 3987 19060 4001
rect 21266 3987 21280 4001
rect 21290 3987 21304 4001
rect 2090 3963 2104 3977
rect 10418 3963 10432 3977
rect 12794 3963 12808 3977
rect 25154 3963 25168 3977
rect 2042 3939 2056 3953
rect 6794 3939 6808 3953
rect 7730 3939 7744 3953
rect 10994 3939 11008 3953
rect 11354 3939 11368 3953
rect 16466 3939 16480 3953
rect 21242 3939 21256 3953
rect 21386 3939 21400 3953
rect 1970 3915 1984 3929
rect 2186 3915 2200 3929
rect 4370 3915 4384 3929
rect 8738 3915 8752 3929
rect 10826 3915 10840 3929
rect 11018 3915 11032 3929
rect 13178 3915 13192 3929
rect 17618 3915 17632 3929
rect 18362 3915 18376 3929
rect 19802 3915 19816 3929
rect 20666 3915 20680 3929
rect 1946 3891 1960 3905
rect 9458 3891 9472 3905
rect 11546 3891 11560 3905
rect 12194 3891 12208 3905
rect 22586 3891 22600 3905
rect 23234 3891 23248 3905
rect 1898 3867 1912 3881
rect 5066 3867 5080 3881
rect 12722 3867 12736 3881
rect 20786 3867 20800 3881
rect 1874 3843 1888 3857
rect 3938 3843 3952 3857
rect 6554 3843 6568 3857
rect 9434 3843 9448 3857
rect 9866 3843 9880 3857
rect 11042 3843 11056 3857
rect 13538 3843 13552 3857
rect 18578 3843 18592 3857
rect 23714 3843 23728 3857
rect 1850 3819 1864 3833
rect 2738 3819 2752 3833
rect 16226 3819 16240 3833
rect 22346 3819 22360 3833
rect 1802 3795 1816 3809
rect 5858 3795 5872 3809
rect 5906 3795 5920 3809
rect 22538 3795 22552 3809
rect 1754 3771 1768 3785
rect 7802 3771 7816 3785
rect 9314 3771 9328 3785
rect 9362 3771 9376 3785
rect 21206 3771 21220 3785
rect 1706 3747 1720 3761
rect 20282 3747 20296 3761
rect 1634 3723 1648 3737
rect 1730 3723 1744 3737
rect 2210 3723 2224 3737
rect 2234 3723 2248 3737
rect 3338 3723 3352 3737
rect 4754 3723 4768 3737
rect 5090 3723 5104 3737
rect 9050 3723 9064 3737
rect 14570 3723 14584 3737
rect 15218 3723 15232 3737
rect 16226 3723 16240 3737
rect 20162 3723 20176 3737
rect 23858 3723 23872 3737
rect 25922 3723 25936 3737
rect 1610 3699 1624 3713
rect 21914 3699 21928 3713
rect 22394 3699 22408 3713
rect 70 3675 84 3689
rect 2378 3675 2392 3689
rect 7370 3675 7384 3689
rect 13082 3675 13096 3689
rect 23906 3675 23920 3689
rect 70 3651 84 3665
rect 13418 3651 13432 3665
rect 13658 3651 13672 3665
rect 17474 3651 17488 3665
rect 18458 3651 18472 3665
rect 19130 3651 19144 3665
rect 20210 3651 20224 3665
rect 23906 3651 23920 3665
rect 24146 3651 24160 3665
rect 1994 3627 2008 3641
rect 18698 3627 18712 3641
rect 2498 3603 2512 3617
rect 4586 3603 4600 3617
rect 4730 3603 4744 3617
rect 5474 3603 5488 3617
rect 5978 3603 5992 3617
rect 15314 3603 15328 3617
rect 18338 3603 18352 3617
rect 18578 3603 18592 3617
rect 18626 3603 18640 3617
rect 18722 3603 18736 3617
rect 18854 3603 18868 3617
rect 2522 3579 2536 3593
rect 9650 3579 9664 3593
rect 9962 3579 9976 3593
rect 14258 3579 14272 3593
rect 14642 3579 14656 3593
rect 18050 3579 18064 3593
rect 19850 3579 19864 3593
rect 24626 3579 24640 3593
rect 2546 3555 2560 3569
rect 19082 3555 19096 3569
rect 2594 3531 2608 3545
rect 4706 3531 4720 3545
rect 5330 3531 5344 3545
rect 6770 3531 6784 3545
rect 14738 3531 14752 3545
rect 22010 3531 22024 3545
rect 2618 3507 2632 3521
rect 4298 3507 4312 3521
rect 4754 3507 4768 3521
rect 6842 3507 6856 3521
rect 11474 3507 11488 3521
rect 14762 3507 14776 3521
rect 14906 3507 14920 3521
rect 25682 3507 25696 3521
rect 2690 3483 2704 3497
rect 15434 3483 15448 3497
rect 15482 3483 15496 3497
rect 15578 3483 15592 3497
rect 16082 3483 16096 3497
rect 16370 3483 16384 3497
rect 16514 3483 16528 3497
rect 24410 3483 24424 3497
rect 2786 3459 2800 3473
rect 18170 3459 18184 3473
rect 18914 3459 18928 3473
rect 2810 3435 2824 3449
rect 6506 3435 6520 3449
rect 24218 3435 24232 3449
rect 2834 3411 2848 3425
rect 13346 3411 13360 3425
rect 16298 3411 16312 3425
rect 17426 3411 17440 3425
rect 18674 3411 18688 3425
rect 19946 3411 19960 3425
rect 2882 3387 2896 3401
rect 14978 3387 14992 3401
rect 22898 3387 22912 3401
rect 23690 3387 23704 3401
rect 24842 3387 24856 3401
rect 2906 3363 2920 3377
rect 3362 3363 3376 3377
rect 11210 3363 11224 3377
rect 13058 3363 13072 3377
rect 15338 3363 15352 3377
rect 16250 3363 16264 3377
rect 16394 3363 16408 3377
rect 2930 3339 2944 3353
rect 4250 3339 4264 3353
rect 5114 3339 5128 3353
rect 5234 3339 5248 3353
rect 8810 3339 8824 3353
rect 9986 3339 10000 3353
rect 15362 3339 15376 3353
rect 15746 3339 15760 3353
rect 17954 3339 17968 3353
rect 20546 3339 20560 3353
rect 21410 3339 21424 3353
rect 24122 3339 24136 3353
rect 3002 3315 3016 3329
rect 3626 3315 3640 3329
rect 5474 3315 5488 3329
rect 5690 3315 5704 3329
rect 7250 3315 7264 3329
rect 7922 3315 7936 3329
rect 11330 3315 11344 3329
rect 12938 3315 12952 3329
rect 16058 3315 16072 3329
rect 17978 3315 17992 3329
rect 18002 3315 18016 3329
rect 19106 3315 19120 3329
rect 24962 3315 24976 3329
rect 3026 3291 3040 3305
rect 3218 3291 3232 3305
rect 11402 3291 11416 3305
rect 13250 3291 13264 3305
rect 18434 3291 18448 3305
rect 22154 3291 22168 3305
rect 22994 3291 23008 3305
rect 3050 3267 3064 3281
rect 15506 3267 15520 3281
rect 23642 3267 23656 3281
rect 3098 3243 3112 3257
rect 4514 3243 4528 3257
rect 6674 3243 6688 3257
rect 19874 3243 19888 3257
rect 3122 3219 3136 3233
rect 6938 3219 6952 3233
rect 14882 3219 14896 3233
rect 19634 3219 19648 3233
rect 21818 3219 21832 3233
rect 3170 3195 3184 3209
rect 9146 3195 9160 3209
rect 22730 3195 22744 3209
rect 3386 3171 3400 3185
rect 10298 3171 10312 3185
rect 15794 3171 15808 3185
rect 18146 3171 18160 3185
rect 19154 3171 19168 3185
rect 20234 3171 20248 3185
rect 24674 3171 24688 3185
rect 3410 3147 3424 3161
rect 14954 3147 14968 3161
rect 18218 3147 18232 3161
rect 3434 3123 3448 3137
rect 9506 3123 9520 3137
rect 9722 3123 9736 3137
rect 14402 3123 14416 3137
rect 14546 3123 14560 3137
rect 15722 3123 15736 3137
rect 17654 3123 17668 3137
rect 20186 3123 20200 3137
rect 21314 3123 21328 3137
rect 3554 3099 3568 3113
rect 18842 3099 18856 3113
rect 3890 3075 3904 3089
rect 6698 3075 6712 3089
rect 9266 3075 9280 3089
rect 10730 3075 10744 3089
rect 10802 3075 10816 3089
rect 11906 3075 11920 3089
rect 12458 3075 12472 3089
rect 13634 3075 13648 3089
rect 17282 3075 17296 3089
rect 18098 3075 18112 3089
rect 19034 3075 19048 3089
rect 21362 3075 21376 3089
rect 3914 3051 3928 3065
rect 8138 3051 8152 3065
rect 8186 3051 8200 3065
rect 9890 3051 9904 3065
rect 9962 3051 9976 3065
rect 17522 3051 17536 3065
rect 21362 3051 21376 3065
rect 21746 3051 21760 3065
rect 4010 3027 4024 3041
rect 5018 3027 5032 3041
rect 5138 3027 5152 3041
rect 17498 3027 17512 3041
rect 4202 3003 4216 3017
rect 15362 3003 15376 3017
rect 15746 3003 15760 3017
rect 15818 3003 15832 3017
rect 17522 3003 17536 3017
rect 17882 3003 17896 3017
rect 4274 2979 4288 2993
rect 6746 2979 6760 2993
rect 6914 2979 6928 2993
rect 8378 2979 8392 2993
rect 15098 2979 15112 2993
rect 15290 2979 15304 2993
rect 19202 2979 19216 2993
rect 20906 2979 20920 2993
rect 22298 2979 22312 2993
rect 22658 2979 22672 2993
rect 4490 2955 4504 2969
rect 25562 2955 25576 2969
rect 4610 2931 4624 2945
rect 7418 2931 7432 2945
rect 9530 2931 9544 2945
rect 10538 2931 10552 2945
rect 10874 2931 10888 2945
rect 11306 2931 11320 2945
rect 15554 2931 15568 2945
rect 17762 2931 17776 2945
rect 21650 2931 21664 2945
rect 22130 2931 22144 2945
rect 22466 2931 22480 2945
rect 24482 2931 24496 2945
rect 4634 2907 4648 2921
rect 21410 2907 21424 2921
rect 22130 2907 22144 2921
rect 22178 2907 22192 2921
rect 4682 2883 4696 2897
rect 26437 2883 26451 2897
rect 4730 2859 4744 2873
rect 20882 2859 20896 2873
rect 25274 2859 25288 2873
rect 4826 2835 4840 2849
rect 7562 2835 7576 2849
rect 10442 2835 10456 2849
rect 11810 2835 11824 2849
rect 22922 2835 22936 2849
rect 23522 2835 23536 2849
rect 4874 2811 4888 2825
rect 6482 2811 6496 2825
rect 13202 2811 13216 2825
rect 14810 2811 14824 2825
rect 20378 2811 20392 2825
rect 22226 2811 22240 2825
rect 24002 2811 24016 2825
rect 25130 2811 25144 2825
rect 4994 2787 5008 2801
rect 25946 2787 25960 2801
rect 5186 2763 5200 2777
rect 14690 2763 14704 2777
rect 18650 2763 18664 2777
rect 20306 2763 20320 2777
rect 23438 2763 23452 2777
rect 25034 2763 25048 2777
rect 5306 2739 5320 2753
rect 9098 2739 9112 2753
rect 17594 2739 17608 2753
rect 19202 2739 19216 2753
rect 20330 2739 20344 2753
rect 20882 2739 20896 2753
rect 20906 2739 20920 2753
rect 22226 2739 22240 2753
rect 22250 2739 22264 2753
rect 5354 2715 5368 2729
rect 9290 2715 9304 2729
rect 15650 2715 15664 2729
rect 17594 2715 17608 2729
rect 17654 2715 17668 2729
rect 5402 2691 5416 2705
rect 6722 2691 6736 2705
rect 9890 2691 9904 2705
rect 23954 2691 23968 2705
rect 5546 2667 5560 2681
rect 9794 2667 9808 2681
rect 11594 2667 11608 2681
rect 16562 2667 16576 2681
rect 17858 2667 17872 2681
rect 21986 2667 22000 2681
rect 5738 2643 5752 2657
rect 6266 2643 6280 2657
rect 14066 2643 14080 2657
rect 21674 2643 21688 2657
rect 25250 2643 25264 2657
rect 5834 2619 5848 2633
rect 10154 2619 10168 2633
rect 10250 2619 10264 2633
rect 11498 2619 11512 2633
rect 11642 2619 11656 2633
rect 26437 2619 26451 2633
rect 6098 2595 6112 2609
rect 13394 2595 13408 2609
rect 13874 2595 13888 2609
rect 14138 2595 14152 2609
rect 24698 2595 24712 2609
rect 6194 2571 6208 2585
rect 14090 2571 14104 2585
rect 14186 2571 14200 2585
rect 14786 2571 14800 2585
rect 15098 2571 15112 2585
rect 24890 2571 24904 2585
rect 6506 2547 6520 2561
rect 6530 2547 6544 2561
rect 6626 2547 6640 2561
rect 9170 2547 9184 2561
rect 17930 2547 17944 2561
rect 23426 2547 23440 2561
rect 6554 2523 6568 2537
rect 11426 2523 11440 2537
rect 12254 2523 12268 2537
rect 22850 2523 22864 2537
rect 6962 2499 6976 2513
rect 15866 2499 15880 2513
rect 19490 2499 19504 2513
rect 6986 2475 7000 2489
rect 16610 2475 16624 2489
rect 7322 2451 7336 2465
rect 7394 2451 7408 2465
rect 7514 2451 7528 2465
rect 8234 2451 8248 2465
rect 8402 2451 8416 2465
rect 23546 2451 23560 2465
rect 7346 2427 7360 2441
rect 19322 2427 19336 2441
rect 7370 2403 7384 2417
rect 9770 2403 9784 2417
rect 9866 2403 9880 2417
rect 12098 2403 12112 2417
rect 12338 2403 12352 2417
rect 13130 2403 13144 2417
rect 13490 2403 13504 2417
rect 14714 2403 14728 2417
rect 15626 2403 15640 2417
rect 15770 2403 15784 2417
rect 16346 2403 16360 2417
rect 16586 2403 16600 2417
rect 18794 2403 18808 2417
rect 22562 2403 22576 2417
rect 7634 2379 7648 2393
rect 17822 2379 17836 2393
rect 20330 2379 20344 2393
rect 23258 2379 23272 2393
rect 7706 2355 7720 2369
rect 7754 2355 7768 2369
rect 7802 2355 7816 2369
rect 10658 2355 10672 2369
rect 10706 2355 10720 2369
rect 20114 2355 20128 2369
rect 22466 2355 22480 2369
rect 7754 2331 7768 2345
rect 15962 2331 15976 2345
rect 23114 2331 23128 2345
rect 7850 2307 7864 2321
rect 21626 2307 21640 2321
rect 25658 2307 25672 2321
rect 7874 2283 7888 2297
rect 26437 2283 26451 2297
rect 8114 2259 8128 2273
rect 21002 2259 21016 2273
rect 25658 2259 25672 2273
rect 25778 2259 25792 2273
rect 8210 2235 8224 2249
rect 15530 2235 15544 2249
rect 22418 2235 22432 2249
rect 8522 2211 8536 2225
rect 24698 2211 24712 2225
rect 8570 2187 8584 2201
rect 8594 2187 8608 2201
rect 8690 2187 8704 2201
rect 18650 2187 18664 2201
rect 24386 2187 24400 2201
rect 8594 2163 8608 2177
rect 13586 2163 13600 2177
rect 13922 2163 13936 2177
rect 15602 2163 15616 2177
rect 15962 2163 15976 2177
rect 16034 2163 16048 2177
rect 16586 2163 16600 2177
rect 17546 2163 17560 2177
rect 8738 2139 8752 2153
rect 23594 2139 23608 2153
rect 8882 2115 8896 2129
rect 8930 2115 8944 2129
rect 8978 2115 8992 2129
rect 15674 2115 15688 2129
rect 23594 2115 23608 2129
rect 23798 2115 23812 2129
rect 8954 2091 8968 2105
rect 13442 2091 13456 2105
rect 14354 2091 14368 2105
rect 20018 2091 20032 2105
rect 9074 2067 9088 2081
rect 15074 2067 15088 2081
rect 9266 2043 9280 2057
rect 10634 2043 10648 2057
rect 16490 2043 16504 2057
rect 18026 2043 18040 2057
rect 18302 2043 18316 2057
rect 21170 2043 21184 2057
rect 23090 2043 23104 2057
rect 25178 2043 25192 2057
rect 9386 2019 9400 2033
rect 18950 2019 18964 2033
rect 19610 2019 19624 2033
rect 19898 2019 19912 2033
rect 20282 2019 20296 2033
rect 23882 2019 23896 2033
rect 25058 2019 25072 2033
rect 25586 2019 25600 2033
rect 9458 1995 9472 2009
rect 12170 1995 12184 2009
rect 12242 1995 12256 2009
rect 18770 1995 18784 2009
rect 25898 1995 25912 2009
rect 9770 1971 9784 1985
rect 12962 1971 12976 1985
rect 13058 1971 13072 1985
rect 13322 1971 13336 1985
rect 13370 1971 13384 1985
rect 23186 1971 23200 1985
rect 10466 1947 10480 1961
rect 21242 1947 21256 1961
rect 23090 1947 23104 1961
rect 24026 1947 24040 1961
rect 10514 1923 10528 1937
rect 15026 1923 15040 1937
rect 21170 1923 21184 1937
rect 21206 1923 21220 1937
rect 10538 1899 10552 1913
rect 10562 1899 10576 1913
rect 10610 1899 10624 1913
rect 17714 1899 17728 1913
rect 22754 1899 22768 1913
rect 10562 1875 10576 1889
rect 11258 1875 11272 1889
rect 14234 1875 14248 1889
rect 15338 1875 15352 1889
rect 24170 1875 24184 1889
rect 24722 1875 24736 1889
rect 10730 1851 10744 1865
rect 10778 1851 10792 1865
rect 10898 1851 10912 1865
rect 17450 1851 17464 1865
rect 22514 1851 22528 1865
rect 22754 1851 22768 1865
rect 24050 1851 24064 1865
rect 10970 1827 10984 1841
rect 25394 1827 25408 1841
rect 11474 1803 11488 1817
rect 11666 1803 11680 1817
rect 11714 1803 11728 1817
rect 11930 1803 11944 1817
rect 12074 1803 12088 1817
rect 12290 1803 12304 1817
rect 16634 1803 16648 1817
rect 11738 1779 11752 1793
rect 24602 1779 24616 1793
rect 13346 1755 13360 1769
rect 21434 1755 21448 1769
rect 24818 1755 24832 1769
rect 11402 922 11416 936
rect 20498 922 20512 936
rect 11210 898 11224 912
rect 13466 898 13480 912
rect 24434 898 24448 912
rect 10442 874 10456 888
rect 15002 874 15016 888
rect 17138 874 17152 888
rect 10298 850 10312 864
rect 20930 850 20944 864
rect 10250 826 10264 840
rect 13322 826 13336 840
rect 13754 826 13768 840
rect 22562 826 22576 840
rect 10082 802 10096 816
rect 15890 802 15904 816
rect 10010 778 10024 792
rect 11594 778 11608 792
rect 12338 778 12352 792
rect 21290 778 21304 792
rect 9914 754 9928 768
rect 14978 754 14992 768
rect 17642 754 17656 768
rect 22250 754 22264 768
rect 9818 730 9832 744
rect 21338 730 21352 744
rect 9194 706 9208 720
rect 15074 706 15088 720
rect 16730 706 16744 720
rect 19610 706 19624 720
rect 20186 706 20200 720
rect 25778 706 25792 720
rect 9026 682 9040 696
rect 18938 682 18952 696
rect 19754 682 19768 696
rect 19874 682 19888 696
rect 20978 682 20992 696
rect 8714 658 8728 672
rect 15578 658 15592 672
rect 16346 658 16360 672
rect 22418 658 22432 672
rect 8666 634 8680 648
rect 15146 634 15160 648
rect 15458 634 15472 648
rect 22178 634 22192 648
rect 8522 610 8536 624
rect 21722 610 21736 624
rect 8426 586 8440 600
rect 22034 586 22048 600
rect 8378 562 8392 576
rect 24818 562 24832 576
rect 8306 538 8320 552
rect 19946 538 19960 552
rect 23810 538 23824 552
rect 8090 514 8104 528
rect 21026 514 21040 528
rect 25754 514 25768 528
rect 25802 514 25816 528
rect 7994 490 8008 504
rect 25514 490 25528 504
rect 25706 490 25720 504
rect 26437 490 26451 504
rect 7682 466 7696 480
rect 11858 466 11872 480
rect 11954 466 11968 480
rect 13034 466 13048 480
rect 13154 466 13168 480
rect 21050 466 21064 480
rect 23162 466 23176 480
rect 25754 466 25768 480
rect 7670 442 7684 456
rect 22346 442 22360 456
rect 7082 418 7096 432
rect 15818 418 15832 432
rect 6722 394 6736 408
rect 6914 394 6928 408
rect 17834 394 17848 408
rect 6314 370 6328 384
rect 21482 370 21496 384
rect 5690 346 5704 360
rect 9626 346 9640 360
rect 9722 346 9736 360
rect 17474 346 17488 360
rect 23546 346 23560 360
rect 5498 322 5512 336
rect 13610 322 13624 336
rect 13778 322 13792 336
rect 14066 322 14080 336
rect 14162 322 14176 336
rect 22922 322 22936 336
rect 5426 298 5440 312
rect 22706 298 22720 312
rect 4946 274 4960 288
rect 7178 274 7192 288
rect 7466 274 7480 288
rect 10490 274 10504 288
rect 10658 274 10672 288
rect 16154 274 16168 288
rect 4898 250 4912 264
rect 11426 250 11440 264
rect 13010 250 13024 264
rect 15242 250 15256 264
rect 4490 226 4504 240
rect 11018 226 11032 240
rect 11138 226 11152 240
rect 24770 226 24784 240
rect 4442 202 4456 216
rect 18818 202 18832 216
rect 4418 178 4432 192
rect 10346 178 10360 192
rect 10418 178 10432 192
rect 12146 178 12160 192
rect 13274 178 13288 192
rect 17906 178 17920 192
rect 2426 154 2440 168
rect 7154 154 7168 168
rect 7490 154 7504 168
rect 12866 154 12880 168
rect 14954 154 14968 168
rect 1658 130 1672 144
rect 9362 130 9376 144
rect 9554 130 9568 144
rect 17954 130 17968 144
rect 1634 106 1648 120
rect 17330 106 17344 120
rect 1610 82 1624 96
rect 2546 82 2560 96
rect 4130 82 4144 96
rect 4394 82 4408 96
rect 5714 82 5728 96
rect 5834 82 5848 96
rect 9578 82 9592 96
rect 9794 82 9808 96
rect 15770 82 15784 96
rect 70 58 84 72
rect 21938 58 21952 72
rect 25802 58 25816 72
rect 26437 58 26451 72
rect 70 34 84 48
rect 1706 34 1720 48
rect 1826 34 1840 48
rect 5042 34 5056 48
rect 5330 34 5344 48
rect 14306 34 14320 48
rect 25754 34 25768 48
rect 26437 34 26451 48
rect 6506 10 6520 24
rect 19898 10 19912 24
rect 25778 10 25792 24
rect 26437 10 26451 24
<< metal2 >>
rect 0 7893 70 7905
rect 0 7869 70 7881
rect 123 7738 323 8060
rect 339 7738 351 8060
rect 363 7738 375 8060
rect 387 7738 399 8060
rect 411 7738 423 8060
rect 2379 7906 2391 8060
rect 1683 7738 1695 7892
rect 2235 7738 2247 7868
rect 3003 7738 3015 7868
rect 3195 7858 3207 8060
rect 3267 7738 3279 7916
rect 3483 7738 3495 7940
rect 3627 7738 3639 7964
rect 4011 7834 4023 8060
rect 4047 7978 4059 8060
rect 5247 7978 5259 8060
rect 5248 7964 5266 7978
rect 5235 7738 5247 7964
rect 5331 7738 5343 7892
rect 5679 7882 5691 8060
rect 7275 7978 7287 8060
rect 6291 7738 6303 7892
rect 6795 7738 6807 7844
rect 7275 7738 7287 7868
rect 8007 7858 8019 8060
rect 8487 8002 8499 8060
rect 9375 8002 9387 8060
rect 8488 7988 8506 8002
rect 9376 7988 9394 8002
rect 8008 7844 8026 7858
rect 7995 7738 8007 7844
rect 8427 7738 8439 7844
rect 8475 7738 8487 7988
rect 9363 7738 9375 7988
rect 10263 7978 10275 8060
rect 11355 7978 11367 8060
rect 12171 8002 12183 8060
rect 10264 7964 10282 7978
rect 9987 7738 9999 7964
rect 10251 7738 10263 7964
rect 12207 7858 12219 8060
rect 11403 7738 11415 7820
rect 11619 7738 11631 7820
rect 12195 7738 12207 7796
rect 12243 7738 12255 7844
rect 12747 7738 12759 8012
rect 13023 7954 13035 8060
rect 13923 7738 13935 7940
rect 14091 7738 14103 7796
rect 14607 7786 14619 8060
rect 14631 7930 14643 8060
rect 14787 7738 14799 7988
rect 15027 7738 15039 7916
rect 15435 7882 15447 8060
rect 16239 7930 16251 8060
rect 17703 8002 17715 8060
rect 17704 7988 17722 8002
rect 15147 7738 15159 7772
rect 15267 7738 15279 7772
rect 16347 7738 16359 7868
rect 17139 7738 17151 7796
rect 17283 7738 17295 7916
rect 17691 7738 17703 7988
rect 17883 7738 17895 7988
rect 18627 7762 18639 8060
rect 18651 7882 18663 8060
rect 19455 8026 19467 8060
rect 21039 8026 21051 8060
rect 21735 8050 21747 8060
rect 21736 8036 21754 8050
rect 20883 7738 20895 7868
rect 21723 7738 21735 8036
rect 21867 7882 21879 8060
rect 22671 7858 22683 8060
rect 23475 7906 23487 8060
rect 24279 7954 24291 8060
rect 23619 7738 23631 7748
rect 24435 7738 24447 8012
rect 24747 7738 24759 7964
rect 25083 7786 25095 8060
rect 25995 7738 26007 7892
rect 26019 7762 26031 7820
rect 26043 7786 26055 7892
rect 26067 7834 26079 7988
rect 26091 7810 26103 7844
rect 26115 7810 26127 7916
rect 26139 7738 26339 8060
rect 26451 7845 26521 7857
rect 26451 7821 26521 7833
rect 26451 7797 26521 7809
rect 26451 7773 26521 7785
rect 26451 7749 26521 7761
rect 0 3676 70 3688
rect 0 3652 70 3664
rect 123 1745 323 6939
rect 339 1745 351 6939
rect 363 1745 375 6939
rect 387 1745 399 6939
rect 411 1745 423 6939
rect 1611 3713 1623 6939
rect 1635 3737 1647 6939
rect 1707 1745 1719 3747
rect 1731 3737 1743 6939
rect 1755 3785 1767 6939
rect 1803 3809 1815 6939
rect 1851 3833 1863 6939
rect 1875 3857 1887 6939
rect 1899 3881 1911 6939
rect 1947 3905 1959 6939
rect 1971 3929 1983 6939
rect 1995 3641 2007 6939
rect 2043 3953 2055 6939
rect 2091 3977 2103 6939
rect 2163 4001 2175 6939
rect 2187 4025 2199 6939
rect 2187 1745 2199 3915
rect 2211 3737 2223 6939
rect 2283 4049 2295 6939
rect 2331 4073 2343 6939
rect 2403 4097 2415 6939
rect 2451 4121 2463 6939
rect 2523 4145 2535 6939
rect 2235 1745 2247 3723
rect 2379 1745 2391 3675
rect 2499 1745 2511 3603
rect 2523 1745 2535 3579
rect 2547 3569 2559 6939
rect 2595 4169 2607 6939
rect 2643 4193 2655 6939
rect 2667 4217 2679 6939
rect 2595 1745 2607 3531
rect 2619 1745 2631 3507
rect 2691 3497 2703 6939
rect 2715 1745 2727 4227
rect 2739 3833 2751 6939
rect 2787 4265 2799 6939
rect 2859 4289 2871 6939
rect 2883 4313 2895 6939
rect 2907 4337 2919 6939
rect 2931 4361 2943 6939
rect 2979 4409 2991 6939
rect 3003 4433 3015 6939
rect 3051 4457 3063 6939
rect 3099 4481 3111 6939
rect 3123 4505 3135 6939
rect 3171 4529 3183 6939
rect 3219 4553 3231 6939
rect 3339 4577 3351 6939
rect 3363 4601 3375 6939
rect 3387 4625 3399 6939
rect 2787 1745 2799 3459
rect 2811 1745 2823 3435
rect 2835 1745 2847 3411
rect 2883 1745 2895 3387
rect 2907 1745 2919 3363
rect 2931 1745 2943 3339
rect 2955 1745 2967 4371
rect 3003 1745 3015 3315
rect 3027 1745 3039 3291
rect 3051 1745 3063 3267
rect 3099 1745 3111 3243
rect 3123 1745 3135 3219
rect 3171 1745 3183 3195
rect 3219 1745 3231 3291
rect 3267 1745 3279 4491
rect 3339 1745 3351 3723
rect 3363 1745 3375 3363
rect 3387 1745 3399 3171
rect 3411 1745 3423 3147
rect 3435 3137 3447 6939
rect 3459 4553 3471 6939
rect 3531 4673 3543 6939
rect 3531 1745 3543 4635
rect 3555 3113 3567 6939
rect 3579 4697 3591 6939
rect 3627 3329 3639 6939
rect 3651 4721 3663 6939
rect 3675 4745 3687 6939
rect 3699 4769 3711 6939
rect 3723 4793 3735 6939
rect 3771 4817 3783 6939
rect 3795 4841 3807 6939
rect 3819 4865 3831 6939
rect 3867 4889 3879 6939
rect 3891 4913 3903 6939
rect 3891 1745 3903 3075
rect 3915 3065 3927 6939
rect 3963 4145 3975 6939
rect 3987 4937 3999 6939
rect 3939 1745 3951 3843
rect 4011 3041 4023 6939
rect 4059 4961 4071 6939
rect 4083 5009 4095 6939
rect 4083 1745 4095 4971
rect 4107 4793 4119 6939
rect 4131 5033 4143 6939
rect 4155 4793 4167 6939
rect 4203 3017 4215 6939
rect 4227 5057 4239 6939
rect 4251 5081 4263 6939
rect 4227 1745 4239 4755
rect 4251 1745 4263 3339
rect 4275 2993 4287 6939
rect 4299 5105 4311 6939
rect 4347 5153 4359 6939
rect 4299 1745 4311 3507
rect 4323 1745 4335 5115
rect 4371 3929 4383 6939
rect 4419 4313 4431 6939
rect 4467 4793 4479 6939
rect 4491 2969 4503 6939
rect 4539 5177 4551 6939
rect 4587 5201 4599 6939
rect 4611 5225 4623 6939
rect 4515 1745 4527 3243
rect 4539 1745 4551 4779
rect 4587 1745 4599 3603
rect 4611 1745 4623 2931
rect 4635 2921 4647 6939
rect 4659 5249 4671 6939
rect 4659 1745 4671 5139
rect 4683 2897 4695 6939
rect 4731 3617 4743 6939
rect 4755 3737 4767 6939
rect 4803 5297 4815 6939
rect 4851 5321 4863 6939
rect 4899 5345 4911 6939
rect 4971 5369 4983 6939
rect 4707 1745 4719 3531
rect 4731 1745 4743 2859
rect 4755 1745 4767 3507
rect 4779 1745 4791 5259
rect 4827 1745 4839 2835
rect 4851 1745 4863 4731
rect 4995 4337 5007 6939
rect 5019 4265 5031 6939
rect 4875 1745 4887 2811
rect 4971 1745 4983 4251
rect 5067 3881 5079 6939
rect 5091 3737 5103 6939
rect 5139 5393 5151 6939
rect 5187 4337 5199 6939
rect 5211 4073 5223 6939
rect 5235 5417 5247 6939
rect 5259 5465 5271 6939
rect 5307 5489 5319 6939
rect 4995 1745 5007 2787
rect 5019 1745 5031 3027
rect 5091 1745 5103 3723
rect 5115 1745 5127 3339
rect 5139 1745 5151 3027
rect 5187 1745 5199 2763
rect 5211 1745 5223 4059
rect 5235 1745 5247 3339
rect 5259 1745 5271 5427
rect 5331 3545 5343 6939
rect 5379 5513 5391 6939
rect 5427 5537 5439 6939
rect 5307 1745 5319 2739
rect 5355 1745 5367 2715
rect 5403 1745 5415 2691
rect 5451 1745 5463 5547
rect 5475 3617 5487 6939
rect 5547 5585 5559 6939
rect 5571 5633 5583 6939
rect 5595 5681 5607 6939
rect 5643 5729 5655 6939
rect 5667 5753 5679 6939
rect 5691 5777 5703 6939
rect 5475 1745 5487 3315
rect 5547 1745 5559 2667
rect 5571 1745 5583 5595
rect 5595 1745 5607 5643
rect 5643 1745 5655 5691
rect 5667 1745 5679 4299
rect 5691 3329 5703 5739
rect 5739 4529 5751 6939
rect 5763 5753 5775 6939
rect 5787 5825 5799 6939
rect 5739 1745 5751 2643
rect 5787 1745 5799 5787
rect 5811 1745 5823 4419
rect 5835 2633 5847 6939
rect 5859 3809 5871 6939
rect 5907 3809 5919 6939
rect 5955 5873 5967 6939
rect 5955 1745 5967 5835
rect 5979 3617 5991 6939
rect 6003 5897 6015 6939
rect 6051 5921 6063 6939
rect 6075 5537 6087 6939
rect 6099 2609 6111 6939
rect 6147 5945 6159 6939
rect 6171 5657 6183 6939
rect 6195 2585 6207 6939
rect 6219 5657 6231 6939
rect 6267 2657 6279 6939
rect 6291 5585 6303 6939
rect 6315 5969 6327 6939
rect 6363 5993 6375 6939
rect 6363 1745 6375 5571
rect 6387 4409 6399 6939
rect 6411 5585 6423 6939
rect 6459 6017 6471 6939
rect 6483 2825 6495 6939
rect 6507 3449 6519 6939
rect 6531 2561 6543 5739
rect 6555 3857 6567 6939
rect 6579 5753 6591 6939
rect 6507 1745 6519 2547
rect 6555 1745 6567 2523
rect 6579 1745 6591 4419
rect 6627 4145 6639 6939
rect 6675 6041 6687 6939
rect 6699 6065 6711 6939
rect 6723 6089 6735 6939
rect 6627 1745 6639 2547
rect 6675 1745 6687 3243
rect 6699 1745 6711 3075
rect 6723 2705 6735 6051
rect 6771 3545 6783 6939
rect 6795 6065 6807 6939
rect 6819 6113 6831 6939
rect 6867 6137 6879 6939
rect 6891 6065 6903 6939
rect 6747 1745 6759 2979
rect 6795 1745 6807 3939
rect 6819 1745 6831 4755
rect 6843 3521 6855 6051
rect 6867 1745 6879 5355
rect 6915 2993 6927 6939
rect 6963 5969 6975 6939
rect 6939 1745 6951 3219
rect 6963 1745 6975 2499
rect 6987 2489 6999 6939
rect 7011 5969 7023 6939
rect 7035 5849 7047 6939
rect 7083 5849 7095 6939
rect 7011 1745 7023 4923
rect 7035 1745 7047 5739
rect 7107 4817 7119 6939
rect 7131 6161 7143 6939
rect 7179 6185 7191 6939
rect 7131 1745 7143 4203
rect 7203 4049 7215 6939
rect 7227 6233 7239 6939
rect 7227 1745 7239 6195
rect 7251 4553 7263 6939
rect 7251 1745 7263 3315
rect 7275 1745 7287 6243
rect 7323 5921 7335 6939
rect 7347 5297 7359 6939
rect 7371 3689 7383 6939
rect 7395 6281 7407 6939
rect 7443 6305 7455 6939
rect 7395 2465 7407 5979
rect 7467 5417 7479 6939
rect 7515 4745 7527 6939
rect 7563 4889 7575 6939
rect 7323 1745 7335 2451
rect 7347 1745 7359 2427
rect 7371 1745 7383 2403
rect 7419 1745 7431 2931
rect 7443 1745 7455 4107
rect 7515 1745 7527 2451
rect 7563 1745 7575 2835
rect 7587 1745 7599 4827
rect 7611 4289 7623 6939
rect 7683 5993 7695 6939
rect 7707 4841 7719 6939
rect 7731 3953 7743 6939
rect 7635 1745 7647 2379
rect 7755 2369 7767 5379
rect 7779 4745 7791 6939
rect 7803 3785 7815 6939
rect 7827 6329 7839 6939
rect 7875 6353 7887 6939
rect 7899 6377 7911 6939
rect 7923 6401 7935 6939
rect 7971 6257 7983 6939
rect 7707 1745 7719 2355
rect 7755 1745 7767 2331
rect 7803 1745 7815 2355
rect 7827 1745 7839 5211
rect 7995 4769 8007 6939
rect 8019 6041 8031 6939
rect 7851 1745 7863 2307
rect 7875 1745 7887 2283
rect 7923 1745 7935 3315
rect 7947 1745 7959 4059
rect 7971 1745 7983 4755
rect 8043 1745 8055 6243
rect 8067 6041 8079 6939
rect 8067 1745 8079 5739
rect 8091 4769 8103 6939
rect 8115 2273 8127 6939
rect 8163 6425 8175 6939
rect 8139 1745 8151 3051
rect 8163 1745 8175 4131
rect 8187 3065 8199 6939
rect 8211 4649 8223 6939
rect 8235 2465 8247 6411
rect 8259 4649 8271 6939
rect 8283 5681 8295 6939
rect 8307 6425 8319 6939
rect 8331 6449 8343 6939
rect 8211 1745 8223 2235
rect 8259 1745 8271 4323
rect 8283 1745 8295 4299
rect 8331 1745 8343 5235
rect 8379 2993 8391 6939
rect 8403 4385 8415 6939
rect 8475 6497 8487 6939
rect 8403 1745 8415 2451
rect 8451 1745 8463 4371
rect 8475 1745 8487 6459
rect 8523 2225 8535 6939
rect 8547 6545 8559 6939
rect 8547 1745 8559 6507
rect 8571 4193 8583 6939
rect 8619 6305 8631 6939
rect 8667 5993 8679 6939
rect 8595 2201 8607 5811
rect 8571 1745 8583 2187
rect 8595 1745 8607 2163
rect 8643 1745 8655 4179
rect 8739 3929 8751 6939
rect 8763 4505 8775 6939
rect 8811 6569 8823 6939
rect 8691 1745 8703 2187
rect 8739 1745 8751 2139
rect 8787 1745 8799 5811
rect 8811 1745 8823 3339
rect 8835 1745 8847 6579
rect 8859 5921 8871 6939
rect 8883 4121 8895 6939
rect 8907 6617 8919 6939
rect 8955 6641 8967 6939
rect 8883 1745 8895 2115
rect 8907 1745 8919 4419
rect 8931 2129 8943 6291
rect 8955 4385 8967 6603
rect 8979 2129 8991 6939
rect 9003 5873 9015 6939
rect 9051 5873 9063 6939
rect 9075 5417 9087 6939
rect 8955 1745 8967 2091
rect 9003 1745 9015 5139
rect 9051 1745 9063 3723
rect 9099 2753 9111 6939
rect 9147 6617 9159 6939
rect 9171 6665 9183 6939
rect 9075 1745 9087 2067
rect 9123 1745 9135 4059
rect 9147 1745 9159 3195
rect 9171 2561 9183 5859
rect 9219 5201 9231 6939
rect 9243 1745 9255 4803
rect 9267 3089 9279 6939
rect 9291 2729 9303 6939
rect 9315 5873 9327 6939
rect 9363 3785 9375 6939
rect 9411 6689 9423 6939
rect 9267 1745 9279 2043
rect 9315 1745 9327 3771
rect 9387 1745 9399 2019
rect 9411 1745 9423 5043
rect 9435 3857 9447 6939
rect 9459 3905 9471 6939
rect 9459 1745 9471 1995
rect 9483 1745 9495 6123
rect 9507 4769 9519 6939
rect 9507 1745 9519 3123
rect 9531 2945 9543 6675
rect 9555 4817 9567 6939
rect 9627 5057 9639 6939
rect 9651 3593 9663 6939
rect 9675 6689 9687 6939
rect 9675 1745 9687 5139
rect 9699 1745 9711 4707
rect 9723 3137 9735 6939
rect 9747 5441 9759 6939
rect 9771 2417 9783 6939
rect 9795 2681 9807 6939
rect 9843 4385 9855 6939
rect 9867 3857 9879 6939
rect 9891 3065 9903 6939
rect 9939 4841 9951 6939
rect 9963 3593 9975 6939
rect 9987 3353 9999 6939
rect 10011 4385 10023 6939
rect 10059 6425 10071 6939
rect 10083 4505 10095 6939
rect 10107 6713 10119 6939
rect 10155 5681 10167 6939
rect 9771 1745 9783 1971
rect 9867 1745 9879 2403
rect 9891 1745 9903 2691
rect 9963 1745 9975 3051
rect 10107 1745 10119 5427
rect 10179 4649 10191 6939
rect 10203 5681 10215 6939
rect 10155 1745 10167 2619
rect 10203 1745 10215 4275
rect 10227 1745 10239 4131
rect 10251 2633 10263 6939
rect 10299 3185 10311 6939
rect 10323 5417 10335 6939
rect 10347 6737 10359 6939
rect 10395 6761 10407 6939
rect 10419 3977 10431 6939
rect 10443 2849 10455 6939
rect 10467 1961 10479 6939
rect 10515 1937 10527 6939
rect 10539 2945 10551 6939
rect 10563 6785 10575 6939
rect 10563 1913 10575 5835
rect 10611 5369 10623 6939
rect 10635 2057 10647 6939
rect 10659 2369 10671 6939
rect 10539 1745 10551 1899
rect 10563 1745 10575 1875
rect 10611 1745 10623 1899
rect 10683 1745 10695 5571
rect 10707 2369 10719 6939
rect 10731 3089 10743 6939
rect 10755 5585 10767 6939
rect 10803 6809 10815 6939
rect 10851 6233 10863 6939
rect 10779 1865 10791 6219
rect 10923 4673 10935 6939
rect 10947 5921 10959 6939
rect 10971 6377 10983 6939
rect 10731 1745 10743 1851
rect 10803 1745 10815 3075
rect 10827 1745 10839 3915
rect 10875 1745 10887 2931
rect 10899 1745 10911 1851
rect 10971 1745 10983 1827
rect 10995 1745 11007 3939
rect 11019 3929 11031 6939
rect 11043 3857 11055 6939
rect 11067 1745 11079 6531
rect 11091 4217 11103 6939
rect 11139 5153 11151 6939
rect 11163 4289 11175 6939
rect 11091 1745 11103 4155
rect 11187 1745 11199 4923
rect 11211 3377 11223 6939
rect 11235 1745 11247 6531
rect 11259 1889 11271 6939
rect 11283 6377 11295 6939
rect 11283 1745 11295 4275
rect 11307 4169 11319 6939
rect 11331 3329 11343 6363
rect 11355 5513 11367 6939
rect 11379 6377 11391 6939
rect 11307 1745 11319 2931
rect 11355 1745 11367 3939
rect 11403 3305 11415 6939
rect 11427 6833 11439 6939
rect 11427 2537 11439 4155
rect 11451 1745 11463 6219
rect 11475 3521 11487 6939
rect 11523 5489 11535 6939
rect 11475 1745 11487 1803
rect 11499 1745 11511 2619
rect 11547 1745 11559 3891
rect 11571 1745 11583 4155
rect 11595 2681 11607 6939
rect 11643 6233 11655 6939
rect 11691 6857 11703 6939
rect 11619 1745 11631 5739
rect 11643 1745 11655 2619
rect 11667 1817 11679 5235
rect 11691 1745 11703 6699
rect 11715 4265 11727 6939
rect 11739 5249 11751 6939
rect 11763 5321 11775 6939
rect 11811 6449 11823 6939
rect 11835 6833 11847 6939
rect 11859 5321 11871 6939
rect 11883 5273 11895 6939
rect 11907 6449 11919 6939
rect 11955 6161 11967 6939
rect 11979 5273 11991 6939
rect 12003 6713 12015 6939
rect 12027 6833 12039 6939
rect 12051 6881 12063 6939
rect 12099 6905 12111 6939
rect 12123 6929 12135 6939
rect 11715 1745 11727 1803
rect 11739 1745 11751 1779
rect 11787 1745 11799 4251
rect 11811 1745 11823 2835
rect 11907 1745 11919 3075
rect 11931 1745 11943 1803
rect 12003 1745 12015 5979
rect 12027 1745 12039 4419
rect 12051 1745 12063 4035
rect 12075 1817 12087 5403
rect 12147 4601 12159 6939
rect 12099 1745 12111 2403
rect 12123 1745 12135 4443
rect 12171 2009 12183 6435
rect 12195 1745 12207 3891
rect 12219 1745 12231 4923
rect 12255 2537 12267 6819
rect 12315 4457 12327 6939
rect 12339 2417 12351 6915
rect 12363 6137 12375 6939
rect 12435 4601 12447 6939
rect 12459 3089 12471 6939
rect 12483 6449 12495 6939
rect 12531 6833 12543 6939
rect 12579 5801 12591 6939
rect 12651 5801 12663 6939
rect 12675 5201 12687 6939
rect 12699 5345 12711 6939
rect 12723 3881 12735 6939
rect 12795 3977 12807 6939
rect 12819 4721 12831 6939
rect 12867 4265 12879 6939
rect 12915 6809 12927 6939
rect 12939 3329 12951 6939
rect 12243 1745 12255 1995
rect 12963 1985 12975 6939
rect 13011 4505 13023 6939
rect 13035 4337 13047 6939
rect 13059 3377 13071 6939
rect 13083 3689 13095 6939
rect 13107 4961 13119 6939
rect 13155 4145 13167 6939
rect 12291 1745 12303 1803
rect 13059 1745 13071 1971
rect 13107 1745 13119 4083
rect 13179 3929 13191 6939
rect 13203 4961 13215 6939
rect 13251 5201 13263 6939
rect 13275 5345 13287 6939
rect 13299 5009 13311 6939
rect 13131 1745 13143 2403
rect 13203 1745 13215 2811
rect 13227 1745 13239 4923
rect 13251 1745 13263 3291
rect 13323 1985 13335 6027
rect 13347 3425 13359 6939
rect 13371 5297 13383 6939
rect 13395 5009 13407 6939
rect 13515 5201 13527 6939
rect 13347 1745 13359 1755
rect 13371 1745 13383 1971
rect 13395 1745 13407 2595
rect 13419 1745 13431 3651
rect 13443 2105 13455 5187
rect 13491 1745 13503 2403
rect 13515 1745 13527 4107
rect 13539 1745 13551 3843
rect 13563 1745 13575 5787
rect 13587 2177 13599 5187
rect 13635 1745 13647 3075
rect 13659 1745 13671 3651
rect 13707 1745 13719 5091
rect 13827 1745 13839 6123
rect 13875 5633 13887 6939
rect 13923 5105 13935 6939
rect 13851 1745 13863 4707
rect 13875 1745 13887 2595
rect 13923 1745 13935 2163
rect 13947 1745 13959 6555
rect 13995 1745 14007 4155
rect 14043 1745 14055 4515
rect 14067 2657 14079 6939
rect 14115 5945 14127 6939
rect 14235 4625 14247 6939
rect 14091 1745 14103 2571
rect 14139 1745 14151 2595
rect 14187 1745 14199 2571
rect 14235 1745 14247 1875
rect 14259 1745 14271 3579
rect 14283 1745 14295 4827
rect 14355 1745 14367 2091
rect 14379 1745 14391 4611
rect 14403 1745 14415 3123
rect 14451 1745 14463 6771
rect 14595 4937 14607 6939
rect 14475 1745 14487 4659
rect 14619 4577 14631 5235
rect 14643 5201 14655 6939
rect 14499 1745 14511 4563
rect 14547 1745 14559 3123
rect 14571 1745 14583 3723
rect 14595 1745 14607 4563
rect 14643 1745 14655 3579
rect 14667 1745 14679 5403
rect 14691 1745 14703 2763
rect 14715 2417 14727 5187
rect 14739 1745 14751 3531
rect 14763 1745 14775 3507
rect 14787 2585 14799 6939
rect 14835 6161 14847 6939
rect 14883 4577 14895 6939
rect 14811 1745 14823 2811
rect 14859 1745 14871 4059
rect 14883 1745 14895 3219
rect 14907 1745 14919 3507
rect 14955 3161 14967 6939
rect 14979 3401 14991 6939
rect 15075 2081 15087 6939
rect 15099 2993 15111 6939
rect 15123 4553 15135 6939
rect 15195 5945 15207 6939
rect 15219 6017 15231 6939
rect 15027 1745 15039 1923
rect 15099 1745 15111 2571
rect 15195 1745 15207 5763
rect 15315 5201 15327 6939
rect 15219 1745 15231 3723
rect 15291 1745 15303 2979
rect 15315 1745 15327 3603
rect 15339 3377 15351 6939
rect 15363 3353 15375 6939
rect 15387 6857 15399 6939
rect 15339 1745 15351 1875
rect 15363 1745 15375 3003
rect 15411 1745 15423 4995
rect 15435 4937 15447 6939
rect 15459 5009 15471 6939
rect 15483 5705 15495 6939
rect 15531 5249 15543 6939
rect 15555 5201 15567 6939
rect 15435 1745 15447 3483
rect 15483 1745 15495 3483
rect 15507 3281 15519 5187
rect 15579 3497 15591 6483
rect 15531 1745 15543 2235
rect 15555 1745 15567 2931
rect 15603 2177 15615 6939
rect 15651 4049 15663 6939
rect 15675 5633 15687 6939
rect 15699 5705 15711 6939
rect 15747 3353 15759 6939
rect 15627 1745 15639 2403
rect 15651 1745 15663 2715
rect 15675 1745 15687 2115
rect 15723 1745 15735 3123
rect 15747 1745 15759 3003
rect 15771 2417 15783 5187
rect 15795 3185 15807 6939
rect 15819 3017 15831 4323
rect 15843 1745 15855 4131
rect 15867 2513 15879 6939
rect 15891 4817 15903 6939
rect 15915 5201 15927 6939
rect 15939 1745 15951 4443
rect 15963 2345 15975 6939
rect 15987 5801 15999 6939
rect 16011 5777 16023 6939
rect 15963 1745 15975 2163
rect 16011 1745 16023 4035
rect 16035 2177 16047 6747
rect 16059 6041 16071 6939
rect 16083 6593 16095 6939
rect 16107 5561 16119 6939
rect 16155 6545 16167 6939
rect 16179 5753 16191 6939
rect 16059 1745 16071 3315
rect 16083 1745 16095 3483
rect 16107 1745 16119 4731
rect 16131 1745 16143 4755
rect 16203 1745 16215 5907
rect 16227 3833 16239 6939
rect 16275 5465 16287 6939
rect 16299 4793 16311 6939
rect 16323 5465 16335 6939
rect 16227 1745 16239 3723
rect 16251 1745 16263 3363
rect 16299 1745 16311 3411
rect 16347 2417 16359 6027
rect 16371 3497 16383 6747
rect 16395 3377 16407 6939
rect 16419 4793 16431 6939
rect 16443 5897 16455 6939
rect 16467 5561 16479 6939
rect 16491 5897 16503 6939
rect 16539 6449 16551 6939
rect 16563 6041 16575 6939
rect 16419 1745 16431 4491
rect 16443 1745 16455 4203
rect 16467 1745 16479 3939
rect 16491 1745 16503 2043
rect 16515 1745 16527 3483
rect 16563 1745 16575 2667
rect 16587 2417 16599 6939
rect 16611 6137 16623 6939
rect 16587 1745 16599 2163
rect 16611 1745 16623 2475
rect 16635 1817 16647 6123
rect 16731 5657 16743 6939
rect 17283 5657 17295 6939
rect 17331 6137 17343 6939
rect 17355 4673 17367 6939
rect 17403 6449 17415 6939
rect 17283 1745 17295 3075
rect 17307 1745 17319 4419
rect 17379 1745 17391 4803
rect 17403 1745 17415 5403
rect 17427 1745 17439 3411
rect 17451 1865 17463 6939
rect 17475 3665 17487 6939
rect 17499 3041 17511 6939
rect 17523 3065 17535 6939
rect 17523 1745 17535 3003
rect 17547 2177 17559 5643
rect 17571 4385 17583 6939
rect 17595 2753 17607 6939
rect 17619 4865 17631 6939
rect 17643 4985 17655 6939
rect 17691 6473 17703 6939
rect 17739 6065 17751 6939
rect 17595 1745 17607 2715
rect 17619 1745 17631 3915
rect 17655 2729 17667 3123
rect 17691 1745 17703 4059
rect 17715 1745 17727 1899
rect 17739 1745 17751 4443
rect 17763 2945 17775 6939
rect 17787 4457 17799 6939
rect 17811 4601 17823 6939
rect 17787 1745 17799 4419
rect 17823 2393 17835 4443
rect 17859 2681 17871 6939
rect 17907 6521 17919 6939
rect 17883 3017 17895 5931
rect 17955 3353 17967 6939
rect 17979 3329 17991 6939
rect 17931 1745 17943 2547
rect 18003 1745 18015 3315
rect 18027 2057 18039 6939
rect 18075 5753 18087 6939
rect 18051 1745 18063 3579
rect 18099 3089 18111 6939
rect 18123 5537 18135 6939
rect 18171 4385 18183 6939
rect 18195 4937 18207 6939
rect 18219 4841 18231 6939
rect 18243 4913 18255 6939
rect 18291 5369 18303 6939
rect 18123 1745 18135 4275
rect 18147 1745 18159 3171
rect 18171 1745 18183 3459
rect 18219 1745 18231 3147
rect 18267 1745 18279 5043
rect 18303 2057 18315 4371
rect 18339 4193 18351 6939
rect 18411 5513 18423 6939
rect 18339 1745 18351 3603
rect 18363 1745 18375 3915
rect 18411 1745 18423 4659
rect 18435 3305 18447 6939
rect 18483 4385 18495 6939
rect 18459 1745 18471 3651
rect 18507 1745 18519 4323
rect 18531 4121 18543 6939
rect 18555 5921 18567 6939
rect 18579 3857 18591 6939
rect 18603 4553 18615 6939
rect 18579 1745 18591 3603
rect 18603 1745 18615 4323
rect 18627 3617 18639 5211
rect 18651 2777 18663 6939
rect 18675 3425 18687 6939
rect 18699 4433 18711 6939
rect 18723 4409 18735 6939
rect 18651 1745 18663 2187
rect 18699 1745 18711 3627
rect 18723 1745 18735 3603
rect 18747 1745 18759 4779
rect 18771 2009 18783 6939
rect 18819 4001 18831 6939
rect 18855 3617 18867 5739
rect 18891 4409 18903 6939
rect 18795 1745 18807 2403
rect 18843 1745 18855 3099
rect 18891 1745 18903 4395
rect 18915 3473 18927 6939
rect 18939 6137 18951 6939
rect 18987 5489 18999 6939
rect 19011 4769 19023 6939
rect 19035 5825 19047 6939
rect 18951 2033 18963 4419
rect 19047 4001 19059 5715
rect 19083 4433 19095 6939
rect 19011 1745 19023 3987
rect 19035 1745 19047 3075
rect 19083 1745 19095 3555
rect 19107 3329 19119 6939
rect 19131 3665 19143 6939
rect 19179 5753 19191 6939
rect 19155 3185 19167 4419
rect 19203 2993 19215 6939
rect 19227 6209 19239 6939
rect 19275 5201 19287 6939
rect 19299 6737 19311 6939
rect 19203 1745 19215 2739
rect 19323 2441 19335 6939
rect 19371 4169 19383 6939
rect 19419 6257 19431 6939
rect 19491 2513 19503 6939
rect 19539 4841 19551 6939
rect 19611 2033 19623 6939
rect 19635 3233 19647 6939
rect 19683 5441 19695 6939
rect 19731 4529 19743 6939
rect 19755 1745 19767 6939
rect 19779 5969 19791 6939
rect 19827 4433 19839 6939
rect 19803 1745 19815 3915
rect 19827 1745 19839 4131
rect 19851 1745 19863 3579
rect 19875 3257 19887 6939
rect 19899 2033 19911 4419
rect 19923 1745 19935 4923
rect 19947 3425 19959 6939
rect 19971 4913 19983 6939
rect 19995 5345 20007 6939
rect 19971 1745 19983 4875
rect 20043 4601 20055 6939
rect 20067 6233 20079 6939
rect 20019 1745 20031 2091
rect 20043 1745 20055 4563
rect 20067 1745 20079 5451
rect 20091 4433 20103 6939
rect 20115 4457 20127 6939
rect 20115 1745 20127 2355
rect 20139 1745 20151 5283
rect 20163 3737 20175 6939
rect 20187 3137 20199 6939
rect 20211 3665 20223 6939
rect 20235 4553 20247 6939
rect 20235 1745 20247 3171
rect 20259 1745 20271 4755
rect 20283 3761 20295 6939
rect 20307 2777 20319 4899
rect 20331 2753 20343 6939
rect 20475 6929 20487 6939
rect 20283 1745 20295 2019
rect 20331 1745 20343 2379
rect 20355 1745 20367 4299
rect 20379 1745 20391 2811
rect 20403 1745 20415 6603
rect 20451 1745 20463 4059
rect 20475 1745 20487 6867
rect 20499 4457 20511 6915
rect 20835 6377 20847 6939
rect 20547 1745 20559 3339
rect 20571 1745 20583 4803
rect 20595 1745 20607 5403
rect 20619 1745 20631 5259
rect 20667 1745 20679 3915
rect 20691 1745 20703 5739
rect 20715 1745 20727 4083
rect 20763 1745 20775 4155
rect 20787 1745 20799 3867
rect 20811 1745 20823 4083
rect 20859 1745 20871 4995
rect 20883 2873 20895 6939
rect 21027 6545 21039 6939
rect 21075 5921 21087 6939
rect 20907 2753 20919 2979
rect 20883 1745 20895 2739
rect 21003 1745 21015 2259
rect 21075 1745 21087 4059
rect 21123 1745 21135 6267
rect 21147 4265 21159 6939
rect 21171 2057 21183 6939
rect 21195 4457 21207 6939
rect 21243 3953 21255 6939
rect 21267 4145 21279 6939
rect 21291 4001 21303 5787
rect 21207 1937 21219 3771
rect 21171 1745 21183 1923
rect 21243 1745 21255 1947
rect 21267 1745 21279 3987
rect 21315 3137 21327 6939
rect 21363 3089 21375 6939
rect 21387 3953 21399 6939
rect 21411 3353 21423 6939
rect 21363 1745 21375 3051
rect 21411 1745 21423 2907
rect 21435 1769 21447 6939
rect 21483 6785 21495 6939
rect 21531 6641 21543 6939
rect 21459 1745 21471 5091
rect 21507 1745 21519 4635
rect 21555 1745 21567 4347
rect 21579 1745 21591 4467
rect 21603 4145 21615 6939
rect 21627 6017 21639 6939
rect 21651 2945 21663 6939
rect 21675 6665 21687 6939
rect 21627 1745 21639 2307
rect 21675 1745 21687 2643
rect 21699 1745 21711 5091
rect 21723 4097 21735 6939
rect 21747 3065 21759 5379
rect 21771 4313 21783 6939
rect 21795 4361 21807 6939
rect 21819 4481 21831 6939
rect 21843 4265 21855 5403
rect 21771 1745 21783 4251
rect 21867 4241 21879 6939
rect 21891 4505 21903 6939
rect 21939 6761 21951 6939
rect 21951 4265 21963 5571
rect 21987 5489 21999 6939
rect 21819 1745 21831 3219
rect 21891 1745 21903 4251
rect 21915 1745 21927 3699
rect 22011 3545 22023 6939
rect 22059 6425 22071 6939
rect 22107 6089 22119 6939
rect 21987 1745 21999 2667
rect 22107 1745 22119 5139
rect 22131 2945 22143 6939
rect 22155 4025 22167 6939
rect 22203 4721 22215 6939
rect 22131 1745 22143 2907
rect 22155 1745 22167 3291
rect 22179 2921 22191 4347
rect 22227 2825 22239 6939
rect 22275 6857 22287 6939
rect 22251 2753 22263 4179
rect 22227 1745 22239 2739
rect 22275 1745 22287 6795
rect 22299 2993 22311 6843
rect 22323 4577 22335 6939
rect 22323 1745 22335 4515
rect 22347 3833 22359 6939
rect 22371 1745 22383 4419
rect 22395 3713 22407 6939
rect 22443 4697 22455 6939
rect 22419 2249 22431 4563
rect 22443 1745 22455 4251
rect 22467 2945 22479 6939
rect 22491 6353 22503 6939
rect 22539 4313 22551 6939
rect 22467 1745 22479 2355
rect 22515 1745 22527 1851
rect 22539 1745 22551 3795
rect 22563 2417 22575 6939
rect 22587 6305 22599 6939
rect 22635 4361 22647 6939
rect 22659 4505 22671 6939
rect 22683 4793 22695 6939
rect 22587 1745 22599 3891
rect 22611 1745 22623 4299
rect 22659 1745 22671 2979
rect 22683 1745 22695 4755
rect 22707 4265 22719 6531
rect 22731 3209 22743 6939
rect 22755 1913 22767 6939
rect 22803 6833 22815 6939
rect 22755 1745 22767 1851
rect 22779 1745 22791 4371
rect 22827 1745 22839 5307
rect 22851 2537 22863 6939
rect 22875 1745 22887 5043
rect 22899 4385 22911 6939
rect 22971 6137 22983 6939
rect 22923 4409 22935 4779
rect 22899 1745 22911 3387
rect 22923 2849 22935 4371
rect 22971 1745 22983 6099
rect 23019 5081 23031 6939
rect 22995 1745 23007 3291
rect 23043 1745 23055 4707
rect 23067 4073 23079 6123
rect 23091 2057 23103 6939
rect 23115 4937 23127 6939
rect 23139 4529 23151 6939
rect 23163 4841 23175 6939
rect 23091 1745 23103 1947
rect 23115 1745 23127 2331
rect 23139 1745 23151 4467
rect 23187 1985 23199 6939
rect 23235 4937 23247 6939
rect 23211 1745 23223 4107
rect 23235 1745 23247 3891
rect 23259 2393 23271 6939
rect 23283 1745 23295 6027
rect 23307 6017 23319 6939
rect 23355 4985 23367 6939
rect 23403 5849 23415 6939
rect 23475 6761 23487 6939
rect 23331 1745 23343 4203
rect 23355 1745 23367 4923
rect 23379 1745 23391 5547
rect 23439 2777 23451 4971
rect 23427 1745 23439 2547
rect 23475 1745 23487 4995
rect 23499 4745 23511 6939
rect 23523 2849 23535 6939
rect 23547 2465 23559 6939
rect 23571 1745 23583 4947
rect 23595 2153 23607 6939
rect 23619 4049 23631 6939
rect 23667 4169 23679 6939
rect 23715 3857 23727 6939
rect 23739 5129 23751 6939
rect 23787 5249 23799 6939
rect 23835 4937 23847 6939
rect 23595 1745 23607 2115
rect 23643 1745 23655 3267
rect 23691 1745 23703 3387
rect 23763 1745 23775 4851
rect 23799 2129 23811 4515
rect 23859 3737 23871 6939
rect 23883 5153 23895 6939
rect 23907 3689 23919 6939
rect 23931 6185 23943 6939
rect 23979 5681 23991 6939
rect 23883 1745 23895 2019
rect 23907 1745 23919 3651
rect 24003 2825 24015 6939
rect 23955 1745 23967 2691
rect 24027 1961 24039 5787
rect 24051 1865 24063 6939
rect 24075 1745 24087 6387
rect 24099 4769 24111 6939
rect 24123 3353 24135 6939
rect 24147 3665 24159 4827
rect 24171 1889 24183 6939
rect 24219 3449 24231 6939
rect 24267 4361 24279 6939
rect 24339 4553 24351 6939
rect 24363 4193 24375 6939
rect 24387 2201 24399 6939
rect 24411 3497 24423 6939
rect 24483 4457 24495 6939
rect 24507 5801 24519 6939
rect 24555 5225 24567 6939
rect 24483 1745 24495 2931
rect 24603 1793 24615 6939
rect 24627 4361 24639 6939
rect 24651 6713 24663 6939
rect 24627 1745 24639 3579
rect 24651 1745 24663 4275
rect 24675 1745 24687 3171
rect 24699 2609 24711 6939
rect 24699 1745 24711 2211
rect 24723 1889 24735 4347
rect 24747 1745 24759 6435
rect 24819 1769 24831 6939
rect 24843 3401 24855 6939
rect 24891 2585 24903 6939
rect 24939 5993 24951 6939
rect 24939 1745 24951 5883
rect 24963 3329 24975 6939
rect 24987 5633 24999 6939
rect 25035 2777 25047 6939
rect 25059 2033 25071 6939
rect 25083 4625 25095 6939
rect 25131 2825 25143 6939
rect 25155 3977 25167 6939
rect 25179 2057 25191 6939
rect 25203 4337 25215 6939
rect 25251 2657 25263 6939
rect 25275 2873 25287 6939
rect 25299 5825 25311 6939
rect 25347 5849 25359 6939
rect 25299 1745 25311 5715
rect 25323 4601 25335 5811
rect 25347 1745 25359 5739
rect 25371 5417 25383 6939
rect 25395 1841 25407 6939
rect 25419 5705 25431 5835
rect 25443 5513 25455 6939
rect 25467 4505 25479 6939
rect 25491 1745 25503 6675
rect 25515 6065 25527 6939
rect 25539 1745 25551 6315
rect 25563 6161 25575 6939
rect 25563 1745 25575 2955
rect 25587 2033 25599 6939
rect 25611 6065 25623 6939
rect 25611 1745 25623 6027
rect 25635 1745 25647 5859
rect 25659 2321 25671 6939
rect 25683 3521 25695 6939
rect 25707 5177 25719 6939
rect 25731 5801 25743 6939
rect 25755 5825 25767 6939
rect 25659 1745 25671 2259
rect 25707 1745 25719 4347
rect 25755 1745 25767 5763
rect 25779 2273 25791 6891
rect 25803 5993 25815 6939
rect 25827 6065 25839 6939
rect 25851 5033 25863 6939
rect 25875 4361 25887 5811
rect 25899 2009 25911 6939
rect 25923 3737 25935 6939
rect 25947 2801 25959 6939
rect 25995 5609 26007 6939
rect 26139 1745 26339 6939
rect 26451 4300 26521 4312
rect 26451 2884 26521 2896
rect 26451 2620 26521 2632
rect 26451 2284 26521 2296
rect 0 59 70 71
rect 0 35 70 47
rect 123 0 323 946
rect 339 0 351 946
rect 363 0 375 946
rect 387 0 399 946
rect 411 0 423 946
rect 1611 96 1623 946
rect 1635 120 1647 946
rect 1659 144 1671 946
rect 1707 48 1719 946
rect 1827 48 1839 946
rect 2427 168 2439 946
rect 2547 96 2559 946
rect 4131 96 4143 946
rect 4395 96 4407 946
rect 4419 192 4431 946
rect 4443 216 4455 946
rect 4491 240 4503 946
rect 4899 264 4911 946
rect 4947 288 4959 946
rect 5043 48 5055 946
rect 5331 48 5343 946
rect 5427 312 5439 946
rect 5499 336 5511 946
rect 5691 360 5703 946
rect 5715 96 5727 946
rect 5835 96 5847 946
rect 6315 384 6327 946
rect 6507 24 6519 946
rect 6723 408 6735 946
rect 6915 408 6927 946
rect 7083 432 7095 946
rect 7155 168 7167 946
rect 7179 288 7191 946
rect 7467 288 7479 946
rect 7491 168 7503 946
rect 7683 480 7695 946
rect 7995 504 8007 946
rect 8091 528 8103 946
rect 8307 552 8319 946
rect 8379 576 8391 946
rect 8427 600 8439 946
rect 8523 624 8535 946
rect 8667 648 8679 946
rect 8715 672 8727 946
rect 9027 696 9039 946
rect 9195 720 9207 946
rect 7671 0 7683 442
rect 9363 144 9375 946
rect 9555 144 9567 946
rect 9579 96 9591 946
rect 9627 360 9639 946
rect 9723 360 9735 946
rect 9795 96 9807 946
rect 9819 744 9831 946
rect 9915 768 9927 946
rect 10011 792 10023 946
rect 10083 816 10095 946
rect 10251 840 10263 946
rect 10299 864 10311 946
rect 10347 192 10359 946
rect 10419 192 10431 946
rect 10443 888 10455 946
rect 10491 288 10503 946
rect 10659 288 10671 946
rect 11019 240 11031 946
rect 11139 240 11151 946
rect 11211 912 11223 946
rect 11403 936 11415 946
rect 11427 264 11439 946
rect 11595 792 11607 946
rect 11859 480 11871 946
rect 11955 480 11967 946
rect 12147 192 12159 946
rect 12339 792 12351 946
rect 12867 168 12879 946
rect 13011 264 13023 946
rect 13035 480 13047 946
rect 13155 480 13167 946
rect 13275 192 13287 946
rect 13323 840 13335 946
rect 13467 912 13479 946
rect 13611 336 13623 946
rect 13755 840 13767 946
rect 14067 336 14079 946
rect 14163 336 14175 946
rect 13779 0 13791 322
rect 14307 48 14319 946
rect 14955 168 14967 946
rect 14979 768 14991 946
rect 15003 888 15015 946
rect 15075 720 15087 946
rect 15147 648 15159 946
rect 15243 264 15255 946
rect 15459 648 15471 946
rect 15579 672 15591 946
rect 15771 96 15783 946
rect 15819 432 15831 946
rect 15891 816 15903 946
rect 16155 288 16167 946
rect 16347 672 16359 946
rect 16731 720 16743 946
rect 17139 888 17151 946
rect 17331 120 17343 946
rect 17475 360 17487 946
rect 17643 768 17655 946
rect 17835 408 17847 946
rect 17907 192 17919 946
rect 17955 144 17967 946
rect 18819 216 18831 946
rect 18939 696 18951 946
rect 19611 720 19623 946
rect 19755 696 19767 946
rect 19875 696 19887 946
rect 19768 682 19786 696
rect 19767 0 19779 682
rect 19947 552 19959 946
rect 20187 720 20199 946
rect 20499 936 20511 946
rect 20931 864 20943 946
rect 20979 696 20991 946
rect 21027 528 21039 946
rect 21051 480 21063 946
rect 21291 792 21303 946
rect 21339 744 21351 946
rect 21483 384 21495 946
rect 21723 624 21735 946
rect 21939 72 21951 946
rect 22035 600 22047 946
rect 22179 648 22191 946
rect 22251 768 22263 946
rect 22347 456 22359 946
rect 22419 672 22431 946
rect 22563 840 22575 946
rect 22707 312 22719 946
rect 22923 336 22935 946
rect 23163 480 23175 946
rect 23547 360 23559 946
rect 23811 552 23823 946
rect 24435 912 24447 946
rect 24771 240 24783 946
rect 24819 576 24831 946
rect 25515 504 25527 946
rect 25707 504 25719 946
rect 25755 528 25767 946
rect 25755 48 25767 466
rect 25779 24 25791 706
rect 25803 72 25815 514
rect 19899 0 19911 10
rect 26139 0 26339 946
rect 26451 491 26521 503
rect 26451 59 26521 71
rect 26451 35 26521 47
rect 26451 11 26521 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 6939
box 0 0 1464 799
use nor2 g8525
timestamp 1386235306
transform 1 0 1587 0 1 6939
box 0 0 120 799
use and2 g8528
timestamp 1386234845
transform 1 0 1707 0 1 6939
box 0 0 120 799
use nand2 g8561
timestamp 1386234792
transform 1 0 1827 0 1 6939
box 0 0 96 799
use nand2 g8448
timestamp 1386234792
transform 1 0 1923 0 1 6939
box 0 0 96 799
use inv g8291
timestamp 1386238110
transform 1 0 2019 0 1 6939
box 0 0 120 799
use nand3 g8445
timestamp 1386234893
transform 1 0 2139 0 1 6939
box 0 0 120 799
use inv g8606
timestamp 1386238110
transform 1 0 2259 0 1 6939
box 0 0 120 799
use inv g8576
timestamp 1386238110
transform 1 0 2379 0 1 6939
box 0 0 120 799
use nor2 g8369
timestamp 1386235306
transform 1 0 2499 0 1 6939
box 0 0 120 799
use nand2 g8541
timestamp 1386234792
transform 1 0 2619 0 1 6939
box 0 0 96 799
use inv g8462
timestamp 1386238110
transform 1 0 2715 0 1 6939
box 0 0 120 799
use nand3 g8469
timestamp 1386234893
transform 1 0 2835 0 1 6939
box 0 0 120 799
use nor2 g8370
timestamp 1386235306
transform 1 0 2955 0 1 6939
box 0 0 120 799
use nor2 g8513
timestamp 1386235306
transform 1 0 3075 0 1 6939
box 0 0 120 799
use inv g8313
timestamp 1386238110
transform 1 0 3195 0 1 6939
box 0 0 120 799
use nand2 g8344
timestamp 1386234792
transform 1 0 3315 0 1 6939
box 0 0 96 799
use nand2 g8314
timestamp 1386234792
transform 1 0 3411 0 1 6939
box 0 0 96 799
use nand2 g8327
timestamp 1386234792
transform 1 0 3507 0 1 6939
box 0 0 96 799
use nand4 g8545
timestamp 1386234936
transform 1 0 3603 0 1 6939
box 0 0 144 799
use nand2 g8477
timestamp 1386234792
transform 1 0 3747 0 1 6939
box 0 0 96 799
use nand2 g8554
timestamp 1386234792
transform 1 0 3843 0 1 6939
box 0 0 96 799
use nand2 g8295
timestamp 1386234792
transform 1 0 3939 0 1 6939
box 0 0 96 799
use nand4 g8287
timestamp 1386234936
transform 1 0 4035 0 1 6939
box 0 0 144 799
use nand4 g8506
timestamp 1386234936
transform 1 0 4179 0 1 6939
box 0 0 144 799
use and2 g8276
timestamp 1386234845
transform 1 0 4323 0 1 6939
box 0 0 120 799
use nor2 g8261
timestamp 1386235306
transform 1 0 4443 0 1 6939
box 0 0 120 799
use nand4 g8567
timestamp 1386234936
transform 1 0 4563 0 1 6939
box 0 0 144 799
use and2 g8318
timestamp 1386234845
transform 1 0 4707 0 1 6939
box 0 0 120 799
use inv g8377
timestamp 1386238110
transform 1 0 4827 0 1 6939
box 0 0 120 799
use nand2 g8474
timestamp 1386234792
transform 1 0 4947 0 1 6939
box 0 0 96 799
use nor2 g8390
timestamp 1386235306
transform 1 0 5043 0 1 6939
box 0 0 120 799
use nand3 g8585
timestamp 1386234893
transform 1 0 5163 0 1 6939
box 0 0 120 799
use nor2 g8603
timestamp 1386235306
transform 1 0 5283 0 1 6939
box 0 0 120 799
use inv g8584
timestamp 1386238110
transform 1 0 5403 0 1 6939
box 0 0 120 799
use nand2 g8597
timestamp 1386234792
transform 1 0 5523 0 1 6939
box 0 0 96 799
use nand2 g8333
timestamp 1386234792
transform 1 0 5619 0 1 6939
box 0 0 96 799
use nand2 g8472
timestamp 1386234792
transform 1 0 5715 0 1 6939
box 0 0 96 799
use nor2 g8338
timestamp 1386235306
transform 1 0 5811 0 1 6939
box 0 0 120 799
use nand2 g8572
timestamp 1386234792
transform 1 0 5931 0 1 6939
box 0 0 96 799
use nand2 g8280
timestamp 1386234792
transform 1 0 6027 0 1 6939
box 0 0 96 799
use nand3 g8310
timestamp 1386234893
transform 1 0 6123 0 1 6939
box 0 0 120 799
use nand2 g8450
timestamp 1386234792
transform 1 0 6243 0 1 6939
box 0 0 96 799
use nand2 g8456
timestamp 1386234792
transform 1 0 6339 0 1 6939
box 0 0 96 799
use nand2 g8589
timestamp 1386234792
transform 1 0 6435 0 1 6939
box 0 0 96 799
use nor2 g8362
timestamp 1386235306
transform 1 0 6531 0 1 6939
box 0 0 120 799
use nand2 g8616
timestamp 1386234792
transform 1 0 6651 0 1 6939
box 0 0 96 799
use nand2 g8366
timestamp 1386234792
transform 1 0 6747 0 1 6939
box 0 0 96 799
use nand2 g8281
timestamp 1386234792
transform 1 0 6843 0 1 6939
box 0 0 96 799
use nand3 g8547
timestamp 1386234893
transform 1 0 6939 0 1 6939
box 0 0 120 799
use nand2 g8269
timestamp 1386234792
transform 1 0 7059 0 1 6939
box 0 0 96 799
use nand4 g8493
timestamp 1386234936
transform 1 0 7155 0 1 6939
box 0 0 144 799
use nand3 g8440
timestamp 1386234893
transform 1 0 7299 0 1 6939
box 0 0 120 799
use nor2 g8504
timestamp 1386235306
transform 1 0 7419 0 1 6939
box 0 0 120 799
use inv g8449
timestamp 1386238110
transform 1 0 7539 0 1 6939
box 0 0 120 799
use nand2 g8414
timestamp 1386234792
transform 1 0 7659 0 1 6939
box 0 0 96 799
use nand2 g8275
timestamp 1386234792
transform 1 0 7755 0 1 6939
box 0 0 96 799
use nand2 g8418
timestamp 1386234792
transform 1 0 7851 0 1 6939
box 0 0 96 799
use nand2 g8483
timestamp 1386234792
transform 1 0 7947 0 1 6939
box 0 0 96 799
use nand2 g8290
timestamp 1386234792
transform 1 0 8043 0 1 6939
box 0 0 96 799
use nand2 g8511
timestamp 1386234792
transform 1 0 8139 0 1 6939
box 0 0 96 799
use nand3 g8334
timestamp 1386234893
transform 1 0 8235 0 1 6939
box 0 0 120 799
use nand2 g8407
timestamp 1386234792
transform 1 0 8355 0 1 6939
box 0 0 96 799
use rowcrosser AluEn
timestamp 1386086759
transform 1 0 8451 0 1 6939
box 0 0 48 799
use nand2 g8486
timestamp 1386234792
transform 1 0 8499 0 1 6939
box 0 0 96 799
use inv g8618
timestamp 1386238110
transform 1 0 8595 0 1 6939
box 0 0 120 799
use nor2 g8562
timestamp 1386235306
transform 1 0 8715 0 1 6939
box 0 0 120 799
use nand2 g8363
timestamp 1386234792
transform 1 0 8835 0 1 6939
box 0 0 96 799
use nand2 g8489
timestamp 1386234792
transform 1 0 8931 0 1 6939
box 0 0 96 799
use nand2 g8381
timestamp 1386234792
transform 1 0 9027 0 1 6939
box 0 0 96 799
use and2 g8403
timestamp 1386234845
transform 1 0 9123 0 1 6939
box 0 0 120 799
use nand2 g8612
timestamp 1386234792
transform 1 0 9243 0 1 6939
box 0 0 96 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 9339 0 1 6939
box 0 0 48 799
use nand2 g8631
timestamp 1386234792
transform 1 0 9387 0 1 6939
box 0 0 96 799
use inv g8357
timestamp 1386238110
transform 1 0 9483 0 1 6939
box 0 0 120 799
use nand2 g8347
timestamp 1386234792
transform 1 0 9603 0 1 6939
box 0 0 96 799
use nand3 g8532
timestamp 1386234893
transform 1 0 9699 0 1 6939
box 0 0 120 799
use nand2 g8529
timestamp 1386234792
transform 1 0 9819 0 1 6939
box 0 0 96 799
use nand3 g8538
timestamp 1386234893
transform 1 0 9915 0 1 6939
box 0 0 120 799
use nand2 g8580
timestamp 1386234792
transform 1 0 10035 0 1 6939
box 0 0 96 799
use nand2 g8594
timestamp 1386234792
transform 1 0 10131 0 1 6939
box 0 0 96 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 10227 0 1 6939
box 0 0 48 799
use nand2 g8386
timestamp 1386234792
transform 1 0 10275 0 1 6939
box 0 0 96 799
use nand3 g8425
timestamp 1386234893
transform 1 0 10371 0 1 6939
box 0 0 120 799
use nand2 g8374
timestamp 1386234792
transform 1 0 10491 0 1 6939
box 0 0 96 799
use nand2 g8320
timestamp 1386234792
transform 1 0 10587 0 1 6939
box 0 0 96 799
use nand2 g8354
timestamp 1386234792
transform 1 0 10683 0 1 6939
box 0 0 96 799
use inv g8524
timestamp 1386238110
transform 1 0 10779 0 1 6939
box 0 0 120 799
use nand2 g8609
timestamp 1386234792
transform 1 0 10899 0 1 6939
box 0 0 96 799
use nor2 g8479
timestamp 1386235306
transform 1 0 10995 0 1 6939
box 0 0 120 799
use and2 g8564
timestamp 1386234845
transform 1 0 11115 0 1 6939
box 0 0 120 799
use nand2 g8533
timestamp 1386234792
transform 1 0 11235 0 1 6939
box 0 0 96 799
use nand3 g8627
timestamp 1386234893
transform 1 0 11331 0 1 6939
box 0 0 120 799
use inv g8306
timestamp 1386238110
transform 1 0 11451 0 1 6939
box 0 0 120 799
use nand2 g8319
timestamp 1386234792
transform 1 0 11571 0 1 6939
box 0 0 96 799
use nand3 g8431
timestamp 1386234893
transform 1 0 11667 0 1 6939
box 0 0 120 799
use nand4 g8392
timestamp 1386234936
transform 1 0 11787 0 1 6939
box 0 0 144 799
use nand4 g8340
timestamp 1386234936
transform 1 0 11931 0 1 6939
box 0 0 144 799
use nand2 rm_assigns_buf_StatusReg_1
timestamp 1386234792
transform 1 0 12075 0 1 6939
box 0 0 96 799
use buffer g8421
timestamp 1386236986
transform 1 0 12171 0 1 6939
box 0 0 120 799
use inv g8399
timestamp 1386238110
transform 1 0 12291 0 1 6939
box 0 0 120 799
use nand2 g8507
timestamp 1386234792
transform 1 0 12411 0 1 6939
box 0 0 96 799
use inv g8268
timestamp 1386238110
transform 1 0 12507 0 1 6939
box 0 0 120 799
use nand4 g8411
timestamp 1386234936
transform 1 0 12627 0 1 6939
box 0 0 144 799
use and2 g8321
timestamp 1386234845
transform 1 0 12771 0 1 6939
box 0 0 120 799
use nand2 g8379
timestamp 1386234792
transform 1 0 12891 0 1 6939
box 0 0 96 799
use nand4 g8553
timestamp 1386234936
transform 1 0 12987 0 1 6939
box 0 0 144 799
use nand2 g8417
timestamp 1386234792
transform 1 0 13131 0 1 6939
box 0 0 96 799
use nand2 g8361
timestamp 1386234792
transform 1 0 13227 0 1 6939
box 0 0 96 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 13323 0 1 6939
box 0 0 96 799
use scandtype g8308
timestamp 1386241841
transform 1 0 13419 0 1 6939
box 0 0 624 799
use nand2 stateSub_reg_91_2_93_
timestamp 1386234792
transform 1 0 14043 0 1 6939
box 0 0 96 799
use scandtype g8546
timestamp 1386241841
transform 1 0 14139 0 1 6939
box 0 0 624 799
use rowcrosser MemEn
timestamp 1386086759
transform 1 0 14763 0 1 6939
box 0 0 48 799
use inv g8372
timestamp 1386238110
transform 1 0 14811 0 1 6939
box 0 0 120 799
use nor2 g8294
timestamp 1386235306
transform 1 0 14931 0 1 6939
box 0 0 120 799
use nand3 g8444
timestamp 1386234893
transform 1 0 15051 0 1 6939
box 0 0 120 799
use and2 g8433
timestamp 1386234845
transform 1 0 15171 0 1 6939
box 0 0 120 799
use nand3 g8468
timestamp 1386234893
transform 1 0 15291 0 1 6939
box 0 0 120 799
use nand2 g8466
timestamp 1386234792
transform 1 0 15411 0 1 6939
box 0 0 96 799
use nor2 g8420
timestamp 1386235306
transform 1 0 15507 0 1 6939
box 0 0 120 799
use nand2 g8624
timestamp 1386234792
transform 1 0 15627 0 1 6939
box 0 0 96 799
use inv g8537
timestamp 1386238110
transform 1 0 15723 0 1 6939
box 0 0 120 799
use nand2 g8304
timestamp 1386234792
transform 1 0 15843 0 1 6939
box 0 0 96 799
use nand2 g8531
timestamp 1386234792
transform 1 0 15939 0 1 6939
box 0 0 96 799
use nand2 g8542
timestamp 1386234792
transform 1 0 16035 0 1 6939
box 0 0 96 799
use nor2 g8277
timestamp 1386235306
transform 1 0 16131 0 1 6939
box 0 0 120 799
use nand3 g8296
timestamp 1386234893
transform 1 0 16251 0 1 6939
box 0 0 120 799
use nand4 g8348
timestamp 1386234936
transform 1 0 16371 0 1 6939
box 0 0 144 799
use nand3 StatusReg_reg_91_1_93_
timestamp 1386234893
transform 1 0 16515 0 1 6939
box 0 0 120 799
use scandtype g8324
timestamp 1386241841
transform 1 0 16635 0 1 6939
box 0 0 624 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 17259 0 1 6939
box 0 0 48 799
use and2 g8293
timestamp 1386234845
transform 1 0 17307 0 1 6939
box 0 0 120 799
use nand3 g8435
timestamp 1386234893
transform 1 0 17427 0 1 6939
box 0 0 120 799
use nand3 g8452
timestamp 1386234893
transform 1 0 17547 0 1 6939
box 0 0 120 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 17667 0 1 6939
box 0 0 48 799
use nand3 g8312
timestamp 1386234893
transform 1 0 17715 0 1 6939
box 0 0 120 799
use nand2 g8610
timestamp 1386234792
transform 1 0 17835 0 1 6939
box 0 0 96 799
use and2 g8604
timestamp 1386234845
transform 1 0 17931 0 1 6939
box 0 0 120 799
use nand2 g8522
timestamp 1386234792
transform 1 0 18051 0 1 6939
box 0 0 96 799
use nand3 g8400
timestamp 1386234893
transform 1 0 18147 0 1 6939
box 0 0 120 799
use inv g8535
timestamp 1386238110
transform 1 0 18267 0 1 6939
box 0 0 120 799
use nor2 g8514
timestamp 1386235306
transform 1 0 18387 0 1 6939
box 0 0 120 799
use nand3 g8516
timestamp 1386234893
transform 1 0 18507 0 1 6939
box 0 0 120 799
use nand3 g8559
timestamp 1386234893
transform 1 0 18627 0 1 6939
box 0 0 120 799
use inv g8356
timestamp 1386238110
transform 1 0 18747 0 1 6939
box 0 0 120 799
use nand2 g8590
timestamp 1386234792
transform 1 0 18867 0 1 6939
box 0 0 96 799
use nand2 g8599
timestamp 1386234792
transform 1 0 18963 0 1 6939
box 0 0 96 799
use nand2 g8480
timestamp 1386234792
transform 1 0 19059 0 1 6939
box 0 0 96 799
use nand2 g8499
timestamp 1386234792
transform 1 0 19155 0 1 6939
box 0 0 96 799
use nand2 g8436
timestamp 1386234792
transform 1 0 19251 0 1 6939
box 0 0 96 799
use inv g8586
timestamp 1386238110
transform 1 0 19347 0 1 6939
box 0 0 120 799
use inv g8548
timestamp 1386238110
transform 1 0 19467 0 1 6939
box 0 0 120 799
use and2 g8332
timestamp 1386234845
transform 1 0 19587 0 1 6939
box 0 0 120 799
use nand2 g8595
timestamp 1386234792
transform 1 0 19707 0 1 6939
box 0 0 96 799
use inv g8573
timestamp 1386238110
transform 1 0 19803 0 1 6939
box 0 0 120 799
use nand2 g8278
timestamp 1386234792
transform 1 0 19923 0 1 6939
box 0 0 96 799
use nand3 g8376
timestamp 1386234893
transform 1 0 20019 0 1 6939
box 0 0 120 799
use nand3 g8630
timestamp 1386234893
transform 1 0 20139 0 1 6939
box 0 0 120 799
use inv StatusReg_reg_91_0_93_
timestamp 1386238110
transform 1 0 20259 0 1 6939
box 0 0 120 799
use scandtype g8591
timestamp 1386241841
transform 1 0 20379 0 1 6939
box 0 0 624 799
use inv g8373
timestamp 1386238110
transform 1 0 21003 0 1 6939
box 0 0 120 799
use nand2 g8443
timestamp 1386234792
transform 1 0 21123 0 1 6939
box 0 0 96 799
use and2 g8427
timestamp 1386234845
transform 1 0 21219 0 1 6939
box 0 0 120 799
use nand3 g8424
timestamp 1386234893
transform 1 0 21339 0 1 6939
box 0 0 120 799
use inv g8432
timestamp 1386238110
transform 1 0 21459 0 1 6939
box 0 0 120 799
use nand3 g8410
timestamp 1386234893
transform 1 0 21579 0 1 6939
box 0 0 120 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 21699 0 1 6939
box 0 0 48 799
use nand2 g8503
timestamp 1386234792
transform 1 0 21747 0 1 6939
box 0 0 96 799
use and2 g8588
timestamp 1386234845
transform 1 0 21843 0 1 6939
box 0 0 120 799
use and2 g8341
timestamp 1386234845
transform 1 0 21963 0 1 6939
box 0 0 120 799
use nand2 g8495
timestamp 1386234792
transform 1 0 22083 0 1 6939
box 0 0 96 799
use nor2 g8406
timestamp 1386235306
transform 1 0 22179 0 1 6939
box 0 0 120 799
use nor2 g8289
timestamp 1386235306
transform 1 0 22299 0 1 6939
box 0 0 120 799
use nand2 g8487
timestamp 1386234792
transform 1 0 22419 0 1 6939
box 0 0 96 799
use nand2 g8397
timestamp 1386234792
transform 1 0 22515 0 1 6939
box 0 0 96 799
use nand2 g8508
timestamp 1386234792
transform 1 0 22611 0 1 6939
box 0 0 96 799
use nor2 g8563
timestamp 1386235306
transform 1 0 22707 0 1 6939
box 0 0 120 799
use inv g8350
timestamp 1386238110
transform 1 0 22827 0 1 6939
box 0 0 120 799
use inv g8439
timestamp 1386238110
transform 1 0 22947 0 1 6939
box 0 0 120 799
use nand4 g8473
timestamp 1386234936
transform 1 0 23067 0 1 6939
box 0 0 144 799
use and2 g8600
timestamp 1386234845
transform 1 0 23211 0 1 6939
box 0 0 120 799
use inv g8387
timestamp 1386238110
transform 1 0 23331 0 1 6939
box 0 0 120 799
use nand3 g8270
timestamp 1386234893
transform 1 0 23451 0 1 6939
box 0 0 120 799
use nor2 g8494
timestamp 1386235306
transform 1 0 23571 0 1 6939
box 0 0 120 799
use nor2 g8465
timestamp 1386235306
transform 1 0 23691 0 1 6939
box 0 0 120 799
use nand4 g8523
timestamp 1386234936
transform 1 0 23811 0 1 6939
box 0 0 144 799
use and2 g8615
timestamp 1386234845
transform 1 0 23955 0 1 6939
box 0 0 120 799
use and2 g8455
timestamp 1386234845
transform 1 0 24075 0 1 6939
box 0 0 120 799
use inv g8273
timestamp 1386238110
transform 1 0 24195 0 1 6939
box 0 0 120 799
use nand4 g8337
timestamp 1386234936
transform 1 0 24315 0 1 6939
box 0 0 144 799
use and2 g8478
timestamp 1386234845
transform 1 0 24459 0 1 6939
box 0 0 120 799
use nand2 g8367
timestamp 1386234792
transform 1 0 24579 0 1 6939
box 0 0 96 799
use inv g8353
timestamp 1386238110
transform 1 0 24675 0 1 6939
box 0 0 120 799
use nor2 g8447
timestamp 1386235306
transform 1 0 24795 0 1 6939
box 0 0 120 799
use nand2 g8575
timestamp 1386234792
transform 1 0 24915 0 1 6939
box 0 0 96 799
use nand2 g8393
timestamp 1386234792
transform 1 0 25011 0 1 6939
box 0 0 96 799
use nand3 g8305
timestamp 1386234893
transform 1 0 25107 0 1 6939
box 0 0 120 799
use nand2 g8382
timestamp 1386234792
transform 1 0 25227 0 1 6939
box 0 0 96 799
use nand2 g8540
timestamp 1386234792
transform 1 0 25323 0 1 6939
box 0 0 96 799
use and2 g8510
timestamp 1386234845
transform 1 0 25419 0 1 6939
box 0 0 120 799
use nand2 g8257
timestamp 1386234792
transform 1 0 25539 0 1 6939
box 0 0 96 799
use nand4 g8451
timestamp 1386234936
transform 1 0 25635 0 1 6939
box 0 0 144 799
use nand2 g8519
timestamp 1386234792
transform 1 0 25779 0 1 6939
box 0 0 96 799
use nand2 LrWe
timestamp 1386234792
transform 1 0 25875 0 1 6939
box 0 0 96 799
use rowcrosser PcEn
timestamp 1386086759
transform 1 0 25971 0 1 6939
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 26019 0 1 6939
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 946
box 0 0 1464 799
use nand2 stateSub_reg_91_0_93_
timestamp 1386234792
transform 1 0 1587 0 1 946
box 0 0 96 799
use rowcrosser SysBus_91_2_93_
timestamp 1386086759
transform 1 0 1683 0 1 946
box 0 0 48 799
use scandtype g8625
timestamp 1386241841
transform 1 0 1731 0 1 946
box 0 0 624 799
use inv g8552
timestamp 1386238110
transform 1 0 2355 0 1 946
box 0 0 120 799
use nand2 g8558
timestamp 1386234792
transform 1 0 2475 0 1 946
box 0 0 96 799
use xor2 g8409
timestamp 1386237344
transform 1 0 2571 0 1 946
box 0 0 192 799
use nand2 g8430
timestamp 1386234792
transform 1 0 2763 0 1 946
box 0 0 96 799
use nand3 g8614
timestamp 1386234893
transform 1 0 2859 0 1 946
box 0 0 120 799
use nand2 g8543
timestamp 1386234792
transform 1 0 2979 0 1 946
box 0 0 96 799
use and2 g8629
timestamp 1386234845
transform 1 0 3075 0 1 946
box 0 0 120 799
use inv g8416
timestamp 1386238110
transform 1 0 3195 0 1 946
box 0 0 120 799
use nand3 state_reg_91_1_93_
timestamp 1386234893
transform 1 0 3315 0 1 946
box 0 0 120 799
use scandtype g8434
timestamp 1386241841
transform 1 0 3435 0 1 946
box 0 0 624 799
use inv g8578
timestamp 1386238110
transform 1 0 4059 0 1 946
box 0 0 120 799
use mux2 g8359
timestamp 1386235218
transform 1 0 4179 0 1 946
box 0 0 192 799
use nand2 g8300
timestamp 1386234792
transform 1 0 4371 0 1 946
box 0 0 96 799
use nand2 g8566
timestamp 1386234792
transform 1 0 4467 0 1 946
box 0 0 96 799
use and2 g8556
timestamp 1386234845
transform 1 0 4563 0 1 946
box 0 0 120 799
use nand3 g8388
timestamp 1386234893
transform 1 0 4683 0 1 946
box 0 0 120 799
use nand3 g8429
timestamp 1386234893
transform 1 0 4803 0 1 946
box 0 0 120 799
use nand4 g8611
timestamp 1386234936
transform 1 0 4923 0 1 946
box 0 0 144 799
use nand2 g8391
timestamp 1386234792
transform 1 0 5067 0 1 946
box 0 0 96 799
use nand3 g8458
timestamp 1386234893
transform 1 0 5163 0 1 946
box 0 0 120 799
use nand2 g8389
timestamp 1386234792
transform 1 0 5283 0 1 946
box 0 0 96 799
use nand4 g8307
timestamp 1386234936
transform 1 0 5379 0 1 946
box 0 0 144 799
use nand2 g8335
timestamp 1386234792
transform 1 0 5523 0 1 946
box 0 0 96 799
use nand4 g8476
timestamp 1386234936
transform 1 0 5619 0 1 946
box 0 0 144 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 5763 0 1 946
box 0 0 96 799
use scandtype g8498
timestamp 1386241841
transform 1 0 5859 0 1 946
box 0 0 624 799
use rowcrosser RegWe
timestamp 1386086759
transform 1 0 6483 0 1 946
box 0 0 48 799
use nor2 g8501
timestamp 1386235306
transform 1 0 6531 0 1 946
box 0 0 120 799
use nand3 g8401
timestamp 1386234893
transform 1 0 6651 0 1 946
box 0 0 120 799
use nor2 g8587
timestamp 1386235306
transform 1 0 6771 0 1 946
box 0 0 120 799
use nand2 g8608
timestamp 1386234792
transform 1 0 6891 0 1 946
box 0 0 96 799
use and2 g8534
timestamp 1386234845
transform 1 0 6987 0 1 946
box 0 0 120 799
use nand2 g8454
timestamp 1386234792
transform 1 0 7107 0 1 946
box 0 0 96 799
use nand2 g8442
timestamp 1386234792
transform 1 0 7203 0 1 946
box 0 0 96 799
use nand2 g8297
timestamp 1386234792
transform 1 0 7299 0 1 946
box 0 0 96 799
use nand4 g8521
timestamp 1386234936
transform 1 0 7395 0 1 946
box 0 0 144 799
use and2 g8328
timestamp 1386234845
transform 1 0 7539 0 1 946
box 0 0 120 799
use nor2 g8303
timestamp 1386235306
transform 1 0 7659 0 1 946
box 0 0 120 799
use nand3 g8394
timestamp 1386234893
transform 1 0 7779 0 1 946
box 0 0 120 799
use nand3 g8395
timestamp 1386234893
transform 1 0 7899 0 1 946
box 0 0 120 799
use nand2 g8453
timestamp 1386234792
transform 1 0 8019 0 1 946
box 0 0 96 799
use and2 g8461
timestamp 1386234845
transform 1 0 8115 0 1 946
box 0 0 120 799
use nand3 g8267
timestamp 1386234893
transform 1 0 8235 0 1 946
box 0 0 120 799
use nand4 g8282
timestamp 1386234936
transform 1 0 8355 0 1 946
box 0 0 144 799
use nand3 g8274
timestamp 1386234893
transform 1 0 8499 0 1 946
box 0 0 120 799
use nand4 g8550
timestamp 1386234936
transform 1 0 8619 0 1 946
box 0 0 144 799
use nand2 g8438
timestamp 1386234792
transform 1 0 8763 0 1 946
box 0 0 96 799
use nor2 g8349
timestamp 1386235306
transform 1 0 8859 0 1 946
box 0 0 120 799
use nand3 g8412
timestamp 1386234893
transform 1 0 8979 0 1 946
box 0 0 120 799
use and2 g8549
timestamp 1386234845
transform 1 0 9099 0 1 946
box 0 0 120 799
use and2 g8481
timestamp 1386234845
transform 1 0 9219 0 1 946
box 0 0 120 799
use nand2 g8365
timestamp 1386234792
transform 1 0 9339 0 1 946
box 0 0 96 799
use nand2 g8457
timestamp 1386234792
transform 1 0 9435 0 1 946
box 0 0 96 799
use and2 g8518
timestamp 1386234845
transform 1 0 9531 0 1 946
box 0 0 120 799
use nand2 g8301
timestamp 1386234792
transform 1 0 9651 0 1 946
box 0 0 96 799
use nand2 g8515
timestamp 1386234792
transform 1 0 9747 0 1 946
box 0 0 96 799
use nand2 g8292
timestamp 1386234792
transform 1 0 9843 0 1 946
box 0 0 96 799
use inv g8496
timestamp 1386238110
transform 1 0 9939 0 1 946
box 0 0 120 799
use nor2 g8484
timestamp 1386235306
transform 1 0 10059 0 1 946
box 0 0 120 799
use nand2 g8470
timestamp 1386234792
transform 1 0 10179 0 1 946
box 0 0 96 799
use inv g8426
timestamp 1386238110
transform 1 0 10275 0 1 946
box 0 0 120 799
use and2 g8574
timestamp 1386234845
transform 1 0 10395 0 1 946
box 0 0 120 799
use and2 g8315
timestamp 1386234845
transform 1 0 10515 0 1 946
box 0 0 120 799
use and2 g8579
timestamp 1386234845
transform 1 0 10635 0 1 946
box 0 0 120 799
use mux2 g8342
timestamp 1386235218
transform 1 0 10755 0 1 946
box 0 0 192 799
use nand2 g8509
timestamp 1386234792
transform 1 0 10947 0 1 946
box 0 0 96 799
use nor2 g8592
timestamp 1386235306
transform 1 0 11043 0 1 946
box 0 0 120 799
use nand2 g8490
timestamp 1386234792
transform 1 0 11163 0 1 946
box 0 0 96 799
use and2 g8279
timestamp 1386234845
transform 1 0 11259 0 1 946
box 0 0 120 799
use nand4 g8259
timestamp 1386234936
transform 1 0 11379 0 1 946
box 0 0 144 799
use nand4 g8500
timestamp 1386234936
transform 1 0 11523 0 1 946
box 0 0 144 799
use nand2 g8375
timestamp 1386234792
transform 1 0 11667 0 1 946
box 0 0 96 799
use and2 g8605
timestamp 1386234845
transform 1 0 11763 0 1 946
box 0 0 120 799
use nand2 g8446
timestamp 1386234792
transform 1 0 11883 0 1 946
box 0 0 96 799
use nand2 g8459
timestamp 1386234792
transform 1 0 11979 0 1 946
box 0 0 96 799
use nand2 g8560
timestamp 1386234792
transform 1 0 12075 0 1 946
box 0 0 96 799
use nand2 IntStatus_reg
timestamp 1386234792
transform 1 0 12171 0 1 946
box 0 0 96 799
use scanreg g8527
timestamp 1386241447
transform 1 0 12267 0 1 946
box 0 0 720 799
use nand2 g8570
timestamp 1386234792
transform 1 0 12987 0 1 946
box 0 0 96 799
use nand2 g8530
timestamp 1386234792
transform 1 0 13083 0 1 946
box 0 0 96 799
use nand3 g8345
timestamp 1386234893
transform 1 0 13179 0 1 946
box 0 0 120 799
use nand4 g8491
timestamp 1386234936
transform 1 0 13299 0 1 946
box 0 0 144 799
use nand4 g8322
timestamp 1386234936
transform 1 0 13443 0 1 946
box 0 0 144 799
use nand2 g8286
timestamp 1386234792
transform 1 0 13587 0 1 946
box 0 0 96 799
use inv g8368
timestamp 1386238110
transform 1 0 13683 0 1 946
box 0 0 120 799
use nand2 g8437
timestamp 1386234792
transform 1 0 13803 0 1 946
box 0 0 96 799
use nor2 g8331
timestamp 1386235306
transform 1 0 13899 0 1 946
box 0 0 120 799
use nand2 g8336
timestamp 1386234792
transform 1 0 14019 0 1 946
box 0 0 96 799
use nand2 g8526
timestamp 1386234792
transform 1 0 14115 0 1 946
box 0 0 96 799
use nand3 g8423
timestamp 1386234893
transform 1 0 14211 0 1 946
box 0 0 120 799
use nand2 g8383
timestamp 1386234792
transform 1 0 14331 0 1 946
box 0 0 96 799
use nand2 g8405
timestamp 1386234792
transform 1 0 14427 0 1 946
box 0 0 96 799
use nand2 g8601
timestamp 1386234792
transform 1 0 14523 0 1 946
box 0 0 96 799
use nand2 g8582
timestamp 1386234792
transform 1 0 14619 0 1 946
box 0 0 96 799
use nor2 g8398
timestamp 1386235306
transform 1 0 14715 0 1 946
box 0 0 120 799
use nand2 g8464
timestamp 1386234792
transform 1 0 14835 0 1 946
box 0 0 96 799
use nand3 g8325
timestamp 1386234893
transform 1 0 14931 0 1 946
box 0 0 120 799
use nor2 g8568
timestamp 1386235306
transform 1 0 15051 0 1 946
box 0 0 120 799
use nand2 g8460
timestamp 1386234792
transform 1 0 15171 0 1 946
box 0 0 96 799
use nand3 g8317
timestamp 1386234893
transform 1 0 15267 0 1 946
box 0 0 120 799
use nand3 g8404
timestamp 1386234893
transform 1 0 15387 0 1 946
box 0 0 120 799
use nand2 g8428
timestamp 1386234792
transform 1 0 15507 0 1 946
box 0 0 96 799
use nand2 g8413
timestamp 1386234792
transform 1 0 15603 0 1 946
box 0 0 96 799
use nand2 g8577
timestamp 1386234792
transform 1 0 15699 0 1 946
box 0 0 96 799
use nor2 g8358
timestamp 1386235306
transform 1 0 15795 0 1 946
box 0 0 120 799
use nor2 g8323
timestamp 1386235306
transform 1 0 15915 0 1 946
box 0 0 120 799
use nand4 g8571
timestamp 1386234936
transform 1 0 16035 0 1 946
box 0 0 144 799
use nand2 g8408
timestamp 1386234792
transform 1 0 16179 0 1 946
box 0 0 96 799
use inv g8380
timestamp 1386238110
transform 1 0 16275 0 1 946
box 0 0 120 799
use nand4 g8309
timestamp 1386234936
transform 1 0 16395 0 1 946
box 0 0 144 799
use nand2 IRQ2_reg
timestamp 1386234792
transform 1 0 16539 0 1 946
box 0 0 96 799
use scandtype g8602
timestamp 1386241841
transform 1 0 16635 0 1 946
box 0 0 624 799
use nand2 g8593
timestamp 1386234792
transform 1 0 17259 0 1 946
box 0 0 96 799
use nand2 g8517
timestamp 1386234792
transform 1 0 17355 0 1 946
box 0 0 96 799
use inv g8402
timestamp 1386238110
transform 1 0 17451 0 1 946
box 0 0 120 799
use nand2 g8422
timestamp 1386234792
transform 1 0 17571 0 1 946
box 0 0 96 799
use nand2 g8622
timestamp 1386234792
transform 1 0 17667 0 1 946
box 0 0 96 799
use inv g8488
timestamp 1386238110
transform 1 0 17763 0 1 946
box 0 0 120 799
use nand2 g8633
timestamp 1386234792
transform 1 0 17883 0 1 946
box 0 0 96 799
use inv g8475
timestamp 1386238110
transform 1 0 17979 0 1 946
box 0 0 120 799
use nand2 g8415
timestamp 1386234792
transform 1 0 18099 0 1 946
box 0 0 96 799
use inv g8555
timestamp 1386238110
transform 1 0 18195 0 1 946
box 0 0 120 799
use and2 g8598
timestamp 1386234845
transform 1 0 18315 0 1 946
box 0 0 120 799
use inv g8299
timestamp 1386238110
transform 1 0 18435 0 1 946
box 0 0 120 799
use and2 g8520
timestamp 1386234845
transform 1 0 18555 0 1 946
box 0 0 120 799
use nand2 g8326
timestamp 1386234792
transform 1 0 18675 0 1 946
box 0 0 96 799
use nand2 g8396
timestamp 1386234792
transform 1 0 18771 0 1 946
box 0 0 96 799
use inv g8617
timestamp 1386238110
transform 1 0 18867 0 1 946
box 0 0 120 799
use nor2 IRQ1_reg
timestamp 1386235306
transform 1 0 18987 0 1 946
box 0 0 120 799
use scandtype g8502
timestamp 1386241841
transform 1 0 19107 0 1 946
box 0 0 624 799
use rowcrosser SysBus_91_3_93_
timestamp 1386086759
transform 1 0 19731 0 1 946
box 0 0 48 799
use nand3 g8505
timestamp 1386234893
transform 1 0 19779 0 1 946
box 0 0 120 799
use nand2 g8419
timestamp 1386234792
transform 1 0 19899 0 1 946
box 0 0 96 799
use nand2 g8329
timestamp 1386234792
transform 1 0 19995 0 1 946
box 0 0 96 799
use and2 g8596
timestamp 1386234845
transform 1 0 20091 0 1 946
box 0 0 120 799
use nand2 g8463
timestamp 1386234792
transform 1 0 20211 0 1 946
box 0 0 96 799
use nand3 g8339
timestamp 1386234893
transform 1 0 20307 0 1 946
box 0 0 120 799
use nand2 g8557
timestamp 1386234792
transform 1 0 20427 0 1 946
box 0 0 96 799
use nand3 g8607
timestamp 1386234893
transform 1 0 20523 0 1 946
box 0 0 120 799
use nand2 g8260
timestamp 1386234792
transform 1 0 20643 0 1 946
box 0 0 96 799
use nand2 g8471
timestamp 1386234792
transform 1 0 20739 0 1 946
box 0 0 96 799
use nor2 g8351
timestamp 1386235306
transform 1 0 20835 0 1 946
box 0 0 120 799
use nand4 g8492
timestamp 1386234936
transform 1 0 20955 0 1 946
box 0 0 144 799
use inv g8343
timestamp 1386238110
transform 1 0 21099 0 1 946
box 0 0 120 799
use nand2 g8288
timestamp 1386234792
transform 1 0 21219 0 1 946
box 0 0 96 799
use nor2 g8583
timestamp 1386235306
transform 1 0 21315 0 1 946
box 0 0 120 799
use nand2 g8384
timestamp 1386234792
transform 1 0 21435 0 1 946
box 0 0 96 799
use and2 g8311
timestamp 1386234845
transform 1 0 21531 0 1 946
box 0 0 120 799
use nand2 g8621
timestamp 1386234792
transform 1 0 21651 0 1 946
box 0 0 96 799
use inv g8298
timestamp 1386238110
transform 1 0 21747 0 1 946
box 0 0 120 799
use nand2 g8346
timestamp 1386234792
transform 1 0 21867 0 1 946
box 0 0 96 799
use inv g8385
timestamp 1386238110
transform 1 0 21963 0 1 946
box 0 0 120 799
use nand3 g8355
timestamp 1386234893
transform 1 0 22083 0 1 946
box 0 0 120 799
use nand2 g8330
timestamp 1386234792
transform 1 0 22203 0 1 946
box 0 0 96 799
use nand2 g8360
timestamp 1386234792
transform 1 0 22299 0 1 946
box 0 0 96 799
use nand2 g8258
timestamp 1386234792
transform 1 0 22395 0 1 946
box 0 0 96 799
use nand4 g8482
timestamp 1386234936
transform 1 0 22491 0 1 946
box 0 0 144 799
use nand2 g8467
timestamp 1386234792
transform 1 0 22635 0 1 946
box 0 0 96 799
use nor2 g8371
timestamp 1386235306
transform 1 0 22731 0 1 946
box 0 0 120 799
use nand2 g8539
timestamp 1386234792
transform 1 0 22851 0 1 946
box 0 0 96 799
use nor2 g8285
timestamp 1386235306
transform 1 0 22947 0 1 946
box 0 0 120 799
use nand3 g8565
timestamp 1386234893
transform 1 0 23067 0 1 946
box 0 0 120 799
use and2 g8551
timestamp 1386234845
transform 1 0 23187 0 1 946
box 0 0 120 799
use nand2 g8497
timestamp 1386234792
transform 1 0 23307 0 1 946
box 0 0 96 799
use inv g8485
timestamp 1386238110
transform 1 0 23403 0 1 946
box 0 0 120 799
use nand2 g8613
timestamp 1386234792
transform 1 0 23523 0 1 946
box 0 0 96 799
use inv g8544
timestamp 1386238110
transform 1 0 23619 0 1 946
box 0 0 120 799
use inv g8569
timestamp 1386238110
transform 1 0 23739 0 1 946
box 0 0 120 799
use and2 state_reg_91_0_93_
timestamp 1386234845
transform 1 0 23859 0 1 946
box 0 0 120 799
use scandtype g8441
timestamp 1386241841
transform 1 0 23979 0 1 946
box 0 0 624 799
use nand3 g8302
timestamp 1386234893
transform 1 0 24603 0 1 946
box 0 0 120 799
use nor2 stateSub_reg_91_1_93_
timestamp 1386235306
transform 1 0 24723 0 1 946
box 0 0 120 799
use scandtype g8316
timestamp 1386241841
transform 1 0 24843 0 1 946
box 0 0 624 799
use nand3 g8378
timestamp 1386234893
transform 1 0 25467 0 1 946
box 0 0 120 799
use nand2 nIRQ
timestamp 1386234792
transform 1 0 25587 0 1 946
box 0 0 96 799
use rowcrosser AluOR_91_0_93_
timestamp 1386086759
transform 1 0 25683 0 1 946
box 0 0 48 799
use rowcrosser g8364
timestamp 1386086759
transform 1 0 25731 0 1 946
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 26019 0 1 946
box 0 0 320 799
<< labels >>
rlabel m2contact 25809 521 25809 521 8 AluOR[0]
rlabel m2contact 25809 65 25809 65 8 AluOR[0]
rlabel m2contact 25785 713 25785 713 8 ENB
rlabel m2contact 25785 17 25785 17 8 ENB
rlabel m2contact 25761 473 25761 473 8 AluOR[1]
rlabel m2contact 25761 41 25761 41 8 AluOR[1]
rlabel m2contact 25761 521 25761 521 8 AluOR[0]
rlabel m2contact 25713 497 25713 497 8 RegWe
rlabel m2contact 25521 497 25521 497 8 n_248
rlabel m2contact 24825 569 24825 569 8 n_318
rlabel m2contact 24777 233 24777 233 8 n_75
rlabel m2contact 24441 905 24441 905 6 n_7
rlabel m2contact 23817 545 23817 545 8 n_114
rlabel m2contact 23553 353 23553 353 8 n_111
rlabel m2contact 23169 473 23169 473 8 AluOR[1]
rlabel m2contact 22929 329 22929 329 8 n_284
rlabel m2contact 22713 305 22713 305 8 n_102
rlabel m2contact 22569 833 22569 833 6 n_313
rlabel m2contact 22425 665 22425 665 8 n_221
rlabel m2contact 22353 449 22353 449 8 SysBus[0]
rlabel m2contact 22257 761 22257 761 8 n_244
rlabel m2contact 22185 641 22185 641 8 n_204
rlabel m2contact 22041 593 22041 593 8 n_331
rlabel m2contact 21945 65 21945 65 8 nWE
rlabel m2contact 21729 617 21729 617 8 n_287
rlabel m2contact 21489 377 21489 377 8 n_480
rlabel m2contact 21345 737 21345 737 8 n_339
rlabel m2contact 21297 785 21297 785 8 n_308
rlabel m2contact 21057 473 21057 473 8 n_54
rlabel m2contact 21033 521 21033 521 8 n_151
rlabel m2contact 20985 689 20985 689 8 n_44
rlabel m2contact 20937 857 20937 857 6 n_120
rlabel m2contact 20505 929 20505 929 6 n_239
rlabel m2contact 20193 713 20193 713 8 ENB
rlabel m2contact 19953 545 19953 545 8 n_114
rlabel m2contact 19905 17 19905 17 8 SysBus[3]
rlabel m2contact 19881 689 19881 689 8 n_44
rlabel metal2 19779 689 19779 689 8 SysBus[2]
rlabel m2contact 19761 689 19761 689 8 SysBus[2]
rlabel m2contact 19617 713 19617 713 8 IRQ1
rlabel m2contact 18945 689 18945 689 8 n_197
rlabel m2contact 18825 209 18825 209 8 n_184
rlabel m2contact 17961 137 17961 137 8 n_101
rlabel m2contact 17913 185 17913 185 8 n_25
rlabel m2contact 17841 401 17841 401 8 n_19
rlabel m2contact 17649 761 17649 761 8 n_244
rlabel m2contact 17481 353 17481 353 8 n_111
rlabel m2contact 17337 113 17337 113 8 n_14
rlabel m2contact 17145 881 17145 881 6 IRQ2
rlabel m2contact 16737 713 16737 713 8 IRQ1
rlabel m2contact 16353 665 16353 665 8 n_221
rlabel m2contact 16161 281 16161 281 8 n_205
rlabel m2contact 15897 809 15897 809 6 n_43
rlabel m2contact 15825 425 15825 425 8 n_22
rlabel m2contact 15777 89 15777 89 8 n_238
rlabel m2contact 15585 665 15585 665 8 n_225
rlabel m2contact 15465 641 15465 641 8 n_204
rlabel m2contact 15249 257 15249 257 8 n_55
rlabel m2contact 15153 641 15153 641 8 n_298
rlabel m2contact 15081 713 15081 713 8 n_240
rlabel m2contact 15009 881 15009 881 6 IRQ2
rlabel m2contact 14985 761 14985 761 8 n_91
rlabel m2contact 14961 161 14961 161 8 IntStatus
rlabel m2contact 14313 41 14313 41 8 n_78
rlabel m2contact 14169 329 14169 329 8 n_284
rlabel m2contact 14073 329 14073 329 8 SysBus[1]
rlabel m2contact 13785 329 13785 329 8 SysBus[1]
rlabel m2contact 13761 833 13761 833 6 n_313
rlabel m2contact 13617 329 13617 329 8 n_140
rlabel m2contact 13473 905 13473 905 4 n_7
rlabel m2contact 13329 833 13329 833 4 n_154
rlabel m2contact 13281 185 13281 185 2 n_25
rlabel m2contact 13161 473 13161 473 2 n_54
rlabel m2contact 13041 473 13041 473 2 n_18
rlabel m2contact 13017 257 13017 257 2 n_55
rlabel m2contact 12873 161 12873 161 2 IntStatus
rlabel m2contact 12345 785 12345 785 2 n_308
rlabel m2contact 12153 185 12153 185 2 n_131
rlabel m2contact 11961 473 11961 473 2 n_18
rlabel m2contact 11865 473 11865 473 2 n_281
rlabel m2contact 11601 785 11601 785 2 n_247
rlabel m2contact 11433 257 11433 257 2 n_200
rlabel m2contact 11409 929 11409 929 4 n_239
rlabel m2contact 11217 905 11217 905 4 n_7
rlabel m2contact 11145 233 11145 233 2 n_75
rlabel m2contact 11025 233 11025 233 2 n_309
rlabel m2contact 10665 281 10665 281 2 n_205
rlabel m2contact 10497 281 10497 281 2 n_163
rlabel m2contact 10449 881 10449 881 4 IRQ2
rlabel m2contact 10425 185 10425 185 2 n_131
rlabel m2contact 10353 185 10353 185 2 n_130
rlabel m2contact 10305 857 10305 857 4 n_120
rlabel m2contact 10257 833 10257 833 4 n_154
rlabel m2contact 10089 809 10089 809 4 n_43
rlabel m2contact 10017 785 10017 785 2 n_247
rlabel m2contact 9921 761 9921 761 2 n_91
rlabel m2contact 9825 737 9825 737 2 n_339
rlabel m2contact 9801 89 9801 89 2 n_238
rlabel m2contact 9729 353 9729 353 2 n_111
rlabel m2contact 9633 353 9633 353 2 n_168
rlabel m2contact 9585 89 9585 89 2 n_143
rlabel m2contact 9561 137 9561 137 2 n_101
rlabel m2contact 9369 137 9369 137 2 n_92
rlabel m2contact 9201 713 9201 713 2 n_240
rlabel m2contact 9033 689 9033 689 2 n_197
rlabel m2contact 8721 665 8721 665 2 n_225
rlabel m2contact 8673 641 8673 641 2 n_298
rlabel m2contact 8529 617 8529 617 2 n_287
rlabel m2contact 8433 593 8433 593 2 n_331
rlabel m2contact 8385 569 8385 569 2 n_318
rlabel m2contact 8313 545 8313 545 2 n_114
rlabel m2contact 8097 521 8097 521 2 n_151
rlabel m2contact 8001 497 8001 497 2 n_248
rlabel m2contact 7689 473 7689 473 2 n_281
rlabel m2contact 7677 449 7677 449 2 SysBus[0]
rlabel m2contact 7497 161 7497 161 2 IntStatus
rlabel m2contact 7473 281 7473 281 2 n_163
rlabel m2contact 7185 281 7185 281 2 n_42
rlabel m2contact 7161 161 7161 161 2 n_4
rlabel m2contact 7089 425 7089 425 2 n_22
rlabel m2contact 6921 401 6921 401 2 n_19
rlabel m2contact 6729 401 6729 401 2 n_19
rlabel m2contact 6513 17 6513 17 2 SysBus[3]
rlabel m2contact 6321 377 6321 377 2 n_480
rlabel m2contact 5841 89 5841 89 2 n_143
rlabel m2contact 5721 89 5721 89 2 n_183
rlabel m2contact 5697 353 5697 353 2 n_168
rlabel m2contact 5505 329 5505 329 2 n_140
rlabel m2contact 5433 305 5433 305 2 n_102
rlabel m2contact 5337 41 5337 41 2 n_78
rlabel m2contact 5049 41 5049 41 2 n_125
rlabel m2contact 4953 281 4953 281 2 n_42
rlabel m2contact 4905 257 4905 257 2 n_200
rlabel m2contact 4497 233 4497 233 2 n_309
rlabel m2contact 4449 209 4449 209 2 n_184
rlabel m2contact 4425 185 4425 185 2 n_130
rlabel m2contact 4401 89 4401 89 2 n_183
rlabel m2contact 4137 89 4137 89 2 n_183
rlabel m2contact 2553 89 2553 89 2 n_57
rlabel m2contact 2433 161 2433 161 2 n_4
rlabel m2contact 1833 41 1833 41 2 n_125
rlabel m2contact 1713 41 1713 41 2 nIRQ
rlabel m2contact 1665 137 1665 137 2 n_92
rlabel m2contact 1641 113 1641 113 2 n_14
rlabel m2contact 1617 89 1617 89 2 n_57
rlabel m2contact 26121 7923 26121 7923 6 Flags[2]
rlabel m2contact 26121 7803 26121 7803 6 Flags[2]
rlabel m2contact 26097 7851 26097 7851 6 CFlag
rlabel m2contact 26097 7803 26097 7803 6 CFlag
rlabel m2contact 26073 7995 26073 7995 6 Flags[3]
rlabel m2contact 26073 7827 26073 7827 6 Flags[3]
rlabel m2contact 26049 7899 26049 7899 6 Flags[1]
rlabel m2contact 26049 7779 26049 7779 6 Flags[1]
rlabel m2contact 26025 7827 26025 7827 6 Flags[0]
rlabel m2contact 26025 7755 26025 7755 6 Flags[0]
rlabel m2contact 26001 7899 26001 7899 6 Flags[1]
rlabel m2contact 25089 7779 25089 7779 6 StatusRegEn
rlabel m2contact 24753 7971 24753 7971 6 LrSel
rlabel m2contact 24441 8019 24441 8019 6 AluWe
rlabel m2contact 24285 7947 24285 7947 6 StatusReg[3]
rlabel m2contact 23625 7755 23625 7755 6 Op1Sel
rlabel m2contact 23481 7899 23481 7899 6 StatusReg[2]
rlabel m2contact 22677 7851 22677 7851 6 StatusReg[1]
rlabel m2contact 21873 7875 21873 7875 6 StatusReg[0]
rlabel metal2 21747 8043 21747 8043 6 AluEn
rlabel m2contact 21729 8043 21729 8043 6 AluEn
rlabel m2contact 21045 8019 21045 8019 6 AluWe
rlabel m2contact 20889 7875 20889 7875 6 StatusReg[0]
rlabel m2contact 19461 8019 19461 8019 6 Op2Sel[1]
rlabel m2contact 18657 7875 18657 7875 6 Op2Sel[0]
rlabel m2contact 18633 7755 18633 7755 6 Op1Sel
rlabel m2contact 17889 7995 17889 7995 6 Flags[3]
rlabel metal2 17715 7995 17715 7995 6 PcEn
rlabel m2contact 17697 7995 17697 7995 6 PcEn
rlabel m2contact 17289 7923 17289 7923 6 Flags[2]
rlabel m2contact 17145 7803 17145 7803 6 CFlag
rlabel m2contact 16353 7875 16353 7875 6 Op2Sel[0]
rlabel m2contact 16245 7923 16245 7923 6 WdSel
rlabel m2contact 15441 7875 15441 7875 6 PcWe
rlabel m2contact 15273 7779 15273 7779 6 StatusRegEn
rlabel m2contact 15153 7779 15153 7779 6 PcSel[1]
rlabel m2contact 15033 7923 15033 7923 6 WdSel
rlabel m2contact 14793 7995 14793 7995 6 LrWe
rlabel m2contact 14637 7923 14637 7923 6 PcSel[2]
rlabel m2contact 14613 7779 14613 7779 6 PcSel[1]
rlabel m2contact 14097 7803 14097 7803 6 CFlag
rlabel m2contact 13929 7947 13929 7947 6 StatusReg[3]
rlabel m2contact 13029 7947 13029 7947 4 PcSel[0]
rlabel m2contact 12753 8019 12753 8019 4 Op2Sel[1]
rlabel m2contact 12249 7851 12249 7851 4 StatusReg[1]
rlabel m2contact 12213 7851 12213 7851 4 LrEn
rlabel m2contact 12201 7803 12201 7803 4 CFlag
rlabel m2contact 12177 7995 12177 7995 4 LrWe
rlabel m2contact 11625 7827 11625 7827 4 Flags[0]
rlabel m2contact 11409 7827 11409 7827 4 OpcodeCondIn[2]
rlabel m2contact 11361 7971 11361 7971 4 LrSel
rlabel metal2 10275 7971 10275 7971 4 ImmSel
rlabel m2contact 10257 7971 10257 7971 4 ImmSel
rlabel m2contact 9993 7971 9993 7971 4 OpcodeCondIn[6]
rlabel metal2 9387 7995 9387 7995 4 IrWe
rlabel m2contact 9369 7995 9369 7995 4 IrWe
rlabel metal2 8499 7995 8499 7995 4 MemEn
rlabel m2contact 8481 7995 8481 7995 4 MemEn
rlabel m2contact 8433 7851 8433 7851 4 LrEn
rlabel metal2 8019 7851 8019 7851 4 OpcodeCondIn[7]
rlabel m2contact 8001 7851 8001 7851 4 OpcodeCondIn[7]
rlabel m2contact 7281 7971 7281 7971 4 OpcodeCondIn[6]
rlabel m2contact 7281 7875 7281 7875 4 PcWe
rlabel m2contact 6801 7851 6801 7851 4 OpcodeCondIn[1]
rlabel m2contact 6297 7899 6297 7899 4 StatusReg[2]
rlabel m2contact 5685 7875 5685 7875 4 OpcodeCondIn[5]
rlabel m2contact 5337 7899 5337 7899 4 OpcodeCondIn[0]
rlabel metal2 5259 7971 5259 7971 4 OpcodeCondIn[4]
rlabel m2contact 5241 7971 5241 7971 4 OpcodeCondIn[4]
rlabel m2contact 4053 7971 4053 7971 4 OpcodeCondIn[3]
rlabel m2contact 4017 7827 4017 7827 4 OpcodeCondIn[2]
rlabel m2contact 3633 7971 3633 7971 4 OpcodeCondIn[3]
rlabel m2contact 3489 7947 3489 7947 4 PcSel[0]
rlabel m2contact 3273 7923 3273 7923 4 PcSel[2]
rlabel m2contact 3201 7851 3201 7851 4 OpcodeCondIn[1]
rlabel m2contact 3009 7875 3009 7875 4 OpcodeCondIn[5]
rlabel m2contact 2385 7899 2385 7899 4 OpcodeCondIn[0]
rlabel m2contact 2241 7875 2241 7875 4 nME
rlabel m2contact 1689 7899 1689 7899 4 ALE
rlabel m2contact 26001 5602 26001 5602 6 Flags[1]
rlabel m2contact 25953 2794 25953 2794 6 n_63
rlabel m2contact 25929 3730 25929 3730 6 stateSub[0]
rlabel m2contact 25905 2002 25905 2002 6 n_32
rlabel m2contact 25881 5818 25881 5818 6 RegWe
rlabel m2contact 25881 4354 25881 4354 6 RegWe
rlabel m2contact 25857 5026 25857 5026 6 n_170
rlabel m2contact 25833 6058 25833 6058 6 n_95
rlabel m2contact 25809 5986 25809 5986 6 n_174
rlabel m2contact 25785 6898 25785 6898 6 n_181
rlabel m2contact 25785 2266 25785 2266 6 n_181
rlabel m2contact 25761 5818 25761 5818 6 RegWe
rlabel m2contact 25761 5770 25761 5770 6 AluOR[0]
rlabel m2contact 25737 5794 25737 5794 6 n_356
rlabel m2contact 25713 4354 25713 4354 6 RegWe
rlabel m2contact 25713 5170 25713 5170 6 n_345
rlabel m2contact 25689 3514 25689 3514 6 n_227
rlabel m2contact 25665 2266 25665 2266 6 n_181
rlabel m2contact 25665 2314 25665 2314 6 n_346
rlabel m2contact 25641 5866 25641 5866 6 n_165
rlabel m2contact 25617 6058 25617 6058 6 n_95
rlabel m2contact 25617 6034 25617 6034 6 n_180
rlabel m2contact 25593 2026 25593 2026 6 n_93
rlabel m2contact 25569 6154 25569 6154 6 n_94
rlabel m2contact 25569 2962 25569 2962 6 n_315
rlabel m2contact 25545 6322 25545 6322 6 n_192
rlabel m2contact 25521 6058 25521 6058 6 n_135
rlabel m2contact 25497 6682 25497 6682 6 n_291
rlabel m2contact 25473 4498 25473 4498 6 n_210
rlabel m2contact 25449 5506 25449 5506 6 n_39
rlabel m2contact 25425 5842 25425 5842 6 n_219
rlabel m2contact 25425 5698 25425 5698 6 n_219
rlabel m2contact 25401 1834 25401 1834 6 n_259
rlabel m2contact 25377 5410 25377 5410 6 OpcodeCondIn[4]
rlabel m2contact 25353 5842 25353 5842 6 n_219
rlabel m2contact 25353 5746 25353 5746 6 stateSub[1]
rlabel m2contact 25329 5818 25329 5818 6 n_292
rlabel m2contact 25329 4594 25329 4594 6 n_292
rlabel m2contact 25305 5818 25305 5818 6 n_292
rlabel m2contact 25305 5722 25305 5722 6 n_10
rlabel m2contact 25281 2866 25281 2866 6 StatusReg[0]
rlabel m2contact 25257 2650 25257 2650 6 n_289
rlabel m2contact 25209 4330 25209 4330 6 n_251
rlabel m2contact 25185 2050 25185 2050 6 n_264
rlabel m2contact 25161 3970 25161 3970 6 n_250
rlabel m2contact 25137 2818 25137 2818 6 n_199
rlabel m2contact 25089 4618 25089 4618 6 n_37
rlabel m2contact 25065 2026 25065 2026 6 n_93
rlabel m2contact 25041 2770 25041 2770 6 n_68
rlabel m2contact 24993 5626 24993 5626 6 n_173
rlabel m2contact 24969 3322 24969 3322 6 OpcodeCondIn[3]
rlabel m2contact 24945 5890 24945 5890 6 n_332
rlabel m2contact 24945 5986 24945 5986 6 n_174
rlabel m2contact 24897 2578 24897 2578 6 n_268
rlabel m2contact 24849 3394 24849 3394 6 n_269
rlabel m2contact 24825 1762 24825 1762 6 n_267
rlabel m2contact 24753 6442 24753 6442 6 n_279
rlabel m2contact 24729 4354 24729 4354 6 n_106
rlabel m2contact 24729 1882 24729 1882 6 n_106
rlabel m2contact 24705 2602 24705 2602 6 n_316
rlabel m2contact 24705 2218 24705 2218 6 n_178
rlabel m2contact 24681 3178 24681 3178 6 n_176
rlabel m2contact 24657 6706 24657 6706 6 n_117
rlabel m2contact 24657 4282 24657 4282 6 n_155
rlabel m2contact 24633 4354 24633 4354 6 n_106
rlabel m2contact 24633 3586 24633 3586 6 n_177
rlabel m2contact 24609 1786 24609 1786 6 n_81
rlabel m2contact 24561 5218 24561 5218 6 n_347
rlabel m2contact 24513 5794 24513 5794 6 n_356
rlabel m2contact 24489 4450 24489 4450 6 n_282
rlabel m2contact 24489 2938 24489 2938 6 state[0]
rlabel m2contact 24417 3490 24417 3490 6 n_209
rlabel m2contact 24393 2194 24393 2194 6 n_358
rlabel m2contact 24369 4186 24369 4186 6 n_359
rlabel m2contact 24345 4546 24345 4546 6 n_262
rlabel m2contact 24273 4354 24273 4354 6 n_193
rlabel m2contact 24225 3442 24225 3442 6 n_157
rlabel m2contact 24177 1882 24177 1882 6 n_106
rlabel m2contact 24153 4834 24153 4834 6 n_172
rlabel m2contact 24153 3658 24153 3658 6 n_172
rlabel m2contact 24129 3346 24129 3346 6 OpcodeCondIn[6]
rlabel m2contact 24105 4762 24105 4762 6 OpcodeCondIn[7]
rlabel m2contact 24081 6394 24081 6394 6 n_333
rlabel m2contact 24057 1858 24057 1858 6 n_79
rlabel m2contact 24033 5794 24033 5794 6 n_356
rlabel m2contact 24033 1954 24033 1954 6 n_356
rlabel m2contact 24009 2818 24009 2818 6 n_199
rlabel m2contact 23985 5674 23985 5674 6 n_48
rlabel m2contact 23961 2698 23961 2698 6 n_139
rlabel m2contact 23937 6178 23937 6178 6 n_124
rlabel m2contact 23913 3658 23913 3658 6 n_172
rlabel m2contact 23913 3682 23913 3682 6 nWait
rlabel m2contact 23889 2026 23889 2026 6 n_93
rlabel m2contact 23889 5146 23889 5146 6 n_203
rlabel m2contact 23865 3730 23865 3730 6 stateSub[0]
rlabel m2contact 23841 4930 23841 4930 6 n_123
rlabel m2contact 23805 4522 23805 4522 6 n_128
rlabel m2contact 23805 2122 23805 2122 6 n_128
rlabel m2contact 23793 5242 23793 5242 6 n_45
rlabel m2contact 23769 4858 23769 4858 6 n_74
rlabel m2contact 23745 5122 23745 5122 6 n_17
rlabel m2contact 23721 3850 23721 3850 6 state[1]
rlabel m2contact 23697 3394 23697 3394 6 n_269
rlabel m2contact 23673 4162 23673 4162 6 n_368
rlabel m2contact 23649 3274 23649 3274 6 n_16
rlabel m2contact 23625 4042 23625 4042 6 Op1Sel
rlabel m2contact 23601 2122 23601 2122 6 n_128
rlabel m2contact 23601 2146 23601 2146 6 n_360
rlabel m2contact 23577 4954 23577 4954 6 n_24
rlabel m2contact 23553 2458 23553 2458 6 n_202
rlabel m2contact 23529 2842 23529 2842 6 n_256
rlabel m2contact 23505 4738 23505 4738 6 n_201
rlabel m2contact 23481 5002 23481 5002 6 n_119
rlabel m2contact 23481 6754 23481 6754 6 n_257
rlabel m2contact 23445 4978 23445 4978 6 n_68
rlabel m2contact 23445 2770 23445 2770 6 n_68
rlabel m2contact 23433 2554 23433 2554 6 n_100
rlabel m2contact 23409 5842 23409 5842 6 n_56
rlabel m2contact 23385 5554 23385 5554 6 n_35
rlabel m2contact 23361 4978 23361 4978 6 n_68
rlabel m2contact 23361 4930 23361 4930 6 n_123
rlabel m2contact 23337 4210 23337 4210 6 n_208
rlabel m2contact 23313 6010 23313 6010 6 n_147
rlabel m2contact 23289 6034 23289 6034 6 n_180
rlabel m2contact 23265 2386 23265 2386 6 n_134
rlabel m2contact 23241 4930 23241 4930 6 n_123
rlabel m2contact 23241 3898 23241 3898 6 n_319
rlabel m2contact 23217 4114 23217 4114 6 n_84
rlabel m2contact 23193 1978 23193 1978 6 n_179
rlabel m2contact 23169 4834 23169 4834 6 n_172
rlabel m2contact 23145 4522 23145 4522 6 n_128
rlabel m2contact 23145 4474 23145 4474 6 n_229
rlabel m2contact 23121 2338 23121 2338 6 n_343
rlabel m2contact 23121 4930 23121 4930 6 n_123
rlabel m2contact 23097 1954 23097 1954 6 n_356
rlabel m2contact 23097 2050 23097 2050 6 n_264
rlabel m2contact 23073 6130 23073 6130 6 n_213
rlabel m2contact 23073 4066 23073 4066 6 n_213
rlabel m2contact 23049 4714 23049 4714 6 n_241
rlabel m2contact 23025 5074 23025 5074 6 n_234
rlabel m2contact 23001 3298 23001 3298 6 OpcodeCondIn[2]
rlabel m2contact 22977 6130 22977 6130 6 n_213
rlabel m2contact 22977 6106 22977 6106 6 n_5
rlabel m2contact 22929 4378 22929 4378 6 n_256
rlabel m2contact 22929 2842 22929 2842 6 n_256
rlabel m2contact 22929 4786 22929 4786 6 n_196
rlabel m2contact 22929 4402 22929 4402 6 n_196
rlabel m2contact 22905 4378 22905 4378 6 n_256
rlabel m2contact 22905 3394 22905 3394 6 n_269
rlabel m2contact 22881 5050 22881 5050 6 n_283
rlabel m2contact 22857 2530 22857 2530 6 n_67
rlabel m2contact 22833 5314 22833 5314 6 n_122
rlabel m2contact 22809 6826 22809 6826 6 n_98
rlabel m2contact 22785 4378 22785 4378 6 n_34
rlabel m2contact 22761 1858 22761 1858 6 n_79
rlabel m2contact 22761 1906 22761 1906 6 n_96
rlabel m2contact 22737 3202 22737 3202 6 n_97
rlabel m2contact 22713 6538 22713 6538 6 n_222
rlabel m2contact 22713 4258 22713 4258 6 n_222
rlabel m2contact 22689 4786 22689 4786 6 n_196
rlabel m2contact 22689 4762 22689 4762 6 OpcodeCondIn[7]
rlabel m2contact 22665 2986 22665 2986 6 n_108
rlabel m2contact 22665 4498 22665 4498 6 n_210
rlabel m2contact 22641 4354 22641 4354 6 n_193
rlabel m2contact 22617 4306 22617 4306 6 Rs1Sel[0]
rlabel m2contact 22593 6298 22593 6298 6 n_158
rlabel m2contact 22593 3898 22593 3898 6 n_319
rlabel m2contact 22569 2410 22569 2410 6 stateSub[2]
rlabel m2contact 22545 3802 22545 3802 6 n_118
rlabel m2contact 22545 4306 22545 4306 6 n_194
rlabel m2contact 22521 1858 22521 1858 6 n_245
rlabel m2contact 22497 6346 22497 6346 6 n_311
rlabel m2contact 22473 2362 22473 2362 6 n_300
rlabel m2contact 22473 2938 22473 2938 6 state[0]
rlabel m2contact 22449 4258 22449 4258 6 n_222
rlabel m2contact 22449 4690 22449 4690 6 n_285
rlabel m2contact 22425 4570 22425 4570 6 n_224
rlabel m2contact 22425 2242 22425 2242 6 n_224
rlabel m2contact 22401 3706 22401 3706 6 n_271
rlabel m2contact 22377 4426 22377 4426 6 n_277
rlabel m2contact 22353 3826 22353 3826 6 n_76
rlabel m2contact 22329 4570 22329 4570 6 n_224
rlabel m2contact 22329 4522 22329 4522 6 n_276
rlabel m2contact 22305 6850 22305 6850 6 n_108
rlabel m2contact 22305 2986 22305 2986 6 n_108
rlabel m2contact 22281 6850 22281 6850 6 n_108
rlabel m2contact 22281 6802 22281 6802 6 n_304
rlabel m2contact 22257 4186 22257 4186 6 n_359
rlabel m2contact 22257 2746 22257 2746 6 n_359
rlabel m2contact 22233 2746 22233 2746 6 n_359
rlabel m2contact 22233 2818 22233 2818 6 n_199
rlabel m2contact 22209 4714 22209 4714 6 n_241
rlabel m2contact 22185 4354 22185 4354 6 n_193
rlabel m2contact 22185 2914 22185 2914 6 n_193
rlabel m2contact 22161 3298 22161 3298 6 OpcodeCondIn[2]
rlabel m2contact 22161 4018 22161 4018 6 n_235
rlabel m2contact 22137 2914 22137 2914 6 n_193
rlabel m2contact 22137 2938 22137 2938 6 state[0]
rlabel m2contact 22113 6082 22113 6082 6 n_182
rlabel m2contact 22113 5146 22113 5146 6 n_203
rlabel m2contact 22065 6418 22065 6418 6 n_40
rlabel m2contact 22017 3538 22017 3538 6 OpcodeCondIn[0]
rlabel m2contact 21993 2674 21993 2674 6 n_336
rlabel m2contact 21993 5482 21993 5482 6 n_12
rlabel m2contact 21957 5578 21957 5578 6 n_301
rlabel m2contact 21957 4258 21957 4258 6 n_301
rlabel m2contact 21945 6754 21945 6754 6 n_257
rlabel m2contact 21921 3706 21921 3706 6 n_271
rlabel m2contact 21897 4258 21897 4258 6 n_301
rlabel m2contact 21897 4498 21897 4498 6 n_210
rlabel m2contact 21873 4234 21873 4234 6 n_15
rlabel m2contact 21849 5410 21849 5410 6 OpcodeCondIn[4]
rlabel m2contact 21849 4258 21849 4258 6 OpcodeCondIn[4]
rlabel m2contact 21825 4474 21825 4474 6 n_229
rlabel m2contact 21825 3226 21825 3226 6 n_59
rlabel m2contact 21801 4354 21801 4354 6 n_193
rlabel m2contact 21777 4258 21777 4258 6 OpcodeCondIn[4]
rlabel m2contact 21777 4306 21777 4306 6 n_194
rlabel m2contact 21753 5386 21753 5386 6 n_310
rlabel m2contact 21753 3058 21753 3058 6 n_310
rlabel m2contact 21729 4090 21729 4090 6 AluEn
rlabel m2contact 21705 5098 21705 5098 6 StatusReg[3]
rlabel m2contact 21681 6658 21681 6658 6 n_159
rlabel m2contact 21681 2650 21681 2650 6 n_289
rlabel m2contact 21657 2938 21657 2938 6 state[0]
rlabel m2contact 21633 2314 21633 2314 6 n_346
rlabel m2contact 21633 6010 21633 6010 6 n_147
rlabel m2contact 21609 4138 21609 4138 6 n_169
rlabel m2contact 21585 4474 21585 4474 6 n_229
rlabel m2contact 21561 4354 21561 4354 6 n_156
rlabel m2contact 21537 6634 21537 6634 6 n_187
rlabel m2contact 21513 4642 21513 4642 6 n_46
rlabel m2contact 21489 6778 21489 6778 6 n_186
rlabel m2contact 21465 5098 21465 5098 6 StatusReg[3]
rlabel m2contact 21441 1762 21441 1762 6 n_267
rlabel m2contact 21417 2914 21417 2914 6 n_351
rlabel m2contact 21417 3346 21417 3346 6 OpcodeCondIn[6]
rlabel m2contact 21393 3946 21393 3946 6 n_207
rlabel m2contact 21369 3058 21369 3058 6 n_310
rlabel m2contact 21369 3082 21369 3082 6 n_217
rlabel m2contact 21321 3130 21321 3130 6 n_243
rlabel m2contact 21297 5794 21297 5794 6 n_356
rlabel m2contact 21297 3994 21297 3994 6 n_356
rlabel m2contact 21273 3994 21273 3994 6 n_356
rlabel m2contact 21273 4138 21273 4138 6 n_169
rlabel m2contact 21249 3946 21249 3946 6 n_207
rlabel m2contact 21249 1954 21249 1954 6 n_258
rlabel m2contact 21213 3778 21213 3778 6 IrWe
rlabel m2contact 21213 1930 21213 1930 6 IrWe
rlabel m2contact 21201 4450 21201 4450 6 n_282
rlabel m2contact 21177 1930 21177 1930 6 IrWe
rlabel m2contact 21177 2050 21177 2050 6 n_264
rlabel m2contact 21153 4258 21153 4258 6 n_280
rlabel m2contact 21129 6274 21129 6274 6 n_115
rlabel m2contact 21081 4066 21081 4066 6 n_213
rlabel m2contact 21081 5914 21081 5914 6 n_89
rlabel m2contact 21033 6538 21033 6538 6 n_222
rlabel m2contact 21009 2266 21009 2266 6 n_116
rlabel m2contact 20913 2986 20913 2986 6 n_108
rlabel m2contact 20913 2746 20913 2746 6 n_108
rlabel m2contact 20889 2746 20889 2746 6 n_108
rlabel m2contact 20889 2866 20889 2866 6 StatusReg[0]
rlabel m2contact 20865 5002 20865 5002 6 n_119
rlabel m2contact 20841 6370 20841 6370 6 n_478
rlabel m2contact 20817 4090 20817 4090 6 AluEn
rlabel m2contact 20793 3874 20793 3874 6 n_354
rlabel m2contact 20769 4162 20769 4162 6 n_368
rlabel m2contact 20721 4090 20721 4090 6 n_27
rlabel m2contact 20697 5746 20697 5746 6 stateSub[1]
rlabel m2contact 20673 3922 20673 3922 6 n_99
rlabel m2contact 20625 5266 20625 5266 6 n_29
rlabel m2contact 20601 5410 20601 5410 6 OpcodeCondIn[4]
rlabel m2contact 20577 4810 20577 4810 6 n_58
rlabel m2contact 20553 3346 20553 3346 6 OpcodeCondIn[6]
rlabel m2contact 20505 6922 20505 6922 6 n_366
rlabel m2contact 20505 4450 20505 4450 6 n_366
rlabel m2contact 20481 6922 20481 6922 6 n_366
rlabel m2contact 20481 6874 20481 6874 6 n_153
rlabel m2contact 20457 4066 20457 4066 6 n_252
rlabel m2contact 20409 6610 20409 6610 6 n_145
rlabel m2contact 20385 2818 20385 2818 6 n_199
rlabel m2contact 20361 4306 20361 4306 6 n_194
rlabel m2contact 20337 2746 20337 2746 6 n_3
rlabel m2contact 20337 2386 20337 2386 6 n_134
rlabel m2contact 20313 4906 20313 4906 6 n_68
rlabel m2contact 20313 2770 20313 2770 6 n_68
rlabel m2contact 20289 2026 20289 2026 6 n_93
rlabel m2contact 20289 3754 20289 3754 6 nIRQ
rlabel m2contact 20265 4762 20265 4762 6 OpcodeCondIn[7]
rlabel m2contact 20241 4546 20241 4546 6 n_262
rlabel m2contact 20241 3178 20241 3178 6 n_176
rlabel m2contact 20217 3658 20217 3658 6 n_28
rlabel m2contact 20193 3130 20193 3130 6 n_243
rlabel m2contact 20169 3730 20169 3730 6 stateSub[0]
rlabel m2contact 20145 5290 20145 5290 6 n_231
rlabel m2contact 20121 4450 20121 4450 6 n_366
rlabel m2contact 20121 2362 20121 2362 6 n_300
rlabel m2contact 20097 4426 20097 4426 6 n_277
rlabel m2contact 20073 5458 20073 5458 6 n_190
rlabel m2contact 20073 6226 20073 6226 6 n_338
rlabel m2contact 20049 4594 20049 4594 6 n_292
rlabel m2contact 20049 4570 20049 4570 6 n_73
rlabel m2contact 20025 2098 20025 2098 6 n_189
rlabel m2contact 20001 5338 20001 5338 6 n_52
rlabel m2contact 19977 4906 19977 4906 6 n_68
rlabel m2contact 19977 4882 19977 4882 6 n_126
rlabel m2contact 19953 3418 19953 3418 6 n_51
rlabel m2contact 19929 4930 19929 4930 6 n_123
rlabel m2contact 19905 4426 19905 4426 6 n_93
rlabel m2contact 19905 2026 19905 2026 6 n_93
rlabel m2contact 19881 3250 19881 3250 6 n_65
rlabel m2contact 19857 3586 19857 3586 6 n_177
rlabel m2contact 19833 4426 19833 4426 6 n_93
rlabel m2contact 19833 4138 19833 4138 6 n_169
rlabel m2contact 19809 3922 19809 3922 6 n_99
rlabel m2contact 19785 5962 19785 5962 6 n_274
rlabel metal2 19761 4162 19761 4162 6 SysBus[2]
rlabel m2contact 19737 4522 19737 4522 6 n_276
rlabel m2contact 19689 5434 19689 5434 6 n_38
rlabel m2contact 19641 3226 19641 3226 6 n_59
rlabel m2contact 19617 2026 19617 2026 6 n_93
rlabel m2contact 19545 4834 19545 4834 6 n_172
rlabel m2contact 19497 2506 19497 2506 6 n_30
rlabel m2contact 19425 6250 19425 6250 6 n_138
rlabel m2contact 19377 4162 19377 4162 6 n_137
rlabel m2contact 19329 2434 19329 2434 6 n_82
rlabel m2contact 19305 6730 19305 6730 6 n_9
rlabel m2contact 19281 5194 19281 5194 6 n_49
rlabel m2contact 19233 6202 19233 6202 6 n_103
rlabel m2contact 19209 2746 19209 2746 6 n_3
rlabel m2contact 19209 2986 19209 2986 6 n_108
rlabel m2contact 19185 5746 19185 5746 6 stateSub[1]
rlabel m2contact 19161 4426 19161 4426 6 n_176
rlabel m2contact 19161 3178 19161 3178 6 n_176
rlabel m2contact 19137 3658 19137 3658 6 n_28
rlabel m2contact 19113 3322 19113 3322 6 OpcodeCondIn[3]
rlabel m2contact 19089 4426 19089 4426 6 n_176
rlabel m2contact 19089 3562 19089 3562 6 n_21
rlabel m2contact 19053 5722 19053 5722 6 n_10
rlabel m2contact 19053 3994 19053 3994 6 n_10
rlabel m2contact 19041 5818 19041 5818 6 n_13
rlabel m2contact 19041 3082 19041 3082 6 n_217
rlabel m2contact 19017 3994 19017 3994 6 n_10
rlabel m2contact 19017 4762 19017 4762 6 OpcodeCondIn[7]
rlabel m2contact 18993 5482 18993 5482 6 n_12
rlabel m2contact 18957 4426 18957 4426 6 n_93
rlabel m2contact 18957 2026 18957 2026 6 n_93
rlabel m2contact 18945 6130 18945 6130 6 n_233
rlabel m2contact 18921 3466 18921 3466 6 n_195
rlabel m2contact 18897 4402 18897 4402 6 n_196
rlabel m2contact 18861 5746 18861 5746 6 stateSub[1]
rlabel m2contact 18861 3610 18861 3610 6 stateSub[1]
rlabel m2contact 18849 3106 18849 3106 6 n_228
rlabel m2contact 18825 3994 18825 3994 6 n_33
rlabel m2contact 18801 2410 18801 2410 6 stateSub[2]
rlabel m2contact 18777 2002 18777 2002 6 n_32
rlabel m2contact 18753 4786 18753 4786 6 n_62
rlabel m2contact 18729 3610 18729 3610 6 stateSub[1]
rlabel m2contact 18729 4402 18729 4402 6 n_104
rlabel m2contact 18705 4426 18705 4426 6 n_93
rlabel m2contact 18705 3634 18705 3634 6 n_31
rlabel m2contact 18681 3418 18681 3418 6 n_51
rlabel m2contact 18657 2194 18657 2194 6 n_358
rlabel m2contact 18657 2770 18657 2770 6 n_68
rlabel m2contact 18633 5218 18633 5218 6 n_347
rlabel m2contact 18633 3610 18633 3610 6 n_347
rlabel m2contact 18609 4330 18609 4330 6 n_251
rlabel m2contact 18609 4546 18609 4546 6 n_325
rlabel m2contact 18585 3610 18585 3610 6 n_347
rlabel m2contact 18585 3850 18585 3850 6 state[1]
rlabel m2contact 18561 5914 18561 5914 6 n_89
rlabel m2contact 18537 4114 18537 4114 6 n_84
rlabel m2contact 18513 4330 18513 4330 6 n_254
rlabel m2contact 18489 4378 18489 4378 6 n_34
rlabel m2contact 18465 3658 18465 3658 6 n_28
rlabel m2contact 18441 3298 18441 3298 6 OpcodeCondIn[2]
rlabel m2contact 18417 5506 18417 5506 6 n_39
rlabel m2contact 18417 4666 18417 4666 6 n_278
rlabel m2contact 18369 3922 18369 3922 6 n_99
rlabel m2contact 18345 4186 18345 4186 6 n_359
rlabel m2contact 18345 3610 18345 3610 6 n_107
rlabel m2contact 18309 4378 18309 4378 6 n_264
rlabel m2contact 18309 2050 18309 2050 6 n_264
rlabel m2contact 18297 5362 18297 5362 6 n_260
rlabel m2contact 18273 5050 18273 5050 6 n_283
rlabel m2contact 18249 4906 18249 4906 6 n_80
rlabel m2contact 18225 4834 18225 4834 6 n_172
rlabel m2contact 18225 3154 18225 3154 6 n_237
rlabel m2contact 18201 4930 18201 4930 6 n_123
rlabel m2contact 18177 4378 18177 4378 6 n_264
rlabel m2contact 18177 3466 18177 3466 6 n_195
rlabel m2contact 18153 3178 18153 3178 6 n_176
rlabel m2contact 18129 5530 18129 5530 6 n_26
rlabel m2contact 18129 4282 18129 4282 6 n_155
rlabel m2contact 18105 3082 18105 3082 6 n_217
rlabel m2contact 18081 5746 18081 5746 6 stateSub[1]
rlabel m2contact 18057 3586 18057 3586 6 n_177
rlabel m2contact 18033 2050 18033 2050 6 n_264
rlabel m2contact 18009 3322 18009 3322 6 OpcodeCondIn[3]
rlabel m2contact 17985 3322 17985 3322 6 OpcodeCondIn[3]
rlabel m2contact 17961 3346 17961 3346 6 OpcodeCondIn[6]
rlabel m2contact 17937 2554 17937 2554 6 n_100
rlabel m2contact 17913 6514 17913 6514 6 n_334
rlabel m2contact 17889 5938 17889 5938 6 n_112
rlabel m2contact 17889 3010 17889 3010 6 n_112
rlabel m2contact 17865 2674 17865 2674 6 n_336
rlabel m2contact 17829 4450 17829 4450 6 n_134
rlabel m2contact 17829 2386 17829 2386 6 n_134
rlabel m2contact 17817 4594 17817 4594 6 n_136
rlabel m2contact 17793 4450 17793 4450 6 n_134
rlabel m2contact 17793 4426 17793 4426 6 OpcodeCondIn[5]
rlabel m2contact 17769 2938 17769 2938 6 state[0]
rlabel m2contact 17745 4450 17745 4450 6 n_273
rlabel m2contact 17745 6058 17745 6058 6 n_135
rlabel m2contact 17721 1906 17721 1906 6 n_96
rlabel m2contact 17697 6466 17697 6466 6 PcEn
rlabel m2contact 17697 4066 17697 4066 6 n_252
rlabel m2contact 17661 3130 17661 3130 6 n_243
rlabel m2contact 17661 2722 17661 2722 6 n_243
rlabel m2contact 17649 4978 17649 4978 6 n_141
rlabel m2contact 17625 4858 17625 4858 6 n_74
rlabel m2contact 17625 3922 17625 3922 6 n_99
rlabel m2contact 17601 2722 17601 2722 6 n_243
rlabel m2contact 17601 2746 17601 2746 6 n_132
rlabel m2contact 17577 4378 17577 4378 6 n_61
rlabel m2contact 17553 5650 17553 5650 6 Flags[2]
rlabel m2contact 17553 2170 17553 2170 6 Flags[2]
rlabel m2contact 17529 3010 17529 3010 6 n_112
rlabel m2contact 17529 3058 17529 3058 6 n_246
rlabel m2contact 17505 3034 17505 3034 6 n_6
rlabel m2contact 17481 3658 17481 3658 6 n_167
rlabel m2contact 17457 1858 17457 1858 6 n_245
rlabel m2contact 17433 3418 17433 3418 6 n_51
rlabel m2contact 17409 6442 17409 6442 6 n_279
rlabel m2contact 17409 5410 17409 5410 6 OpcodeCondIn[4]
rlabel m2contact 17385 4810 17385 4810 6 n_58
rlabel m2contact 17361 4666 17361 4666 6 n_278
rlabel m2contact 17337 6130 17337 6130 6 n_233
rlabel m2contact 17313 4426 17313 4426 6 OpcodeCondIn[5]
rlabel m2contact 17289 5650 17289 5650 6 Flags[2]
rlabel m2contact 17289 3082 17289 3082 6 n_217
rlabel m2contact 16737 5650 16737 5650 6 n_365
rlabel m2contact 16641 6130 16641 6130 6 n_185
rlabel m2contact 16641 1810 16641 1810 6 n_185
rlabel m2contact 16617 6130 16617 6130 6 n_185
rlabel m2contact 16617 2482 16617 2482 6 n_335
rlabel m2contact 16593 2170 16593 2170 6 Flags[2]
rlabel m2contact 16593 2410 16593 2410 6 stateSub[2]
rlabel m2contact 16569 6034 16569 6034 6 n_180
rlabel m2contact 16569 2674 16569 2674 6 n_336
rlabel m2contact 16545 6442 16545 6442 6 n_166
rlabel m2contact 16521 3490 16521 3490 6 n_209
rlabel m2contact 16497 5890 16497 5890 6 n_332
rlabel m2contact 16497 2050 16497 2050 6 n_264
rlabel m2contact 16473 5554 16473 5554 6 n_35
rlabel m2contact 16473 3946 16473 3946 6 n_207
rlabel m2contact 16449 5890 16449 5890 6 n_295
rlabel m2contact 16449 4210 16449 4210 6 n_208
rlabel m2contact 16425 4786 16425 4786 6 n_62
rlabel m2contact 16425 4498 16425 4498 6 n_210
rlabel m2contact 16401 3370 16401 3370 6 n_72
rlabel m2contact 16377 6754 16377 6754 6 n_257
rlabel m2contact 16377 3490 16377 3490 6 n_257
rlabel m2contact 16353 6034 16353 6034 6 stateSub[2]
rlabel m2contact 16353 2410 16353 2410 6 stateSub[2]
rlabel m2contact 16329 5458 16329 5458 6 n_190
rlabel m2contact 16305 4786 16305 4786 6 n_324
rlabel m2contact 16305 3418 16305 3418 6 n_220
rlabel m2contact 16281 5458 16281 5458 6 n_255
rlabel m2contact 16257 3370 16257 3370 6 n_72
rlabel m2contact 16233 3826 16233 3826 6 n_76
rlabel m2contact 16233 3730 16233 3730 6 stateSub[0]
rlabel m2contact 16209 5914 16209 5914 6 n_89
rlabel m2contact 16185 5746 16185 5746 6 stateSub[1]
rlabel m2contact 16161 6538 16161 6538 6 n_222
rlabel m2contact 16137 4762 16137 4762 6 OpcodeCondIn[7]
rlabel m2contact 16113 5554 16113 5554 6 n_86
rlabel m2contact 16113 4738 16113 4738 6 n_201
rlabel m2contact 16089 3490 16089 3490 6 n_257
rlabel m2contact 16089 6586 16089 6586 6 n_36
rlabel m2contact 16065 6034 16065 6034 6 stateSub[2]
rlabel m2contact 16065 3322 16065 3322 6 OpcodeCondIn[3]
rlabel m2contact 16041 6754 16041 6754 6 n_257
rlabel m2contact 16041 2170 16041 2170 6 n_257
rlabel m2contact 16017 4042 16017 4042 6 Op1Sel
rlabel m2contact 16017 5770 16017 5770 6 AluOR[0]
rlabel m2contact 15993 5794 15993 5794 6 n_356
rlabel m2contact 15969 2170 15969 2170 6 n_257
rlabel m2contact 15969 2338 15969 2338 6 n_343
rlabel m2contact 15945 4450 15945 4450 6 n_273
rlabel m2contact 15921 5194 15921 5194 6 n_49
rlabel m2contact 15897 4810 15897 4810 6 n_58
rlabel m2contact 15873 2506 15873 2506 6 n_30
rlabel m2contact 15849 4138 15849 4138 6 n_169
rlabel m2contact 15825 4330 15825 4330 6 n_254
rlabel m2contact 15825 3010 15825 3010 6 n_254
rlabel m2contact 15801 3178 15801 3178 6 n_176
rlabel m2contact 15777 5194 15777 5194 6 stateSub[2]
rlabel m2contact 15777 2410 15777 2410 6 stateSub[2]
rlabel m2contact 15753 3010 15753 3010 6 n_254
rlabel m2contact 15753 3346 15753 3346 6 OpcodeCondIn[6]
rlabel m2contact 15729 3130 15729 3130 6 n_243
rlabel m2contact 15705 5698 15705 5698 6 n_219
rlabel m2contact 15681 5626 15681 5626 6 n_173
rlabel m2contact 15681 2122 15681 2122 6 n_162
rlabel m2contact 15657 2722 15657 2722 6 n_161
rlabel m2contact 15657 4042 15657 4042 6 n_218
rlabel m2contact 15633 2410 15633 2410 6 stateSub[2]
rlabel m2contact 15609 2170 15609 2170 6 n_85
rlabel m2contact 15585 6490 15585 6490 6 MemEn
rlabel m2contact 15585 3490 15585 3490 6 MemEn
rlabel m2contact 15561 5194 15561 5194 6 stateSub[2]
rlabel m2contact 15561 2938 15561 2938 6 state[0]
rlabel m2contact 15537 5242 15537 5242 6 n_45
rlabel m2contact 15537 2242 15537 2242 6 n_224
rlabel m2contact 15513 5194 15513 5194 6 n_16
rlabel m2contact 15513 3274 15513 3274 6 n_16
rlabel m2contact 15489 3490 15489 3490 6 MemEn
rlabel m2contact 15489 5698 15489 5698 6 n_121
rlabel m2contact 15465 5002 15465 5002 6 n_119
rlabel m2contact 15441 4930 15441 4930 6 n_123
rlabel m2contact 15441 3490 15441 3490 6 n_266
rlabel m2contact 15417 5002 15417 5002 6 n_232
rlabel m2contact 15393 6850 15393 6850 6 n_212
rlabel m2contact 15369 3010 15369 3010 6 n_109
rlabel m2contact 15369 3346 15369 3346 6 OpcodeCondIn[6]
rlabel m2contact 15345 1882 15345 1882 6 n_106
rlabel m2contact 15345 3370 15345 3370 6 n_214
rlabel m2contact 15321 5194 15321 5194 6 n_16
rlabel m2contact 15321 3610 15321 3610 6 n_107
rlabel m2contact 15297 2986 15297 2986 6 n_108
rlabel m2contact 15225 6010 15225 6010 6 n_147
rlabel m2contact 15225 3730 15225 3730 6 stateSub[0]
rlabel m2contact 15201 5938 15201 5938 6 n_112
rlabel m2contact 15201 5770 15201 5770 6 n_11
rlabel m2contact 15129 4546 15129 4546 6 n_325
rlabel m2contact 15105 2578 15105 2578 6 n_268
rlabel m2contact 15105 2986 15105 2986 6 n_329
rlabel m2contact 15081 2074 15081 2074 6 n_294
rlabel m2contact 15033 1930 15033 1930 6 n_144
rlabel m2contact 14985 3394 14985 3394 6 n_269
rlabel m2contact 14961 3154 14961 3154 6 n_237
rlabel m2contact 14913 3514 14913 3514 6 n_227
rlabel m2contact 14889 4570 14889 4570 6 n_73
rlabel m2contact 14889 3226 14889 3226 6 n_59
rlabel m2contact 14865 4066 14865 4066 6 n_252
rlabel m2contact 14841 6154 14841 6154 6 n_94
rlabel m2contact 14817 2818 14817 2818 6 n_199
rlabel m2contact 14793 2578 14793 2578 6 LrWe
rlabel m2contact 14769 3514 14769 3514 6 OpcodeCondIn[1]
rlabel m2contact 14745 3538 14745 3538 6 OpcodeCondIn[0]
rlabel m2contact 14721 5194 14721 5194 6 stateSub[2]
rlabel m2contact 14721 2410 14721 2410 6 stateSub[2]
rlabel m2contact 14697 2770 14697 2770 6 n_68
rlabel m2contact 14673 5410 14673 5410 6 OpcodeCondIn[4]
rlabel m2contact 14649 5194 14649 5194 6 stateSub[2]
rlabel m2contact 14649 3586 14649 3586 6 n_177
rlabel m2contact 14625 5242 14625 5242 6 n_242
rlabel m2contact 14625 4570 14625 4570 6 n_242
rlabel m2contact 14601 4570 14601 4570 6 n_242
rlabel m2contact 14601 4930 14601 4930 6 n_123
rlabel m2contact 14577 3730 14577 3730 6 stateSub[0]
rlabel m2contact 14553 3130 14553 3130 6 n_243
rlabel m2contact 14505 4570 14505 4570 6 n_206
rlabel m2contact 14481 4666 14481 4666 6 n_278
rlabel m2contact 14457 6778 14457 6778 6 n_186
rlabel m2contact 14409 3130 14409 3130 6 n_188
rlabel m2contact 14385 4618 14385 4618 6 n_37
rlabel m2contact 14361 2098 14361 2098 6 n_189
rlabel m2contact 14289 4834 14289 4834 6 n_172
rlabel m2contact 14265 3586 14265 3586 6 n_177
rlabel m2contact 14241 1882 14241 1882 6 n_106
rlabel m2contact 14241 4618 14241 4618 6 n_286
rlabel m2contact 14193 2578 14193 2578 6 LrWe
rlabel m2contact 14145 2602 14145 2602 6 n_316
rlabel m2contact 14121 5938 14121 5938 6 n_290
rlabel m2contact 14097 2578 14097 2578 6 n_275
rlabel m2contact 14073 2650 14073 2650 6 n_289
rlabel m2contact 14049 4522 14049 4522 6 n_276
rlabel m2contact 14001 4162 14001 4162 6 n_137
rlabel m2contact 13953 6562 13953 6562 6 n_20
rlabel m2contact 13929 2170 13929 2170 6 n_85
rlabel m2contact 13929 5098 13929 5098 6 StatusReg[3]
rlabel m2contact 13881 2602 13881 2602 6 n_316
rlabel m2contact 13881 5626 13881 5626 6 n_479
rlabel m2contact 13857 4714 13857 4714 6 n_241
rlabel m2contact 13833 6130 13833 6130 6 n_302
rlabel m2contact 13713 5098 13713 5098 6 n_299
rlabel m2contact 13665 3658 13665 3658 6 n_167
rlabel m2contact 13641 3082 13641 3082 6 n_217
rlabel m2contact 13593 5194 13593 5194 6 n_361
rlabel m2contact 13593 2170 13593 2170 6 n_361
rlabel m2contact 13569 5794 13569 5794 4 n_356
rlabel m2contact 13545 3850 13545 3850 4 state[1]
rlabel m2contact 13521 5194 13521 5194 4 n_361
rlabel m2contact 13521 4114 13521 4114 4 n_84
rlabel m2contact 13497 2410 13497 2410 4 stateSub[2]
rlabel m2contact 13449 5194 13449 5194 4 n_189
rlabel m2contact 13449 2098 13449 2098 4 n_189
rlabel m2contact 13425 3658 13425 3658 4 nOE
rlabel m2contact 13401 5002 13401 5002 4 n_232
rlabel m2contact 13401 2602 13401 2602 4 n_71
rlabel m2contact 13377 1978 13377 1978 4 n_179
rlabel m2contact 13377 5290 13377 5290 4 n_231
rlabel m2contact 13353 1762 13353 1762 4 n_267
rlabel m2contact 13353 3418 13353 3418 4 n_220
rlabel m2contact 13329 6034 13329 6034 4 n_77
rlabel m2contact 13329 1978 13329 1978 4 n_77
rlabel m2contact 13305 5002 13305 5002 4 n_191
rlabel m2contact 13281 5338 13281 5338 4 n_52
rlabel m2contact 13257 5194 13257 5194 4 n_189
rlabel m2contact 13257 3298 13257 3298 4 OpcodeCondIn[2]
rlabel m2contact 13233 4930 13233 4930 4 n_123
rlabel m2contact 13209 4954 13209 4954 4 n_24
rlabel m2contact 13209 2818 13209 2818 4 n_199
rlabel m2contact 13185 3922 13185 3922 4 n_99
rlabel m2contact 13161 4138 13161 4138 4 n_169
rlabel m2contact 13137 2410 13137 2410 4 stateSub[2]
rlabel m2contact 13113 4954 13113 4954 4 n_211
rlabel m2contact 13113 4090 13113 4090 4 n_27
rlabel m2contact 13089 3682 13089 3682 4 nWait
rlabel m2contact 13065 1978 13065 1978 4 n_77
rlabel m2contact 13065 3370 13065 3370 4 n_214
rlabel m2contact 13041 4330 13041 4330 4 n_254
rlabel m2contact 13017 4498 13017 4498 4 n_210
rlabel m2contact 12969 1978 12969 1978 4 n_312
rlabel m2contact 12945 3322 12945 3322 4 OpcodeCondIn[3]
rlabel m2contact 12921 6802 12921 6802 4 n_304
rlabel m2contact 12873 4258 12873 4258 4 n_280
rlabel m2contact 12825 4714 12825 4714 4 n_241
rlabel m2contact 12801 3970 12801 3970 4 n_250
rlabel m2contact 12729 3874 12729 3874 4 n_354
rlabel m2contact 12705 5338 12705 5338 4 n_323
rlabel m2contact 12681 5194 12681 5194 4 n_355
rlabel m2contact 12657 5794 12657 5794 4 n_356
rlabel m2contact 12585 5794 12585 5794 4 n_113
rlabel m2contact 12537 6826 12537 6826 4 n_98
rlabel m2contact 12489 6442 12489 6442 4 n_166
rlabel m2contact 12465 3082 12465 3082 4 n_217
rlabel m2contact 12441 4594 12441 4594 4 n_136
rlabel m2contact 12369 6130 12369 6130 4 n_302
rlabel m2contact 12345 6922 12345 6922 4 stateSub[2]
rlabel m2contact 12345 2410 12345 2410 4 stateSub[2]
rlabel m2contact 12321 4450 12321 4450 4 n_273
rlabel m2contact 12297 1810 12297 1810 4 n_185
rlabel m2contact 12261 6826 12261 6826 4 n_67
rlabel m2contact 12261 2530 12261 2530 4 n_67
rlabel m2contact 12249 2002 12249 2002 4 n_32
rlabel m2contact 12225 4930 12225 4930 4 n_123
rlabel m2contact 12201 3898 12201 3898 4 n_319
rlabel m2contact 12177 6442 12177 6442 4 n_160
rlabel m2contact 12177 2002 12177 2002 4 n_160
rlabel m2contact 12153 4594 12153 4594 4 n_236
rlabel m2contact 12129 6922 12129 6922 4 stateSub[2]
rlabel m2contact 12129 4450 12129 4450 4 n_105
rlabel m2contact 12105 6898 12105 6898 4 n_181
rlabel m2contact 12105 2410 12105 2410 4 stateSub[2]
rlabel m2contact 12081 5410 12081 5410 4 OpcodeCondIn[4]
rlabel m2contact 12081 1810 12081 1810 4 OpcodeCondIn[4]
rlabel m2contact 12057 6874 12057 6874 4 n_153
rlabel m2contact 12057 4042 12057 4042 4 n_218
rlabel m2contact 12033 6826 12033 6826 4 n_67
rlabel m2contact 12033 4426 12033 4426 4 OpcodeCondIn[5]
rlabel m2contact 12009 6706 12009 6706 4 n_117
rlabel m2contact 12009 5986 12009 5986 4 n_174
rlabel m2contact 11985 5266 11985 5266 4 n_29
rlabel m2contact 11961 6154 11961 6154 4 n_94
rlabel m2contact 11937 1810 11937 1810 4 OpcodeCondIn[4]
rlabel m2contact 11913 6442 11913 6442 4 n_160
rlabel m2contact 11913 3082 11913 3082 4 n_217
rlabel m2contact 11889 5266 11889 5266 4 n_8
rlabel m2contact 11865 5314 11865 5314 4 n_122
rlabel m2contact 11841 6826 11841 6826 4 n_53
rlabel m2contact 11817 6442 11817 6442 4 n_64
rlabel m2contact 11817 2842 11817 2842 4 n_256
rlabel m2contact 11793 4258 11793 4258 4 n_280
rlabel m2contact 11769 5314 11769 5314 4 n_314
rlabel m2contact 11745 1786 11745 1786 4 n_81
rlabel m2contact 11745 5242 11745 5242 4 n_242
rlabel m2contact 11721 1810 11721 1810 4 OpcodeCondIn[4]
rlabel m2contact 11721 4258 11721 4258 4 n_261
rlabel m2contact 11697 6850 11697 6850 4 n_212
rlabel m2contact 11697 6706 11697 6706 4 n_41
rlabel m2contact 11673 5242 11673 5242 4 n_341
rlabel m2contact 11673 1810 11673 1810 4 n_341
rlabel m2contact 11649 2626 11649 2626 4 RwSel[0]
rlabel m2contact 11649 6226 11649 6226 4 n_338
rlabel m2contact 11625 5746 11625 5746 4 stateSub[1]
rlabel m2contact 11601 2674 11601 2674 4 n_336
rlabel m2contact 11577 4162 11577 4162 4 n_137
rlabel m2contact 11553 3898 11553 3898 4 n_319
rlabel m2contact 11529 5482 11529 5482 4 n_12
rlabel m2contact 11505 2626 11505 2626 4 ImmSel
rlabel m2contact 11481 1810 11481 1810 4 n_341
rlabel m2contact 11481 3514 11481 3514 4 OpcodeCondIn[1]
rlabel m2contact 11457 6226 11457 6226 4 n_305
rlabel m2contact 11433 6826 11433 6826 4 n_53
rlabel m2contact 11433 4162 11433 4162 4 n_67
rlabel m2contact 11433 2530 11433 2530 4 n_67
rlabel m2contact 11409 3298 11409 3298 4 OpcodeCondIn[2]
rlabel m2contact 11385 6370 11385 6370 4 n_478
rlabel m2contact 11361 3946 11361 3946 4 n_207
rlabel m2contact 11361 5506 11361 5506 4 n_39
rlabel m2contact 11337 6370 11337 6370 4 OpcodeCondIn[3]
rlabel m2contact 11337 3322 11337 3322 4 OpcodeCondIn[3]
rlabel m2contact 11313 4162 11313 4162 4 n_67
rlabel m2contact 11313 2938 11313 2938 4 state[0]
rlabel m2contact 11289 6370 11289 6370 4 OpcodeCondIn[3]
rlabel m2contact 11289 4282 11289 4282 4 n_155
rlabel m2contact 11265 1882 11265 1882 4 n_106
rlabel m2contact 11241 6538 11241 6538 4 n_222
rlabel m2contact 11217 3370 11217 3370 4 n_214
rlabel m2contact 11193 4930 11193 4930 4 n_123
rlabel m2contact 11169 4282 11169 4282 4 n_155
rlabel m2contact 11145 5146 11145 5146 4 n_203
rlabel m2contact 11097 4210 11097 4210 4 n_208
rlabel m2contact 11097 4162 11097 4162 4 n_50
rlabel m2contact 11073 6538 11073 6538 4 n_222
rlabel m2contact 11049 3850 11049 3850 4 state[1]
rlabel m2contact 11025 3922 11025 3922 4 n_99
rlabel m2contact 11001 3946 11001 3946 4 n_226
rlabel m2contact 10977 1834 10977 1834 4 n_259
rlabel m2contact 10977 6370 10977 6370 4 n_90
rlabel m2contact 10953 5914 10953 5914 4 n_89
rlabel m2contact 10929 4666 10929 4666 4 n_278
rlabel m2contact 10905 1858 10905 1858 4 n_245
rlabel m2contact 10881 2938 10881 2938 4 state[0]
rlabel m2contact 10857 6226 10857 6226 4 n_305
rlabel m2contact 10833 3922 10833 3922 4 n_99
rlabel m2contact 10809 6802 10809 6802 4 n_304
rlabel m2contact 10809 3082 10809 3082 4 n_217
rlabel m2contact 10785 6226 10785 6226 4 n_263
rlabel m2contact 10785 1858 10785 1858 4 n_263
rlabel m2contact 10761 5578 10761 5578 4 n_301
rlabel m2contact 10737 1858 10737 1858 4 n_263
rlabel m2contact 10737 3082 10737 3082 4 n_217
rlabel m2contact 10713 2362 10713 2362 4 n_300
rlabel m2contact 10689 5578 10689 5578 4 n_171
rlabel m2contact 10665 2362 10665 2362 4 n_265
rlabel m2contact 10641 2050 10641 2050 4 n_264
rlabel m2contact 10617 1906 10617 1906 4 n_96
rlabel m2contact 10617 5362 10617 5362 4 n_260
rlabel m2contact 10569 1882 10569 1882 4 n_106
rlabel m2contact 10569 6778 10569 6778 4 n_186
rlabel m2contact 10569 5842 10569 5842 4 n_56
rlabel m2contact 10569 1906 10569 1906 4 n_56
rlabel m2contact 10545 1906 10545 1906 4 n_56
rlabel m2contact 10545 2938 10545 2938 4 state[0]
rlabel m2contact 10521 1930 10521 1930 4 n_144
rlabel m2contact 10473 1954 10473 1954 4 n_258
rlabel m2contact 10449 2842 10449 2842 4 n_256
rlabel m2contact 10425 3970 10425 3970 4 n_250
rlabel m2contact 10401 6754 10401 6754 4 n_257
rlabel m2contact 10353 6730 10353 6730 4 n_9
rlabel m2contact 10329 5410 10329 5410 4 OpcodeCondIn[4]
rlabel m2contact 10305 3178 10305 3178 4 n_176
rlabel m2contact 10257 2626 10257 2626 4 ImmSel
rlabel m2contact 10233 4138 10233 4138 4 n_169
rlabel m2contact 10209 5674 10209 5674 4 n_48
rlabel m2contact 10209 4282 10209 4282 4 n_155
rlabel m2contact 10185 4642 10185 4642 4 n_46
rlabel m2contact 10161 2626 10161 2626 4 n_83
rlabel m2contact 10161 5674 10161 5674 4 n_47
rlabel m2contact 10113 6706 10113 6706 4 n_41
rlabel m2contact 10113 5434 10113 5434 4 n_38
rlabel m2contact 10089 4498 10089 4498 4 n_210
rlabel m2contact 10065 6418 10065 6418 4 n_40
rlabel m2contact 10017 4378 10017 4378 4 n_61
rlabel m2contact 9993 3346 9993 3346 4 OpcodeCondIn[6]
rlabel m2contact 9969 3058 9969 3058 4 n_246
rlabel m2contact 9969 3586 9969 3586 4 n_177
rlabel m2contact 9945 4834 9945 4834 4 n_172
rlabel m2contact 9897 3058 9897 3058 4 n_88
rlabel m2contact 9897 2698 9897 2698 4 n_139
rlabel m2contact 9873 2410 9873 2410 4 stateSub[2]
rlabel m2contact 9873 3850 9873 3850 4 state[1]
rlabel m2contact 9849 4378 9849 4378 4 n_87
rlabel m2contact 9801 2674 9801 2674 4 n_336
rlabel m2contact 9777 1978 9777 1978 4 n_312
rlabel m2contact 9777 2410 9777 2410 4 n_175
rlabel m2contact 9753 5434 9753 5434 4 n_253
rlabel m2contact 9729 3130 9729 3130 4 n_188
rlabel m2contact 9705 4714 9705 4714 4 n_241
rlabel m2contact 9681 6682 9681 6682 4 n_291
rlabel m2contact 9681 5146 9681 5146 4 n_203
rlabel m2contact 9657 3586 9657 3586 4 n_177
rlabel m2contact 9633 5050 9633 5050 4 n_283
rlabel m2contact 9561 4810 9561 4810 4 n_58
rlabel m2contact 9537 6682 9537 6682 4 state[0]
rlabel m2contact 9537 2938 9537 2938 4 state[0]
rlabel m2contact 9513 4762 9513 4762 4 OpcodeCondIn[7]
rlabel m2contact 9513 3130 9513 3130 4 n_303
rlabel m2contact 9489 6130 9489 6130 4 n_302
rlabel m2contact 9465 2002 9465 2002 4 n_160
rlabel m2contact 9465 3898 9465 3898 4 n_319
rlabel m2contact 9441 3850 9441 3850 4 state[1]
rlabel m2contact 9417 6682 9417 6682 4 state[0]
rlabel m2contact 9417 5050 9417 5050 4 n_129
rlabel m2contact 9393 2026 9393 2026 4 n_93
rlabel m2contact 9369 3778 9369 3778 4 IrWe
rlabel m2contact 9321 5866 9321 5866 4 n_165
rlabel m2contact 9321 3778 9321 3778 4 n_69
rlabel m2contact 9297 2722 9297 2722 4 n_161
rlabel m2contact 9273 2050 9273 2050 4 n_264
rlabel m2contact 9273 3082 9273 3082 4 n_217
rlabel m2contact 9249 4810 9249 4810 4 n_58
rlabel m2contact 9225 5194 9225 5194 4 n_355
rlabel m2contact 9177 6658 9177 6658 4 n_159
rlabel m2contact 9177 5866 9177 5866 4 n_100
rlabel m2contact 9177 2554 9177 2554 4 n_100
rlabel m2contact 9153 6610 9153 6610 4 n_145
rlabel m2contact 9153 3202 9153 3202 4 n_97
rlabel m2contact 9129 4066 9129 4066 4 n_252
rlabel m2contact 9105 2746 9105 2746 4 n_132
rlabel m2contact 9081 2074 9081 2074 4 n_294
rlabel m2contact 9081 5410 9081 5410 4 OpcodeCondIn[4]
rlabel m2contact 9057 5866 9057 5866 4 n_100
rlabel m2contact 9057 3730 9057 3730 4 stateSub[0]
rlabel m2contact 9009 5866 9009 5866 4 n_230
rlabel m2contact 9009 5146 9009 5146 4 n_203
rlabel m2contact 8985 2122 8985 2122 4 n_162
rlabel m2contact 8961 6634 8961 6634 4 n_187
rlabel m2contact 8961 2098 8961 2098 4 n_189
rlabel m2contact 8961 6610 8961 6610 4 n_87
rlabel m2contact 8961 4378 8961 4378 4 n_87
rlabel m2contact 8937 6298 8937 6298 4 n_158
rlabel m2contact 8937 2122 8937 2122 4 n_158
rlabel m2contact 8913 6610 8913 6610 4 n_87
rlabel m2contact 8913 4426 8913 4426 4 OpcodeCondIn[5]
rlabel m2contact 8889 2122 8889 2122 4 n_158
rlabel m2contact 8889 4114 8889 4114 4 n_84
rlabel m2contact 8865 5914 8865 5914 4 n_89
rlabel m2contact 8841 6586 8841 6586 4 n_36
rlabel m2contact 8817 6562 8817 6562 4 n_20
rlabel m2contact 8817 3346 8817 3346 4 OpcodeCondIn[6]
rlabel m2contact 8793 5818 8793 5818 4 n_13
rlabel m2contact 8769 4498 8769 4498 4 n_210
rlabel m2contact 8745 2146 8745 2146 4 n_360
rlabel m2contact 8745 3922 8745 3922 4 n_99
rlabel m2contact 8697 2194 8697 2194 4 n_358
rlabel m2contact 8673 5986 8673 5986 4 n_174
rlabel m2contact 8649 4186 8649 4186 4 n_359
rlabel m2contact 8625 6298 8625 6298 4 n_158
rlabel m2contact 8601 2170 8601 2170 4 n_361
rlabel m2contact 8601 5818 8601 5818 4 n_297
rlabel m2contact 8601 2194 8601 2194 4 n_297
rlabel m2contact 8577 2194 8577 2194 4 n_297
rlabel m2contact 8577 4186 8577 4186 4 n_223
rlabel m2contact 8553 6538 8553 6538 4 n_222
rlabel m2contact 8553 6514 8553 6514 4 n_334
rlabel m2contact 8529 2218 8529 2218 4 n_178
rlabel m2contact 8481 6490 8481 6490 4 MemEn
rlabel m2contact 8481 6466 8481 6466 4 PcEn
rlabel m2contact 8457 4378 8457 4378 4 n_87
rlabel m2contact 8409 2458 8409 2458 4 n_202
rlabel m2contact 8409 4378 8409 4378 4 n_215
rlabel m2contact 8385 2986 8385 2986 4 n_329
rlabel m2contact 8337 6442 8337 6442 4 n_64
rlabel m2contact 8337 5242 8337 5242 4 n_341
rlabel m2contact 8313 6418 8313 6418 4 n_40
rlabel m2contact 8289 5674 8289 5674 4 n_47
rlabel m2contact 8289 4306 8289 4306 4 n_194
rlabel m2contact 8265 4642 8265 4642 4 n_46
rlabel m2contact 8265 4330 8265 4330 4 n_254
rlabel m2contact 8241 6418 8241 6418 4 n_216
rlabel m2contact 8241 2458 8241 2458 4 n_216
rlabel m2contact 8217 2242 8217 2242 4 n_224
rlabel m2contact 8217 4642 8217 4642 4 n_249
rlabel m2contact 8193 3058 8193 3058 4 n_88
rlabel m2contact 8169 6418 8169 6418 4 n_216
rlabel m2contact 8169 4138 8169 4138 4 n_169
rlabel m2contact 8145 3058 8145 3058 4 n_142
rlabel m2contact 8121 2266 8121 2266 4 n_116
rlabel m2contact 8097 4762 8097 4762 4 OpcodeCondIn[7]
rlabel m2contact 8073 6034 8073 6034 4 n_77
rlabel m2contact 8073 5746 8073 5746 4 stateSub[1]
rlabel m2contact 8049 6250 8049 6250 4 n_138
rlabel m2contact 8025 6034 8025 6034 4 n_164
rlabel m2contact 8001 4762 8001 4762 4 OpcodeCondIn[7]
rlabel m2contact 7977 6250 7977 6250 4 n_133
rlabel m2contact 7977 4762 7977 4762 4 OpcodeCondIn[7]
rlabel m2contact 7953 4066 7953 4066 4 n_252
rlabel m2contact 7929 6394 7929 6394 4 n_333
rlabel m2contact 7929 3322 7929 3322 4 OpcodeCondIn[3]
rlabel m2contact 7905 6370 7905 6370 4 n_90
rlabel m2contact 7881 6346 7881 6346 4 n_311
rlabel m2contact 7881 2290 7881 2290 4 RwSel[1]
rlabel m2contact 7857 2314 7857 2314 4 n_346
rlabel m2contact 7833 6322 7833 6322 4 n_192
rlabel m2contact 7833 5218 7833 5218 4 n_347
rlabel m2contact 7809 2362 7809 2362 4 n_265
rlabel m2contact 7809 3778 7809 3778 4 n_69
rlabel m2contact 7785 4738 7785 4738 4 n_201
rlabel m2contact 7761 2338 7761 2338 4 n_343
rlabel m2contact 7761 5386 7761 5386 4 n_310
rlabel m2contact 7761 2362 7761 2362 4 n_310
rlabel m2contact 7737 3946 7737 3946 4 n_226
rlabel m2contact 7713 2362 7713 2362 4 n_310
rlabel m2contact 7713 4834 7713 4834 4 n_172
rlabel m2contact 7689 5986 7689 5986 4 n_174
rlabel m2contact 7641 2386 7641 2386 4 n_134
rlabel m2contact 7617 4282 7617 4282 4 n_155
rlabel m2contact 7593 4834 7593 4834 4 n_172
rlabel m2contact 7569 2842 7569 2842 4 n_256
rlabel m2contact 7569 4882 7569 4882 4 n_126
rlabel m2contact 7521 2458 7521 2458 4 n_216
rlabel m2contact 7521 4738 7521 4738 4 n_201
rlabel m2contact 7473 5410 7473 5410 4 OpcodeCondIn[4]
rlabel m2contact 7449 6298 7449 6298 4 n_158
rlabel m2contact 7449 4114 7449 4114 4 n_84
rlabel m2contact 7425 2938 7425 2938 4 state[0]
rlabel m2contact 7401 6274 7401 6274 4 n_115
rlabel m2contact 7401 5986 7401 5986 4 n_174
rlabel m2contact 7401 2458 7401 2458 4 n_174
rlabel m2contact 7377 2410 7377 2410 4 n_175
rlabel m2contact 7377 3682 7377 3682 4 nWait
rlabel m2contact 7353 2434 7353 2434 4 n_82
rlabel m2contact 7353 5290 7353 5290 4 n_231
rlabel m2contact 7329 2458 7329 2458 4 n_174
rlabel m2contact 7329 5914 7329 5914 4 n_89
rlabel m2contact 7281 6250 7281 6250 4 n_133
rlabel m2contact 7257 4546 7257 4546 4 n_325
rlabel m2contact 7257 3322 7257 3322 4 OpcodeCondIn[3]
rlabel m2contact 7233 6226 7233 6226 4 n_263
rlabel m2contact 7233 6202 7233 6202 4 n_103
rlabel m2contact 7209 4042 7209 4042 4 n_218
rlabel m2contact 7185 6178 7185 6178 4 n_124
rlabel m2contact 7137 6154 7137 6154 4 n_94
rlabel m2contact 7137 4210 7137 4210 4 n_208
rlabel m2contact 7113 4810 7113 4810 4 n_58
rlabel m2contact 7089 5842 7089 5842 4 n_56
rlabel m2contact 7041 5746 7041 5746 4 stateSub[1]
rlabel m2contact 7041 5842 7041 5842 4 n_362
rlabel m2contact 7017 5962 7017 5962 4 n_274
rlabel m2contact 7017 4930 7017 4930 4 n_123
rlabel m2contact 6993 2482 6993 2482 4 n_335
rlabel m2contact 6969 2506 6969 2506 4 n_30
rlabel m2contact 6969 5962 6969 5962 4 n_288
rlabel m2contact 6945 3226 6945 3226 4 n_59
rlabel m2contact 6921 2986 6921 2986 4 n_329
rlabel m2contact 6897 6058 6897 6058 4 n_135
rlabel m2contact 6873 6130 6873 6130 4 n_302
rlabel m2contact 6873 5362 6873 5362 4 n_260
rlabel m2contact 6849 6058 6849 6058 4 OpcodeCondIn[1]
rlabel m2contact 6849 3514 6849 3514 4 OpcodeCondIn[1]
rlabel m2contact 6825 6106 6825 6106 4 n_5
rlabel m2contact 6825 4762 6825 4762 4 OpcodeCondIn[7]
rlabel m2contact 6801 6058 6801 6058 4 OpcodeCondIn[1]
rlabel m2contact 6801 3946 6801 3946 4 n_226
rlabel m2contact 6777 3538 6777 3538 4 OpcodeCondIn[0]
rlabel m2contact 6753 2986 6753 2986 4 n_66
rlabel m2contact 6729 6082 6729 6082 4 n_182
rlabel m2contact 6729 6058 6729 6058 4 n_139
rlabel m2contact 6729 2698 6729 2698 4 n_139
rlabel m2contact 6705 6058 6705 6058 4 n_139
rlabel m2contact 6705 3082 6705 3082 4 n_217
rlabel m2contact 6681 6034 6681 6034 4 n_164
rlabel m2contact 6681 3250 6681 3250 4 n_65
rlabel m2contact 6633 2554 6633 2554 4 n_100
rlabel m2contact 6633 4138 6633 4138 4 n_169
rlabel m2contact 6585 5746 6585 5746 4 stateSub[1]
rlabel m2contact 6585 4426 6585 4426 4 OpcodeCondIn[5]
rlabel m2contact 6561 2530 6561 2530 4 n_67
rlabel m2contact 6561 3850 6561 3850 4 state[1]
rlabel m2contact 6537 5746 6537 5746 4 SysBus[3]
rlabel m2contact 6537 2554 6537 2554 4 SysBus[3]
rlabel m2contact 6513 2554 6513 2554 4 SysBus[3]
rlabel m2contact 6513 3442 6513 3442 4 n_157
rlabel m2contact 6489 2818 6489 2818 4 n_199
rlabel m2contact 6465 6010 6465 6010 4 n_147
rlabel m2contact 6417 5578 6417 5578 4 n_171
rlabel m2contact 6393 4402 6393 4402 4 n_104
rlabel m2contact 6369 5986 6369 5986 4 n_174
rlabel m2contact 6369 5578 6369 5578 4 StatusReg[2]
rlabel m2contact 6321 5962 6321 5962 4 n_288
rlabel m2contact 6297 5578 6297 5578 4 StatusReg[2]
rlabel m2contact 6273 2650 6273 2650 4 n_289
rlabel m2contact 6225 5650 6225 5650 4 n_365
rlabel m2contact 6201 2578 6201 2578 4 n_275
rlabel m2contact 6177 5650 6177 5650 4 n_337
rlabel m2contact 6153 5938 6153 5938 4 n_290
rlabel m2contact 6105 2602 6105 2602 4 n_71
rlabel m2contact 6081 5530 6081 5530 4 n_26
rlabel m2contact 6057 5914 6057 5914 4 n_89
rlabel m2contact 6009 5890 6009 5890 4 n_295
rlabel m2contact 5985 3610 5985 3610 4 n_107
rlabel m2contact 5961 5866 5961 5866 4 n_230
rlabel m2contact 5961 5842 5961 5842 4 n_362
rlabel m2contact 5913 3802 5913 3802 4 n_118
rlabel m2contact 5865 3802 5865 3802 4 n_70
rlabel m2contact 5841 2626 5841 2626 4 n_83
rlabel m2contact 5817 4426 5817 4426 4 OpcodeCondIn[5]
rlabel m2contact 5793 5818 5793 5818 4 n_297
rlabel m2contact 5793 5794 5793 5794 4 n_113
rlabel m2contact 5769 5746 5769 5746 4 SysBus[3]
rlabel m2contact 5745 2650 5745 2650 4 n_289
rlabel m2contact 5745 4522 5745 4522 4 n_276
rlabel m2contact 5697 5770 5697 5770 4 n_11
rlabel m2contact 5697 5746 5697 5746 4 OpcodeCondIn[3]
rlabel m2contact 5697 3322 5697 3322 4 OpcodeCondIn[3]
rlabel m2contact 5673 5746 5673 5746 4 OpcodeCondIn[3]
rlabel m2contact 5673 4306 5673 4306 4 n_194
rlabel m2contact 5649 5722 5649 5722 4 n_10
rlabel m2contact 5649 5698 5649 5698 4 n_121
rlabel m2contact 5601 5674 5601 5674 4 n_47
rlabel m2contact 5601 5650 5601 5650 4 n_337
rlabel m2contact 5577 5626 5577 5626 4 n_479
rlabel m2contact 5577 5602 5577 5602 4 Flags[1]
rlabel m2contact 5553 5578 5553 5578 4 StatusReg[2]
rlabel m2contact 5553 2674 5553 2674 4 n_336
rlabel m2contact 5481 3322 5481 3322 4 OpcodeCondIn[3]
rlabel m2contact 5481 3610 5481 3610 4 n_107
rlabel m2contact 5457 5554 5457 5554 4 n_86
rlabel m2contact 5433 5530 5433 5530 4 n_26
rlabel m2contact 5409 2698 5409 2698 4 n_139
rlabel m2contact 5385 5506 5385 5506 4 n_39
rlabel m2contact 5361 2722 5361 2722 4 n_161
rlabel m2contact 5337 3538 5337 3538 4 OpcodeCondIn[0]
rlabel m2contact 5313 5482 5313 5482 4 n_12
rlabel m2contact 5313 2746 5313 2746 4 n_132
rlabel m2contact 5265 5458 5265 5458 4 n_255
rlabel m2contact 5265 5434 5265 5434 4 n_253
rlabel m2contact 5241 5410 5241 5410 4 OpcodeCondIn[4]
rlabel m2contact 5241 3346 5241 3346 4 OpcodeCondIn[6]
rlabel m2contact 5217 4066 5217 4066 4 n_252
rlabel m2contact 5193 2770 5193 2770 4 n_68
rlabel m2contact 5193 4330 5193 4330 4 n_254
rlabel m2contact 5145 5386 5145 5386 4 n_310
rlabel m2contact 5145 3034 5145 3034 4 n_6
rlabel m2contact 5121 3346 5121 3346 4 OpcodeCondIn[6]
rlabel m2contact 5097 3730 5097 3730 4 stateSub[0]
rlabel m2contact 5073 3874 5073 3874 4 n_354
rlabel m2contact 5025 4258 5025 4258 4 n_261
rlabel m2contact 5025 3034 5025 3034 4 n_23
rlabel m2contact 5001 2794 5001 2794 4 n_63
rlabel m2contact 5001 4330 5001 4330 4 n_254
rlabel m2contact 4977 5362 4977 5362 4 n_260
rlabel m2contact 4977 4258 4977 4258 4 n_60
rlabel m2contact 4905 5338 4905 5338 4 n_323
rlabel m2contact 4881 2818 4881 2818 4 n_199
rlabel m2contact 4857 5314 4857 5314 4 n_314
rlabel m2contact 4857 4738 4857 4738 4 n_201
rlabel m2contact 4833 2842 4833 2842 4 n_256
rlabel m2contact 4809 5290 4809 5290 4 n_231
rlabel m2contact 4785 5266 4785 5266 4 n_8
rlabel m2contact 4761 3514 4761 3514 4 OpcodeCondIn[1]
rlabel m2contact 4761 3730 4761 3730 4 stateSub[0]
rlabel m2contact 4737 2866 4737 2866 4 StatusReg[0]
rlabel m2contact 4737 3610 4737 3610 4 n_107
rlabel m2contact 4713 3538 4713 3538 4 OpcodeCondIn[0]
rlabel m2contact 4689 2890 4689 2890 4 Rs1Sel[1]
rlabel m2contact 4665 5242 4665 5242 4 n_341
rlabel m2contact 4665 5146 4665 5146 4 n_203
rlabel m2contact 4641 2914 4641 2914 4 n_351
rlabel m2contact 4617 5218 4617 5218 4 n_347
rlabel m2contact 4617 2938 4617 2938 4 state[0]
rlabel m2contact 4593 5194 4593 5194 4 n_355
rlabel m2contact 4593 3610 4593 3610 4 n_107
rlabel m2contact 4545 5170 4545 5170 4 n_345
rlabel m2contact 4545 4786 4545 4786 4 n_324
rlabel m2contact 4521 3250 4521 3250 4 n_65
rlabel m2contact 4497 2962 4497 2962 4 n_315
rlabel m2contact 4473 4786 4473 4786 4 n_296
rlabel m2contact 4425 4306 4425 4306 4 n_194
rlabel m2contact 4377 3922 4377 3922 4 n_99
rlabel m2contact 4353 5146 4353 5146 4 n_203
rlabel m2contact 4329 5122 4329 5122 4 n_17
rlabel m2contact 4305 5098 4305 5098 4 n_299
rlabel m2contact 4305 3514 4305 3514 4 OpcodeCondIn[1]
rlabel m2contact 4281 2986 4281 2986 4 n_66
rlabel m2contact 4257 5074 4257 5074 4 n_234
rlabel m2contact 4257 3346 4257 3346 4 OpcodeCondIn[6]
rlabel m2contact 4233 5050 4233 5050 4 n_129
rlabel m2contact 4233 4762 4233 4762 4 OpcodeCondIn[7]
rlabel m2contact 4209 3010 4209 3010 4 n_109
rlabel m2contact 4161 4786 4161 4786 4 n_296
rlabel m2contact 4137 5026 4137 5026 4 n_170
rlabel m2contact 4113 4786 4113 4786 4 n_198
rlabel m2contact 4089 5002 4089 5002 4 n_191
rlabel m2contact 4089 4978 4089 4978 4 n_141
rlabel m2contact 4065 4954 4065 4954 4 n_211
rlabel m2contact 4017 3034 4017 3034 4 n_23
rlabel m2contact 3993 4930 3993 4930 4 n_123
rlabel m2contact 3969 4138 3969 4138 4 n_169
rlabel m2contact 3945 3850 3945 3850 4 state[1]
rlabel m2contact 3921 3058 3921 3058 4 n_142
rlabel m2contact 3897 4906 3897 4906 4 n_80
rlabel m2contact 3897 3082 3897 3082 4 n_217
rlabel m2contact 3873 4882 3873 4882 4 n_126
rlabel m2contact 3825 4858 3825 4858 4 n_74
rlabel m2contact 3801 4834 3801 4834 4 n_172
rlabel m2contact 3777 4810 3777 4810 4 n_58
rlabel m2contact 3729 4786 3729 4786 4 n_198
rlabel m2contact 3705 4762 3705 4762 4 OpcodeCondIn[7]
rlabel m2contact 3681 4738 3681 4738 4 n_201
rlabel m2contact 3657 4714 3657 4714 4 n_241
rlabel m2contact 3633 3322 3633 3322 4 OpcodeCondIn[3]
rlabel m2contact 3585 4690 3585 4690 4 n_285
rlabel m2contact 3561 3106 3561 3106 4 n_228
rlabel m2contact 3537 4666 3537 4666 4 n_278
rlabel m2contact 3537 4642 3537 4642 4 n_249
rlabel m2contact 3465 4546 3465 4546 4 n_325
rlabel m2contact 3441 3130 3441 3130 4 n_303
rlabel m2contact 3417 3154 3417 3154 4 n_237
rlabel m2contact 3393 4618 3393 4618 4 n_286
rlabel m2contact 3393 3178 3393 3178 4 n_176
rlabel m2contact 3369 4594 3369 4594 4 n_236
rlabel m2contact 3369 3370 3369 3370 4 n_214
rlabel m2contact 3345 4570 3345 4570 4 n_206
rlabel m2contact 3345 3730 3345 3730 4 stateSub[0]
rlabel m2contact 3273 4498 3273 4498 4 n_210
rlabel m2contact 3225 4546 3225 4546 4 n_325
rlabel m2contact 3225 3298 3225 3298 4 OpcodeCondIn[2]
rlabel m2contact 3177 4522 3177 4522 4 n_276
rlabel m2contact 3177 3202 3177 3202 4 n_97
rlabel m2contact 3129 4498 3129 4498 4 n_210
rlabel m2contact 3129 3226 3129 3226 4 n_59
rlabel m2contact 3105 4474 3105 4474 4 n_229
rlabel m2contact 3105 3250 3105 3250 4 n_65
rlabel m2contact 3057 4450 3057 4450 4 n_105
rlabel m2contact 3057 3274 3057 3274 4 n_16
rlabel m2contact 3033 3298 3033 3298 4 OpcodeCondIn[2]
rlabel m2contact 3009 4426 3009 4426 4 OpcodeCondIn[5]
rlabel m2contact 3009 3322 3009 3322 4 OpcodeCondIn[3]
rlabel m2contact 2985 4402 2985 4402 4 n_104
rlabel m2contact 2961 4378 2961 4378 4 n_215
rlabel m2contact 2937 4354 2937 4354 4 n_156
rlabel m2contact 2937 3346 2937 3346 4 OpcodeCondIn[6]
rlabel m2contact 2913 4330 2913 4330 4 n_254
rlabel m2contact 2913 3370 2913 3370 4 n_214
rlabel m2contact 2889 4306 2889 4306 4 n_194
rlabel m2contact 2889 3394 2889 3394 4 n_269
rlabel m2contact 2865 4282 2865 4282 4 n_155
rlabel m2contact 2841 3418 2841 3418 4 n_220
rlabel m2contact 2817 3442 2817 3442 4 n_157
rlabel m2contact 2793 4258 2793 4258 4 n_60
rlabel m2contact 2793 3466 2793 3466 4 n_195
rlabel m2contact 2745 3826 2745 3826 4 n_76
rlabel m2contact 2721 4234 2721 4234 4 n_15
rlabel m2contact 2697 3490 2697 3490 4 n_266
rlabel m2contact 2673 4210 2673 4210 4 n_208
rlabel m2contact 2649 4186 2649 4186 4 n_223
rlabel m2contact 2625 3514 2625 3514 4 OpcodeCondIn[1]
rlabel m2contact 2601 4162 2601 4162 4 n_50
rlabel m2contact 2601 3538 2601 3538 4 OpcodeCondIn[0]
rlabel m2contact 2553 3562 2553 3562 4 n_21
rlabel m2contact 2529 4138 2529 4138 4 n_169
rlabel m2contact 2529 3586 2529 3586 4 n_177
rlabel m2contact 2505 3610 2505 3610 4 n_107
rlabel m2contact 2457 4114 2457 4114 4 n_84
rlabel m2contact 2409 4090 2409 4090 4 n_27
rlabel m2contact 2385 3682 2385 3682 4 nWait
rlabel m2contact 2337 4066 2337 4066 4 n_252
rlabel m2contact 2289 4042 2289 4042 4 n_218
rlabel m2contact 2241 3730 2241 3730 4 stateSub[0]
rlabel m2contact 2217 3730 2217 3730 4 stateSub[0]
rlabel m2contact 2193 4018 2193 4018 4 n_235
rlabel m2contact 2193 3922 2193 3922 4 n_99
rlabel m2contact 2169 3994 2169 3994 4 n_33
rlabel m2contact 2097 3970 2097 3970 4 n_250
rlabel m2contact 2049 3946 2049 3946 4 n_226
rlabel m2contact 2001 3634 2001 3634 4 n_31
rlabel m2contact 1977 3922 1977 3922 4 n_99
rlabel m2contact 1953 3898 1953 3898 4 n_319
rlabel m2contact 1905 3874 1905 3874 4 n_354
rlabel m2contact 1881 3850 1881 3850 4 state[1]
rlabel m2contact 1857 3826 1857 3826 4 n_76
rlabel m2contact 1809 3802 1809 3802 4 n_70
rlabel m2contact 1761 3778 1761 3778 4 n_69
rlabel m2contact 1737 3730 1737 3730 4 stateSub[0]
rlabel m2contact 1713 3754 1713 3754 4 nIRQ
rlabel m2contact 1641 3730 1641 3730 4 stateSub[0]
rlabel m2contact 1617 3706 1617 3706 4 n_271
rlabel metal2 25083 8060 25095 8060 6 StatusRegEn
rlabel metal2 24279 8060 24291 8060 6 StatusReg[3]
rlabel metal2 23475 8060 23487 8060 6 StatusReg[2]
rlabel metal2 22671 8060 22683 8060 6 StatusReg[1]
rlabel metal2 21867 8060 21879 8060 6 StatusReg[0]
rlabel metal2 21735 8060 21747 8060 6 AluEn
rlabel metal2 21039 8060 21051 8060 6 AluWe
rlabel metal2 19455 8060 19467 8060 6 Op2Sel[1]
rlabel metal2 18651 8060 18663 8060 6 Op2Sel[0]
rlabel metal2 18627 8060 18639 8060 6 Op1Sel
rlabel metal2 17703 8060 17715 8060 6 PcEn
rlabel metal2 16239 8060 16251 8060 6 WdSel
rlabel metal2 15435 8060 15447 8060 6 PcWe
rlabel metal2 14631 8060 14643 8060 6 PcSel[2]
rlabel metal2 14607 8060 14619 8060 6 PcSel[1]
rlabel metal2 13023 8060 13035 8060 4 PcSel[0]
rlabel metal2 12207 8060 12219 8060 4 LrEn
rlabel metal2 12171 8060 12183 8060 4 LrWe
rlabel metal2 11355 8060 11367 8060 4 LrSel
rlabel metal2 10263 8060 10275 8060 4 ImmSel
rlabel metal2 9375 8060 9387 8060 4 IrWe
rlabel metal2 8487 8060 8499 8060 4 MemEn
rlabel metal2 8007 8060 8019 8060 4 OpcodeCondIn[7]
rlabel metal2 7275 8060 7287 8060 4 OpcodeCondIn[6]
rlabel metal2 5679 8060 5691 8060 4 OpcodeCondIn[5]
rlabel metal2 5247 8060 5259 8060 4 OpcodeCondIn[4]
rlabel metal2 4047 8060 4059 8060 4 OpcodeCondIn[3]
rlabel metal2 4011 8060 4023 8060 4 OpcodeCondIn[2]
rlabel metal2 3195 8060 3207 8060 4 OpcodeCondIn[1]
rlabel metal2 2379 8060 2391 8060 4 OpcodeCondIn[0]
rlabel metal2 19899 0 19911 0 8 SysBus[3]
rlabel metal2 19767 0 19779 0 8 SysBus[2]
rlabel metal2 13779 0 13791 0 8 SysBus[1]
rlabel metal2 7671 0 7683 0 2 SysBus[0]
rlabel metal2 26521 491 26521 503 8 RegWe
rlabel metal2 26521 59 26521 71 8 AluOR[0]
rlabel metal2 26521 35 26521 47 8 AluOR[1]
rlabel metal2 26521 11 26521 23 8 ENB
rlabel metal2 26521 4300 26521 4312 6 Rs1Sel[0]
rlabel metal2 26521 2884 26521 2896 6 Rs1Sel[1]
rlabel metal2 26521 2620 26521 2632 6 RwSel[0]
rlabel metal2 26521 2284 26521 2296 6 RwSel[1]
rlabel metal2 26521 7845 26521 7857 6 CFlag
rlabel metal2 26521 7821 26521 7833 6 Flags[3]
rlabel metal2 26521 7797 26521 7809 6 Flags[2]
rlabel metal2 26521 7773 26521 7785 6 Flags[1]
rlabel metal2 26521 7749 26521 7761 6 Flags[0]
rlabel metal2 26139 8060 26339 8060 5 GND!
rlabel metal2 26139 0 26339 0 1 GND!
rlabel metal2 0 59 0 71 2 nWE
rlabel metal2 0 35 0 47 2 nIRQ
rlabel metal2 0 3676 0 3688 4 nWait
rlabel metal2 0 3652 0 3664 4 nOE
rlabel metal2 0 7893 0 7905 4 ALE
rlabel metal2 0 7869 0 7881 4 nME
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 123 8060 323 8060 5 Vdd!
rlabel metal2 339 8060 351 8060 5 SDO
rlabel metal2 363 8060 375 8060 5 Test
rlabel metal2 387 8060 399 8060 5 Clock
rlabel metal2 411 8060 423 8060 5 nReset
<< end >>
