magic
tech c035u
timestamp 1395339964
<< nwell >>
rect 1464 684 3720 1082
rect 15289 684 15912 1082
rect 23568 684 24336 1082
<< pwell >>
rect 1464 283 3720 684
rect 15289 290 15912 684
rect 23568 283 24336 684
<< pohmic >>
rect 1464 359 1470 369
rect 3714 359 3720 369
rect 15289 359 15294 369
rect 15906 359 15912 369
rect 23568 359 23572 369
rect 24330 359 24336 369
<< nohmic >>
rect 1464 1019 1470 1029
rect 3716 1019 3720 1029
rect 15289 1019 15294 1029
rect 15906 1019 15912 1029
rect 23568 1019 23572 1029
rect 24330 1019 24336 1029
<< psubstratetap >>
rect 1470 359 3714 375
rect 15294 359 15906 375
rect 23572 359 24330 375
<< nsubstratetap >>
rect 1470 1013 3716 1029
rect 15294 1013 15906 1029
rect 23572 1013 24330 1029
<< metal1 >>
rect 4621 1286 5807 1296
rect 4669 1264 5759 1274
rect 6014 1268 6072 1278
rect 4285 1242 5375 1252
rect 5990 1246 6072 1256
rect 4237 1220 5423 1230
rect 5461 1220 5567 1230
rect 5653 1220 5976 1230
rect 6037 1223 6072 1233
rect 3805 1198 5039 1208
rect 5077 1198 5183 1208
rect 5269 1198 6000 1208
rect 15289 1197 15912 1207
rect 3853 1176 4991 1186
rect 5173 1176 5543 1186
rect 5557 1176 5927 1186
rect 15289 1175 15912 1185
rect 4021 1154 4391 1164
rect 4405 1154 4775 1164
rect 4981 1154 5351 1164
rect 5365 1154 5735 1164
rect 5845 1154 5951 1164
rect 15289 1153 15912 1163
rect 4117 1132 6072 1142
rect 15289 1131 15912 1141
rect 3877 1110 4031 1120
rect 4309 1110 4415 1120
rect 4501 1110 6072 1120
rect 15289 1109 15912 1119
rect 3781 1088 4199 1098
rect 4213 1088 4583 1098
rect 4693 1087 4799 1097
rect 4885 1087 6072 1097
rect 15289 1087 15912 1097
rect 1464 1065 3720 1075
rect 15289 1065 15912 1075
rect 23568 1065 24336 1075
rect 1464 1042 3720 1052
rect 15289 1042 15912 1052
rect 23568 1042 24336 1052
rect 1464 1013 1470 1029
rect 3716 1013 3720 1029
rect 1464 1004 3720 1013
rect 15289 1013 15294 1029
rect 15906 1013 15912 1029
rect 15289 1004 15912 1013
rect 23568 1013 23572 1029
rect 24330 1013 24336 1029
rect 23568 1004 24336 1013
rect 1464 375 3720 384
rect 1464 359 1470 375
rect 3714 359 3720 375
rect 15289 375 15912 384
rect 15289 359 15294 375
rect 15906 359 15912 375
rect 23568 375 24336 384
rect 23568 359 23572 375
rect 24330 359 24336 375
rect 1464 336 3720 346
rect 15289 336 15912 346
rect 1464 313 3720 323
rect 15289 313 15912 323
rect 1464 290 3720 300
rect 15289 290 15912 300
rect 21349 7 21383 17
rect 21397 7 21431 17
rect 21445 7 21479 17
rect 21493 7 21527 17
rect 21541 7 21575 17
rect 21589 7 21623 17
rect 21637 7 21671 17
rect 21685 7 21983 17
rect 21997 7 22031 17
rect 22045 7 22079 17
rect 22093 7 22127 17
rect 22141 7 22439 17
rect 22453 7 22487 17
rect 22501 7 22799 17
<< m2contact >>
rect 4607 1284 4621 1298
rect 5807 1284 5821 1298
rect 4655 1262 4669 1276
rect 5759 1262 5773 1276
rect 6000 1266 6014 1280
rect 4271 1240 4285 1254
rect 5375 1240 5389 1254
rect 5976 1245 5990 1259
rect 4223 1218 4237 1232
rect 5423 1218 5437 1232
rect 5447 1218 5461 1232
rect 5567 1218 5581 1232
rect 5639 1218 5653 1232
rect 5976 1218 5990 1232
rect 6023 1221 6037 1235
rect 3791 1197 3805 1211
rect 5039 1196 5053 1210
rect 5063 1196 5077 1210
rect 5183 1196 5197 1210
rect 5255 1196 5269 1210
rect 6000 1196 6014 1210
rect 3839 1174 3853 1188
rect 4991 1174 5005 1188
rect 5159 1174 5173 1188
rect 5543 1174 5557 1188
rect 5927 1174 5941 1188
rect 4007 1152 4021 1166
rect 4391 1152 4405 1166
rect 4775 1152 4789 1166
rect 4967 1152 4981 1166
rect 5351 1152 5365 1166
rect 5735 1152 5749 1166
rect 5831 1152 5845 1166
rect 5951 1152 5965 1166
rect 4103 1130 4117 1144
rect 3863 1108 3877 1122
rect 4031 1108 4045 1122
rect 4295 1108 4309 1122
rect 4415 1108 4429 1122
rect 4487 1108 4501 1122
rect 3767 1086 3781 1100
rect 4199 1086 4213 1100
rect 4583 1086 4597 1100
rect 4679 1085 4693 1099
rect 4799 1085 4813 1099
rect 4871 1085 4885 1099
rect 21335 5 21349 19
rect 21383 5 21397 19
rect 21431 5 21445 19
rect 21479 5 21493 19
rect 21527 5 21541 19
rect 21575 5 21589 19
rect 21623 5 21637 19
rect 21671 5 21685 19
rect 21983 4 21997 18
rect 22031 4 22045 18
rect 22079 4 22093 18
rect 22127 4 22141 18
rect 22439 5 22453 19
rect 22487 5 22501 19
rect 22799 5 22813 19
<< metal2 >>
rect 0 1082 200 1321
rect 216 1082 228 1321
rect 240 1082 252 1321
rect 264 1082 276 1321
rect 288 1082 300 1321
rect 3768 1100 3780 1321
rect 3792 1211 3804 1321
rect 3768 1082 3780 1086
rect 3792 1082 3804 1197
rect 3840 1188 3852 1321
rect 3840 1082 3852 1174
rect 4008 1166 4020 1321
rect 4224 1232 4236 1321
rect 4272 1254 4284 1321
rect 4608 1298 4620 1321
rect 3864 1082 3876 1108
rect 4008 1082 4020 1152
rect 4032 1082 4044 1108
rect 4104 1082 4116 1130
rect 4200 1082 4212 1086
rect 4224 1082 4236 1218
rect 4272 1082 4284 1240
rect 4296 1082 4308 1108
rect 4392 1082 4404 1152
rect 4416 1082 4428 1108
rect 4488 1082 4500 1108
rect 4584 1082 4596 1086
rect 4608 1082 4620 1284
rect 4656 1276 4668 1321
rect 4656 1082 4668 1262
rect 4968 1166 4980 1321
rect 4680 1082 4692 1085
rect 4776 1082 4788 1152
rect 4800 1082 4812 1085
rect 4872 1082 4884 1085
rect 4968 1082 4980 1152
rect 4992 1082 5004 1174
rect 5040 1082 5052 1196
rect 5064 1082 5076 1196
rect 5160 1188 5172 1321
rect 6194 1309 6206 1321
rect 6748 1309 6760 1321
rect 6772 1309 6784 1321
rect 6796 1309 6808 1321
rect 14185 1309 14197 1321
rect 14209 1309 14221 1321
rect 14401 1309 14413 1321
rect 14449 1309 14461 1321
rect 14593 1309 14605 1321
rect 14785 1309 14797 1321
rect 14977 1309 14989 1321
rect 15169 1309 15181 1321
rect 5160 1082 5172 1174
rect 5184 1082 5196 1196
rect 5256 1082 5268 1196
rect 5352 1082 5364 1152
rect 5376 1082 5388 1240
rect 5424 1082 5436 1218
rect 5448 1082 5460 1218
rect 5544 1082 5556 1174
rect 5568 1082 5580 1218
rect 5640 1082 5652 1218
rect 5736 1082 5748 1152
rect 5760 1082 5772 1262
rect 5808 1082 5820 1284
rect 5977 1232 5989 1245
rect 6001 1210 6013 1266
rect 16968 1258 16980 1321
rect 17160 1258 17172 1321
rect 17232 1258 17244 1321
rect 17328 1258 17340 1321
rect 21984 1258 21996 1321
rect 22176 1258 22188 1321
rect 22296 1258 22308 1321
rect 22416 1258 22428 1321
rect 23496 1258 23508 1321
rect 5832 1082 5844 1152
rect 5928 1082 5940 1174
rect 5952 1082 5964 1152
rect 6024 1082 6036 1221
rect 24456 1082 24656 1321
rect 0 0 200 283
rect 216 0 228 283
rect 240 0 252 283
rect 264 0 276 283
rect 288 0 300 283
rect 3936 273 3948 283
rect 4080 273 4092 283
rect 4320 273 4332 274
rect 4464 273 4476 283
rect 4848 273 4860 283
rect 5232 273 5244 283
rect 5472 273 5484 274
rect 5616 273 5628 283
rect 6000 273 6012 283
rect 3936 261 6012 273
rect 6144 0 6156 178
rect 6888 0 6900 178
rect 7104 0 7116 178
rect 7296 0 7308 178
rect 8040 0 8052 178
rect 8256 0 8268 178
rect 8448 0 8460 178
rect 9192 0 9204 178
rect 9408 0 9420 178
rect 9600 0 9612 178
rect 10344 0 10356 178
rect 10560 0 10572 178
rect 10752 0 10764 178
rect 11496 0 11508 178
rect 11712 0 11724 178
rect 11904 0 11916 178
rect 12648 0 12660 178
rect 12864 0 12876 178
rect 13056 0 13068 178
rect 13800 0 13812 178
rect 14016 0 14028 178
rect 14208 0 14220 178
rect 14952 0 14964 178
rect 15168 0 15180 178
rect 15984 0 15996 19
rect 16248 0 16260 19
rect 16416 0 16428 19
rect 16584 0 16596 19
rect 16608 0 16620 19
rect 16680 0 16692 19
rect 16896 0 16908 19
rect 17040 0 17052 19
rect 17376 0 17388 19
rect 17736 0 17748 19
rect 18144 0 18156 19
rect 18480 0 18492 19
rect 18792 0 18804 19
rect 19128 0 19140 19
rect 19248 0 19260 19
rect 19296 0 19308 19
rect 19464 0 19476 19
rect 21264 0 21276 19
rect 21289 0 21301 19
rect 21336 0 21348 5
rect 21384 0 21396 5
rect 21432 0 21444 5
rect 21480 0 21492 5
rect 21528 0 21540 5
rect 21576 0 21588 5
rect 21624 0 21636 5
rect 21672 0 21684 5
rect 21912 0 21924 19
rect 21984 0 21996 4
rect 22032 0 22044 4
rect 22080 0 22092 4
rect 22128 0 22140 4
rect 22368 0 22380 19
rect 22440 0 22452 5
rect 22488 0 22500 5
rect 22728 0 22740 19
rect 22800 0 22812 5
rect 23088 0 23100 19
rect 23256 0 23268 19
rect 23496 7 24228 19
rect 24216 0 24228 7
rect 24456 0 24656 283
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 0 0 1 283
box 0 0 1464 799
use mux2 mux2_6
timestamp 1386235218
transform 1 0 3720 0 1 283
box 0 0 192 799
use tiehigh tiehigh_3
timestamp 1386086759
transform 1 0 3912 0 1 283
box 0 0 48 799
use mux2 mux2_7
timestamp 1386235218
transform 1 0 3960 0 1 283
box 0 0 192 799
use mux2 mux2_8
timestamp 1386235218
transform 1 0 4152 0 1 283
box 0 0 192 799
use mux2 mux2_9
timestamp 1386235218
transform 1 0 4344 0 1 283
box 0 0 192 799
use mux2 mux2_10
timestamp 1386235218
transform 1 0 4536 0 1 283
box 0 0 192 799
use mux2 mux2_11
timestamp 1386235218
transform 1 0 4728 0 1 283
box 0 0 192 799
use mux2 mux2_4
timestamp 1386235218
transform 1 0 4920 0 1 283
box 0 0 192 799
use mux2 mux2_5
timestamp 1386235218
transform 1 0 5112 0 1 283
box 0 0 192 799
use mux2 mux2_2
timestamp 1386235218
transform 1 0 5304 0 1 283
box 0 0 192 799
use mux2 mux2_3
timestamp 1386235218
transform 1 0 5496 0 1 283
box 0 0 192 799
use mux2 mux2_1
timestamp 1386235218
transform 1 0 5688 0 1 283
box 0 0 192 799
use mux2 mux2_0
timestamp 1386235218
transform 1 0 5880 0 1 283
box 0 0 192 799
use regBlock_decoder regBlock_decoder_0
timestamp 1395339189
transform 1 0 6072 0 1 178
box 0 0 9217 1131
use ALUDecoder_new ALUDecoder_new_0
timestamp 1395338636
transform 1 0 15912 0 1 19
box 0 0 7656 1239
use rightend rightend_0
timestamp 1386235834
transform 1 0 24336 0 1 283
box 0 0 320 799
<< labels >>
rlabel metal1 6069 1228 6069 1228 1 Rw0
rlabel metal1 6068 1250 6068 1250 1 Rw1
rlabel metal1 6063 1270 6063 1270 1 Rw2
rlabel metal1 15877 1090 15877 1090 1 AOp0
rlabel metal1 15878 1112 15878 1112 1 AOp1
rlabel metal1 15878 1133 15878 1133 1 AOp2
rlabel metal1 15878 1158 15878 1158 1 AOp3
rlabel metal1 15877 1178 15877 1178 1 AOp4
rlabel metal1 15876 1201 15876 1201 1 ACin
rlabel metal2 4272 1321 4284 1321 5 Ir[6]
rlabel metal2 4224 1321 4236 1321 5 Ir[9]
rlabel metal2 3840 1321 3852 1321 5 Ir[7]
rlabel metal2 3792 1321 3804 1321 5 Ir[10]
rlabel metal2 4008 1321 4020 1321 5 Rs1Sel[1]
rlabel metal2 3768 1321 3780 1321 5 Rs1Sel[0]
rlabel metal2 4608 1321 4620 1321 5 Ir[8]
rlabel metal2 4656 1321 4668 1321 5 Ir[5]
rlabel metal2 4968 1321 4980 1321 5 RwSel[0]
rlabel metal2 5160 1321 5172 1321 5 RwSel[1]
rlabel metal2 14185 1321 14197 1321 1 AluOR[1]
rlabel metal2 14209 1321 14221 1321 5 Ir[15]
rlabel metal2 14401 1321 14413 1321 5 Ir[14]
rlabel metal2 14449 1321 14461 1321 1 AluOR[0]
rlabel metal2 14593 1321 14605 1321 5 Ir[13]
rlabel metal2 14785 1321 14797 1321 5 Ir[12]
rlabel metal2 14977 1321 14989 1321 5 Ir[11]
rlabel metal2 15169 1321 15181 1321 5 Cin
rlabel metal2 6796 1321 6808 1321 5 Ir[4]
rlabel metal2 6772 1321 6784 1321 5 Ir[3]
rlabel metal2 6748 1321 6760 1321 5 Ir[2]
rlabel metal2 23496 1321 23508 1321 5 ALUOutEn
rlabel metal2 6194 1321 6206 1321 5 RegWe
rlabel metal2 240 1321 252 1321 1 Test
rlabel metal2 264 1321 276 1321 1 Clock
rlabel metal2 288 1321 300 1321 1 nReset
rlabel metal2 0 1321 200 1321 5 Vdd!
rlabel metal2 216 1321 228 1321 5 SDO
rlabel metal2 24456 1321 24656 1321 1 GND!
rlabel metal2 17232 1321 17244 1321 5 Flags[3]
rlabel metal2 17160 1321 17172 1321 5 Flags[1]
rlabel metal2 16968 1321 16980 1321 5 Flags[2]
rlabel metal2 21984 1321 21996 1321 5 Ir[3]
rlabel metal2 22176 1321 22188 1321 5 Ir[2]
rlabel metal2 22296 1321 22308 1321 5 Ir[1]
rlabel metal2 22416 1321 22428 1321 5 Ir[0]
rlabel metal2 17328 1321 17340 1321 5 Flags[0]
rlabel metal2 22728 0 22740 0 1 Sh1
rlabel metal2 22368 0 22380 0 1 Sh2
rlabel metal2 21912 0 21924 0 1 Sh4
rlabel metal2 24216 0 24228 0 1 ALUOutEn
rlabel metal2 22800 0 22812 0 1 ShiftIn
rlabel metal2 22488 0 22500 0 1 ShiftIn
rlabel metal2 22440 0 22452 0 1 ShiftIn
rlabel metal2 22128 0 22140 0 1 ShiftIn
rlabel metal2 22080 0 22092 0 1 ShiftIn
rlabel metal2 22032 0 22044 0 1 ShiftIn
rlabel metal2 21984 0 21996 0 1 ShiftIn
rlabel metal2 21672 0 21684 0 1 ShiftIn
rlabel metal2 21624 0 21636 0 1 ShiftIn
rlabel metal2 21576 0 21588 0 1 ShiftIn
rlabel metal2 21528 0 21540 0 1 ShiftIn
rlabel metal2 21480 0 21492 0 1 ShiftIn
rlabel metal2 21432 0 21444 0 1 ShiftIn
rlabel metal2 21384 0 21396 0 1 ShiftIn
rlabel metal2 21336 0 21348 0 1 ShiftIn
rlabel metal2 0 0 200 0 1 Vdd!
rlabel metal2 288 0 300 0 1 nReset
rlabel metal2 264 0 276 0 1 Clock
rlabel metal2 240 0 252 0 1 Test
rlabel metal2 216 0 228 0 1 SDI
rlabel metal2 10560 0 10572 0 1 Rs2[3]
rlabel metal2 8040 0 8052 0 1 Rs1[1]
rlabel metal2 7296 0 7308 0 1 Rw[1]
rlabel metal2 15168 0 15180 0 1 Rs2[7]
rlabel metal2 14952 0 14964 0 1 Rs1[7]
rlabel metal2 14208 0 14220 0 1 Rw[7]
rlabel metal2 14016 0 14028 0 1 Rs2[6]
rlabel metal2 13800 0 13812 0 1 Rs1[6]
rlabel metal2 13056 0 13068 0 1 Rw[6]
rlabel metal2 12864 0 12876 0 1 Rs2[5]
rlabel metal2 12648 0 12660 0 1 Rs1[5]
rlabel metal2 11904 0 11916 0 1 Rw[5]
rlabel metal2 11712 0 11724 0 1 Rs2[4]
rlabel metal2 11496 0 11508 0 1 Rs1[4]
rlabel metal2 10752 0 10764 0 1 Rw[4]
rlabel metal2 10344 0 10356 0 1 Rs1[3]
rlabel metal2 9600 0 9612 0 1 Rw[3]
rlabel metal2 9408 0 9420 0 1 Rs2[2]
rlabel metal2 9192 0 9204 0 1 Rs1[2]
rlabel metal2 8448 0 8460 0 1 Rw[2]
rlabel metal2 8256 0 8268 0 1 Rs2[1]
rlabel metal2 7104 0 7116 0 1 Rs2[0]
rlabel metal2 6888 0 6900 0 1 Rs1[0]
rlabel metal2 6144 0 6156 0 1 Rw[0]
rlabel metal2 24458 0 24656 0 1 GND!
rlabel metal2 18792 0 18804 0 1 NAND
rlabel metal2 16248 0 16260 0 1 SUB
rlabel metal2 16416 0 16428 0 1 CIn_slice
rlabel metal2 16584 0 16596 0 1 LastCIn
rlabel metal2 16608 0 16620 0 1 COut
rlabel metal2 16896 0 16908 0 1 nZ
rlabel metal2 17040 0 17052 0 1 FAOut
rlabel metal2 17376 0 17388 0 1 AND
rlabel metal2 17736 0 17748 0 1 OR
rlabel metal2 18144 0 18156 0 1 XOR
rlabel metal2 18480 0 18492 0 1 NOT
rlabel metal2 19464 0 19476 0 1 ShL
rlabel metal2 19248 0 19260 0 1 ASign
rlabel metal2 19296 0 19308 0 1 ShB
rlabel metal2 19128 0 19140 0 1 NOR
rlabel metal2 21289 0 21301 0 1 ShR
rlabel metal2 23088 0 23100 0 1 ShOut
rlabel metal2 23256 0 23268 0 1 LLI
rlabel metal2 15984 0 15996 0 1 ZeroA
rlabel metal2 16680 0 16692 0 1 Flags[3]
rlabel metal2 21264 0 21276 0 1 Sh8
<< end >>
