magic
tech c035u
timestamp 1395354352
<< metal1 >>
rect 6912 44410 6922 44462
rect 6960 44410 6970 44462
rect 6912 44400 6970 44410
rect 5828 43440 5890 43450
rect 5880 43426 5890 43440
rect 6912 43429 6922 44400
rect 7008 43429 7018 44462
rect 11280 44266 11290 44462
rect 11328 44293 11338 44462
rect 15744 44437 15754 44462
rect 15792 44437 15802 44462
rect 20232 44437 20242 44462
rect 20280 44437 20290 44462
rect 20424 44437 20434 44462
rect 29160 44437 29170 44462
rect 29208 44437 29218 44462
rect 29352 44410 29362 44462
rect 33648 44437 33658 44462
rect 33696 44437 33706 44462
rect 33840 44437 33850 44462
rect 38112 44437 38122 44462
rect 12936 44400 29362 44410
rect 12936 44386 12946 44400
rect 38160 44410 38170 44462
rect 38304 44410 38314 44462
rect 29389 44400 38170 44410
rect 38184 44400 38314 44410
rect 12912 44376 12946 44386
rect 12912 44365 12922 44376
rect 12973 44376 29207 44386
rect 29245 44376 33647 44386
rect 33661 44376 38111 44386
rect 38184 44386 38194 44400
rect 38136 44376 38194 44386
rect 12936 44352 15791 44362
rect 12936 44338 12946 44352
rect 15829 44352 33839 44362
rect 38136 44362 38146 44376
rect 33864 44352 38146 44362
rect 12888 44328 12946 44338
rect 12888 44293 12898 44328
rect 12997 44328 33695 44338
rect 33864 44338 33874 44352
rect 33720 44328 33874 44338
rect 33720 44314 33730 44328
rect 12936 44304 33730 44314
rect 12936 44293 12946 44304
rect 13021 44280 29375 44290
rect 11280 44256 15743 44266
rect 11328 43429 11338 44231
rect 5880 43416 5903 43426
rect 12864 43402 12874 44256
rect 15781 44256 20231 44266
rect 20245 44256 29159 44266
rect 29173 44256 29231 44266
rect 13032 44232 20423 44242
rect 5828 43392 12874 43402
rect 5880 38317 5890 43392
rect 5904 38314 5914 43367
rect 6912 40042 6922 43367
rect 7008 40069 7018 43367
rect 11328 40069 11338 43367
rect 12888 40213 12898 44231
rect 12912 40213 12922 44231
rect 12936 40213 12946 44231
rect 12960 40186 12970 44231
rect 12984 40189 12994 44231
rect 13008 40189 13018 44231
rect 13032 40189 13042 44232
rect 13056 44208 20279 44218
rect 13056 40189 13066 44208
rect 13080 44184 15815 44194
rect 13080 40189 13090 44184
rect 13104 44160 15767 44170
rect 12853 40176 12970 40186
rect 12829 40152 12935 40162
rect 13104 40162 13114 44160
rect 38112 43621 38122 44327
rect 43776 43632 43840 43642
rect 43776 43621 43786 43632
rect 12960 40152 13114 40162
rect 13128 43584 43840 43594
rect 12960 40138 12970 40152
rect 12792 40128 12970 40138
rect 12792 40117 12802 40128
rect 13128 40138 13138 43584
rect 38112 43477 38122 43559
rect 43776 43477 43786 43559
rect 13104 40128 13138 40138
rect 13152 43440 43840 43450
rect 13080 40114 13090 40127
rect 13104 40117 13114 40128
rect 12864 40104 13090 40114
rect 12840 40090 12850 40103
rect 12864 40093 12874 40104
rect 13152 40114 13162 43440
rect 13141 40104 13162 40114
rect 12781 40080 12850 40090
rect 12936 40080 13162 40090
rect 12888 40066 12898 40079
rect 12936 40069 12946 40080
rect 12757 40056 12898 40066
rect 12973 40056 13055 40066
rect 13080 40056 13103 40066
rect 6912 40032 13055 40042
rect 12709 40008 12815 40018
rect 13080 40018 13090 40056
rect 13128 40042 13138 40055
rect 12853 40008 13090 40018
rect 13104 40032 13138 40042
rect 7008 39809 7018 40007
rect 11328 39833 11338 40007
rect 12672 39984 12743 39994
rect 12672 39857 12682 39984
rect 13104 39994 13114 40032
rect 12829 39984 13114 39994
rect 12720 39960 13031 39970
rect 12720 39920 12730 39960
rect 12744 39936 13007 39946
rect 12744 39920 12754 39936
rect 12888 39912 12983 39922
rect 12888 39902 12898 39912
rect 13056 39922 13066 39959
rect 13152 39946 13162 40080
rect 13152 39936 13258 39946
rect 13248 39922 13258 39936
rect 38112 39922 38122 43415
rect 43776 39922 43786 43415
rect 13056 39912 13234 39922
rect 13248 39912 13354 39922
rect 38112 39912 43786 39922
rect 13224 39901 13234 39912
rect 13344 39901 13354 39912
rect 12672 39847 12983 39857
rect 40237 39847 40402 39857
rect 11328 39823 12983 39833
rect 7008 39799 12983 39809
rect 40237 39799 40343 39809
rect 40237 39775 40378 39785
rect 5904 38304 5938 38314
rect 5828 38280 5914 38290
rect 5880 38242 5890 38255
rect 5828 38232 5890 38242
rect 5880 33157 5890 38232
rect 5904 35232 5914 38280
rect 5928 35256 5938 38304
rect 12696 35317 12706 39767
rect 12720 35317 12730 39767
rect 12744 35317 12754 39767
rect 12768 35317 12778 39767
rect 12792 35317 12802 39767
rect 12816 35317 12826 39767
rect 12840 35317 12850 39767
rect 12864 35317 12874 39767
rect 12888 35317 12898 39767
rect 12912 35317 12922 39767
rect 12936 35290 12946 39767
rect 12960 35293 12970 39767
rect 40237 39751 40330 39761
rect 40237 39727 40306 39737
rect 40237 39703 40282 39713
rect 40237 39679 40258 39689
rect 40248 36517 40258 39679
rect 40272 36514 40282 39703
rect 40296 36541 40306 39727
rect 40320 36541 40330 39751
rect 40344 36541 40354 39743
rect 40368 36541 40378 39775
rect 40392 36541 40402 39847
rect 43776 38482 43786 39912
rect 43776 38472 43840 38482
rect 43776 38461 43786 38472
rect 43752 38424 43840 38434
rect 43752 38341 43762 38424
rect 43776 38314 43786 38399
rect 43728 38304 43786 38314
rect 40272 36504 40426 36514
rect 40237 36480 40282 36490
rect 12685 35280 12946 35290
rect 5928 35246 12983 35256
rect 5904 35222 12983 35232
rect 12949 35199 12983 35209
rect 12672 33130 12682 35197
rect 5828 33120 12682 33130
rect 5880 33082 5890 33095
rect 5828 33072 5890 33082
rect 5880 30922 5890 33072
rect 12696 31885 12706 35197
rect 12720 31885 12730 35197
rect 12744 31858 12754 35197
rect 12768 31861 12778 35197
rect 12792 35184 12802 35197
rect 12792 35174 12983 35184
rect 12792 31861 12802 35174
rect 12816 31861 12826 35141
rect 12840 31861 12850 35141
rect 12864 31861 12874 35141
rect 12685 31848 12754 31858
rect 12888 31834 12898 35141
rect 12912 31837 12922 35141
rect 12936 31837 12946 35141
rect 12960 31837 12970 35141
rect 40248 33709 40258 36455
rect 40272 33709 40282 36480
rect 40296 33706 40306 36479
rect 40320 33733 40330 36479
rect 40344 33733 40354 36479
rect 40368 33733 40378 36479
rect 40392 33733 40402 36479
rect 40416 33733 40426 36504
rect 40296 33696 40439 33706
rect 40237 33663 40295 33673
rect 40357 33672 40474 33682
rect 40237 33639 40354 33649
rect 12661 31824 12898 31834
rect 12637 31800 12863 31810
rect 12901 31800 12983 31810
rect 12600 31776 12839 31786
rect 12600 31522 12610 31776
rect 12877 31776 12983 31786
rect 40248 31765 40258 33611
rect 40272 31765 40282 33611
rect 12744 31752 12983 31762
rect 12624 31525 12634 31751
rect 12648 31525 12658 31751
rect 12672 31525 12682 31751
rect 12696 31525 12706 31751
rect 12720 31525 12730 31751
rect 12744 31525 12754 31752
rect 40296 31762 40306 33611
rect 40320 31789 40330 33611
rect 40344 31786 40354 33639
rect 40368 31813 40378 33647
rect 40392 31810 40402 33647
rect 40416 31837 40426 33647
rect 40440 31837 40450 33647
rect 40464 31837 40474 33672
rect 43728 33322 43738 38304
rect 43776 38280 43840 38290
rect 43752 33349 43762 38279
rect 43776 33349 43786 38280
rect 43728 33312 43840 33322
rect 43728 33301 43738 33312
rect 43704 33264 43840 33274
rect 43704 33157 43714 33264
rect 43728 33157 43738 33239
rect 43752 33157 43762 33239
rect 43776 33157 43786 33239
rect 43680 33120 43840 33130
rect 40392 31800 40487 31810
rect 40344 31776 40511 31786
rect 40296 31752 40546 31762
rect 40536 31741 40546 31752
rect 12840 31728 12983 31738
rect 12768 31525 12778 31727
rect 12792 31525 12802 31727
rect 12816 31525 12826 31727
rect 12840 31525 12850 31728
rect 40237 31728 40402 31738
rect 40392 31717 40402 31728
rect 12864 31546 12874 31703
rect 12888 31573 12898 31703
rect 12912 31573 12922 31703
rect 12936 31573 12946 31703
rect 12960 31573 12970 31703
rect 40237 31704 40343 31714
rect 40464 31714 40474 31727
rect 40464 31704 40559 31714
rect 40237 31680 40463 31690
rect 40501 31680 40594 31690
rect 40584 31669 40594 31680
rect 40237 31656 40487 31666
rect 40237 31632 40618 31642
rect 40237 31608 40295 31618
rect 40608 31618 40618 31632
rect 40608 31608 40631 31618
rect 43680 31597 43690 33120
rect 40261 31584 40679 31594
rect 43704 31570 43714 33095
rect 40261 31560 43714 31570
rect 12864 31536 12983 31546
rect 24480 31546 24490 31559
rect 13021 31536 24490 31546
rect 24504 31536 27575 31546
rect 24504 31525 24514 31536
rect 27613 31536 40271 31546
rect 12552 31512 12610 31522
rect 12552 31501 12562 31512
rect 12877 31512 24479 31522
rect 40320 31522 40330 31535
rect 24541 31512 40330 31522
rect 40392 31498 40402 31535
rect 12589 31488 40402 31498
rect 12541 31464 12719 31474
rect 12853 31464 13055 31474
rect 13093 31464 23423 31474
rect 23485 31464 40367 31474
rect 12517 31440 12671 31450
rect 12733 31440 13369 31450
rect 13408 31440 13463 31450
rect 13501 31440 20471 31450
rect 20509 31440 38159 31450
rect 12493 31416 12743 31426
rect 12853 31416 23423 31426
rect 40416 31426 40426 31535
rect 23461 31416 40426 31426
rect 12469 31392 12647 31402
rect 12685 31392 21959 31402
rect 40440 31402 40450 31535
rect 21997 31392 40450 31402
rect 40464 31381 40474 31535
rect 12445 31368 12767 31378
rect 12901 31368 13103 31378
rect 13141 31368 32246 31378
rect 32317 31368 33743 31378
rect 35221 31368 38111 31378
rect 12408 31344 12551 31354
rect 12408 31309 12418 31344
rect 40488 31354 40498 31535
rect 12613 31344 40498 31354
rect 40512 31333 40522 31535
rect 12552 31320 40463 31330
rect 12552 31309 12562 31320
rect 40536 31306 40546 31535
rect 12661 31296 40546 31306
rect 12397 31272 12815 31282
rect 12901 31272 30791 31282
rect 30829 31272 40511 31282
rect 12360 31248 12647 31258
rect 12360 31237 12370 31248
rect 12757 31248 24935 31258
rect 24960 31248 26423 31258
rect 24960 31237 24970 31248
rect 26461 31248 32270 31258
rect 37765 31248 38087 31258
rect 12648 31224 24935 31234
rect 12504 31210 12514 31223
rect 12648 31213 12658 31224
rect 40560 31234 40570 31535
rect 24997 31224 40570 31234
rect 12349 31200 12514 31210
rect 12768 31200 29327 31210
rect 12696 31186 12706 31199
rect 12768 31189 12778 31200
rect 40584 31210 40594 31535
rect 40632 31213 40642 31535
rect 40680 31213 40690 31535
rect 43680 31213 43690 31535
rect 43728 31213 43738 33095
rect 43752 31213 43762 33095
rect 29365 31200 40594 31210
rect 12325 31176 12706 31186
rect 12829 31176 13394 31186
rect 43776 31186 43786 33095
rect 13512 31176 43786 31186
rect 12277 31152 12455 31162
rect 12517 31152 13426 31162
rect 13416 31141 13426 31152
rect 13464 31141 13474 31175
rect 13488 31141 13498 31175
rect 13512 31141 13522 31176
rect 13536 31152 40631 31162
rect 12240 31128 12623 31138
rect 12240 31093 12250 31128
rect 12709 31128 13391 31138
rect 13536 31114 13546 31152
rect 43752 31138 43762 31151
rect 13621 31128 43762 31138
rect 12288 31104 13546 31114
rect 13560 31104 19007 31114
rect 12288 31093 12298 31104
rect 12469 31080 13511 31090
rect 13560 31090 13570 31104
rect 19045 31104 23471 31114
rect 23509 31104 26447 31114
rect 26472 31104 29327 31114
rect 13549 31080 13570 31090
rect 26472 31090 26482 31104
rect 29389 31104 40679 31114
rect 13597 31080 26482 31090
rect 27589 31080 32303 31090
rect 12216 31056 12479 31066
rect 12216 31018 12226 31056
rect 12637 31056 13127 31066
rect 43680 31066 43690 31103
rect 13189 31056 43690 31066
rect 12493 31032 13607 31042
rect 17160 31032 23447 31042
rect 12216 31008 13127 31018
rect 13152 31008 13535 31018
rect 12216 30984 12527 30994
rect 12216 30949 12226 30984
rect 13152 30994 13162 31008
rect 13560 31008 13583 31018
rect 13045 30984 13162 30994
rect 13406 30984 13487 30994
rect 13560 30994 13570 31008
rect 13512 30984 13570 30994
rect 13176 30970 13186 30983
rect 12528 30960 13186 30970
rect 12528 30949 12538 30960
rect 5880 30912 13162 30922
rect 12216 30637 12226 30887
rect 12240 30637 12250 30887
rect 12264 30637 12274 30887
rect 12288 30637 12298 30887
rect 12312 30637 12322 30887
rect 12336 30637 12346 30887
rect 12360 30637 12370 30887
rect 12384 30637 12394 30887
rect 12408 30637 12418 30887
rect 12432 30610 12442 30887
rect 12456 30613 12466 30887
rect 12480 30613 12490 30887
rect 12504 30613 12514 30887
rect 12528 30613 12538 30887
rect 12552 30613 12562 30887
rect 12576 30613 12586 30887
rect 12600 30613 12610 30887
rect 12624 30613 12634 30887
rect 12648 30613 12658 30887
rect 12672 30613 12682 30887
rect 12696 30613 12706 30887
rect 12720 30613 12730 30887
rect 12744 30613 12754 30887
rect 12768 30613 12778 30887
rect 12792 30613 12802 30887
rect 12816 30613 12826 30887
rect 12840 30613 12850 30887
rect 12864 30613 12874 30887
rect 12888 30613 12898 30887
rect 12205 30600 12442 30610
rect 12912 30586 12922 30887
rect 12936 30589 12946 30887
rect 12960 30589 12970 30887
rect 12984 30589 12994 30887
rect 13008 30589 13018 30887
rect 13032 30589 13042 30887
rect 13056 30589 13066 30887
rect 12181 30576 12922 30586
rect 12157 30552 12599 30562
rect 13080 30562 13090 30887
rect 12925 30552 13090 30562
rect 12120 30528 12959 30538
rect 12120 30517 12130 30528
rect 12997 30528 13079 30538
rect 13104 30538 13114 30887
rect 13128 30562 13138 30887
rect 13152 30586 13162 30912
rect 13224 30610 13234 30983
rect 13344 30634 13354 30959
rect 13368 30658 13378 30983
rect 13512 30970 13522 30984
rect 13429 30960 13522 30970
rect 13440 30682 13450 30935
rect 13464 30706 13474 30935
rect 13464 30696 13487 30706
rect 13440 30672 13681 30682
rect 13368 30648 13633 30658
rect 13623 30637 13633 30648
rect 13344 30624 13598 30634
rect 13671 30613 13681 30672
rect 13224 30600 13463 30610
rect 13501 30600 13646 30610
rect 15432 30610 15442 31031
rect 17160 30637 17170 31032
rect 23485 31032 23495 31042
rect 23520 31032 24527 31042
rect 23520 31018 23530 31032
rect 24552 31032 24983 31042
rect 24552 31018 24562 31032
rect 27576 31032 27599 31042
rect 17400 31008 23530 31018
rect 23544 31008 24562 31018
rect 17400 30637 17410 31008
rect 17533 30984 20495 30994
rect 20520 30984 21983 30994
rect 18360 30960 19031 30970
rect 18360 30637 18370 30960
rect 20520 30970 20530 30984
rect 23544 30994 23554 31008
rect 24949 31008 24959 31018
rect 22008 30984 23554 30994
rect 22008 30970 22018 30984
rect 24493 30984 24503 30994
rect 19056 30960 20530 30970
rect 20544 30960 22018 30970
rect 19056 30946 19066 30960
rect 20544 30946 20554 30960
rect 23437 30960 23471 30970
rect 18552 30936 19066 30946
rect 19584 30936 20554 30946
rect 18552 30637 18562 30936
rect 19584 30637 19594 30936
rect 27576 30637 27586 31032
rect 27840 31032 29375 31042
rect 27840 30637 27850 31032
rect 29400 31032 30815 31042
rect 28560 31008 29351 31018
rect 28560 30637 28570 31008
rect 29400 31018 29410 31032
rect 29376 31008 29410 31018
rect 29376 30994 29386 31008
rect 29341 30984 29386 30994
rect 38088 30946 38098 31031
rect 38112 30973 38122 31031
rect 38136 30973 38146 31031
rect 38160 30973 38170 31031
rect 38088 30936 38183 30946
rect 39960 30922 39970 31031
rect 37920 30912 39970 30922
rect 15432 30600 30418 30610
rect 30408 30586 30418 30600
rect 13152 30576 30394 30586
rect 30408 30576 30610 30586
rect 13128 30552 30359 30562
rect 30384 30562 30394 30576
rect 30600 30562 30610 30576
rect 30384 30552 30586 30562
rect 30600 30552 30671 30562
rect 13104 30528 30551 30538
rect 30576 30538 30586 30552
rect 37920 30541 37930 30912
rect 38088 30541 38098 30912
rect 38112 30541 38122 30887
rect 38136 30541 38146 30887
rect 38160 30541 38170 30887
rect 38184 30541 38194 30887
rect 40248 30541 40258 31031
rect 40296 30541 40306 31031
rect 30576 30528 30743 30538
rect 40344 30514 40354 31031
rect 12432 30504 40354 30514
rect 12216 30490 12226 30503
rect 12432 30493 12442 30504
rect 12096 30480 12226 30490
rect 12096 30469 12106 30480
rect 12613 30480 13031 30490
rect 13093 30480 30623 30490
rect 30661 30480 30719 30490
rect 30757 30480 37919 30490
rect 38101 30480 38207 30490
rect 40296 30466 40306 30479
rect 12229 30456 40306 30466
rect 12072 30432 12551 30442
rect 5828 28008 5890 28018
rect 5880 22981 5890 28008
rect 12072 27658 12082 30432
rect 12973 30432 13007 30442
rect 13069 30432 30647 30442
rect 30685 30432 38087 30442
rect 40248 30418 40258 30431
rect 12552 30408 40258 30418
rect 12096 27685 12106 30407
rect 12120 27685 12130 30407
rect 12144 27685 12154 30407
rect 12168 27685 12178 30407
rect 12192 27685 12202 30407
rect 12216 27685 12226 30407
rect 12240 27685 12250 30407
rect 12264 27685 12274 30407
rect 12288 27685 12298 30407
rect 12312 27685 12322 30407
rect 12336 27685 12346 30407
rect 12360 27685 12370 30407
rect 12384 27685 12394 30407
rect 12408 27685 12418 30407
rect 12432 27685 12442 30407
rect 12456 27685 12466 30407
rect 12480 27685 12490 30407
rect 12504 27685 12514 30407
rect 12528 27685 12538 30407
rect 12552 27685 12562 30408
rect 12576 27685 12586 30383
rect 12600 27685 12610 30383
rect 12624 27685 12634 30383
rect 12648 27685 12658 30383
rect 12672 27685 12682 30383
rect 12696 27685 12706 30383
rect 12720 27685 12730 30383
rect 12744 27685 12754 30383
rect 12768 27685 12778 30383
rect 12792 27685 12802 30383
rect 12816 27685 12826 30383
rect 12840 27685 12850 30383
rect 12864 27685 12874 30383
rect 12888 27685 12898 30383
rect 12912 27685 12922 30383
rect 12936 27685 12946 30383
rect 12960 27685 12970 30383
rect 12072 27652 12994 27658
rect 12072 27648 13008 27652
rect 12984 27642 13008 27648
rect 12096 27610 12106 27623
rect 12984 27610 13008 27620
rect 12096 27600 12994 27610
rect 12133 27576 13008 27586
rect 12144 26482 12154 27551
rect 12168 26509 12178 27551
rect 12192 26509 12202 27551
rect 12216 26509 12226 27551
rect 12240 26509 12250 27551
rect 12264 26509 12274 27551
rect 12288 26509 12298 27551
rect 12312 26509 12322 27551
rect 12336 26509 12346 27551
rect 12360 26509 12370 27551
rect 12384 26509 12394 27551
rect 12408 26509 12418 27551
rect 12432 26509 12442 27551
rect 12456 26509 12466 27551
rect 12480 26509 12490 27551
rect 12504 26509 12514 27551
rect 12528 26509 12538 27551
rect 12552 26509 12562 27551
rect 12576 26509 12586 27551
rect 12600 26509 12610 27551
rect 12624 26509 12634 27551
rect 12648 26509 12658 27551
rect 12672 26509 12682 27551
rect 12696 26509 12706 27551
rect 12720 26509 12730 27551
rect 12744 26509 12754 27551
rect 12768 26509 12778 27551
rect 12792 26509 12802 27551
rect 12816 26509 12826 27551
rect 12840 26509 12850 27551
rect 12864 26509 12874 27551
rect 12888 26509 12898 27551
rect 12912 26509 12922 27551
rect 12936 26509 12946 27551
rect 12960 26509 12970 27551
rect 12144 26476 12994 26482
rect 12144 26472 13008 26476
rect 12984 26466 13008 26472
rect 12168 26434 12178 26447
rect 12984 26434 13008 26444
rect 12168 26424 12994 26434
rect 12205 26400 13008 26410
rect 12216 25306 12226 26375
rect 12240 25333 12250 26375
rect 12264 25333 12274 26375
rect 12288 25333 12298 26375
rect 12312 25333 12322 26375
rect 12336 25333 12346 26375
rect 12360 25333 12370 26375
rect 12384 25333 12394 26375
rect 12408 25333 12418 26375
rect 12432 25333 12442 26375
rect 12456 25333 12466 26375
rect 12480 25333 12490 26375
rect 12504 25333 12514 26375
rect 12528 25333 12538 26375
rect 12552 25333 12562 26375
rect 12576 25333 12586 26375
rect 12600 25333 12610 26375
rect 12624 25333 12634 26375
rect 12648 25333 12658 26375
rect 12672 25333 12682 26375
rect 12696 25333 12706 26375
rect 12720 25333 12730 26375
rect 12744 25333 12754 26375
rect 12768 25333 12778 26375
rect 12792 25333 12802 26375
rect 12816 25333 12826 26375
rect 12840 25333 12850 26375
rect 12864 25333 12874 26375
rect 12888 25333 12898 26375
rect 12912 25333 12922 26375
rect 12936 25333 12946 26375
rect 12960 25333 12970 26375
rect 12216 25300 12994 25306
rect 12216 25296 13008 25300
rect 12984 25290 13008 25296
rect 12240 25258 12250 25271
rect 12984 25258 13008 25268
rect 12240 25248 12994 25258
rect 12277 25224 13008 25234
rect 12288 24130 12298 25199
rect 12312 24157 12322 25199
rect 12336 24157 12346 25199
rect 12360 24157 12370 25199
rect 12384 24157 12394 25199
rect 12408 24157 12418 25199
rect 12432 24157 12442 25199
rect 12456 24157 12466 25199
rect 12480 24157 12490 25199
rect 12504 24157 12514 25199
rect 12528 24157 12538 25199
rect 12552 24157 12562 25199
rect 12576 24157 12586 25199
rect 12600 24157 12610 25199
rect 12624 24157 12634 25199
rect 12648 24157 12658 25199
rect 12672 24157 12682 25199
rect 12696 24157 12706 25199
rect 12720 24157 12730 25199
rect 12744 24157 12754 25199
rect 12768 24157 12778 25199
rect 12792 24157 12802 25199
rect 12816 24157 12826 25199
rect 12840 24157 12850 25199
rect 12864 24157 12874 25199
rect 12888 24157 12898 25199
rect 12912 24157 12922 25199
rect 12936 24157 12946 25199
rect 12960 24157 12970 25199
rect 12288 24124 12994 24130
rect 12288 24120 13008 24124
rect 12984 24114 13008 24120
rect 12312 24082 12322 24095
rect 12984 24082 13008 24092
rect 12312 24072 12994 24082
rect 12349 24048 13008 24058
rect 12360 22954 12370 24023
rect 12384 22981 12394 24023
rect 12408 22981 12418 24023
rect 12432 22981 12442 24023
rect 12456 22981 12466 24023
rect 12480 22981 12490 24023
rect 12504 22981 12514 24023
rect 12528 22981 12538 24023
rect 12552 22981 12562 24023
rect 12576 22981 12586 24023
rect 12600 22981 12610 24023
rect 12624 22981 12634 24023
rect 12648 22981 12658 24023
rect 12672 22981 12682 24023
rect 12696 22981 12706 24023
rect 12720 22981 12730 24023
rect 12744 22981 12754 24023
rect 12768 22981 12778 24023
rect 12792 22981 12802 24023
rect 12816 22981 12826 24023
rect 12840 22981 12850 24023
rect 12864 22981 12874 24023
rect 12888 22981 12898 24023
rect 12912 22981 12922 24023
rect 12936 22981 12946 24023
rect 12960 22981 12970 24023
rect 5828 22944 5914 22954
rect 12360 22948 12994 22954
rect 12360 22944 13008 22948
rect 5880 17821 5890 22919
rect 5904 17821 5914 22944
rect 12984 22938 13008 22944
rect 12384 22906 12394 22919
rect 12984 22906 13008 22916
rect 12384 22896 12994 22906
rect 12421 22872 13008 22882
rect 12432 21778 12442 22847
rect 12456 21805 12466 22847
rect 12480 21805 12490 22847
rect 12504 21805 12514 22847
rect 12528 21805 12538 22847
rect 12552 21805 12562 22847
rect 12576 21805 12586 22847
rect 12600 21805 12610 22847
rect 12624 21805 12634 22847
rect 12648 21805 12658 22847
rect 12672 21805 12682 22847
rect 12696 21805 12706 22847
rect 12720 21805 12730 22847
rect 12744 21805 12754 22847
rect 12768 21805 12778 22847
rect 12792 21805 12802 22847
rect 12816 21805 12826 22847
rect 12840 21805 12850 22847
rect 12864 21805 12874 22847
rect 12888 21805 12898 22847
rect 12912 21805 12922 22847
rect 12936 21805 12946 22847
rect 12960 21805 12970 22847
rect 12432 21772 12994 21778
rect 12432 21768 13008 21772
rect 12984 21762 13008 21768
rect 12456 21730 12466 21743
rect 12984 21730 13008 21740
rect 12456 21720 12994 21730
rect 12493 21696 13008 21706
rect 12504 20602 12514 21671
rect 12528 20629 12538 21671
rect 12552 20629 12562 21671
rect 12576 20629 12586 21671
rect 12600 20629 12610 21671
rect 12624 20629 12634 21671
rect 12648 20629 12658 21671
rect 12672 20629 12682 21671
rect 12696 20629 12706 21671
rect 12720 20629 12730 21671
rect 12744 20629 12754 21671
rect 12768 20629 12778 21671
rect 12792 20629 12802 21671
rect 12816 20629 12826 21671
rect 12840 20629 12850 21671
rect 12864 20629 12874 21671
rect 12888 20629 12898 21671
rect 12912 20629 12922 21671
rect 12936 20629 12946 21671
rect 12960 20629 12970 21671
rect 12504 20596 12994 20602
rect 12504 20592 13008 20596
rect 12984 20586 13008 20592
rect 12528 20554 12538 20567
rect 12984 20554 13008 20564
rect 12528 20544 12994 20554
rect 12565 20520 13008 20530
rect 12576 19426 12586 20495
rect 12600 19453 12610 20495
rect 12624 19453 12634 20495
rect 12648 19453 12658 20495
rect 12672 19453 12682 20495
rect 12696 19453 12706 20495
rect 12720 19453 12730 20495
rect 12744 19453 12754 20495
rect 12768 19453 12778 20495
rect 12792 19453 12802 20495
rect 12816 19453 12826 20495
rect 12840 19453 12850 20495
rect 12864 19453 12874 20495
rect 12888 19453 12898 20495
rect 12912 19453 12922 20495
rect 12936 19453 12946 20495
rect 12960 19453 12970 20495
rect 12576 19420 12994 19426
rect 12576 19416 13008 19420
rect 12984 19410 13008 19416
rect 12589 19392 12887 19402
rect 12552 19368 12671 19378
rect 12552 18253 12562 19368
rect 12984 19378 13008 19388
rect 12901 19368 12994 19378
rect 12672 19344 13008 19354
rect 12576 18253 12586 19343
rect 12600 18253 12610 19343
rect 12624 18253 12634 19343
rect 12648 18253 12658 19343
rect 12672 18253 12682 19344
rect 12696 18253 12706 19319
rect 12720 18253 12730 19319
rect 12744 18226 12754 19319
rect 12768 18229 12778 19319
rect 12792 18229 12802 19319
rect 12816 18229 12826 19319
rect 12840 18229 12850 19319
rect 12864 18229 12874 19319
rect 12888 18229 12898 19319
rect 12912 18229 12922 19319
rect 12936 18229 12946 19319
rect 12960 18229 12970 19319
rect 12541 18216 12754 18226
rect 12504 18192 12719 18202
rect 12504 17794 12514 18192
rect 12984 18202 13008 18212
rect 12757 18192 12994 18202
rect 12720 18168 13008 18178
rect 5828 17784 12514 17794
rect 5880 12661 5890 17759
rect 5904 12661 5914 17759
rect 12528 17077 12538 18167
rect 12552 17077 12562 18167
rect 12576 17077 12586 18167
rect 12600 17077 12610 18167
rect 12624 17077 12634 18167
rect 12648 17077 12658 18167
rect 12672 17077 12682 18167
rect 12696 17077 12706 18167
rect 12720 17077 12730 18168
rect 12744 17077 12754 18143
rect 12768 17077 12778 18143
rect 12792 17077 12802 18143
rect 12816 17077 12826 18143
rect 12840 17077 12850 18143
rect 12864 17077 12874 18143
rect 12888 17077 12898 18143
rect 12912 17050 12922 18143
rect 12936 17053 12946 18143
rect 12960 17053 12970 18143
rect 12517 17040 12922 17050
rect 12480 17016 12839 17026
rect 12480 15901 12490 17016
rect 12984 17026 13008 17036
rect 12925 17016 12994 17026
rect 12840 16992 13008 17002
rect 12504 15901 12514 16991
rect 12528 15901 12538 16991
rect 12552 15901 12562 16991
rect 12576 15901 12586 16991
rect 12600 15901 12610 16991
rect 12624 15901 12634 16991
rect 12648 15901 12658 16991
rect 12672 15901 12682 16991
rect 12696 15901 12706 16991
rect 12720 15901 12730 16991
rect 12744 15901 12754 16991
rect 12768 15901 12778 16991
rect 12792 15901 12802 16991
rect 12816 15901 12826 16991
rect 12840 15901 12850 16992
rect 12864 15901 12874 16967
rect 12888 15901 12898 16967
rect 12912 15874 12922 16967
rect 12936 15877 12946 16967
rect 12960 15877 12970 16967
rect 12469 15864 12922 15874
rect 12432 15840 12863 15850
rect 12432 14749 12442 15840
rect 12984 15850 13008 15860
rect 12925 15840 12994 15850
rect 12864 15816 13008 15826
rect 12456 14749 12466 15815
rect 12480 14749 12490 15815
rect 12504 14749 12514 15815
rect 12528 14749 12538 15815
rect 12552 14749 12562 15815
rect 12576 14749 12586 15815
rect 12600 14749 12610 15815
rect 12624 14749 12634 15815
rect 12648 14749 12658 15815
rect 12672 14749 12682 15815
rect 12696 14749 12706 15815
rect 12720 14749 12730 15815
rect 12744 14749 12754 15815
rect 12768 14749 12778 15815
rect 12792 14749 12802 15815
rect 12816 14749 12826 15815
rect 12840 14749 12850 15815
rect 12864 14749 12874 15816
rect 12888 14722 12898 15791
rect 12912 14725 12922 15791
rect 12936 14725 12946 15791
rect 12421 14712 12898 14722
rect 12960 14698 12970 15791
rect 12384 14688 12970 14698
rect 12384 13549 12394 14688
rect 12984 14674 13008 14684
rect 12888 14664 12994 14674
rect 12408 13549 12418 14663
rect 12432 13549 12442 14663
rect 12456 13549 12466 14663
rect 12480 13549 12490 14663
rect 12504 13549 12514 14663
rect 12528 13549 12538 14663
rect 12552 13549 12562 14663
rect 12576 13549 12586 14663
rect 12600 13549 12610 14663
rect 12624 13549 12634 14663
rect 12648 13549 12658 14663
rect 12672 13549 12682 14663
rect 12696 13549 12706 14663
rect 12720 13549 12730 14663
rect 12744 13549 12754 14663
rect 12768 13549 12778 14663
rect 12792 13549 12802 14663
rect 12816 13549 12826 14663
rect 12840 13549 12850 14663
rect 12864 13522 12874 14663
rect 12888 13525 12898 14664
rect 12960 14640 13008 14650
rect 12912 13525 12922 14639
rect 12936 13525 12946 14639
rect 12960 13525 12970 14640
rect 12373 13512 12874 13522
rect 12336 13488 12815 13498
rect 12336 12634 12346 13488
rect 12984 13498 13008 13508
rect 12877 13488 12994 13498
rect 12816 13464 13008 13474
rect 5828 12624 12346 12634
rect 5880 7501 5890 12599
rect 5904 9202 5914 12599
rect 12360 12397 12370 13463
rect 12384 12397 12394 13463
rect 12408 12370 12418 13463
rect 12432 12373 12442 13463
rect 12456 12373 12466 13463
rect 12480 12373 12490 13463
rect 12504 12373 12514 13463
rect 12528 12373 12538 13463
rect 12552 12373 12562 13463
rect 12576 12373 12586 13463
rect 12600 12373 12610 13463
rect 12624 12373 12634 13463
rect 12648 12373 12658 13463
rect 12672 12373 12682 13463
rect 12696 12373 12706 13463
rect 12720 12373 12730 13463
rect 12744 12373 12754 13463
rect 12768 12373 12778 13463
rect 12792 12373 12802 13463
rect 12816 12373 12826 13464
rect 12840 12373 12850 13439
rect 12864 12373 12874 13439
rect 12349 12360 12418 12370
rect 12888 12346 12898 13439
rect 12912 12349 12922 13439
rect 12936 12349 12946 13439
rect 12960 12349 12970 13439
rect 12312 12336 12898 12346
rect 12312 11197 12322 12336
rect 12984 12322 13008 12332
rect 12408 12312 12994 12322
rect 12336 11170 12346 12311
rect 12360 11173 12370 12311
rect 12384 11173 12394 12311
rect 12408 11173 12418 12312
rect 12888 12288 13008 12298
rect 12432 11173 12442 12287
rect 12456 11173 12466 12287
rect 12480 11173 12490 12287
rect 12504 11173 12514 12287
rect 12528 11173 12538 12287
rect 12552 11173 12562 12287
rect 12576 11173 12586 12287
rect 12600 11173 12610 12287
rect 12624 11173 12634 12287
rect 12648 11173 12658 12287
rect 12672 11173 12682 12287
rect 12696 11173 12706 12287
rect 12720 11173 12730 12287
rect 12744 11173 12754 12287
rect 12768 11173 12778 12287
rect 12792 11173 12802 12287
rect 12816 11173 12826 12287
rect 12840 11173 12850 12287
rect 12864 11173 12874 12287
rect 12888 11173 12898 12288
rect 12912 11173 12922 12263
rect 12936 11173 12946 12263
rect 12960 11173 12970 12263
rect 12288 11160 12346 11170
rect 12288 11146 12298 11160
rect 12264 11136 12298 11146
rect 12264 10021 12274 11136
rect 12984 11146 13008 11156
rect 12349 11136 12994 11146
rect 12288 11112 13008 11122
rect 12288 10021 12298 11112
rect 12312 10021 12322 11087
rect 12336 10021 12346 11087
rect 12360 10021 12370 11087
rect 12384 10021 12394 11087
rect 12408 10021 12418 11087
rect 12432 10021 12442 11087
rect 12456 10021 12466 11087
rect 12480 10021 12490 11087
rect 12504 10021 12514 11087
rect 12528 10021 12538 11087
rect 12552 10021 12562 11087
rect 12576 10021 12586 11087
rect 12600 10021 12610 11087
rect 12624 10021 12634 11087
rect 12648 10021 12658 11087
rect 12672 10021 12682 11087
rect 12696 10021 12706 11087
rect 12720 10021 12730 11087
rect 12744 10021 12754 11087
rect 12768 10021 12778 11087
rect 12792 10021 12802 11087
rect 12816 10021 12826 11087
rect 12840 10021 12850 11087
rect 12864 10021 12874 11087
rect 12888 9994 12898 11087
rect 12912 9997 12922 11087
rect 12936 9997 12946 11087
rect 12960 9997 12970 11087
rect 12253 9984 12898 9994
rect 12216 9960 12839 9970
rect 12216 9754 12226 9960
rect 12984 9970 13008 9980
rect 12901 9960 12994 9970
rect 12840 9936 13008 9946
rect 12240 9781 12250 9935
rect 12264 9781 12274 9935
rect 12288 9781 12298 9935
rect 12312 9781 12322 9935
rect 12336 9781 12346 9935
rect 12360 9781 12370 9935
rect 12384 9781 12394 9935
rect 12408 9781 12418 9935
rect 12432 9781 12442 9935
rect 12456 9781 12466 9935
rect 12480 9781 12490 9935
rect 12504 9781 12514 9935
rect 12528 9781 12538 9935
rect 12552 9781 12562 9935
rect 12576 9781 12586 9935
rect 12600 9781 12610 9935
rect 12624 9781 12634 9935
rect 12648 9781 12658 9935
rect 12672 9781 12682 9935
rect 12696 9781 12706 9935
rect 12720 9781 12730 9935
rect 12744 9781 12754 9935
rect 12768 9781 12778 9935
rect 12792 9781 12802 9935
rect 12816 9781 12826 9935
rect 12840 9781 12850 9936
rect 12864 9781 12874 9911
rect 12888 9781 12898 9911
rect 12912 9781 12922 9911
rect 12936 9781 12946 9911
rect 12960 9781 12970 9911
rect 38088 9781 38098 30383
rect 38112 9778 38122 30383
rect 38136 9805 38146 30383
rect 38160 9805 38170 30383
rect 38184 9805 38194 30383
rect 38208 28042 38218 30383
rect 43728 28069 43738 31103
rect 38208 28032 43799 28042
rect 43728 17842 43738 28007
rect 43728 17832 43840 17842
rect 43776 17821 43786 17832
rect 43752 17784 43840 17794
rect 43752 17677 43762 17784
rect 43776 17677 43786 17759
rect 43728 17640 43840 17650
rect 43728 12661 43738 17640
rect 43752 12661 43762 17615
rect 43776 12682 43786 17615
rect 43776 12672 43840 12682
rect 43776 12661 43786 12672
rect 43704 12624 43840 12634
rect 43704 12541 43714 12624
rect 43728 12514 43738 12599
rect 43752 12517 43762 12599
rect 43776 12517 43786 12599
rect 43680 12504 43738 12514
rect 38112 9768 38218 9778
rect 12216 9744 38111 9754
rect 12253 9720 13007 9730
rect 13117 9720 15983 9730
rect 38208 9730 38218 9768
rect 16021 9720 38218 9730
rect 43680 9706 43690 12504
rect 43728 12480 43840 12490
rect 12277 9696 43690 9706
rect 12301 9672 13031 9682
rect 13128 9672 13463 9682
rect 12325 9648 13055 9658
rect 13104 9637 13114 9671
rect 13128 9637 13138 9672
rect 13501 9672 13679 9682
rect 13717 9672 15959 9682
rect 16045 9672 38183 9682
rect 13152 9648 13607 9658
rect 13152 9637 13162 9648
rect 13645 9648 17999 9658
rect 18037 9648 29159 9658
rect 36877 9648 38159 9658
rect 12349 9624 13079 9634
rect 13189 9624 28919 9634
rect 37621 9624 38087 9634
rect 38125 9624 38170 9634
rect 38160 9613 38170 9624
rect 12373 9600 38087 9610
rect 38125 9600 38135 9610
rect 12397 9576 13103 9586
rect 43704 9586 43714 12479
rect 13237 9576 43714 9586
rect 12421 9552 13103 9562
rect 13213 9552 18191 9562
rect 18253 9552 38111 9562
rect 38149 9552 38159 9562
rect 12445 9528 16487 9538
rect 16525 9528 18191 9538
rect 43728 9538 43738 12480
rect 18229 9528 43738 9538
rect 12469 9504 38122 9514
rect 38112 9493 38122 9504
rect 12493 9480 16703 9490
rect 16741 9480 17447 9490
rect 17485 9480 19151 9490
rect 19189 9480 28727 9490
rect 12517 9456 16511 9466
rect 43752 9466 43762 12455
rect 16549 9456 43762 9466
rect 12541 9432 18407 9442
rect 18445 9432 19319 9442
rect 12565 9408 19175 9418
rect 12589 9384 17615 9394
rect 17640 9384 18023 9394
rect 17640 9370 17650 9384
rect 18048 9384 18239 9394
rect 12613 9360 17650 9370
rect 18048 9370 18058 9384
rect 18264 9384 18431 9394
rect 17677 9360 18058 9370
rect 18072 9360 18215 9370
rect 12637 9336 13703 9346
rect 18072 9346 18082 9360
rect 18264 9370 18274 9384
rect 18240 9360 18274 9370
rect 13728 9336 18082 9346
rect 12781 9312 13631 9322
rect 13728 9322 13738 9336
rect 18240 9346 18250 9360
rect 18205 9336 18250 9346
rect 13656 9312 13738 9322
rect 13752 9312 16535 9322
rect 12648 9274 12658 9311
rect 12781 9288 13487 9298
rect 13656 9298 13666 9312
rect 13752 9298 13762 9312
rect 16573 9312 17471 9322
rect 17496 9312 17663 9322
rect 13512 9288 13666 9298
rect 13680 9288 13762 9298
rect 12648 9264 13199 9274
rect 13512 9274 13522 9288
rect 13680 9274 13690 9288
rect 17496 9298 17506 9312
rect 14965 9288 17506 9298
rect 13261 9264 13522 9274
rect 13536 9264 13690 9274
rect 13536 9250 13546 9264
rect 15157 9264 16031 9274
rect 16069 9264 16727 9274
rect 12685 9240 13546 9250
rect 15949 9240 16007 9250
rect 16045 9240 16559 9250
rect 12709 9216 13175 9226
rect 13200 9216 13223 9226
rect 5904 9192 13151 9202
rect 13200 9202 13210 9216
rect 15973 9216 16055 9226
rect 13248 9202 13258 9215
rect 13176 9192 13210 9202
rect 13224 9192 13258 9202
rect 13176 9178 13186 9192
rect 13224 9178 13234 9192
rect 15997 9192 16031 9202
rect 12733 9168 13186 9178
rect 13200 9168 13234 9178
rect 12997 9144 13127 9154
rect 13200 9154 13210 9168
rect 13152 9144 13210 9154
rect 12744 9130 12754 9143
rect 13152 9130 13162 9144
rect 12744 9120 13162 9130
rect 12768 7474 12778 9095
rect 5828 7464 12778 7474
rect 5880 6562 5890 7439
rect 12792 6658 12802 9095
rect 12816 6685 12826 9095
rect 12840 6685 12850 9095
rect 12864 6685 12874 9095
rect 12888 6685 12898 9095
rect 12912 6685 12922 9095
rect 12936 6685 12946 9095
rect 12960 6685 12970 9095
rect 12984 6685 12994 9095
rect 13008 6685 13018 9095
rect 13032 6685 13042 9095
rect 13056 6682 13066 9095
rect 13080 6706 13090 9095
rect 13104 6730 13114 9095
rect 13104 6720 15850 6730
rect 13080 6696 15815 6706
rect 15840 6706 15850 6720
rect 15840 6696 15983 6706
rect 13056 6672 20303 6682
rect 12792 6648 16007 6658
rect 12792 6610 12802 6648
rect 16021 6648 20458 6658
rect 13021 6624 20423 6634
rect 20448 6634 20458 6648
rect 20448 6624 20471 6634
rect 20485 6624 29255 6634
rect 11557 6600 12802 6610
rect 12816 6610 12826 6623
rect 12816 6600 29375 6610
rect 38088 6589 38098 9431
rect 38112 7330 38122 9431
rect 38136 7474 38146 9431
rect 43776 7522 43786 12455
rect 43776 7512 43840 7522
rect 38136 7464 43840 7474
rect 38112 7320 43840 7330
rect 11509 6576 12839 6586
rect 12877 6576 29231 6586
rect 29269 6576 29423 6586
rect 29437 6576 33730 6586
rect 5880 6552 6911 6562
rect 11365 6552 12887 6562
rect 12925 6552 13007 6562
rect 13045 6552 15959 6562
rect 15997 6552 20279 6562
rect 20317 6552 33695 6562
rect 33720 6562 33730 6576
rect 33720 6552 33874 6562
rect 6888 6528 12935 6538
rect 6888 6514 6898 6528
rect 12973 6528 33839 6538
rect 33864 6538 33874 6552
rect 33888 6552 38207 6562
rect 33888 6541 33898 6552
rect 33864 6528 33887 6538
rect 38101 6528 38327 6538
rect 6864 6504 6898 6514
rect 6864 6450 6874 6504
rect 6925 6504 12983 6514
rect 6912 6450 6922 6503
rect 6960 6450 6970 6504
rect 13021 6504 38194 6514
rect 11352 6450 11362 6479
rect 11496 6450 11506 6479
rect 11544 6450 11554 6479
rect 15816 6450 15826 6479
rect 15960 6450 15970 6479
rect 16008 6450 16018 6479
rect 20280 6450 20290 6479
rect 20424 6450 20434 6479
rect 20472 6450 20482 6479
rect 29232 6450 29242 6479
rect 29376 6450 29386 6479
rect 29424 6450 29434 6479
rect 33696 6450 33706 6479
rect 33840 6450 33850 6479
rect 33888 6450 33898 6479
rect 38184 6450 38194 6504
rect 38221 6504 38386 6514
rect 38328 6450 38338 6479
rect 38376 6450 38386 6504
<< m2contact >>
rect 15743 44423 15757 44437
rect 15791 44423 15805 44437
rect 20231 44423 20245 44437
rect 20279 44423 20293 44437
rect 20423 44423 20437 44437
rect 29159 44423 29173 44437
rect 29207 44423 29221 44437
rect 33647 44423 33661 44437
rect 33695 44423 33709 44437
rect 33839 44423 33853 44437
rect 38111 44423 38125 44437
rect 29375 44399 29389 44413
rect 12959 44375 12973 44389
rect 29207 44375 29221 44389
rect 29231 44375 29245 44389
rect 33647 44375 33661 44389
rect 38111 44375 38125 44389
rect 12911 44351 12925 44365
rect 15791 44351 15805 44365
rect 15815 44351 15829 44365
rect 33839 44351 33853 44365
rect 12983 44327 12997 44341
rect 33695 44327 33709 44341
rect 38111 44327 38125 44341
rect 11327 44279 11341 44293
rect 12887 44279 12901 44293
rect 12935 44279 12949 44293
rect 13007 44279 13021 44293
rect 29375 44279 29389 44293
rect 11327 44231 11341 44245
rect 5903 43415 5917 43429
rect 6911 43415 6925 43429
rect 7007 43415 7021 43429
rect 11327 43415 11341 43429
rect 15743 44255 15757 44269
rect 15767 44255 15781 44269
rect 20231 44255 20245 44269
rect 29159 44255 29173 44269
rect 29231 44255 29245 44269
rect 12887 44231 12901 44245
rect 12911 44231 12925 44245
rect 12935 44231 12949 44245
rect 12959 44231 12973 44245
rect 12983 44231 12997 44245
rect 13007 44231 13021 44245
rect 5903 43367 5917 43381
rect 6911 43367 6925 43381
rect 7007 43367 7021 43381
rect 11327 43367 11341 43381
rect 5879 38303 5893 38317
rect 12887 40199 12901 40213
rect 12911 40199 12925 40213
rect 12935 40199 12949 40213
rect 12839 40175 12853 40189
rect 20423 44231 20437 44245
rect 20279 44207 20293 44221
rect 15815 44183 15829 44197
rect 12983 40175 12997 40189
rect 13007 40175 13021 40189
rect 13031 40175 13045 40189
rect 13055 40175 13069 40189
rect 13079 40175 13093 40189
rect 12815 40151 12829 40165
rect 12935 40151 12949 40165
rect 15767 44159 15781 44173
rect 38111 43607 38125 43621
rect 43775 43607 43789 43621
rect 13079 40127 13093 40141
rect 38111 43559 38125 43573
rect 43775 43559 43789 43573
rect 38111 43463 38125 43477
rect 43775 43463 43789 43477
rect 12791 40103 12805 40117
rect 12839 40103 12853 40117
rect 12767 40079 12781 40093
rect 13103 40103 13117 40117
rect 13127 40103 13141 40117
rect 38111 43415 38125 43429
rect 43775 43415 43789 43429
rect 12863 40079 12877 40093
rect 12887 40079 12901 40093
rect 7007 40055 7021 40069
rect 11327 40055 11341 40069
rect 12743 40055 12757 40069
rect 12935 40055 12949 40069
rect 12959 40055 12973 40069
rect 13055 40055 13069 40069
rect 13055 40031 13069 40045
rect 7007 40007 7021 40021
rect 11327 40007 11341 40021
rect 12695 40007 12709 40021
rect 12815 40007 12829 40021
rect 12839 40007 12853 40021
rect 13103 40055 13117 40069
rect 13127 40055 13141 40069
rect 12743 39983 12757 39997
rect 12815 39983 12829 39997
rect 13031 39959 13045 39973
rect 13055 39959 13069 39973
rect 13007 39935 13021 39949
rect 12719 39906 12733 39920
rect 12743 39906 12757 39920
rect 12983 39911 12997 39925
rect 12887 39888 12901 39902
rect 13223 39887 13237 39901
rect 13343 39887 13357 39901
rect 12983 39846 12997 39860
rect 40223 39846 40237 39860
rect 12983 39822 12997 39836
rect 12983 39798 12997 39812
rect 40223 39798 40237 39812
rect 40343 39798 40357 39812
rect 12695 39767 12709 39781
rect 12719 39767 12733 39781
rect 12743 39767 12757 39781
rect 12767 39767 12781 39781
rect 12791 39767 12805 39781
rect 12815 39767 12829 39781
rect 12839 39767 12853 39781
rect 12863 39767 12877 39781
rect 12887 39767 12901 39781
rect 12911 39767 12925 39781
rect 12935 39767 12949 39781
rect 12959 39767 12973 39781
rect 40223 39774 40237 39788
rect 5879 38255 5893 38269
rect 12695 35303 12709 35317
rect 12719 35303 12733 35317
rect 12743 35303 12757 35317
rect 12767 35303 12781 35317
rect 12791 35303 12805 35317
rect 12815 35303 12829 35317
rect 12839 35303 12853 35317
rect 12863 35303 12877 35317
rect 12887 35303 12901 35317
rect 12911 35303 12925 35317
rect 12671 35279 12685 35293
rect 40223 39750 40237 39764
rect 40223 39726 40237 39740
rect 40223 39702 40237 39716
rect 40223 39678 40237 39692
rect 40247 36503 40261 36517
rect 40343 39743 40357 39757
rect 43775 38447 43789 38461
rect 43775 38399 43789 38413
rect 43751 38327 43765 38341
rect 40295 36527 40309 36541
rect 40319 36527 40333 36541
rect 40343 36527 40357 36541
rect 40367 36527 40381 36541
rect 40391 36527 40405 36541
rect 40223 36479 40237 36493
rect 40247 36455 40261 36469
rect 12959 35279 12973 35293
rect 12983 35245 12997 35259
rect 12983 35221 12997 35235
rect 12671 35197 12685 35211
rect 12695 35197 12709 35211
rect 12719 35197 12733 35211
rect 12743 35197 12757 35211
rect 12767 35197 12781 35211
rect 12791 35197 12805 35211
rect 12935 35198 12949 35212
rect 12983 35197 12997 35211
rect 5879 33143 5893 33157
rect 5879 33095 5893 33109
rect 12695 31871 12709 31885
rect 12719 31871 12733 31885
rect 12671 31847 12685 31861
rect 12983 35173 12997 35187
rect 12815 35141 12829 35155
rect 12839 35141 12853 35155
rect 12863 35141 12877 35155
rect 12887 35141 12901 35155
rect 12911 35141 12925 35155
rect 12935 35141 12949 35155
rect 12959 35141 12973 35155
rect 12767 31847 12781 31861
rect 12791 31847 12805 31861
rect 12815 31847 12829 31861
rect 12839 31847 12853 31861
rect 12863 31847 12877 31861
rect 12647 31823 12661 31837
rect 40295 36479 40309 36493
rect 40319 36479 40333 36493
rect 40343 36479 40357 36493
rect 40367 36479 40381 36493
rect 40391 36479 40405 36493
rect 40247 33695 40261 33709
rect 40271 33695 40285 33709
rect 40319 33719 40333 33733
rect 40343 33719 40357 33733
rect 40367 33719 40381 33733
rect 40391 33719 40405 33733
rect 40415 33719 40429 33733
rect 40439 33695 40453 33709
rect 40223 33662 40237 33676
rect 40295 33662 40309 33676
rect 40343 33671 40357 33685
rect 40223 33638 40237 33652
rect 40367 33647 40381 33661
rect 40391 33647 40405 33661
rect 40415 33647 40429 33661
rect 40439 33647 40453 33661
rect 40247 33611 40261 33625
rect 40271 33611 40285 33625
rect 40295 33611 40309 33625
rect 40319 33611 40333 33625
rect 12911 31823 12925 31837
rect 12935 31823 12949 31837
rect 12959 31823 12973 31837
rect 12623 31799 12637 31813
rect 12863 31799 12877 31813
rect 12887 31799 12901 31813
rect 12983 31797 12997 31811
rect 12839 31775 12853 31789
rect 12863 31775 12877 31789
rect 12983 31773 12997 31787
rect 12623 31751 12637 31765
rect 12647 31751 12661 31765
rect 12671 31751 12685 31765
rect 12695 31751 12709 31765
rect 12719 31751 12733 31765
rect 12983 31749 12997 31763
rect 40247 31751 40261 31765
rect 40271 31751 40285 31765
rect 40319 31775 40333 31789
rect 40367 31799 40381 31813
rect 43751 38279 43765 38293
rect 43751 33335 43765 33349
rect 43775 33335 43789 33349
rect 43727 33287 43741 33301
rect 43727 33239 43741 33253
rect 43751 33239 43765 33253
rect 43775 33239 43789 33253
rect 43703 33143 43717 33157
rect 43727 33143 43741 33157
rect 43751 33143 43765 33157
rect 43775 33143 43789 33157
rect 40415 31823 40429 31837
rect 40439 31823 40453 31837
rect 40463 31823 40477 31837
rect 40487 31799 40501 31813
rect 40511 31775 40525 31789
rect 12767 31727 12781 31741
rect 12791 31727 12805 31741
rect 12815 31727 12829 31741
rect 12983 31725 12997 31739
rect 40223 31724 40237 31738
rect 40463 31727 40477 31741
rect 40535 31727 40549 31741
rect 12863 31703 12877 31717
rect 12887 31703 12901 31717
rect 12911 31703 12925 31717
rect 12935 31703 12949 31717
rect 12959 31703 12973 31717
rect 40223 31700 40237 31714
rect 40343 31703 40357 31717
rect 40391 31703 40405 31717
rect 40559 31703 40573 31717
rect 40223 31676 40237 31690
rect 40463 31679 40477 31693
rect 40487 31679 40501 31693
rect 40223 31652 40237 31666
rect 40487 31655 40501 31669
rect 40583 31655 40597 31669
rect 40223 31628 40237 31642
rect 40223 31604 40237 31618
rect 40295 31607 40309 31621
rect 40631 31607 40645 31621
rect 43703 33095 43717 33109
rect 43727 33095 43741 33109
rect 43751 33095 43765 33109
rect 43775 33095 43789 33109
rect 40247 31583 40261 31597
rect 40679 31583 40693 31597
rect 43679 31583 43693 31597
rect 12887 31559 12901 31573
rect 12911 31559 12925 31573
rect 12935 31559 12949 31573
rect 12959 31559 12973 31573
rect 24479 31559 24493 31573
rect 40247 31559 40261 31573
rect 12983 31535 12997 31549
rect 13007 31535 13021 31549
rect 27575 31535 27589 31549
rect 27599 31535 27613 31549
rect 40271 31535 40285 31549
rect 40319 31535 40333 31549
rect 40391 31535 40405 31549
rect 40415 31535 40429 31549
rect 40439 31535 40453 31549
rect 40463 31535 40477 31549
rect 40487 31535 40501 31549
rect 40511 31535 40525 31549
rect 40535 31535 40549 31549
rect 40559 31535 40573 31549
rect 40583 31535 40597 31549
rect 40631 31535 40645 31549
rect 40679 31535 40693 31549
rect 43679 31535 43693 31549
rect 12623 31511 12637 31525
rect 12647 31511 12661 31525
rect 12671 31511 12685 31525
rect 12695 31511 12709 31525
rect 12719 31511 12733 31525
rect 12743 31511 12757 31525
rect 12767 31511 12781 31525
rect 12791 31511 12805 31525
rect 12815 31511 12829 31525
rect 12839 31511 12853 31525
rect 12863 31511 12877 31525
rect 24479 31511 24493 31525
rect 24503 31511 24517 31525
rect 24527 31511 24541 31525
rect 12551 31487 12565 31501
rect 12575 31487 12589 31501
rect 12527 31463 12541 31477
rect 12719 31463 12733 31477
rect 12839 31463 12853 31477
rect 13055 31463 13069 31477
rect 13079 31463 13093 31477
rect 23423 31463 23437 31477
rect 23471 31463 23485 31477
rect 40367 31463 40381 31477
rect 12503 31439 12517 31453
rect 12671 31439 12685 31453
rect 12719 31439 12733 31453
rect 13369 31439 13383 31453
rect 13394 31439 13408 31453
rect 13463 31439 13477 31453
rect 13487 31439 13501 31453
rect 20471 31439 20485 31453
rect 20495 31439 20509 31453
rect 38159 31439 38173 31453
rect 12479 31415 12493 31429
rect 12743 31415 12757 31429
rect 12839 31415 12853 31429
rect 23423 31415 23437 31429
rect 23447 31415 23461 31429
rect 12455 31391 12469 31405
rect 12647 31391 12661 31405
rect 12671 31391 12685 31405
rect 21959 31391 21973 31405
rect 21983 31391 21997 31405
rect 12431 31367 12445 31381
rect 12767 31367 12781 31381
rect 12887 31367 12901 31381
rect 13103 31367 13117 31381
rect 13127 31367 13141 31381
rect 32246 31367 32260 31381
rect 32303 31367 32317 31381
rect 33743 31367 33757 31381
rect 35207 31367 35221 31381
rect 38111 31367 38125 31381
rect 40463 31367 40477 31381
rect 12551 31343 12565 31357
rect 12599 31343 12613 31357
rect 40463 31319 40477 31333
rect 40511 31319 40525 31333
rect 12407 31295 12421 31309
rect 12551 31295 12565 31309
rect 12647 31295 12661 31309
rect 12383 31271 12397 31285
rect 12815 31271 12829 31285
rect 12887 31271 12901 31285
rect 30791 31271 30805 31285
rect 30815 31271 30829 31285
rect 40511 31271 40525 31285
rect 12647 31247 12661 31261
rect 12743 31247 12757 31261
rect 24935 31247 24949 31261
rect 26423 31247 26437 31261
rect 26447 31247 26461 31261
rect 32270 31247 32284 31261
rect 37751 31247 37765 31261
rect 38087 31247 38101 31261
rect 12359 31223 12373 31237
rect 12503 31223 12517 31237
rect 12335 31199 12349 31213
rect 24935 31223 24949 31237
rect 24959 31223 24973 31237
rect 24983 31223 24997 31237
rect 12647 31199 12661 31213
rect 12695 31199 12709 31213
rect 12311 31175 12325 31189
rect 29327 31199 29341 31213
rect 29351 31199 29365 31213
rect 40631 31199 40645 31213
rect 40679 31199 40693 31213
rect 43679 31199 43693 31213
rect 43727 31199 43741 31213
rect 43751 31199 43765 31213
rect 12767 31175 12781 31189
rect 12815 31175 12829 31189
rect 13394 31175 13408 31189
rect 13463 31175 13477 31189
rect 13487 31175 13501 31189
rect 12263 31151 12277 31165
rect 12455 31151 12469 31165
rect 12503 31151 12517 31165
rect 12623 31127 12637 31141
rect 12695 31127 12709 31141
rect 13391 31127 13405 31141
rect 13415 31127 13429 31141
rect 13463 31127 13477 31141
rect 13487 31127 13501 31141
rect 13511 31127 13525 31141
rect 40631 31151 40645 31165
rect 43751 31151 43765 31165
rect 13607 31127 13621 31141
rect 12239 31079 12253 31093
rect 12287 31079 12301 31093
rect 12455 31079 12469 31093
rect 13511 31079 13525 31093
rect 13535 31079 13549 31093
rect 19007 31103 19021 31117
rect 19031 31103 19045 31117
rect 23471 31103 23485 31117
rect 23495 31103 23509 31117
rect 26447 31103 26461 31117
rect 13583 31079 13597 31093
rect 29327 31103 29341 31117
rect 29375 31103 29389 31117
rect 40679 31103 40693 31117
rect 43679 31103 43693 31117
rect 43727 31103 43741 31117
rect 27575 31079 27589 31093
rect 32303 31079 32317 31093
rect 12479 31055 12493 31069
rect 12623 31055 12637 31069
rect 13127 31055 13141 31069
rect 13175 31055 13189 31069
rect 12479 31031 12493 31045
rect 13607 31031 13621 31045
rect 15431 31031 15445 31045
rect 13127 31007 13141 31021
rect 12527 30983 12541 30997
rect 13031 30983 13045 30997
rect 13535 31007 13549 31021
rect 13175 30983 13189 30997
rect 13223 30983 13237 30997
rect 13368 30983 13382 30997
rect 13392 30983 13406 30997
rect 13487 30983 13501 30997
rect 13583 31007 13597 31021
rect 12215 30935 12229 30949
rect 12527 30935 12541 30949
rect 12215 30887 12229 30901
rect 12239 30887 12253 30901
rect 12263 30887 12277 30901
rect 12287 30887 12301 30901
rect 12311 30887 12325 30901
rect 12335 30887 12349 30901
rect 12359 30887 12373 30901
rect 12383 30887 12397 30901
rect 12407 30887 12421 30901
rect 12431 30887 12445 30901
rect 12455 30887 12469 30901
rect 12479 30887 12493 30901
rect 12503 30887 12517 30901
rect 12527 30887 12541 30901
rect 12551 30887 12565 30901
rect 12575 30887 12589 30901
rect 12599 30887 12613 30901
rect 12623 30887 12637 30901
rect 12647 30887 12661 30901
rect 12671 30887 12685 30901
rect 12695 30887 12709 30901
rect 12719 30887 12733 30901
rect 12743 30887 12757 30901
rect 12767 30887 12781 30901
rect 12791 30887 12805 30901
rect 12815 30887 12829 30901
rect 12839 30887 12853 30901
rect 12863 30887 12877 30901
rect 12887 30887 12901 30901
rect 12911 30887 12925 30901
rect 12935 30887 12949 30901
rect 12959 30887 12973 30901
rect 12983 30887 12997 30901
rect 13007 30887 13021 30901
rect 13031 30887 13045 30901
rect 13055 30887 13069 30901
rect 13079 30887 13093 30901
rect 13103 30887 13117 30901
rect 13127 30887 13141 30901
rect 12215 30623 12229 30637
rect 12239 30623 12253 30637
rect 12263 30623 12277 30637
rect 12287 30623 12301 30637
rect 12311 30623 12325 30637
rect 12335 30623 12349 30637
rect 12359 30623 12373 30637
rect 12383 30623 12397 30637
rect 12407 30623 12421 30637
rect 12191 30599 12205 30613
rect 12455 30599 12469 30613
rect 12479 30599 12493 30613
rect 12503 30599 12517 30613
rect 12527 30599 12541 30613
rect 12551 30599 12565 30613
rect 12575 30599 12589 30613
rect 12599 30599 12613 30613
rect 12623 30599 12637 30613
rect 12647 30599 12661 30613
rect 12671 30599 12685 30613
rect 12695 30599 12709 30613
rect 12719 30599 12733 30613
rect 12743 30599 12757 30613
rect 12767 30599 12781 30613
rect 12791 30599 12805 30613
rect 12815 30599 12829 30613
rect 12839 30599 12853 30613
rect 12863 30599 12877 30613
rect 12887 30599 12901 30613
rect 12167 30575 12181 30589
rect 12935 30575 12949 30589
rect 12959 30575 12973 30589
rect 12983 30575 12997 30589
rect 13007 30575 13021 30589
rect 13031 30575 13045 30589
rect 13055 30575 13069 30589
rect 12143 30551 12157 30565
rect 12599 30551 12613 30565
rect 12911 30551 12925 30565
rect 12959 30527 12973 30541
rect 12983 30527 12997 30541
rect 13079 30527 13093 30541
rect 13343 30959 13357 30973
rect 13415 30959 13429 30973
rect 13439 30935 13453 30949
rect 13463 30935 13477 30949
rect 13487 30695 13501 30709
rect 13598 30623 13612 30637
rect 13622 30623 13636 30637
rect 13463 30599 13477 30613
rect 13487 30599 13501 30613
rect 13646 30599 13660 30613
rect 13670 30599 13684 30613
rect 23447 31031 23461 31045
rect 23471 31031 23485 31045
rect 23495 31031 23509 31045
rect 24527 31031 24541 31045
rect 24983 31031 24997 31045
rect 17519 30983 17533 30997
rect 20495 30983 20509 30997
rect 19031 30959 19045 30973
rect 21983 30983 21997 30997
rect 24935 31007 24949 31021
rect 24959 31007 24973 31021
rect 24479 30983 24493 30997
rect 24503 30983 24517 30997
rect 23423 30959 23437 30973
rect 23471 30959 23485 30973
rect 27599 31031 27613 31045
rect 29375 31031 29389 31045
rect 29351 31007 29365 31021
rect 30815 31031 30829 31045
rect 38087 31031 38101 31045
rect 38111 31031 38125 31045
rect 38135 31031 38149 31045
rect 38159 31031 38173 31045
rect 39959 31031 39973 31045
rect 40247 31031 40261 31045
rect 40295 31031 40309 31045
rect 40343 31031 40357 31045
rect 29327 30983 29341 30997
rect 38111 30959 38125 30973
rect 38135 30959 38149 30973
rect 38159 30959 38173 30973
rect 38183 30935 38197 30949
rect 17159 30623 17173 30637
rect 17399 30623 17413 30637
rect 18359 30623 18373 30637
rect 18551 30623 18565 30637
rect 19583 30623 19597 30637
rect 27575 30623 27589 30637
rect 27839 30623 27853 30637
rect 28559 30623 28573 30637
rect 30359 30551 30373 30565
rect 30551 30527 30565 30541
rect 30671 30551 30685 30565
rect 38111 30887 38125 30901
rect 38135 30887 38149 30901
rect 38159 30887 38173 30901
rect 38183 30887 38197 30901
rect 30743 30527 30757 30541
rect 37919 30527 37933 30541
rect 38087 30527 38101 30541
rect 38111 30527 38125 30541
rect 38135 30527 38149 30541
rect 38159 30527 38173 30541
rect 38183 30527 38197 30541
rect 40247 30527 40261 30541
rect 40295 30527 40309 30541
rect 12119 30503 12133 30517
rect 12215 30503 12229 30517
rect 12431 30479 12445 30493
rect 12599 30479 12613 30493
rect 13031 30479 13045 30493
rect 13079 30479 13093 30493
rect 30623 30479 30637 30493
rect 30647 30479 30661 30493
rect 30719 30479 30733 30493
rect 30743 30479 30757 30493
rect 37919 30479 37933 30493
rect 38087 30479 38101 30493
rect 38207 30479 38221 30493
rect 40295 30479 40309 30493
rect 12095 30455 12109 30469
rect 12215 30455 12229 30469
rect 12551 30431 12565 30445
rect 12959 30431 12973 30445
rect 13007 30431 13021 30445
rect 13055 30431 13069 30445
rect 30647 30431 30661 30445
rect 30671 30431 30685 30445
rect 38087 30431 38101 30445
rect 40247 30431 40261 30445
rect 12095 30407 12109 30421
rect 12119 30407 12133 30421
rect 12143 30407 12157 30421
rect 12167 30407 12181 30421
rect 12191 30407 12205 30421
rect 12215 30407 12229 30421
rect 12239 30407 12253 30421
rect 12263 30407 12277 30421
rect 12287 30407 12301 30421
rect 12311 30407 12325 30421
rect 12335 30407 12349 30421
rect 12359 30407 12373 30421
rect 12383 30407 12397 30421
rect 12407 30407 12421 30421
rect 12431 30407 12445 30421
rect 12455 30407 12469 30421
rect 12479 30407 12493 30421
rect 12503 30407 12517 30421
rect 12527 30407 12541 30421
rect 12575 30383 12589 30397
rect 12599 30383 12613 30397
rect 12623 30383 12637 30397
rect 12647 30383 12661 30397
rect 12671 30383 12685 30397
rect 12695 30383 12709 30397
rect 12719 30383 12733 30397
rect 12743 30383 12757 30397
rect 12767 30383 12781 30397
rect 12791 30383 12805 30397
rect 12815 30383 12829 30397
rect 12839 30383 12853 30397
rect 12863 30383 12877 30397
rect 12887 30383 12901 30397
rect 12911 30383 12925 30397
rect 12935 30383 12949 30397
rect 12959 30383 12973 30397
rect 38087 30383 38101 30397
rect 38111 30383 38125 30397
rect 38135 30383 38149 30397
rect 38159 30383 38173 30397
rect 38183 30383 38197 30397
rect 38207 30383 38221 30397
rect 12095 27671 12109 27685
rect 12119 27671 12133 27685
rect 12143 27671 12157 27685
rect 12167 27671 12181 27685
rect 12191 27671 12205 27685
rect 12215 27671 12229 27685
rect 12239 27671 12253 27685
rect 12263 27671 12277 27685
rect 12287 27671 12301 27685
rect 12311 27671 12325 27685
rect 12335 27671 12349 27685
rect 12359 27671 12373 27685
rect 12383 27671 12397 27685
rect 12407 27671 12421 27685
rect 12431 27671 12445 27685
rect 12455 27671 12469 27685
rect 12479 27671 12493 27685
rect 12503 27671 12517 27685
rect 12527 27671 12541 27685
rect 12551 27671 12565 27685
rect 12575 27671 12589 27685
rect 12599 27671 12613 27685
rect 12623 27671 12637 27685
rect 12647 27671 12661 27685
rect 12671 27671 12685 27685
rect 12695 27671 12709 27685
rect 12719 27671 12733 27685
rect 12743 27671 12757 27685
rect 12767 27671 12781 27685
rect 12791 27671 12805 27685
rect 12815 27671 12829 27685
rect 12839 27671 12853 27685
rect 12863 27671 12877 27685
rect 12887 27671 12901 27685
rect 12911 27671 12925 27685
rect 12935 27671 12949 27685
rect 12959 27671 12973 27685
rect 12095 27623 12109 27637
rect 12119 27575 12133 27589
rect 12143 27551 12157 27565
rect 12167 27551 12181 27565
rect 12191 27551 12205 27565
rect 12215 27551 12229 27565
rect 12239 27551 12253 27565
rect 12263 27551 12277 27565
rect 12287 27551 12301 27565
rect 12311 27551 12325 27565
rect 12335 27551 12349 27565
rect 12359 27551 12373 27565
rect 12383 27551 12397 27565
rect 12407 27551 12421 27565
rect 12431 27551 12445 27565
rect 12455 27551 12469 27565
rect 12479 27551 12493 27565
rect 12503 27551 12517 27565
rect 12527 27551 12541 27565
rect 12551 27551 12565 27565
rect 12575 27551 12589 27565
rect 12599 27551 12613 27565
rect 12623 27551 12637 27565
rect 12647 27551 12661 27565
rect 12671 27551 12685 27565
rect 12695 27551 12709 27565
rect 12719 27551 12733 27565
rect 12743 27551 12757 27565
rect 12767 27551 12781 27565
rect 12791 27551 12805 27565
rect 12815 27551 12829 27565
rect 12839 27551 12853 27565
rect 12863 27551 12877 27565
rect 12887 27551 12901 27565
rect 12911 27551 12925 27565
rect 12935 27551 12949 27565
rect 12959 27551 12973 27565
rect 12167 26495 12181 26509
rect 12191 26495 12205 26509
rect 12215 26495 12229 26509
rect 12239 26495 12253 26509
rect 12263 26495 12277 26509
rect 12287 26495 12301 26509
rect 12311 26495 12325 26509
rect 12335 26495 12349 26509
rect 12359 26495 12373 26509
rect 12383 26495 12397 26509
rect 12407 26495 12421 26509
rect 12431 26495 12445 26509
rect 12455 26495 12469 26509
rect 12479 26495 12493 26509
rect 12503 26495 12517 26509
rect 12527 26495 12541 26509
rect 12551 26495 12565 26509
rect 12575 26495 12589 26509
rect 12599 26495 12613 26509
rect 12623 26495 12637 26509
rect 12647 26495 12661 26509
rect 12671 26495 12685 26509
rect 12695 26495 12709 26509
rect 12719 26495 12733 26509
rect 12743 26495 12757 26509
rect 12767 26495 12781 26509
rect 12791 26495 12805 26509
rect 12815 26495 12829 26509
rect 12839 26495 12853 26509
rect 12863 26495 12877 26509
rect 12887 26495 12901 26509
rect 12911 26495 12925 26509
rect 12935 26495 12949 26509
rect 12959 26495 12973 26509
rect 12167 26447 12181 26461
rect 12191 26399 12205 26413
rect 12215 26375 12229 26389
rect 12239 26375 12253 26389
rect 12263 26375 12277 26389
rect 12287 26375 12301 26389
rect 12311 26375 12325 26389
rect 12335 26375 12349 26389
rect 12359 26375 12373 26389
rect 12383 26375 12397 26389
rect 12407 26375 12421 26389
rect 12431 26375 12445 26389
rect 12455 26375 12469 26389
rect 12479 26375 12493 26389
rect 12503 26375 12517 26389
rect 12527 26375 12541 26389
rect 12551 26375 12565 26389
rect 12575 26375 12589 26389
rect 12599 26375 12613 26389
rect 12623 26375 12637 26389
rect 12647 26375 12661 26389
rect 12671 26375 12685 26389
rect 12695 26375 12709 26389
rect 12719 26375 12733 26389
rect 12743 26375 12757 26389
rect 12767 26375 12781 26389
rect 12791 26375 12805 26389
rect 12815 26375 12829 26389
rect 12839 26375 12853 26389
rect 12863 26375 12877 26389
rect 12887 26375 12901 26389
rect 12911 26375 12925 26389
rect 12935 26375 12949 26389
rect 12959 26375 12973 26389
rect 12239 25319 12253 25333
rect 12263 25319 12277 25333
rect 12287 25319 12301 25333
rect 12311 25319 12325 25333
rect 12335 25319 12349 25333
rect 12359 25319 12373 25333
rect 12383 25319 12397 25333
rect 12407 25319 12421 25333
rect 12431 25319 12445 25333
rect 12455 25319 12469 25333
rect 12479 25319 12493 25333
rect 12503 25319 12517 25333
rect 12527 25319 12541 25333
rect 12551 25319 12565 25333
rect 12575 25319 12589 25333
rect 12599 25319 12613 25333
rect 12623 25319 12637 25333
rect 12647 25319 12661 25333
rect 12671 25319 12685 25333
rect 12695 25319 12709 25333
rect 12719 25319 12733 25333
rect 12743 25319 12757 25333
rect 12767 25319 12781 25333
rect 12791 25319 12805 25333
rect 12815 25319 12829 25333
rect 12839 25319 12853 25333
rect 12863 25319 12877 25333
rect 12887 25319 12901 25333
rect 12911 25319 12925 25333
rect 12935 25319 12949 25333
rect 12959 25319 12973 25333
rect 12239 25271 12253 25285
rect 12263 25223 12277 25237
rect 12287 25199 12301 25213
rect 12311 25199 12325 25213
rect 12335 25199 12349 25213
rect 12359 25199 12373 25213
rect 12383 25199 12397 25213
rect 12407 25199 12421 25213
rect 12431 25199 12445 25213
rect 12455 25199 12469 25213
rect 12479 25199 12493 25213
rect 12503 25199 12517 25213
rect 12527 25199 12541 25213
rect 12551 25199 12565 25213
rect 12575 25199 12589 25213
rect 12599 25199 12613 25213
rect 12623 25199 12637 25213
rect 12647 25199 12661 25213
rect 12671 25199 12685 25213
rect 12695 25199 12709 25213
rect 12719 25199 12733 25213
rect 12743 25199 12757 25213
rect 12767 25199 12781 25213
rect 12791 25199 12805 25213
rect 12815 25199 12829 25213
rect 12839 25199 12853 25213
rect 12863 25199 12877 25213
rect 12887 25199 12901 25213
rect 12911 25199 12925 25213
rect 12935 25199 12949 25213
rect 12959 25199 12973 25213
rect 12311 24143 12325 24157
rect 12335 24143 12349 24157
rect 12359 24143 12373 24157
rect 12383 24143 12397 24157
rect 12407 24143 12421 24157
rect 12431 24143 12445 24157
rect 12455 24143 12469 24157
rect 12479 24143 12493 24157
rect 12503 24143 12517 24157
rect 12527 24143 12541 24157
rect 12551 24143 12565 24157
rect 12575 24143 12589 24157
rect 12599 24143 12613 24157
rect 12623 24143 12637 24157
rect 12647 24143 12661 24157
rect 12671 24143 12685 24157
rect 12695 24143 12709 24157
rect 12719 24143 12733 24157
rect 12743 24143 12757 24157
rect 12767 24143 12781 24157
rect 12791 24143 12805 24157
rect 12815 24143 12829 24157
rect 12839 24143 12853 24157
rect 12863 24143 12877 24157
rect 12887 24143 12901 24157
rect 12911 24143 12925 24157
rect 12935 24143 12949 24157
rect 12959 24143 12973 24157
rect 12311 24095 12325 24109
rect 12335 24047 12349 24061
rect 12359 24023 12373 24037
rect 12383 24023 12397 24037
rect 12407 24023 12421 24037
rect 12431 24023 12445 24037
rect 12455 24023 12469 24037
rect 12479 24023 12493 24037
rect 12503 24023 12517 24037
rect 12527 24023 12541 24037
rect 12551 24023 12565 24037
rect 12575 24023 12589 24037
rect 12599 24023 12613 24037
rect 12623 24023 12637 24037
rect 12647 24023 12661 24037
rect 12671 24023 12685 24037
rect 12695 24023 12709 24037
rect 12719 24023 12733 24037
rect 12743 24023 12757 24037
rect 12767 24023 12781 24037
rect 12791 24023 12805 24037
rect 12815 24023 12829 24037
rect 12839 24023 12853 24037
rect 12863 24023 12877 24037
rect 12887 24023 12901 24037
rect 12911 24023 12925 24037
rect 12935 24023 12949 24037
rect 12959 24023 12973 24037
rect 5879 22967 5893 22981
rect 12383 22967 12397 22981
rect 12407 22967 12421 22981
rect 12431 22967 12445 22981
rect 12455 22967 12469 22981
rect 12479 22967 12493 22981
rect 12503 22967 12517 22981
rect 12527 22967 12541 22981
rect 12551 22967 12565 22981
rect 12575 22967 12589 22981
rect 12599 22967 12613 22981
rect 12623 22967 12637 22981
rect 12647 22967 12661 22981
rect 12671 22967 12685 22981
rect 12695 22967 12709 22981
rect 12719 22967 12733 22981
rect 12743 22967 12757 22981
rect 12767 22967 12781 22981
rect 12791 22967 12805 22981
rect 12815 22967 12829 22981
rect 12839 22967 12853 22981
rect 12863 22967 12877 22981
rect 12887 22967 12901 22981
rect 12911 22967 12925 22981
rect 12935 22967 12949 22981
rect 12959 22967 12973 22981
rect 5879 22919 5893 22933
rect 12383 22919 12397 22933
rect 12407 22871 12421 22885
rect 12431 22847 12445 22861
rect 12455 22847 12469 22861
rect 12479 22847 12493 22861
rect 12503 22847 12517 22861
rect 12527 22847 12541 22861
rect 12551 22847 12565 22861
rect 12575 22847 12589 22861
rect 12599 22847 12613 22861
rect 12623 22847 12637 22861
rect 12647 22847 12661 22861
rect 12671 22847 12685 22861
rect 12695 22847 12709 22861
rect 12719 22847 12733 22861
rect 12743 22847 12757 22861
rect 12767 22847 12781 22861
rect 12791 22847 12805 22861
rect 12815 22847 12829 22861
rect 12839 22847 12853 22861
rect 12863 22847 12877 22861
rect 12887 22847 12901 22861
rect 12911 22847 12925 22861
rect 12935 22847 12949 22861
rect 12959 22847 12973 22861
rect 12455 21791 12469 21805
rect 12479 21791 12493 21805
rect 12503 21791 12517 21805
rect 12527 21791 12541 21805
rect 12551 21791 12565 21805
rect 12575 21791 12589 21805
rect 12599 21791 12613 21805
rect 12623 21791 12637 21805
rect 12647 21791 12661 21805
rect 12671 21791 12685 21805
rect 12695 21791 12709 21805
rect 12719 21791 12733 21805
rect 12743 21791 12757 21805
rect 12767 21791 12781 21805
rect 12791 21791 12805 21805
rect 12815 21791 12829 21805
rect 12839 21791 12853 21805
rect 12863 21791 12877 21805
rect 12887 21791 12901 21805
rect 12911 21791 12925 21805
rect 12935 21791 12949 21805
rect 12959 21791 12973 21805
rect 12455 21743 12469 21757
rect 12479 21695 12493 21709
rect 12503 21671 12517 21685
rect 12527 21671 12541 21685
rect 12551 21671 12565 21685
rect 12575 21671 12589 21685
rect 12599 21671 12613 21685
rect 12623 21671 12637 21685
rect 12647 21671 12661 21685
rect 12671 21671 12685 21685
rect 12695 21671 12709 21685
rect 12719 21671 12733 21685
rect 12743 21671 12757 21685
rect 12767 21671 12781 21685
rect 12791 21671 12805 21685
rect 12815 21671 12829 21685
rect 12839 21671 12853 21685
rect 12863 21671 12877 21685
rect 12887 21671 12901 21685
rect 12911 21671 12925 21685
rect 12935 21671 12949 21685
rect 12959 21671 12973 21685
rect 12527 20615 12541 20629
rect 12551 20615 12565 20629
rect 12575 20615 12589 20629
rect 12599 20615 12613 20629
rect 12623 20615 12637 20629
rect 12647 20615 12661 20629
rect 12671 20615 12685 20629
rect 12695 20615 12709 20629
rect 12719 20615 12733 20629
rect 12743 20615 12757 20629
rect 12767 20615 12781 20629
rect 12791 20615 12805 20629
rect 12815 20615 12829 20629
rect 12839 20615 12853 20629
rect 12863 20615 12877 20629
rect 12887 20615 12901 20629
rect 12911 20615 12925 20629
rect 12935 20615 12949 20629
rect 12959 20615 12973 20629
rect 12527 20567 12541 20581
rect 12551 20519 12565 20533
rect 12575 20495 12589 20509
rect 12599 20495 12613 20509
rect 12623 20495 12637 20509
rect 12647 20495 12661 20509
rect 12671 20495 12685 20509
rect 12695 20495 12709 20509
rect 12719 20495 12733 20509
rect 12743 20495 12757 20509
rect 12767 20495 12781 20509
rect 12791 20495 12805 20509
rect 12815 20495 12829 20509
rect 12839 20495 12853 20509
rect 12863 20495 12877 20509
rect 12887 20495 12901 20509
rect 12911 20495 12925 20509
rect 12935 20495 12949 20509
rect 12959 20495 12973 20509
rect 12599 19439 12613 19453
rect 12623 19439 12637 19453
rect 12647 19439 12661 19453
rect 12671 19439 12685 19453
rect 12695 19439 12709 19453
rect 12719 19439 12733 19453
rect 12743 19439 12757 19453
rect 12767 19439 12781 19453
rect 12791 19439 12805 19453
rect 12815 19439 12829 19453
rect 12839 19439 12853 19453
rect 12863 19439 12877 19453
rect 12887 19439 12901 19453
rect 12911 19439 12925 19453
rect 12935 19439 12949 19453
rect 12959 19439 12973 19453
rect 12575 19391 12589 19405
rect 12887 19391 12901 19405
rect 12671 19367 12685 19381
rect 12887 19367 12901 19381
rect 12575 19343 12589 19357
rect 12599 19343 12613 19357
rect 12623 19343 12637 19357
rect 12647 19343 12661 19357
rect 12695 19319 12709 19333
rect 12719 19319 12733 19333
rect 12743 19319 12757 19333
rect 12767 19319 12781 19333
rect 12791 19319 12805 19333
rect 12815 19319 12829 19333
rect 12839 19319 12853 19333
rect 12863 19319 12877 19333
rect 12887 19319 12901 19333
rect 12911 19319 12925 19333
rect 12935 19319 12949 19333
rect 12959 19319 12973 19333
rect 12551 18239 12565 18253
rect 12575 18239 12589 18253
rect 12599 18239 12613 18253
rect 12623 18239 12637 18253
rect 12647 18239 12661 18253
rect 12671 18239 12685 18253
rect 12695 18239 12709 18253
rect 12719 18239 12733 18253
rect 12527 18215 12541 18229
rect 12767 18215 12781 18229
rect 12791 18215 12805 18229
rect 12815 18215 12829 18229
rect 12839 18215 12853 18229
rect 12863 18215 12877 18229
rect 12887 18215 12901 18229
rect 12911 18215 12925 18229
rect 12935 18215 12949 18229
rect 12959 18215 12973 18229
rect 5879 17807 5893 17821
rect 5903 17807 5917 17821
rect 12719 18191 12733 18205
rect 12743 18191 12757 18205
rect 12527 18167 12541 18181
rect 12551 18167 12565 18181
rect 12575 18167 12589 18181
rect 12599 18167 12613 18181
rect 12623 18167 12637 18181
rect 12647 18167 12661 18181
rect 12671 18167 12685 18181
rect 12695 18167 12709 18181
rect 5879 17759 5893 17773
rect 5903 17759 5917 17773
rect 12743 18143 12757 18157
rect 12767 18143 12781 18157
rect 12791 18143 12805 18157
rect 12815 18143 12829 18157
rect 12839 18143 12853 18157
rect 12863 18143 12877 18157
rect 12887 18143 12901 18157
rect 12911 18143 12925 18157
rect 12935 18143 12949 18157
rect 12959 18143 12973 18157
rect 12527 17063 12541 17077
rect 12551 17063 12565 17077
rect 12575 17063 12589 17077
rect 12599 17063 12613 17077
rect 12623 17063 12637 17077
rect 12647 17063 12661 17077
rect 12671 17063 12685 17077
rect 12695 17063 12709 17077
rect 12719 17063 12733 17077
rect 12743 17063 12757 17077
rect 12767 17063 12781 17077
rect 12791 17063 12805 17077
rect 12815 17063 12829 17077
rect 12839 17063 12853 17077
rect 12863 17063 12877 17077
rect 12887 17063 12901 17077
rect 12503 17039 12517 17053
rect 12935 17039 12949 17053
rect 12959 17039 12973 17053
rect 12839 17015 12853 17029
rect 12911 17015 12925 17029
rect 12503 16991 12517 17005
rect 12527 16991 12541 17005
rect 12551 16991 12565 17005
rect 12575 16991 12589 17005
rect 12599 16991 12613 17005
rect 12623 16991 12637 17005
rect 12647 16991 12661 17005
rect 12671 16991 12685 17005
rect 12695 16991 12709 17005
rect 12719 16991 12733 17005
rect 12743 16991 12757 17005
rect 12767 16991 12781 17005
rect 12791 16991 12805 17005
rect 12815 16991 12829 17005
rect 12863 16967 12877 16981
rect 12887 16967 12901 16981
rect 12911 16967 12925 16981
rect 12935 16967 12949 16981
rect 12959 16967 12973 16981
rect 12479 15887 12493 15901
rect 12503 15887 12517 15901
rect 12527 15887 12541 15901
rect 12551 15887 12565 15901
rect 12575 15887 12589 15901
rect 12599 15887 12613 15901
rect 12623 15887 12637 15901
rect 12647 15887 12661 15901
rect 12671 15887 12685 15901
rect 12695 15887 12709 15901
rect 12719 15887 12733 15901
rect 12743 15887 12757 15901
rect 12767 15887 12781 15901
rect 12791 15887 12805 15901
rect 12815 15887 12829 15901
rect 12839 15887 12853 15901
rect 12863 15887 12877 15901
rect 12887 15887 12901 15901
rect 12455 15863 12469 15877
rect 12935 15863 12949 15877
rect 12959 15863 12973 15877
rect 12863 15839 12877 15853
rect 12911 15839 12925 15853
rect 12455 15815 12469 15829
rect 12479 15815 12493 15829
rect 12503 15815 12517 15829
rect 12527 15815 12541 15829
rect 12551 15815 12565 15829
rect 12575 15815 12589 15829
rect 12599 15815 12613 15829
rect 12623 15815 12637 15829
rect 12647 15815 12661 15829
rect 12671 15815 12685 15829
rect 12695 15815 12709 15829
rect 12719 15815 12733 15829
rect 12743 15815 12757 15829
rect 12767 15815 12781 15829
rect 12791 15815 12805 15829
rect 12815 15815 12829 15829
rect 12839 15815 12853 15829
rect 12887 15791 12901 15805
rect 12911 15791 12925 15805
rect 12935 15791 12949 15805
rect 12959 15791 12973 15805
rect 12431 14735 12445 14749
rect 12455 14735 12469 14749
rect 12479 14735 12493 14749
rect 12503 14735 12517 14749
rect 12527 14735 12541 14749
rect 12551 14735 12565 14749
rect 12575 14735 12589 14749
rect 12599 14735 12613 14749
rect 12623 14735 12637 14749
rect 12647 14735 12661 14749
rect 12671 14735 12685 14749
rect 12695 14735 12709 14749
rect 12719 14735 12733 14749
rect 12743 14735 12757 14749
rect 12767 14735 12781 14749
rect 12791 14735 12805 14749
rect 12815 14735 12829 14749
rect 12839 14735 12853 14749
rect 12863 14735 12877 14749
rect 12407 14711 12421 14725
rect 12911 14711 12925 14725
rect 12935 14711 12949 14725
rect 12407 14663 12421 14677
rect 12431 14663 12445 14677
rect 12455 14663 12469 14677
rect 12479 14663 12493 14677
rect 12503 14663 12517 14677
rect 12527 14663 12541 14677
rect 12551 14663 12565 14677
rect 12575 14663 12589 14677
rect 12599 14663 12613 14677
rect 12623 14663 12637 14677
rect 12647 14663 12661 14677
rect 12671 14663 12685 14677
rect 12695 14663 12709 14677
rect 12719 14663 12733 14677
rect 12743 14663 12757 14677
rect 12767 14663 12781 14677
rect 12791 14663 12805 14677
rect 12815 14663 12829 14677
rect 12839 14663 12853 14677
rect 12863 14663 12877 14677
rect 12383 13535 12397 13549
rect 12407 13535 12421 13549
rect 12431 13535 12445 13549
rect 12455 13535 12469 13549
rect 12479 13535 12493 13549
rect 12503 13535 12517 13549
rect 12527 13535 12541 13549
rect 12551 13535 12565 13549
rect 12575 13535 12589 13549
rect 12599 13535 12613 13549
rect 12623 13535 12637 13549
rect 12647 13535 12661 13549
rect 12671 13535 12685 13549
rect 12695 13535 12709 13549
rect 12719 13535 12733 13549
rect 12743 13535 12757 13549
rect 12767 13535 12781 13549
rect 12791 13535 12805 13549
rect 12815 13535 12829 13549
rect 12839 13535 12853 13549
rect 12359 13511 12373 13525
rect 12911 14639 12925 14653
rect 12935 14639 12949 14653
rect 12887 13511 12901 13525
rect 12911 13511 12925 13525
rect 12935 13511 12949 13525
rect 12959 13511 12973 13525
rect 5879 12647 5893 12661
rect 5903 12647 5917 12661
rect 12815 13487 12829 13501
rect 12863 13487 12877 13501
rect 12359 13463 12373 13477
rect 12383 13463 12397 13477
rect 12407 13463 12421 13477
rect 12431 13463 12445 13477
rect 12455 13463 12469 13477
rect 12479 13463 12493 13477
rect 12503 13463 12517 13477
rect 12527 13463 12541 13477
rect 12551 13463 12565 13477
rect 12575 13463 12589 13477
rect 12599 13463 12613 13477
rect 12623 13463 12637 13477
rect 12647 13463 12661 13477
rect 12671 13463 12685 13477
rect 12695 13463 12709 13477
rect 12719 13463 12733 13477
rect 12743 13463 12757 13477
rect 12767 13463 12781 13477
rect 12791 13463 12805 13477
rect 5879 12599 5893 12613
rect 5903 12599 5917 12613
rect 12359 12383 12373 12397
rect 12383 12383 12397 12397
rect 12335 12359 12349 12373
rect 12839 13439 12853 13453
rect 12863 13439 12877 13453
rect 12887 13439 12901 13453
rect 12911 13439 12925 13453
rect 12935 13439 12949 13453
rect 12959 13439 12973 13453
rect 12431 12359 12445 12373
rect 12455 12359 12469 12373
rect 12479 12359 12493 12373
rect 12503 12359 12517 12373
rect 12527 12359 12541 12373
rect 12551 12359 12565 12373
rect 12575 12359 12589 12373
rect 12599 12359 12613 12373
rect 12623 12359 12637 12373
rect 12647 12359 12661 12373
rect 12671 12359 12685 12373
rect 12695 12359 12709 12373
rect 12719 12359 12733 12373
rect 12743 12359 12757 12373
rect 12767 12359 12781 12373
rect 12791 12359 12805 12373
rect 12815 12359 12829 12373
rect 12839 12359 12853 12373
rect 12863 12359 12877 12373
rect 12911 12335 12925 12349
rect 12935 12335 12949 12349
rect 12959 12335 12973 12349
rect 12335 12311 12349 12325
rect 12359 12311 12373 12325
rect 12383 12311 12397 12325
rect 12311 11183 12325 11197
rect 12431 12287 12445 12301
rect 12455 12287 12469 12301
rect 12479 12287 12493 12301
rect 12503 12287 12517 12301
rect 12527 12287 12541 12301
rect 12551 12287 12565 12301
rect 12575 12287 12589 12301
rect 12599 12287 12613 12301
rect 12623 12287 12637 12301
rect 12647 12287 12661 12301
rect 12671 12287 12685 12301
rect 12695 12287 12709 12301
rect 12719 12287 12733 12301
rect 12743 12287 12757 12301
rect 12767 12287 12781 12301
rect 12791 12287 12805 12301
rect 12815 12287 12829 12301
rect 12839 12287 12853 12301
rect 12863 12287 12877 12301
rect 12911 12263 12925 12277
rect 12935 12263 12949 12277
rect 12959 12263 12973 12277
rect 12359 11159 12373 11173
rect 12383 11159 12397 11173
rect 12407 11159 12421 11173
rect 12431 11159 12445 11173
rect 12455 11159 12469 11173
rect 12479 11159 12493 11173
rect 12503 11159 12517 11173
rect 12527 11159 12541 11173
rect 12551 11159 12565 11173
rect 12575 11159 12589 11173
rect 12599 11159 12613 11173
rect 12623 11159 12637 11173
rect 12647 11159 12661 11173
rect 12671 11159 12685 11173
rect 12695 11159 12709 11173
rect 12719 11159 12733 11173
rect 12743 11159 12757 11173
rect 12767 11159 12781 11173
rect 12791 11159 12805 11173
rect 12815 11159 12829 11173
rect 12839 11159 12853 11173
rect 12863 11159 12877 11173
rect 12887 11159 12901 11173
rect 12911 11159 12925 11173
rect 12935 11159 12949 11173
rect 12959 11159 12973 11173
rect 12335 11135 12349 11149
rect 12311 11087 12325 11101
rect 12335 11087 12349 11101
rect 12359 11087 12373 11101
rect 12383 11087 12397 11101
rect 12407 11087 12421 11101
rect 12431 11087 12445 11101
rect 12455 11087 12469 11101
rect 12479 11087 12493 11101
rect 12503 11087 12517 11101
rect 12527 11087 12541 11101
rect 12551 11087 12565 11101
rect 12575 11087 12589 11101
rect 12599 11087 12613 11101
rect 12623 11087 12637 11101
rect 12647 11087 12661 11101
rect 12671 11087 12685 11101
rect 12695 11087 12709 11101
rect 12719 11087 12733 11101
rect 12743 11087 12757 11101
rect 12767 11087 12781 11101
rect 12791 11087 12805 11101
rect 12815 11087 12829 11101
rect 12839 11087 12853 11101
rect 12863 11087 12877 11101
rect 12887 11087 12901 11101
rect 12911 11087 12925 11101
rect 12935 11087 12949 11101
rect 12959 11087 12973 11101
rect 12263 10007 12277 10021
rect 12287 10007 12301 10021
rect 12311 10007 12325 10021
rect 12335 10007 12349 10021
rect 12359 10007 12373 10021
rect 12383 10007 12397 10021
rect 12407 10007 12421 10021
rect 12431 10007 12445 10021
rect 12455 10007 12469 10021
rect 12479 10007 12493 10021
rect 12503 10007 12517 10021
rect 12527 10007 12541 10021
rect 12551 10007 12565 10021
rect 12575 10007 12589 10021
rect 12599 10007 12613 10021
rect 12623 10007 12637 10021
rect 12647 10007 12661 10021
rect 12671 10007 12685 10021
rect 12695 10007 12709 10021
rect 12719 10007 12733 10021
rect 12743 10007 12757 10021
rect 12767 10007 12781 10021
rect 12791 10007 12805 10021
rect 12815 10007 12829 10021
rect 12839 10007 12853 10021
rect 12863 10007 12877 10021
rect 12239 9983 12253 9997
rect 12911 9983 12925 9997
rect 12935 9983 12949 9997
rect 12959 9983 12973 9997
rect 12839 9959 12853 9973
rect 12887 9959 12901 9973
rect 12239 9935 12253 9949
rect 12263 9935 12277 9949
rect 12287 9935 12301 9949
rect 12311 9935 12325 9949
rect 12335 9935 12349 9949
rect 12359 9935 12373 9949
rect 12383 9935 12397 9949
rect 12407 9935 12421 9949
rect 12431 9935 12445 9949
rect 12455 9935 12469 9949
rect 12479 9935 12493 9949
rect 12503 9935 12517 9949
rect 12527 9935 12541 9949
rect 12551 9935 12565 9949
rect 12575 9935 12589 9949
rect 12599 9935 12613 9949
rect 12623 9935 12637 9949
rect 12647 9935 12661 9949
rect 12671 9935 12685 9949
rect 12695 9935 12709 9949
rect 12719 9935 12733 9949
rect 12743 9935 12757 9949
rect 12767 9935 12781 9949
rect 12791 9935 12805 9949
rect 12815 9935 12829 9949
rect 12863 9911 12877 9925
rect 12887 9911 12901 9925
rect 12911 9911 12925 9925
rect 12935 9911 12949 9925
rect 12959 9911 12973 9925
rect 12239 9767 12253 9781
rect 12263 9767 12277 9781
rect 12287 9767 12301 9781
rect 12311 9767 12325 9781
rect 12335 9767 12349 9781
rect 12359 9767 12373 9781
rect 12383 9767 12397 9781
rect 12407 9767 12421 9781
rect 12431 9767 12445 9781
rect 12455 9767 12469 9781
rect 12479 9767 12493 9781
rect 12503 9767 12517 9781
rect 12527 9767 12541 9781
rect 12551 9767 12565 9781
rect 12575 9767 12589 9781
rect 12599 9767 12613 9781
rect 12623 9767 12637 9781
rect 12647 9767 12661 9781
rect 12671 9767 12685 9781
rect 12695 9767 12709 9781
rect 12719 9767 12733 9781
rect 12743 9767 12757 9781
rect 12767 9767 12781 9781
rect 12791 9767 12805 9781
rect 12815 9767 12829 9781
rect 12839 9767 12853 9781
rect 12863 9767 12877 9781
rect 12887 9767 12901 9781
rect 12911 9767 12925 9781
rect 12935 9767 12949 9781
rect 12959 9767 12973 9781
rect 38087 9767 38101 9781
rect 43727 28055 43741 28069
rect 43799 28031 43813 28045
rect 43727 28007 43741 28021
rect 43775 17807 43789 17821
rect 43775 17759 43789 17773
rect 43751 17663 43765 17677
rect 43775 17663 43789 17677
rect 43751 17615 43765 17629
rect 43775 17615 43789 17629
rect 43727 12647 43741 12661
rect 43751 12647 43765 12661
rect 43775 12647 43789 12661
rect 43727 12599 43741 12613
rect 43751 12599 43765 12613
rect 43775 12599 43789 12613
rect 43703 12527 43717 12541
rect 38135 9791 38149 9805
rect 38159 9791 38173 9805
rect 38183 9791 38197 9805
rect 38111 9743 38125 9757
rect 12239 9719 12253 9733
rect 13007 9719 13021 9733
rect 13103 9719 13117 9733
rect 15983 9719 15997 9733
rect 16007 9719 16021 9733
rect 12263 9695 12277 9709
rect 43751 12503 43765 12517
rect 43775 12503 43789 12517
rect 43703 12479 43717 12493
rect 12287 9671 12301 9685
rect 13031 9671 13045 9685
rect 13103 9671 13117 9685
rect 12311 9647 12325 9661
rect 13055 9647 13069 9661
rect 13463 9671 13477 9685
rect 13487 9671 13501 9685
rect 13679 9671 13693 9685
rect 13703 9671 13717 9685
rect 15959 9671 15973 9685
rect 16031 9671 16045 9685
rect 38183 9671 38197 9685
rect 13607 9647 13621 9661
rect 13631 9647 13645 9661
rect 17999 9647 18013 9661
rect 18023 9647 18037 9661
rect 29159 9647 29173 9661
rect 36863 9647 36877 9661
rect 38159 9647 38173 9661
rect 12335 9623 12349 9637
rect 13079 9623 13093 9637
rect 13103 9623 13117 9637
rect 13127 9623 13141 9637
rect 13151 9623 13165 9637
rect 13175 9623 13189 9637
rect 28919 9623 28933 9637
rect 37607 9623 37621 9637
rect 38087 9623 38101 9637
rect 38111 9623 38125 9637
rect 12359 9599 12373 9613
rect 38087 9599 38101 9613
rect 38111 9599 38125 9613
rect 38135 9599 38149 9613
rect 38159 9599 38173 9613
rect 12383 9575 12397 9589
rect 13103 9575 13117 9589
rect 13223 9575 13237 9589
rect 12407 9551 12421 9565
rect 13103 9551 13117 9565
rect 13199 9551 13213 9565
rect 18191 9551 18205 9565
rect 18239 9551 18253 9565
rect 38111 9551 38125 9565
rect 38135 9551 38149 9565
rect 38159 9551 38173 9565
rect 12431 9527 12445 9541
rect 16487 9527 16501 9541
rect 16511 9527 16525 9541
rect 18191 9527 18205 9541
rect 18215 9527 18229 9541
rect 43751 12455 43765 12469
rect 43775 12455 43789 12469
rect 12455 9503 12469 9517
rect 12479 9479 12493 9493
rect 16703 9479 16717 9493
rect 16727 9479 16741 9493
rect 17447 9479 17461 9493
rect 17471 9479 17485 9493
rect 19151 9479 19165 9493
rect 19175 9479 19189 9493
rect 28727 9479 28741 9493
rect 38111 9479 38125 9493
rect 12503 9455 12517 9469
rect 16511 9455 16525 9469
rect 16535 9455 16549 9469
rect 12527 9431 12541 9445
rect 18407 9431 18421 9445
rect 18431 9431 18445 9445
rect 19319 9431 19333 9445
rect 38087 9431 38101 9445
rect 38111 9431 38125 9445
rect 38135 9431 38149 9445
rect 12551 9407 12565 9421
rect 19175 9407 19189 9421
rect 12575 9383 12589 9397
rect 17615 9383 17629 9397
rect 12599 9359 12613 9373
rect 18023 9383 18037 9397
rect 17663 9359 17677 9373
rect 18239 9383 18253 9397
rect 12623 9335 12637 9349
rect 13703 9335 13717 9349
rect 18215 9359 18229 9373
rect 18431 9383 18445 9397
rect 12647 9311 12661 9325
rect 12767 9311 12781 9325
rect 13631 9311 13645 9325
rect 18191 9335 18205 9349
rect 12767 9287 12781 9301
rect 13487 9287 13501 9301
rect 16535 9311 16549 9325
rect 16559 9311 16573 9325
rect 17471 9311 17485 9325
rect 13199 9263 13213 9277
rect 13247 9263 13261 9277
rect 14951 9287 14965 9301
rect 17663 9311 17677 9325
rect 12671 9239 12685 9253
rect 15143 9263 15157 9277
rect 16031 9263 16045 9277
rect 16055 9263 16069 9277
rect 16727 9263 16741 9277
rect 15935 9239 15949 9253
rect 16007 9239 16021 9253
rect 16031 9239 16045 9253
rect 16559 9239 16573 9253
rect 12695 9215 12709 9229
rect 13175 9215 13189 9229
rect 13151 9191 13165 9205
rect 13223 9215 13237 9229
rect 13247 9215 13261 9229
rect 15959 9215 15973 9229
rect 16055 9215 16069 9229
rect 12719 9167 12733 9181
rect 15983 9191 15997 9205
rect 16031 9191 16045 9205
rect 12743 9143 12757 9157
rect 12983 9143 12997 9157
rect 13127 9143 13141 9157
rect 12767 9095 12781 9109
rect 12791 9095 12805 9109
rect 12815 9095 12829 9109
rect 12839 9095 12853 9109
rect 12863 9095 12877 9109
rect 12887 9095 12901 9109
rect 12911 9095 12925 9109
rect 12935 9095 12949 9109
rect 12959 9095 12973 9109
rect 12983 9095 12997 9109
rect 13007 9095 13021 9109
rect 13031 9095 13045 9109
rect 13055 9095 13069 9109
rect 13079 9095 13093 9109
rect 13103 9095 13117 9109
rect 5879 7487 5893 7501
rect 5879 7439 5893 7453
rect 12815 6671 12829 6685
rect 12839 6671 12853 6685
rect 12863 6671 12877 6685
rect 12887 6671 12901 6685
rect 12911 6671 12925 6685
rect 12935 6671 12949 6685
rect 12959 6671 12973 6685
rect 12983 6671 12997 6685
rect 13007 6671 13021 6685
rect 13031 6671 13045 6685
rect 15815 6695 15829 6709
rect 15983 6695 15997 6709
rect 20303 6671 20317 6685
rect 11543 6599 11557 6613
rect 16007 6647 16021 6661
rect 12815 6623 12829 6637
rect 13007 6623 13021 6637
rect 20423 6623 20437 6637
rect 20471 6623 20485 6637
rect 29255 6623 29269 6637
rect 29375 6599 29389 6613
rect 11495 6575 11509 6589
rect 12839 6575 12853 6589
rect 12863 6575 12877 6589
rect 29231 6575 29245 6589
rect 29255 6575 29269 6589
rect 29423 6575 29437 6589
rect 6911 6551 6925 6565
rect 11351 6551 11365 6565
rect 12887 6551 12901 6565
rect 12911 6551 12925 6565
rect 13007 6551 13021 6565
rect 13031 6551 13045 6565
rect 15959 6551 15973 6565
rect 15983 6551 15997 6565
rect 20279 6551 20293 6565
rect 20303 6551 20317 6565
rect 33695 6551 33709 6565
rect 38087 6575 38101 6589
rect 12935 6527 12949 6541
rect 12959 6527 12973 6541
rect 33839 6527 33853 6541
rect 38207 6551 38221 6565
rect 33887 6527 33901 6541
rect 38087 6527 38101 6541
rect 38327 6527 38341 6541
rect 6911 6503 6925 6517
rect 12983 6503 12997 6517
rect 13007 6503 13021 6517
rect 11351 6479 11365 6493
rect 11495 6479 11509 6493
rect 11543 6479 11557 6493
rect 15815 6479 15829 6493
rect 15959 6479 15973 6493
rect 16007 6479 16021 6493
rect 20279 6479 20293 6493
rect 20423 6479 20437 6493
rect 20471 6479 20485 6493
rect 29231 6479 29245 6493
rect 29375 6479 29389 6493
rect 29423 6479 29437 6493
rect 33695 6479 33709 6493
rect 33839 6479 33853 6493
rect 33887 6479 33901 6493
rect 38207 6503 38221 6517
rect 38327 6479 38341 6493
<< metal2 >>
rect 11328 44245 11340 44279
rect 12888 44245 12900 44279
rect 12912 44245 12924 44351
rect 12936 44245 12948 44279
rect 12960 44245 12972 44375
rect 12984 44245 12996 44327
rect 13008 44245 13020 44279
rect 15744 44269 15756 44423
rect 15792 44365 15804 44423
rect 15768 44173 15780 44255
rect 15816 44197 15828 44351
rect 20232 44269 20244 44423
rect 20280 44221 20292 44423
rect 20424 44245 20436 44423
rect 29160 44269 29172 44423
rect 29208 44389 29220 44423
rect 29232 44269 29244 44375
rect 29376 44293 29388 44399
rect 33648 44389 33660 44423
rect 33696 44341 33708 44423
rect 33840 44365 33852 44423
rect 38112 44389 38124 44423
rect 38112 44341 38124 44375
rect 38112 43573 38124 43607
rect 43776 43573 43788 43607
rect 38112 43429 38124 43463
rect 43776 43429 43788 43463
rect 5904 43381 5916 43415
rect 6912 43381 6924 43415
rect 7008 43381 7020 43415
rect 11328 43381 11340 43415
rect 7008 40021 7020 40055
rect 11328 40021 11340 40055
rect 12696 39781 12708 40007
rect 12744 39997 12756 40055
rect 12720 39781 12732 39906
rect 12744 39781 12756 39906
rect 12768 39781 12780 40079
rect 12792 39781 12804 40103
rect 12816 40021 12828 40151
rect 12840 40117 12852 40175
rect 12888 40093 12900 40199
rect 12816 39781 12828 39983
rect 12840 39781 12852 40007
rect 12864 39781 12876 40079
rect 12888 39781 12900 39888
rect 12912 39781 12924 40199
rect 12936 40165 12948 40199
rect 12936 39781 12948 40055
rect 12960 39781 12972 40055
rect 12984 39925 12996 40175
rect 13008 39949 13020 40175
rect 13032 39973 13044 40175
rect 13056 40069 13068 40175
rect 13080 40141 13092 40175
rect 13104 40069 13116 40103
rect 13128 40069 13140 40103
rect 13056 39973 13068 40031
rect 13357 39887 13359 39901
rect 13224 39870 13236 39887
rect 13347 39870 13359 39887
rect 12997 39847 13008 39859
rect 40191 39847 40223 39859
rect 12997 39823 13008 39835
rect 12997 39799 13008 39811
rect 40191 39799 40223 39811
rect 40191 39775 40223 39787
rect 40191 39751 40223 39763
rect 40344 39757 40356 39798
rect 40191 39727 40223 39739
rect 40191 39703 40223 39715
rect 40191 39679 40223 39691
rect 43776 38413 43788 38447
rect 5880 38269 5892 38303
rect 43752 38293 43764 38327
rect 40191 36479 40223 36482
rect 40191 36470 40237 36479
rect 40248 36469 40260 36503
rect 40296 36493 40308 36527
rect 40320 36493 40332 36527
rect 40344 36493 40356 36527
rect 40368 36493 40380 36527
rect 40392 36493 40404 36527
rect 12672 35211 12684 35279
rect 12696 35211 12708 35303
rect 12720 35211 12732 35303
rect 12744 35211 12756 35303
rect 12768 35211 12780 35303
rect 12792 35211 12804 35303
rect 12816 35155 12828 35303
rect 12840 35155 12852 35303
rect 12864 35155 12876 35303
rect 12888 35155 12900 35303
rect 12912 35155 12924 35303
rect 12936 35155 12948 35198
rect 12960 35155 12972 35279
rect 12997 35246 13008 35258
rect 12997 35222 13008 35234
rect 12997 35198 13008 35210
rect 12997 35174 13008 35186
rect 40191 33662 40223 33674
rect 40191 33638 40223 33650
rect 40248 33625 40260 33695
rect 40272 33625 40284 33695
rect 40296 33625 40308 33662
rect 40320 33625 40332 33719
rect 40344 33685 40356 33719
rect 40368 33661 40380 33719
rect 40392 33661 40404 33719
rect 40416 33661 40428 33719
rect 40440 33661 40452 33695
rect 43728 33253 43740 33287
rect 43752 33253 43764 33335
rect 43776 33253 43788 33335
rect 5880 33109 5892 33143
rect 43704 33109 43716 33143
rect 43728 33109 43740 33143
rect 43752 33109 43764 33143
rect 43776 33109 43788 33143
rect 12624 31765 12636 31799
rect 12648 31765 12660 31823
rect 12672 31765 12684 31847
rect 12696 31765 12708 31871
rect 12720 31765 12732 31871
rect 12768 31741 12780 31847
rect 12792 31741 12804 31847
rect 12816 31741 12828 31847
rect 12840 31789 12852 31847
rect 12864 31813 12876 31847
rect 12864 31717 12876 31775
rect 12888 31717 12900 31799
rect 12912 31717 12924 31823
rect 12936 31717 12948 31823
rect 12960 31717 12972 31823
rect 12997 31797 13008 31809
rect 12997 31773 13008 31785
rect 12997 31749 13008 31761
rect 12997 31725 13008 31737
rect 40191 31725 40223 31737
rect 40191 31701 40223 31713
rect 40191 31677 40223 31689
rect 40191 31653 40223 31665
rect 40191 31629 40223 31641
rect 40191 31605 40223 31617
rect 40248 31597 40260 31751
rect 12216 30901 12228 30935
rect 12240 30901 12252 31079
rect 12264 30901 12276 31151
rect 12288 30901 12300 31079
rect 12312 30901 12324 31175
rect 12336 30901 12348 31199
rect 12360 30901 12372 31223
rect 12384 30901 12396 31271
rect 12408 30901 12420 31295
rect 12432 30901 12444 31367
rect 12456 31165 12468 31391
rect 12456 30901 12468 31079
rect 12480 31069 12492 31415
rect 12504 31237 12516 31439
rect 12480 30901 12492 31031
rect 12504 30901 12516 31151
rect 12528 30997 12540 31463
rect 12552 31357 12564 31487
rect 12528 30901 12540 30935
rect 12552 30901 12564 31295
rect 12576 30901 12588 31487
rect 12600 30901 12612 31343
rect 12624 31141 12636 31511
rect 12648 31405 12660 31511
rect 12672 31453 12684 31511
rect 12648 31261 12660 31295
rect 12624 30901 12636 31055
rect 12648 30901 12660 31199
rect 12672 30901 12684 31391
rect 12696 31213 12708 31511
rect 12720 31477 12732 31511
rect 12696 30901 12708 31127
rect 12720 30901 12732 31439
rect 12744 31429 12756 31511
rect 12768 31381 12780 31511
rect 12744 30901 12756 31247
rect 12768 30901 12780 31175
rect 12792 30901 12804 31511
rect 12816 31285 12828 31511
rect 12840 31477 12852 31511
rect 12816 30901 12828 31175
rect 12840 30901 12852 31415
rect 12864 30901 12876 31511
rect 12888 31381 12900 31559
rect 12888 30901 12900 31271
rect 12912 30901 12924 31559
rect 12936 30901 12948 31559
rect 12960 30901 12972 31559
rect 12984 30901 12996 31535
rect 13008 30901 13020 31535
rect 13032 30901 13044 30983
rect 13056 30901 13068 31463
rect 13080 30901 13092 31463
rect 13104 30901 13116 31367
rect 13128 31069 13140 31367
rect 13128 30901 13140 31007
rect 13176 30997 13188 31055
rect 13224 30997 13236 31594
rect 13347 31586 13359 31594
rect 13346 31574 13359 31586
rect 13346 30985 13358 31574
rect 13371 31453 13383 31594
rect 13395 31453 13407 31594
rect 13369 30997 13381 31439
rect 13395 31189 13407 31439
rect 13419 31188 13431 31594
rect 15423 31572 15435 31594
rect 17523 31572 17535 31594
rect 15423 31560 15444 31572
rect 13464 31189 13476 31439
rect 13488 31189 13500 31439
rect 13419 31176 13452 31188
rect 13393 30997 13405 31127
rect 13343 30973 13358 30985
rect 13416 30973 13428 31127
rect 13440 30949 13452 31176
rect 13464 30949 13476 31127
rect 13488 30997 13500 31127
rect 13512 31093 13524 31127
rect 13536 31021 13548 31079
rect 13584 31021 13596 31079
rect 13608 31045 13620 31127
rect 15432 31045 15444 31560
rect 17520 31560 17535 31572
rect 18999 31572 19011 31594
rect 20475 31572 20487 31594
rect 18999 31560 19020 31572
rect 17520 30997 17532 31560
rect 19008 31117 19020 31560
rect 20472 31560 20487 31572
rect 21951 31572 21963 31594
rect 23427 31572 23439 31594
rect 21951 31560 21972 31572
rect 20472 31453 20484 31560
rect 19032 30973 19044 31103
rect 20496 30997 20508 31439
rect 21960 31405 21972 31560
rect 23424 31560 23439 31572
rect 24471 31573 24483 31594
rect 23424 31477 23436 31560
rect 24471 31559 24479 31573
rect 24939 31572 24951 31594
rect 24936 31560 24951 31572
rect 26415 31572 26427 31594
rect 29319 31572 29331 31594
rect 30783 31572 30795 31594
rect 26415 31560 26436 31572
rect 29319 31560 29340 31572
rect 30783 31560 30804 31572
rect 21984 30997 21996 31391
rect 23424 30973 23436 31415
rect 23448 31045 23460 31415
rect 23472 31117 23484 31463
rect 23496 31045 23508 31103
rect 23472 30973 23484 31031
rect 24480 30997 24492 31511
rect 24504 30997 24516 31511
rect 24528 31045 24540 31511
rect 24936 31261 24948 31560
rect 26424 31261 26436 31560
rect 24936 31021 24948 31223
rect 24960 31021 24972 31223
rect 24984 31045 24996 31223
rect 26448 31117 26460 31247
rect 27576 31093 27588 31535
rect 27600 31045 27612 31535
rect 29328 31213 29340 31560
rect 30792 31285 30804 31560
rect 32247 31381 32259 31594
rect 29328 30997 29340 31103
rect 29352 31021 29364 31199
rect 29376 31045 29388 31103
rect 30816 31045 30828 31271
rect 32271 31261 32283 31594
rect 33735 31572 33747 31594
rect 35199 31572 35211 31594
rect 37743 31572 37755 31594
rect 38127 31572 38139 31594
rect 33735 31560 33756 31572
rect 35199 31560 35220 31572
rect 37743 31560 37764 31572
rect 38127 31560 38148 31572
rect 33744 31381 33756 31560
rect 35208 31381 35220 31560
rect 32304 31093 32316 31367
rect 37752 31261 37764 31560
rect 38088 31045 38100 31247
rect 38112 31045 38124 31367
rect 38136 31045 38148 31560
rect 38160 31045 38172 31439
rect 39960 31045 39972 31594
rect 40248 31045 40260 31559
rect 40272 31549 40284 31751
rect 40296 31045 40308 31607
rect 40320 31549 40332 31775
rect 40344 31045 40356 31703
rect 40368 31477 40380 31799
rect 40392 31549 40404 31703
rect 40416 31549 40428 31823
rect 40440 31549 40452 31823
rect 40464 31741 40476 31823
rect 40488 31693 40500 31799
rect 40464 31549 40476 31679
rect 40488 31549 40500 31655
rect 40512 31549 40524 31775
rect 40536 31549 40548 31727
rect 40560 31549 40572 31703
rect 40584 31549 40596 31655
rect 40632 31549 40644 31607
rect 40680 31549 40692 31583
rect 43680 31549 43692 31583
rect 40464 31333 40476 31367
rect 40512 31285 40524 31319
rect 40632 31165 40644 31199
rect 40680 31117 40692 31199
rect 43680 31117 43692 31199
rect 43728 31117 43740 31199
rect 43752 31165 43764 31199
rect 38112 30901 38124 30959
rect 38136 30901 38148 30959
rect 38160 30901 38172 30959
rect 38184 30901 38196 30935
rect 12096 30421 12108 30455
rect 12120 30421 12132 30503
rect 12144 30421 12156 30551
rect 12168 30421 12180 30575
rect 12192 30421 12204 30599
rect 12216 30517 12228 30623
rect 12216 30421 12228 30455
rect 12240 30421 12252 30623
rect 12264 30421 12276 30623
rect 12288 30421 12300 30623
rect 12312 30421 12324 30623
rect 12336 30421 12348 30623
rect 12360 30421 12372 30623
rect 12384 30421 12396 30623
rect 12408 30421 12420 30623
rect 13488 30613 13500 30695
rect 12432 30421 12444 30479
rect 12456 30421 12468 30599
rect 12480 30421 12492 30599
rect 12504 30421 12516 30599
rect 12528 30421 12540 30599
rect 12552 30445 12564 30599
rect 12576 30397 12588 30599
rect 12600 30565 12612 30599
rect 12600 30397 12612 30479
rect 12624 30397 12636 30599
rect 12648 30397 12660 30599
rect 12672 30397 12684 30599
rect 12696 30397 12708 30599
rect 12720 30397 12732 30599
rect 12744 30397 12756 30599
rect 12768 30397 12780 30599
rect 12792 30397 12804 30599
rect 12816 30397 12828 30599
rect 12840 30397 12852 30599
rect 12864 30397 12876 30599
rect 12888 30397 12900 30599
rect 12912 30397 12924 30551
rect 12936 30397 12948 30575
rect 12960 30541 12972 30575
rect 12984 30541 12996 30575
rect 13008 30445 13020 30575
rect 13032 30493 13044 30575
rect 13056 30445 13068 30575
rect 13080 30493 13092 30527
rect 12960 30397 12972 30431
rect 13464 30364 13476 30599
rect 13599 30364 13611 30623
rect 13623 30364 13635 30623
rect 13647 30364 13659 30599
rect 13671 30364 13683 30599
rect 17160 30396 17172 30623
rect 17400 30396 17412 30623
rect 18360 30396 18372 30623
rect 18552 30396 18564 30623
rect 19584 30396 19596 30623
rect 27576 30396 27588 30623
rect 27840 30396 27852 30623
rect 28560 30396 28572 30623
rect 30360 30396 30372 30551
rect 30552 30396 30564 30527
rect 30624 30396 30636 30479
rect 30648 30445 30660 30479
rect 30672 30445 30684 30551
rect 30744 30493 30756 30527
rect 37920 30493 37932 30527
rect 38088 30493 38100 30527
rect 30720 30396 30732 30479
rect 17151 30384 17172 30396
rect 17391 30384 17412 30396
rect 18351 30384 18372 30396
rect 18543 30384 18564 30396
rect 19577 30384 19596 30396
rect 27568 30384 27588 30396
rect 27832 30384 27852 30396
rect 28552 30384 28572 30396
rect 30351 30384 30372 30396
rect 30543 30384 30564 30396
rect 30615 30384 30636 30396
rect 30711 30384 30732 30396
rect 17151 30364 17163 30384
rect 17391 30364 17403 30384
rect 18351 30364 18363 30384
rect 18543 30364 18555 30384
rect 19577 30364 19589 30384
rect 27568 30364 27580 30384
rect 27832 30364 27844 30384
rect 28552 30364 28564 30384
rect 30351 30364 30363 30384
rect 30543 30364 30555 30384
rect 30615 30364 30627 30384
rect 30711 30364 30723 30384
rect 37920 30364 37932 30479
rect 38088 30397 38100 30431
rect 38112 30397 38124 30527
rect 38136 30397 38148 30527
rect 38160 30397 38172 30527
rect 38184 30397 38196 30527
rect 38208 30397 38220 30479
rect 40248 30445 40260 30527
rect 40296 30493 40308 30527
rect 43728 28021 43740 28055
rect 43813 28032 43840 28044
rect 12096 27637 12108 27671
rect 12120 27589 12132 27671
rect 12144 27565 12156 27671
rect 12168 27565 12180 27671
rect 12192 27565 12204 27671
rect 12216 27565 12228 27671
rect 12240 27565 12252 27671
rect 12264 27565 12276 27671
rect 12288 27565 12300 27671
rect 12312 27565 12324 27671
rect 12336 27565 12348 27671
rect 12360 27565 12372 27671
rect 12384 27565 12396 27671
rect 12408 27565 12420 27671
rect 12432 27565 12444 27671
rect 12456 27565 12468 27671
rect 12480 27565 12492 27671
rect 12504 27565 12516 27671
rect 12528 27565 12540 27671
rect 12552 27565 12564 27671
rect 12576 27565 12588 27671
rect 12600 27565 12612 27671
rect 12624 27565 12636 27671
rect 12648 27565 12660 27671
rect 12672 27565 12684 27671
rect 12696 27565 12708 27671
rect 12720 27565 12732 27671
rect 12744 27565 12756 27671
rect 12768 27565 12780 27671
rect 12792 27565 12804 27671
rect 12816 27565 12828 27671
rect 12840 27565 12852 27671
rect 12864 27565 12876 27671
rect 12888 27565 12900 27671
rect 12912 27565 12924 27671
rect 12936 27565 12948 27671
rect 12960 27565 12972 27671
rect 12168 26461 12180 26495
rect 12192 26413 12204 26495
rect 12216 26389 12228 26495
rect 12240 26389 12252 26495
rect 12264 26389 12276 26495
rect 12288 26389 12300 26495
rect 12312 26389 12324 26495
rect 12336 26389 12348 26495
rect 12360 26389 12372 26495
rect 12384 26389 12396 26495
rect 12408 26389 12420 26495
rect 12432 26389 12444 26495
rect 12456 26389 12468 26495
rect 12480 26389 12492 26495
rect 12504 26389 12516 26495
rect 12528 26389 12540 26495
rect 12552 26389 12564 26495
rect 12576 26389 12588 26495
rect 12600 26389 12612 26495
rect 12624 26389 12636 26495
rect 12648 26389 12660 26495
rect 12672 26389 12684 26495
rect 12696 26389 12708 26495
rect 12720 26389 12732 26495
rect 12744 26389 12756 26495
rect 12768 26389 12780 26495
rect 12792 26389 12804 26495
rect 12816 26389 12828 26495
rect 12840 26389 12852 26495
rect 12864 26389 12876 26495
rect 12888 26389 12900 26495
rect 12912 26389 12924 26495
rect 12936 26389 12948 26495
rect 12960 26389 12972 26495
rect 12240 25285 12252 25319
rect 12264 25237 12276 25319
rect 12288 25213 12300 25319
rect 12312 25213 12324 25319
rect 12336 25213 12348 25319
rect 12360 25213 12372 25319
rect 12384 25213 12396 25319
rect 12408 25213 12420 25319
rect 12432 25213 12444 25319
rect 12456 25213 12468 25319
rect 12480 25213 12492 25319
rect 12504 25213 12516 25319
rect 12528 25213 12540 25319
rect 12552 25213 12564 25319
rect 12576 25213 12588 25319
rect 12600 25213 12612 25319
rect 12624 25213 12636 25319
rect 12648 25213 12660 25319
rect 12672 25213 12684 25319
rect 12696 25213 12708 25319
rect 12720 25213 12732 25319
rect 12744 25213 12756 25319
rect 12768 25213 12780 25319
rect 12792 25213 12804 25319
rect 12816 25213 12828 25319
rect 12840 25213 12852 25319
rect 12864 25213 12876 25319
rect 12888 25213 12900 25319
rect 12912 25213 12924 25319
rect 12936 25213 12948 25319
rect 12960 25213 12972 25319
rect 12312 24109 12324 24143
rect 12336 24061 12348 24143
rect 12360 24037 12372 24143
rect 12384 24037 12396 24143
rect 12408 24037 12420 24143
rect 12432 24037 12444 24143
rect 12456 24037 12468 24143
rect 12480 24037 12492 24143
rect 12504 24037 12516 24143
rect 12528 24037 12540 24143
rect 12552 24037 12564 24143
rect 12576 24037 12588 24143
rect 12600 24037 12612 24143
rect 12624 24037 12636 24143
rect 12648 24037 12660 24143
rect 12672 24037 12684 24143
rect 12696 24037 12708 24143
rect 12720 24037 12732 24143
rect 12744 24037 12756 24143
rect 12768 24037 12780 24143
rect 12792 24037 12804 24143
rect 12816 24037 12828 24143
rect 12840 24037 12852 24143
rect 12864 24037 12876 24143
rect 12888 24037 12900 24143
rect 12912 24037 12924 24143
rect 12936 24037 12948 24143
rect 12960 24037 12972 24143
rect 5880 22933 5892 22967
rect 12384 22933 12396 22967
rect 12408 22885 12420 22967
rect 12432 22861 12444 22967
rect 12456 22861 12468 22967
rect 12480 22861 12492 22967
rect 12504 22861 12516 22967
rect 12528 22861 12540 22967
rect 12552 22861 12564 22967
rect 12576 22861 12588 22967
rect 12600 22861 12612 22967
rect 12624 22861 12636 22967
rect 12648 22861 12660 22967
rect 12672 22861 12684 22967
rect 12696 22861 12708 22967
rect 12720 22861 12732 22967
rect 12744 22861 12756 22967
rect 12768 22861 12780 22967
rect 12792 22861 12804 22967
rect 12816 22861 12828 22967
rect 12840 22861 12852 22967
rect 12864 22861 12876 22967
rect 12888 22861 12900 22967
rect 12912 22861 12924 22967
rect 12936 22861 12948 22967
rect 12960 22861 12972 22967
rect 12456 21757 12468 21791
rect 12480 21709 12492 21791
rect 12504 21685 12516 21791
rect 12528 21685 12540 21791
rect 12552 21685 12564 21791
rect 12576 21685 12588 21791
rect 12600 21685 12612 21791
rect 12624 21685 12636 21791
rect 12648 21685 12660 21791
rect 12672 21685 12684 21791
rect 12696 21685 12708 21791
rect 12720 21685 12732 21791
rect 12744 21685 12756 21791
rect 12768 21685 12780 21791
rect 12792 21685 12804 21791
rect 12816 21685 12828 21791
rect 12840 21685 12852 21791
rect 12864 21685 12876 21791
rect 12888 21685 12900 21791
rect 12912 21685 12924 21791
rect 12936 21685 12948 21791
rect 12960 21685 12972 21791
rect 12528 20581 12540 20615
rect 12552 20533 12564 20615
rect 12576 20509 12588 20615
rect 12600 20509 12612 20615
rect 12624 20509 12636 20615
rect 12648 20509 12660 20615
rect 12672 20509 12684 20615
rect 12696 20509 12708 20615
rect 12720 20509 12732 20615
rect 12744 20509 12756 20615
rect 12768 20509 12780 20615
rect 12792 20509 12804 20615
rect 12816 20509 12828 20615
rect 12840 20509 12852 20615
rect 12864 20509 12876 20615
rect 12888 20509 12900 20615
rect 12912 20509 12924 20615
rect 12936 20509 12948 20615
rect 12960 20509 12972 20615
rect 12576 19357 12588 19391
rect 12600 19357 12612 19439
rect 12624 19357 12636 19439
rect 12648 19357 12660 19439
rect 12672 19381 12684 19439
rect 12696 19333 12708 19439
rect 12720 19333 12732 19439
rect 12744 19333 12756 19439
rect 12768 19333 12780 19439
rect 12792 19333 12804 19439
rect 12816 19333 12828 19439
rect 12840 19333 12852 19439
rect 12864 19333 12876 19439
rect 12888 19405 12900 19439
rect 12888 19333 12900 19367
rect 12912 19333 12924 19439
rect 12936 19333 12948 19439
rect 12960 19333 12972 19439
rect 12528 18181 12540 18215
rect 12552 18181 12564 18239
rect 12576 18181 12588 18239
rect 12600 18181 12612 18239
rect 12624 18181 12636 18239
rect 12648 18181 12660 18239
rect 12672 18181 12684 18239
rect 12696 18181 12708 18239
rect 12720 18205 12732 18239
rect 12744 18157 12756 18191
rect 12768 18157 12780 18215
rect 12792 18157 12804 18215
rect 12816 18157 12828 18215
rect 12840 18157 12852 18215
rect 12864 18157 12876 18215
rect 12888 18157 12900 18215
rect 12912 18157 12924 18215
rect 12936 18157 12948 18215
rect 12960 18157 12972 18215
rect 5880 17773 5892 17807
rect 5904 17773 5916 17807
rect 43776 17773 43788 17807
rect 43752 17629 43764 17663
rect 43776 17629 43788 17663
rect 12504 17005 12516 17039
rect 12528 17005 12540 17063
rect 12552 17005 12564 17063
rect 12576 17005 12588 17063
rect 12600 17005 12612 17063
rect 12624 17005 12636 17063
rect 12648 17005 12660 17063
rect 12672 17005 12684 17063
rect 12696 17005 12708 17063
rect 12720 17005 12732 17063
rect 12744 17005 12756 17063
rect 12768 17005 12780 17063
rect 12792 17005 12804 17063
rect 12816 17005 12828 17063
rect 12840 17029 12852 17063
rect 12864 16981 12876 17063
rect 12888 16981 12900 17063
rect 12912 16981 12924 17015
rect 12936 16981 12948 17039
rect 12960 16981 12972 17039
rect 12456 15829 12468 15863
rect 12480 15829 12492 15887
rect 12504 15829 12516 15887
rect 12528 15829 12540 15887
rect 12552 15829 12564 15887
rect 12576 15829 12588 15887
rect 12600 15829 12612 15887
rect 12624 15829 12636 15887
rect 12648 15829 12660 15887
rect 12672 15829 12684 15887
rect 12696 15829 12708 15887
rect 12720 15829 12732 15887
rect 12744 15829 12756 15887
rect 12768 15829 12780 15887
rect 12792 15829 12804 15887
rect 12816 15829 12828 15887
rect 12840 15829 12852 15887
rect 12864 15853 12876 15887
rect 12888 15805 12900 15887
rect 12912 15805 12924 15839
rect 12936 15805 12948 15863
rect 12960 15805 12972 15863
rect 12408 14677 12420 14711
rect 12432 14677 12444 14735
rect 12456 14677 12468 14735
rect 12480 14677 12492 14735
rect 12504 14677 12516 14735
rect 12528 14677 12540 14735
rect 12552 14677 12564 14735
rect 12576 14677 12588 14735
rect 12600 14677 12612 14735
rect 12624 14677 12636 14735
rect 12648 14677 12660 14735
rect 12672 14677 12684 14735
rect 12696 14677 12708 14735
rect 12720 14677 12732 14735
rect 12744 14677 12756 14735
rect 12768 14677 12780 14735
rect 12792 14677 12804 14735
rect 12816 14677 12828 14735
rect 12840 14677 12852 14735
rect 12864 14677 12876 14735
rect 12912 14653 12924 14711
rect 12936 14653 12948 14711
rect 12360 13477 12372 13511
rect 12384 13477 12396 13535
rect 12408 13477 12420 13535
rect 12432 13477 12444 13535
rect 12456 13477 12468 13535
rect 12480 13477 12492 13535
rect 12504 13477 12516 13535
rect 12528 13477 12540 13535
rect 12552 13477 12564 13535
rect 12576 13477 12588 13535
rect 12600 13477 12612 13535
rect 12624 13477 12636 13535
rect 12648 13477 12660 13535
rect 12672 13477 12684 13535
rect 12696 13477 12708 13535
rect 12720 13477 12732 13535
rect 12744 13477 12756 13535
rect 12768 13477 12780 13535
rect 12792 13477 12804 13535
rect 12816 13501 12828 13535
rect 12840 13453 12852 13535
rect 12864 13453 12876 13487
rect 12888 13453 12900 13511
rect 12912 13453 12924 13511
rect 12936 13453 12948 13511
rect 12960 13453 12972 13511
rect 5880 12613 5892 12647
rect 5904 12613 5916 12647
rect 43728 12613 43740 12647
rect 43752 12613 43764 12647
rect 43776 12613 43788 12647
rect 43704 12493 43716 12527
rect 43752 12469 43764 12503
rect 43776 12469 43788 12503
rect 12336 12325 12348 12359
rect 12360 12325 12372 12383
rect 12384 12325 12396 12383
rect 12432 12301 12444 12359
rect 12456 12301 12468 12359
rect 12480 12301 12492 12359
rect 12504 12301 12516 12359
rect 12528 12301 12540 12359
rect 12552 12301 12564 12359
rect 12576 12301 12588 12359
rect 12600 12301 12612 12359
rect 12624 12301 12636 12359
rect 12648 12301 12660 12359
rect 12672 12301 12684 12359
rect 12696 12301 12708 12359
rect 12720 12301 12732 12359
rect 12744 12301 12756 12359
rect 12768 12301 12780 12359
rect 12792 12301 12804 12359
rect 12816 12301 12828 12359
rect 12840 12301 12852 12359
rect 12864 12301 12876 12359
rect 12912 12277 12924 12335
rect 12936 12277 12948 12335
rect 12960 12277 12972 12335
rect 12312 11101 12324 11183
rect 12336 11101 12348 11135
rect 12360 11101 12372 11159
rect 12384 11101 12396 11159
rect 12408 11101 12420 11159
rect 12432 11101 12444 11159
rect 12456 11101 12468 11159
rect 12480 11101 12492 11159
rect 12504 11101 12516 11159
rect 12528 11101 12540 11159
rect 12552 11101 12564 11159
rect 12576 11101 12588 11159
rect 12600 11101 12612 11159
rect 12624 11101 12636 11159
rect 12648 11101 12660 11159
rect 12672 11101 12684 11159
rect 12696 11101 12708 11159
rect 12720 11101 12732 11159
rect 12744 11101 12756 11159
rect 12768 11101 12780 11159
rect 12792 11101 12804 11159
rect 12816 11101 12828 11159
rect 12840 11101 12852 11159
rect 12864 11101 12876 11159
rect 12888 11101 12900 11159
rect 12912 11101 12924 11159
rect 12936 11101 12948 11159
rect 12960 11101 12972 11159
rect 12240 9949 12252 9983
rect 12264 9949 12276 10007
rect 12288 9949 12300 10007
rect 12312 9949 12324 10007
rect 12336 9949 12348 10007
rect 12360 9949 12372 10007
rect 12384 9949 12396 10007
rect 12408 9949 12420 10007
rect 12432 9949 12444 10007
rect 12456 9949 12468 10007
rect 12480 9949 12492 10007
rect 12504 9949 12516 10007
rect 12528 9949 12540 10007
rect 12552 9949 12564 10007
rect 12576 9949 12588 10007
rect 12600 9949 12612 10007
rect 12624 9949 12636 10007
rect 12648 9949 12660 10007
rect 12672 9949 12684 10007
rect 12696 9949 12708 10007
rect 12720 9949 12732 10007
rect 12744 9949 12756 10007
rect 12768 9949 12780 10007
rect 12792 9949 12804 10007
rect 12816 9949 12828 10007
rect 12840 9973 12852 10007
rect 12864 9925 12876 10007
rect 12888 9925 12900 9959
rect 12912 9925 12924 9983
rect 12936 9925 12948 9983
rect 12960 9925 12972 9983
rect 12240 9733 12252 9767
rect 12264 9709 12276 9767
rect 12288 9685 12300 9767
rect 12312 9661 12324 9767
rect 12336 9637 12348 9767
rect 12360 9613 12372 9767
rect 12384 9589 12396 9767
rect 12408 9565 12420 9767
rect 12432 9541 12444 9767
rect 12456 9517 12468 9767
rect 12480 9493 12492 9767
rect 12504 9469 12516 9767
rect 12528 9445 12540 9767
rect 12552 9421 12564 9767
rect 12576 9397 12588 9767
rect 12600 9373 12612 9767
rect 12624 9349 12636 9767
rect 12648 9325 12660 9767
rect 12672 9253 12684 9767
rect 12696 9229 12708 9767
rect 12720 9181 12732 9767
rect 12744 9157 12756 9767
rect 12768 9325 12780 9767
rect 12768 9109 12780 9287
rect 12792 9109 12804 9767
rect 12816 9109 12828 9767
rect 12840 9109 12852 9767
rect 12864 9109 12876 9767
rect 12888 9109 12900 9767
rect 12912 9109 12924 9767
rect 12936 9109 12948 9767
rect 12960 9109 12972 9767
rect 12984 9109 12996 9143
rect 13008 9109 13020 9719
rect 13104 9685 13116 9719
rect 13464 9685 13476 9792
rect 13599 9780 13611 9792
rect 13671 9780 13683 9792
rect 14943 9780 14955 9792
rect 15135 9780 15147 9792
rect 15927 9780 15939 9792
rect 16479 9780 16491 9792
rect 16695 9780 16707 9792
rect 17439 9780 17451 9792
rect 17607 9780 17619 9792
rect 17991 9780 18003 9792
rect 18183 9780 18195 9792
rect 18399 9780 18411 9792
rect 19143 9780 19155 9792
rect 19311 9780 19323 9792
rect 28719 9780 28731 9792
rect 28911 9780 28923 9792
rect 29151 9780 29163 9792
rect 36855 9780 36867 9792
rect 37599 9780 37611 9792
rect 13599 9768 13620 9780
rect 13671 9768 13692 9780
rect 14943 9768 14964 9780
rect 15135 9768 15156 9780
rect 15927 9768 15948 9780
rect 16479 9768 16500 9780
rect 16695 9768 16716 9780
rect 17439 9768 17460 9780
rect 17607 9768 17628 9780
rect 17991 9768 18012 9780
rect 18183 9768 18204 9780
rect 18399 9768 18420 9780
rect 19143 9768 19164 9780
rect 19311 9768 19332 9780
rect 28719 9768 28740 9780
rect 28911 9768 28932 9780
rect 29151 9768 29172 9780
rect 36855 9768 36876 9780
rect 37599 9768 37620 9780
rect 13032 9109 13044 9671
rect 13056 9109 13068 9647
rect 13080 9109 13092 9623
rect 13104 9589 13116 9623
rect 13104 9109 13116 9551
rect 13128 9157 13140 9623
rect 13152 9205 13164 9623
rect 13176 9229 13188 9623
rect 13200 9277 13212 9551
rect 13224 9229 13236 9575
rect 13488 9301 13500 9671
rect 13608 9661 13620 9768
rect 13680 9685 13692 9768
rect 13632 9325 13644 9647
rect 13704 9349 13716 9671
rect 14952 9301 14964 9768
rect 15144 9277 15156 9768
rect 13248 9229 13260 9263
rect 15936 9253 15948 9768
rect 15960 9229 15972 9671
rect 15984 9205 15996 9719
rect 16008 9253 16020 9719
rect 16032 9277 16044 9671
rect 16488 9541 16500 9768
rect 16512 9469 16524 9527
rect 16704 9493 16716 9768
rect 17448 9493 17460 9768
rect 16536 9325 16548 9455
rect 16032 9205 16044 9239
rect 16056 9229 16068 9263
rect 16560 9253 16572 9311
rect 16728 9277 16740 9479
rect 17472 9325 17484 9479
rect 17616 9397 17628 9768
rect 18000 9661 18012 9768
rect 18024 9397 18036 9647
rect 18192 9565 18204 9768
rect 17664 9325 17676 9359
rect 18192 9349 18204 9527
rect 18216 9373 18228 9527
rect 18240 9397 18252 9551
rect 18408 9445 18420 9768
rect 19152 9493 19164 9768
rect 18432 9397 18444 9431
rect 19176 9421 19188 9479
rect 19320 9445 19332 9768
rect 28728 9493 28740 9768
rect 28920 9637 28932 9768
rect 29160 9661 29172 9768
rect 36864 9661 36876 9768
rect 37608 9637 37620 9768
rect 38088 9637 38100 9767
rect 38112 9637 38124 9743
rect 38136 9613 38148 9791
rect 38160 9661 38172 9791
rect 38184 9685 38196 9791
rect 38088 9445 38100 9599
rect 38112 9565 38124 9599
rect 38160 9565 38172 9599
rect 38112 9445 38124 9479
rect 38136 9445 38148 9551
rect 5880 7453 5892 7487
rect 12816 6637 12828 6671
rect 6912 6517 6924 6551
rect 11352 6493 11364 6551
rect 11496 6493 11508 6575
rect 11544 6493 11556 6599
rect 12840 6589 12852 6671
rect 12864 6589 12876 6671
rect 12888 6565 12900 6671
rect 12912 6565 12924 6671
rect 12936 6541 12948 6671
rect 12960 6541 12972 6671
rect 12984 6517 12996 6671
rect 13008 6637 13020 6671
rect 13032 6565 13044 6671
rect 13008 6517 13020 6551
rect 15816 6493 15828 6695
rect 15984 6565 15996 6695
rect 15960 6493 15972 6551
rect 16008 6493 16020 6647
rect 20304 6565 20316 6671
rect 20280 6493 20292 6551
rect 20424 6493 20436 6623
rect 20472 6493 20484 6623
rect 29256 6589 29268 6623
rect 29232 6493 29244 6575
rect 29376 6493 29388 6599
rect 29424 6493 29436 6575
rect 33696 6493 33708 6551
rect 38088 6541 38100 6575
rect 33840 6493 33852 6527
rect 33888 6493 33900 6527
rect 38208 6517 38220 6551
rect 38328 6493 38340 6527
<< metal4 >>
rect 6166 49274 7726 50834
rect 10638 49274 12198 50834
rect 15110 49274 16670 50834
rect 19582 49274 21142 50834
rect 24054 49274 25614 50834
rect 28526 49274 30086 50834
rect 32998 49274 34558 50834
rect 37470 49274 39030 50834
rect 41942 49274 43502 50834
rect -544 42736 1016 44296
rect 48652 42736 50212 44296
rect -544 37576 1016 39136
rect 48652 37576 50212 39136
rect -544 32416 1016 33976
rect 48652 32416 50212 33976
rect -544 27256 1016 28816
rect 48652 27256 50212 28816
rect -544 22096 1016 23656
rect 48652 22096 50212 23656
rect -544 16936 1016 18496
rect 48652 16936 50212 18496
rect -544 11776 1016 13336
rect 48652 11776 50212 13336
rect -544 6616 1016 8176
rect 48652 6616 50212 8176
rect 6166 78 7726 1638
rect 10638 78 12198 1638
rect 15110 78 16670 1638
rect 19582 78 21142 1638
rect 24054 78 25614 1638
rect 28526 78 30086 1638
rect 32998 78 34558 1638
rect 37470 78 39030 1638
rect 41942 78 43502 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 -622 -1 0 50912
box 0 0 6450 6450
use fillpp_mt fillpp_mt_805
timestamp 1300117811
transform 0 -1 5914 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_804
timestamp 1300117811
transform 0 -1 6000 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_803
timestamp 1300117811
transform 0 -1 6086 1 0 44462
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 7806 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_802
timestamp 1300117811
transform 0 -1 7892 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_801
timestamp 1300117811
transform 0 -1 7978 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_800
timestamp 1300117811
transform 0 -1 8064 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_799
timestamp 1300117811
transform 0 -1 8150 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_798
timestamp 1300117811
transform 0 -1 8236 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_797
timestamp 1300117811
transform 0 -1 8322 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_796
timestamp 1300117811
transform 0 -1 8408 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_795
timestamp 1300117811
transform 0 -1 8494 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_794
timestamp 1300117811
transform 0 -1 8580 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_793
timestamp 1300117811
transform 0 -1 8666 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_792
timestamp 1300117811
transform 0 -1 8752 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_791
timestamp 1300117811
transform 0 -1 8838 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_790
timestamp 1300117811
transform 0 -1 8924 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_789
timestamp 1300117811
transform 0 -1 9010 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_788
timestamp 1300117811
transform 0 -1 9096 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform 0 -1 9182 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform 0 -1 9268 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform 0 -1 9354 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform 0 -1 9440 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform 0 -1 9526 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform 0 -1 9612 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform 0 -1 9698 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform 0 -1 9784 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform 0 -1 9870 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform 0 -1 9956 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform 0 -1 10042 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform 0 -1 10128 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform 0 -1 10214 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform 0 -1 10300 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform 0 -1 10386 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform 0 -1 10472 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform 0 -1 10558 1 0 44462
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 12278 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform 0 -1 12364 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform 0 -1 12450 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform 0 -1 12536 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform 0 -1 12622 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform 0 -1 12708 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform 0 -1 12794 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform 0 -1 12880 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform 0 -1 12966 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform 0 -1 13052 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform 0 -1 13138 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform 0 -1 13224 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform 0 -1 13310 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform 0 -1 13396 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform 0 -1 13482 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform 0 -1 13568 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform 0 -1 13654 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform 0 -1 13740 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform 0 -1 13826 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform 0 -1 13912 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform 0 -1 13998 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform 0 -1 14084 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform 0 -1 14170 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform 0 -1 14256 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform 0 -1 14342 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform 0 -1 14428 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform 0 -1 14514 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform 0 -1 14600 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform 0 -1 14686 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform 0 -1 14772 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform 0 -1 14858 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform 0 -1 14944 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform 0 -1 15030 1 0 44462
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 16750 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform 0 -1 16836 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform 0 -1 16922 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform 0 -1 17008 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform 0 -1 17094 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform 0 -1 17180 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform 0 -1 17266 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform 0 -1 17352 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform 0 -1 17438 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform 0 -1 17524 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform 0 -1 17610 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform 0 -1 17696 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform 0 -1 17782 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform 0 -1 17868 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform 0 -1 17954 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform 0 -1 18040 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform 0 -1 18126 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform 0 -1 18212 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform 0 -1 18298 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform 0 -1 18384 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform 0 -1 18470 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform 0 -1 18556 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform 0 -1 18642 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform 0 -1 18728 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform 0 -1 18814 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform 0 -1 18900 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform 0 -1 18986 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform 0 -1 19072 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform 0 -1 19158 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform 0 -1 19244 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform 0 -1 19330 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform 0 -1 19416 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform 0 -1 19502 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 21222 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform 0 -1 21308 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform 0 -1 21394 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform 0 -1 21480 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform 0 -1 21566 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform 0 -1 21652 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform 0 -1 21738 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform 0 -1 21824 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform 0 -1 21910 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform 0 -1 21996 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform 0 -1 22082 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform 0 -1 22168 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform 0 -1 22254 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform 0 -1 22340 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform 0 -1 22426 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform 0 -1 22512 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform 0 -1 22598 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform 0 -1 22684 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform 0 -1 22770 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform 0 -1 22856 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform 0 -1 22942 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform 0 -1 23028 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform 0 -1 23114 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform 0 -1 23200 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform 0 -1 23286 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform 0 -1 23372 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform 0 -1 23458 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform 0 -1 23544 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform 0 -1 23630 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform 0 -1 23716 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform 0 -1 23802 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform 0 -1 23888 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform 0 -1 23974 1 0 44462
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 25694 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform 0 -1 25780 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform 0 -1 25866 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform 0 -1 25952 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform 0 -1 26038 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform 0 -1 26124 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform 0 -1 26210 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform 0 -1 26296 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform 0 -1 26382 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform 0 -1 26468 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform 0 -1 26554 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform 0 -1 26640 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform 0 -1 26726 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform 0 -1 26812 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform 0 -1 26898 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform 0 -1 26984 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform 0 -1 27070 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform 0 -1 27156 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform 0 -1 27242 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform 0 -1 27328 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform 0 -1 27414 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform 0 -1 27500 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform 0 -1 27586 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform 0 -1 27672 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform 0 -1 27758 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform 0 -1 27844 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform 0 -1 27930 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform 0 -1 28016 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform 0 -1 28102 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform 0 -1 28188 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform 0 -1 28274 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform 0 -1 28360 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform 0 -1 28446 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 30166 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform 0 -1 30252 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform 0 -1 30338 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform 0 -1 30424 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform 0 -1 30510 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform 0 -1 30596 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform 0 -1 30682 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform 0 -1 30768 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform 0 -1 30854 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform 0 -1 30940 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform 0 -1 31026 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform 0 -1 31112 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform 0 -1 31198 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform 0 -1 31284 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform 0 -1 31370 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform 0 -1 31456 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform 0 -1 31542 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform 0 -1 31628 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform 0 -1 31714 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform 0 -1 31800 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform 0 -1 31886 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform 0 -1 31972 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform 0 -1 32058 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform 0 -1 32144 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform 0 -1 32230 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform 0 -1 32316 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform 0 -1 32402 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform 0 -1 32488 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform 0 -1 32574 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform 0 -1 32660 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform 0 -1 32746 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform 0 -1 32832 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform 0 -1 32918 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 34638 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform 0 -1 34724 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform 0 -1 34810 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform 0 -1 34896 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform 0 -1 34982 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform 0 -1 35068 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform 0 -1 35154 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform 0 -1 35240 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform 0 -1 35326 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform 0 -1 35412 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform 0 -1 35498 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform 0 -1 35584 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform 0 -1 35670 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform 0 -1 35756 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform 0 -1 35842 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform 0 -1 35928 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform 0 -1 36014 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform 0 -1 36100 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform 0 -1 36186 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform 0 -1 36272 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform 0 -1 36358 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform 0 -1 36444 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform 0 -1 36530 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform 0 -1 36616 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform 0 -1 36702 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform 0 -1 36788 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform 0 -1 36874 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform 0 -1 36960 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform 0 -1 37046 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform 0 -1 37132 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform 0 -1 37218 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform 0 -1 37304 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform 0 -1 37390 1 0 44462
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 39110 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform 0 -1 39196 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform 0 -1 39282 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform 0 -1 39368 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform 0 -1 39454 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform 0 -1 39540 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform 0 -1 39626 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform 0 -1 39712 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform 0 -1 39798 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform 0 -1 39884 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform 0 -1 39970 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform 0 -1 40056 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform 0 -1 40142 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform 0 -1 40228 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform 0 -1 40314 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform 0 -1 40400 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 40486 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 40572 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 40658 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 40744 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 40830 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 40916 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 41002 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 41088 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 41174 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 41260 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 41346 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 41432 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 41518 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 41604 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 41690 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 41776 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 41862 1 0 44462
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 43582 1 0 44462
box 0 0 6450 1720
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 43668 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 43754 1 0 44462
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 43840 1 0 44462
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 50290 0 -1 50912
box 0 0 6450 6450
use fillpp_mt fillpp_mt_806
timestamp 1300117811
transform -1 0 5828 0 -1 44462
box 0 0 6450 86
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 5828 0 -1 44376
box 0 0 6450 1720
use fillpp_mt fillpp_mt_807
timestamp 1300117811
transform -1 0 5828 0 -1 42656
box 0 0 6450 86
use fillpp_mt fillpp_mt_808
timestamp 1300117811
transform -1 0 5828 0 -1 42570
box 0 0 6450 86
use fillpp_mt fillpp_mt_809
timestamp 1300117811
transform -1 0 5828 0 -1 42484
box 0 0 6450 86
use fillpp_mt fillpp_mt_810
timestamp 1300117811
transform -1 0 5828 0 -1 42398
box 0 0 6450 86
use fillpp_mt fillpp_mt_811
timestamp 1300117811
transform -1 0 5828 0 -1 42312
box 0 0 6450 86
use fillpp_mt fillpp_mt_812
timestamp 1300117811
transform -1 0 5828 0 -1 42226
box 0 0 6450 86
use fillpp_mt fillpp_mt_813
timestamp 1300117811
transform -1 0 5828 0 -1 42140
box 0 0 6450 86
use fillpp_mt fillpp_mt_814
timestamp 1300117811
transform -1 0 5828 0 -1 42054
box 0 0 6450 86
use fillpp_mt fillpp_mt_815
timestamp 1300117811
transform -1 0 5828 0 -1 41968
box 0 0 6450 86
use fillpp_mt fillpp_mt_816
timestamp 1300117811
transform -1 0 5828 0 -1 41882
box 0 0 6450 86
use fillpp_mt fillpp_mt_817
timestamp 1300117811
transform -1 0 5828 0 -1 41796
box 0 0 6450 86
use fillpp_mt fillpp_mt_818
timestamp 1300117811
transform -1 0 5828 0 -1 41710
box 0 0 6450 86
use fillpp_mt fillpp_mt_819
timestamp 1300117811
transform -1 0 5828 0 -1 41624
box 0 0 6450 86
use fillpp_mt fillpp_mt_820
timestamp 1300117811
transform -1 0 5828 0 -1 41538
box 0 0 6450 86
use fillpp_mt fillpp_mt_821
timestamp 1300117811
transform -1 0 5828 0 -1 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_822
timestamp 1300117811
transform -1 0 5828 0 -1 41366
box 0 0 6450 86
use fillpp_mt fillpp_mt_823
timestamp 1300117811
transform -1 0 5828 0 -1 41280
box 0 0 6450 86
use fillpp_mt fillpp_mt_824
timestamp 1300117811
transform -1 0 5828 0 -1 41194
box 0 0 6450 86
use fillpp_mt fillpp_mt_825
timestamp 1300117811
transform -1 0 5828 0 -1 41108
box 0 0 6450 86
use fillpp_mt fillpp_mt_826
timestamp 1300117811
transform -1 0 5828 0 -1 41022
box 0 0 6450 86
use fillpp_mt fillpp_mt_827
timestamp 1300117811
transform -1 0 5828 0 -1 40936
box 0 0 6450 86
use fillpp_mt fillpp_mt_828
timestamp 1300117811
transform -1 0 5828 0 -1 40850
box 0 0 6450 86
use fillpp_mt fillpp_mt_829
timestamp 1300117811
transform -1 0 5828 0 -1 40764
box 0 0 6450 86
use fillpp_mt fillpp_mt_830
timestamp 1300117811
transform -1 0 5828 0 -1 40678
box 0 0 6450 86
use fillpp_mt fillpp_mt_831
timestamp 1300117811
transform -1 0 5828 0 -1 40592
box 0 0 6450 86
use fillpp_mt fillpp_mt_832
timestamp 1300117811
transform -1 0 5828 0 -1 40506
box 0 0 6450 86
use fillpp_mt fillpp_mt_833
timestamp 1300117811
transform -1 0 5828 0 -1 40420
box 0 0 6450 86
use fillpp_mt fillpp_mt_834
timestamp 1300117811
transform -1 0 5828 0 -1 40334
box 0 0 6450 86
use fillpp_mt fillpp_mt_835
timestamp 1300117811
transform -1 0 5828 0 -1 40248
box 0 0 6450 86
use fillpp_mt fillpp_mt_836
timestamp 1300117811
transform -1 0 5828 0 -1 40162
box 0 0 6450 86
use fillpp_mt fillpp_mt_837
timestamp 1300117811
transform -1 0 5828 0 -1 40076
box 0 0 6450 86
use fillpp_mt fillpp_mt_838
timestamp 1300117811
transform -1 0 5828 0 -1 39990
box 0 0 6450 86
use fillpp_mt fillpp_mt_839
timestamp 1300117811
transform -1 0 5828 0 -1 39904
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 1 0 43840 0 1 44376
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 43840 0 1 42656
box 0 0 6450 1720
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 1 0 43840 0 1 42570
box 0 0 6450 86
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 1 0 43840 0 1 42484
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 1 0 43840 0 1 42398
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 1 0 43840 0 1 42312
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 1 0 43840 0 1 42226
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 1 0 43840 0 1 42140
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 1 0 43840 0 1 42054
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 1 0 43840 0 1 41968
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 1 0 43840 0 1 41882
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 1 0 43840 0 1 41796
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 1 0 43840 0 1 41710
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 1 0 43840 0 1 41624
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 1 0 43840 0 1 41538
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 1 0 43840 0 1 41452
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 1 0 43840 0 1 41366
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 1 0 43840 0 1 41280
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 1 0 43840 0 1 41194
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 1 0 43840 0 1 41108
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 1 0 43840 0 1 41022
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 1 0 43840 0 1 40936
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 1 0 43840 0 1 40850
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 1 0 43840 0 1 40764
box 0 0 6450 86
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 1 0 43840 0 1 40678
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 1 0 43840 0 1 40592
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 1 0 43840 0 1 40506
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 1 0 43840 0 1 40420
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 1 0 43840 0 1 40334
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 1 0 43840 0 1 40248
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 1 0 43840 0 1 40162
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 1 0 43840 0 1 40076
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 1 0 43840 0 1 39990
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 1 0 43840 0 1 39904
box 0 0 6450 86
use fillpp_mt fillpp_mt_840
timestamp 1300117811
transform -1 0 5828 0 -1 39818
box 0 0 6450 86
use fillpp_mt fillpp_mt_841
timestamp 1300117811
transform -1 0 5828 0 -1 39732
box 0 0 6450 86
use fillpp_mt fillpp_mt_842
timestamp 1300117811
transform -1 0 5828 0 -1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_843
timestamp 1300117811
transform -1 0 5828 0 -1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_844
timestamp 1300117811
transform -1 0 5828 0 -1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_845
timestamp 1300117811
transform -1 0 5828 0 -1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_846
timestamp 1300117811
transform -1 0 5828 0 -1 39302
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 5828 0 -1 39216
box 0 0 6450 1720
use fillpp_mt fillpp_mt_847
timestamp 1300117811
transform -1 0 5828 0 -1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_848
timestamp 1300117811
transform -1 0 5828 0 -1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_849
timestamp 1300117811
transform -1 0 5828 0 -1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_850
timestamp 1300117811
transform -1 0 5828 0 -1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_851
timestamp 1300117811
transform -1 0 5828 0 -1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_852
timestamp 1300117811
transform -1 0 5828 0 -1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_853
timestamp 1300117811
transform -1 0 5828 0 -1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_854
timestamp 1300117811
transform -1 0 5828 0 -1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_855
timestamp 1300117811
transform -1 0 5828 0 -1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_856
timestamp 1300117811
transform -1 0 5828 0 -1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_857
timestamp 1300117811
transform -1 0 5828 0 -1 36636
box 0 0 6450 86
use fillpp_mt fillpp_mt_858
timestamp 1300117811
transform -1 0 5828 0 -1 36550
box 0 0 6450 86
use fillpp_mt fillpp_mt_859
timestamp 1300117811
transform -1 0 5828 0 -1 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_860
timestamp 1300117811
transform -1 0 5828 0 -1 36378
box 0 0 6450 86
use fillpp_mt fillpp_mt_861
timestamp 1300117811
transform -1 0 5828 0 -1 36292
box 0 0 6450 86
use fillpp_mt fillpp_mt_862
timestamp 1300117811
transform -1 0 5828 0 -1 36206
box 0 0 6450 86
use fillpp_mt fillpp_mt_863
timestamp 1300117811
transform -1 0 5828 0 -1 36120
box 0 0 6450 86
use fillpp_mt fillpp_mt_864
timestamp 1300117811
transform -1 0 5828 0 -1 36034
box 0 0 6450 86
use fillpp_mt fillpp_mt_865
timestamp 1300117811
transform -1 0 5828 0 -1 35948
box 0 0 6450 86
use fillpp_mt fillpp_mt_866
timestamp 1300117811
transform -1 0 5828 0 -1 35862
box 0 0 6450 86
use fillpp_mt fillpp_mt_867
timestamp 1300117811
transform -1 0 5828 0 -1 35776
box 0 0 6450 86
use fillpp_mt fillpp_mt_868
timestamp 1300117811
transform -1 0 5828 0 -1 35690
box 0 0 6450 86
use fillpp_mt fillpp_mt_869
timestamp 1300117811
transform -1 0 5828 0 -1 35604
box 0 0 6450 86
use fillpp_mt fillpp_mt_870
timestamp 1300117811
transform -1 0 5828 0 -1 35518
box 0 0 6450 86
use fillpp_mt fillpp_mt_871
timestamp 1300117811
transform -1 0 5828 0 -1 35432
box 0 0 6450 86
use fillpp_mt fillpp_mt_872
timestamp 1300117811
transform -1 0 5828 0 -1 35346
box 0 0 6450 86
use fillpp_mt fillpp_mt_873
timestamp 1300117811
transform -1 0 5828 0 -1 35260
box 0 0 6450 86
use fillpp_mt fillpp_mt_874
timestamp 1300117811
transform -1 0 5828 0 -1 35174
box 0 0 6450 86
use fillpp_mt fillpp_mt_875
timestamp 1300117811
transform -1 0 5828 0 -1 35088
box 0 0 6450 86
use fillpp_mt fillpp_mt_876
timestamp 1300117811
transform -1 0 5828 0 -1 35002
box 0 0 6450 86
use fillpp_mt fillpp_mt_877
timestamp 1300117811
transform -1 0 5828 0 -1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_878
timestamp 1300117811
transform -1 0 5828 0 -1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_879
timestamp 1300117811
transform -1 0 5828 0 -1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_880
timestamp 1300117811
transform -1 0 5828 0 -1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_881
timestamp 1300117811
transform -1 0 5828 0 -1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_882
timestamp 1300117811
transform -1 0 5828 0 -1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_883
timestamp 1300117811
transform -1 0 5828 0 -1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_884
timestamp 1300117811
transform -1 0 5828 0 -1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_885
timestamp 1300117811
transform -1 0 5828 0 -1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_886
timestamp 1300117811
transform -1 0 5828 0 -1 34142
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 5828 0 -1 34056
box 0 0 6450 1720
use fillpp_mt fillpp_mt_887
timestamp 1300117811
transform -1 0 5828 0 -1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_888
timestamp 1300117811
transform -1 0 5828 0 -1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_889
timestamp 1300117811
transform -1 0 5828 0 -1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_890
timestamp 1300117811
transform -1 0 5828 0 -1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_891
timestamp 1300117811
transform -1 0 5828 0 -1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_892
timestamp 1300117811
transform -1 0 5828 0 -1 31906
box 0 0 6450 86
use fillpp_mt fillpp_mt_893
timestamp 1300117811
transform -1 0 5828 0 -1 31820
box 0 0 6450 86
use fillpp_mt fillpp_mt_894
timestamp 1300117811
transform -1 0 5828 0 -1 31734
box 0 0 6450 86
use fillpp_mt fillpp_mt_895
timestamp 1300117811
transform -1 0 5828 0 -1 31648
box 0 0 6450 86
use control control_0
timestamp 1395354352
transform 1 0 14508 0 1 31594
box -1500 0 25683 8276
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 1 0 43840 0 1 39818
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 1 0 43840 0 1 39732
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 1 0 43840 0 1 39646
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 1 0 43840 0 1 39560
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 1 0 43840 0 1 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 1 0 43840 0 1 39388
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 1 0 43840 0 1 39302
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 1 0 43840 0 1 39216
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 43840 0 1 37496
box 0 0 6450 1720
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 1 0 43840 0 1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 1 0 43840 0 1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 1 0 43840 0 1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 1 0 43840 0 1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 1 0 43840 0 1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 1 0 43840 0 1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 1 0 43840 0 1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 1 0 43840 0 1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 1 0 43840 0 1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 1 0 43840 0 1 36636
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 1 0 43840 0 1 36550
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 1 0 43840 0 1 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 1 0 43840 0 1 36378
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 1 0 43840 0 1 36292
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 1 0 43840 0 1 36206
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 1 0 43840 0 1 36120
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 1 0 43840 0 1 36034
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 1 0 43840 0 1 35948
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 1 0 43840 0 1 35862
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 1 0 43840 0 1 35776
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 1 0 43840 0 1 35690
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 1 0 43840 0 1 35604
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 1 0 43840 0 1 35518
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 1 0 43840 0 1 35432
box 0 0 6450 86
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 1 0 43840 0 1 35346
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 1 0 43840 0 1 35260
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 1 0 43840 0 1 35174
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 1 0 43840 0 1 35088
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 1 0 43840 0 1 35002
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 1 0 43840 0 1 34916
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 1 0 43840 0 1 34830
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 1 0 43840 0 1 34744
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 1 0 43840 0 1 34658
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 1 0 43840 0 1 34572
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 1 0 43840 0 1 34486
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 1 0 43840 0 1 34400
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 1 0 43840 0 1 34314
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 1 0 43840 0 1 34228
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 1 0 43840 0 1 34142
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 1 0 43840 0 1 34056
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 43840 0 1 32336
box 0 0 6450 1720
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 1 0 43840 0 1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 1 0 43840 0 1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 1 0 43840 0 1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 1 0 43840 0 1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 1 0 43840 0 1 31906
box 0 0 6450 86
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 1 0 43840 0 1 31820
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 1 0 43840 0 1 31734
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 1 0 43840 0 1 31648
box 0 0 6450 86
use fillpp_mt fillpp_mt_896
timestamp 1300117811
transform -1 0 5828 0 -1 31562
box 0 0 6450 86
use fillpp_mt fillpp_mt_897
timestamp 1300117811
transform -1 0 5828 0 -1 31476
box 0 0 6450 86
use fillpp_mt fillpp_mt_898
timestamp 1300117811
transform -1 0 5828 0 -1 31390
box 0 0 6450 86
use fillpp_mt fillpp_mt_899
timestamp 1300117811
transform -1 0 5828 0 -1 31304
box 0 0 6450 86
use fillpp_mt fillpp_mt_900
timestamp 1300117811
transform -1 0 5828 0 -1 31218
box 0 0 6450 86
use fillpp_mt fillpp_mt_901
timestamp 1300117811
transform -1 0 5828 0 -1 31132
box 0 0 6450 86
use fillpp_mt fillpp_mt_902
timestamp 1300117811
transform -1 0 5828 0 -1 31046
box 0 0 6450 86
use fillpp_mt fillpp_mt_903
timestamp 1300117811
transform -1 0 5828 0 -1 30960
box 0 0 6450 86
use fillpp_mt fillpp_mt_904
timestamp 1300117811
transform -1 0 5828 0 -1 30874
box 0 0 6450 86
use fillpp_mt fillpp_mt_905
timestamp 1300117811
transform -1 0 5828 0 -1 30788
box 0 0 6450 86
use fillpp_mt fillpp_mt_906
timestamp 1300117811
transform -1 0 5828 0 -1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_907
timestamp 1300117811
transform -1 0 5828 0 -1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_908
timestamp 1300117811
transform -1 0 5828 0 -1 30530
box 0 0 6450 86
use fillpp_mt fillpp_mt_909
timestamp 1300117811
transform -1 0 5828 0 -1 30444
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 1 0 43840 0 1 31562
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 1 0 43840 0 1 31476
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 1 0 43840 0 1 31390
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 1 0 43840 0 1 31304
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 1 0 43840 0 1 31218
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 1 0 43840 0 1 31132
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 1 0 43840 0 1 31046
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 1 0 43840 0 1 30960
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 1 0 43840 0 1 30874
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 1 0 43840 0 1 30788
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 1 0 43840 0 1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 1 0 43840 0 1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 1 0 43840 0 1 30530
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 1 0 43840 0 1 30444
box 0 0 6450 86
use fillpp_mt fillpp_mt_910
timestamp 1300117811
transform -1 0 5828 0 -1 30358
box 0 0 6450 86
use fillpp_mt fillpp_mt_911
timestamp 1300117811
transform -1 0 5828 0 -1 30272
box 0 0 6450 86
use fillpp_mt fillpp_mt_912
timestamp 1300117811
transform -1 0 5828 0 -1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_913
timestamp 1300117811
transform -1 0 5828 0 -1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_914
timestamp 1300117811
transform -1 0 5828 0 -1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_915
timestamp 1300117811
transform -1 0 5828 0 -1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_916
timestamp 1300117811
transform -1 0 5828 0 -1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_917
timestamp 1300117811
transform -1 0 5828 0 -1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_918
timestamp 1300117811
transform -1 0 5828 0 -1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_919
timestamp 1300117811
transform -1 0 5828 0 -1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_920
timestamp 1300117811
transform -1 0 5828 0 -1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_921
timestamp 1300117811
transform -1 0 5828 0 -1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_922
timestamp 1300117811
transform -1 0 5828 0 -1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_923
timestamp 1300117811
transform -1 0 5828 0 -1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_924
timestamp 1300117811
transform -1 0 5828 0 -1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_925
timestamp 1300117811
transform -1 0 5828 0 -1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_926
timestamp 1300117811
transform -1 0 5828 0 -1 28982
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 5828 0 -1 28896
box 0 0 6450 1720
use fillpp_mt fillpp_mt_927
timestamp 1300117811
transform -1 0 5828 0 -1 27176
box 0 0 6450 86
use fillpp_mt fillpp_mt_928
timestamp 1300117811
transform -1 0 5828 0 -1 27090
box 0 0 6450 86
use fillpp_mt fillpp_mt_929
timestamp 1300117811
transform -1 0 5828 0 -1 27004
box 0 0 6450 86
use fillpp_mt fillpp_mt_930
timestamp 1300117811
transform -1 0 5828 0 -1 26918
box 0 0 6450 86
use fillpp_mt fillpp_mt_931
timestamp 1300117811
transform -1 0 5828 0 -1 26832
box 0 0 6450 86
use fillpp_mt fillpp_mt_932
timestamp 1300117811
transform -1 0 5828 0 -1 26746
box 0 0 6450 86
use fillpp_mt fillpp_mt_933
timestamp 1300117811
transform -1 0 5828 0 -1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_934
timestamp 1300117811
transform -1 0 5828 0 -1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_935
timestamp 1300117811
transform -1 0 5828 0 -1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_936
timestamp 1300117811
transform -1 0 5828 0 -1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_937
timestamp 1300117811
transform -1 0 5828 0 -1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_938
timestamp 1300117811
transform -1 0 5828 0 -1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_939
timestamp 1300117811
transform -1 0 5828 0 -1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_940
timestamp 1300117811
transform -1 0 5828 0 -1 26058
box 0 0 6450 86
use fillpp_mt fillpp_mt_941
timestamp 1300117811
transform -1 0 5828 0 -1 25972
box 0 0 6450 86
use fillpp_mt fillpp_mt_942
timestamp 1300117811
transform -1 0 5828 0 -1 25886
box 0 0 6450 86
use fillpp_mt fillpp_mt_943
timestamp 1300117811
transform -1 0 5828 0 -1 25800
box 0 0 6450 86
use fillpp_mt fillpp_mt_944
timestamp 1300117811
transform -1 0 5828 0 -1 25714
box 0 0 6450 86
use fillpp_mt fillpp_mt_945
timestamp 1300117811
transform -1 0 5828 0 -1 25628
box 0 0 6450 86
use fillpp_mt fillpp_mt_946
timestamp 1300117811
transform -1 0 5828 0 -1 25542
box 0 0 6450 86
use fillpp_mt fillpp_mt_947
timestamp 1300117811
transform -1 0 5828 0 -1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_948
timestamp 1300117811
transform -1 0 5828 0 -1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_949
timestamp 1300117811
transform -1 0 5828 0 -1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_950
timestamp 1300117811
transform -1 0 5828 0 -1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_951
timestamp 1300117811
transform -1 0 5828 0 -1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_952
timestamp 1300117811
transform -1 0 5828 0 -1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_953
timestamp 1300117811
transform -1 0 5828 0 -1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_954
timestamp 1300117811
transform -1 0 5828 0 -1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_955
timestamp 1300117811
transform -1 0 5828 0 -1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_956
timestamp 1300117811
transform -1 0 5828 0 -1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_957
timestamp 1300117811
transform -1 0 5828 0 -1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_958
timestamp 1300117811
transform -1 0 5828 0 -1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_959
timestamp 1300117811
transform -1 0 5828 0 -1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_960
timestamp 1300117811
transform -1 0 5828 0 -1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_961
timestamp 1300117811
transform -1 0 5828 0 -1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_962
timestamp 1300117811
transform -1 0 5828 0 -1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_963
timestamp 1300117811
transform -1 0 5828 0 -1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_964
timestamp 1300117811
transform -1 0 5828 0 -1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_965
timestamp 1300117811
transform -1 0 5828 0 -1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_966
timestamp 1300117811
transform -1 0 5828 0 -1 23822
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 5828 0 -1 23736
box 0 0 6450 1720
use fillpp_mt fillpp_mt_967
timestamp 1300117811
transform -1 0 5828 0 -1 22016
box 0 0 6450 86
use fillpp_mt fillpp_mt_968
timestamp 1300117811
transform -1 0 5828 0 -1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_969
timestamp 1300117811
transform -1 0 5828 0 -1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_970
timestamp 1300117811
transform -1 0 5828 0 -1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_971
timestamp 1300117811
transform -1 0 5828 0 -1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_972
timestamp 1300117811
transform -1 0 5828 0 -1 21586
box 0 0 6450 86
use fillpp_mt fillpp_mt_973
timestamp 1300117811
transform -1 0 5828 0 -1 21500
box 0 0 6450 86
use fillpp_mt fillpp_mt_974
timestamp 1300117811
transform -1 0 5828 0 -1 21414
box 0 0 6450 86
use fillpp_mt fillpp_mt_975
timestamp 1300117811
transform -1 0 5828 0 -1 21328
box 0 0 6450 86
use fillpp_mt fillpp_mt_976
timestamp 1300117811
transform -1 0 5828 0 -1 21242
box 0 0 6450 86
use fillpp_mt fillpp_mt_977
timestamp 1300117811
transform -1 0 5828 0 -1 21156
box 0 0 6450 86
use fillpp_mt fillpp_mt_978
timestamp 1300117811
transform -1 0 5828 0 -1 21070
box 0 0 6450 86
use fillpp_mt fillpp_mt_979
timestamp 1300117811
transform -1 0 5828 0 -1 20984
box 0 0 6450 86
use fillpp_mt fillpp_mt_980
timestamp 1300117811
transform -1 0 5828 0 -1 20898
box 0 0 6450 86
use fillpp_mt fillpp_mt_981
timestamp 1300117811
transform -1 0 5828 0 -1 20812
box 0 0 6450 86
use fillpp_mt fillpp_mt_982
timestamp 1300117811
transform -1 0 5828 0 -1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_983
timestamp 1300117811
transform -1 0 5828 0 -1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_984
timestamp 1300117811
transform -1 0 5828 0 -1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_985
timestamp 1300117811
transform -1 0 5828 0 -1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_986
timestamp 1300117811
transform -1 0 5828 0 -1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_987
timestamp 1300117811
transform -1 0 5828 0 -1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_988
timestamp 1300117811
transform -1 0 5828 0 -1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_989
timestamp 1300117811
transform -1 0 5828 0 -1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_990
timestamp 1300117811
transform -1 0 5828 0 -1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_991
timestamp 1300117811
transform -1 0 5828 0 -1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_992
timestamp 1300117811
transform -1 0 5828 0 -1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_993
timestamp 1300117811
transform -1 0 5828 0 -1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_994
timestamp 1300117811
transform -1 0 5828 0 -1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_995
timestamp 1300117811
transform -1 0 5828 0 -1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_996
timestamp 1300117811
transform -1 0 5828 0 -1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_997
timestamp 1300117811
transform -1 0 5828 0 -1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_998
timestamp 1300117811
transform -1 0 5828 0 -1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_999
timestamp 1300117811
transform -1 0 5828 0 -1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_1000
timestamp 1300117811
transform -1 0 5828 0 -1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_1001
timestamp 1300117811
transform -1 0 5828 0 -1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_1002
timestamp 1300117811
transform -1 0 5828 0 -1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_1003
timestamp 1300117811
transform -1 0 5828 0 -1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_1004
timestamp 1300117811
transform -1 0 5828 0 -1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_1005
timestamp 1300117811
transform -1 0 5828 0 -1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_1006
timestamp 1300117811
transform -1 0 5828 0 -1 18662
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 5828 0 -1 18576
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1007
timestamp 1300117811
transform -1 0 5828 0 -1 16856
box 0 0 6450 86
use fillpp_mt fillpp_mt_1008
timestamp 1300117811
transform -1 0 5828 0 -1 16770
box 0 0 6450 86
use fillpp_mt fillpp_mt_1009
timestamp 1300117811
transform -1 0 5828 0 -1 16684
box 0 0 6450 86
use fillpp_mt fillpp_mt_1010
timestamp 1300117811
transform -1 0 5828 0 -1 16598
box 0 0 6450 86
use fillpp_mt fillpp_mt_1011
timestamp 1300117811
transform -1 0 5828 0 -1 16512
box 0 0 6450 86
use fillpp_mt fillpp_mt_1012
timestamp 1300117811
transform -1 0 5828 0 -1 16426
box 0 0 6450 86
use fillpp_mt fillpp_mt_1013
timestamp 1300117811
transform -1 0 5828 0 -1 16340
box 0 0 6450 86
use fillpp_mt fillpp_mt_1014
timestamp 1300117811
transform -1 0 5828 0 -1 16254
box 0 0 6450 86
use fillpp_mt fillpp_mt_1015
timestamp 1300117811
transform -1 0 5828 0 -1 16168
box 0 0 6450 86
use fillpp_mt fillpp_mt_1016
timestamp 1300117811
transform -1 0 5828 0 -1 16082
box 0 0 6450 86
use fillpp_mt fillpp_mt_1017
timestamp 1300117811
transform -1 0 5828 0 -1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_1018
timestamp 1300117811
transform -1 0 5828 0 -1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_1019
timestamp 1300117811
transform -1 0 5828 0 -1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_1020
timestamp 1300117811
transform -1 0 5828 0 -1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_1021
timestamp 1300117811
transform -1 0 5828 0 -1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_1022
timestamp 1300117811
transform -1 0 5828 0 -1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_1023
timestamp 1300117811
transform -1 0 5828 0 -1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_1024
timestamp 1300117811
transform -1 0 5828 0 -1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_1025
timestamp 1300117811
transform -1 0 5828 0 -1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_1026
timestamp 1300117811
transform -1 0 5828 0 -1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_1027
timestamp 1300117811
transform -1 0 5828 0 -1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_1028
timestamp 1300117811
transform -1 0 5828 0 -1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_1029
timestamp 1300117811
transform -1 0 5828 0 -1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_1030
timestamp 1300117811
transform -1 0 5828 0 -1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_1031
timestamp 1300117811
transform -1 0 5828 0 -1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_1032
timestamp 1300117811
transform -1 0 5828 0 -1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_1033
timestamp 1300117811
transform -1 0 5828 0 -1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_1034
timestamp 1300117811
transform -1 0 5828 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_1035
timestamp 1300117811
transform -1 0 5828 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_1036
timestamp 1300117811
transform -1 0 5828 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_1037
timestamp 1300117811
transform -1 0 5828 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_1038
timestamp 1300117811
transform -1 0 5828 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_1039
timestamp 1300117811
transform -1 0 5828 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_1040
timestamp 1300117811
transform -1 0 5828 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_1041
timestamp 1300117811
transform -1 0 5828 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_1042
timestamp 1300117811
transform -1 0 5828 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_1043
timestamp 1300117811
transform -1 0 5828 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_1044
timestamp 1300117811
transform -1 0 5828 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_1045
timestamp 1300117811
transform -1 0 5828 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_1046
timestamp 1300117811
transform -1 0 5828 0 -1 13502
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 5828 0 -1 13416
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1047
timestamp 1300117811
transform -1 0 5828 0 -1 11696
box 0 0 6450 86
use fillpp_mt fillpp_mt_1048
timestamp 1300117811
transform -1 0 5828 0 -1 11610
box 0 0 6450 86
use fillpp_mt fillpp_mt_1049
timestamp 1300117811
transform -1 0 5828 0 -1 11524
box 0 0 6450 86
use fillpp_mt fillpp_mt_1050
timestamp 1300117811
transform -1 0 5828 0 -1 11438
box 0 0 6450 86
use fillpp_mt fillpp_mt_1051
timestamp 1300117811
transform -1 0 5828 0 -1 11352
box 0 0 6450 86
use fillpp_mt fillpp_mt_1052
timestamp 1300117811
transform -1 0 5828 0 -1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_1053
timestamp 1300117811
transform -1 0 5828 0 -1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_1054
timestamp 1300117811
transform -1 0 5828 0 -1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_1055
timestamp 1300117811
transform -1 0 5828 0 -1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_1056
timestamp 1300117811
transform -1 0 5828 0 -1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_1057
timestamp 1300117811
transform -1 0 5828 0 -1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_1058
timestamp 1300117811
transform -1 0 5828 0 -1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_1059
timestamp 1300117811
transform -1 0 5828 0 -1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_1060
timestamp 1300117811
transform -1 0 5828 0 -1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_1061
timestamp 1300117811
transform -1 0 5828 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_1062
timestamp 1300117811
transform -1 0 5828 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_1063
timestamp 1300117811
transform -1 0 5828 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_1064
timestamp 1300117811
transform -1 0 5828 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_1065
timestamp 1300117811
transform -1 0 5828 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_1066
timestamp 1300117811
transform -1 0 5828 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_1067
timestamp 1300117811
transform -1 0 5828 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_1068
timestamp 1300117811
transform -1 0 5828 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_1069
timestamp 1300117811
transform -1 0 5828 0 -1 9804
box 0 0 6450 86
use datapath datapath_0
timestamp 1395340701
transform 1 0 12594 0 1 9749
box 414 43 25445 20615
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 1 0 43840 0 1 30358
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 1 0 43840 0 1 30272
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 1 0 43840 0 1 30186
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 1 0 43840 0 1 30100
box 0 0 6450 86
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 1 0 43840 0 1 30014
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 1 0 43840 0 1 29928
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 1 0 43840 0 1 29842
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 1 0 43840 0 1 29756
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 1 0 43840 0 1 29670
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 1 0 43840 0 1 29584
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 1 0 43840 0 1 29498
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 1 0 43840 0 1 29412
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 1 0 43840 0 1 29326
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 1 0 43840 0 1 29240
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 1 0 43840 0 1 29154
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 1 0 43840 0 1 29068
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 1 0 43840 0 1 28982
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 1 0 43840 0 1 28896
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 43840 0 1 27176
box 0 0 6450 1720
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 1 0 43840 0 1 27090
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 1 0 43840 0 1 27004
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 1 0 43840 0 1 26918
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 1 0 43840 0 1 26832
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 1 0 43840 0 1 26746
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 1 0 43840 0 1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 1 0 43840 0 1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 1 0 43840 0 1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 1 0 43840 0 1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 1 0 43840 0 1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 1 0 43840 0 1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 1 0 43840 0 1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 1 0 43840 0 1 26058
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 1 0 43840 0 1 25972
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 1 0 43840 0 1 25886
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 1 0 43840 0 1 25800
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 1 0 43840 0 1 25714
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 1 0 43840 0 1 25628
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 1 0 43840 0 1 25542
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 1 0 43840 0 1 25456
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 1 0 43840 0 1 25370
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 1 0 43840 0 1 25284
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 1 0 43840 0 1 25198
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 1 0 43840 0 1 25112
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 1 0 43840 0 1 25026
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 1 0 43840 0 1 24940
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 1 0 43840 0 1 24854
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 1 0 43840 0 1 24768
box 0 0 6450 86
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 1 0 43840 0 1 24682
box 0 0 6450 86
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 43840 0 1 24596
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 43840 0 1 24510
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 43840 0 1 24424
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 43840 0 1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 43840 0 1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 43840 0 1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 43840 0 1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 43840 0 1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 43840 0 1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 43840 0 1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 43840 0 1 23736
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 43840 0 1 22016
box 0 0 6450 1720
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 43840 0 1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 43840 0 1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 43840 0 1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 43840 0 1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 43840 0 1 21586
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 43840 0 1 21500
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 43840 0 1 21414
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 43840 0 1 21328
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 43840 0 1 21242
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 43840 0 1 21156
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 43840 0 1 21070
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 43840 0 1 20984
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 43840 0 1 20898
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 43840 0 1 20812
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 43840 0 1 20726
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 43840 0 1 20640
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 43840 0 1 20554
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 43840 0 1 20468
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 43840 0 1 20382
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 43840 0 1 20296
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 43840 0 1 20210
box 0 0 6450 86
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 43840 0 1 20124
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 43840 0 1 20038
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 43840 0 1 19952
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 43840 0 1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 43840 0 1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 43840 0 1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 43840 0 1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 43840 0 1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 43840 0 1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 43840 0 1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 43840 0 1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 43840 0 1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 43840 0 1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 43840 0 1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 43840 0 1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 43840 0 1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 43840 0 1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 43840 0 1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 43840 0 1 18576
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 43840 0 1 16856
box 0 0 6450 1720
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 43840 0 1 16770
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 43840 0 1 16684
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 43840 0 1 16598
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 43840 0 1 16512
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 43840 0 1 16426
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 43840 0 1 16340
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 43840 0 1 16254
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 43840 0 1 16168
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 43840 0 1 16082
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 43840 0 1 15996
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 43840 0 1 15910
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 43840 0 1 15824
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 43840 0 1 15738
box 0 0 6450 86
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 43840 0 1 15652
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 43840 0 1 15566
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 43840 0 1 15480
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 43840 0 1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 43840 0 1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 43840 0 1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 43840 0 1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 43840 0 1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 43840 0 1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 43840 0 1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 43840 0 1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 43840 0 1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 43840 0 1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 43840 0 1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 43840 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 43840 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 43840 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 43840 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 43840 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 43840 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 43840 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 43840 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 43840 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 43840 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 43840 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 43840 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 43840 0 1 13416
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 43840 0 1 11696
box 0 0 6450 1720
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 43840 0 1 11610
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 43840 0 1 11524
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 43840 0 1 11438
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 43840 0 1 11352
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 43840 0 1 11266
box 0 0 6450 86
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 43840 0 1 11180
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 43840 0 1 11094
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 43840 0 1 11008
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 43840 0 1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 43840 0 1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 43840 0 1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 43840 0 1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 43840 0 1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 43840 0 1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 43840 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 43840 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 43840 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 43840 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 43840 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 43840 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 43840 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 43840 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_1070
timestamp 1300117811
transform -1 0 5828 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_1071
timestamp 1300117811
transform -1 0 5828 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_1072
timestamp 1300117811
transform -1 0 5828 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_1073
timestamp 1300117811
transform -1 0 5828 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_1074
timestamp 1300117811
transform -1 0 5828 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_1075
timestamp 1300117811
transform -1 0 5828 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_1076
timestamp 1300117811
transform -1 0 5828 0 -1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_1077
timestamp 1300117811
transform -1 0 5828 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_1078
timestamp 1300117811
transform -1 0 5828 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_1079
timestamp 1300117811
transform -1 0 5828 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_1080
timestamp 1300117811
transform -1 0 5828 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_1081
timestamp 1300117811
transform -1 0 5828 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_1082
timestamp 1300117811
transform -1 0 5828 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_1083
timestamp 1300117811
transform -1 0 5828 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_1084
timestamp 1300117811
transform -1 0 5828 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_1085
timestamp 1300117811
transform -1 0 5828 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_1086
timestamp 1300117811
transform -1 0 5828 0 -1 8342
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 5828 0 -1 8256
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1087
timestamp 1300117811
transform -1 0 5828 0 -1 6536
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 43840 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 43840 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 43840 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 43840 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 43840 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 43840 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 43840 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 43840 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 43840 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 43840 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 43840 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 43840 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 43840 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 43840 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 43840 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 43840 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 43840 0 1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 43840 0 1 8256
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 43840 0 1 6536
box 0 0 6450 1720
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 43840 0 1 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 -622 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 5828 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 5914 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 6000 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6086 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 7806 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 7892 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 7978 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8064 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8150 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8236 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8322 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 8408 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 8494 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 8580 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 8666 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 8752 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 8838 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 8924 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9010 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9096 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9182 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9268 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9354 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 9440 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 9526 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 9612 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 9698 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 9784 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 9870 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 9956 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 10042 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 10128 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 10214 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 10300 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 10386 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 10472 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10558 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12278 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12364 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 12450 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 12536 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 12622 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 12708 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 12794 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 12880 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 12966 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 13052 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 13138 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 13224 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 13310 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 13396 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 13482 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 13568 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 13654 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 13740 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 13826 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 13912 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 13998 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 14084 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 14170 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 14256 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 14342 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 14428 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 14514 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 14600 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 14686 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 14772 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 14858 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 14944 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 15030 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 16750 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 16836 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 16922 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 17008 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 17094 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 17180 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 17266 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 17352 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 17438 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 17524 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 17610 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 17696 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 17782 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 17868 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 17954 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 18040 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 18126 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 18212 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 18298 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 18384 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 18470 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 18556 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 18642 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 18728 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 18814 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 18900 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 18986 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 19072 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 19158 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 19244 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 19330 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 19416 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 19502 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 21222 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 21308 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 21394 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 21480 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 21566 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 21652 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 21738 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 21824 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 21910 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 21996 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 22082 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 22168 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 22254 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 22340 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 22426 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 22512 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 22598 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 22684 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 22770 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 22856 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 22942 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 23028 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 23114 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 23200 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 23286 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 23372 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 23458 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 23544 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 23630 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 23716 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 23802 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 23888 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 23974 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 25694 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 25780 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 25866 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 25952 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 26038 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 26124 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 26210 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 26296 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 26382 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 26468 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 26554 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 26640 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 26726 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 26812 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 26898 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 26984 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 27070 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 27156 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 27242 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 27328 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 27414 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 27500 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 27586 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 27672 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 27758 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 27844 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 27930 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 28016 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 28102 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 28188 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 28274 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 28360 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 28446 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 30166 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 30252 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 30338 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 30424 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 30510 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 30596 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 30682 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 0 1 30768 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 0 1 30854 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 0 1 30940 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 0 1 31026 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 0 1 31112 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 0 1 31198 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 0 1 31284 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 0 1 31370 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 0 1 31456 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 0 1 31542 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 0 1 31628 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 0 1 31714 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 0 1 31800 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 0 1 31886 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 0 1 31972 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 0 1 32058 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 0 1 32144 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 0 1 32230 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 0 1 32316 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 0 1 32402 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 0 1 32488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 0 1 32574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 0 1 32660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 0 1 32746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 0 1 32832 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 32918 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 0 1 34638 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 0 1 34724 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 0 1 34810 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 0 1 34896 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 0 1 34982 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 0 1 35068 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 0 1 35154 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 0 1 35240 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 0 1 35326 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 0 1 35412 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 0 1 35498 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 0 1 35584 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 0 1 35670 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 0 1 35756 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 0 1 35842 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 0 1 35928 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 0 1 36014 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 0 1 36100 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 0 1 36186 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 0 1 36272 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 0 1 36358 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 0 1 36444 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 0 1 36530 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 0 1 36616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 0 1 36702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 0 1 36788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 0 1 36874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 0 1 36960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 0 1 37046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 0 1 37132 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 0 1 37218 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 0 1 37304 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 37390 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 0 1 39110 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 0 1 39196 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 0 1 39282 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 0 1 39368 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 0 1 39454 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 0 1 39540 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 0 1 39626 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 0 1 39712 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 0 1 39798 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 0 1 39884 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 0 1 39970 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 0 1 40056 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 0 1 40142 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 0 1 40228 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 0 1 40314 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 0 1 40400 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 0 1 40486 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 0 1 40572 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 0 1 40658 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 0 1 40744 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 0 1 40830 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 0 1 40916 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 0 1 41002 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 0 1 41088 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 0 1 41174 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 0 1 41260 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 0 1 41346 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 0 1 41432 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 0 1 41518 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 0 1 41604 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 0 1 41690 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 0 1 41776 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 41862 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 0 1 43582 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 0 1 43668 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 0 1 43754 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 50290 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 -544 6616 1016 8176 0 nReset
rlabel metal4 -544 11776 1016 13336 0 Clock
rlabel metal4 -544 16936 1016 18496 0 Test
rlabel metal4 -544 22096 1016 23656 0 SDI
rlabel metal4 -544 27256 1016 28816 0 Vdd!
rlabel metal4 -544 32416 1016 33976 0 SDO
rlabel metal4 -544 37576 1016 39136 0 RnW
rlabel metal4 -544 42736 1016 44296 0 nOE
rlabel metal4 6166 49274 7726 50834 0 nWait
rlabel metal4 10638 49274 12198 50834 0 nME
rlabel metal4 15110 49274 16670 50834 0 ALE
rlabel metal4 19582 49274 21142 50834 0 Data[15]
rlabel metal4 24054 49274 25614 50834 0 gnde!
rlabel metal4 28526 49274 30086 50834 0 Data[14]
rlabel metal4 32998 49274 34558 50834 0 Data[13]
rlabel metal4 37470 49274 39030 50834 0 Data[12]
rlabel metal4 41942 49274 43502 50834 0 vdde!
rlabel metal4 48652 42736 50212 44296 0 Data[11]
rlabel metal4 48652 37576 50212 39136 0 Data[10]
rlabel metal4 48652 32416 50212 33976 0 Data[9]
rlabel metal4 48652 27256 50212 28816 0 GND!
rlabel metal4 48652 22096 50212 23656 0 gnde!
rlabel metal4 48652 16936 50212 18496 0 Data[8]
rlabel metal4 48652 11776 50212 13336 0 Data[7]
rlabel metal4 48652 6616 50212 8176 0 Data[6]
rlabel metal4 41942 78 43502 1638 0 gnde!
rlabel metal4 37470 78 39030 1638 0 Data[5]
rlabel metal4 32998 78 34558 1638 0 Data[4]
rlabel metal4 28526 78 30086 1638 0 Data[3]
rlabel metal4 24054 78 25614 1638 0 vdde!
rlabel metal4 19582 78 21142 1638 0 Data[2]
rlabel metal4 15110 78 16670 1638 0 Data[1]
rlabel metal4 10638 78 12198 1638 0 Data[0]
rlabel metal4 6166 78 7726 1638 0 nIRQ
<< end >>
