magic
tech c035u
timestamp 1395431750
<< metal1 >>
rect 14464 8146 14482 8160
rect 18184 8148 18314 8158
rect 20560 8146 20578 8160
rect 22216 8146 22234 8160
rect 12880 8124 25694 8134
rect 4120 8100 18194 8110
rect 19720 8100 27178 8110
rect 3280 8076 4622 8086
rect 6904 8074 6922 8088
rect 10648 8076 19946 8086
rect 19960 8076 26090 8086
rect 2896 8052 22694 8062
rect 84 8028 8762 8038
rect 9136 8028 23738 8038
rect 24112 8028 24194 8038
rect 27033 8028 27565 8038
rect 84 8004 1730 8014
rect 2320 8004 27047 8014
rect 27112 8004 27146 8014
rect 27160 8004 27565 8014
rect 84 7980 10130 7990
rect 10720 7980 15194 7990
rect 18184 7980 27020 7990
rect 27139 7980 27565 7990
rect 3088 7956 23978 7966
rect 27061 7956 27565 7966
rect 3712 7932 27154 7942
rect 27192 7932 27565 7942
rect 4600 7908 7826 7918
rect 8896 7908 12182 7918
rect 12376 7908 27565 7918
rect 12160 7884 16658 7894
rect 18376 7884 27125 7894
rect 27168 7884 27565 7894
rect 14896 7051 14954 7061
rect 23944 7051 26138 7061
rect 13528 7027 24290 7037
rect 13432 7003 13706 7013
rect 13912 7003 14138 7013
rect 14512 7003 24122 7013
rect 12832 6979 24434 6989
rect 11992 6955 12842 6965
rect 13144 6955 23930 6965
rect 11944 6931 12386 6941
rect 12712 6931 13142 6941
rect 13288 6931 13970 6941
rect 13984 6931 17954 6941
rect 17968 6931 18722 6941
rect 11752 6907 11786 6917
rect 11896 6907 11954 6917
rect 12016 6907 12890 6917
rect 13096 6907 13898 6917
rect 13912 6907 17978 6917
rect 10432 6883 10826 6893
rect 11656 6883 16682 6893
rect 10216 6859 10466 6869
rect 10480 6859 12434 6869
rect 12448 6859 20018 6869
rect 20032 6859 24986 6869
rect 10120 6835 10514 6845
rect 11272 6835 13754 6845
rect 14272 6835 14330 6845
rect 14416 6835 14474 6845
rect 14560 6835 26234 6845
rect 10096 6811 17162 6821
rect 18568 6811 18866 6821
rect 9952 6787 24314 6797
rect 24328 6787 27218 6797
rect 9904 6763 11426 6773
rect 11608 6763 20690 6773
rect 9880 6739 14426 6749
rect 14440 6739 25010 6749
rect 9856 6715 13850 6725
rect 13864 6715 22754 6725
rect 23272 6715 26066 6725
rect 9760 6691 15410 6701
rect 15424 6691 18554 6701
rect 18568 6691 25394 6701
rect 9736 6667 10370 6677
rect 10384 6667 11834 6677
rect 11848 6667 22874 6677
rect 22888 6667 24242 6677
rect 9688 6643 10562 6653
rect 10816 6643 11618 6653
rect 11680 6643 11714 6653
rect 11824 6643 14210 6653
rect 14224 6643 18050 6653
rect 18064 6643 24146 6653
rect 9640 6619 14306 6629
rect 14392 6619 23570 6629
rect 9352 6595 11306 6605
rect 11320 6595 14882 6605
rect 14896 6595 17234 6605
rect 17248 6595 23258 6605
rect 9088 6571 15602 6581
rect 9064 6547 21050 6557
rect 21064 6547 27050 6557
rect 8968 6523 11090 6533
rect 11104 6523 12818 6533
rect 12832 6523 20378 6533
rect 20392 6523 23306 6533
rect 8944 6499 10298 6509
rect 10312 6499 12482 6509
rect 12496 6499 13730 6509
rect 13744 6499 18482 6509
rect 18496 6499 18842 6509
rect 18856 6499 21026 6509
rect 21040 6499 23330 6509
rect 8848 6475 23858 6485
rect 8752 6451 21530 6461
rect 8680 6427 16418 6437
rect 26368 6427 26594 6437
rect 8656 6403 26354 6413
rect 26368 6403 27170 6413
rect 8560 6379 14690 6389
rect 14848 6379 16778 6389
rect 20152 6379 24530 6389
rect 8536 6355 25346 6365
rect 8200 6331 11258 6341
rect 11272 6331 20210 6341
rect 20224 6331 21554 6341
rect 21568 6331 21986 6341
rect 22000 6331 25634 6341
rect 8080 6307 10586 6317
rect 10744 6307 21098 6317
rect 7792 6283 19826 6293
rect 20104 6283 20354 6293
rect 7624 6259 14834 6269
rect 15736 6259 15806 6269
rect 16552 6259 16658 6269
rect 19888 6259 19922 6269
rect 20008 6259 20282 6269
rect 21448 6259 21698 6269
rect 7600 6235 11306 6245
rect 11512 6235 14906 6245
rect 14920 6235 20114 6245
rect 20128 6235 25058 6245
rect 7432 6211 21434 6221
rect 7408 6187 17642 6197
rect 19792 6187 21218 6197
rect 21856 6187 21878 6197
rect 7312 6163 10322 6173
rect 10336 6163 23594 6173
rect 7216 6139 7706 6149
rect 7720 6139 14810 6149
rect 14824 6139 15722 6149
rect 15736 6139 18290 6149
rect 18304 6139 21650 6149
rect 21664 6139 21842 6149
rect 7048 6115 11042 6125
rect 11128 6115 14306 6125
rect 14320 6115 23786 6125
rect 7000 6091 18410 6101
rect 19648 6091 20666 6101
rect 6784 6067 7778 6077
rect 7792 6067 11234 6077
rect 11248 6067 11738 6077
rect 11752 6067 13658 6077
rect 13672 6067 13778 6077
rect 14128 6067 17090 6077
rect 17104 6067 22130 6077
rect 22144 6067 22646 6077
rect 6520 6043 6530 6053
rect 6592 6043 20954 6053
rect 6328 6019 12194 6029
rect 12280 6019 13286 6029
rect 13336 6019 13610 6029
rect 14080 6019 20522 6029
rect 6304 5995 11138 6005
rect 11224 5995 11282 6005
rect 11368 5995 23210 6005
rect 6064 5971 10226 5981
rect 10240 5971 22322 5981
rect 5968 5947 22586 5957
rect 22600 5947 25826 5957
rect 5872 5923 26738 5933
rect 5800 5899 6218 5909
rect 6232 5899 9890 5909
rect 9904 5899 11666 5909
rect 11680 5899 20450 5909
rect 24472 5899 25154 5909
rect 5728 5875 13586 5885
rect 13840 5875 14570 5885
rect 16408 5875 19970 5885
rect 20056 5875 26474 5885
rect 5632 5851 13538 5861
rect 13648 5851 17042 5861
rect 17056 5851 17594 5861
rect 17608 5851 23138 5861
rect 23152 5851 25106 5861
rect 5680 5827 21914 5837
rect 21928 5827 23450 5837
rect 23464 5827 25202 5837
rect 5512 5803 11858 5813
rect 11872 5803 12458 5813
rect 12472 5803 12986 5813
rect 13000 5803 16538 5813
rect 16552 5803 16802 5813
rect 19576 5803 24458 5813
rect 5464 5779 8642 5789
rect 8656 5779 8978 5789
rect 8992 5779 9290 5789
rect 9304 5779 16514 5789
rect 17392 5779 25778 5789
rect 5416 5755 7586 5765
rect 7600 5755 20594 5765
rect 5368 5731 10274 5741
rect 10288 5731 15746 5741
rect 15760 5731 16418 5741
rect 16432 5731 26690 5741
rect 5272 5707 24602 5717
rect 5224 5683 14522 5693
rect 16336 5683 16370 5693
rect 17368 5683 20210 5693
rect 26200 5683 26330 5693
rect 5200 5659 5834 5669
rect 5848 5659 6818 5669
rect 6832 5659 6914 5669
rect 6928 5659 26186 5669
rect 5176 5635 8330 5645
rect 8344 5635 21266 5645
rect 5104 5611 8570 5621
rect 8584 5611 13490 5621
rect 13504 5611 24242 5621
rect 24256 5611 25466 5621
rect 5008 5587 8402 5597
rect 8464 5587 15050 5597
rect 15592 5587 22730 5597
rect 4984 5563 10634 5573
rect 10648 5563 19322 5573
rect 19432 5563 24578 5573
rect 4888 5539 8306 5549
rect 8320 5539 10874 5549
rect 10888 5539 13922 5549
rect 13936 5539 18386 5549
rect 18400 5539 22706 5549
rect 22720 5539 24362 5549
rect 24376 5539 27122 5549
rect 4864 5515 9818 5525
rect 9832 5515 10850 5525
rect 10864 5515 11186 5525
rect 11200 5515 12938 5525
rect 12952 5515 13514 5525
rect 13528 5515 14078 5525
rect 14092 5515 17618 5525
rect 17632 5515 19298 5525
rect 19312 5515 20570 5525
rect 20584 5515 21194 5525
rect 21208 5515 22490 5525
rect 22504 5515 24338 5525
rect 4672 5491 9650 5501
rect 9664 5491 25730 5501
rect 26464 5491 26666 5501
rect 4600 5467 7538 5477
rect 7552 5467 21938 5477
rect 21952 5467 26450 5477
rect 4384 5443 26018 5453
rect 4312 5419 12674 5429
rect 12928 5419 13538 5429
rect 13552 5419 18002 5429
rect 18904 5419 21458 5429
rect 21472 5419 24074 5429
rect 4288 5395 16442 5405
rect 16840 5395 16874 5405
rect 16936 5395 17066 5405
rect 17296 5395 19034 5405
rect 19240 5395 20714 5405
rect 20896 5395 21674 5405
rect 4264 5371 4490 5381
rect 4504 5371 9938 5381
rect 9952 5371 11210 5381
rect 11224 5371 12962 5381
rect 12976 5371 14234 5381
rect 14248 5371 18818 5381
rect 18832 5371 18890 5381
rect 18904 5371 21122 5381
rect 21136 5371 25010 5381
rect 4072 5347 10658 5357
rect 10672 5347 18218 5357
rect 19144 5347 23690 5357
rect 4000 5323 7322 5333
rect 7336 5323 8618 5333
rect 8632 5323 11762 5333
rect 11776 5323 11882 5333
rect 11896 5323 12794 5333
rect 12808 5323 14402 5333
rect 14416 5323 22250 5333
rect 22264 5323 22466 5333
rect 3976 5299 6794 5309
rect 6808 5299 12770 5309
rect 12784 5299 20642 5309
rect 20656 5299 21818 5309
rect 21832 5299 23522 5309
rect 3904 5275 6146 5285
rect 6160 5275 10058 5285
rect 10072 5275 13034 5285
rect 13048 5275 13346 5285
rect 13360 5275 16706 5285
rect 16720 5275 20090 5285
rect 20104 5275 20462 5285
rect 20476 5275 20738 5285
rect 20752 5275 22346 5285
rect 22360 5275 25730 5285
rect 25744 5275 25970 5285
rect 3760 5251 14594 5261
rect 14752 5251 22994 5261
rect 3664 5227 10610 5237
rect 10624 5227 20978 5237
rect 3568 5203 6650 5213
rect 6664 5203 23006 5213
rect 3544 5179 22850 5189
rect 3496 5155 4778 5165
rect 4792 5155 11354 5165
rect 11416 5155 12578 5165
rect 12664 5155 23306 5165
rect 23416 5155 23486 5165
rect 3448 5131 10922 5141
rect 10984 5131 23834 5141
rect 3376 5107 26546 5117
rect 3352 5083 4706 5093
rect 4720 5083 7850 5093
rect 7864 5083 8162 5093
rect 8176 5083 14282 5093
rect 14296 5083 16154 5093
rect 16168 5083 16826 5093
rect 16840 5083 18626 5093
rect 18640 5083 21290 5093
rect 21304 5083 22274 5093
rect 22288 5083 23402 5093
rect 23416 5083 27146 5093
rect 3328 5059 7466 5069
rect 7480 5059 7922 5069
rect 8056 5059 10586 5069
rect 10600 5059 13682 5069
rect 13696 5059 18818 5069
rect 18832 5059 19682 5069
rect 19768 5059 22418 5069
rect 3256 5035 21962 5045
rect 21976 5035 23234 5045
rect 3232 5011 3794 5021
rect 3880 5011 10346 5021
rect 10360 5011 21290 5021
rect 21304 5011 26402 5021
rect 3136 4987 17762 4997
rect 18184 4987 18242 4997
rect 18328 4987 18338 4997
rect 19072 4987 21002 4997
rect 21328 4987 26762 4997
rect 3112 4963 9986 4973
rect 10072 4963 11786 4973
rect 11800 4963 20498 4973
rect 20848 4963 21578 4973
rect 21592 4963 25970 4973
rect 3016 4939 18770 4949
rect 18784 4939 19610 4949
rect 19672 4939 22034 4949
rect 22216 4939 25154 4949
rect 2968 4915 7802 4925
rect 7816 4915 8426 4925
rect 8440 4915 25250 4925
rect 2920 4891 14786 4901
rect 15568 4891 21350 4901
rect 22168 4891 22466 4901
rect 2824 4867 16610 4877
rect 16912 4867 16970 4877
rect 17128 4867 18458 4877
rect 19000 4867 23186 4877
rect 2776 4843 7682 4853
rect 7768 4843 8234 4853
rect 8248 4843 8258 4853
rect 8272 4843 23714 4853
rect 23728 4843 23906 4853
rect 2704 4819 10778 4829
rect 10792 4819 13418 4829
rect 13432 4819 16754 4829
rect 16768 4819 22562 4829
rect 2680 4795 8786 4805
rect 8800 4795 14162 4805
rect 14176 4795 17474 4805
rect 17488 4795 20162 4805
rect 20176 4795 24026 4805
rect 2632 4771 9410 4781
rect 9472 4771 15806 4781
rect 16288 4771 16850 4781
rect 16864 4771 19946 4781
rect 19960 4771 22538 4781
rect 2584 4747 10442 4757
rect 10504 4747 25682 4757
rect 2536 4723 20402 4733
rect 20776 4723 23162 4733
rect 2512 4699 10802 4709
rect 10816 4699 22514 4709
rect 2488 4675 6266 4685
rect 6280 4675 21386 4685
rect 21400 4675 24050 4685
rect 24064 4675 25130 4685
rect 2416 4651 18458 4661
rect 18472 4651 23378 4661
rect 2368 4627 13010 4637
rect 13072 4627 13442 4637
rect 13576 4627 26402 4637
rect 2296 4603 3674 4613
rect 3688 4603 9194 4613
rect 9208 4603 10634 4613
rect 10720 4603 26570 4613
rect 2248 4579 3194 4589
rect 3208 4579 18314 4589
rect 18664 4579 22430 4589
rect 2248 4555 25322 4565
rect 2224 4531 7730 4541
rect 7744 4531 11426 4541
rect 11440 4531 23954 4541
rect 2152 4507 3266 4517
rect 3280 4507 5930 4517
rect 5944 4507 7154 4517
rect 7168 4507 15866 4517
rect 15880 4507 16034 4517
rect 16048 4507 16922 4517
rect 16936 4507 18434 4517
rect 18448 4507 22058 4517
rect 22072 4507 23090 4517
rect 23104 4507 23546 4517
rect 2128 4483 24482 4493
rect 24880 4483 24890 4493
rect 1960 4459 3410 4469
rect 3424 4459 18194 4469
rect 18520 4459 26090 4469
rect 1912 4435 4826 4445
rect 4840 4435 5354 4445
rect 5368 4435 8282 4445
rect 8296 4435 13202 4445
rect 13216 4435 13874 4445
rect 14032 4435 18914 4445
rect 18928 4435 22010 4445
rect 22024 4435 26594 4445
rect 1888 4411 13178 4421
rect 13192 4411 24386 4421
rect 1840 4387 8714 4397
rect 8776 4387 19466 4397
rect 20080 4387 22802 4397
rect 22816 4387 25874 4397
rect 1816 4363 21602 4373
rect 21616 4363 22082 4373
rect 22096 4363 22610 4373
rect 22624 4363 22826 4373
rect 22840 4363 25226 4373
rect 1696 4339 17186 4349
rect 17776 4339 18338 4349
rect 18424 4339 18722 4349
rect 18856 4339 27098 4349
rect 1672 4315 4514 4325
rect 4528 4315 11330 4325
rect 11344 4315 16610 4325
rect 16768 4315 16778 4325
rect 17056 4315 19514 4325
rect 20656 4315 20666 4325
rect 21208 4315 21554 4325
rect 21640 4315 26786 4325
rect 1624 4291 2306 4301
rect 2320 4291 6650 4301
rect 6664 4291 8426 4301
rect 8440 4291 11930 4301
rect 11944 4291 12770 4301
rect 12784 4291 14258 4301
rect 14272 4291 19370 4301
rect 21280 4291 21650 4301
rect 22288 4291 22322 4301
rect 22624 4291 22646 4301
rect 22840 4291 23006 4301
rect 23536 4291 23570 4301
rect 84 4267 21770 4277
rect 84 4243 22226 4253
rect 84 4219 1994 4229
rect 2056 4219 19298 4229
rect 84 4195 14738 4205
rect 14944 4195 23666 4205
rect 1744 4171 6506 4181
rect 6688 4171 14186 4181
rect 14200 4171 15650 4181
rect 15808 4171 19202 4181
rect 19216 4171 25922 4181
rect 1792 4147 22634 4157
rect 2056 4123 4442 4133
rect 4456 4123 7514 4133
rect 7528 4123 16058 4133
rect 16072 4123 16730 4133
rect 16744 4123 23090 4133
rect 23104 4123 23690 4133
rect 23704 4123 26162 4133
rect 2104 4099 5690 4109
rect 5704 4099 7274 4109
rect 7288 4099 9866 4109
rect 9880 4099 12146 4109
rect 12160 4099 12698 4109
rect 12712 4099 14354 4109
rect 14368 4099 15962 4109
rect 15976 4099 21506 4109
rect 21520 4099 23066 4109
rect 23080 4099 26882 4109
rect 2176 4075 14690 4085
rect 16336 4075 25538 4085
rect 25552 4075 27098 4085
rect 2272 4051 14618 4061
rect 14728 4051 17522 4061
rect 17920 4051 18362 4061
rect 19024 4051 21794 4061
rect 23080 4051 23138 4061
rect 2296 4027 6866 4037
rect 6880 4027 22298 4037
rect 22312 4027 22394 4037
rect 2416 4003 7322 4013
rect 7336 4003 8210 4013
rect 8224 4003 11018 4013
rect 11032 4003 13802 4013
rect 13816 4003 14858 4013
rect 14872 4003 19994 4013
rect 20008 4003 20954 4013
rect 20968 4003 22706 4013
rect 22720 4003 24098 4013
rect 24112 4003 26306 4013
rect 26320 4003 26642 4013
rect 2512 3979 2594 3989
rect 2608 3979 5282 3989
rect 5296 3979 6578 3989
rect 6592 3979 6986 3989
rect 7000 3979 8834 3989
rect 8848 3979 9674 3989
rect 9688 3979 11162 3989
rect 11176 3979 16130 3989
rect 16144 3979 26498 3989
rect 26512 3979 26978 3989
rect 2536 3955 4610 3965
rect 4624 3955 4994 3965
rect 5008 3955 7058 3965
rect 7072 3955 7130 3965
rect 7144 3955 7874 3965
rect 7888 3955 8954 3965
rect 8968 3955 12002 3965
rect 12016 3955 12122 3965
rect 12136 3955 12242 3965
rect 12256 3955 17018 3965
rect 17032 3955 22106 3965
rect 22120 3955 22970 3965
rect 22984 3955 24866 3965
rect 24880 3955 25946 3965
rect 25960 3955 27002 3965
rect 2584 3931 7610 3941
rect 7624 3931 9506 3941
rect 9520 3931 10034 3941
rect 10048 3931 10754 3941
rect 10768 3931 15938 3941
rect 15952 3931 16898 3941
rect 18136 3931 20546 3941
rect 22408 3931 22430 3941
rect 2632 3907 3578 3917
rect 3592 3907 5570 3917
rect 5584 3907 13142 3917
rect 13156 3907 23810 3917
rect 23824 3907 25298 3917
rect 2728 3883 12602 3893
rect 12736 3883 17138 3893
rect 2776 3859 2882 3869
rect 2944 3859 6842 3869
rect 6952 3859 13370 3869
rect 13576 3859 19898 3869
rect 3064 3835 10418 3845
rect 10552 3835 24194 3845
rect 3088 3811 3626 3821
rect 3688 3811 16874 3821
rect 16888 3811 18602 3821
rect 18616 3811 19874 3821
rect 19888 3811 24914 3821
rect 24928 3811 25658 3821
rect 3184 3787 13058 3797
rect 13120 3787 14138 3797
rect 14152 3787 21878 3797
rect 21892 3787 23138 3797
rect 3328 3763 6122 3773
rect 6136 3763 7898 3773
rect 7912 3763 9530 3773
rect 9544 3763 10946 3773
rect 10960 3763 11978 3773
rect 11992 3763 18530 3773
rect 18544 3763 25754 3773
rect 3472 3739 3842 3749
rect 3856 3739 5810 3749
rect 5824 3739 7130 3749
rect 7144 3739 22778 3749
rect 22792 3739 26858 3749
rect 3544 3715 19082 3725
rect 19912 3715 19970 3725
rect 3616 3691 21722 3701
rect 3760 3667 19130 3677
rect 19144 3667 20186 3677
rect 20200 3667 21050 3677
rect 3808 3643 4178 3653
rect 4192 3643 11906 3653
rect 11920 3643 12170 3653
rect 12184 3643 12410 3653
rect 12424 3643 15770 3653
rect 15784 3643 16442 3653
rect 16456 3643 18746 3653
rect 18760 3643 21146 3653
rect 21160 3643 25610 3653
rect 25624 3643 26282 3653
rect 3832 3619 5138 3629
rect 5152 3619 6362 3629
rect 6376 3619 7490 3629
rect 7504 3619 7946 3629
rect 7960 3619 9842 3629
rect 9856 3619 10994 3629
rect 11008 3619 11546 3629
rect 11560 3619 12746 3629
rect 12760 3619 17066 3629
rect 17080 3619 17498 3629
rect 17512 3619 17570 3629
rect 17584 3619 20810 3629
rect 20824 3619 21242 3629
rect 21256 3619 22010 3629
rect 22024 3619 25778 3629
rect 25792 3619 26210 3629
rect 26296 3619 26474 3629
rect 3904 3595 4082 3605
rect 4192 3595 13466 3605
rect 13480 3595 18170 3605
rect 18184 3595 19922 3605
rect 19936 3595 23594 3605
rect 3928 3571 22994 3581
rect 3952 3547 12506 3557
rect 12520 3547 13394 3557
rect 13408 3547 23162 3557
rect 3976 3523 11474 3533
rect 11560 3523 13706 3533
rect 13720 3523 16562 3533
rect 16576 3523 23018 3533
rect 4000 3499 23642 3509
rect 4024 3475 9746 3485
rect 9976 3475 12050 3485
rect 12064 3475 14666 3485
rect 14680 3475 16346 3485
rect 16360 3475 26378 3485
rect 4048 3451 9266 3461
rect 9280 3451 9986 3461
rect 10000 3451 12218 3461
rect 12232 3451 12434 3461
rect 12448 3451 16586 3461
rect 18760 3451 19034 3461
rect 20200 3451 20462 3461
rect 4096 3427 4154 3437
rect 4216 3427 12626 3437
rect 12808 3427 16658 3437
rect 4264 3403 13442 3413
rect 13456 3403 18674 3413
rect 4288 3379 6530 3389
rect 6544 3379 7418 3389
rect 7432 3379 8354 3389
rect 8368 3379 10178 3389
rect 10192 3379 11282 3389
rect 11296 3379 13994 3389
rect 14008 3379 26426 3389
rect 4360 3355 6362 3365
rect 6424 3355 6434 3365
rect 6496 3355 8186 3365
rect 8200 3355 12890 3365
rect 12904 3355 14042 3365
rect 14176 3355 14210 3365
rect 14368 3355 14426 3365
rect 14584 3355 26810 3365
rect 4360 3331 12026 3341
rect 12040 3331 19538 3341
rect 4384 3307 6002 3317
rect 6016 3307 6338 3317
rect 6352 3307 12290 3317
rect 12304 3307 13322 3317
rect 13336 3307 16082 3317
rect 16096 3307 20306 3317
rect 20320 3307 20498 3317
rect 20512 3307 21410 3317
rect 21424 3307 23042 3317
rect 23056 3307 26618 3317
rect 4408 3283 12674 3293
rect 12688 3283 24650 3293
rect 4432 3259 12122 3269
rect 12184 3259 12362 3269
rect 12640 3259 12866 3269
rect 12976 3259 13286 3269
rect 13648 3259 13946 3269
rect 14008 3259 14078 3269
rect 20320 3259 20570 3269
rect 4480 3235 22418 3245
rect 4480 3211 4754 3221
rect 4768 3211 7250 3221
rect 7264 3211 10298 3221
rect 10312 3211 11474 3221
rect 11488 3211 12554 3221
rect 12568 3211 20234 3221
rect 20248 3211 24170 3221
rect 24184 3211 25202 3221
rect 4552 3187 5282 3197
rect 5392 3187 10514 3197
rect 10528 3187 12098 3197
rect 12112 3187 12530 3197
rect 12544 3187 16298 3197
rect 16312 3187 16490 3197
rect 16504 3187 21074 3197
rect 21088 3187 21146 3197
rect 4552 3163 9770 3173
rect 9976 3163 11714 3173
rect 11728 3163 19394 3173
rect 19408 3163 20330 3173
rect 20344 3163 24890 3173
rect 4624 3139 15002 3149
rect 21088 3139 21350 3149
rect 4672 3115 6554 3125
rect 6568 3115 13610 3125
rect 4816 3091 11402 3101
rect 11416 3091 13226 3101
rect 4840 3067 20354 3077
rect 4888 3043 4898 3053
rect 4912 3043 20282 3053
rect 4936 3019 7394 3029
rect 7408 3019 11954 3029
rect 11968 3019 20618 3029
rect 20632 3019 20858 3029
rect 20872 3019 20906 3029
rect 20920 3019 21314 3029
rect 21328 3019 23618 3029
rect 4960 2995 15458 3005
rect 5056 2971 21338 2981
rect 5080 2947 6026 2957
rect 6040 2947 26258 2957
rect 26272 2947 26522 2957
rect 5128 2923 9554 2933
rect 9568 2923 23486 2933
rect 5200 2899 9146 2909
rect 9160 2899 21482 2909
rect 5272 2875 20258 2885
rect 5320 2851 12074 2861
rect 12328 2851 20378 2861
rect 5320 2827 6890 2837
rect 6976 2827 14474 2837
rect 5416 2803 18362 2813
rect 18376 2803 22682 2813
rect 5752 2779 20714 2789
rect 22696 2779 23018 2789
rect 5920 2755 7562 2765
rect 7648 2755 23426 2765
rect 6088 2731 17834 2741
rect 6136 2707 8498 2717
rect 8512 2707 18578 2717
rect 18592 2707 24266 2717
rect 6184 2683 6410 2693
rect 6736 2683 18938 2693
rect 18952 2683 26330 2693
rect 6352 2659 6434 2669
rect 6760 2659 24818 2669
rect 6400 2635 16850 2645
rect 6448 2611 24698 2621
rect 7096 2587 17810 2597
rect 7096 2563 19178 2573
rect 19192 2563 20426 2573
rect 20440 2563 21866 2573
rect 7216 2539 9098 2549
rect 9112 2539 9386 2549
rect 9520 2539 22946 2549
rect 22960 2539 24770 2549
rect 7240 2515 7994 2525
rect 8008 2515 10394 2525
rect 10408 2515 12146 2525
rect 12160 2515 17882 2525
rect 7264 2491 16970 2501
rect 7360 2467 12554 2477
rect 12880 2467 22922 2477
rect 7360 2443 19490 2453
rect 7456 2419 14786 2429
rect 7528 2395 7586 2405
rect 7648 2395 7730 2405
rect 7744 2395 8738 2405
rect 8752 2395 10826 2405
rect 10840 2395 12362 2405
rect 12376 2395 22898 2405
rect 22912 2395 24554 2405
rect 24568 2395 26498 2405
rect 7672 2371 25058 2381
rect 7672 2347 9434 2357
rect 9616 2347 12290 2357
rect 13024 2347 21170 2357
rect 21184 2347 22370 2357
rect 22384 2347 26930 2357
rect 7888 2323 11450 2333
rect 11464 2323 14066 2333
rect 14080 2323 18698 2333
rect 18712 2323 19154 2333
rect 22384 2323 22538 2333
rect 22912 2323 23138 2333
rect 8104 2299 12842 2309
rect 12856 2299 19274 2309
rect 8128 2275 18794 2285
rect 8320 2251 8330 2261
rect 8416 2251 12386 2261
rect 13192 2251 13490 2261
rect 8464 2227 14330 2237
rect 8584 2203 21698 2213
rect 8728 2179 8786 2189
rect 8872 2179 17426 2189
rect 17440 2179 21746 2189
rect 8824 2155 18506 2165
rect 9016 2131 12338 2141
rect 13264 2131 14642 2141
rect 14656 2131 27194 2141
rect 9784 2107 16994 2117
rect 17008 2107 26666 2117
rect 10096 2083 10130 2093
rect 10144 2083 23474 2093
rect 10168 2059 10682 2069
rect 10696 2059 16634 2069
rect 16648 2059 17738 2069
rect 17752 2059 18866 2069
rect 18880 2059 24794 2069
rect 10216 2035 14450 2045
rect 16648 2035 16682 2045
rect 10288 2011 10322 2021
rect 10408 2011 18242 2021
rect 18256 2011 24170 2021
rect 10336 1987 11522 1997
rect 11608 1987 23114 1997
rect 10672 1963 27565 1973
rect 10984 1939 14762 1949
rect 27232 1939 27565 1949
rect 11032 1915 14954 1925
rect 27208 1915 27565 1925
rect 11056 1891 11690 1901
rect 11776 1891 23354 1901
rect 27112 1891 27565 1901
rect 11152 1867 11234 1877
rect 11392 1867 18962 1877
rect 18976 1867 20594 1877
rect 20608 1867 20930 1877
rect 27184 1867 27565 1877
rect 11656 1843 16946 1853
rect 20944 1843 21458 1853
rect 27160 1843 27565 1853
rect 16960 1819 17090 1829
rect 27136 1819 27565 1829
rect 26547 1790 27123 1800
rect 26547 1767 27123 1777
rect 26547 1729 27123 1754
rect 26547 1084 27123 1109
rect 12592 986 22082 996
rect 12400 962 16994 972
rect 12256 938 16250 948
rect 19096 938 23954 948
rect 11824 914 20546 924
rect 11704 890 25370 900
rect 10048 866 10850 876
rect 10864 866 23714 876
rect 8512 842 22922 852
rect 8392 818 19178 828
rect 20128 818 22178 828
rect 8224 794 15602 804
rect 15616 794 18074 804
rect 18280 794 23018 804
rect 8008 770 13754 780
rect 14224 770 25130 780
rect 7984 746 8810 756
rect 8824 746 10466 756
rect 10480 746 11906 756
rect 11920 746 14090 756
rect 14104 746 16130 756
rect 16144 746 16730 756
rect 16744 746 23354 756
rect 23368 746 26330 756
rect 7552 722 16466 732
rect 17536 722 20834 732
rect 7312 698 10754 708
rect 11104 698 11786 708
rect 12112 698 20450 708
rect 20776 698 21698 708
rect 7048 674 16706 684
rect 17176 674 19706 684
rect 19720 674 20810 684
rect 6832 650 9098 660
rect 9808 650 15842 660
rect 15856 650 22034 660
rect 6808 626 20858 636
rect 6784 602 14522 612
rect 15904 602 22154 612
rect 22984 602 23114 612
rect 6712 578 19850 588
rect 19864 578 25034 588
rect 6568 554 26306 564
rect 6496 530 16082 540
rect 16816 530 22322 540
rect 22504 530 23762 540
rect 6472 506 8978 516
rect 9712 506 10922 516
rect 10936 506 26042 516
rect 5560 482 17858 492
rect 5512 458 22538 468
rect 5488 434 6602 444
rect 6688 434 12842 444
rect 12856 434 25250 444
rect 5248 410 23210 420
rect 5032 386 7010 396
rect 7024 386 7826 396
rect 7840 386 14354 396
rect 14368 386 22298 396
rect 22312 386 22802 396
rect 22816 386 23282 396
rect 23296 386 26306 396
rect 4600 362 16370 372
rect 4504 338 12914 348
rect 13456 338 26210 348
rect 4312 314 13610 324
rect 13672 314 24002 324
rect 4216 290 17714 300
rect 4168 266 13706 276
rect 14488 266 15410 276
rect 16000 266 22202 276
rect 3880 242 4682 252
rect 4696 242 8186 252
rect 8200 242 20258 252
rect 20272 242 26354 252
rect 3496 218 13466 228
rect 13696 218 14018 228
rect 14512 218 17570 228
rect 2680 194 4562 204
rect 4744 194 19034 204
rect 19048 194 24050 204
rect 2464 170 12938 180
rect 12952 170 13778 180
rect 2392 146 14114 156
rect 26392 146 27565 156
rect 84 122 3602 132
rect 3712 122 8642 132
rect 8656 122 8858 132
rect 8872 122 11282 132
rect 11296 122 25226 132
rect 25240 122 26402 132
rect 84 98 2642 108
rect 2728 98 23642 108
rect 23656 98 25106 108
rect 26368 98 27565 108
rect 84 74 5594 84
rect 6280 74 8882 84
rect 8944 74 13802 84
rect 26344 74 27565 84
rect 84 50 2234 60
rect 2344 50 23186 60
rect 26320 50 27565 60
rect 5368 26 26378 36
rect 26416 26 27565 36
rect 9976 2 27565 12
<< m2contact >>
rect 14450 8146 14464 8160
rect 18170 8146 18184 8160
rect 18314 8146 18328 8160
rect 20546 8146 20560 8160
rect 22202 8146 22216 8160
rect 12866 8122 12880 8136
rect 25694 8122 25708 8136
rect 4106 8098 4120 8112
rect 18194 8098 18208 8112
rect 19706 8098 19720 8112
rect 27178 8098 27192 8112
rect 3266 8074 3280 8088
rect 4622 8074 4636 8088
rect 6890 8074 6904 8088
rect 10634 8074 10648 8088
rect 19946 8074 19960 8088
rect 26090 8074 26104 8088
rect 2882 8050 2896 8064
rect 22694 8050 22708 8064
rect 70 8026 84 8040
rect 8762 8026 8776 8040
rect 9122 8026 9136 8040
rect 23738 8026 23752 8040
rect 24098 8026 24112 8040
rect 24194 8026 24208 8040
rect 27019 8026 27033 8040
rect 27565 8026 27579 8040
rect 70 8002 84 8016
rect 1730 8002 1744 8016
rect 2306 8002 2320 8016
rect 27047 8002 27061 8016
rect 27098 8002 27112 8016
rect 27146 8002 27160 8016
rect 27565 8002 27579 8016
rect 70 7978 84 7992
rect 10130 7978 10144 7992
rect 10706 7978 10720 7992
rect 15194 7978 15208 7992
rect 18170 7978 18184 7992
rect 27020 7978 27034 7993
rect 27125 7978 27139 7992
rect 27565 7978 27579 7992
rect 3074 7954 3088 7968
rect 23978 7954 23992 7968
rect 27047 7954 27061 7968
rect 27565 7954 27579 7968
rect 3698 7930 3712 7944
rect 27154 7930 27168 7944
rect 27178 7930 27192 7944
rect 27565 7930 27579 7944
rect 4586 7906 4600 7920
rect 7826 7906 7840 7920
rect 8882 7906 8896 7920
rect 12182 7906 12196 7920
rect 12362 7906 12376 7920
rect 27565 7906 27579 7920
rect 12146 7882 12160 7896
rect 16658 7882 16672 7896
rect 18362 7882 18376 7896
rect 27125 7882 27139 7896
rect 27154 7882 27168 7896
rect 27565 7882 27579 7896
rect 14882 7049 14896 7063
rect 14954 7049 14968 7063
rect 23930 7049 23944 7063
rect 26138 7049 26152 7063
rect 13514 7025 13528 7039
rect 24290 7025 24304 7039
rect 13418 7001 13432 7015
rect 13706 7001 13720 7015
rect 13898 7001 13912 7015
rect 14138 7001 14152 7015
rect 14498 7001 14512 7015
rect 24122 7001 24136 7015
rect 12818 6977 12832 6991
rect 24434 6977 24448 6991
rect 11978 6953 11992 6967
rect 12842 6953 12856 6967
rect 13130 6953 13144 6967
rect 23930 6953 23944 6967
rect 11930 6929 11944 6943
rect 12386 6929 12400 6943
rect 12698 6929 12712 6943
rect 13142 6929 13156 6943
rect 13274 6929 13288 6943
rect 13970 6929 13984 6943
rect 17954 6929 17968 6943
rect 18722 6929 18736 6943
rect 11738 6905 11752 6919
rect 11786 6905 11800 6919
rect 11882 6905 11896 6919
rect 11954 6905 11968 6919
rect 12002 6905 12016 6919
rect 12890 6905 12904 6919
rect 13082 6905 13096 6919
rect 13898 6905 13912 6919
rect 17978 6905 17992 6919
rect 10418 6881 10432 6895
rect 10826 6881 10840 6895
rect 11642 6881 11656 6895
rect 16682 6881 16696 6895
rect 10202 6857 10216 6871
rect 10466 6857 10480 6871
rect 12434 6857 12448 6871
rect 20018 6857 20032 6871
rect 24986 6857 25000 6871
rect 10106 6833 10120 6847
rect 10514 6833 10528 6847
rect 11258 6833 11272 6847
rect 13754 6833 13768 6847
rect 14258 6833 14272 6847
rect 14330 6833 14344 6847
rect 14402 6833 14416 6847
rect 14474 6833 14488 6847
rect 14546 6833 14560 6847
rect 26234 6833 26248 6847
rect 10082 6809 10096 6823
rect 17162 6809 17176 6823
rect 18554 6809 18568 6823
rect 18866 6809 18880 6823
rect 9938 6785 9952 6799
rect 24314 6785 24328 6799
rect 27218 6785 27232 6799
rect 9890 6761 9904 6775
rect 11426 6761 11440 6775
rect 11594 6761 11608 6775
rect 20690 6761 20704 6775
rect 9866 6737 9880 6751
rect 14426 6737 14440 6751
rect 25010 6737 25024 6751
rect 9842 6713 9856 6727
rect 13850 6713 13864 6727
rect 22754 6713 22768 6727
rect 23258 6713 23272 6727
rect 26066 6713 26080 6727
rect 9746 6689 9760 6703
rect 15410 6689 15424 6703
rect 18554 6689 18568 6703
rect 25394 6689 25408 6703
rect 9722 6665 9736 6679
rect 10370 6665 10384 6679
rect 11834 6665 11848 6679
rect 22874 6665 22888 6679
rect 24242 6665 24256 6679
rect 9674 6641 9688 6655
rect 10562 6641 10576 6655
rect 10802 6641 10816 6655
rect 11618 6641 11632 6655
rect 11666 6641 11680 6655
rect 11714 6641 11728 6655
rect 11810 6641 11824 6655
rect 14210 6641 14224 6655
rect 18050 6641 18064 6655
rect 24146 6641 24160 6655
rect 9626 6617 9640 6631
rect 14306 6617 14320 6631
rect 14378 6617 14392 6631
rect 23570 6617 23584 6631
rect 9338 6593 9352 6607
rect 11306 6593 11320 6607
rect 14882 6593 14896 6607
rect 17234 6593 17248 6607
rect 23258 6593 23272 6607
rect 9074 6569 9088 6583
rect 15602 6569 15616 6583
rect 9050 6545 9064 6559
rect 21050 6545 21064 6559
rect 27050 6545 27064 6559
rect 8954 6521 8968 6535
rect 11090 6521 11104 6535
rect 12818 6521 12832 6535
rect 20378 6521 20392 6535
rect 23306 6521 23320 6535
rect 8930 6497 8944 6511
rect 10298 6497 10312 6511
rect 12482 6497 12496 6511
rect 13730 6497 13744 6511
rect 18482 6497 18496 6511
rect 18842 6497 18856 6511
rect 21026 6497 21040 6511
rect 23330 6497 23344 6511
rect 8834 6473 8848 6487
rect 23858 6473 23872 6487
rect 8738 6449 8752 6463
rect 21530 6449 21544 6463
rect 8666 6425 8680 6439
rect 16418 6425 16432 6439
rect 26354 6425 26368 6439
rect 26594 6425 26608 6439
rect 8642 6401 8656 6415
rect 26354 6401 26368 6415
rect 27170 6401 27184 6415
rect 8546 6377 8560 6391
rect 14690 6377 14704 6391
rect 14834 6377 14848 6391
rect 16778 6377 16792 6391
rect 20138 6377 20152 6391
rect 24530 6377 24544 6391
rect 8522 6353 8536 6367
rect 25346 6353 25360 6367
rect 8186 6329 8200 6343
rect 11258 6329 11272 6343
rect 20210 6329 20224 6343
rect 21554 6329 21568 6343
rect 21986 6329 22000 6343
rect 25634 6329 25648 6343
rect 8066 6305 8080 6319
rect 10586 6305 10600 6319
rect 10730 6305 10744 6319
rect 21098 6305 21112 6319
rect 7778 6281 7792 6295
rect 19826 6281 19840 6295
rect 20090 6281 20104 6295
rect 20354 6281 20368 6295
rect 7610 6257 7624 6271
rect 14834 6257 14848 6271
rect 15722 6257 15736 6271
rect 15806 6257 15820 6271
rect 16538 6257 16552 6271
rect 16658 6257 16672 6271
rect 19874 6257 19888 6271
rect 19922 6257 19936 6271
rect 19994 6257 20008 6271
rect 20282 6257 20296 6271
rect 21434 6257 21448 6271
rect 21698 6257 21712 6271
rect 7586 6233 7600 6247
rect 11306 6233 11320 6247
rect 11498 6233 11512 6247
rect 14906 6233 14920 6247
rect 20114 6233 20128 6247
rect 25058 6233 25072 6247
rect 7418 6209 7432 6223
rect 21434 6209 21448 6223
rect 7394 6185 7408 6199
rect 17642 6185 17656 6199
rect 19778 6185 19792 6199
rect 21218 6185 21232 6199
rect 21842 6185 21856 6199
rect 21878 6185 21892 6199
rect 7298 6161 7312 6175
rect 10322 6161 10336 6175
rect 23594 6161 23608 6175
rect 7202 6137 7216 6151
rect 7706 6137 7720 6151
rect 14810 6137 14824 6151
rect 15722 6137 15736 6151
rect 18290 6137 18304 6151
rect 21650 6137 21664 6151
rect 21842 6137 21856 6151
rect 7034 6113 7048 6127
rect 11042 6113 11056 6127
rect 11114 6113 11128 6127
rect 14306 6113 14320 6127
rect 23786 6113 23800 6127
rect 6986 6089 7000 6103
rect 18410 6089 18424 6103
rect 19634 6089 19648 6103
rect 20666 6089 20680 6103
rect 6770 6065 6784 6079
rect 7778 6065 7792 6079
rect 11234 6065 11248 6079
rect 11738 6065 11752 6079
rect 13658 6065 13672 6079
rect 13778 6065 13792 6079
rect 14114 6065 14128 6079
rect 17090 6065 17104 6079
rect 22130 6065 22144 6079
rect 22646 6065 22660 6079
rect 6506 6041 6520 6055
rect 6530 6041 6544 6055
rect 6578 6041 6592 6055
rect 20954 6041 20968 6055
rect 6314 6017 6328 6031
rect 12194 6017 12208 6031
rect 12266 6017 12280 6031
rect 13286 6017 13300 6031
rect 13322 6017 13336 6031
rect 13610 6017 13624 6031
rect 14066 6017 14080 6031
rect 20522 6017 20536 6031
rect 6290 5993 6304 6007
rect 11138 5993 11152 6007
rect 11210 5993 11224 6007
rect 11282 5993 11296 6007
rect 11354 5993 11368 6007
rect 23210 5993 23224 6007
rect 6050 5969 6064 5983
rect 10226 5969 10240 5983
rect 22322 5969 22336 5983
rect 5954 5945 5968 5959
rect 22586 5945 22600 5959
rect 25826 5945 25840 5959
rect 5858 5921 5872 5935
rect 26738 5921 26752 5935
rect 5786 5897 5800 5911
rect 6218 5897 6232 5911
rect 9890 5897 9904 5911
rect 11666 5897 11680 5911
rect 20450 5897 20464 5911
rect 24458 5897 24472 5911
rect 25154 5897 25168 5911
rect 5714 5873 5728 5887
rect 13586 5873 13600 5887
rect 13826 5873 13840 5887
rect 14570 5873 14584 5887
rect 16394 5873 16408 5887
rect 19970 5873 19984 5887
rect 20042 5873 20056 5887
rect 26474 5873 26488 5887
rect 5618 5849 5632 5863
rect 13538 5849 13552 5863
rect 13634 5849 13648 5863
rect 17042 5849 17056 5863
rect 17594 5849 17608 5863
rect 23138 5849 23152 5863
rect 25106 5849 25120 5863
rect 5666 5825 5680 5839
rect 21914 5825 21928 5839
rect 23450 5825 23464 5839
rect 25202 5825 25216 5839
rect 5498 5801 5512 5815
rect 11858 5801 11872 5815
rect 12458 5801 12472 5815
rect 12986 5801 13000 5815
rect 16538 5801 16552 5815
rect 16802 5801 16816 5815
rect 19562 5801 19576 5815
rect 24458 5801 24472 5815
rect 5450 5777 5464 5791
rect 8642 5777 8656 5791
rect 8978 5777 8992 5791
rect 9290 5777 9304 5791
rect 16514 5777 16528 5791
rect 17378 5777 17392 5791
rect 25778 5777 25792 5791
rect 5402 5753 5416 5767
rect 7586 5753 7600 5767
rect 20594 5753 20608 5767
rect 5354 5729 5368 5743
rect 10274 5729 10288 5743
rect 15746 5729 15760 5743
rect 16418 5729 16432 5743
rect 26690 5729 26704 5743
rect 5258 5705 5272 5719
rect 24602 5705 24616 5719
rect 5210 5681 5224 5695
rect 14522 5681 14536 5695
rect 16322 5681 16336 5695
rect 16370 5681 16384 5695
rect 17354 5681 17368 5695
rect 20210 5681 20224 5695
rect 26186 5681 26200 5695
rect 26330 5681 26344 5695
rect 5186 5657 5200 5671
rect 5834 5657 5848 5671
rect 6818 5657 6832 5671
rect 6914 5657 6928 5671
rect 26186 5657 26200 5671
rect 5162 5633 5176 5647
rect 8330 5633 8344 5647
rect 21266 5633 21280 5647
rect 5090 5609 5104 5623
rect 8570 5609 8584 5623
rect 13490 5609 13504 5623
rect 24242 5609 24256 5623
rect 25466 5609 25480 5623
rect 4994 5585 5008 5599
rect 8402 5585 8416 5599
rect 8450 5585 8464 5599
rect 15050 5585 15064 5599
rect 15578 5585 15592 5599
rect 22730 5585 22744 5599
rect 4970 5561 4984 5575
rect 10634 5561 10648 5575
rect 19322 5561 19336 5575
rect 19418 5561 19432 5575
rect 24578 5561 24592 5575
rect 4874 5537 4888 5551
rect 8306 5537 8320 5551
rect 10874 5537 10888 5551
rect 13922 5537 13936 5551
rect 18386 5537 18400 5551
rect 22706 5537 22720 5551
rect 24362 5537 24376 5551
rect 27122 5537 27136 5551
rect 4850 5513 4864 5527
rect 9818 5513 9832 5527
rect 10850 5513 10864 5527
rect 11186 5513 11200 5527
rect 12938 5513 12952 5527
rect 13514 5513 13528 5527
rect 14078 5513 14092 5527
rect 17618 5513 17632 5527
rect 19298 5513 19312 5527
rect 20570 5513 20584 5527
rect 21194 5513 21208 5527
rect 22490 5513 22504 5527
rect 24338 5513 24352 5527
rect 4658 5489 4672 5503
rect 9650 5489 9664 5503
rect 25730 5489 25744 5503
rect 26450 5489 26464 5503
rect 26666 5489 26680 5503
rect 4586 5465 4600 5479
rect 7538 5465 7552 5479
rect 21938 5465 21952 5479
rect 26450 5465 26464 5479
rect 4370 5441 4384 5455
rect 26018 5441 26032 5455
rect 4298 5417 4312 5431
rect 12674 5417 12688 5431
rect 12914 5417 12928 5431
rect 13538 5417 13552 5431
rect 18002 5417 18016 5431
rect 18890 5417 18904 5431
rect 21458 5417 21472 5431
rect 24074 5417 24088 5431
rect 4274 5393 4288 5407
rect 16442 5393 16456 5407
rect 16826 5393 16840 5407
rect 16874 5393 16888 5407
rect 16922 5393 16936 5407
rect 17066 5393 17080 5407
rect 17282 5393 17296 5407
rect 19034 5393 19048 5407
rect 19226 5393 19240 5407
rect 20714 5393 20728 5407
rect 20882 5393 20896 5407
rect 21674 5393 21688 5407
rect 4250 5369 4264 5383
rect 4490 5369 4504 5383
rect 9938 5369 9952 5383
rect 11210 5369 11224 5383
rect 12962 5369 12976 5383
rect 14234 5369 14248 5383
rect 18818 5369 18832 5383
rect 18890 5369 18904 5383
rect 21122 5369 21136 5383
rect 25010 5369 25024 5383
rect 4058 5345 4072 5359
rect 10658 5345 10672 5359
rect 18218 5345 18232 5359
rect 19130 5345 19144 5359
rect 23690 5345 23704 5359
rect 3986 5321 4000 5335
rect 7322 5321 7336 5335
rect 8618 5321 8632 5335
rect 11762 5321 11776 5335
rect 11882 5321 11896 5335
rect 12794 5321 12808 5335
rect 14402 5321 14416 5335
rect 22250 5321 22264 5335
rect 22466 5321 22480 5335
rect 3962 5297 3976 5311
rect 6794 5297 6808 5311
rect 12770 5297 12784 5311
rect 20642 5297 20656 5311
rect 21818 5297 21832 5311
rect 23522 5297 23536 5311
rect 3890 5273 3904 5287
rect 6146 5273 6160 5287
rect 10058 5273 10072 5287
rect 13034 5273 13048 5287
rect 13346 5273 13360 5287
rect 16706 5273 16720 5287
rect 20090 5273 20104 5287
rect 20462 5273 20476 5287
rect 20738 5273 20752 5287
rect 22346 5273 22360 5287
rect 25730 5273 25744 5287
rect 25970 5273 25984 5287
rect 3746 5249 3760 5263
rect 14594 5249 14608 5263
rect 14738 5249 14752 5263
rect 22994 5249 23008 5263
rect 3650 5225 3664 5239
rect 10610 5225 10624 5239
rect 20978 5225 20992 5239
rect 3554 5201 3568 5215
rect 6650 5201 6664 5215
rect 23006 5201 23020 5215
rect 3530 5177 3544 5191
rect 22850 5177 22864 5191
rect 3482 5153 3496 5167
rect 4778 5153 4792 5167
rect 11354 5153 11368 5167
rect 11402 5153 11416 5167
rect 12578 5153 12592 5167
rect 12650 5153 12664 5167
rect 23306 5153 23320 5167
rect 23402 5153 23416 5167
rect 23486 5153 23500 5167
rect 3434 5129 3448 5143
rect 10922 5129 10936 5143
rect 10970 5129 10984 5143
rect 23834 5129 23848 5143
rect 3362 5105 3376 5119
rect 26546 5105 26560 5119
rect 3338 5081 3352 5095
rect 4706 5081 4720 5095
rect 7850 5081 7864 5095
rect 8162 5081 8176 5095
rect 14282 5081 14296 5095
rect 16154 5081 16168 5095
rect 16826 5081 16840 5095
rect 18626 5081 18640 5095
rect 21290 5081 21304 5095
rect 22274 5081 22288 5095
rect 23402 5081 23416 5095
rect 27146 5081 27160 5095
rect 3314 5057 3328 5071
rect 7466 5057 7480 5071
rect 7922 5057 7936 5071
rect 8042 5057 8056 5071
rect 10586 5057 10600 5071
rect 13682 5057 13696 5071
rect 18818 5057 18832 5071
rect 19682 5057 19696 5071
rect 19754 5057 19768 5071
rect 22418 5057 22432 5071
rect 3242 5033 3256 5047
rect 21962 5033 21976 5047
rect 23234 5033 23248 5047
rect 3218 5009 3232 5023
rect 3794 5009 3808 5023
rect 3866 5009 3880 5023
rect 10346 5009 10360 5023
rect 21290 5009 21304 5023
rect 26402 5009 26416 5023
rect 3122 4985 3136 4999
rect 17762 4985 17776 4999
rect 18170 4985 18184 4999
rect 18242 4985 18256 4999
rect 18314 4985 18328 4999
rect 18338 4985 18352 4999
rect 19058 4985 19072 4999
rect 21002 4985 21016 4999
rect 21314 4985 21328 4999
rect 26762 4985 26776 4999
rect 3098 4961 3112 4975
rect 9986 4961 10000 4975
rect 10058 4961 10072 4975
rect 11786 4961 11800 4975
rect 20498 4961 20512 4975
rect 20834 4961 20848 4975
rect 21578 4961 21592 4975
rect 25970 4961 25984 4975
rect 3002 4937 3016 4951
rect 18770 4937 18784 4951
rect 19610 4937 19624 4951
rect 19658 4937 19672 4951
rect 22034 4937 22048 4951
rect 22202 4937 22216 4951
rect 25154 4937 25168 4951
rect 2954 4913 2968 4927
rect 7802 4913 7816 4927
rect 8426 4913 8440 4927
rect 25250 4913 25264 4927
rect 2906 4889 2920 4903
rect 14786 4889 14800 4903
rect 15554 4889 15568 4903
rect 21350 4889 21364 4903
rect 22154 4889 22168 4903
rect 22466 4889 22480 4903
rect 2810 4865 2824 4879
rect 16610 4865 16624 4879
rect 16898 4865 16912 4879
rect 16970 4865 16984 4879
rect 17114 4865 17128 4879
rect 18458 4865 18472 4879
rect 18986 4865 19000 4879
rect 23186 4865 23200 4879
rect 2762 4841 2776 4855
rect 7682 4841 7696 4855
rect 7754 4841 7768 4855
rect 8234 4841 8248 4855
rect 8258 4841 8272 4855
rect 23714 4841 23728 4855
rect 23906 4841 23920 4855
rect 2690 4817 2704 4831
rect 10778 4817 10792 4831
rect 13418 4817 13432 4831
rect 16754 4817 16768 4831
rect 22562 4817 22576 4831
rect 2666 4793 2680 4807
rect 8786 4793 8800 4807
rect 14162 4793 14176 4807
rect 17474 4793 17488 4807
rect 20162 4793 20176 4807
rect 24026 4793 24040 4807
rect 2618 4769 2632 4783
rect 9410 4769 9424 4783
rect 9458 4769 9472 4783
rect 15806 4769 15820 4783
rect 16274 4769 16288 4783
rect 16850 4769 16864 4783
rect 19946 4769 19960 4783
rect 22538 4769 22552 4783
rect 2570 4745 2584 4759
rect 10442 4745 10456 4759
rect 10490 4745 10504 4759
rect 25682 4745 25696 4759
rect 2522 4721 2536 4735
rect 20402 4721 20416 4735
rect 20762 4721 20776 4735
rect 23162 4721 23176 4735
rect 2498 4697 2512 4711
rect 10802 4697 10816 4711
rect 22514 4697 22528 4711
rect 2474 4673 2488 4687
rect 6266 4673 6280 4687
rect 21386 4673 21400 4687
rect 24050 4673 24064 4687
rect 25130 4673 25144 4687
rect 2402 4649 2416 4663
rect 18458 4649 18472 4663
rect 23378 4649 23392 4663
rect 2354 4625 2368 4639
rect 13010 4625 13024 4639
rect 13058 4625 13072 4639
rect 13442 4625 13456 4639
rect 13562 4625 13576 4639
rect 26402 4625 26416 4639
rect 2282 4601 2296 4615
rect 3674 4601 3688 4615
rect 9194 4601 9208 4615
rect 10634 4601 10648 4615
rect 10706 4601 10720 4615
rect 26570 4601 26584 4615
rect 2234 4577 2248 4591
rect 3194 4577 3208 4591
rect 18314 4577 18328 4591
rect 18650 4577 18664 4591
rect 22430 4577 22444 4591
rect 2234 4553 2248 4567
rect 25322 4553 25336 4567
rect 2210 4529 2224 4543
rect 7730 4529 7744 4543
rect 11426 4529 11440 4543
rect 23954 4529 23968 4543
rect 2138 4505 2152 4519
rect 3266 4505 3280 4519
rect 5930 4505 5944 4519
rect 7154 4505 7168 4519
rect 15866 4505 15880 4519
rect 16034 4505 16048 4519
rect 16922 4505 16936 4519
rect 18434 4505 18448 4519
rect 22058 4505 22072 4519
rect 23090 4505 23104 4519
rect 23546 4505 23560 4519
rect 2114 4481 2128 4495
rect 24482 4481 24496 4495
rect 24866 4481 24880 4495
rect 24890 4481 24904 4495
rect 1946 4457 1960 4471
rect 3410 4457 3424 4471
rect 18194 4457 18208 4471
rect 18506 4457 18520 4471
rect 26090 4457 26104 4471
rect 1898 4433 1912 4447
rect 4826 4433 4840 4447
rect 5354 4433 5368 4447
rect 8282 4433 8296 4447
rect 13202 4433 13216 4447
rect 13874 4433 13888 4447
rect 14018 4433 14032 4447
rect 18914 4433 18928 4447
rect 22010 4433 22024 4447
rect 26594 4433 26608 4447
rect 1874 4409 1888 4423
rect 13178 4409 13192 4423
rect 24386 4409 24400 4423
rect 1826 4385 1840 4399
rect 8714 4385 8728 4399
rect 8762 4385 8776 4399
rect 19466 4385 19480 4399
rect 20066 4385 20080 4399
rect 22802 4385 22816 4399
rect 25874 4385 25888 4399
rect 1802 4361 1816 4375
rect 21602 4361 21616 4375
rect 22082 4361 22096 4375
rect 22610 4361 22624 4375
rect 22826 4361 22840 4375
rect 25226 4361 25240 4375
rect 1682 4337 1696 4351
rect 17186 4337 17200 4351
rect 17762 4337 17776 4351
rect 18338 4337 18352 4351
rect 18410 4337 18424 4351
rect 18722 4337 18736 4351
rect 18842 4337 18856 4351
rect 27098 4337 27112 4351
rect 1658 4313 1672 4327
rect 4514 4313 4528 4327
rect 11330 4313 11344 4327
rect 16610 4313 16624 4327
rect 16754 4313 16768 4327
rect 16778 4313 16792 4327
rect 17042 4313 17056 4327
rect 19514 4313 19528 4327
rect 20642 4313 20656 4327
rect 20666 4313 20680 4327
rect 21194 4313 21208 4327
rect 21554 4313 21568 4327
rect 21626 4313 21640 4327
rect 26786 4313 26800 4327
rect 1610 4289 1624 4303
rect 2306 4289 2320 4303
rect 6650 4289 6664 4303
rect 8426 4289 8440 4303
rect 11930 4289 11944 4303
rect 12770 4289 12784 4303
rect 14258 4289 14272 4303
rect 19370 4289 19384 4303
rect 21266 4289 21280 4303
rect 21650 4289 21664 4303
rect 22274 4289 22288 4303
rect 22322 4289 22336 4303
rect 22610 4289 22624 4303
rect 22646 4289 22660 4303
rect 22826 4289 22840 4303
rect 23006 4289 23020 4303
rect 23522 4289 23536 4303
rect 23570 4289 23584 4303
rect 70 4265 84 4279
rect 21770 4265 21784 4279
rect 70 4241 84 4255
rect 22226 4241 22240 4255
rect 70 4217 84 4231
rect 1994 4217 2008 4231
rect 2042 4217 2056 4231
rect 19298 4217 19312 4231
rect 70 4193 84 4207
rect 14738 4193 14752 4207
rect 14930 4193 14944 4207
rect 23666 4193 23680 4207
rect 1730 4169 1744 4183
rect 6506 4169 6520 4183
rect 6674 4169 6688 4183
rect 14186 4169 14200 4183
rect 15650 4169 15664 4183
rect 15794 4169 15808 4183
rect 19202 4169 19216 4183
rect 25922 4169 25936 4183
rect 1778 4145 1792 4159
rect 22634 4145 22648 4159
rect 2042 4121 2056 4135
rect 4442 4121 4456 4135
rect 7514 4121 7528 4135
rect 16058 4121 16072 4135
rect 16730 4121 16744 4135
rect 23090 4121 23104 4135
rect 23690 4121 23704 4135
rect 26162 4121 26176 4135
rect 2090 4097 2104 4111
rect 5690 4097 5704 4111
rect 7274 4097 7288 4111
rect 9866 4097 9880 4111
rect 12146 4097 12160 4111
rect 12698 4097 12712 4111
rect 14354 4097 14368 4111
rect 15962 4097 15976 4111
rect 21506 4097 21520 4111
rect 23066 4097 23080 4111
rect 26882 4097 26896 4111
rect 2162 4073 2176 4087
rect 14690 4073 14704 4087
rect 16322 4073 16336 4087
rect 25538 4073 25552 4087
rect 27098 4073 27112 4087
rect 2258 4049 2272 4063
rect 14618 4049 14632 4063
rect 14714 4049 14728 4063
rect 17522 4049 17536 4063
rect 17906 4049 17920 4063
rect 18362 4049 18376 4063
rect 19010 4049 19024 4063
rect 21794 4049 21808 4063
rect 23066 4049 23080 4063
rect 23138 4049 23152 4063
rect 2282 4025 2296 4039
rect 6866 4025 6880 4039
rect 22298 4025 22312 4039
rect 22394 4025 22408 4039
rect 2402 4001 2416 4015
rect 7322 4001 7336 4015
rect 8210 4001 8224 4015
rect 11018 4001 11032 4015
rect 13802 4001 13816 4015
rect 14858 4001 14872 4015
rect 19994 4001 20008 4015
rect 20954 4001 20968 4015
rect 22706 4001 22720 4015
rect 24098 4001 24112 4015
rect 26306 4001 26320 4015
rect 26642 4001 26656 4015
rect 2498 3977 2512 3991
rect 2594 3977 2608 3991
rect 5282 3977 5296 3991
rect 6578 3977 6592 3991
rect 6986 3977 7000 3991
rect 8834 3977 8848 3991
rect 9674 3977 9688 3991
rect 11162 3977 11176 3991
rect 16130 3977 16144 3991
rect 26498 3977 26512 3991
rect 26978 3977 26992 3991
rect 2522 3953 2536 3967
rect 4610 3953 4624 3967
rect 4994 3953 5008 3967
rect 7058 3953 7072 3967
rect 7130 3953 7144 3967
rect 7874 3953 7888 3967
rect 8954 3953 8968 3967
rect 12002 3953 12016 3967
rect 12122 3953 12136 3967
rect 12242 3953 12256 3967
rect 17018 3953 17032 3967
rect 22106 3953 22120 3967
rect 22970 3953 22984 3967
rect 24866 3953 24880 3967
rect 25946 3953 25960 3967
rect 27002 3953 27016 3967
rect 2570 3929 2584 3943
rect 7610 3929 7624 3943
rect 9506 3929 9520 3943
rect 10034 3929 10048 3943
rect 10754 3929 10768 3943
rect 15938 3929 15952 3943
rect 16898 3929 16912 3943
rect 18122 3929 18136 3943
rect 20546 3929 20560 3943
rect 22394 3929 22408 3943
rect 22430 3929 22444 3943
rect 2618 3905 2632 3919
rect 3578 3905 3592 3919
rect 5570 3905 5584 3919
rect 13142 3905 13156 3919
rect 23810 3905 23824 3919
rect 25298 3905 25312 3919
rect 2714 3881 2728 3895
rect 12602 3881 12616 3895
rect 12722 3881 12736 3895
rect 17138 3881 17152 3895
rect 2762 3857 2776 3871
rect 2882 3857 2896 3871
rect 2930 3857 2944 3871
rect 6842 3857 6856 3871
rect 6938 3857 6952 3871
rect 13370 3857 13384 3871
rect 13562 3857 13576 3871
rect 19898 3857 19912 3871
rect 3050 3833 3064 3847
rect 10418 3833 10432 3847
rect 10538 3833 10552 3847
rect 24194 3833 24208 3847
rect 3074 3809 3088 3823
rect 3626 3809 3640 3823
rect 3674 3809 3688 3823
rect 16874 3809 16888 3823
rect 18602 3809 18616 3823
rect 19874 3809 19888 3823
rect 24914 3809 24928 3823
rect 25658 3809 25672 3823
rect 3170 3785 3184 3799
rect 13058 3785 13072 3799
rect 13106 3785 13120 3799
rect 14138 3785 14152 3799
rect 21878 3785 21892 3799
rect 23138 3785 23152 3799
rect 3314 3761 3328 3775
rect 6122 3761 6136 3775
rect 7898 3761 7912 3775
rect 9530 3761 9544 3775
rect 10946 3761 10960 3775
rect 11978 3761 11992 3775
rect 18530 3761 18544 3775
rect 25754 3761 25768 3775
rect 3458 3737 3472 3751
rect 3842 3737 3856 3751
rect 5810 3737 5824 3751
rect 7130 3737 7144 3751
rect 22778 3737 22792 3751
rect 26858 3737 26872 3751
rect 3530 3713 3544 3727
rect 19082 3713 19096 3727
rect 19898 3713 19912 3727
rect 19970 3713 19984 3727
rect 3602 3689 3616 3703
rect 21722 3689 21736 3703
rect 3746 3665 3760 3679
rect 19130 3665 19144 3679
rect 20186 3665 20200 3679
rect 21050 3665 21064 3679
rect 3794 3641 3808 3655
rect 4178 3641 4192 3655
rect 11906 3641 11920 3655
rect 12170 3641 12184 3655
rect 12410 3641 12424 3655
rect 15770 3641 15784 3655
rect 16442 3641 16456 3655
rect 18746 3641 18760 3655
rect 21146 3641 21160 3655
rect 25610 3641 25624 3655
rect 26282 3641 26296 3655
rect 3818 3617 3832 3631
rect 5138 3617 5152 3631
rect 6362 3617 6376 3631
rect 7490 3617 7504 3631
rect 7946 3617 7960 3631
rect 9842 3617 9856 3631
rect 10994 3617 11008 3631
rect 11546 3617 11560 3631
rect 12746 3617 12760 3631
rect 17066 3617 17080 3631
rect 17498 3617 17512 3631
rect 17570 3617 17584 3631
rect 20810 3617 20824 3631
rect 21242 3617 21256 3631
rect 22010 3617 22024 3631
rect 25778 3617 25792 3631
rect 26210 3617 26224 3631
rect 26282 3617 26296 3631
rect 26474 3617 26488 3631
rect 3890 3593 3904 3607
rect 4082 3593 4096 3607
rect 4178 3593 4192 3607
rect 13466 3593 13480 3607
rect 18170 3593 18184 3607
rect 19922 3593 19936 3607
rect 23594 3593 23608 3607
rect 3914 3569 3928 3583
rect 22994 3569 23008 3583
rect 3938 3545 3952 3559
rect 12506 3545 12520 3559
rect 13394 3545 13408 3559
rect 23162 3545 23176 3559
rect 3962 3521 3976 3535
rect 11474 3521 11488 3535
rect 11546 3521 11560 3535
rect 13706 3521 13720 3535
rect 16562 3521 16576 3535
rect 23018 3521 23032 3535
rect 3986 3497 4000 3511
rect 23642 3497 23656 3511
rect 4010 3473 4024 3487
rect 9746 3473 9760 3487
rect 9962 3473 9976 3487
rect 12050 3473 12064 3487
rect 14666 3473 14680 3487
rect 16346 3473 16360 3487
rect 26378 3473 26392 3487
rect 4034 3449 4048 3463
rect 9266 3449 9280 3463
rect 9986 3449 10000 3463
rect 12218 3449 12232 3463
rect 12434 3449 12448 3463
rect 16586 3449 16600 3463
rect 18746 3449 18760 3463
rect 19034 3449 19048 3463
rect 20186 3449 20200 3463
rect 20462 3449 20476 3463
rect 4082 3425 4096 3439
rect 4154 3425 4168 3439
rect 4202 3425 4216 3439
rect 12626 3425 12640 3439
rect 12794 3425 12808 3439
rect 16658 3425 16672 3439
rect 4250 3401 4264 3415
rect 13442 3401 13456 3415
rect 18674 3401 18688 3415
rect 4274 3377 4288 3391
rect 6530 3377 6544 3391
rect 7418 3377 7432 3391
rect 8354 3377 8368 3391
rect 10178 3377 10192 3391
rect 11282 3377 11296 3391
rect 13994 3377 14008 3391
rect 26426 3377 26440 3391
rect 4346 3353 4360 3367
rect 6362 3353 6376 3367
rect 6410 3353 6424 3367
rect 6434 3353 6448 3367
rect 6482 3353 6496 3367
rect 8186 3353 8200 3367
rect 12890 3353 12904 3367
rect 14042 3353 14056 3367
rect 14162 3353 14176 3367
rect 14210 3353 14224 3367
rect 14354 3353 14368 3367
rect 14426 3353 14440 3367
rect 14570 3353 14584 3367
rect 26810 3353 26824 3367
rect 4346 3329 4360 3343
rect 12026 3329 12040 3343
rect 19538 3329 19552 3343
rect 4370 3305 4384 3319
rect 6002 3305 6016 3319
rect 6338 3305 6352 3319
rect 12290 3305 12304 3319
rect 13322 3305 13336 3319
rect 16082 3305 16096 3319
rect 20306 3305 20320 3319
rect 20498 3305 20512 3319
rect 21410 3305 21424 3319
rect 23042 3305 23056 3319
rect 26618 3305 26632 3319
rect 4394 3281 4408 3295
rect 12674 3281 12688 3295
rect 24650 3281 24664 3295
rect 4418 3257 4432 3271
rect 12122 3257 12136 3271
rect 12170 3257 12184 3271
rect 12362 3257 12376 3271
rect 12626 3257 12640 3271
rect 12866 3257 12880 3271
rect 12962 3257 12976 3271
rect 13286 3257 13300 3271
rect 13634 3257 13648 3271
rect 13946 3257 13960 3271
rect 13994 3257 14008 3271
rect 14078 3257 14092 3271
rect 20306 3257 20320 3271
rect 20570 3257 20584 3271
rect 4466 3233 4480 3247
rect 22418 3233 22432 3247
rect 4466 3209 4480 3223
rect 4754 3209 4768 3223
rect 7250 3209 7264 3223
rect 10298 3209 10312 3223
rect 11474 3209 11488 3223
rect 12554 3209 12568 3223
rect 20234 3209 20248 3223
rect 24170 3209 24184 3223
rect 25202 3209 25216 3223
rect 4538 3185 4552 3199
rect 5282 3185 5296 3199
rect 5378 3185 5392 3199
rect 10514 3185 10528 3199
rect 12098 3185 12112 3199
rect 12530 3185 12544 3199
rect 16298 3185 16312 3199
rect 16490 3185 16504 3199
rect 21074 3185 21088 3199
rect 21146 3185 21160 3199
rect 4538 3161 4552 3175
rect 9770 3161 9784 3175
rect 9962 3161 9976 3175
rect 11714 3161 11728 3175
rect 19394 3161 19408 3175
rect 20330 3161 20344 3175
rect 24890 3161 24904 3175
rect 4610 3137 4624 3151
rect 15002 3137 15016 3151
rect 21074 3137 21088 3151
rect 21350 3137 21364 3151
rect 4658 3113 4672 3127
rect 6554 3113 6568 3127
rect 13610 3113 13624 3127
rect 4802 3089 4816 3103
rect 11402 3089 11416 3103
rect 13226 3089 13240 3103
rect 4826 3065 4840 3079
rect 20354 3065 20368 3079
rect 4874 3041 4888 3055
rect 4898 3041 4912 3055
rect 20282 3041 20296 3055
rect 4922 3017 4936 3031
rect 7394 3017 7408 3031
rect 11954 3017 11968 3031
rect 20618 3017 20632 3031
rect 20858 3017 20872 3031
rect 20906 3017 20920 3031
rect 21314 3017 21328 3031
rect 23618 3017 23632 3031
rect 4946 2993 4960 3007
rect 15458 2993 15472 3007
rect 5042 2969 5056 2983
rect 21338 2969 21352 2983
rect 5066 2945 5080 2959
rect 6026 2945 6040 2959
rect 26258 2945 26272 2959
rect 26522 2945 26536 2959
rect 5114 2921 5128 2935
rect 9554 2921 9568 2935
rect 23486 2921 23500 2935
rect 5186 2897 5200 2911
rect 9146 2897 9160 2911
rect 21482 2897 21496 2911
rect 5258 2873 5272 2887
rect 20258 2873 20272 2887
rect 5306 2849 5320 2863
rect 12074 2849 12088 2863
rect 12314 2849 12328 2863
rect 20378 2849 20392 2863
rect 5306 2825 5320 2839
rect 6890 2825 6904 2839
rect 6962 2825 6976 2839
rect 14474 2825 14488 2839
rect 5402 2801 5416 2815
rect 18362 2801 18376 2815
rect 22682 2801 22696 2815
rect 5738 2777 5752 2791
rect 20714 2777 20728 2791
rect 22682 2777 22696 2791
rect 23018 2777 23032 2791
rect 5906 2753 5920 2767
rect 7562 2753 7576 2767
rect 7634 2753 7648 2767
rect 23426 2753 23440 2767
rect 6074 2729 6088 2743
rect 17834 2729 17848 2743
rect 6122 2705 6136 2719
rect 8498 2705 8512 2719
rect 18578 2705 18592 2719
rect 24266 2705 24280 2719
rect 6170 2681 6184 2695
rect 6410 2681 6424 2695
rect 6722 2681 6736 2695
rect 18938 2681 18952 2695
rect 26330 2681 26344 2695
rect 6338 2657 6352 2671
rect 6434 2657 6448 2671
rect 6746 2657 6760 2671
rect 24818 2657 24832 2671
rect 6386 2633 6400 2647
rect 16850 2633 16864 2647
rect 6434 2609 6448 2623
rect 24698 2609 24712 2623
rect 7082 2585 7096 2599
rect 17810 2585 17824 2599
rect 7082 2561 7096 2575
rect 19178 2561 19192 2575
rect 20426 2561 20440 2575
rect 21866 2561 21880 2575
rect 7202 2537 7216 2551
rect 9098 2537 9112 2551
rect 9386 2537 9400 2551
rect 9506 2537 9520 2551
rect 22946 2537 22960 2551
rect 24770 2537 24784 2551
rect 7226 2513 7240 2527
rect 7994 2513 8008 2527
rect 10394 2513 10408 2527
rect 12146 2513 12160 2527
rect 17882 2513 17896 2527
rect 7250 2489 7264 2503
rect 16970 2489 16984 2503
rect 7346 2465 7360 2479
rect 12554 2465 12568 2479
rect 12866 2465 12880 2479
rect 22922 2465 22936 2479
rect 7346 2441 7360 2455
rect 19490 2441 19504 2455
rect 7442 2417 7456 2431
rect 14786 2417 14800 2431
rect 7514 2393 7528 2407
rect 7586 2393 7600 2407
rect 7634 2393 7648 2407
rect 7730 2393 7744 2407
rect 8738 2393 8752 2407
rect 10826 2393 10840 2407
rect 12362 2393 12376 2407
rect 22898 2393 22912 2407
rect 24554 2393 24568 2407
rect 26498 2393 26512 2407
rect 7658 2369 7672 2383
rect 25058 2369 25072 2383
rect 7658 2345 7672 2359
rect 9434 2345 9448 2359
rect 9602 2345 9616 2359
rect 12290 2345 12304 2359
rect 13010 2345 13024 2359
rect 21170 2345 21184 2359
rect 22370 2345 22384 2359
rect 26930 2345 26944 2359
rect 7874 2321 7888 2335
rect 11450 2321 11464 2335
rect 14066 2321 14080 2335
rect 18698 2321 18712 2335
rect 19154 2321 19168 2335
rect 22370 2321 22384 2335
rect 22538 2321 22552 2335
rect 22898 2321 22912 2335
rect 23138 2321 23152 2335
rect 8090 2297 8104 2311
rect 12842 2297 12856 2311
rect 19274 2297 19288 2311
rect 8114 2273 8128 2287
rect 18794 2273 18808 2287
rect 8306 2249 8320 2263
rect 8330 2249 8344 2263
rect 8402 2249 8416 2263
rect 12386 2249 12400 2263
rect 13178 2249 13192 2263
rect 13490 2249 13504 2263
rect 8450 2225 8464 2239
rect 14330 2225 14344 2239
rect 8570 2201 8584 2215
rect 21698 2201 21712 2215
rect 8714 2177 8728 2191
rect 8786 2177 8800 2191
rect 8858 2177 8872 2191
rect 17426 2177 17440 2191
rect 21746 2177 21760 2191
rect 8810 2153 8824 2167
rect 18506 2153 18520 2167
rect 9002 2129 9016 2143
rect 12338 2129 12352 2143
rect 13250 2129 13264 2143
rect 14642 2129 14656 2143
rect 27194 2129 27208 2143
rect 9770 2105 9784 2119
rect 16994 2105 17008 2119
rect 26666 2105 26680 2119
rect 10082 2081 10096 2095
rect 10130 2081 10144 2095
rect 23474 2081 23488 2095
rect 10154 2057 10168 2071
rect 10682 2057 10696 2071
rect 16634 2057 16648 2071
rect 17738 2057 17752 2071
rect 18866 2057 18880 2071
rect 24794 2057 24808 2071
rect 10202 2033 10216 2047
rect 14450 2033 14464 2047
rect 16634 2033 16648 2047
rect 16682 2033 16696 2047
rect 10274 2009 10288 2023
rect 10322 2009 10336 2023
rect 10394 2009 10408 2023
rect 18242 2009 18256 2023
rect 24170 2009 24184 2023
rect 10322 1985 10336 1999
rect 11522 1985 11536 1999
rect 11594 1985 11608 1999
rect 23114 1985 23128 1999
rect 10658 1961 10672 1975
rect 27565 1961 27579 1975
rect 10970 1937 10984 1951
rect 14762 1937 14776 1951
rect 27218 1937 27232 1951
rect 27565 1937 27579 1951
rect 11018 1913 11032 1927
rect 14954 1913 14968 1927
rect 27194 1913 27208 1927
rect 27565 1913 27579 1927
rect 11042 1889 11056 1903
rect 11690 1889 11704 1903
rect 11762 1889 11776 1903
rect 23354 1889 23368 1903
rect 27098 1889 27112 1903
rect 27565 1889 27579 1903
rect 11138 1865 11152 1879
rect 11234 1865 11248 1879
rect 11378 1865 11392 1879
rect 18962 1865 18976 1879
rect 20594 1865 20608 1879
rect 20930 1865 20944 1879
rect 27170 1865 27184 1879
rect 27565 1865 27579 1879
rect 11642 1841 11656 1855
rect 16946 1841 16960 1855
rect 20930 1841 20944 1855
rect 21458 1841 21472 1855
rect 27146 1841 27160 1855
rect 27565 1841 27579 1855
rect 16946 1817 16960 1831
rect 17090 1817 17104 1831
rect 27122 1817 27136 1831
rect 27565 1817 27579 1831
rect 12578 984 12592 998
rect 22082 984 22096 998
rect 12386 960 12400 974
rect 16994 960 17008 974
rect 12242 936 12256 950
rect 16250 936 16264 950
rect 19082 936 19096 950
rect 23954 936 23968 950
rect 11810 912 11824 926
rect 20546 912 20560 926
rect 11690 888 11704 902
rect 25370 888 25384 902
rect 10034 864 10048 878
rect 10850 864 10864 878
rect 23714 864 23728 878
rect 8498 840 8512 854
rect 22922 840 22936 854
rect 8378 816 8392 830
rect 19178 816 19192 830
rect 20114 816 20128 830
rect 22178 816 22192 830
rect 8210 792 8224 806
rect 15602 792 15616 806
rect 18074 792 18088 806
rect 18266 792 18280 806
rect 23018 792 23032 806
rect 7994 768 8008 782
rect 13754 768 13768 782
rect 14210 768 14224 782
rect 25130 768 25144 782
rect 7970 744 7984 758
rect 8810 744 8824 758
rect 10466 744 10480 758
rect 11906 744 11920 758
rect 14090 744 14104 758
rect 16130 744 16144 758
rect 16730 744 16744 758
rect 23354 744 23368 758
rect 26330 744 26344 758
rect 7538 720 7552 734
rect 16466 720 16480 734
rect 17522 720 17536 734
rect 20834 720 20848 734
rect 7298 696 7312 710
rect 10754 696 10768 710
rect 11090 696 11104 710
rect 11786 696 11800 710
rect 12098 696 12112 710
rect 20450 696 20464 710
rect 20762 696 20776 710
rect 21698 696 21712 710
rect 7034 672 7048 686
rect 16706 672 16720 686
rect 17162 672 17176 686
rect 19706 672 19720 686
rect 20810 672 20824 686
rect 6818 648 6832 662
rect 9098 648 9112 662
rect 9794 648 9808 662
rect 15842 648 15856 662
rect 22034 648 22048 662
rect 6794 624 6808 638
rect 20858 624 20872 638
rect 6770 600 6784 614
rect 14522 600 14536 614
rect 15890 600 15904 614
rect 22154 600 22168 614
rect 22970 600 22984 614
rect 23114 600 23128 614
rect 6698 576 6712 590
rect 19850 576 19864 590
rect 25034 576 25048 590
rect 6554 552 6568 566
rect 26306 552 26320 566
rect 6482 528 6496 542
rect 16082 528 16096 542
rect 16802 528 16816 542
rect 22322 528 22336 542
rect 22490 528 22504 542
rect 23762 528 23776 542
rect 6458 504 6472 518
rect 8978 504 8992 518
rect 9698 504 9712 518
rect 10922 504 10936 518
rect 26042 504 26056 518
rect 5546 480 5560 494
rect 17858 480 17872 494
rect 5498 456 5512 470
rect 22538 456 22552 470
rect 5474 432 5488 446
rect 6602 432 6616 446
rect 6674 432 6688 446
rect 12842 432 12856 446
rect 25250 432 25264 446
rect 5234 408 5248 422
rect 23210 408 23224 422
rect 5018 384 5032 398
rect 7010 384 7024 398
rect 7826 384 7840 398
rect 14354 384 14368 398
rect 22298 384 22312 398
rect 22802 384 22816 398
rect 23282 384 23296 398
rect 26306 384 26320 398
rect 4586 360 4600 374
rect 16370 360 16384 374
rect 4490 336 4504 350
rect 12914 336 12928 350
rect 13442 336 13456 350
rect 26210 336 26224 350
rect 4298 312 4312 326
rect 13610 312 13624 326
rect 13658 312 13672 326
rect 24002 312 24016 326
rect 4202 288 4216 302
rect 17714 288 17728 302
rect 4154 264 4168 278
rect 13706 264 13720 278
rect 14474 264 14488 278
rect 15410 264 15424 278
rect 15986 264 16000 278
rect 22202 264 22216 278
rect 3866 240 3880 254
rect 4682 240 4696 254
rect 8186 240 8200 254
rect 20258 240 20272 254
rect 26354 240 26368 254
rect 3482 216 3496 230
rect 13466 216 13480 230
rect 13682 216 13696 230
rect 14018 216 14032 230
rect 14498 216 14512 230
rect 17570 216 17584 230
rect 2666 192 2680 206
rect 4562 192 4576 206
rect 4730 192 4744 206
rect 19034 192 19048 206
rect 24050 192 24064 206
rect 2450 168 2464 182
rect 12938 168 12952 182
rect 13778 168 13792 182
rect 2378 144 2392 158
rect 14114 144 14128 158
rect 26378 144 26392 158
rect 27565 144 27579 158
rect 70 120 84 134
rect 3602 120 3616 134
rect 3698 120 3712 134
rect 8642 120 8656 134
rect 8858 120 8872 134
rect 11282 120 11296 134
rect 25226 120 25240 134
rect 26402 120 26416 134
rect 70 96 84 110
rect 2642 96 2656 110
rect 2714 96 2728 110
rect 23642 96 23656 110
rect 25106 96 25120 110
rect 26354 96 26368 110
rect 27565 96 27579 110
rect 70 72 84 86
rect 5594 72 5608 86
rect 6266 72 6280 86
rect 8882 72 8896 86
rect 8930 72 8944 86
rect 13802 72 13816 86
rect 26330 72 26344 86
rect 27565 72 27579 86
rect 70 48 84 62
rect 2234 48 2248 62
rect 2330 48 2344 62
rect 23186 48 23200 62
rect 26306 48 26320 62
rect 27565 48 27579 62
rect 5354 24 5368 38
rect 26378 24 26392 38
rect 26402 24 26416 38
rect 27565 24 27579 38
rect 9962 0 9976 14
rect 27565 0 27579 14
<< metal2 >>
rect 0 8027 70 8039
rect 0 8003 70 8015
rect 0 7979 70 7991
rect 123 7872 323 8170
rect 339 7872 351 8170
rect 363 7872 375 8170
rect 387 7872 399 8170
rect 411 7872 423 8170
rect 1731 7872 1743 8002
rect 2307 7872 2319 8002
rect 2883 7872 2895 8050
rect 3075 7968 3087 8170
rect 3267 7872 3279 8074
rect 3699 7872 3711 7930
rect 4107 7872 4119 8098
rect 4587 7920 4599 8170
rect 4623 8088 4635 8170
rect 6903 8088 6915 8170
rect 6904 8074 6922 8088
rect 6891 7872 6903 8074
rect 9123 8040 9135 8170
rect 10635 8088 10647 8170
rect 7827 7872 7839 7906
rect 8763 7872 8775 8026
rect 8883 7872 8895 7906
rect 10131 7872 10143 7978
rect 10707 7872 10719 7978
rect 12147 7896 12159 8170
rect 12183 7920 12195 8170
rect 14463 8160 14475 8170
rect 14464 8146 14482 8160
rect 12363 7872 12375 7906
rect 12867 7872 12879 8122
rect 14451 7872 14463 8146
rect 15195 7992 15207 8170
rect 18171 8160 18183 8170
rect 18195 8112 18207 8170
rect 20559 8160 20571 8170
rect 22215 8160 22227 8170
rect 20560 8146 20578 8160
rect 22216 8146 22234 8160
rect 16659 7872 16671 7882
rect 18171 7872 18183 7978
rect 18315 7872 18327 8146
rect 18363 7872 18375 7882
rect 19707 7872 19719 8098
rect 19947 7872 19959 8074
rect 20547 7872 20559 8146
rect 22203 7872 22215 8146
rect 22695 8064 22707 8170
rect 24195 8040 24207 8170
rect 25695 8136 25707 8170
rect 23739 7872 23751 8026
rect 23979 7872 23991 7954
rect 24099 7872 24111 8026
rect 26091 7872 26103 8074
rect 27020 7993 27032 8026
rect 27048 7968 27060 8002
rect 27099 7872 27111 8002
rect 27126 7896 27138 7978
rect 27179 7944 27191 8098
rect 27155 7896 27167 7930
rect 27243 7872 27443 8170
rect 27579 8027 27649 8039
rect 27579 8003 27649 8015
rect 27579 7979 27649 7991
rect 27579 7955 27649 7967
rect 27579 7931 27649 7943
rect 27579 7907 27649 7919
rect 27579 7883 27649 7895
rect 0 4266 70 4278
rect 0 4242 70 4254
rect 0 4218 70 4230
rect 0 4194 70 4206
rect 123 1807 323 7073
rect 339 1807 351 7073
rect 363 1807 375 7073
rect 387 1807 399 7073
rect 411 1807 423 7073
rect 1611 4303 1623 7073
rect 1659 4327 1671 7073
rect 1683 1807 1695 4337
rect 1731 4183 1743 7073
rect 1779 4159 1791 7073
rect 1803 4375 1815 7073
rect 1827 4399 1839 7073
rect 1875 4423 1887 7073
rect 1899 4447 1911 7073
rect 1947 4471 1959 7073
rect 1995 4231 2007 7073
rect 2043 4231 2055 7073
rect 2115 4495 2127 7073
rect 2139 4519 2151 7073
rect 2043 1807 2055 4121
rect 2091 1807 2103 4097
rect 2163 4087 2175 7073
rect 2211 4543 2223 7073
rect 2235 4591 2247 7073
rect 2235 1807 2247 4553
rect 2259 4063 2271 7073
rect 2283 4615 2295 7073
rect 2355 4639 2367 7073
rect 2403 4663 2415 7073
rect 2475 4687 2487 7073
rect 2499 4711 2511 7073
rect 2523 4735 2535 7073
rect 2571 4759 2583 7073
rect 2283 1807 2295 4025
rect 2307 1807 2319 4289
rect 2403 1807 2415 4001
rect 2595 3991 2607 7073
rect 2619 4783 2631 7073
rect 2667 4807 2679 7073
rect 2691 4831 2703 7073
rect 2499 1807 2511 3977
rect 2523 1807 2535 3953
rect 2571 1807 2583 3929
rect 2619 1807 2631 3905
rect 2715 3895 2727 7073
rect 2763 4855 2775 7073
rect 2811 4879 2823 7073
rect 2883 3871 2895 7073
rect 2763 1807 2775 3857
rect 2907 1807 2919 4889
rect 2931 3871 2943 7073
rect 2955 4927 2967 7073
rect 3003 4951 3015 7073
rect 3051 3847 3063 7073
rect 3075 3823 3087 7073
rect 3099 4975 3111 7073
rect 3123 4999 3135 7073
rect 3171 3799 3183 7073
rect 3195 4591 3207 7073
rect 3219 5023 3231 7073
rect 3243 5047 3255 7073
rect 3315 5071 3327 7073
rect 3339 5095 3351 7073
rect 3363 5119 3375 7073
rect 3267 1807 3279 4505
rect 3411 4471 3423 7073
rect 3435 5143 3447 7073
rect 3483 5167 3495 7073
rect 3531 5191 3543 7073
rect 3555 5215 3567 7073
rect 3315 1807 3327 3761
rect 3459 1807 3471 3737
rect 3531 1807 3543 3713
rect 3579 1807 3591 3905
rect 3603 3703 3615 7073
rect 3651 5239 3663 7073
rect 3675 4615 3687 7073
rect 3747 5263 3759 7073
rect 3795 5023 3807 7073
rect 3867 5023 3879 7073
rect 3891 5287 3903 7073
rect 3627 1807 3639 3809
rect 3675 1807 3687 3809
rect 3747 1807 3759 3665
rect 3795 1807 3807 3641
rect 3819 1807 3831 3617
rect 3843 1807 3855 3737
rect 3891 1807 3903 3593
rect 3915 3583 3927 7073
rect 3963 5311 3975 7073
rect 3987 5335 3999 7073
rect 3939 1807 3951 3545
rect 3963 1807 3975 3521
rect 3987 1807 3999 3497
rect 4011 3487 4023 7073
rect 4059 5359 4071 7073
rect 4083 3607 4095 7073
rect 4035 1807 4047 3449
rect 4155 3439 4167 7073
rect 4179 3655 4191 7073
rect 4083 1807 4095 3425
rect 4179 1807 4191 3593
rect 4203 3439 4215 7073
rect 4251 5383 4263 7073
rect 4275 5407 4287 7073
rect 4299 5431 4311 7073
rect 4251 1807 4263 3401
rect 4275 1807 4287 3377
rect 4347 3367 4359 7073
rect 4371 5455 4383 7073
rect 4347 1807 4359 3329
rect 4371 1807 4383 3305
rect 4395 1807 4407 3281
rect 4419 3271 4431 7073
rect 4443 1807 4455 4121
rect 4467 3247 4479 7073
rect 4491 5383 4503 7073
rect 4515 4327 4527 7073
rect 4467 1807 4479 3209
rect 4539 3199 4551 7073
rect 4587 5479 4599 7073
rect 4611 3967 4623 7073
rect 4659 5503 4671 7073
rect 4707 5095 4719 7073
rect 4755 3223 4767 7073
rect 4539 1807 4551 3161
rect 4611 1807 4623 3137
rect 4659 1807 4671 3113
rect 4779 1807 4791 5153
rect 4827 4447 4839 7073
rect 4851 5527 4863 7073
rect 4875 5551 4887 7073
rect 4803 1807 4815 3089
rect 4827 1807 4839 3065
rect 4899 3055 4911 7073
rect 4875 1807 4887 3041
rect 4923 1807 4935 3017
rect 4947 3007 4959 7073
rect 4971 5575 4983 7073
rect 4995 5599 5007 7073
rect 4995 1807 5007 3953
rect 5043 2983 5055 7073
rect 5091 5623 5103 7073
rect 5163 5647 5175 7073
rect 5187 5671 5199 7073
rect 5211 5695 5223 7073
rect 5259 5719 5271 7073
rect 5283 3991 5295 7073
rect 5067 1807 5079 2945
rect 5115 1807 5127 2921
rect 5139 1807 5151 3617
rect 5187 1807 5199 2897
rect 5259 1807 5271 2873
rect 5283 1807 5295 3185
rect 5307 2863 5319 7073
rect 5355 5743 5367 7073
rect 5307 1807 5319 2825
rect 5355 1807 5367 4433
rect 5379 3199 5391 7073
rect 5403 5767 5415 7073
rect 5451 5791 5463 7073
rect 5499 5815 5511 7073
rect 5571 3919 5583 7073
rect 5403 1807 5415 2801
rect 5595 1807 5607 7073
rect 5619 5863 5631 7073
rect 5667 5839 5679 7073
rect 5691 4111 5703 7073
rect 5715 1807 5727 5873
rect 5739 2791 5751 7073
rect 5787 5911 5799 7073
rect 5811 3751 5823 7073
rect 5835 5671 5847 7073
rect 5859 5935 5871 7073
rect 5907 2767 5919 7073
rect 5931 4519 5943 7073
rect 5955 5959 5967 7073
rect 6003 3319 6015 7073
rect 6027 2959 6039 7073
rect 6051 5983 6063 7073
rect 6075 2743 6087 7073
rect 6123 3775 6135 7073
rect 6147 5287 6159 7073
rect 6123 1807 6135 2705
rect 6171 2695 6183 7073
rect 6219 5911 6231 7073
rect 6267 4687 6279 7073
rect 6291 1807 6303 5993
rect 6315 1807 6327 6017
rect 6339 3319 6351 7073
rect 6363 3631 6375 7073
rect 6339 1807 6351 2657
rect 6363 1807 6375 3353
rect 6387 2647 6399 7073
rect 6411 3367 6423 7073
rect 6483 3367 6495 7073
rect 6507 6055 6519 7073
rect 6411 1807 6423 2681
rect 6435 2671 6447 3353
rect 6435 1807 6447 2609
rect 6507 1807 6519 4169
rect 6531 3391 6543 6041
rect 6555 3127 6567 7073
rect 6579 6055 6591 7073
rect 6651 5215 6663 7073
rect 6579 1807 6591 3977
rect 6651 1807 6663 4289
rect 6675 4183 6687 7073
rect 6723 2695 6735 7073
rect 6771 6079 6783 7073
rect 6795 5311 6807 7073
rect 6819 5671 6831 7073
rect 6843 3871 6855 7073
rect 6747 1807 6759 2657
rect 6867 1807 6879 4025
rect 6891 2839 6903 7073
rect 6915 1807 6927 5657
rect 6939 3871 6951 7073
rect 6963 2839 6975 7073
rect 6987 6103 6999 7073
rect 7035 6127 7047 7073
rect 6987 1807 6999 3977
rect 7059 3967 7071 7073
rect 7083 2599 7095 7073
rect 7131 3967 7143 7073
rect 7155 4519 7167 7073
rect 7203 6151 7215 7073
rect 7083 1807 7095 2561
rect 7131 1807 7143 3737
rect 7251 3223 7263 7073
rect 7275 4111 7287 7073
rect 7299 6175 7311 7073
rect 7323 5335 7335 7073
rect 7203 1807 7215 2537
rect 7227 1807 7239 2513
rect 7251 1807 7263 2489
rect 7323 1807 7335 4001
rect 7347 2479 7359 7073
rect 7395 6199 7407 7073
rect 7419 6223 7431 7073
rect 7347 1807 7359 2441
rect 7395 1807 7407 3017
rect 7419 1807 7431 3377
rect 7443 2431 7455 7073
rect 7467 1807 7479 5057
rect 7491 3631 7503 7073
rect 7515 4135 7527 7073
rect 7539 5479 7551 7073
rect 7587 6247 7599 7073
rect 7611 6271 7623 7073
rect 7515 1807 7527 2393
rect 7563 1807 7575 2753
rect 7587 2407 7599 5753
rect 7611 1807 7623 3929
rect 7635 2767 7647 7073
rect 7635 1807 7647 2393
rect 7659 2383 7671 7073
rect 7683 4855 7695 7073
rect 7659 1807 7671 2345
rect 7707 1807 7719 6137
rect 7731 4543 7743 7073
rect 7755 4855 7767 7073
rect 7779 6295 7791 7073
rect 7731 1807 7743 2393
rect 7779 1807 7791 6065
rect 7803 4927 7815 7073
rect 7851 1807 7863 5081
rect 7875 3967 7887 7073
rect 7899 3775 7911 7073
rect 7875 1807 7887 2321
rect 7923 1807 7935 5057
rect 7947 1807 7959 3617
rect 7995 2527 8007 7073
rect 8067 6319 8079 7073
rect 8043 1807 8055 5057
rect 8091 1807 8103 2297
rect 8115 2287 8127 7073
rect 8187 6343 8199 7073
rect 8163 1807 8175 5081
rect 8211 4015 8223 7073
rect 8235 4855 8247 7073
rect 8187 1807 8199 3353
rect 8259 1807 8271 4841
rect 8283 4447 8295 7073
rect 8307 5551 8319 7073
rect 8331 2263 8343 5633
rect 8355 3391 8367 7073
rect 8403 5599 8415 7073
rect 8427 4927 8439 7073
rect 8451 5599 8463 7073
rect 8307 1807 8319 2249
rect 8403 1807 8415 2249
rect 8427 1807 8439 4289
rect 8499 2719 8511 7073
rect 8451 1807 8463 2225
rect 8523 1807 8535 6353
rect 8547 1807 8559 6377
rect 8571 5623 8583 7073
rect 8643 6415 8655 7073
rect 8571 1807 8583 2201
rect 8619 1807 8631 5321
rect 8643 1807 8655 5777
rect 8667 1807 8679 6425
rect 8715 4399 8727 7073
rect 8739 6463 8751 7073
rect 8715 1807 8727 2177
rect 8739 1807 8751 2393
rect 8763 1807 8775 4385
rect 8787 2191 8799 4793
rect 8811 2167 8823 7073
rect 8835 6487 8847 7073
rect 8835 1807 8847 3977
rect 8859 2191 8871 7073
rect 8931 6511 8943 7073
rect 8955 6535 8967 7073
rect 8979 5791 8991 7073
rect 8955 1807 8967 3953
rect 9003 2143 9015 7073
rect 9051 6559 9063 7073
rect 9075 6583 9087 7073
rect 9099 2551 9111 7073
rect 9147 2911 9159 7073
rect 9195 4615 9207 7073
rect 9267 3463 9279 7073
rect 9291 5791 9303 7073
rect 9339 6607 9351 7073
rect 9387 2551 9399 7073
rect 9411 4783 9423 7073
rect 9435 2359 9447 7073
rect 9459 4783 9471 7073
rect 9507 3943 9519 7073
rect 9531 3775 9543 7073
rect 9555 2935 9567 7073
rect 9507 1807 9519 2537
rect 9603 2359 9615 7073
rect 9627 6631 9639 7073
rect 9675 6655 9687 7073
rect 9723 6679 9735 7073
rect 9747 6703 9759 7073
rect 9651 1807 9663 5489
rect 9675 1807 9687 3977
rect 9747 1807 9759 3473
rect 9771 3175 9783 7073
rect 9819 5527 9831 7073
rect 9843 6727 9855 7073
rect 9867 6751 9879 7073
rect 9891 6775 9903 7073
rect 9939 6799 9951 7073
rect 9771 1807 9783 2105
rect 9843 1807 9855 3617
rect 9867 1807 9879 4097
rect 9891 1807 9903 5897
rect 9939 1807 9951 5369
rect 9963 3487 9975 7073
rect 9987 4975 9999 7073
rect 10035 3943 10047 7073
rect 10059 5287 10071 7073
rect 10083 6823 10095 7073
rect 9963 1807 9975 3161
rect 9987 1807 9999 3449
rect 10059 1807 10071 4961
rect 10083 1807 10095 2081
rect 10107 1807 10119 6833
rect 10131 2095 10143 7073
rect 10179 3391 10191 7073
rect 10203 6871 10215 7073
rect 10227 5983 10239 7073
rect 10275 5743 10287 7073
rect 10299 6511 10311 7073
rect 10155 1807 10167 2057
rect 10203 1807 10215 2033
rect 10275 1807 10287 2009
rect 10299 1807 10311 3209
rect 10323 2023 10335 6161
rect 10347 5023 10359 7073
rect 10323 1807 10335 1985
rect 10371 1807 10383 6665
rect 10395 2527 10407 7073
rect 10419 6895 10431 7073
rect 10443 4759 10455 7073
rect 10395 1807 10407 2009
rect 10419 1807 10431 3833
rect 10467 1807 10479 6857
rect 10491 4759 10503 7073
rect 10515 6847 10527 7073
rect 10539 3847 10551 7073
rect 10563 6655 10575 7073
rect 10587 6319 10599 7073
rect 10635 5575 10647 7073
rect 10659 5359 10671 7073
rect 10515 1807 10527 3185
rect 10587 1807 10599 5057
rect 10611 1807 10623 5225
rect 10635 1807 10647 4601
rect 10683 2071 10695 7073
rect 10659 1807 10671 1961
rect 10707 1807 10719 4601
rect 10731 1807 10743 6305
rect 10755 3943 10767 7073
rect 10779 4831 10791 7073
rect 10803 6655 10815 7073
rect 10803 1807 10815 4697
rect 10827 2407 10839 6881
rect 10851 5527 10863 7073
rect 10875 5551 10887 7073
rect 10923 5143 10935 7073
rect 10971 5143 10983 7073
rect 10947 1807 10959 3761
rect 10995 3631 11007 7073
rect 11019 4015 11031 7073
rect 11043 6127 11055 7073
rect 11091 6535 11103 7073
rect 11115 6127 11127 7073
rect 11139 6007 11151 7073
rect 11187 5527 11199 7073
rect 11211 6007 11223 7073
rect 11259 6847 11271 7073
rect 11307 6607 11319 7073
rect 10971 1807 10983 1937
rect 11019 1807 11031 1913
rect 11043 1807 11055 1889
rect 11139 1807 11151 1865
rect 11163 1807 11175 3977
rect 11211 1807 11223 5369
rect 11235 1879 11247 6065
rect 11259 1807 11271 6329
rect 11283 3391 11295 5993
rect 11307 1807 11319 6233
rect 11331 4327 11343 7073
rect 11355 6007 11367 7073
rect 11403 5167 11415 7073
rect 11427 6775 11439 7073
rect 11355 1807 11367 5153
rect 11379 1807 11391 1865
rect 11403 1807 11415 3089
rect 11427 1807 11439 4529
rect 11451 2335 11463 7073
rect 11475 3535 11487 7073
rect 11475 1807 11487 3209
rect 11499 1807 11511 6233
rect 11523 1999 11535 7073
rect 11547 3631 11559 7073
rect 11595 6775 11607 7073
rect 11643 6895 11655 7073
rect 11667 6655 11679 7073
rect 11547 1807 11559 3521
rect 11595 1807 11607 1985
rect 11619 1807 11631 6641
rect 11643 1807 11655 1841
rect 11667 1807 11679 5897
rect 11691 1903 11703 7073
rect 11739 6919 11751 7073
rect 11715 3175 11727 6641
rect 11739 1807 11751 6065
rect 11763 5335 11775 7073
rect 11787 4975 11799 6905
rect 11811 6655 11823 7073
rect 11763 1807 11775 1889
rect 11835 1807 11847 6665
rect 11859 5815 11871 7073
rect 11883 6919 11895 7073
rect 11883 1807 11895 5321
rect 11907 3655 11919 7073
rect 11931 6943 11943 7073
rect 11979 6967 11991 7073
rect 12003 6919 12015 7073
rect 11931 1807 11943 4289
rect 11955 3031 11967 6905
rect 11979 1807 11991 3761
rect 12003 1807 12015 3953
rect 12051 3487 12063 7073
rect 12027 1807 12039 3329
rect 12099 3199 12111 7073
rect 12123 3967 12135 7073
rect 12147 4111 12159 7073
rect 12171 3655 12183 7073
rect 12195 6031 12207 7073
rect 12243 3967 12255 7073
rect 12267 6031 12279 7073
rect 12075 1807 12087 2849
rect 12123 1807 12135 3257
rect 12147 1807 12159 2513
rect 12171 1807 12183 3257
rect 12219 1807 12231 3449
rect 12291 3319 12303 7073
rect 12315 2863 12327 7073
rect 12363 3271 12375 7073
rect 12291 1807 12303 2345
rect 12339 1807 12351 2129
rect 12363 1807 12375 2393
rect 12387 2263 12399 6929
rect 12411 3655 12423 7073
rect 12435 6871 12447 7073
rect 12483 6511 12495 7073
rect 12435 1807 12447 3449
rect 12459 1807 12471 5801
rect 12507 1807 12519 3545
rect 12531 3199 12543 7073
rect 12555 3223 12567 7073
rect 12579 5167 12591 7073
rect 12555 1807 12567 2465
rect 12603 1807 12615 3881
rect 12627 3439 12639 7073
rect 12651 5167 12663 7073
rect 12675 5431 12687 7073
rect 12699 6943 12711 7073
rect 12627 1807 12639 3257
rect 12675 1807 12687 3281
rect 12699 1807 12711 4097
rect 12723 1807 12735 3881
rect 12747 3631 12759 7073
rect 12771 5311 12783 7073
rect 12795 5335 12807 7073
rect 12819 6991 12831 7073
rect 12771 1807 12783 4289
rect 12795 1807 12807 3425
rect 12819 1807 12831 6521
rect 12843 2311 12855 6953
rect 12867 3271 12879 7073
rect 12891 3367 12903 6905
rect 12915 5431 12927 7073
rect 12939 5527 12951 7073
rect 12963 5383 12975 7073
rect 12987 5815 12999 7073
rect 13011 4639 13023 7073
rect 12867 1807 12879 2465
rect 12963 1807 12975 3257
rect 13011 1807 13023 2345
rect 13035 1807 13047 5273
rect 13059 4639 13071 7073
rect 13083 6919 13095 7073
rect 13131 6967 13143 7073
rect 13143 3919 13155 6929
rect 13179 4423 13191 7073
rect 13203 4447 13215 7073
rect 13059 1807 13071 3785
rect 13107 1807 13119 3785
rect 13227 3103 13239 7073
rect 13275 6943 13287 7073
rect 13323 6031 13335 7073
rect 13287 3271 13299 6017
rect 13179 1807 13191 2249
rect 13251 1807 13263 2129
rect 13323 1807 13335 3305
rect 13347 1807 13359 5273
rect 13371 1807 13383 3857
rect 13395 3559 13407 7073
rect 13419 7015 13431 7073
rect 13419 1807 13431 4817
rect 13443 3415 13455 4625
rect 13467 3607 13479 7073
rect 13515 7039 13527 7073
rect 13539 5863 13551 7073
rect 13491 2263 13503 5609
rect 13515 1807 13527 5513
rect 13539 1807 13551 5417
rect 13563 4639 13575 7073
rect 13587 5887 13599 7073
rect 13563 1807 13575 3857
rect 13611 3127 13623 6017
rect 13635 5863 13647 7073
rect 13659 6079 13671 7073
rect 13683 5071 13695 7073
rect 13707 3535 13719 7001
rect 13731 6511 13743 7073
rect 13755 6847 13767 7073
rect 13779 6079 13791 7073
rect 13803 4015 13815 7073
rect 13827 5887 13839 7073
rect 13635 1807 13647 3257
rect 13851 1807 13863 6713
rect 13875 4447 13887 7073
rect 13899 7015 13911 7073
rect 13899 1807 13911 6905
rect 13923 5551 13935 7073
rect 13947 3271 13959 7073
rect 13971 1807 13983 6929
rect 13995 3391 14007 7073
rect 14019 4447 14031 7073
rect 14043 3367 14055 7073
rect 14067 6031 14079 7073
rect 14115 6079 14127 7073
rect 14079 3271 14091 5513
rect 14139 3799 14151 7001
rect 14163 4807 14175 7073
rect 13995 1807 14007 3257
rect 14067 1807 14079 2321
rect 14163 1807 14175 3353
rect 14187 1807 14199 4169
rect 14211 3367 14223 6641
rect 14235 5383 14247 7073
rect 14259 6847 14271 7073
rect 14307 6631 14319 7073
rect 14259 1807 14271 4289
rect 14283 1807 14295 5081
rect 14307 1807 14319 6113
rect 14331 2239 14343 6833
rect 14355 4111 14367 7073
rect 14379 6631 14391 7073
rect 14403 6847 14415 7073
rect 14355 1807 14367 3353
rect 14403 1807 14415 5321
rect 14427 3367 14439 6737
rect 14451 2047 14463 7073
rect 14499 7015 14511 7073
rect 14475 2839 14487 6833
rect 14523 5695 14535 7073
rect 14547 6847 14559 7073
rect 14571 5887 14583 7073
rect 14595 5263 14607 7073
rect 14571 1807 14583 3353
rect 14619 1807 14631 4049
rect 14643 2143 14655 7073
rect 14667 3487 14679 7073
rect 14691 6391 14703 7073
rect 14739 5263 14751 7073
rect 14691 1807 14703 4073
rect 14715 1807 14727 4049
rect 14739 1807 14751 4193
rect 14763 1951 14775 7073
rect 14787 4903 14799 7073
rect 14835 6391 14847 7073
rect 14787 1807 14799 2417
rect 14811 1807 14823 6137
rect 14835 1807 14847 6257
rect 14859 4015 14871 7073
rect 14883 7063 14895 7073
rect 14883 1807 14895 6593
rect 14907 1807 14919 6233
rect 14931 1807 14943 4193
rect 14955 1927 14967 7049
rect 15003 3151 15015 7073
rect 15411 6703 15423 7073
rect 15051 1807 15063 5585
rect 15555 4903 15567 7073
rect 15579 5599 15591 7073
rect 15603 6583 15615 7073
rect 15723 6271 15735 7073
rect 15459 1807 15471 2993
rect 15651 1807 15663 4169
rect 15723 1807 15735 6137
rect 15747 1807 15759 5729
rect 15807 4783 15819 6257
rect 15771 1807 15783 3641
rect 15795 1807 15807 4169
rect 15867 1807 15879 4505
rect 15939 1807 15951 3929
rect 15963 1807 15975 4097
rect 16035 1807 16047 4505
rect 16059 1807 16071 4121
rect 16083 3319 16095 7073
rect 16131 3991 16143 7073
rect 16155 1807 16167 5081
rect 16275 4783 16287 7073
rect 16299 3199 16311 7073
rect 16323 5695 16335 7073
rect 16371 5695 16383 7073
rect 16395 5887 16407 7073
rect 16419 6439 16431 7073
rect 16323 1807 16335 4073
rect 16347 1807 16359 3473
rect 16419 1807 16431 5729
rect 16443 5407 16455 7073
rect 16443 1807 16455 3641
rect 16491 3199 16503 7073
rect 16515 5791 16527 7073
rect 16539 6271 16551 7073
rect 16539 1807 16551 5801
rect 16563 1807 16575 3521
rect 16587 3463 16599 7073
rect 16611 4879 16623 7073
rect 16611 1807 16623 4313
rect 16635 2071 16647 7073
rect 16659 3439 16671 6257
rect 16683 2047 16695 6881
rect 16707 5287 16719 7073
rect 16731 4135 16743 7073
rect 16755 4831 16767 7073
rect 16779 4327 16791 6377
rect 16803 5815 16815 7073
rect 16827 5407 16839 7073
rect 16635 1807 16647 2033
rect 16755 1807 16767 4313
rect 16827 1807 16839 5081
rect 16851 4783 16863 7073
rect 16875 3823 16887 5393
rect 16899 4879 16911 7073
rect 16923 5407 16935 7073
rect 16851 1807 16863 2633
rect 16899 1807 16911 3929
rect 16923 1807 16935 4505
rect 16947 1855 16959 7073
rect 16971 2503 16983 4865
rect 16995 2119 17007 7073
rect 17043 5863 17055 7073
rect 16947 1807 16959 1817
rect 17019 1807 17031 3953
rect 17043 1807 17055 4313
rect 17067 3631 17079 5393
rect 17091 1831 17103 6065
rect 17115 4879 17127 7073
rect 17139 3895 17151 7073
rect 17163 6823 17175 7073
rect 17187 4351 17199 7073
rect 17235 6607 17247 7073
rect 17283 5407 17295 7073
rect 17355 5695 17367 7073
rect 17379 5791 17391 7073
rect 17427 2191 17439 7073
rect 17475 4807 17487 7073
rect 17499 3631 17511 7073
rect 17523 4063 17535 7073
rect 17571 3631 17583 7073
rect 17595 5863 17607 7073
rect 17619 5527 17631 7073
rect 17643 6199 17655 7073
rect 17763 4999 17775 7073
rect 17739 1807 17751 2057
rect 17763 1807 17775 4337
rect 17811 1807 17823 2585
rect 17835 1807 17847 2729
rect 17883 1807 17895 2513
rect 17907 1807 17919 4049
rect 17955 1807 17967 6929
rect 17979 1807 17991 6905
rect 18003 1807 18015 5417
rect 18051 1807 18063 6641
rect 18171 4999 18183 7073
rect 18123 1807 18135 3929
rect 18171 1807 18183 3593
rect 18195 1807 18207 4457
rect 18219 1807 18231 5345
rect 18243 2023 18255 4985
rect 18291 1807 18303 6137
rect 18315 4999 18327 7073
rect 18315 1807 18327 4577
rect 18339 4351 18351 4985
rect 18363 4063 18375 7073
rect 18411 6103 18423 7073
rect 18363 1807 18375 2801
rect 18387 1807 18399 5537
rect 18435 4519 18447 7073
rect 18459 4879 18471 7073
rect 18411 1807 18423 4337
rect 18459 1807 18471 4649
rect 18483 1807 18495 6497
rect 18507 4471 18519 7073
rect 18531 3775 18543 7073
rect 18555 6823 18567 7073
rect 18507 1807 18519 2153
rect 18555 1807 18567 6689
rect 18603 3823 18615 7073
rect 18627 5095 18639 7073
rect 18651 4591 18663 7073
rect 18579 1807 18591 2705
rect 18675 1807 18687 3401
rect 18699 2335 18711 7073
rect 18723 4351 18735 6929
rect 18747 3655 18759 7073
rect 18819 5383 18831 7073
rect 18843 6511 18855 7073
rect 18747 1807 18759 3449
rect 18771 1807 18783 4937
rect 18795 1807 18807 2273
rect 18819 1807 18831 5057
rect 18843 1807 18855 4337
rect 18867 2071 18879 6809
rect 18891 5431 18903 7073
rect 18891 1807 18903 5369
rect 18915 1807 18927 4433
rect 18939 2695 18951 7073
rect 18987 4879 18999 7073
rect 18963 1807 18975 1865
rect 19011 1807 19023 4049
rect 19035 3463 19047 5393
rect 19059 4999 19071 7073
rect 19083 3727 19095 7073
rect 19131 5359 19143 7073
rect 19131 1807 19143 3665
rect 19179 2575 19191 7073
rect 19203 4183 19215 7073
rect 19227 5407 19239 7073
rect 19155 1807 19167 2321
rect 19275 2311 19287 7073
rect 19299 5527 19311 7073
rect 19323 5575 19335 7073
rect 19371 4303 19383 7073
rect 19299 1807 19311 4217
rect 19395 3175 19407 7073
rect 19419 5575 19431 7073
rect 19467 4399 19479 7073
rect 19491 2455 19503 7073
rect 19515 4327 19527 7073
rect 19539 3343 19551 7073
rect 19563 5815 19575 7073
rect 19611 4951 19623 7073
rect 19635 6103 19647 7073
rect 19659 4951 19671 7073
rect 19683 5071 19695 7073
rect 19755 5071 19767 7073
rect 19779 6199 19791 7073
rect 19827 6295 19839 7073
rect 19875 6271 19887 7073
rect 19899 3871 19911 7073
rect 19995 6271 20007 7073
rect 20019 6871 20031 7073
rect 19875 1807 19887 3809
rect 19899 1807 19911 3713
rect 19923 3607 19935 6257
rect 20043 5887 20055 7073
rect 20091 6295 20103 7073
rect 20115 6247 20127 7073
rect 20139 6391 20151 7073
rect 19947 1807 19959 4769
rect 19971 3727 19983 5873
rect 19995 1807 20007 4001
rect 20067 1807 20079 4385
rect 20091 1807 20103 5273
rect 20163 1807 20175 4793
rect 20187 3679 20199 7073
rect 20211 6343 20223 7073
rect 20187 1807 20199 3449
rect 20211 1807 20223 5681
rect 20235 3223 20247 7073
rect 20259 2887 20271 7073
rect 20283 3055 20295 6257
rect 20307 3319 20319 7073
rect 20307 1807 20319 3257
rect 20331 3175 20343 7073
rect 20379 6535 20391 7073
rect 20355 3079 20367 6281
rect 20379 1807 20391 2849
rect 20403 1807 20415 4721
rect 20427 2575 20439 7073
rect 20451 5911 20463 7073
rect 20463 3463 20475 5273
rect 20499 4975 20511 7073
rect 20499 1807 20511 3305
rect 20523 1807 20535 6017
rect 20547 3943 20559 7073
rect 20595 5767 20607 7073
rect 20571 3271 20583 5513
rect 20643 5311 20655 7073
rect 20667 4327 20679 6089
rect 20595 1807 20607 1865
rect 20619 1807 20631 3017
rect 20643 1807 20655 4313
rect 20691 1807 20703 6761
rect 20715 5407 20727 7073
rect 20739 5287 20751 7073
rect 20763 4735 20775 7073
rect 20811 3631 20823 7073
rect 20835 4975 20847 7073
rect 20859 3031 20871 7073
rect 20883 5407 20895 7073
rect 20715 1807 20727 2777
rect 20907 1807 20919 3017
rect 20931 1879 20943 7073
rect 20955 6055 20967 7073
rect 20931 1807 20943 1841
rect 20955 1807 20967 4001
rect 20979 1807 20991 5225
rect 21003 4999 21015 7073
rect 21051 6559 21063 7073
rect 21027 1807 21039 6497
rect 21051 1807 21063 3665
rect 21075 3199 21087 7073
rect 21099 6319 21111 7073
rect 21075 1807 21087 3137
rect 21123 1807 21135 5369
rect 21147 3655 21159 7073
rect 21147 1807 21159 3185
rect 21171 2359 21183 7073
rect 21195 5527 21207 7073
rect 21219 6199 21231 7073
rect 21267 5647 21279 7073
rect 21291 5095 21303 7073
rect 21195 1807 21207 4313
rect 21243 1807 21255 3617
rect 21267 1807 21279 4289
rect 21291 1807 21303 5009
rect 21315 4999 21327 7073
rect 21435 6271 21447 7073
rect 21351 3151 21363 4889
rect 21315 1807 21327 3017
rect 21339 1807 21351 2969
rect 21387 1807 21399 4673
rect 21411 1807 21423 3305
rect 21435 1807 21447 6209
rect 21459 1855 21471 5417
rect 21483 1807 21495 2897
rect 21507 1807 21519 4097
rect 21531 1807 21543 6449
rect 21555 4327 21567 6329
rect 21579 1807 21591 4961
rect 21603 1807 21615 4361
rect 21627 1807 21639 4313
rect 21651 4303 21663 6137
rect 21675 1807 21687 5393
rect 21699 2215 21711 6257
rect 21723 1807 21735 3689
rect 21747 1807 21759 2177
rect 21771 1807 21783 4265
rect 21795 4063 21807 7073
rect 21843 6199 21855 7073
rect 21987 6343 21999 7073
rect 21819 1807 21831 5297
rect 21843 1807 21855 6137
rect 21879 3799 21891 6185
rect 21867 1807 21879 2561
rect 21915 1807 21927 5825
rect 21939 1807 21951 5465
rect 21963 1807 21975 5033
rect 22011 4447 22023 7073
rect 22035 4951 22047 7073
rect 22011 1807 22023 3617
rect 22059 1807 22071 4505
rect 22083 4375 22095 7073
rect 22107 3967 22119 7073
rect 22131 1807 22143 6065
rect 22155 4903 22167 7073
rect 22203 4951 22215 7073
rect 22251 5335 22263 7073
rect 22275 5095 22287 7073
rect 22227 1807 22239 4241
rect 22275 1807 22287 4289
rect 22299 4039 22311 7073
rect 22323 4303 22335 5969
rect 22347 5287 22359 7073
rect 22371 2359 22383 7073
rect 22395 4039 22407 7073
rect 22419 5071 22431 7073
rect 22467 5335 22479 7073
rect 22491 5527 22503 7073
rect 22431 3943 22443 4577
rect 22371 1807 22383 2321
rect 22395 1807 22407 3929
rect 22419 1807 22431 3233
rect 22467 1807 22479 4889
rect 22515 4711 22527 7073
rect 22563 4831 22575 7073
rect 22539 2335 22551 4769
rect 22587 1807 22599 5945
rect 22611 4375 22623 7073
rect 22647 4303 22659 6065
rect 22611 1807 22623 4289
rect 22635 1807 22647 4145
rect 22683 2815 22695 7073
rect 22707 5551 22719 7073
rect 22755 6727 22767 7073
rect 22683 1807 22695 2777
rect 22707 1807 22719 4001
rect 22731 1807 22743 5585
rect 22803 4399 22815 7073
rect 22827 4375 22839 7073
rect 22851 5191 22863 7073
rect 22779 1807 22791 3737
rect 22827 1807 22839 4289
rect 22875 1807 22887 6665
rect 22899 2407 22911 7073
rect 22923 2479 22935 7073
rect 22947 2551 22959 7073
rect 22971 3967 22983 7073
rect 22995 5263 23007 7073
rect 23007 4303 23019 5201
rect 22899 1807 22911 2321
rect 22995 1807 23007 3569
rect 23019 2791 23031 3521
rect 23043 3319 23055 7073
rect 23067 4111 23079 7073
rect 23091 4519 23103 7073
rect 23067 1807 23079 4049
rect 23091 1807 23103 4121
rect 23115 1999 23127 7073
rect 23139 4063 23151 5849
rect 23163 4735 23175 7073
rect 23187 4879 23199 7073
rect 23211 6007 23223 7073
rect 23235 5047 23247 7073
rect 23259 6727 23271 7073
rect 23139 2335 23151 3785
rect 23163 1807 23175 3545
rect 23259 1807 23271 6593
rect 23307 6535 23319 7073
rect 23331 6511 23343 7073
rect 23307 1807 23319 5153
rect 23355 1903 23367 7073
rect 23403 5167 23415 7073
rect 23451 5839 23463 7073
rect 23523 5311 23535 7073
rect 23379 1807 23391 4649
rect 23403 1807 23415 5081
rect 23487 2935 23499 5153
rect 23547 4519 23559 7073
rect 23571 4303 23583 6617
rect 23595 6175 23607 7073
rect 23427 1807 23439 2753
rect 23475 1807 23487 2081
rect 23523 1807 23535 4289
rect 23595 1807 23607 3593
rect 23643 3511 23655 7073
rect 23667 4207 23679 7073
rect 23691 5359 23703 7073
rect 23715 4855 23727 7073
rect 23787 6127 23799 7073
rect 23835 5143 23847 7073
rect 23619 1807 23631 3017
rect 23691 1807 23703 4121
rect 23811 1807 23823 3905
rect 23859 1807 23871 6473
rect 23907 4855 23919 7073
rect 23931 7063 23943 7073
rect 23931 1807 23943 6953
rect 23955 4543 23967 7073
rect 24027 4807 24039 7073
rect 24051 4687 24063 7073
rect 24075 1807 24087 5417
rect 24099 1807 24111 4001
rect 24123 1807 24135 7001
rect 24147 6655 24159 7073
rect 24171 3223 24183 7073
rect 24195 3847 24207 7073
rect 24243 6679 24255 7073
rect 24171 1807 24183 2009
rect 24243 1807 24255 5609
rect 24267 2719 24279 7073
rect 24291 7039 24303 7073
rect 24315 1807 24327 6785
rect 24339 5527 24351 7073
rect 24363 5551 24375 7073
rect 24387 4423 24399 7073
rect 24435 6991 24447 7073
rect 24459 5911 24471 7073
rect 24459 1807 24471 5801
rect 24483 4495 24495 7073
rect 24531 6391 24543 7073
rect 24555 2407 24567 7073
rect 24579 5575 24591 7073
rect 24603 5719 24615 7073
rect 24651 3295 24663 7073
rect 24699 2623 24711 7073
rect 24771 2551 24783 7073
rect 24795 2071 24807 7073
rect 24819 2671 24831 7073
rect 24867 4495 24879 7073
rect 24867 1807 24879 3953
rect 24891 3175 24903 4481
rect 24915 3823 24927 7073
rect 24987 6871 24999 7073
rect 25011 6751 25023 7073
rect 25059 6247 25071 7073
rect 25107 5863 25119 7073
rect 25011 1807 25023 5369
rect 25131 4687 25143 7073
rect 25155 5911 25167 7073
rect 25203 5839 25215 7073
rect 25059 1807 25071 2369
rect 25155 1807 25167 4937
rect 25227 4375 25239 7073
rect 25251 4927 25263 7073
rect 25299 3919 25311 7073
rect 25323 4567 25335 7073
rect 25347 6367 25359 7073
rect 25395 6703 25407 7073
rect 25467 5623 25479 7073
rect 25539 4087 25551 7073
rect 25611 3655 25623 7073
rect 25635 6343 25647 7073
rect 25659 3823 25671 7073
rect 25683 4759 25695 7073
rect 25731 5503 25743 7073
rect 25203 1807 25215 3209
rect 25731 1807 25743 5273
rect 25755 3775 25767 7073
rect 25779 5791 25791 7073
rect 25827 5959 25839 7073
rect 25875 4399 25887 7073
rect 25779 1807 25791 3617
rect 25923 1807 25935 4169
rect 25947 3967 25959 7073
rect 25971 5287 25983 7073
rect 26019 5455 26031 7073
rect 26067 6727 26079 7073
rect 26139 7063 26151 7073
rect 26187 5695 26199 7073
rect 25971 1807 25983 4961
rect 26091 1807 26103 4457
rect 26163 1807 26175 4121
rect 26187 1807 26199 5657
rect 26211 3631 26223 7073
rect 26235 6847 26247 7073
rect 26283 3655 26295 7073
rect 26307 4015 26319 7073
rect 26355 6439 26367 7073
rect 26259 1807 26271 2945
rect 26283 1807 26295 3617
rect 26331 2695 26343 5681
rect 26355 1807 26367 6401
rect 26403 5023 26415 7073
rect 26379 1807 26391 3473
rect 26403 1807 26415 4625
rect 26427 3391 26439 7073
rect 26451 5503 26463 7073
rect 26451 1807 26463 5465
rect 26475 3631 26487 5873
rect 26499 3991 26511 7073
rect 26523 2959 26535 7073
rect 26547 5119 26559 7073
rect 26571 4615 26583 7073
rect 26595 4447 26607 6425
rect 26619 3319 26631 7073
rect 26643 4015 26655 7073
rect 26691 5743 26703 7073
rect 26739 5935 26751 7073
rect 26499 1807 26511 2393
rect 26667 2119 26679 5489
rect 26763 4999 26775 7073
rect 26787 4327 26799 7073
rect 26811 3367 26823 7073
rect 26859 3751 26871 7073
rect 26883 4111 26895 7073
rect 26931 2359 26943 7073
rect 26979 3991 26991 7073
rect 27003 3967 27015 7073
rect 27051 6559 27063 7073
rect 27099 4351 27111 7073
rect 27099 1903 27111 4073
rect 27123 1831 27135 5537
rect 27147 1855 27159 5081
rect 27171 1879 27183 6401
rect 27195 1927 27207 2129
rect 27219 1951 27231 6785
rect 27243 1807 27443 7073
rect 27579 1962 27649 1974
rect 27579 1938 27649 1950
rect 27579 1914 27649 1926
rect 27579 1890 27649 1902
rect 27579 1866 27649 1878
rect 27579 1842 27649 1854
rect 27579 1818 27649 1830
rect 0 121 70 133
rect 0 97 70 109
rect 0 73 70 85
rect 0 49 70 61
rect 124 0 324 1008
rect 339 0 351 1008
rect 363 0 375 1008
rect 387 0 399 1008
rect 411 0 423 1008
rect 2235 62 2247 1008
rect 2331 62 2343 1008
rect 2379 158 2391 1008
rect 2451 182 2463 1008
rect 2643 110 2655 1008
rect 2667 206 2679 1008
rect 2715 110 2727 1008
rect 3483 230 3495 1008
rect 3603 134 3615 1008
rect 3699 134 3711 1008
rect 3867 254 3879 1008
rect 4155 278 4167 1008
rect 4203 302 4215 1008
rect 4299 326 4311 1008
rect 4491 350 4503 1008
rect 4563 206 4575 1008
rect 4587 374 4599 1008
rect 4683 254 4695 1008
rect 4731 206 4743 1008
rect 5019 398 5031 1008
rect 5235 422 5247 1008
rect 5355 38 5367 1008
rect 5475 446 5487 1008
rect 5499 470 5511 1008
rect 5547 494 5559 1008
rect 5595 86 5607 1008
rect 6267 86 6279 1008
rect 6459 518 6471 1008
rect 6483 542 6495 1008
rect 6555 566 6567 1008
rect 6603 446 6615 1008
rect 6675 446 6687 1008
rect 6699 590 6711 1008
rect 6771 614 6783 1008
rect 6795 638 6807 1008
rect 6819 662 6831 1008
rect 7011 398 7023 1008
rect 7035 686 7047 1008
rect 7299 710 7311 1008
rect 7539 734 7551 1008
rect 7827 398 7839 1008
rect 7971 758 7983 1008
rect 7995 782 8007 1008
rect 8187 254 8199 1008
rect 8211 806 8223 1008
rect 8379 830 8391 1008
rect 8499 854 8511 1008
rect 8643 134 8655 1008
rect 8811 758 8823 1008
rect 8859 134 8871 1008
rect 8883 86 8895 1008
rect 8931 86 8943 1008
rect 8979 518 8991 1008
rect 9099 662 9111 1008
rect 9699 518 9711 1008
rect 9795 662 9807 1008
rect 9963 14 9975 1008
rect 10035 878 10047 1008
rect 10467 758 10479 1008
rect 10755 710 10767 1008
rect 10851 878 10863 1008
rect 10923 518 10935 1008
rect 11091 710 11103 1008
rect 11283 134 11295 1008
rect 11691 902 11703 1008
rect 11787 710 11799 1008
rect 11811 926 11823 1008
rect 11907 758 11919 1008
rect 12099 710 12111 1008
rect 12243 950 12255 1008
rect 12387 974 12399 1008
rect 12579 998 12591 1008
rect 12843 446 12855 1008
rect 12915 350 12927 1008
rect 12939 182 12951 1008
rect 13443 350 13455 1008
rect 13467 230 13479 1008
rect 13611 326 13623 1008
rect 13659 326 13671 1008
rect 13683 230 13695 1008
rect 13707 278 13719 1008
rect 13755 782 13767 1008
rect 13779 182 13791 1008
rect 13803 86 13815 1008
rect 14019 230 14031 1008
rect 14091 758 14103 1008
rect 14115 158 14127 1008
rect 14211 782 14223 1008
rect 14355 398 14367 1008
rect 14475 278 14487 1008
rect 14499 230 14511 1008
rect 14523 614 14535 1008
rect 15411 278 15423 1008
rect 15603 806 15615 1008
rect 15843 662 15855 1008
rect 15891 614 15903 1008
rect 15987 278 15999 1008
rect 16083 542 16095 1008
rect 16131 758 16143 1008
rect 16251 950 16263 1008
rect 16371 374 16383 1008
rect 16467 734 16479 1008
rect 16707 686 16719 1008
rect 16731 758 16743 1008
rect 16803 542 16815 1008
rect 16995 974 17007 1008
rect 17163 686 17175 1008
rect 17523 734 17535 1008
rect 17571 230 17583 1008
rect 17715 302 17727 1008
rect 17859 494 17871 1008
rect 18075 806 18087 1008
rect 18267 806 18279 1008
rect 19035 206 19047 1008
rect 19083 950 19095 1008
rect 19179 830 19191 1008
rect 19707 686 19719 1008
rect 19851 590 19863 1008
rect 20115 830 20127 1008
rect 20259 254 20271 1008
rect 20451 710 20463 1008
rect 20547 926 20559 1008
rect 20763 710 20775 1008
rect 20811 686 20823 1008
rect 20835 734 20847 1008
rect 20859 638 20871 1008
rect 21699 710 21711 1008
rect 22035 662 22047 1008
rect 22083 998 22095 1008
rect 22155 614 22167 1008
rect 22179 830 22191 1008
rect 22203 278 22215 1008
rect 22299 398 22311 1008
rect 22323 542 22335 1008
rect 22491 542 22503 1008
rect 22539 470 22551 1008
rect 22803 398 22815 1008
rect 22923 854 22935 1008
rect 22971 614 22983 1008
rect 23019 806 23031 1008
rect 23115 614 23127 1008
rect 23187 62 23199 1008
rect 23211 422 23223 1008
rect 23283 398 23295 1008
rect 23355 758 23367 1008
rect 23643 110 23655 1008
rect 23715 878 23727 1008
rect 23763 542 23775 1008
rect 23955 950 23967 1008
rect 24003 326 24015 1008
rect 24051 206 24063 1008
rect 25035 590 25047 1008
rect 25107 110 25119 1008
rect 25131 782 25143 1008
rect 25227 134 25239 1008
rect 25251 446 25263 1008
rect 25371 902 25383 1008
rect 26043 518 26055 1008
rect 26211 350 26223 1008
rect 26307 566 26319 1008
rect 26307 62 26319 384
rect 26331 86 26343 744
rect 26355 110 26367 240
rect 26379 38 26391 144
rect 26403 38 26415 120
rect 27243 0 27443 1008
rect 27579 145 27649 157
rect 27579 97 27649 109
rect 27579 73 27649 85
rect 27579 49 27649 61
rect 27579 25 27649 37
rect 27579 1 27649 13
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7073
box 0 0 1464 799
use inv g8182
timestamp 1386238110
transform 1 0 1587 0 1 7073
box 0 0 120 799
use rowcrosser Rs1Sel_91_0_93_
timestamp 1386086759
transform 1 0 1707 0 1 7073
box 0 0 48 799
use nand2 g8369
timestamp 1386234792
transform 1 0 1755 0 1 7073
box 0 0 96 799
use nor2 g8462
timestamp 1386235306
transform 1 0 1851 0 1 7073
box 0 0 120 799
use inv g8169
timestamp 1386238110
transform 1 0 1971 0 1 7073
box 0 0 120 799
use nand2 g8107
timestamp 1386234792
transform 1 0 2091 0 1 7073
box 0 0 96 799
use nand4 g8229
timestamp 1386234936
transform 1 0 2187 0 1 7073
box 0 0 144 799
use inv g8370
timestamp 1386238110
transform 1 0 2331 0 1 7073
box 0 0 120 799
use nand2 g8313
timestamp 1386234792
transform 1 0 2451 0 1 7073
box 0 0 96 799
use nand2 g8344
timestamp 1386234792
transform 1 0 2547 0 1 7073
box 0 0 96 799
use nand2 g8123
timestamp 1386234792
transform 1 0 2643 0 1 7073
box 0 0 96 799
use inv g8222
timestamp 1386238110
transform 1 0 2739 0 1 7073
box 0 0 120 799
use rowcrosser PcSel_91_2_93_
timestamp 1386086759
transform 1 0 2859 0 1 7073
box 0 0 48 799
use and2 g8102
timestamp 1386234845
transform 1 0 2907 0 1 7073
box 0 0 120 799
use nand3 g8098
timestamp 1386234893
transform 1 0 3027 0 1 7073
box 0 0 120 799
use nand4 g8314
timestamp 1386234936
transform 1 0 3147 0 1 7073
box 0 0 144 799
use nand2 g8327
timestamp 1386234792
transform 1 0 3291 0 1 7073
box 0 0 96 799
use nor2 g8187
timestamp 1386235306
transform 1 0 3387 0 1 7073
box 0 0 120 799
use and2 g8171
timestamp 1386234845
transform 1 0 3507 0 1 7073
box 0 0 120 799
use nand2 g8135
timestamp 1386234792
transform 1 0 3627 0 1 7073
box 0 0 96 799
use inv g8295
timestamp 1386238110
transform 1 0 3723 0 1 7073
box 0 0 120 799
use nand2 g8287
timestamp 1386234792
transform 1 0 3843 0 1 7073
box 0 0 96 799
use nand2 g8154
timestamp 1386234792
transform 1 0 3939 0 1 7073
box 0 0 96 799
use nand2 g8276
timestamp 1386234792
transform 1 0 4035 0 1 7073
box 0 0 96 799
use nand2 g8261
timestamp 1386234792
transform 1 0 4131 0 1 7073
box 0 0 96 799
use nand2 g8130
timestamp 1386234792
transform 1 0 4227 0 1 7073
box 0 0 96 799
use nor2 g8318
timestamp 1386235306
transform 1 0 4323 0 1 7073
box 0 0 120 799
use nand3 g8377
timestamp 1386234893
transform 1 0 4443 0 1 7073
box 0 0 120 799
use nor2 g8474
timestamp 1386235306
transform 1 0 4563 0 1 7073
box 0 0 120 799
use inv g8390
timestamp 1386238110
transform 1 0 4683 0 1 7073
box 0 0 120 799
use nand3 g8168
timestamp 1386234893
transform 1 0 4803 0 1 7073
box 0 0 120 799
use nand2 g8238
timestamp 1386234792
transform 1 0 4923 0 1 7073
box 0 0 96 799
use inv g8225
timestamp 1386238110
transform 1 0 5019 0 1 7073
box 0 0 120 799
use nand2 g8143
timestamp 1386234792
transform 1 0 5139 0 1 7073
box 0 0 96 799
use nand2 g8333
timestamp 1386234792
transform 1 0 5235 0 1 7073
box 0 0 96 799
use nand2 g8472
timestamp 1386234792
transform 1 0 5331 0 1 7073
box 0 0 96 799
use inv g8149
timestamp 1386238110
transform 1 0 5427 0 1 7073
box 0 0 120 799
use nand2 g8338
timestamp 1386234792
transform 1 0 5547 0 1 7073
box 0 0 96 799
use and2 g8280
timestamp 1386234845
transform 1 0 5643 0 1 7073
box 0 0 120 799
use nand3 g8249
timestamp 1386234893
transform 1 0 5763 0 1 7073
box 0 0 120 799
use nand2 g8310
timestamp 1386234792
transform 1 0 5883 0 1 7073
box 0 0 96 799
use nand3 g8450
timestamp 1386234893
transform 1 0 5979 0 1 7073
box 0 0 120 799
use nand2 g8456
timestamp 1386234792
transform 1 0 6099 0 1 7073
box 0 0 96 799
use inv g8235
timestamp 1386238110
transform 1 0 6195 0 1 7073
box 0 0 120 799
use nand3 g8362
timestamp 1386234893
transform 1 0 6315 0 1 7073
box 0 0 120 799
use mux2 g8214
timestamp 1386235218
transform 1 0 6435 0 1 7073
box 0 0 192 799
use nor2 g8281
timestamp 1386235306
transform 1 0 6627 0 1 7073
box 0 0 120 799
use nand3 g8366
timestamp 1386234893
transform 1 0 6747 0 1 7073
box 0 0 120 799
use rowcrosser LrSel
timestamp 1386086759
transform 1 0 6867 0 1 7073
box 0 0 48 799
use nand2 g8269
timestamp 1386234792
transform 1 0 6915 0 1 7073
box 0 0 96 799
use nand2 g8440
timestamp 1386234792
transform 1 0 7011 0 1 7073
box 0 0 96 799
use and2 g8183
timestamp 1386234845
transform 1 0 7107 0 1 7073
box 0 0 120 799
use nand4 g8170
timestamp 1386234936
transform 1 0 7227 0 1 7073
box 0 0 144 799
use nand2 g8449
timestamp 1386234792
transform 1 0 7371 0 1 7073
box 0 0 96 799
use nand2 g8124
timestamp 1386234792
transform 1 0 7467 0 1 7073
box 0 0 96 799
use nand4 g8106
timestamp 1386234936
transform 1 0 7563 0 1 7073
box 0 0 144 799
use nand4 g8414
timestamp 1386234936
transform 1 0 7707 0 1 7073
box 0 0 144 799
use xor2 g8119
timestamp 1386237344
transform 1 0 7851 0 1 7073
box 0 0 192 799
use inv g8275
timestamp 1386238110
transform 1 0 8043 0 1 7073
box 0 0 120 799
use nand2 g8418
timestamp 1386234792
transform 1 0 8163 0 1 7073
box 0 0 96 799
use nor2 g8146
timestamp 1386235306
transform 1 0 8259 0 1 7073
box 0 0 120 799
use nand2 g477
timestamp 1386234792
transform 1 0 8379 0 1 7073
box 0 0 96 799
use trisbuf g8155
timestamp 1386237216
transform 1 0 8475 0 1 7073
box 0 0 216 799
use nand2 g8127
timestamp 1386234792
transform 1 0 8691 0 1 7073
box 0 0 96 799
use nand3 g8290
timestamp 1386234893
transform 1 0 8787 0 1 7073
box 0 0 120 799
use nand3 g8252
timestamp 1386234893
transform 1 0 8907 0 1 7073
box 0 0 120 799
use nand2 g8334
timestamp 1386234792
transform 1 0 9027 0 1 7073
box 0 0 96 799
use inv g8244
timestamp 1386238110
transform 1 0 9123 0 1 7073
box 0 0 120 799
use nor2 g8240
timestamp 1386235306
transform 1 0 9243 0 1 7073
box 0 0 120 799
use nand3 g8407
timestamp 1386234893
transform 1 0 9363 0 1 7073
box 0 0 120 799
use nand2 g8139
timestamp 1386234792
transform 1 0 9483 0 1 7073
box 0 0 96 799
use nor2 g8118
timestamp 1386235306
transform 1 0 9579 0 1 7073
box 0 0 120 799
use nand2 g8363
timestamp 1386234792
transform 1 0 9699 0 1 7073
box 0 0 96 799
use nand3 g8111
timestamp 1386234893
transform 1 0 9795 0 1 7073
box 0 0 120 799
use nand2 g8381
timestamp 1386234792
transform 1 0 9915 0 1 7073
box 0 0 96 799
use nand2 g8403
timestamp 1386234792
transform 1 0 10011 0 1 7073
box 0 0 96 799
use rowcrosser MemEn
timestamp 1386086759
transform 1 0 10107 0 1 7073
box 0 0 48 799
use nand2 g8357
timestamp 1386234792
transform 1 0 10155 0 1 7073
box 0 0 96 799
use and2 g8347
timestamp 1386234845
transform 1 0 10251 0 1 7073
box 0 0 120 799
use nand2 g8120
timestamp 1386234792
transform 1 0 10371 0 1 7073
box 0 0 96 799
use nand4 g8134
timestamp 1386234936
transform 1 0 10467 0 1 7073
box 0 0 144 799
use nand3 g8386
timestamp 1386234893
transform 1 0 10611 0 1 7073
box 0 0 120 799
use nand2 g8425
timestamp 1386234792
transform 1 0 10731 0 1 7073
box 0 0 96 799
use nor2 g8320
timestamp 1386235306
transform 1 0 10827 0 1 7073
box 0 0 120 799
use nand3 g8354
timestamp 1386234893
transform 1 0 10947 0 1 7073
box 0 0 120 799
use nand2 g8374
timestamp 1386234792
transform 1 0 11067 0 1 7073
box 0 0 96 799
use and2 g8218
timestamp 1386234845
transform 1 0 11163 0 1 7073
box 0 0 120 799
use nand2 g8284
timestamp 1386234792
transform 1 0 11283 0 1 7073
box 0 0 96 799
use nand3 g8198
timestamp 1386234893
transform 1 0 11379 0 1 7073
box 0 0 120 799
use nor2 g8272
timestamp 1386235306
transform 1 0 11499 0 1 7073
box 0 0 120 799
use nand2 g8199
timestamp 1386234792
transform 1 0 11619 0 1 7073
box 0 0 96 799
use and2 g8306
timestamp 1386234845
transform 1 0 11715 0 1 7073
box 0 0 120 799
use nand3 g8221
timestamp 1386234893
transform 1 0 11835 0 1 7073
box 0 0 120 799
use and2 g8319
timestamp 1386234845
transform 1 0 11955 0 1 7073
box 0 0 120 799
use nand4 g8220
timestamp 1386234936
transform 1 0 12075 0 1 7073
box 0 0 144 799
use nand3 g8392
timestamp 1386234893
transform 1 0 12219 0 1 7073
box 0 0 120 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 12339 0 1 7073
box 0 0 48 799
use and2 g8431
timestamp 1386234845
transform 1 0 12387 0 1 7073
box 0 0 120 799
use nand2 g8194
timestamp 1386234792
transform 1 0 12507 0 1 7073
box 0 0 96 799
use nand3 g8271
timestamp 1386234893
transform 1 0 12603 0 1 7073
box 0 0 120 799
use nand3 g8230
timestamp 1386234893
transform 1 0 12723 0 1 7073
box 0 0 120 799
use rowcrosser RegWe
timestamp 1386086759
transform 1 0 12843 0 1 7073
box 0 0 48 799
use nand4 g8340
timestamp 1386234936
transform 1 0 12891 0 1 7073
box 0 0 144 799
use nor2 g8399
timestamp 1386235306
transform 1 0 13035 0 1 7073
box 0 0 120 799
use nand2 g8421
timestamp 1386234792
transform 1 0 13155 0 1 7073
box 0 0 96 799
use inv g8209
timestamp 1386238110
transform 1 0 13251 0 1 7073
box 0 0 120 799
use and2 g8103
timestamp 1386234845
transform 1 0 13371 0 1 7073
box 0 0 120 799
use nand3 g8268
timestamp 1386234893
transform 1 0 13491 0 1 7073
box 0 0 120 799
use nand2 g8283
timestamp 1386234792
transform 1 0 13611 0 1 7073
box 0 0 96 799
use nand4 g8411
timestamp 1386234936
transform 1 0 13707 0 1 7073
box 0 0 144 799
use nand3 g8321
timestamp 1386234893
transform 1 0 13851 0 1 7073
box 0 0 120 799
use nand3 g8379
timestamp 1386234893
transform 1 0 13971 0 1 7073
box 0 0 120 799
use inv g8180
timestamp 1386238110
transform 1 0 14091 0 1 7073
box 0 0 120 799
use and2 g8417
timestamp 1386234845
transform 1 0 14211 0 1 7073
box 0 0 120 799
use nand2 g8136
timestamp 1386234792
transform 1 0 14331 0 1 7073
box 0 0 96 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 14427 0 1 7073
box 0 0 48 799
use nand4 g8110
timestamp 1386234936
transform 1 0 14475 0 1 7073
box 0 0 144 799
use nand2 g8153
timestamp 1386234792
transform 1 0 14619 0 1 7073
box 0 0 96 799
use nand2 g8361
timestamp 1386234792
transform 1 0 14715 0 1 7073
box 0 0 96 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 14811 0 1 7073
box 0 0 96 799
use scandtype g8308
timestamp 1386241841
transform 1 0 14907 0 1 7073
box 0 0 624 799
use nand2 stateSub_reg_91_2_93_
timestamp 1386234792
transform 1 0 15531 0 1 7073
box 0 0 96 799
use scandtype g8372
timestamp 1386241841
transform 1 0 15627 0 1 7073
box 0 0 624 799
use nand2 g8294
timestamp 1386234792
transform 1 0 16251 0 1 7073
box 0 0 96 799
use nand3 g8444
timestamp 1386234893
transform 1 0 16347 0 1 7073
box 0 0 120 799
use nand2 g8099
timestamp 1386234792
transform 1 0 16467 0 1 7073
box 0 0 96 799
use nand3 g8433
timestamp 1386234893
transform 1 0 16563 0 1 7073
box 0 0 120 799
use nand2 g8420
timestamp 1386234792
transform 1 0 16683 0 1 7073
box 0 0 96 799
use nand2 g8190
timestamp 1386234792
transform 1 0 16779 0 1 7073
box 0 0 96 799
use nand2 g8304
timestamp 1386234792
transform 1 0 16875 0 1 7073
box 0 0 96 799
use inv g8277
timestamp 1386238110
transform 1 0 16971 0 1 7073
box 0 0 120 799
use nand3 g8243
timestamp 1386234893
transform 1 0 17091 0 1 7073
box 0 0 120 799
use inv g8296
timestamp 1386238110
transform 1 0 17211 0 1 7073
box 0 0 120 799
use and2 g8348
timestamp 1386234845
transform 1 0 17331 0 1 7073
box 0 0 120 799
use nand2 g8234
timestamp 1386234792
transform 1 0 17451 0 1 7073
box 0 0 96 799
use nand3 StatusReg_reg_91_1_93_
timestamp 1386234893
transform 1 0 17547 0 1 7073
box 0 0 120 799
use scandtype g8324
timestamp 1386241841
transform 1 0 17667 0 1 7073
box 0 0 624 799
use rowcrosser stateSub_reg_91_0_93_
timestamp 1386086759
transform 1 0 18291 0 1 7073
box 0 0 48 799
use rowcrosser Op2Sel_91_0_93_
timestamp 1386086759
transform 1 0 18339 0 1 7073
box 0 0 48 799
use nand2 g8293
timestamp 1386234792
transform 1 0 18387 0 1 7073
box 0 0 96 799
use nand2 g8435
timestamp 1386234792
transform 1 0 18483 0 1 7073
box 0 0 96 799
use nand2 g8452
timestamp 1386234792
transform 1 0 18579 0 1 7073
box 0 0 96 799
use inv g8312
timestamp 1386238110
transform 1 0 18675 0 1 7073
box 0 0 120 799
use and2 g8213
timestamp 1386234845
transform 1 0 18795 0 1 7073
box 0 0 120 799
use inv g8212
timestamp 1386238110
transform 1 0 18915 0 1 7073
box 0 0 120 799
use nor2 g8265
timestamp 1386235306
transform 1 0 19035 0 1 7073
box 0 0 120 799
use nand2 g8200
timestamp 1386234792
transform 1 0 19155 0 1 7073
box 0 0 96 799
use nand2 g8400
timestamp 1386234792
transform 1 0 19251 0 1 7073
box 0 0 96 799
use nand2 g8108
timestamp 1386234792
transform 1 0 19347 0 1 7073
box 0 0 96 799
use nand4 g8159
timestamp 1386234936
transform 1 0 19443 0 1 7073
box 0 0 144 799
use nand4 g8144
timestamp 1386234936
transform 1 0 19587 0 1 7073
box 0 0 144 799
use and2 g8177
timestamp 1386234845
transform 1 0 19731 0 1 7073
box 0 0 120 799
use and2 g8356
timestamp 1386234845
transform 1 0 19851 0 1 7073
box 0 0 120 799
use nand2 g8251
timestamp 1386234792
transform 1 0 19971 0 1 7073
box 0 0 96 799
use nand2 g8226
timestamp 1386234792
transform 1 0 20067 0 1 7073
box 0 0 96 799
use nand3 g8436
timestamp 1386234893
transform 1 0 20163 0 1 7073
box 0 0 120 799
use nor2 g8264
timestamp 1386235306
transform 1 0 20283 0 1 7073
box 0 0 120 799
use nor2 g8332
timestamp 1386235306
transform 1 0 20403 0 1 7073
box 0 0 120 799
use rowcrosser LrWe
timestamp 1386086759
transform 1 0 20523 0 1 7073
box 0 0 48 799
use inv g8206
timestamp 1386238110
transform 1 0 20571 0 1 7073
box 0 0 120 799
use nand2 g8237
timestamp 1386234792
transform 1 0 20691 0 1 7073
box 0 0 96 799
use nand3 g8278
timestamp 1386234893
transform 1 0 20787 0 1 7073
box 0 0 120 799
use and2 g8376
timestamp 1386234845
transform 1 0 20907 0 1 7073
box 0 0 120 799
use nand2 g8181
timestamp 1386234792
transform 1 0 21027 0 1 7073
box 0 0 96 799
use nand3 g8216
timestamp 1386234893
transform 1 0 21123 0 1 7073
box 0 0 120 799
use nand2 StatusReg_reg_91_0_93_
timestamp 1386234792
transform 1 0 21243 0 1 7073
box 0 0 96 799
use scandtype g8253
timestamp 1386241841
transform 1 0 21339 0 1 7073
box 0 0 624 799
use nand2 g8373
timestamp 1386234792
transform 1 0 21963 0 1 7073
box 0 0 96 799
use nor2 g8443
timestamp 1386235306
transform 1 0 22059 0 1 7073
box 0 0 120 799
use rowcrosser nWait
timestamp 1386086759
transform 1 0 22179 0 1 7073
box 0 0 48 799
use nand2 g8186
timestamp 1386234792
transform 1 0 22227 0 1 7073
box 0 0 96 799
use nand3 g8427
timestamp 1386234893
transform 1 0 22323 0 1 7073
box 0 0 120 799
use nand2 g8432
timestamp 1386234792
transform 1 0 22443 0 1 7073
box 0 0 96 799
use inv g8424
timestamp 1386238110
transform 1 0 22539 0 1 7073
box 0 0 120 799
use nor2 g8223
timestamp 1386235306
transform 1 0 22659 0 1 7073
box 0 0 120 799
use nand2 g8195
timestamp 1386234792
transform 1 0 22779 0 1 7073
box 0 0 96 799
use nand4 g8410
timestamp 1386234936
transform 1 0 22875 0 1 7073
box 0 0 144 799
use nand3 g8133
timestamp 1386234893
transform 1 0 23019 0 1 7073
box 0 0 120 799
use nand4 g8341
timestamp 1386234936
transform 1 0 23139 0 1 7073
box 0 0 144 799
use nand2 g8406
timestamp 1386234792
transform 1 0 23283 0 1 7073
box 0 0 96 799
use inv g8289
timestamp 1386238110
transform 1 0 23379 0 1 7073
box 0 0 120 799
use and2 g8128
timestamp 1386234845
transform 1 0 23499 0 1 7073
box 0 0 120 799
use nand4 g8397
timestamp 1386234936
transform 1 0 23619 0 1 7073
box 0 0 144 799
use inv g8100
timestamp 1386238110
transform 1 0 23763 0 1 7073
box 0 0 120 799
use nand3 g8350
timestamp 1386234893
transform 1 0 23883 0 1 7073
box 0 0 120 799
use and2 g8167
timestamp 1386234845
transform 1 0 24003 0 1 7073
box 0 0 120 799
use nand2 g8117
timestamp 1386234792
transform 1 0 24123 0 1 7073
box 0 0 96 799
use nand2 g8439
timestamp 1386234792
transform 1 0 24219 0 1 7073
box 0 0 96 799
use nand2 g8227
timestamp 1386234792
transform 1 0 24315 0 1 7073
box 0 0 96 799
use nand2 g8191
timestamp 1386234792
transform 1 0 24411 0 1 7073
box 0 0 96 799
use nand3 g8387
timestamp 1386234893
transform 1 0 24507 0 1 7073
box 0 0 120 799
use inv g8270
timestamp 1386238110
transform 1 0 24627 0 1 7073
box 0 0 120 799
use nand2 g8465
timestamp 1386234792
transform 1 0 24747 0 1 7073
box 0 0 96 799
use inv g8455
timestamp 1386238110
transform 1 0 24843 0 1 7073
box 0 0 120 799
use and2 g8273
timestamp 1386234845
transform 1 0 24963 0 1 7073
box 0 0 120 799
use nand2 g8337
timestamp 1386234792
transform 1 0 25083 0 1 7073
box 0 0 96 799
use nand2 g8147
timestamp 1386234792
transform 1 0 25179 0 1 7073
box 0 0 96 799
use nand2 g1
timestamp 1386234792
transform 1 0 25275 0 1 7073
box 0 0 96 799
use trisbuf g8217
timestamp 1386237216
transform 1 0 25371 0 1 7073
box 0 0 216 799
use nand3 g8353
timestamp 1386234893
transform 1 0 25587 0 1 7073
box 0 0 120 799
use nand2 g8248
timestamp 1386234792
transform 1 0 25707 0 1 7073
box 0 0 96 799
use inv g8447
timestamp 1386238110
transform 1 0 25803 0 1 7073
box 0 0 120 799
use nor2 g8114
timestamp 1386235306
transform 1 0 25923 0 1 7073
box 0 0 120 799
use nor2 g8174
timestamp 1386235306
transform 1 0 26043 0 1 7073
box 0 0 120 799
use nand2 g8393
timestamp 1386234792
transform 1 0 26163 0 1 7073
box 0 0 96 799
use and2 g8305
timestamp 1386234845
transform 1 0 26259 0 1 7073
box 0 0 120 799
use nand2 g8241
timestamp 1386234792
transform 1 0 26379 0 1 7073
box 0 0 96 799
use nand3 g8382
timestamp 1386234893
transform 1 0 26475 0 1 7073
box 0 0 120 799
use and2 g8158
timestamp 1386234845
transform 1 0 26595 0 1 7073
box 0 0 120 799
use nand3 g8257
timestamp 1386234893
transform 1 0 26715 0 1 7073
box 0 0 120 799
use and2 g8451
timestamp 1386234845
transform 1 0 26835 0 1 7073
box 0 0 120 799
use and2 RwSel_91_0_93_
timestamp 1386234845
transform 1 0 26955 0 1 7073
box 0 0 120 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 27075 0 1 7073
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27123 0 1 7073
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 1008
box 0 0 1464 799
use scandtype g8409
timestamp 1386241841
transform 1 0 1587 0 1 1008
box 0 0 624 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 2211 0 1 1008
box 0 0 48 799
use nand2 g8352
timestamp 1386234792
transform 1 0 2259 0 1 1008
box 0 0 96 799
use and2 g8430
timestamp 1386234845
transform 1 0 2355 0 1 1008
box 0 0 120 799
use nor2 g8150
timestamp 1386235306
transform 1 0 2475 0 1 1008
box 0 0 120 799
use nand2 g8178
timestamp 1386234792
transform 1 0 2595 0 1 1008
box 0 0 96 799
use inv state_reg_91_1_93_
timestamp 1386238110
transform 1 0 2691 0 1 1008
box 0 0 120 799
use scandtype g8250
timestamp 1386241841
transform 1 0 2811 0 1 1008
box 0 0 624 799
use and2 g8148
timestamp 1386234845
transform 1 0 3435 0 1 1008
box 0 0 120 799
use nand2 g8434
timestamp 1386234792
transform 1 0 3555 0 1 1008
box 0 0 96 799
use and2 g8196
timestamp 1386234845
transform 1 0 3651 0 1 1008
box 0 0 120 799
use nand4 g8211
timestamp 1386234936
transform 1 0 3771 0 1 1008
box 0 0 144 799
use nand2 g8300
timestamp 1386234792
transform 1 0 3915 0 1 1008
box 0 0 96 799
use inv g8175
timestamp 1386238110
transform 1 0 4011 0 1 1008
box 0 0 120 799
use nand2 g8359
timestamp 1386234792
transform 1 0 4131 0 1 1008
box 0 0 96 799
use nand2 g8388
timestamp 1386234792
transform 1 0 4227 0 1 1008
box 0 0 96 799
use nand2 g8429
timestamp 1386234792
transform 1 0 4323 0 1 1008
box 0 0 96 799
use nand2 g8104
timestamp 1386234792
transform 1 0 4419 0 1 1008
box 0 0 96 799
use nand3 g8391
timestamp 1386234893
transform 1 0 4515 0 1 1008
box 0 0 120 799
use and2 g8307
timestamp 1386234845
transform 1 0 4635 0 1 1008
box 0 0 120 799
use nand2 g8389
timestamp 1386234792
transform 1 0 4755 0 1 1008
box 0 0 96 799
use inv g8458
timestamp 1386238110
transform 1 0 4851 0 1 1008
box 0 0 120 799
use and2 g8335
timestamp 1386234845
transform 1 0 4971 0 1 1008
box 0 0 120 799
use nor2 g8160
timestamp 1386235306
transform 1 0 5091 0 1 1008
box 0 0 120 799
use nand3 g8476
timestamp 1386234893
transform 1 0 5211 0 1 1008
box 0 0 120 799
use inv g8224
timestamp 1386238110
transform 1 0 5331 0 1 1008
box 0 0 120 799
use and2 StatusReg_reg_91_2_93_
timestamp 1386234845
transform 1 0 5451 0 1 1008
box 0 0 120 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 5571 0 1 1008
box 0 0 48 799
use scandtype g8161
timestamp 1386241841
transform 1 0 5619 0 1 1008
box 0 0 624 799
use nand4 g8121
timestamp 1386234936
transform 1 0 6243 0 1 1008
box 0 0 144 799
use nand4 g8266
timestamp 1386234936
transform 1 0 6387 0 1 1008
box 0 0 144 799
use nand2 g8401
timestamp 1386234792
transform 1 0 6531 0 1 1008
box 0 0 96 799
use nand2 g8189
timestamp 1386234792
transform 1 0 6627 0 1 1008
box 0 0 96 799
use nand3 g8442
timestamp 1386234893
transform 1 0 6723 0 1 1008
box 0 0 120 799
use inv g8454
timestamp 1386238110
transform 1 0 6843 0 1 1008
box 0 0 120 799
use nand2 g8297
timestamp 1386234792
transform 1 0 6963 0 1 1008
box 0 0 96 799
use inv g8232
timestamp 1386238110
transform 1 0 7059 0 1 1008
box 0 0 120 799
use nand2 g8152
timestamp 1386234792
transform 1 0 7179 0 1 1008
box 0 0 96 799
use nand2 g8328
timestamp 1386234792
transform 1 0 7275 0 1 1008
box 0 0 96 799
use nor2 g8303
timestamp 1386235306
transform 1 0 7371 0 1 1008
box 0 0 120 799
use nand2 g8394
timestamp 1386234792
transform 1 0 7491 0 1 1008
box 0 0 96 799
use nand2 g8395
timestamp 1386234792
transform 1 0 7587 0 1 1008
box 0 0 96 799
use and2 g8453
timestamp 1386234845
transform 1 0 7683 0 1 1008
box 0 0 120 799
use nand2 g8282
timestamp 1386234792
transform 1 0 7803 0 1 1008
box 0 0 96 799
use nand3 g8267
timestamp 1386234893
transform 1 0 7899 0 1 1008
box 0 0 120 799
use inv g8461
timestamp 1386238110
transform 1 0 8019 0 1 1008
box 0 0 120 799
use nand2 g8274
timestamp 1386234792
transform 1 0 8139 0 1 1008
box 0 0 96 799
use inv g8236
timestamp 1386238110
transform 1 0 8235 0 1 1008
box 0 0 120 799
use nand3 g8101
timestamp 1386234893
transform 1 0 8355 0 1 1008
box 0 0 120 799
use nand3 g8438
timestamp 1386234893
transform 1 0 8475 0 1 1008
box 0 0 120 799
use nand2 g8349
timestamp 1386234792
transform 1 0 8595 0 1 1008
box 0 0 96 799
use nand2 g8412
timestamp 1386234792
transform 1 0 8691 0 1 1008
box 0 0 96 799
use nand3 g8185
timestamp 1386234893
transform 1 0 8787 0 1 1008
box 0 0 120 799
use nand2 IntReq_reg
timestamp 1386234792
transform 1 0 8907 0 1 1008
box 0 0 96 799
use scandtype g8365
timestamp 1386241841
transform 1 0 9003 0 1 1008
box 0 0 624 799
use nand2 g8255
timestamp 1386234792
transform 1 0 9627 0 1 1008
box 0 0 96 799
use nand2 g8457
timestamp 1386234792
transform 1 0 9723 0 1 1008
box 0 0 96 799
use nand2 g8301
timestamp 1386234792
transform 1 0 9819 0 1 1008
box 0 0 96 799
use nand2 g8192
timestamp 1386234792
transform 1 0 9915 0 1 1008
box 0 0 96 799
use nand3 g8292
timestamp 1386234893
transform 1 0 10011 0 1 1008
box 0 0 120 799
use inv g8254
timestamp 1386238110
transform 1 0 10131 0 1 1008
box 0 0 120 799
use nand2 g8116
timestamp 1386234792
transform 1 0 10251 0 1 1008
box 0 0 96 799
use nand2 g8470
timestamp 1386234792
transform 1 0 10347 0 1 1008
box 0 0 96 799
use inv g8145
timestamp 1386238110
transform 1 0 10443 0 1 1008
box 0 0 120 799
use nand3 g8166
timestamp 1386234893
transform 1 0 10563 0 1 1008
box 0 0 120 799
use nand2 g8426
timestamp 1386234792
transform 1 0 10683 0 1 1008
box 0 0 96 799
use inv g8315
timestamp 1386238110
transform 1 0 10779 0 1 1008
box 0 0 120 799
use nand2 g8228
timestamp 1386234792
transform 1 0 10899 0 1 1008
box 0 0 96 799
use and2 g8342
timestamp 1386234845
transform 1 0 10995 0 1 1008
box 0 0 120 799
use and2 g8279
timestamp 1386234845
transform 1 0 11115 0 1 1008
box 0 0 120 799
use nand2 g8259
timestamp 1386234792
transform 1 0 11235 0 1 1008
box 0 0 96 799
use nand3 g8375
timestamp 1386234893
transform 1 0 11331 0 1 1008
box 0 0 120 799
use and2 g8122
timestamp 1386234845
transform 1 0 11451 0 1 1008
box 0 0 120 799
use nand4 g8129
timestamp 1386234936
transform 1 0 11571 0 1 1008
box 0 0 144 799
use nand4 g8446
timestamp 1386234936
transform 1 0 11715 0 1 1008
box 0 0 144 799
use nand2 g8459
timestamp 1386234792
transform 1 0 11859 0 1 1008
box 0 0 96 799
use nand2 g8097
timestamp 1386234792
transform 1 0 11955 0 1 1008
box 0 0 96 799
use nand4 g8247
timestamp 1386234936
transform 1 0 12051 0 1 1008
box 0 0 144 799
use nor2 g8263
timestamp 1386235306
transform 1 0 12195 0 1 1008
box 0 0 120 799
use nand2 g8256
timestamp 1386234792
transform 1 0 12315 0 1 1008
box 0 0 96 799
use nor2 g8131
timestamp 1386235306
transform 1 0 12411 0 1 1008
box 0 0 120 799
use nand3 g8345
timestamp 1386234893
transform 1 0 12531 0 1 1008
box 0 0 120 799
use nand2 g8322
timestamp 1386234792
transform 1 0 12651 0 1 1008
box 0 0 96 799
use nand4 g8286
timestamp 1386234936
transform 1 0 12747 0 1 1008
box 0 0 144 799
use nand2 g8201
timestamp 1386234792
transform 1 0 12891 0 1 1008
box 0 0 96 799
use nand2 g479
timestamp 1386234792
transform 1 0 12987 0 1 1008
box 0 0 96 799
use trisbuf g8437
timestamp 1386237216
transform 1 0 13083 0 1 1008
box 0 0 216 799
use nand2 g8331
timestamp 1386234792
transform 1 0 13299 0 1 1008
box 0 0 96 799
use nand2 g8336
timestamp 1386234792
transform 1 0 13395 0 1 1008
box 0 0 96 799
use nand2 g8242
timestamp 1386234792
transform 1 0 13491 0 1 1008
box 0 0 96 799
use nand4 g8207
timestamp 1386234936
transform 1 0 13587 0 1 1008
box 0 0 144 799
use nand2 g8423
timestamp 1386234792
transform 1 0 13731 0 1 1008
box 0 0 96 799
use inv g8383
timestamp 1386238110
transform 1 0 13827 0 1 1008
box 0 0 120 799
use nand2 g8405
timestamp 1386234792
transform 1 0 13947 0 1 1008
box 0 0 96 799
use nand2 g8173
timestamp 1386234792
transform 1 0 14043 0 1 1008
box 0 0 96 799
use nand2 g8398
timestamp 1386234792
transform 1 0 14139 0 1 1008
box 0 0 96 799
use nand2 g8464
timestamp 1386234792
transform 1 0 14235 0 1 1008
box 0 0 96 799
use inv g8325
timestamp 1386238110
transform 1 0 14331 0 1 1008
box 0 0 120 799
use nand2 g8157
timestamp 1386234792
transform 1 0 14451 0 1 1008
box 0 0 96 799
use inv g8140
timestamp 1386238110
transform 1 0 14547 0 1 1008
box 0 0 120 799
use nand2 g8141
timestamp 1386234792
transform 1 0 14667 0 1 1008
box 0 0 96 799
use nand2 g8210
timestamp 1386234792
transform 1 0 14763 0 1 1008
box 0 0 96 799
use nand2 InISR_reg
timestamp 1386234792
transform 1 0 14859 0 1 1008
box 0 0 96 799
use scandtype g8460
timestamp 1386241841
transform 1 0 14955 0 1 1008
box 0 0 624 799
use inv g8317
timestamp 1386238110
transform 1 0 15579 0 1 1008
box 0 0 120 799
use nand3 g8203
timestamp 1386234893
transform 1 0 15699 0 1 1008
box 0 0 120 799
use nand2 g8404
timestamp 1386234792
transform 1 0 15819 0 1 1008
box 0 0 96 799
use nand2 g8428
timestamp 1386234792
transform 1 0 15915 0 1 1008
box 0 0 96 799
use nand2 g8413
timestamp 1386234792
transform 1 0 16011 0 1 1008
box 0 0 96 799
use xor2 g8113
timestamp 1386237344
transform 1 0 16107 0 1 1008
box 0 0 192 799
use nand2 g8358
timestamp 1386234792
transform 1 0 16299 0 1 1008
box 0 0 96 799
use nand2 g8323
timestamp 1386234792
transform 1 0 16395 0 1 1008
box 0 0 96 799
use mux2 g8408
timestamp 1386235218
transform 1 0 16491 0 1 1008
box 0 0 192 799
use nand2 g8309
timestamp 1386234792
transform 1 0 16683 0 1 1008
box 0 0 96 799
use nand2 g8380
timestamp 1386234792
transform 1 0 16779 0 1 1008
box 0 0 96 799
use nand2 g8233
timestamp 1386234792
transform 1 0 16875 0 1 1008
box 0 0 96 799
use nand2 IRQ2_reg
timestamp 1386234792
transform 1 0 16971 0 1 1008
box 0 0 96 799
use scandtype g8151
timestamp 1386241841
transform 1 0 17067 0 1 1008
box 0 0 624 799
use nand2 g8138
timestamp 1386234792
transform 1 0 17691 0 1 1008
box 0 0 96 799
use nand4 g8402
timestamp 1386234936
transform 1 0 17787 0 1 1008
box 0 0 144 799
use nand2 g8188
timestamp 1386234792
transform 1 0 17931 0 1 1008
box 0 0 96 799
use and2 g8176
timestamp 1386234845
transform 1 0 18027 0 1 1008
box 0 0 120 799
use nand2 g8172
timestamp 1386234792
transform 1 0 18147 0 1 1008
box 0 0 96 799
use nand2 g8422
timestamp 1386234792
transform 1 0 18243 0 1 1008
box 0 0 96 799
use nand2 g8162
timestamp 1386234792
transform 1 0 18339 0 1 1008
box 0 0 96 799
use nand2 g8415
timestamp 1386234792
transform 1 0 18435 0 1 1008
box 0 0 96 799
use xor2 g8095
timestamp 1386237344
transform 1 0 18531 0 1 1008
box 0 0 192 799
use nand4 g8299
timestamp 1386234936
transform 1 0 18723 0 1 1008
box 0 0 144 799
use and2 g8326
timestamp 1386234845
transform 1 0 18867 0 1 1008
box 0 0 120 799
use and2 g8396
timestamp 1386234845
transform 1 0 18987 0 1 1008
box 0 0 120 799
use nand2 IRQ1_reg
timestamp 1386234792
transform 1 0 19107 0 1 1008
box 0 0 96 799
use scandtype g8329
timestamp 1386241841
transform 1 0 19203 0 1 1008
box 0 0 624 799
use nand2 g8419
timestamp 1386234792
transform 1 0 19827 0 1 1008
box 0 0 96 799
use inv g8205
timestamp 1386238110
transform 1 0 19923 0 1 1008
box 0 0 120 799
use nand2 g8339
timestamp 1386234792
transform 1 0 20043 0 1 1008
box 0 0 96 799
use nand2 g8463
timestamp 1386234792
transform 1 0 20139 0 1 1008
box 0 0 96 799
use inv g8164
timestamp 1386238110
transform 1 0 20235 0 1 1008
box 0 0 120 799
use and2 g8245
timestamp 1386234845
transform 1 0 20355 0 1 1008
box 0 0 120 799
use nand2 g8260
timestamp 1386234792
transform 1 0 20475 0 1 1008
box 0 0 96 799
use nand2 g8165
timestamp 1386234792
transform 1 0 20571 0 1 1008
box 0 0 96 799
use nor2 g8351
timestamp 1386235306
transform 1 0 20667 0 1 1008
box 0 0 120 799
use nand2 g8215
timestamp 1386234792
transform 1 0 20787 0 1 1008
box 0 0 96 799
use nand3 g8343
timestamp 1386234893
transform 1 0 20883 0 1 1008
box 0 0 120 799
use nand2 g8288
timestamp 1386234792
transform 1 0 21003 0 1 1008
box 0 0 96 799
use and2 g8239
timestamp 1386234845
transform 1 0 21099 0 1 1008
box 0 0 120 799
use nand4 g8384
timestamp 1386234936
transform 1 0 21219 0 1 1008
box 0 0 144 799
use nand2 g8311
timestamp 1386234792
transform 1 0 21363 0 1 1008
box 0 0 96 799
use nand2 g8262
timestamp 1386234792
transform 1 0 21459 0 1 1008
box 0 0 96 799
use nand2 g8109
timestamp 1386234792
transform 1 0 21555 0 1 1008
box 0 0 96 799
use nand4 g8298
timestamp 1386234936
transform 1 0 21651 0 1 1008
box 0 0 144 799
use nand2 g8346
timestamp 1386234792
transform 1 0 21795 0 1 1008
box 0 0 96 799
use nand2 g8184
timestamp 1386234792
transform 1 0 21891 0 1 1008
box 0 0 96 799
use nand3 g8132
timestamp 1386234893
transform 1 0 21987 0 1 1008
box 0 0 120 799
use nand4 g8355
timestamp 1386234936
transform 1 0 22107 0 1 1008
box 0 0 144 799
use nand2 g8385
timestamp 1386234792
transform 1 0 22251 0 1 1008
box 0 0 96 799
use nand2 g8330
timestamp 1386234792
transform 1 0 22347 0 1 1008
box 0 0 96 799
use nor2 g8219
timestamp 1386235306
transform 1 0 22443 0 1 1008
box 0 0 120 799
use nand2 g8360
timestamp 1386234792
transform 1 0 22563 0 1 1008
box 0 0 96 799
use nand2 g8258
timestamp 1386234792
transform 1 0 22659 0 1 1008
box 0 0 96 799
use nand2 g8115
timestamp 1386234792
transform 1 0 22755 0 1 1008
box 0 0 96 799
use nand2 g8202
timestamp 1386234792
transform 1 0 22851 0 1 1008
box 0 0 96 799
use nand2 g8246
timestamp 1386234792
transform 1 0 22947 0 1 1008
box 0 0 96 799
use nand2 g8208
timestamp 1386234792
transform 1 0 23043 0 1 1008
box 0 0 96 799
use nand2 g8231
timestamp 1386234792
transform 1 0 23139 0 1 1008
box 0 0 96 799
use nand2 g8156
timestamp 1386234792
transform 1 0 23235 0 1 1008
box 0 0 96 799
use nand3 g8467
timestamp 1386234893
transform 1 0 23331 0 1 1008
box 0 0 120 799
use inv g8179
timestamp 1386238110
transform 1 0 23451 0 1 1008
box 0 0 120 799
use nand2 g8371
timestamp 1386234792
transform 1 0 23571 0 1 1008
box 0 0 96 799
use nor2 g8193
timestamp 1386235306
transform 1 0 23667 0 1 1008
box 0 0 120 799
use inv g8285
timestamp 1386238110
transform 1 0 23787 0 1 1008
box 0 0 120 799
use nor2 g8204
timestamp 1386235306
transform 1 0 23907 0 1 1008
box 0 0 120 799
use nand3 g478
timestamp 1386234893
transform 1 0 24027 0 1 1008
box 0 0 120 799
use trisbuf state_reg_91_0_93_
timestamp 1386237216
transform 1 0 24147 0 1 1008
box 0 0 216 799
use scandtype g8302
timestamp 1386241841
transform 1 0 24363 0 1 1008
box 0 0 624 799
use nand2 g8142
timestamp 1386234792
transform 1 0 24987 0 1 1008
box 0 0 96 799
use nand2 g8441
timestamp 1386234792
transform 1 0 25083 0 1 1008
box 0 0 96 799
use nand2 stateSub_reg_91_1_93_
timestamp 1386234792
transform 1 0 25179 0 1 1008
box 0 0 96 799
use scandtype g8316
timestamp 1386241841
transform 1 0 25275 0 1 1008
box 0 0 624 799
use inv g8364
timestamp 1386238110
transform 1 0 25899 0 1 1008
box 0 0 120 799
use inv g8378
timestamp 1386238110
transform 1 0 26019 0 1 1008
box 0 0 120 799
use nand2 g8291
timestamp 1386234792
transform 1 0 26139 0 1 1008
box 0 0 96 799
use nand2 g8112
timestamp 1386234792
transform 1 0 26235 0 1 1008
box 0 0 96 799
use nand2 g8448
timestamp 1386234792
transform 1 0 26331 0 1 1008
box 0 0 96 799
use inv Flags_91_0_93_
timestamp 1386238110
transform 1 0 26427 0 1 1008
box 0 0 120 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27123 0 1 1008
box 0 0 320 799
<< labels >>
rlabel m2contact 26409 127 26409 127 8 OpcodeCondIn[4]
rlabel m2contact 26409 31 26409 31 8 OpcodeCondIn[4]
rlabel m2contact 26385 151 26385 151 8 OpcodeCondIn[0]
rlabel m2contact 26385 31 26385 31 8 OpcodeCondIn[0]
rlabel m2contact 26361 247 26361 247 8 OpcodeCondIn[2]
rlabel m2contact 26361 103 26361 103 8 OpcodeCondIn[2]
rlabel m2contact 26337 751 26337 751 8 OpcodeCondIn[7]
rlabel m2contact 26337 79 26337 79 8 OpcodeCondIn[7]
rlabel m2contact 26313 391 26313 391 8 OpcodeCondIn[6]
rlabel m2contact 26313 55 26313 55 8 OpcodeCondIn[6]
rlabel m2contact 26313 559 26313 559 8 n_126
rlabel m2contact 26217 343 26217 343 8 n_56
rlabel m2contact 26049 511 26049 511 8 n_108
rlabel m2contact 25377 895 25377 895 6 n_313
rlabel m2contact 25257 439 25257 439 8 n_52
rlabel m2contact 25233 127 25233 127 8 OpcodeCondIn[4]
rlabel m2contact 25137 775 25137 775 8 n_309
rlabel m2contact 25113 103 25113 103 8 n_306
rlabel m2contact 25041 583 25041 583 8 n_97
rlabel m2contact 24057 199 24057 199 8 n_118
rlabel m2contact 24009 319 24009 319 8 n_155
rlabel m2contact 23961 943 23961 943 6 n_119
rlabel m2contact 23769 535 23769 535 8 n_60
rlabel m2contact 23721 871 23721 871 6 n_58
rlabel m2contact 23649 103 23649 103 8 n_306
rlabel m2contact 23361 751 23361 751 8 OpcodeCondIn[7]
rlabel m2contact 23289 391 23289 391 8 OpcodeCondIn[6]
rlabel m2contact 23217 415 23217 415 8 n_233
rlabel m2contact 23193 55 23193 55 8 n_50
rlabel m2contact 23121 607 23121 607 8 n_216
rlabel m2contact 23025 799 23025 799 6 n_255
rlabel m2contact 22977 607 22977 607 8 n_216
rlabel m2contact 22929 847 22929 847 6 n_279
rlabel m2contact 22809 391 22809 391 8 OpcodeCondIn[6]
rlabel m2contact 22545 463 22545 463 8 n_117
rlabel m2contact 22497 535 22497 535 8 n_60
rlabel m2contact 22329 535 22329 535 8 n_66
rlabel m2contact 22305 391 22305 391 8 OpcodeCondIn[6]
rlabel m2contact 22209 271 22209 271 8 n_31
rlabel m2contact 22185 823 22185 823 6 n_252
rlabel m2contact 22161 607 22161 607 8 n_254
rlabel m2contact 22089 991 22089 991 6 n_289
rlabel m2contact 22041 655 22041 655 8 n_253
rlabel m2contact 21705 703 21705 703 8 n_295
rlabel m2contact 20865 631 20865 631 8 n_111
rlabel m2contact 20841 727 20841 727 8 n_476
rlabel m2contact 20817 679 20817 679 8 IRQ1
rlabel m2contact 20769 703 20769 703 8 n_295
rlabel m2contact 20553 919 20553 919 6 n_173
rlabel m2contact 20457 703 20457 703 8 n_197
rlabel m2contact 20265 247 20265 247 8 OpcodeCondIn[2]
rlabel m2contact 20121 823 20121 823 6 n_252
rlabel m2contact 19857 583 19857 583 8 n_97
rlabel m2contact 19713 679 19713 679 8 IRQ1
rlabel m2contact 19185 823 19185 823 6 n_48
rlabel m2contact 19089 943 19089 943 6 n_119
rlabel m2contact 19041 199 19041 199 8 n_118
rlabel m2contact 18273 799 18273 799 6 n_255
rlabel m2contact 18081 799 18081 799 6 n_9
rlabel m2contact 17865 487 17865 487 8 n_180
rlabel m2contact 17721 295 17721 295 8 n_293
rlabel m2contact 17577 223 17577 223 8 IRQ2
rlabel m2contact 17529 727 17529 727 8 n_476
rlabel m2contact 17169 679 17169 679 8 IRQ1
rlabel m2contact 17001 967 17001 967 6 n_146
rlabel m2contact 16809 535 16809 535 8 n_66
rlabel m2contact 16737 751 16737 751 8 OpcodeCondIn[7]
rlabel m2contact 16713 679 16713 679 8 n_4
rlabel m2contact 16473 727 16473 727 8 n_110
rlabel m2contact 16377 367 16377 367 8 n_315
rlabel m2contact 16257 943 16257 943 6 n_17
rlabel m2contact 16137 751 16137 751 8 OpcodeCondIn[7]
rlabel m2contact 16089 535 16089 535 8 n_20
rlabel m2contact 15993 271 15993 271 8 n_31
rlabel m2contact 15897 607 15897 607 8 n_254
rlabel m2contact 15849 655 15849 655 8 n_253
rlabel m2contact 15609 799 15609 799 6 n_9
rlabel m2contact 15417 271 15417 271 8 n_478
rlabel m2contact 14529 607 14529 607 8 n_100
rlabel m2contact 14505 223 14505 223 8 IRQ2
rlabel m2contact 14481 271 14481 271 8 n_478
rlabel m2contact 14361 391 14361 391 8 OpcodeCondIn[6]
rlabel m2contact 14217 775 14217 775 8 n_309
rlabel m2contact 14121 151 14121 151 8 n_30
rlabel m2contact 14097 751 14097 751 8 OpcodeCondIn[7]
rlabel m2contact 14025 223 14025 223 2 n_39
rlabel m2contact 13809 79 13809 79 2 n_163
rlabel m2contact 13785 175 13785 175 2 n_127
rlabel m2contact 13761 775 13761 775 2 n_143
rlabel m2contact 13713 271 13713 271 2 n_218
rlabel m2contact 13689 223 13689 223 2 n_39
rlabel m2contact 13665 319 13665 319 2 n_155
rlabel m2contact 13617 319 13617 319 2 n_46
rlabel m2contact 13473 223 13473 223 2 n_116
rlabel m2contact 13449 343 13449 343 2 n_56
rlabel m2contact 12945 175 12945 175 2 n_127
rlabel m2contact 12921 343 12921 343 2 n_5
rlabel m2contact 12849 439 12849 439 2 n_52
rlabel m2contact 12585 991 12585 991 4 n_289
rlabel m2contact 12393 967 12393 967 4 n_146
rlabel m2contact 12249 943 12249 943 4 n_17
rlabel m2contact 12105 703 12105 703 2 n_197
rlabel m2contact 11913 751 11913 751 2 OpcodeCondIn[7]
rlabel m2contact 11817 919 11817 919 4 n_173
rlabel m2contact 11793 703 11793 703 2 n_160
rlabel m2contact 11697 895 11697 895 4 n_313
rlabel m2contact 11289 127 11289 127 2 OpcodeCondIn[4]
rlabel m2contact 11097 703 11097 703 2 n_160
rlabel m2contact 10929 511 10929 511 2 n_108
rlabel m2contact 10857 871 10857 871 4 n_58
rlabel m2contact 10761 703 10761 703 2 n_241
rlabel m2contact 10473 751 10473 751 2 OpcodeCondIn[7]
rlabel m2contact 10041 871 10041 871 4 n_58
rlabel m2contact 9969 7 9969 7 2 OpcodeCondIn[5]
rlabel m2contact 9801 655 9801 655 2 n_253
rlabel m2contact 9705 511 9705 511 2 n_108
rlabel m2contact 9105 655 9105 655 2 n_234
rlabel m2contact 8985 511 8985 511 2 n_207
rlabel m2contact 8937 79 8937 79 2 n_163
rlabel m2contact 8889 79 8889 79 2 n_18
rlabel m2contact 8865 127 8865 127 2 OpcodeCondIn[4]
rlabel m2contact 8817 751 8817 751 2 OpcodeCondIn[7]
rlabel m2contact 8649 127 8649 127 2 OpcodeCondIn[4]
rlabel m2contact 8505 847 8505 847 4 n_279
rlabel m2contact 8385 823 8385 823 4 n_48
rlabel m2contact 8217 799 8217 799 4 n_9
rlabel m2contact 8193 247 8193 247 2 OpcodeCondIn[2]
rlabel m2contact 8001 775 8001 775 2 n_143
rlabel m2contact 7977 751 7977 751 2 OpcodeCondIn[7]
rlabel m2contact 7833 391 7833 391 2 OpcodeCondIn[6]
rlabel m2contact 7545 727 7545 727 2 n_110
rlabel m2contact 7305 703 7305 703 2 n_241
rlabel m2contact 7041 679 7041 679 2 n_4
rlabel m2contact 7017 391 7017 391 2 OpcodeCondIn[6]
rlabel m2contact 6825 655 6825 655 2 n_234
rlabel m2contact 6801 631 6801 631 2 n_111
rlabel m2contact 6777 607 6777 607 2 n_100
rlabel m2contact 6705 583 6705 583 2 n_97
rlabel m2contact 6681 439 6681 439 2 n_52
rlabel m2contact 6609 439 6609 439 2 n_157
rlabel m2contact 6561 559 6561 559 2 n_126
rlabel m2contact 6489 535 6489 535 2 n_20
rlabel m2contact 6465 511 6465 511 2 n_207
rlabel m2contact 6273 79 6273 79 2 n_18
rlabel m2contact 5601 79 5601 79 2 Flags[2]
rlabel m2contact 5553 487 5553 487 2 n_180
rlabel m2contact 5505 463 5505 463 2 n_117
rlabel m2contact 5481 439 5481 439 2 n_157
rlabel m2contact 5361 31 5361 31 2 OpcodeCondIn[0]
rlabel m2contact 5241 415 5241 415 2 n_233
rlabel m2contact 5025 391 5025 391 2 OpcodeCondIn[6]
rlabel m2contact 4737 199 4737 199 2 n_118
rlabel m2contact 4689 247 4689 247 2 OpcodeCondIn[2]
rlabel m2contact 4593 367 4593 367 2 n_315
rlabel m2contact 4569 199 4569 199 2 n_331
rlabel m2contact 4497 343 4497 343 2 n_5
rlabel m2contact 4305 319 4305 319 2 n_46
rlabel m2contact 4209 295 4209 295 2 n_293
rlabel m2contact 4161 271 4161 271 2 n_218
rlabel m2contact 3873 247 3873 247 2 OpcodeCondIn[2]
rlabel m2contact 3705 127 3705 127 2 OpcodeCondIn[4]
rlabel m2contact 3609 127 3609 127 2 Flags[1]
rlabel m2contact 3489 223 3489 223 2 n_116
rlabel m2contact 2721 103 2721 103 2 n_306
rlabel m2contact 2673 199 2673 199 2 n_331
rlabel m2contact 2649 103 2649 103 2 Flags[3]
rlabel m2contact 2457 175 2457 175 2 n_127
rlabel m2contact 2385 151 2385 151 2 n_30
rlabel m2contact 2337 55 2337 55 2 n_50
rlabel m2contact 2241 55 2241 55 2 Flags[0]
rlabel m2contact 26097 8081 26097 8081 6 Op1Sel
rlabel m2contact 25701 8129 25701 8129 6 MemEn
rlabel m2contact 24201 8033 24201 8033 6 IrWe
rlabel m2contact 24105 8033 24105 8033 6 IrWe
rlabel m2contact 23985 7961 23985 7961 6 AluEn
rlabel m2contact 23745 8033 23745 8033 6 ImmSel
rlabel m2contact 22701 8057 22701 8057 6 LrSel
rlabel metal2 22227 8153 22227 8153 6 LrWe
rlabel m2contact 22209 8153 22209 8153 6 LrWe
rlabel metal2 20571 8153 20571 8153 6 WdSel
rlabel m2contact 20553 8153 20553 8153 6 WdSel
rlabel m2contact 19953 8081 19953 8081 6 Op1Sel
rlabel m2contact 19713 8105 19713 8105 6 RwSel[1]
rlabel m2contact 18369 7889 18369 7889 6 RwSel[0]
rlabel m2contact 18321 8153 18321 8153 6 PcSel[0]
rlabel m2contact 18201 8105 18201 8105 6 LrEn
rlabel m2contact 18177 7985 18177 7985 6 CFlag
rlabel m2contact 18177 8153 18177 8153 6 PcSel[0]
rlabel m2contact 16665 7889 16665 7889 6 PcWe
rlabel m2contact 15201 7985 15201 7985 6 PcSel[1]
rlabel metal2 14475 8153 14475 8153 6 PcSel[2]
rlabel m2contact 14457 8153 14457 8153 6 PcSel[2]
rlabel m2contact 12873 8129 12873 8129 4 MemEn
rlabel m2contact 12369 7913 12369 7913 4 Rs1Sel[0]
rlabel m2contact 12189 7913 12189 7913 4 PcEn
rlabel m2contact 12153 7889 12153 7889 4 PcWe
rlabel m2contact 10713 7985 10713 7985 4 PcSel[1]
rlabel m2contact 10641 8081 10641 8081 4 Op1Sel
rlabel m2contact 10137 7985 10137 7985 4 nWait
rlabel m2contact 9129 8033 9129 8033 4 ImmSel
rlabel m2contact 8889 7913 8889 7913 4 PcEn
rlabel m2contact 8769 8033 8769 8033 4 ALE
rlabel m2contact 7833 7913 7833 7913 4 AluWe
rlabel metal2 6915 8081 6915 8081 4 Op2Sel[0]
rlabel m2contact 6897 8081 6897 8081 4 Op2Sel[0]
rlabel m2contact 4629 8081 4629 8081 4 Op2Sel[1]
rlabel m2contact 4593 7913 4593 7913 4 AluWe
rlabel m2contact 4113 8105 4113 8105 4 LrEn
rlabel m2contact 3705 7937 3705 7937 4 AluOR[0]
rlabel m2contact 3273 8081 3273 8081 4 Op2Sel[1]
rlabel m2contact 3081 7961 3081 7961 4 AluEn
rlabel m2contact 2889 8057 2889 8057 4 LrSel
rlabel m2contact 2313 8009 2313 8009 4 Rs1Sel[1]
rlabel m2contact 1737 8009 1737 8009 4 nME
rlabel m2contact 27225 6792 27225 6792 6 SysBus[1]
rlabel m2contact 27225 1944 27225 1944 6 SysBus[1]
rlabel m2contact 27201 2136 27201 2136 6 SysBus[0]
rlabel m2contact 27201 1920 27201 1920 6 SysBus[0]
rlabel m2contact 27177 6408 27177 6408 6 SysBus[2]
rlabel m2contact 27177 1872 27177 1872 6 SysBus[2]
rlabel m2contact 27153 5088 27153 5088 6 OpcodeCondIn[3]
rlabel m2contact 27153 1848 27153 1848 6 OpcodeCondIn[3]
rlabel m2contact 27129 5544 27129 5544 6 OpcodeCondIn[1]
rlabel m2contact 27129 1824 27129 1824 6 OpcodeCondIn[1]
rlabel m2contact 27105 4080 27105 4080 6 SysBus[3]
rlabel m2contact 27105 1896 27105 1896 6 SysBus[3]
rlabel m2contact 27105 4344 27105 4344 6 RegWe
rlabel m2contact 27057 6552 27057 6552 6 n_21
rlabel m2contact 27009 3960 27009 3960 6 state[0]
rlabel m2contact 26985 3984 26985 3984 6 stateSub[2]
rlabel m2contact 26937 2352 26937 2352 6 n_303
rlabel m2contact 26889 4104 26889 4104 6 stateSub[0]
rlabel m2contact 26865 3744 26865 3744 6 n_258
rlabel m2contact 26817 3360 26817 3360 6 n_314
rlabel m2contact 26793 4320 26793 4320 6 n_186
rlabel m2contact 26769 4992 26769 4992 6 n_249
rlabel m2contact 26745 5928 26745 5928 6 n_265
rlabel m2contact 26697 5736 26697 5736 6 n_115
rlabel m2contact 26673 5496 26673 5496 6 n_166
rlabel m2contact 26673 2112 26673 2112 6 n_166
rlabel m2contact 26649 4008 26649 4008 6 n_202
rlabel m2contact 26625 3312 26625 3312 6 n_172
rlabel m2contact 26601 6432 26601 6432 6 n_151
rlabel m2contact 26601 4440 26601 4440 6 n_151
rlabel m2contact 26577 4608 26577 4608 6 n_194
rlabel m2contact 26553 5112 26553 5112 6 n_134
rlabel m2contact 26529 2952 26529 2952 6 n_125
rlabel m2contact 26505 2400 26505 2400 6 n_145
rlabel m2contact 26505 3984 26505 3984 6 stateSub[2]
rlabel m2contact 26481 5880 26481 5880 6 n_74
rlabel m2contact 26481 3624 26481 3624 6 n_74
rlabel m2contact 26457 5496 26457 5496 6 n_166
rlabel m2contact 26457 5472 26457 5472 6 n_40
rlabel m2contact 26433 3384 26433 3384 6 n_130
rlabel m2contact 26409 4632 26409 4632 6 n_316
rlabel m2contact 26409 5016 26409 5016 6 n_152
rlabel m2contact 26385 3480 26385 3480 6 n_317
rlabel m2contact 26361 6432 26361 6432 6 n_151
rlabel m2contact 26361 6408 26361 6408 6 SysBus[2]
rlabel m2contact 26337 5688 26337 5688 6 n_296
rlabel m2contact 26337 2688 26337 2688 6 n_296
rlabel m2contact 26313 4008 26313 4008 6 n_202
rlabel m2contact 26289 3624 26289 3624 6 n_74
rlabel m2contact 26289 3648 26289 3648 6 n_259
rlabel m2contact 26265 2952 26265 2952 6 n_125
rlabel m2contact 26241 6840 26241 6840 6 n_327
rlabel m2contact 26217 3624 26217 3624 6 stateSub[1]
rlabel m2contact 26193 5688 26193 5688 6 n_296
rlabel m2contact 26193 5664 26193 5664 6 n_243
rlabel m2contact 26169 4128 26169 4128 6 n_59
rlabel m2contact 26145 7056 26145 7056 6 n_358
rlabel m2contact 26097 4464 26097 4464 6 n_109
rlabel m2contact 26073 6720 26073 6720 6 n_349
rlabel m2contact 26025 5448 26025 5448 6 n_11
rlabel m2contact 25977 4968 25977 4968 6 n_185
rlabel m2contact 25977 5280 25977 5280 6 n_280
rlabel m2contact 25953 3960 25953 3960 6 state[0]
rlabel m2contact 25929 4176 25929 4176 6 n_147
rlabel m2contact 25881 4392 25881 4392 6 n_247
rlabel m2contact 25833 5952 25833 5952 6 n_214
rlabel m2contact 25785 5784 25785 5784 6 n_82
rlabel m2contact 25785 3624 25785 3624 6 stateSub[1]
rlabel m2contact 25761 3768 25761 3768 6 state[1]
rlabel m2contact 25737 5496 25737 5496 6 n_79
rlabel m2contact 25737 5280 25737 5280 6 n_280
rlabel m2contact 25689 4752 25689 4752 6 n_200
rlabel m2contact 25665 3816 25665 3816 6 n_96
rlabel m2contact 25641 6336 25641 6336 6 n_198
rlabel m2contact 25617 3648 25617 3648 6 n_259
rlabel m2contact 25545 4080 25545 4080 6 SysBus[3]
rlabel m2contact 25473 5616 25473 5616 6 n_235
rlabel m2contact 25401 6696 25401 6696 6 StatusReg[3]
rlabel m2contact 25353 6360 25353 6360 6 n_335
rlabel m2contact 25329 4560 25329 4560 6 Flags[0]
rlabel m2contact 25305 3912 25305 3912 6 n_333
rlabel m2contact 25257 4920 25257 4920 6 n_346
rlabel m2contact 25233 4368 25233 4368 6 n_246
rlabel m2contact 25209 5832 25209 5832 6 n_93
rlabel m2contact 25209 3216 25209 3216 6 n_237
rlabel m2contact 25161 5904 25161 5904 6 n_206
rlabel m2contact 25161 4944 25161 4944 6 LrWe
rlabel m2contact 25137 4680 25137 4680 6 n_106
rlabel m2contact 25113 5856 25113 5856 6 n_215
rlabel m2contact 25065 6240 25065 6240 6 n_170
rlabel m2contact 25065 2376 25065 2376 6 n_150
rlabel m2contact 25017 6744 25017 6744 6 OpcodeCondIn[6]
rlabel m2contact 25017 5376 25017 5376 6 n_187
rlabel m2contact 24993 6864 24993 6864 6 OpcodeCondIn[7]
rlabel m2contact 24921 3816 24921 3816 6 n_96
rlabel m2contact 24897 4488 24897 4488 6 OpcodeCondIn[5]
rlabel m2contact 24897 3168 24897 3168 6 OpcodeCondIn[5]
rlabel m2contact 24873 4488 24873 4488 6 OpcodeCondIn[5]
rlabel m2contact 24873 3960 24873 3960 6 state[0]
rlabel m2contact 24825 2664 24825 2664 6 n_184
rlabel m2contact 24801 2064 24801 2064 6 n_339
rlabel m2contact 24777 2544 24777 2544 6 IntReq
rlabel m2contact 24705 2616 24705 2616 6 n_33
rlabel m2contact 24657 3288 24657 3288 6 n_32
rlabel m2contact 24609 5712 24609 5712 6 n_204
rlabel m2contact 24585 5568 24585 5568 6 n_53
rlabel m2contact 24561 2400 24561 2400 6 n_145
rlabel m2contact 24537 6384 24537 6384 6 n_171
rlabel m2contact 24489 4488 24489 4488 6 n_242
rlabel m2contact 24465 5904 24465 5904 6 n_206
rlabel m2contact 24465 5808 24465 5808 6 n_338
rlabel m2contact 24441 6984 24441 6984 6 n_179
rlabel m2contact 24393 4416 24393 4416 6 n_43
rlabel m2contact 24369 5544 24369 5544 6 OpcodeCondIn[1]
rlabel m2contact 24345 5520 24345 5520 6 n_282
rlabel m2contact 24321 6792 24321 6792 6 SysBus[1]
rlabel m2contact 24297 7032 24297 7032 6 n_275
rlabel m2contact 24273 2712 24273 2712 6 StatusReg[2]
rlabel m2contact 24249 6672 24249 6672 6 n_277
rlabel m2contact 24249 5616 24249 5616 6 n_235
rlabel m2contact 24201 3840 24201 3840 6 n_312
rlabel m2contact 24177 2016 24177 2016 6 CFlag
rlabel m2contact 24177 3216 24177 3216 6 n_237
rlabel m2contact 24153 6648 24153 6648 6 n_308
rlabel m2contact 24129 7008 24129 7008 6 n_203
rlabel m2contact 24105 4008 24105 4008 6 n_202
rlabel m2contact 24081 5424 24081 5424 6 n_201
rlabel m2contact 24057 4680 24057 4680 6 n_106
rlabel m2contact 24033 4800 24033 4800 6 n_91
rlabel m2contact 23961 4536 23961 4536 6 n_365
rlabel m2contact 23937 7056 23937 7056 6 n_358
rlabel m2contact 23937 6960 23937 6960 6 n_70
rlabel m2contact 23913 4848 23913 4848 6 n_364
rlabel m2contact 23865 6480 23865 6480 6 n_321
rlabel m2contact 23841 5136 23841 5136 6 n_76
rlabel m2contact 23817 3912 23817 3912 6 n_333
rlabel m2contact 23793 6120 23793 6120 6 n_75
rlabel m2contact 23721 4848 23721 4848 6 n_364
rlabel m2contact 23697 5352 23697 5352 6 n_273
rlabel m2contact 23697 4128 23697 4128 6 n_59
rlabel m2contact 23673 4200 23673 4200 6 n_231
rlabel m2contact 23649 3504 23649 3504 6 n_230
rlabel m2contact 23625 3024 23625 3024 6 n_220
rlabel m2contact 23601 6168 23601 6168 6 n_212
rlabel m2contact 23601 3600 23601 3600 6 n_292
rlabel m2contact 23577 6624 23577 6624 6 n_1
rlabel m2contact 23577 4296 23577 4296 6 n_1
rlabel m2contact 23553 4512 23553 4512 6 n_288
rlabel m2contact 23529 4296 23529 4296 6 n_1
rlabel m2contact 23529 5304 23529 5304 6 n_178
rlabel m2contact 23493 5160 23493 5160 6 n_51
rlabel m2contact 23493 2928 23493 2928 6 n_51
rlabel m2contact 23481 2088 23481 2088 6 nWait
rlabel m2contact 23457 5832 23457 5832 6 n_93
rlabel m2contact 23433 2760 23433 2760 6 n_250
rlabel m2contact 23409 5160 23409 5160 6 n_51
rlabel m2contact 23409 5088 23409 5088 6 OpcodeCondIn[3]
rlabel m2contact 23385 4656 23385 4656 6 n_223
rlabel m2contact 23361 1896 23361 1896 6 n_90
rlabel m2contact 23337 6504 23337 6504 6 n_148
rlabel m2contact 23313 5160 23313 5160 6 n_222
rlabel m2contact 23313 6528 23313 6528 6 n_89
rlabel m2contact 23265 6720 23265 6720 6 n_349
rlabel m2contact 23265 6600 23265 6600 6 n_227
rlabel m2contact 23241 5040 23241 5040 6 n_348
rlabel m2contact 23217 6000 23217 6000 6 n_228
rlabel m2contact 23193 4872 23193 4872 6 n_297
rlabel m2contact 23169 4728 23169 4728 6 n_251
rlabel m2contact 23169 3552 23169 3552 6 n_232
rlabel m2contact 23145 5856 23145 5856 6 n_215
rlabel m2contact 23145 4056 23145 4056 6 n_215
rlabel m2contact 23145 3792 23145 3792 6 StatusReg[0]
rlabel m2contact 23145 2328 23145 2328 6 StatusReg[0]
rlabel m2contact 23121 1992 23121 1992 6 n_25
rlabel m2contact 23097 4512 23097 4512 6 n_288
rlabel m2contact 23097 4128 23097 4128 6 n_59
rlabel m2contact 23073 4056 23073 4056 6 n_215
rlabel m2contact 23073 4104 23073 4104 6 stateSub[0]
rlabel m2contact 23049 3312 23049 3312 6 n_172
rlabel m2contact 23025 3528 23025 3528 6 n_102
rlabel m2contact 23025 2784 23025 2784 6 n_102
rlabel m2contact 23013 5208 23013 5208 6 n_272
rlabel m2contact 23013 4296 23013 4296 6 n_272
rlabel m2contact 23001 5256 23001 5256 6 n_139
rlabel m2contact 23001 3576 23001 3576 6 n_153
rlabel m2contact 22977 3960 22977 3960 6 state[0]
rlabel m2contact 22953 2544 22953 2544 6 IntReq
rlabel m2contact 22929 2472 22929 2472 6 n_72
rlabel m2contact 22905 2328 22905 2328 6 StatusReg[0]
rlabel m2contact 22905 2400 22905 2400 6 n_145
rlabel m2contact 22881 6672 22881 6672 6 n_277
rlabel m2contact 22857 5184 22857 5184 6 n_248
rlabel m2contact 22833 4296 22833 4296 6 n_272
rlabel m2contact 22833 4368 22833 4368 6 n_246
rlabel m2contact 22809 4392 22809 4392 6 n_247
rlabel m2contact 22785 3744 22785 3744 6 n_258
rlabel m2contact 22761 6720 22761 6720 6 n_29
rlabel m2contact 22737 5592 22737 5592 6 n_64
rlabel m2contact 22713 5544 22713 5544 6 OpcodeCondIn[1]
rlabel m2contact 22713 4008 22713 4008 6 n_202
rlabel m2contact 22689 2784 22689 2784 6 n_102
rlabel m2contact 22689 2808 22689 2808 6 n_8
rlabel m2contact 22653 6072 22653 6072 6 n_225
rlabel m2contact 22653 4296 22653 4296 6 n_225
rlabel m2contact 22641 4152 22641 4152 6 n_226
rlabel m2contact 22617 4296 22617 4296 6 n_225
rlabel m2contact 22617 4368 22617 4368 6 n_246
rlabel m2contact 22593 5952 22593 5952 6 n_214
rlabel m2contact 22569 4824 22569 4824 6 n_85
rlabel m2contact 22545 4776 22545 4776 6 n_36
rlabel m2contact 22545 2328 22545 2328 6 n_36
rlabel m2contact 22521 4704 22521 4704 6 n_28
rlabel m2contact 22497 5520 22497 5520 6 n_282
rlabel m2contact 22473 4896 22473 4896 6 n_57
rlabel m2contact 22473 5328 22473 5328 6 n_236
rlabel m2contact 22437 4584 22437 4584 6 n_15
rlabel m2contact 22437 3936 22437 3936 6 n_15
rlabel m2contact 22425 5064 22425 5064 6 n_304
rlabel m2contact 22425 3240 22425 3240 6 n_37
rlabel m2contact 22401 3936 22401 3936 6 n_15
rlabel m2contact 22401 4032 22401 4032 6 n_49
rlabel m2contact 22377 2328 22377 2328 6 n_36
rlabel m2contact 22377 2352 22377 2352 6 n_303
rlabel m2contact 22353 5280 22353 5280 6 n_280
rlabel m2contact 22329 5976 22329 5976 6 n_65
rlabel m2contact 22329 4296 22329 4296 6 n_65
rlabel m2contact 22305 4032 22305 4032 6 n_49
rlabel m2contact 22281 4296 22281 4296 6 n_65
rlabel m2contact 22281 5088 22281 5088 6 OpcodeCondIn[3]
rlabel m2contact 22257 5328 22257 5328 6 n_236
rlabel m2contact 22233 4248 22233 4248 6 nWE
rlabel m2contact 22209 4944 22209 4944 6 LrWe
rlabel m2contact 22161 4896 22161 4896 6 n_57
rlabel m2contact 22137 6072 22137 6072 6 n_225
rlabel m2contact 22113 3960 22113 3960 6 state[0]
rlabel m2contact 22089 4368 22089 4368 6 n_246
rlabel m2contact 22065 4512 22065 4512 6 n_288
rlabel m2contact 22041 4944 22041 4944 6 n_191
rlabel m2contact 22017 4440 22017 4440 6 n_151
rlabel m2contact 22017 3624 22017 3624 6 stateSub[1]
rlabel m2contact 21993 6336 21993 6336 6 n_198
rlabel m2contact 21969 5040 21969 5040 6 n_348
rlabel m2contact 21945 5472 21945 5472 6 n_40
rlabel m2contact 21921 5832 21921 5832 6 n_93
rlabel m2contact 21885 6192 21885 6192 6 StatusReg[0]
rlabel m2contact 21885 3792 21885 3792 6 StatusReg[0]
rlabel m2contact 21873 2568 21873 2568 6 n_209
rlabel m2contact 21849 6192 21849 6192 6 StatusReg[0]
rlabel m2contact 21849 6144 21849 6144 6 n_310
rlabel m2contact 21825 5304 21825 5304 6 n_178
rlabel m2contact 21801 4056 21801 4056 6 n_477
rlabel m2contact 21777 4272 21777 4272 6 nOE
rlabel m2contact 21753 2184 21753 2184 6 n_350
rlabel m2contact 21729 3696 21729 3696 6 n_299
rlabel m2contact 21705 6264 21705 6264 6 n_368
rlabel m2contact 21705 2208 21705 2208 6 n_368
rlabel m2contact 21681 5400 21681 5400 6 n_221
rlabel m2contact 21657 6144 21657 6144 6 n_310
rlabel m2contact 21657 4296 21657 4296 6 n_310
rlabel m2contact 21633 4320 21633 4320 6 n_186
rlabel m2contact 21609 4368 21609 4368 6 n_246
rlabel m2contact 21585 4968 21585 4968 6 n_185
rlabel m2contact 21561 6336 21561 6336 6 n_198
rlabel m2contact 21561 4320 21561 4320 6 n_198
rlabel m2contact 21537 6456 21537 6456 6 n_122
rlabel m2contact 21513 4104 21513 4104 6 stateSub[0]
rlabel m2contact 21489 2904 21489 2904 6 n_95
rlabel m2contact 21465 5424 21465 5424 6 n_201
rlabel m2contact 21465 1848 21465 1848 6 n_201
rlabel m2contact 21441 6264 21441 6264 6 n_368
rlabel m2contact 21441 6216 21441 6216 6 n_54
rlabel m2contact 21417 3312 21417 3312 6 n_172
rlabel m2contact 21393 4680 21393 4680 6 n_106
rlabel m2contact 21357 4896 21357 4896 6 n_88
rlabel m2contact 21357 3144 21357 3144 6 n_88
rlabel m2contact 21345 2976 21345 2976 6 n_174
rlabel m2contact 21321 4992 21321 4992 6 n_249
rlabel m2contact 21321 3024 21321 3024 6 n_220
rlabel m2contact 21297 5016 21297 5016 6 n_152
rlabel m2contact 21297 5088 21297 5088 6 OpcodeCondIn[3]
rlabel m2contact 21273 4296 21273 4296 6 n_310
rlabel m2contact 21273 5640 21273 5640 6 n_244
rlabel m2contact 21249 3624 21249 3624 6 stateSub[1]
rlabel m2contact 21225 6192 21225 6192 6 n_305
rlabel m2contact 21201 4320 21201 4320 6 n_198
rlabel m2contact 21201 5520 21201 5520 6 n_282
rlabel m2contact 21177 2352 21177 2352 6 n_303
rlabel m2contact 21153 3192 21153 3192 6 n_114
rlabel m2contact 21153 3648 21153 3648 6 n_259
rlabel m2contact 21129 5376 21129 5376 6 n_187
rlabel m2contact 21105 6312 21105 6312 6 n_22
rlabel m2contact 21081 3144 21081 3144 6 n_88
rlabel m2contact 21081 3192 21081 3192 6 n_114
rlabel m2contact 21057 6552 21057 6552 6 n_21
rlabel m2contact 21057 3672 21057 3672 6 n_87
rlabel m2contact 21033 6504 21033 6504 6 n_148
rlabel m2contact 21009 4992 21009 4992 6 n_183
rlabel m2contact 20985 5232 20985 5232 6 n_266
rlabel m2contact 20961 6048 20961 6048 6 n_80
rlabel m2contact 20961 4008 20961 4008 6 n_202
rlabel m2contact 20937 1848 20937 1848 6 n_201
rlabel m2contact 20937 1872 20937 1872 6 n_189
rlabel m2contact 20913 3024 20913 3024 6 n_220
rlabel m2contact 20889 5400 20889 5400 6 n_221
rlabel m2contact 20865 3024 20865 3024 6 n_220
rlabel m2contact 20841 4968 20841 4968 6 n_185
rlabel m2contact 20817 3624 20817 3624 6 stateSub[1]
rlabel m2contact 20769 4728 20769 4728 6 n_251
rlabel m2contact 20745 5280 20745 5280 6 n_280
rlabel m2contact 20721 5400 20721 5400 6 n_210
rlabel m2contact 20721 2784 20721 2784 6 n_94
rlabel m2contact 20697 6768 20697 6768 6 n_257
rlabel m2contact 20673 6096 20673 6096 6 n_190
rlabel m2contact 20673 4320 20673 4320 6 n_190
rlabel m2contact 20649 4320 20649 4320 6 n_190
rlabel m2contact 20649 5304 20649 5304 6 n_178
rlabel m2contact 20625 3024 20625 3024 6 n_220
rlabel m2contact 20601 1872 20601 1872 6 n_189
rlabel m2contact 20601 5760 20601 5760 6 n_129
rlabel m2contact 20577 5520 20577 5520 6 n_282
rlabel m2contact 20577 3264 20577 3264 6 n_282
rlabel m2contact 20553 3936 20553 3936 6 WdSel
rlabel m2contact 20529 6024 20529 6024 6 n_131
rlabel m2contact 20505 4968 20505 4968 6 n_256
rlabel m2contact 20505 3312 20505 3312 6 n_172
rlabel m2contact 20469 5280 20469 5280 6 n_280
rlabel m2contact 20469 3456 20469 3456 6 n_280
rlabel m2contact 20457 5904 20457 5904 6 n_264
rlabel m2contact 20433 2568 20433 2568 6 n_209
rlabel m2contact 20409 4728 20409 4728 6 n_42
rlabel m2contact 20385 2856 20385 2856 6 n_161
rlabel m2contact 20385 6528 20385 6528 6 n_89
rlabel m2contact 20361 6288 20361 6288 6 n_138
rlabel m2contact 20361 3072 20361 3072 6 n_138
rlabel m2contact 20337 3168 20337 3168 6 OpcodeCondIn[5]
rlabel m2contact 20313 3264 20313 3264 6 n_282
rlabel m2contact 20313 3312 20313 3312 6 n_172
rlabel m2contact 20289 6264 20289 6264 6 n_55
rlabel m2contact 20289 3048 20289 3048 6 n_55
rlabel m2contact 20265 2880 20265 2880 6 n_199
rlabel m2contact 20241 3216 20241 3216 6 n_237
rlabel m2contact 20217 5688 20217 5688 6 n_92
rlabel m2contact 20217 6336 20217 6336 6 n_198
rlabel m2contact 20193 3456 20193 3456 6 n_280
rlabel m2contact 20193 3672 20193 3672 6 n_87
rlabel m2contact 20169 4800 20169 4800 6 n_91
rlabel m2contact 20145 6384 20145 6384 6 n_171
rlabel m2contact 20121 6240 20121 6240 6 n_170
rlabel m2contact 20097 6288 20097 6288 6 n_138
rlabel m2contact 20097 5280 20097 5280 6 n_280
rlabel m2contact 20073 4392 20073 4392 6 n_247
rlabel m2contact 20049 5880 20049 5880 6 n_74
rlabel m2contact 20025 6864 20025 6864 6 OpcodeCondIn[7]
rlabel m2contact 20001 6264 20001 6264 6 n_55
rlabel m2contact 20001 4008 20001 4008 6 n_202
rlabel m2contact 19977 5880 19977 5880 6 n_98
rlabel m2contact 19977 3720 19977 3720 6 n_98
rlabel m2contact 19953 4776 19953 4776 6 n_36
rlabel m2contact 19929 6264 19929 6264 6 n_292
rlabel m2contact 19929 3600 19929 3600 6 n_292
rlabel m2contact 19905 3720 19905 3720 6 n_98
rlabel m2contact 19905 3864 19905 3864 6 n_113
rlabel m2contact 19881 6264 19881 6264 6 n_292
rlabel m2contact 19881 3816 19881 3816 6 n_96
rlabel m2contact 19833 6288 19833 6288 6 n_336
rlabel m2contact 19785 6192 19785 6192 6 n_305
rlabel m2contact 19761 5064 19761 5064 6 n_304
rlabel m2contact 19689 5064 19689 5064 6 n_300
rlabel m2contact 19665 4944 19665 4944 6 n_191
rlabel m2contact 19641 6096 19641 6096 6 n_190
rlabel m2contact 19617 4944 19617 4944 6 n_301
rlabel m2contact 19569 5808 19569 5808 6 n_338
rlabel m2contact 19545 3336 19545 3336 6 n_23
rlabel m2contact 19521 4320 19521 4320 6 n_177
rlabel m2contact 19497 2448 19497 2448 6 n_276
rlabel m2contact 19473 4392 19473 4392 6 n_83
rlabel m2contact 19425 5568 19425 5568 6 n_53
rlabel m2contact 19401 3168 19401 3168 6 OpcodeCondIn[5]
rlabel m2contact 19377 4296 19377 4296 6 n_71
rlabel m2contact 19329 5568 19329 5568 6 n_328
rlabel m2contact 19305 5520 19305 5520 6 n_282
rlabel m2contact 19305 4224 19305 4224 6 n_3
rlabel m2contact 19281 2304 19281 2304 6 n_270
rlabel m2contact 19233 5400 19233 5400 6 n_210
rlabel m2contact 19209 4176 19209 4176 6 n_147
rlabel m2contact 19185 2568 19185 2568 6 n_209
rlabel m2contact 19161 2328 19161 2328 6 n_47
rlabel m2contact 19137 5352 19137 5352 6 n_273
rlabel m2contact 19137 3672 19137 3672 6 n_87
rlabel m2contact 19089 3720 19089 3720 6 n_239
rlabel m2contact 19065 4992 19065 4992 6 n_183
rlabel m2contact 19041 5400 19041 5400 6 n_217
rlabel m2contact 19041 3456 19041 3456 6 n_217
rlabel m2contact 19017 4056 19017 4056 6 n_477
rlabel m2contact 18993 4872 18993 4872 6 n_297
rlabel m2contact 18969 1872 18969 1872 6 n_189
rlabel m2contact 18945 2688 18945 2688 6 n_296
rlabel m2contact 18921 4440 18921 4440 6 n_151
rlabel m2contact 18897 5424 18897 5424 6 n_201
rlabel m2contact 18897 5376 18897 5376 6 n_187
rlabel m2contact 18873 6816 18873 6816 6 n_339
rlabel m2contact 18873 2064 18873 2064 6 n_339
rlabel m2contact 18849 4344 18849 4344 6 RegWe
rlabel m2contact 18849 6504 18849 6504 6 n_148
rlabel m2contact 18825 5064 18825 5064 6 n_300
rlabel m2contact 18825 5376 18825 5376 6 n_187
rlabel m2contact 18801 2280 18801 2280 6 n_352
rlabel m2contact 18777 4944 18777 4944 6 n_301
rlabel m2contact 18753 3456 18753 3456 6 n_217
rlabel m2contact 18753 3648 18753 3648 6 n_259
rlabel m2contact 18729 6936 18729 6936 6 n_38
rlabel m2contact 18729 4344 18729 4344 6 n_38
rlabel m2contact 18705 2328 18705 2328 6 n_47
rlabel m2contact 18681 3408 18681 3408 6 n_45
rlabel m2contact 18657 4584 18657 4584 6 n_15
rlabel m2contact 18633 5088 18633 5088 6 OpcodeCondIn[3]
rlabel m2contact 18609 3816 18609 3816 6 n_96
rlabel m2contact 18585 2712 18585 2712 6 StatusReg[2]
rlabel m2contact 18561 6816 18561 6816 6 n_339
rlabel m2contact 18561 6696 18561 6696 6 StatusReg[3]
rlabel m2contact 18537 3768 18537 3768 6 state[1]
rlabel m2contact 18513 4464 18513 4464 6 n_109
rlabel m2contact 18513 2160 18513 2160 6 n_224
rlabel m2contact 18489 6504 18489 6504 6 n_148
rlabel m2contact 18465 4872 18465 4872 6 n_101
rlabel m2contact 18465 4656 18465 4656 6 n_223
rlabel m2contact 18441 4512 18441 4512 6 n_288
rlabel m2contact 18417 4344 18417 4344 6 n_38
rlabel m2contact 18417 6096 18417 6096 6 n_44
rlabel m2contact 18393 5544 18393 5544 6 OpcodeCondIn[1]
rlabel m2contact 18369 4056 18369 4056 6 RwSel[0]
rlabel m2contact 18369 2808 18369 2808 6 n_8
rlabel m2contact 18345 4992 18345 4992 6 PcSel[0]
rlabel m2contact 18345 4344 18345 4344 6 PcSel[0]
rlabel m2contact 18321 4992 18321 4992 6 PcSel[0]
rlabel m2contact 18321 4584 18321 4584 6 n_361
rlabel m2contact 18297 6144 18297 6144 6 n_310
rlabel m2contact 18249 4992 18249 4992 6 CFlag
rlabel m2contact 18249 2016 18249 2016 6 CFlag
rlabel m2contact 18225 5352 18225 5352 6 n_324
rlabel m2contact 18201 4464 18201 4464 6 n_99
rlabel m2contact 18177 4992 18177 4992 6 CFlag
rlabel m2contact 18177 3600 18177 3600 6 n_292
rlabel m2contact 18129 3936 18129 3936 6 WdSel
rlabel m2contact 18057 6648 18057 6648 6 n_308
rlabel m2contact 18009 5424 18009 5424 6 n_112
rlabel m2contact 17985 6912 17985 6912 6 n_69
rlabel m2contact 17961 6936 17961 6936 6 n_38
rlabel m2contact 17913 4056 17913 4056 6 RwSel[0]
rlabel m2contact 17889 2520 17889 2520 6 n_268
rlabel m2contact 17841 2736 17841 2736 6 n_104
rlabel m2contact 17817 2592 17817 2592 6 n_156
rlabel m2contact 17769 4344 17769 4344 6 PcSel[0]
rlabel m2contact 17769 4992 17769 4992 6 n_363
rlabel m2contact 17745 2064 17745 2064 6 n_339
rlabel m2contact 17649 6192 17649 6192 6 n_240
rlabel m2contact 17625 5520 17625 5520 6 n_282
rlabel m2contact 17601 5856 17601 5856 6 n_215
rlabel m2contact 17577 3624 17577 3624 6 stateSub[1]
rlabel m2contact 17529 4056 17529 4056 6 n_84
rlabel m2contact 17505 3624 17505 3624 6 stateSub[1]
rlabel m2contact 17481 4800 17481 4800 6 n_91
rlabel m2contact 17433 2184 17433 2184 6 n_350
rlabel m2contact 17385 5784 17385 5784 6 n_82
rlabel m2contact 17361 5688 17361 5688 6 n_92
rlabel m2contact 17289 5400 17289 5400 6 n_217
rlabel m2contact 17241 6600 17241 6600 6 n_227
rlabel m2contact 17193 4344 17193 4344 6 n_144
rlabel m2contact 17169 6816 17169 6816 6 n_27
rlabel m2contact 17145 3888 17145 3888 6 n_68
rlabel m2contact 17121 4872 17121 4872 6 n_101
rlabel m2contact 17097 6072 17097 6072 6 n_225
rlabel m2contact 17097 1824 17097 1824 6 n_225
rlabel m2contact 17073 5400 17073 5400 6 stateSub[1]
rlabel m2contact 17073 3624 17073 3624 6 stateSub[1]
rlabel m2contact 17049 4320 17049 4320 6 n_177
rlabel m2contact 17049 5856 17049 5856 6 n_215
rlabel m2contact 17025 3960 17025 3960 6 state[0]
rlabel m2contact 17001 2112 17001 2112 6 n_166
rlabel m2contact 16977 4872 16977 4872 6 n_196
rlabel m2contact 16977 2496 16977 2496 6 n_196
rlabel m2contact 16953 1824 16953 1824 6 n_225
rlabel m2contact 16953 1848 16953 1848 6 n_263
rlabel m2contact 16929 5400 16929 5400 6 stateSub[1]
rlabel m2contact 16929 4512 16929 4512 6 n_288
rlabel m2contact 16905 4872 16905 4872 6 n_196
rlabel m2contact 16905 3936 16905 3936 6 n_34
rlabel m2contact 16881 5400 16881 5400 6 n_96
rlabel m2contact 16881 3816 16881 3816 6 n_96
rlabel m2contact 16857 4776 16857 4776 6 n_36
rlabel m2contact 16857 2640 16857 2640 6 n_123
rlabel m2contact 16833 5400 16833 5400 6 n_96
rlabel m2contact 16833 5088 16833 5088 6 OpcodeCondIn[3]
rlabel m2contact 16809 5808 16809 5808 6 n_158
rlabel m2contact 16785 6384 16785 6384 6 n_24
rlabel m2contact 16785 4320 16785 4320 6 n_24
rlabel m2contact 16761 4320 16761 4320 6 n_24
rlabel m2contact 16761 4824 16761 4824 6 n_85
rlabel m2contact 16737 4128 16737 4128 6 n_59
rlabel m2contact 16713 5280 16713 5280 6 n_280
rlabel m2contact 16689 6888 16689 6888 6 n_103
rlabel m2contact 16689 2040 16689 2040 6 n_103
rlabel m2contact 16665 6264 16665 6264 6 n_12
rlabel m2contact 16665 3432 16665 3432 6 n_12
rlabel m2contact 16641 2040 16641 2040 6 n_103
rlabel m2contact 16641 2064 16641 2064 6 n_339
rlabel m2contact 16617 4872 16617 4872 6 n_367
rlabel m2contact 16617 4320 16617 4320 6 n_164
rlabel m2contact 16593 3456 16593 3456 6 n_193
rlabel m2contact 16569 3528 16569 3528 6 n_102
rlabel m2contact 16545 6264 16545 6264 6 n_12
rlabel m2contact 16545 5808 16545 5808 6 n_158
rlabel m2contact 16521 5784 16521 5784 6 OpcodeCondIn[4]
rlabel m2contact 16497 3192 16497 3192 6 n_114
rlabel m2contact 16449 5400 16449 5400 6 n_154
rlabel m2contact 16449 3648 16449 3648 6 n_259
rlabel m2contact 16425 6432 16425 6432 6 n_13
rlabel m2contact 16425 5736 16425 5736 6 n_115
rlabel m2contact 16401 5880 16401 5880 6 n_98
rlabel m2contact 16377 5688 16377 5688 6 n_41
rlabel m2contact 16353 3480 16353 3480 6 n_317
rlabel m2contact 16329 4080 16329 4080 6 SysBus[3]
rlabel m2contact 16329 5688 16329 5688 6 n_41
rlabel m2contact 16305 3192 16305 3192 6 n_114
rlabel m2contact 16281 4776 16281 4776 6 n_36
rlabel m2contact 16161 5088 16161 5088 6 OpcodeCondIn[3]
rlabel m2contact 16137 3984 16137 3984 6 stateSub[2]
rlabel m2contact 16089 3312 16089 3312 6 n_172
rlabel m2contact 16065 4128 16065 4128 6 n_59
rlabel m2contact 16041 4512 16041 4512 6 n_288
rlabel m2contact 15969 4104 15969 4104 6 stateSub[0]
rlabel m2contact 15945 3936 15945 3936 6 n_34
rlabel m2contact 15873 4512 15873 4512 6 n_288
rlabel m2contact 15813 6264 15813 6264 6 n_219
rlabel m2contact 15813 4776 15813 4776 6 n_219
rlabel m2contact 15801 4176 15801 4176 6 n_147
rlabel m2contact 15777 3648 15777 3648 6 n_259
rlabel m2contact 15753 5736 15753 5736 6 n_115
rlabel m2contact 15729 6264 15729 6264 6 n_219
rlabel m2contact 15729 6144 15729 6144 6 n_310
rlabel m2contact 15657 4176 15657 4176 6 n_271
rlabel m2contact 15609 6576 15609 6576 6 n_135
rlabel m2contact 15585 5592 15585 5592 6 n_64
rlabel m2contact 15561 4896 15561 4896 6 n_88
rlabel m2contact 15465 3000 15465 3000 6 InISR
rlabel m2contact 15417 6696 15417 6696 6 StatusReg[3]
rlabel m2contact 15057 5592 15057 5592 6 n_347
rlabel m2contact 15009 3144 15009 3144 6 n_356
rlabel m2contact 14961 7056 14961 7056 6 n_63
rlabel m2contact 14961 1920 14961 1920 6 n_63
rlabel m2contact 14937 4200 14937 4200 6 n_231
rlabel m2contact 14913 6240 14913 6240 6 n_170
rlabel m2contact 14889 7056 14889 7056 6 n_63
rlabel m2contact 14889 6600 14889 6600 6 n_227
rlabel m2contact 14865 4008 14865 4008 6 n_202
rlabel m2contact 14841 6384 14841 6384 6 n_24
rlabel m2contact 14841 6264 14841 6264 6 n_319
rlabel m2contact 14817 6144 14817 6144 6 n_310
rlabel m2contact 14793 2424 14793 2424 6 n_294
rlabel m2contact 14793 4896 14793 4896 6 n_162
rlabel m2contact 14769 1944 14769 1944 6 n_132
rlabel m2contact 14745 5256 14745 5256 6 n_139
rlabel m2contact 14745 4200 14745 4200 6 ENB
rlabel m2contact 14721 4056 14721 4056 6 n_84
rlabel m2contact 14697 6384 14697 6384 6 n_320
rlabel m2contact 14697 4080 14697 4080 6 n_311
rlabel m2contact 14673 3480 14673 3480 6 n_317
rlabel m2contact 14649 2136 14649 2136 6 SysBus[0]
rlabel m2contact 14625 4056 14625 4056 6 n_330
rlabel m2contact 14601 5256 14601 5256 6 n_353
rlabel m2contact 14577 3360 14577 3360 6 n_314
rlabel m2contact 14577 5880 14577 5880 6 n_142
rlabel m2contact 14553 6840 14553 6840 6 n_327
rlabel m2contact 14529 5688 14529 5688 6 n_245
rlabel m2contact 14505 7008 14505 7008 6 n_203
rlabel m2contact 14481 6840 14481 6840 6 n_7
rlabel m2contact 14481 2832 14481 2832 6 n_7
rlabel m2contact 14457 2040 14457 2040 6 PcSel[2]
rlabel m2contact 14433 6744 14433 6744 6 OpcodeCondIn[6]
rlabel m2contact 14433 3360 14433 3360 6 OpcodeCondIn[6]
rlabel m2contact 14409 6840 14409 6840 6 n_7
rlabel m2contact 14409 5328 14409 5328 6 n_236
rlabel m2contact 14385 6624 14385 6624 6 n_1
rlabel m2contact 14361 3360 14361 3360 6 OpcodeCondIn[6]
rlabel m2contact 14361 4104 14361 4104 6 stateSub[0]
rlabel m2contact 14337 6840 14337 6840 6 n_175
rlabel m2contact 14337 2232 14337 2232 6 n_175
rlabel m2contact 14313 6120 14313 6120 6 n_75
rlabel m2contact 14313 6624 14313 6624 6 n_211
rlabel m2contact 14289 5088 14289 5088 6 OpcodeCondIn[3]
rlabel m2contact 14265 6840 14265 6840 6 n_175
rlabel m2contact 14265 4296 14265 4296 6 n_71
rlabel m2contact 14241 5376 14241 5376 6 n_187
rlabel m2contact 14217 6648 14217 6648 6 n_308
rlabel m2contact 14217 3360 14217 3360 6 n_308
rlabel m2contact 14193 4176 14193 4176 6 n_271
rlabel m2contact 14169 3360 14169 3360 6 n_308
rlabel m2contact 14169 4800 14169 4800 6 n_91
rlabel m2contact 14145 7008 14145 7008 6 StatusReg[0]
rlabel m2contact 14145 3792 14145 3792 6 StatusReg[0]
rlabel m2contact 14121 6072 14121 6072 6 n_225
rlabel m2contact 14085 5520 14085 5520 6 n_282
rlabel m2contact 14085 3264 14085 3264 6 n_282
rlabel m2contact 14073 6024 14073 6024 6 n_131
rlabel m2contact 14073 2328 14073 2328 6 n_47
rlabel m2contact 14049 3360 14049 3360 6 OpcodeCondIn[2]
rlabel m2contact 14025 4440 14025 4440 4 n_151
rlabel m2contact 14001 3264 14001 3264 4 n_282
rlabel m2contact 14001 3384 14001 3384 4 n_130
rlabel m2contact 13977 6936 13977 6936 4 n_38
rlabel m2contact 13953 3264 13953 3264 4 n_19
rlabel m2contact 13929 5544 13929 5544 4 OpcodeCondIn[1]
rlabel m2contact 13905 7008 13905 7008 4 StatusReg[0]
rlabel m2contact 13905 6912 13905 6912 4 n_69
rlabel m2contact 13881 4440 13881 4440 4 OpcodeCondIn[0]
rlabel m2contact 13857 6720 13857 6720 4 n_29
rlabel m2contact 13833 5880 13833 5880 4 n_142
rlabel m2contact 13809 4008 13809 4008 4 n_202
rlabel m2contact 13785 6072 13785 6072 4 n_208
rlabel m2contact 13761 6840 13761 6840 4 n_26
rlabel m2contact 13737 6504 13737 6504 4 n_148
rlabel m2contact 13713 7008 13713 7008 4 n_102
rlabel m2contact 13713 3528 13713 3528 4 n_102
rlabel m2contact 13689 5064 13689 5064 4 n_300
rlabel m2contact 13665 6072 13665 6072 4 n_208
rlabel m2contact 13641 3264 13641 3264 4 n_19
rlabel m2contact 13641 5856 13641 5856 4 n_215
rlabel m2contact 13617 6024 13617 6024 4 n_78
rlabel m2contact 13617 3120 13617 3120 4 n_78
rlabel m2contact 13593 5880 13593 5880 4 n_359
rlabel m2contact 13569 3864 13569 3864 4 n_113
rlabel m2contact 13569 4632 13569 4632 4 n_316
rlabel m2contact 13545 5424 13545 5424 4 n_112
rlabel m2contact 13545 5856 13545 5856 4 n_332
rlabel m2contact 13521 7032 13521 7032 4 n_275
rlabel m2contact 13521 5520 13521 5520 4 n_282
rlabel m2contact 13497 5616 13497 5616 4 n_235
rlabel m2contact 13497 2256 13497 2256 4 n_235
rlabel m2contact 13473 3600 13473 3600 4 n_292
rlabel m2contact 13449 4632 13449 4632 4 n_45
rlabel m2contact 13449 3408 13449 3408 4 n_45
rlabel m2contact 13425 7008 13425 7008 4 n_102
rlabel m2contact 13425 4824 13425 4824 4 n_85
rlabel m2contact 13401 3552 13401 3552 4 n_232
rlabel m2contact 13377 3864 13377 3864 4 n_14
rlabel m2contact 13353 5280 13353 5280 4 n_280
rlabel m2contact 13329 6024 13329 6024 4 n_78
rlabel m2contact 13329 3312 13329 3312 4 n_172
rlabel m2contact 13293 6024 13293 6024 4 n_128
rlabel m2contact 13293 3264 13293 3264 4 n_128
rlabel m2contact 13281 6936 13281 6936 4 n_38
rlabel m2contact 13257 2136 13257 2136 4 SysBus[0]
rlabel m2contact 13233 3096 13233 3096 4 n_136
rlabel m2contact 13209 4440 13209 4440 4 OpcodeCondIn[0]
rlabel m2contact 13185 2256 13185 2256 4 n_235
rlabel m2contact 13185 4416 13185 4416 4 n_43
rlabel m2contact 13149 6936 13149 6936 4 n_333
rlabel m2contact 13149 3912 13149 3912 4 n_333
rlabel m2contact 13137 6960 13137 6960 4 n_70
rlabel m2contact 13113 3792 13113 3792 4 StatusReg[0]
rlabel m2contact 13089 6912 13089 6912 4 n_69
rlabel m2contact 13065 4632 13065 4632 4 n_45
rlabel m2contact 13065 3792 13065 3792 4 n_281
rlabel m2contact 13041 5280 13041 5280 4 n_280
rlabel m2contact 13017 2352 13017 2352 4 n_303
rlabel m2contact 13017 4632 13017 4632 4 n_159
rlabel m2contact 12993 5808 12993 5808 4 n_158
rlabel m2contact 12969 3264 12969 3264 4 n_128
rlabel m2contact 12969 5376 12969 5376 4 n_187
rlabel m2contact 12945 5520 12945 5520 4 n_282
rlabel m2contact 12921 5424 12921 5424 4 n_112
rlabel m2contact 12897 6912 12897 6912 4 OpcodeCondIn[2]
rlabel m2contact 12897 3360 12897 3360 4 OpcodeCondIn[2]
rlabel m2contact 12873 2472 12873 2472 4 n_72
rlabel m2contact 12873 3264 12873 3264 4 MemEn
rlabel m2contact 12849 6960 12849 6960 4 n_270
rlabel m2contact 12849 2304 12849 2304 4 n_270
rlabel m2contact 12825 6984 12825 6984 4 n_179
rlabel m2contact 12825 6528 12825 6528 4 n_89
rlabel m2contact 12801 3432 12801 3432 4 n_12
rlabel m2contact 12801 5328 12801 5328 4 n_236
rlabel m2contact 12777 5304 12777 5304 4 n_178
rlabel m2contact 12777 4296 12777 4296 4 n_71
rlabel m2contact 12753 3624 12753 3624 4 stateSub[1]
rlabel m2contact 12729 3888 12729 3888 4 n_68
rlabel m2contact 12705 6936 12705 6936 4 n_333
rlabel m2contact 12705 4104 12705 4104 4 stateSub[0]
rlabel m2contact 12681 3288 12681 3288 4 n_32
rlabel m2contact 12681 5424 12681 5424 4 n_188
rlabel m2contact 12657 5160 12657 5160 4 n_222
rlabel m2contact 12633 3264 12633 3264 4 MemEn
rlabel m2contact 12633 3432 12633 3432 4 n_205
rlabel m2contact 12609 3888 12609 3888 4 n_86
rlabel m2contact 12585 5160 12585 5160 4 n_6
rlabel m2contact 12561 2472 12561 2472 4 n_238
rlabel m2contact 12561 3216 12561 3216 4 n_237
rlabel m2contact 12537 3192 12537 3192 4 n_114
rlabel m2contact 12513 3552 12513 3552 4 n_232
rlabel m2contact 12489 6504 12489 6504 4 n_148
rlabel m2contact 12465 5808 12465 5808 4 n_158
rlabel m2contact 12441 6864 12441 6864 4 OpcodeCondIn[7]
rlabel m2contact 12441 3456 12441 3456 4 n_193
rlabel m2contact 12417 3648 12417 3648 4 n_259
rlabel m2contact 12393 6936 12393 6936 4 n_124
rlabel m2contact 12393 2256 12393 2256 4 n_124
rlabel m2contact 12369 3264 12369 3264 4 Rs1Sel[0]
rlabel m2contact 12369 2400 12369 2400 4 n_145
rlabel m2contact 12345 2136 12345 2136 4 n_105
rlabel m2contact 12321 2856 12321 2856 4 n_161
rlabel m2contact 12297 2352 12297 2352 4 n_192
rlabel m2contact 12297 3312 12297 3312 4 n_172
rlabel m2contact 12273 6024 12273 6024 4 n_128
rlabel m2contact 12249 3960 12249 3960 4 state[0]
rlabel m2contact 12225 3456 12225 3456 4 n_193
rlabel m2contact 12201 6024 12201 6024 4 n_73
rlabel m2contact 12177 3264 12177 3264 4 Rs1Sel[0]
rlabel m2contact 12177 3648 12177 3648 4 n_259
rlabel m2contact 12153 2520 12153 2520 4 n_268
rlabel m2contact 12153 4104 12153 4104 4 stateSub[0]
rlabel m2contact 12129 3264 12129 3264 4 n_291
rlabel m2contact 12129 3960 12129 3960 4 state[0]
rlabel m2contact 12105 3192 12105 3192 4 n_114
rlabel m2contact 12081 2856 12081 2856 4 n_261
rlabel m2contact 12057 3480 12057 3480 4 n_317
rlabel m2contact 12033 3336 12033 3336 4 n_23
rlabel m2contact 12009 6912 12009 6912 4 OpcodeCondIn[2]
rlabel m2contact 12009 3960 12009 3960 4 state[0]
rlabel m2contact 11985 6960 11985 6960 4 n_270
rlabel m2contact 11985 3768 11985 3768 4 state[1]
rlabel m2contact 11961 6912 11961 6912 4 n_220
rlabel m2contact 11961 3024 11961 3024 4 n_220
rlabel m2contact 11937 6936 11937 6936 4 n_124
rlabel m2contact 11937 4296 11937 4296 4 n_71
rlabel m2contact 11913 3648 11913 3648 4 n_259
rlabel m2contact 11889 6912 11889 6912 4 n_220
rlabel m2contact 11889 5328 11889 5328 4 n_236
rlabel m2contact 11865 5808 11865 5808 4 n_158
rlabel m2contact 11841 6672 11841 6672 4 n_277
rlabel m2contact 11817 6648 11817 6648 4 n_308
rlabel m2contact 11793 6912 11793 6912 4 n_256
rlabel m2contact 11793 4968 11793 4968 4 n_256
rlabel m2contact 11769 1896 11769 1896 4 n_90
rlabel m2contact 11769 5328 11769 5328 4 n_236
rlabel m2contact 11745 6912 11745 6912 4 n_256
rlabel m2contact 11745 6072 11745 6072 4 n_208
rlabel m2contact 11721 6648 11721 6648 4 OpcodeCondIn[5]
rlabel m2contact 11721 3168 11721 3168 4 OpcodeCondIn[5]
rlabel m2contact 11697 1896 11697 1896 4 n_140
rlabel m2contact 11673 6648 11673 6648 4 OpcodeCondIn[5]
rlabel m2contact 11673 5904 11673 5904 4 n_264
rlabel m2contact 11649 1848 11649 1848 4 n_263
rlabel m2contact 11649 6888 11649 6888 4 n_103
rlabel m2contact 11625 6648 11625 6648 4 n_35
rlabel m2contact 11601 1992 11601 1992 4 n_25
rlabel m2contact 11601 6768 11601 6768 4 n_257
rlabel m2contact 11553 3528 11553 3528 4 n_102
rlabel m2contact 11553 3624 11553 3624 4 stateSub[1]
rlabel m2contact 11529 1992 11529 1992 4 n_213
rlabel m2contact 11505 6240 11505 6240 4 n_170
rlabel m2contact 11481 3216 11481 3216 4 n_237
rlabel m2contact 11481 3528 11481 3528 4 n_141
rlabel m2contact 11457 2328 11457 2328 4 n_47
rlabel m2contact 11433 6768 11433 6768 4 n_62
rlabel m2contact 11433 4536 11433 4536 4 n_365
rlabel m2contact 11409 5160 11409 5160 4 n_6
rlabel m2contact 11409 3096 11409 3096 4 n_136
rlabel m2contact 11385 1872 11385 1872 4 n_189
rlabel m2contact 11361 6000 11361 6000 4 n_228
rlabel m2contact 11361 5160 11361 5160 4 n_137
rlabel m2contact 11337 4320 11337 4320 4 n_164
rlabel m2contact 11313 6600 11313 6600 4 n_227
rlabel m2contact 11313 6240 11313 6240 4 n_182
rlabel m2contact 11289 6000 11289 6000 4 n_130
rlabel m2contact 11289 3384 11289 3384 4 n_130
rlabel m2contact 11265 6840 11265 6840 4 n_26
rlabel m2contact 11265 6336 11265 6336 4 n_198
rlabel m2contact 11241 6072 11241 6072 4 n_208
rlabel m2contact 11241 1872 11241 1872 4 n_208
rlabel m2contact 11217 6000 11217 6000 4 n_130
rlabel m2contact 11217 5376 11217 5376 4 n_187
rlabel m2contact 11193 5520 11193 5520 4 n_282
rlabel m2contact 11169 3984 11169 3984 4 stateSub[2]
rlabel m2contact 11145 1872 11145 1872 4 n_208
rlabel m2contact 11145 6000 11145 6000 4 n_81
rlabel m2contact 11121 6120 11121 6120 4 n_75
rlabel m2contact 11097 6528 11097 6528 4 n_89
rlabel m2contact 11049 1896 11049 1896 4 n_140
rlabel m2contact 11049 6120 11049 6120 4 n_120
rlabel m2contact 11025 1920 11025 1920 4 n_63
rlabel m2contact 11025 4008 11025 4008 4 n_202
rlabel m2contact 11001 3624 11001 3624 4 stateSub[1]
rlabel m2contact 10977 1944 10977 1944 4 n_132
rlabel m2contact 10977 5136 10977 5136 4 n_76
rlabel m2contact 10953 3768 10953 3768 4 state[1]
rlabel m2contact 10929 5136 10929 5136 4 n_16
rlabel m2contact 10881 5544 10881 5544 4 OpcodeCondIn[1]
rlabel m2contact 10857 5520 10857 5520 4 n_282
rlabel m2contact 10833 6888 10833 6888 4 n_145
rlabel m2contact 10833 2400 10833 2400 4 n_145
rlabel m2contact 10809 6648 10809 6648 4 n_35
rlabel m2contact 10809 4704 10809 4704 4 n_28
rlabel m2contact 10785 4824 10785 4824 4 n_85
rlabel m2contact 10761 3936 10761 3936 4 n_34
rlabel m2contact 10737 6312 10737 6312 4 n_22
rlabel m2contact 10713 4608 10713 4608 4 n_194
rlabel m2contact 10689 2064 10689 2064 4 n_339
rlabel m2contact 10665 1968 10665 1968 4 AluOR[1]
rlabel m2contact 10665 5352 10665 5352 4 n_324
rlabel m2contact 10641 5568 10641 5568 4 n_328
rlabel m2contact 10641 4608 10641 4608 4 n_286
rlabel m2contact 10617 5232 10617 5232 4 n_266
rlabel m2contact 10593 5064 10593 5064 4 n_300
rlabel m2contact 10593 6312 10593 6312 4 n_345
rlabel m2contact 10569 6648 10569 6648 4 n_262
rlabel m2contact 10545 3840 10545 3840 4 n_312
rlabel m2contact 10521 6840 10521 6840 4 n_283
rlabel m2contact 10521 3192 10521 3192 4 n_114
rlabel m2contact 10497 4752 10497 4752 4 n_200
rlabel m2contact 10473 6864 10473 6864 4 OpcodeCondIn[7]
rlabel m2contact 10449 4752 10449 4752 4 n_67
rlabel m2contact 10425 6888 10425 6888 4 n_145
rlabel m2contact 10425 3840 10425 3840 4 n_278
rlabel m2contact 10401 2016 10401 2016 4 CFlag
rlabel m2contact 10401 2520 10401 2520 4 n_268
rlabel m2contact 10377 6672 10377 6672 4 n_277
rlabel m2contact 10353 5016 10353 5016 4 n_152
rlabel m2contact 10329 1992 10329 1992 4 n_213
rlabel m2contact 10329 6168 10329 6168 4 n_212
rlabel m2contact 10329 2016 10329 2016 4 n_212
rlabel m2contact 10305 6504 10305 6504 4 n_148
rlabel m2contact 10305 3216 10305 3216 4 n_237
rlabel m2contact 10281 2016 10281 2016 4 n_212
rlabel m2contact 10281 5736 10281 5736 4 n_115
rlabel m2contact 10233 5976 10233 5976 4 n_65
rlabel m2contact 10209 2040 10209 2040 4 PcSel[2]
rlabel m2contact 10209 6864 10209 6864 4 OpcodeCondIn[7]
rlabel m2contact 10185 3384 10185 3384 4 n_130
rlabel m2contact 10161 2064 10161 2064 4 n_339
rlabel m2contact 10137 2088 10137 2088 4 nWait
rlabel m2contact 10113 6840 10113 6840 4 n_283
rlabel m2contact 10089 6816 10089 6816 4 n_27
rlabel m2contact 10089 2088 10089 2088 4 nWait
rlabel m2contact 10065 4968 10065 4968 4 n_256
rlabel m2contact 10065 5280 10065 5280 4 n_280
rlabel m2contact 10041 3936 10041 3936 4 n_34
rlabel m2contact 9993 3456 9993 3456 4 n_193
rlabel m2contact 9993 4968 9993 4968 4 n_318
rlabel m2contact 9969 3168 9969 3168 4 OpcodeCondIn[5]
rlabel m2contact 9969 3480 9969 3480 4 n_317
rlabel m2contact 9945 6792 9945 6792 4 SysBus[1]
rlabel m2contact 9945 5376 9945 5376 4 n_187
rlabel m2contact 9897 6768 9897 6768 4 n_62
rlabel m2contact 9897 5904 9897 5904 4 n_264
rlabel m2contact 9873 6744 9873 6744 4 OpcodeCondIn[6]
rlabel m2contact 9873 4104 9873 4104 4 stateSub[0]
rlabel m2contact 9849 6720 9849 6720 4 n_29
rlabel m2contact 9849 3624 9849 3624 4 stateSub[1]
rlabel m2contact 9825 5520 9825 5520 4 n_282
rlabel m2contact 9777 2112 9777 2112 4 n_166
rlabel m2contact 9777 3168 9777 3168 4 n_274
rlabel m2contact 9753 6696 9753 6696 4 StatusReg[3]
rlabel m2contact 9753 3480 9753 3480 4 n_169
rlabel m2contact 9729 6672 9729 6672 4 n_277
rlabel m2contact 9681 6648 9681 6648 4 n_262
rlabel m2contact 9681 3984 9681 3984 4 stateSub[2]
rlabel m2contact 9657 5496 9657 5496 4 n_79
rlabel m2contact 9633 6624 9633 6624 4 n_211
rlabel m2contact 9609 2352 9609 2352 4 n_192
rlabel m2contact 9561 2928 9561 2928 4 n_51
rlabel m2contact 9537 3768 9537 3768 4 state[1]
rlabel m2contact 9513 2544 9513 2544 4 IntReq
rlabel m2contact 9513 3936 9513 3936 4 n_34
rlabel m2contact 9465 4776 9465 4776 4 n_219
rlabel m2contact 9441 2352 9441 2352 4 n_77
rlabel m2contact 9417 4776 9417 4776 4 n_121
rlabel m2contact 9393 2544 9393 2544 4 n_195
rlabel m2contact 9345 6600 9345 6600 4 n_227
rlabel m2contact 9297 5784 9297 5784 4 OpcodeCondIn[4]
rlabel m2contact 9273 3456 9273 3456 4 n_193
rlabel m2contact 9201 4608 9201 4608 4 n_286
rlabel m2contact 9153 2904 9153 2904 4 n_95
rlabel m2contact 9105 2544 9105 2544 4 n_195
rlabel m2contact 9081 6576 9081 6576 4 n_135
rlabel m2contact 9057 6552 9057 6552 4 n_21
rlabel m2contact 9009 2136 9009 2136 4 n_105
rlabel m2contact 8985 5784 8985 5784 4 OpcodeCondIn[4]
rlabel m2contact 8961 6528 8961 6528 4 n_89
rlabel m2contact 8961 3960 8961 3960 4 state[0]
rlabel m2contact 8937 6504 8937 6504 4 n_148
rlabel m2contact 8865 2184 8865 2184 4 n_350
rlabel m2contact 8841 6480 8841 6480 4 n_321
rlabel m2contact 8841 3984 8841 3984 4 stateSub[2]
rlabel m2contact 8817 2160 8817 2160 4 n_224
rlabel m2contact 8793 4800 8793 4800 4 n_91
rlabel m2contact 8793 2184 8793 2184 4 n_91
rlabel m2contact 8769 4392 8769 4392 4 n_83
rlabel m2contact 8745 6456 8745 6456 4 n_122
rlabel m2contact 8745 2400 8745 2400 4 n_145
rlabel m2contact 8721 2184 8721 2184 4 n_91
rlabel m2contact 8721 4392 8721 4392 4 n_290
rlabel m2contact 8673 6432 8673 6432 4 n_13
rlabel m2contact 8649 6408 8649 6408 4 SysBus[2]
rlabel m2contact 8649 5784 8649 5784 4 OpcodeCondIn[4]
rlabel m2contact 8625 5328 8625 5328 4 n_236
rlabel m2contact 8577 2208 8577 2208 4 n_368
rlabel m2contact 8577 5616 8577 5616 4 n_235
rlabel m2contact 8553 6384 8553 6384 4 n_320
rlabel m2contact 8529 6360 8529 6360 4 n_335
rlabel m2contact 8505 2712 8505 2712 4 StatusReg[2]
rlabel m2contact 8457 2232 8457 2232 4 n_175
rlabel m2contact 8457 5592 8457 5592 4 n_347
rlabel m2contact 8433 4920 8433 4920 4 n_346
rlabel m2contact 8433 4296 8433 4296 4 n_71
rlabel m2contact 8409 2256 8409 2256 4 n_124
rlabel m2contact 8409 5592 8409 5592 4 n_329
rlabel m2contact 8361 3384 8361 3384 4 n_130
rlabel m2contact 8337 5640 8337 5640 4 n_244
rlabel m2contact 8337 2256 8337 2256 4 n_244
rlabel m2contact 8313 2256 8313 2256 4 n_244
rlabel m2contact 8313 5544 8313 5544 4 OpcodeCondIn[1]
rlabel m2contact 8289 4440 8289 4440 4 OpcodeCondIn[0]
rlabel m2contact 8265 4848 8265 4848 4 n_364
rlabel m2contact 8241 4848 8241 4848 4 n_364
rlabel m2contact 8217 4008 8217 4008 4 n_202
rlabel m2contact 8193 6336 8193 6336 4 n_198
rlabel m2contact 8193 3360 8193 3360 4 OpcodeCondIn[2]
rlabel m2contact 8169 5088 8169 5088 4 OpcodeCondIn[3]
rlabel m2contact 8121 2280 8121 2280 4 n_352
rlabel m2contact 8097 2304 8097 2304 4 n_270
rlabel m2contact 8073 6312 8073 6312 4 n_345
rlabel m2contact 8049 5064 8049 5064 4 n_300
rlabel m2contact 8001 2520 8001 2520 4 n_268
rlabel m2contact 7953 3624 7953 3624 4 stateSub[1]
rlabel m2contact 7929 5064 7929 5064 4 n_133
rlabel m2contact 7905 3768 7905 3768 4 state[1]
rlabel m2contact 7881 2328 7881 2328 4 n_47
rlabel m2contact 7881 3960 7881 3960 4 state[0]
rlabel m2contact 7857 5088 7857 5088 4 OpcodeCondIn[3]
rlabel m2contact 7809 4920 7809 4920 4 n_346
rlabel m2contact 7785 6288 7785 6288 4 n_336
rlabel m2contact 7785 6072 7785 6072 4 n_208
rlabel m2contact 7761 4848 7761 4848 4 n_364
rlabel m2contact 7737 2400 7737 2400 4 n_145
rlabel m2contact 7737 4536 7737 4536 4 n_365
rlabel m2contact 7713 6144 7713 6144 4 n_310
rlabel m2contact 7689 4848 7689 4848 4 n_355
rlabel m2contact 7665 2352 7665 2352 4 n_77
rlabel m2contact 7665 2376 7665 2376 4 n_150
rlabel m2contact 7641 2400 7641 2400 4 n_145
rlabel m2contact 7641 2760 7641 2760 4 n_250
rlabel m2contact 7617 6264 7617 6264 4 n_319
rlabel m2contact 7617 3936 7617 3936 4 n_34
rlabel m2contact 7593 6240 7593 6240 4 n_182
rlabel m2contact 7593 5760 7593 5760 4 n_129
rlabel m2contact 7593 2400 7593 2400 4 n_129
rlabel m2contact 7569 2760 7569 2760 4 n_149
rlabel m2contact 7545 5472 7545 5472 4 n_40
rlabel m2contact 7521 2400 7521 2400 4 n_129
rlabel m2contact 7521 4128 7521 4128 4 n_59
rlabel m2contact 7497 3624 7497 3624 4 stateSub[1]
rlabel m2contact 7473 5064 7473 5064 4 n_133
rlabel m2contact 7449 2424 7449 2424 4 n_294
rlabel m2contact 7425 6216 7425 6216 4 n_54
rlabel m2contact 7425 3384 7425 3384 4 n_130
rlabel m2contact 7401 6192 7401 6192 4 n_240
rlabel m2contact 7401 3024 7401 3024 4 n_220
rlabel m2contact 7353 2448 7353 2448 4 n_276
rlabel m2contact 7353 2472 7353 2472 4 n_238
rlabel m2contact 7329 5328 7329 5328 4 n_236
rlabel m2contact 7329 4008 7329 4008 4 n_202
rlabel m2contact 7305 6168 7305 6168 4 n_212
rlabel m2contact 7281 4104 7281 4104 4 stateSub[0]
rlabel m2contact 7257 2496 7257 2496 4 n_196
rlabel m2contact 7257 3216 7257 3216 4 n_237
rlabel m2contact 7233 2520 7233 2520 4 n_268
rlabel m2contact 7209 2544 7209 2544 4 n_195
rlabel m2contact 7209 6144 7209 6144 4 n_310
rlabel m2contact 7161 4512 7161 4512 4 n_288
rlabel m2contact 7137 3744 7137 3744 4 n_258
rlabel m2contact 7137 3960 7137 3960 4 state[0]
rlabel m2contact 7089 2568 7089 2568 4 n_209
rlabel m2contact 7089 2592 7089 2592 4 n_156
rlabel m2contact 7065 3960 7065 3960 4 state[0]
rlabel m2contact 7041 6120 7041 6120 4 n_120
rlabel m2contact 6993 6096 6993 6096 4 n_44
rlabel m2contact 6993 3984 6993 3984 4 stateSub[2]
rlabel m2contact 6969 2832 6969 2832 4 n_7
rlabel m2contact 6945 3864 6945 3864 4 n_14
rlabel m2contact 6921 5664 6921 5664 4 n_243
rlabel m2contact 6897 2832 6897 2832 4 Op2Sel[0]
rlabel m2contact 6873 4032 6873 4032 4 n_49
rlabel m2contact 6849 3864 6849 3864 4 n_181
rlabel m2contact 6825 5664 6825 5664 4 n_243
rlabel m2contact 6801 5304 6801 5304 4 n_178
rlabel m2contact 6777 6072 6777 6072 4 n_208
rlabel m2contact 6753 2664 6753 2664 4 n_184
rlabel m2contact 6729 2688 6729 2688 4 n_296
rlabel m2contact 6681 4176 6681 4176 4 n_271
rlabel m2contact 6657 5208 6657 5208 4 n_272
rlabel m2contact 6657 4296 6657 4296 4 n_71
rlabel m2contact 6585 6048 6585 6048 4 n_80
rlabel m2contact 6585 3984 6585 3984 4 stateSub[2]
rlabel m2contact 6561 3120 6561 3120 4 n_78
rlabel m2contact 6537 6048 6537 6048 4 n_130
rlabel m2contact 6537 3384 6537 3384 4 n_130
rlabel m2contact 6513 6048 6513 6048 4 n_130
rlabel m2contact 6513 4176 6513 4176 4 nME
rlabel m2contact 6489 3360 6489 3360 4 OpcodeCondIn[2]
rlabel m2contact 6441 2616 6441 2616 4 n_33
rlabel m2contact 6441 3360 6441 3360 4 n_176
rlabel m2contact 6441 2664 6441 2664 4 n_176
rlabel m2contact 6417 3360 6417 3360 4 n_176
rlabel m2contact 6417 2688 6417 2688 4 n_10
rlabel m2contact 6393 2640 6393 2640 4 n_123
rlabel m2contact 6369 3360 6369 3360 4 n_229
rlabel m2contact 6369 3624 6369 3624 4 stateSub[1]
rlabel m2contact 6345 2664 6345 2664 4 n_176
rlabel m2contact 6345 3312 6345 3312 4 n_172
rlabel m2contact 6321 6024 6321 6024 4 n_73
rlabel m2contact 6297 6000 6297 6000 4 n_81
rlabel m2contact 6273 4680 6273 4680 4 n_106
rlabel m2contact 6225 5904 6225 5904 4 n_264
rlabel m2contact 6177 2688 6177 2688 4 n_10
rlabel m2contact 6153 5280 6153 5280 4 n_280
rlabel m2contact 6129 2712 6129 2712 4 StatusReg[2]
rlabel m2contact 6129 3768 6129 3768 4 state[1]
rlabel m2contact 6081 2736 6081 2736 4 n_104
rlabel m2contact 6057 5976 6057 5976 4 n_65
rlabel m2contact 6033 2952 6033 2952 4 n_125
rlabel m2contact 6009 3312 6009 3312 4 n_172
rlabel m2contact 5961 5952 5961 5952 4 n_214
rlabel m2contact 5937 4512 5937 4512 4 n_288
rlabel m2contact 5913 2760 5913 2760 4 n_149
rlabel m2contact 5865 5928 5865 5928 4 n_265
rlabel m2contact 5841 5664 5841 5664 4 n_243
rlabel m2contact 5817 3744 5817 3744 4 n_258
rlabel m2contact 5793 5904 5793 5904 4 n_264
rlabel m2contact 5745 2784 5745 2784 4 n_94
rlabel m2contact 5721 5880 5721 5880 4 n_359
rlabel m2contact 5697 4104 5697 4104 4 stateSub[0]
rlabel m2contact 5673 5832 5673 5832 4 n_93
rlabel m2contact 5625 5856 5625 5856 4 n_332
rlabel metal2 5601 5832 5601 5832 4 Flags[2]
rlabel m2contact 5577 3912 5577 3912 4 n_333
rlabel m2contact 5505 5808 5505 5808 4 n_158
rlabel m2contact 5457 5784 5457 5784 4 OpcodeCondIn[4]
rlabel m2contact 5409 2808 5409 2808 4 n_8
rlabel m2contact 5409 5760 5409 5760 4 n_129
rlabel m2contact 5385 3192 5385 3192 4 n_114
rlabel m2contact 5361 5736 5361 5736 4 n_115
rlabel m2contact 5361 4440 5361 4440 4 OpcodeCondIn[0]
rlabel m2contact 5313 2832 5313 2832 4 Op2Sel[0]
rlabel m2contact 5313 2856 5313 2856 4 n_261
rlabel m2contact 5289 3192 5289 3192 4 n_165
rlabel m2contact 5289 3984 5289 3984 4 stateSub[2]
rlabel m2contact 5265 2880 5265 2880 4 n_199
rlabel m2contact 5265 5712 5265 5712 4 n_204
rlabel m2contact 5217 5688 5217 5688 4 n_245
rlabel m2contact 5193 2904 5193 2904 4 n_95
rlabel m2contact 5193 5664 5193 5664 4 n_243
rlabel m2contact 5169 5640 5169 5640 4 n_244
rlabel m2contact 5145 3624 5145 3624 4 stateSub[1]
rlabel m2contact 5121 2928 5121 2928 4 n_51
rlabel m2contact 5097 5616 5097 5616 4 n_235
rlabel m2contact 5073 2952 5073 2952 4 n_125
rlabel m2contact 5049 2976 5049 2976 4 n_174
rlabel m2contact 5001 5592 5001 5592 4 n_329
rlabel m2contact 5001 3960 5001 3960 4 state[0]
rlabel m2contact 4977 5568 4977 5568 4 n_328
rlabel m2contact 4953 3000 4953 3000 4 InISR
rlabel m2contact 4929 3024 4929 3024 4 n_220
rlabel m2contact 4905 3048 4905 3048 4 n_55
rlabel m2contact 4881 3048 4881 3048 4 n_55
rlabel m2contact 4881 5544 4881 5544 4 OpcodeCondIn[1]
rlabel m2contact 4857 5520 4857 5520 4 n_282
rlabel m2contact 4833 3072 4833 3072 4 n_138
rlabel m2contact 4833 4440 4833 4440 4 OpcodeCondIn[0]
rlabel m2contact 4809 3096 4809 3096 4 n_136
rlabel m2contact 4785 5160 4785 5160 4 n_137
rlabel m2contact 4761 3216 4761 3216 4 n_237
rlabel m2contact 4713 5088 4713 5088 4 OpcodeCondIn[3]
rlabel m2contact 4665 3120 4665 3120 4 n_78
rlabel m2contact 4665 5496 4665 5496 4 n_79
rlabel m2contact 4617 3144 4617 3144 4 n_356
rlabel m2contact 4617 3960 4617 3960 4 state[0]
rlabel m2contact 4593 5472 4593 5472 4 n_40
rlabel m2contact 4545 3168 4545 3168 4 n_274
rlabel m2contact 4545 3192 4545 3192 4 n_165
rlabel m2contact 4521 4320 4521 4320 4 n_164
rlabel m2contact 4497 5376 4497 5376 4 n_187
rlabel m2contact 4473 3216 4473 3216 4 n_237
rlabel m2contact 4473 3240 4473 3240 4 n_37
rlabel m2contact 4449 4128 4449 4128 4 n_59
rlabel m2contact 4425 3264 4425 3264 4 n_291
rlabel m2contact 4401 3288 4401 3288 4 n_32
rlabel m2contact 4377 3312 4377 3312 4 n_172
rlabel m2contact 4377 5448 4377 5448 4 n_11
rlabel m2contact 4353 3336 4353 3336 4 n_23
rlabel m2contact 4353 3360 4353 3360 4 n_229
rlabel m2contact 4305 5424 4305 5424 4 n_188
rlabel m2contact 4281 3384 4281 3384 4 n_130
rlabel m2contact 4281 5400 4281 5400 4 n_154
rlabel m2contact 4257 3408 4257 3408 4 n_45
rlabel m2contact 4257 5376 4257 5376 4 n_187
rlabel m2contact 4209 3432 4209 3432 4 n_205
rlabel m2contact 4185 3600 4185 3600 4 n_292
rlabel m2contact 4185 3648 4185 3648 4 n_259
rlabel m2contact 4161 3432 4161 3432 4 n_167
rlabel m2contact 4089 3432 4089 3432 4 n_167
rlabel m2contact 4089 3600 4089 3600 4 n_260
rlabel m2contact 4065 5352 4065 5352 4 n_324
rlabel m2contact 4041 3456 4041 3456 4 n_193
rlabel m2contact 4017 3480 4017 3480 4 n_169
rlabel m2contact 3993 3504 3993 3504 4 n_230
rlabel m2contact 3993 5328 3993 5328 4 n_236
rlabel m2contact 3969 3528 3969 3528 4 n_141
rlabel m2contact 3969 5304 3969 5304 4 n_178
rlabel m2contact 3945 3552 3945 3552 4 n_232
rlabel m2contact 3921 3576 3921 3576 4 n_153
rlabel m2contact 3897 3600 3897 3600 4 n_260
rlabel m2contact 3897 5280 3897 5280 4 n_280
rlabel m2contact 3873 5016 3873 5016 4 n_152
rlabel m2contact 3849 3744 3849 3744 4 n_258
rlabel m2contact 3825 3624 3825 3624 4 stateSub[1]
rlabel m2contact 3801 3648 3801 3648 4 n_259
rlabel m2contact 3801 5016 3801 5016 4 n_360
rlabel m2contact 3753 3672 3753 3672 4 n_87
rlabel m2contact 3753 5256 3753 5256 4 n_353
rlabel m2contact 3681 3816 3681 3816 4 n_96
rlabel m2contact 3681 4608 3681 4608 4 n_286
rlabel m2contact 3657 5232 3657 5232 4 n_266
rlabel m2contact 3633 3816 3633 3816 4 n_334
rlabel m2contact 3609 3696 3609 3696 4 n_299
rlabel m2contact 3585 3912 3585 3912 4 n_333
rlabel m2contact 3561 5208 3561 5208 4 n_272
rlabel m2contact 3537 3720 3537 3720 4 n_239
rlabel m2contact 3537 5184 3537 5184 4 n_248
rlabel m2contact 3489 5160 3489 5160 4 n_137
rlabel m2contact 3465 3744 3465 3744 4 n_258
rlabel m2contact 3441 5136 3441 5136 4 n_16
rlabel m2contact 3417 4464 3417 4464 4 n_99
rlabel m2contact 3369 5112 3369 5112 4 n_134
rlabel m2contact 3345 5088 3345 5088 4 OpcodeCondIn[3]
rlabel m2contact 3321 3768 3321 3768 4 state[1]
rlabel m2contact 3321 5064 3321 5064 4 n_133
rlabel m2contact 3273 4512 3273 4512 4 n_288
rlabel m2contact 3249 5040 3249 5040 4 n_348
rlabel m2contact 3225 5016 3225 5016 4 n_360
rlabel m2contact 3201 4584 3201 4584 4 n_361
rlabel m2contact 3177 3792 3177 3792 4 n_281
rlabel m2contact 3129 4992 3129 4992 4 n_363
rlabel m2contact 3105 4968 3105 4968 4 n_318
rlabel m2contact 3081 3816 3081 3816 4 n_334
rlabel m2contact 3057 3840 3057 3840 4 n_278
rlabel m2contact 3009 4944 3009 4944 4 n_301
rlabel m2contact 2961 4920 2961 4920 4 n_346
rlabel m2contact 2937 3864 2937 3864 4 n_181
rlabel m2contact 2913 4896 2913 4896 4 n_162
rlabel m2contact 2889 3864 2889 3864 4 LrSel
rlabel m2contact 2817 4872 2817 4872 4 n_367
rlabel m2contact 2769 3864 2769 3864 4 LrSel
rlabel m2contact 2769 4848 2769 4848 4 n_355
rlabel m2contact 2721 3888 2721 3888 4 n_86
rlabel m2contact 2697 4824 2697 4824 4 n_85
rlabel m2contact 2673 4800 2673 4800 4 n_91
rlabel m2contact 2625 3912 2625 3912 4 n_333
rlabel m2contact 2625 4776 2625 4776 4 n_121
rlabel m2contact 2601 3984 2601 3984 4 stateSub[2]
rlabel m2contact 2577 3936 2577 3936 4 n_34
rlabel m2contact 2577 4752 2577 4752 4 n_67
rlabel m2contact 2529 4728 2529 4728 4 n_42
rlabel m2contact 2529 3960 2529 3960 4 state[0]
rlabel m2contact 2505 4704 2505 4704 4 n_28
rlabel m2contact 2505 3984 2505 3984 4 stateSub[2]
rlabel m2contact 2481 4680 2481 4680 4 n_106
rlabel m2contact 2409 4656 2409 4656 4 n_223
rlabel m2contact 2409 4008 2409 4008 4 n_202
rlabel m2contact 2361 4632 2361 4632 4 n_159
rlabel m2contact 2313 4296 2313 4296 4 n_71
rlabel m2contact 2289 4608 2289 4608 4 n_286
rlabel m2contact 2289 4032 2289 4032 4 n_49
rlabel m2contact 2265 4056 2265 4056 4 n_330
rlabel m2contact 2241 4584 2241 4584 4 n_361
rlabel m2contact 2241 4560 2241 4560 4 Flags[0]
rlabel m2contact 2217 4536 2217 4536 4 n_365
rlabel m2contact 2169 4080 2169 4080 4 n_311
rlabel m2contact 2145 4512 2145 4512 4 n_288
rlabel m2contact 2121 4488 2121 4488 4 n_242
rlabel m2contact 2097 4104 2097 4104 4 stateSub[0]
rlabel m2contact 2049 4128 2049 4128 4 n_59
rlabel m2contact 2049 4224 2049 4224 4 n_3
rlabel m2contact 2001 4224 2001 4224 4 nIRQ
rlabel m2contact 1953 4464 1953 4464 4 n_99
rlabel m2contact 1905 4440 1905 4440 4 OpcodeCondIn[0]
rlabel m2contact 1881 4416 1881 4416 4 n_43
rlabel m2contact 1833 4392 1833 4392 4 n_290
rlabel m2contact 1809 4368 1809 4368 4 n_246
rlabel m2contact 1785 4152 1785 4152 4 n_226
rlabel m2contact 1737 4176 1737 4176 4 nME
rlabel m2contact 1689 4344 1689 4344 4 n_144
rlabel m2contact 1665 4320 1665 4320 4 n_164
rlabel m2contact 1617 4296 1617 4296 4 n_71
rlabel metal2 25695 8170 25707 8170 6 MemEn
rlabel metal2 24195 8170 24207 8170 6 IrWe
rlabel metal2 22695 8170 22707 8170 6 LrSel
rlabel metal2 22215 8170 22227 8170 6 LrWe
rlabel metal2 20559 8170 20571 8170 6 WdSel
rlabel metal2 18195 8170 18207 8170 6 LrEn
rlabel metal2 18171 8170 18183 8170 6 PcSel[0]
rlabel metal2 15195 8170 15207 8170 6 PcSel[1]
rlabel metal2 14463 8170 14475 8170 6 PcSel[2]
rlabel metal2 12183 8170 12195 8170 4 PcEn
rlabel metal2 12147 8170 12159 8170 4 PcWe
rlabel metal2 10635 8170 10647 8170 4 Op1Sel
rlabel metal2 9123 8170 9135 8170 4 ImmSel
rlabel metal2 6903 8170 6915 8170 4 Op2Sel[0]
rlabel metal2 4623 8170 4635 8170 4 Op2Sel[1]
rlabel metal2 4587 8170 4599 8170 4 AluWe
rlabel metal2 3075 8170 3087 8170 4 AluEn
rlabel metal2 27649 145 27649 157 8 OpcodeCondIn[0]
rlabel metal2 27649 97 27649 109 8 OpcodeCondIn[2]
rlabel metal2 27649 73 27649 85 8 OpcodeCondIn[7]
rlabel metal2 27649 49 27649 61 8 OpcodeCondIn[6]
rlabel metal2 27649 25 27649 37 8 OpcodeCondIn[4]
rlabel metal2 27649 1 27649 13 8 OpcodeCondIn[5]
rlabel metal2 27649 1962 27649 1974 6 AluOR[1]
rlabel metal2 27649 1938 27649 1950 6 SysBus[1]
rlabel metal2 27649 1914 27649 1926 6 SysBus[0]
rlabel metal2 27649 1890 27649 1902 6 SysBus[3]
rlabel metal2 27649 1866 27649 1878 6 SysBus[2]
rlabel metal2 27649 1842 27649 1854 6 OpcodeCondIn[3]
rlabel metal2 27649 1818 27649 1830 6 OpcodeCondIn[1]
rlabel metal2 27649 8027 27649 8039 6 CFlag
rlabel metal2 27649 8003 27649 8015 6 RegWe
rlabel metal2 27649 7979 27649 7991 6 RwSel[0]
rlabel metal2 27649 7955 27649 7967 6 Rs1Sel[1]
rlabel metal2 27649 7931 27649 7943 6 RwSel[1]
rlabel metal2 27649 7907 27649 7919 6 Rs1Sel[0]
rlabel metal2 27649 7883 27649 7895 6 AluOR[0]
rlabel m2contact 27054 7961 27054 7961 6 Rs1Sel[1]
rlabel m2contact 27054 8009 27054 8009 6 Rs1Sel[1]
rlabel m2contact 27105 8009 27105 8009 6 RegWe
rlabel m2contact 27153 8009 27153 8009 6 RegWe
rlabel m2contact 27026 8033 27026 8033 6 CFlag
rlabel m2contact 27027 7985 27027 7985 6 CFlag
rlabel m2contact 27132 7889 27132 7889 6 RwSel[0]
rlabel m2contact 27132 7985 27132 7985 6 RwSel[0]
rlabel m2contact 27161 7937 27161 7937 6 AluOR[0]
rlabel m2contact 27161 7889 27161 7889 6 AluOR[0]
rlabel m2contact 27185 7937 27185 7937 6 RwSel[1]
rlabel m2contact 27185 8105 27185 8105 6 RwSel[1]
rlabel metal2 27243 8170 27443 8170 5 GND!
rlabel metal2 27243 0 27443 0 1 GND!
rlabel metal2 0 121 0 133 2 Flags[1]
rlabel metal2 0 97 0 109 2 Flags[3]
rlabel metal2 0 73 0 85 2 Flags[2]
rlabel metal2 0 49 0 61 2 Flags[0]
rlabel metal2 0 4266 0 4278 4 nOE
rlabel metal2 0 4242 0 4254 4 nWE
rlabel metal2 0 4218 0 4230 4 nIRQ
rlabel metal2 0 4194 0 4206 4 ENB
rlabel metal2 0 8027 0 8039 4 ALE
rlabel metal2 0 8003 0 8015 4 nME
rlabel metal2 0 7979 0 7991 4 nWait
rlabel metal2 124 0 324 0 1 Vdd!
rlabel metal2 123 8170 323 8170 5 Vdd!
rlabel metal2 339 8170 351 8170 5 SDO
rlabel metal2 363 8170 375 8170 5 Test
rlabel metal2 387 8170 399 8170 5 Clock
rlabel metal2 411 8170 423 8170 5 nReset
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 339 0 351 0 1 SDI
<< end >>
