magic
tech c035u
timestamp 1393514645
<< metal1 >>
rect 614 1144 743 1154
rect 757 1144 1895 1154
rect 1909 1144 3047 1154
rect 3062 1144 4199 1154
rect 4213 1144 5351 1154
rect 5365 1144 6503 1154
rect 6517 1144 7654 1154
rect 7669 1144 8807 1154
rect 1332 1094 1463 1104
rect 1477 1094 1679 1104
rect 2484 1094 2615 1104
rect 2629 1094 2831 1104
rect 3636 1094 3767 1104
rect 3781 1094 3983 1104
rect 4788 1094 4919 1104
rect 4933 1094 5135 1104
rect 5940 1094 6071 1104
rect 6085 1094 6287 1104
rect 7092 1094 7223 1104
rect 7237 1094 7439 1104
rect 8244 1094 8375 1104
rect 8389 1094 8591 1104
rect 9396 1094 9527 1104
rect 9541 1094 9743 1104
rect 0 75 23 85
rect 37 75 9937 85
rect 0 40 1606 50
rect 1621 40 2758 50
rect 2773 40 3910 50
rect 3925 40 5063 50
rect 5078 40 6213 50
rect 6231 40 7365 50
rect 7383 40 8517 50
rect 8535 40 9671 50
rect 9685 40 9952 50
rect 0 5 1823 15
rect 1837 5 2975 15
rect 2989 5 4127 15
rect 4141 5 5279 15
rect 5294 5 6430 15
rect 6448 5 7582 15
rect 7600 5 8734 15
rect 8752 5 9887 15
rect 9901 5 9917 15
<< m2contact >>
rect 598 1139 614 1155
rect 743 1141 757 1155
rect 1895 1143 1909 1157
rect 3047 1143 3062 1157
rect 4199 1143 4213 1157
rect 5351 1143 5365 1157
rect 6503 1143 6517 1157
rect 7654 1142 7669 1156
rect 8807 1143 8822 1158
rect 1318 1092 1332 1106
rect 1463 1091 1477 1105
rect 1679 1091 1693 1105
rect 2470 1092 2484 1106
rect 2615 1091 2629 1105
rect 2831 1092 2845 1106
rect 3622 1092 3636 1106
rect 3767 1091 3781 1105
rect 3983 1092 3997 1106
rect 4774 1092 4788 1106
rect 4919 1091 4933 1105
rect 5135 1092 5149 1106
rect 5926 1092 5940 1106
rect 6071 1091 6085 1105
rect 6287 1092 6301 1106
rect 7078 1092 7092 1106
rect 7223 1091 7237 1105
rect 7439 1092 7453 1106
rect 8230 1092 8244 1106
rect 8375 1091 8389 1105
rect 8591 1092 8605 1106
rect 9382 1092 9396 1106
rect 9527 1091 9541 1105
rect 9743 1092 9757 1106
rect 23 74 37 88
rect 1606 38 1621 52
rect 2758 38 2773 52
rect 3910 38 3925 52
rect 5063 38 5078 53
rect 6213 38 6231 53
rect 7365 38 7383 53
rect 8517 38 8535 53
rect 9671 37 9685 52
rect 1823 4 1837 18
rect 2975 4 2989 18
rect 4127 4 4141 18
rect 5279 3 5294 18
rect 6430 0 6448 15
rect 7582 0 7600 15
rect 8734 0 8752 15
rect 9887 3 9901 18
<< metal2 >>
rect 24 1068 36 1194
rect 72 1068 84 1194
rect 600 1068 612 1139
rect 744 1068 756 1141
rect 792 1068 804 1194
rect 1320 1068 1332 1092
rect 1464 1068 1476 1091
rect 1536 1068 1548 1194
rect 1608 1068 1620 1194
rect 1680 1068 1692 1091
rect 1752 1068 1764 1194
rect 1824 1068 1836 1194
rect 1896 1068 1908 1143
rect 1944 1068 1956 1194
rect 2472 1068 2484 1092
rect 2616 1068 2628 1091
rect 2688 1068 2700 1194
rect 2760 1068 2772 1194
rect 2832 1068 2844 1092
rect 2904 1068 2916 1194
rect 2976 1068 2988 1194
rect 3048 1068 3060 1143
rect 3096 1068 3108 1194
rect 3624 1068 3636 1092
rect 3768 1068 3780 1091
rect 3840 1068 3852 1194
rect 3912 1068 3924 1194
rect 3984 1068 3996 1092
rect 4056 1068 4068 1194
rect 4128 1068 4140 1194
rect 4200 1068 4212 1143
rect 4248 1068 4260 1194
rect 4776 1068 4788 1092
rect 4920 1068 4932 1091
rect 4992 1068 5004 1194
rect 5064 1068 5076 1194
rect 5136 1068 5148 1092
rect 5208 1068 5220 1194
rect 5280 1068 5292 1194
rect 5352 1068 5364 1143
rect 5400 1068 5412 1194
rect 5928 1068 5940 1092
rect 6072 1068 6084 1091
rect 6144 1068 6156 1194
rect 6216 1068 6228 1194
rect 6288 1068 6300 1092
rect 6360 1068 6372 1194
rect 6432 1068 6444 1194
rect 6504 1068 6516 1143
rect 6552 1068 6564 1194
rect 7080 1068 7092 1092
rect 7224 1068 7236 1091
rect 7296 1068 7308 1194
rect 7368 1068 7380 1194
rect 7440 1068 7452 1092
rect 7512 1068 7524 1194
rect 7584 1068 7596 1194
rect 7656 1068 7668 1142
rect 7704 1068 7716 1194
rect 8232 1068 8244 1092
rect 8376 1068 8388 1091
rect 8448 1068 8460 1194
rect 8520 1068 8532 1194
rect 8592 1068 8604 1092
rect 8664 1068 8676 1194
rect 8736 1068 8748 1194
rect 8808 1068 8820 1143
rect 8856 1068 8868 1194
rect 9384 1068 9396 1092
rect 9528 1068 9540 1091
rect 9600 1068 9612 1194
rect 9672 1068 9684 1194
rect 9744 1068 9756 1092
rect 9816 1068 9828 1194
rect 9888 1068 9900 1194
rect 24 88 36 269
rect 1608 52 1620 269
rect 1824 18 1836 269
rect 2760 52 2772 269
rect 2976 18 2988 269
rect 3912 52 3924 269
rect 4128 18 4140 269
rect 5064 53 5076 269
rect 5280 18 5292 269
rect 6216 53 6228 269
rect 6432 15 6444 269
rect 7368 53 7380 269
rect 7584 15 7596 269
rect 8520 53 8532 269
rect 8736 15 8748 269
rect 9672 52 9684 269
rect 9888 18 9900 269
use scanreg scanreg_0
timestamp 1386241447
transform 1 0 0 0 1 269
box 0 0 720 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 720 0 1 269
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 1440 0 1 269
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 1656 0 1 269
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 1872 0 1 269
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 2592 0 1 269
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2808 0 1 269
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 3024 0 1 269
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3744 0 1 269
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3960 0 1 269
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 4176 0 1 269
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4896 0 1 269
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 5112 0 1 269
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 5328 0 1 269
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 6048 0 1 269
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 6264 0 1 269
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 6480 0 1 269
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 7200 0 1 269
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 7416 0 1 269
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 7632 0 1 269
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 8352 0 1 269
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 8568 0 1 269
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 8784 0 1 269
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 9504 0 1 269
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9720 0 1 269
box 0 0 216 799
<< labels >>
rlabel metal2 72 1194 84 1194 5 IRWc
rlabel metal2 792 1194 804 1194 5 WData[0]
rlabel metal2 1944 1194 1956 1194 5 WData[1]
rlabel metal2 3096 1194 3108 1194 5 WData[2]
rlabel metal2 4248 1194 4260 1194 5 WData[3]
rlabel metal2 5400 1194 5412 1194 5 WData[4]
rlabel metal2 6552 1194 6564 1194 5 WData[5]
rlabel metal2 7704 1194 7716 1194 5 WData[6]
rlabel metal2 8856 1194 8868 1194 5 WData[7]
<< end >>
