../behavioural/cpu_core.sv