../../../Design/Implementation/verilog/behavioural/io_switches.sv