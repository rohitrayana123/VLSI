magic
tech c035u
timestamp 1395929667
<< metal4 >>
rect 6616 44286 8176 45846
rect 10142 44286 11702 45846
rect 13668 44286 15228 45846
rect 17194 44286 18754 45846
rect 20720 44286 22280 45846
rect 24246 44286 25806 45846
rect 27772 44286 29332 45846
rect 31298 44286 32858 45846
rect 34824 44286 36384 45846
rect 78 37834 1638 39394
rect 41362 37834 42922 39394
rect 78 33362 1638 34922
rect 41362 33362 42922 34922
rect 78 28890 1638 30450
rect 41362 28890 42922 30450
rect 78 24418 1638 25978
rect 41362 24418 42922 25978
rect 78 19946 1638 21506
rect 41362 19946 42922 21506
rect 78 15474 1638 17034
rect 41362 15474 42922 17034
rect 78 11002 1638 12562
rect 41362 11002 42922 12562
rect 78 6530 1638 8090
rect 41362 6530 42922 8090
rect 6616 78 8176 1638
rect 10142 78 11702 1638
rect 13668 78 15228 1638
rect 17194 78 18754 1638
rect 20720 78 22280 1638
rect 24246 78 25806 1638
rect 27772 78 29332 1638
rect 31298 78 32858 1638
rect 34824 78 36384 1638
use corns_clamp_mt CORNER_3
timestamp 1300118495
transform 0 1 0 -1 0 45924
box 0 0 6450 6450
use fillpp_mt fillpp_mt_563
timestamp 1300117811
transform 0 -1 6536 1 0 39474
box 0 0 6450 86
use ibacx6c3_mt nWait
timestamp 1300117536
transform 0 -1 8256 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_562
timestamp 1300117811
transform 0 -1 8342 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_561
timestamp 1300117811
transform 0 -1 8428 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_560
timestamp 1300117811
transform 0 -1 8514 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_559
timestamp 1300117811
transform 0 -1 8600 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_558
timestamp 1300117811
transform 0 -1 8686 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_557
timestamp 1300117811
transform 0 -1 8772 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_556
timestamp 1300117811
transform 0 -1 8858 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_555
timestamp 1300117811
transform 0 -1 8944 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_554
timestamp 1300117811
transform 0 -1 9030 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_553
timestamp 1300117811
transform 0 -1 9116 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_552
timestamp 1300117811
transform 0 -1 9202 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_551
timestamp 1300117811
transform 0 -1 9288 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_550
timestamp 1300117811
transform 0 -1 9374 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_549
timestamp 1300117811
transform 0 -1 9460 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_548
timestamp 1300117811
transform 0 -1 9546 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_547
timestamp 1300117811
transform 0 -1 9632 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_546
timestamp 1300117811
transform 0 -1 9718 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_545
timestamp 1300117811
transform 0 -1 9804 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_544
timestamp 1300117811
transform 0 -1 9890 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_543
timestamp 1300117811
transform 0 -1 9976 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_542
timestamp 1300117811
transform 0 -1 10062 1 0 39474
box 0 0 6450 86
use obaxxcsxe04_mt nME
timestamp 1300117393
transform 0 -1 11782 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_541
timestamp 1300117811
transform 0 -1 11868 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_540
timestamp 1300117811
transform 0 -1 11954 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_539
timestamp 1300117811
transform 0 -1 12040 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_538
timestamp 1300117811
transform 0 -1 12126 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_537
timestamp 1300117811
transform 0 -1 12212 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_536
timestamp 1300117811
transform 0 -1 12298 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_535
timestamp 1300117811
transform 0 -1 12384 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_534
timestamp 1300117811
transform 0 -1 12470 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_533
timestamp 1300117811
transform 0 -1 12556 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_532
timestamp 1300117811
transform 0 -1 12642 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_531
timestamp 1300117811
transform 0 -1 12728 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_530
timestamp 1300117811
transform 0 -1 12814 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_529
timestamp 1300117811
transform 0 -1 12900 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_528
timestamp 1300117811
transform 0 -1 12986 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_527
timestamp 1300117811
transform 0 -1 13072 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_526
timestamp 1300117811
transform 0 -1 13158 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_525
timestamp 1300117811
transform 0 -1 13244 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_524
timestamp 1300117811
transform 0 -1 13330 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_523
timestamp 1300117811
transform 0 -1 13416 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_522
timestamp 1300117811
transform 0 -1 13502 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_521
timestamp 1300117811
transform 0 -1 13588 1 0 39474
box 0 0 6450 86
use obaxxcsxe04_mt ALE
timestamp 1300117393
transform 0 -1 15308 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_520
timestamp 1300117811
transform 0 -1 15394 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_519
timestamp 1300117811
transform 0 -1 15480 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_518
timestamp 1300117811
transform 0 -1 15566 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_517
timestamp 1300117811
transform 0 -1 15652 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_516
timestamp 1300117811
transform 0 -1 15738 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_515
timestamp 1300117811
transform 0 -1 15824 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_514
timestamp 1300117811
transform 0 -1 15910 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_513
timestamp 1300117811
transform 0 -1 15996 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_512
timestamp 1300117811
transform 0 -1 16082 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_511
timestamp 1300117811
transform 0 -1 16168 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_510
timestamp 1300117811
transform 0 -1 16254 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_509
timestamp 1300117811
transform 0 -1 16340 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_508
timestamp 1300117811
transform 0 -1 16426 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_507
timestamp 1300117811
transform 0 -1 16512 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_506
timestamp 1300117811
transform 0 -1 16598 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_505
timestamp 1300117811
transform 0 -1 16684 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_504
timestamp 1300117811
transform 0 -1 16770 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_503
timestamp 1300117811
transform 0 -1 16856 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_502
timestamp 1300117811
transform 0 -1 16942 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_501
timestamp 1300117811
transform 0 -1 17028 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_500
timestamp 1300117811
transform 0 -1 17114 1 0 39474
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_15
timestamp 1300115302
transform 0 -1 18834 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_499
timestamp 1300117811
transform 0 -1 18920 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_498
timestamp 1300117811
transform 0 -1 19006 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_497
timestamp 1300117811
transform 0 -1 19092 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_496
timestamp 1300117811
transform 0 -1 19178 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_495
timestamp 1300117811
transform 0 -1 19264 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_494
timestamp 1300117811
transform 0 -1 19350 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_493
timestamp 1300117811
transform 0 -1 19436 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_492
timestamp 1300117811
transform 0 -1 19522 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_491
timestamp 1300117811
transform 0 -1 19608 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_490
timestamp 1300117811
transform 0 -1 19694 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_489
timestamp 1300117811
transform 0 -1 19780 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_488
timestamp 1300117811
transform 0 -1 19866 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_487
timestamp 1300117811
transform 0 -1 19952 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_486
timestamp 1300117811
transform 0 -1 20038 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_485
timestamp 1300117811
transform 0 -1 20124 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_484
timestamp 1300117811
transform 0 -1 20210 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_483
timestamp 1300117811
transform 0 -1 20296 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_482
timestamp 1300117811
transform 0 -1 20382 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_481
timestamp 1300117811
transform 0 -1 20468 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_480
timestamp 1300117811
transform 0 -1 20554 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_479
timestamp 1300117811
transform 0 -1 20640 1 0 39474
box 0 0 6450 86
use zgppxpg_mt VSSpads_0
timestamp 1300122446
transform 0 -1 22360 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_478
timestamp 1300117811
transform 0 -1 22446 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_477
timestamp 1300117811
transform 0 -1 22532 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_476
timestamp 1300117811
transform 0 -1 22618 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_475
timestamp 1300117811
transform 0 -1 22704 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_474
timestamp 1300117811
transform 0 -1 22790 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_473
timestamp 1300117811
transform 0 -1 22876 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_472
timestamp 1300117811
transform 0 -1 22962 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_471
timestamp 1300117811
transform 0 -1 23048 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_470
timestamp 1300117811
transform 0 -1 23134 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_469
timestamp 1300117811
transform 0 -1 23220 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_468
timestamp 1300117811
transform 0 -1 23306 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_467
timestamp 1300117811
transform 0 -1 23392 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_466
timestamp 1300117811
transform 0 -1 23478 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_465
timestamp 1300117811
transform 0 -1 23564 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_464
timestamp 1300117811
transform 0 -1 23650 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_463
timestamp 1300117811
transform 0 -1 23736 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_462
timestamp 1300117811
transform 0 -1 23822 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_461
timestamp 1300117811
transform 0 -1 23908 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_460
timestamp 1300117811
transform 0 -1 23994 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_459
timestamp 1300117811
transform 0 -1 24080 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_458
timestamp 1300117811
transform 0 -1 24166 1 0 39474
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_14
timestamp 1300115302
transform 0 -1 25886 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_457
timestamp 1300117811
transform 0 -1 25972 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_456
timestamp 1300117811
transform 0 -1 26058 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_455
timestamp 1300117811
transform 0 -1 26144 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_454
timestamp 1300117811
transform 0 -1 26230 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_453
timestamp 1300117811
transform 0 -1 26316 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_452
timestamp 1300117811
transform 0 -1 26402 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_451
timestamp 1300117811
transform 0 -1 26488 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_450
timestamp 1300117811
transform 0 -1 26574 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_449
timestamp 1300117811
transform 0 -1 26660 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_448
timestamp 1300117811
transform 0 -1 26746 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_447
timestamp 1300117811
transform 0 -1 26832 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_446
timestamp 1300117811
transform 0 -1 26918 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_445
timestamp 1300117811
transform 0 -1 27004 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_444
timestamp 1300117811
transform 0 -1 27090 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_443
timestamp 1300117811
transform 0 -1 27176 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_442
timestamp 1300117811
transform 0 -1 27262 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_441
timestamp 1300117811
transform 0 -1 27348 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_440
timestamp 1300117811
transform 0 -1 27434 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_439
timestamp 1300117811
transform 0 -1 27520 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_438
timestamp 1300117811
transform 0 -1 27606 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_437
timestamp 1300117811
transform 0 -1 27692 1 0 39474
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_13
timestamp 1300115302
transform 0 -1 29412 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_436
timestamp 1300117811
transform 0 -1 29498 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_435
timestamp 1300117811
transform 0 -1 29584 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_434
timestamp 1300117811
transform 0 -1 29670 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_433
timestamp 1300117811
transform 0 -1 29756 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_432
timestamp 1300117811
transform 0 -1 29842 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_431
timestamp 1300117811
transform 0 -1 29928 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_430
timestamp 1300117811
transform 0 -1 30014 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_429
timestamp 1300117811
transform 0 -1 30100 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_428
timestamp 1300117811
transform 0 -1 30186 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_427
timestamp 1300117811
transform 0 -1 30272 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_426
timestamp 1300117811
transform 0 -1 30358 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_425
timestamp 1300117811
transform 0 -1 30444 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_424
timestamp 1300117811
transform 0 -1 30530 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_423
timestamp 1300117811
transform 0 -1 30616 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_422
timestamp 1300117811
transform 0 -1 30702 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_421
timestamp 1300117811
transform 0 -1 30788 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_420
timestamp 1300117811
transform 0 -1 30874 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_419
timestamp 1300117811
transform 0 -1 30960 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_418
timestamp 1300117811
transform 0 -1 31046 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_417
timestamp 1300117811
transform 0 -1 31132 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_416
timestamp 1300117811
transform 0 -1 31218 1 0 39474
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_12
timestamp 1300115302
transform 0 -1 32938 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_415
timestamp 1300117811
transform 0 -1 33024 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_414
timestamp 1300117811
transform 0 -1 33110 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_413
timestamp 1300117811
transform 0 -1 33196 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_412
timestamp 1300117811
transform 0 -1 33282 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_411
timestamp 1300117811
transform 0 -1 33368 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_410
timestamp 1300117811
transform 0 -1 33454 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_409
timestamp 1300117811
transform 0 -1 33540 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_408
timestamp 1300117811
transform 0 -1 33626 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_407
timestamp 1300117811
transform 0 -1 33712 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_406
timestamp 1300117811
transform 0 -1 33798 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_405
timestamp 1300117811
transform 0 -1 33884 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_404
timestamp 1300117811
transform 0 -1 33970 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_403
timestamp 1300117811
transform 0 -1 34056 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_402
timestamp 1300117811
transform 0 -1 34142 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_401
timestamp 1300117811
transform 0 -1 34228 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_400
timestamp 1300117811
transform 0 -1 34314 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_399
timestamp 1300117811
transform 0 -1 34400 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_398
timestamp 1300117811
transform 0 -1 34486 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_397
timestamp 1300117811
transform 0 -1 34572 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_396
timestamp 1300117811
transform 0 -1 34658 1 0 39474
box 0 0 6450 86
use fillpp_mt fillpp_mt_395
timestamp 1300117811
transform 0 -1 34744 1 0 39474
box 0 0 6450 86
use zgppxpp_mt VDDPads_1
timestamp 1300121810
transform 0 -1 36464 1 0 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_394
timestamp 1300117811
transform 0 -1 36550 1 0 39474
box 0 0 6450 86
use corns_clamp_mt CORNER_2
timestamp 1300118495
transform -1 0 43000 0 -1 45924
box 0 0 6450 6450
use obaxxcsxe04_mt nOE
timestamp 1300117393
transform -1 0 6450 0 -1 39474
box 0 0 6450 1720
use fillpp_mt fillpp_mt_564
timestamp 1300117811
transform -1 0 6450 0 -1 37754
box 0 0 6450 86
use fillpp_mt fillpp_mt_565
timestamp 1300117811
transform -1 0 6450 0 -1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_566
timestamp 1300117811
transform -1 0 6450 0 -1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_567
timestamp 1300117811
transform -1 0 6450 0 -1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_568
timestamp 1300117811
transform -1 0 6450 0 -1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_569
timestamp 1300117811
transform -1 0 6450 0 -1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_570
timestamp 1300117811
transform -1 0 6450 0 -1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_571
timestamp 1300117811
transform -1 0 6450 0 -1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_572
timestamp 1300117811
transform -1 0 6450 0 -1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_573
timestamp 1300117811
transform -1 0 6450 0 -1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_574
timestamp 1300117811
transform -1 0 6450 0 -1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_575
timestamp 1300117811
transform -1 0 6450 0 -1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_576
timestamp 1300117811
transform -1 0 6450 0 -1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_577
timestamp 1300117811
transform -1 0 6450 0 -1 36636
box 0 0 6450 86
use fillpp_mt fillpp_mt_578
timestamp 1300117811
transform -1 0 6450 0 -1 36550
box 0 0 6450 86
use fillpp_mt fillpp_mt_579
timestamp 1300117811
transform -1 0 6450 0 -1 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_580
timestamp 1300117811
transform -1 0 6450 0 -1 36378
box 0 0 6450 86
use fillpp_mt fillpp_mt_581
timestamp 1300117811
transform -1 0 6450 0 -1 36292
box 0 0 6450 86
use fillpp_mt fillpp_mt_582
timestamp 1300117811
transform -1 0 6450 0 -1 36206
box 0 0 6450 86
use fillpp_mt fillpp_mt_583
timestamp 1300117811
transform -1 0 6450 0 -1 36120
box 0 0 6450 86
use fillpp_mt fillpp_mt_584
timestamp 1300117811
transform -1 0 6450 0 -1 36034
box 0 0 6450 86
use fillpp_mt fillpp_mt_585
timestamp 1300117811
transform -1 0 6450 0 -1 35948
box 0 0 6450 86
use fillpp_mt fillpp_mt_586
timestamp 1300117811
transform -1 0 6450 0 -1 35862
box 0 0 6450 86
use fillpp_mt fillpp_mt_587
timestamp 1300117811
transform -1 0 6450 0 -1 35776
box 0 0 6450 86
use fillpp_mt fillpp_mt_588
timestamp 1300117811
transform -1 0 6450 0 -1 35690
box 0 0 6450 86
use fillpp_mt fillpp_mt_589
timestamp 1300117811
transform -1 0 6450 0 -1 35604
box 0 0 6450 86
use fillpp_mt fillpp_mt_590
timestamp 1300117811
transform -1 0 6450 0 -1 35518
box 0 0 6450 86
use fillpp_mt fillpp_mt_591
timestamp 1300117811
transform -1 0 6450 0 -1 35432
box 0 0 6450 86
use fillpp_mt fillpp_mt_592
timestamp 1300117811
transform -1 0 6450 0 -1 35346
box 0 0 6450 86
use fillpp_mt fillpp_mt_593
timestamp 1300117811
transform -1 0 6450 0 -1 35260
box 0 0 6450 86
use fillpp_mt fillpp_mt_594
timestamp 1300117811
transform -1 0 6450 0 -1 35174
box 0 0 6450 86
use fillpp_mt fillpp_mt_595
timestamp 1300117811
transform -1 0 6450 0 -1 35088
box 0 0 6450 86
use obaxxcsxe04_mt RnW
timestamp 1300117393
transform -1 0 6450 0 -1 35002
box 0 0 6450 1720
use fillpp_mt fillpp_mt_596
timestamp 1300117811
transform -1 0 6450 0 -1 33282
box 0 0 6450 86
use fillpp_mt fillpp_mt_597
timestamp 1300117811
transform -1 0 6450 0 -1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_598
timestamp 1300117811
transform -1 0 6450 0 -1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_599
timestamp 1300117811
transform -1 0 6450 0 -1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_600
timestamp 1300117811
transform -1 0 6450 0 -1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_601
timestamp 1300117811
transform -1 0 6450 0 -1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_602
timestamp 1300117811
transform -1 0 6450 0 -1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_603
timestamp 1300117811
transform -1 0 6450 0 -1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_604
timestamp 1300117811
transform -1 0 6450 0 -1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_605
timestamp 1300117811
transform -1 0 6450 0 -1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_606
timestamp 1300117811
transform -1 0 6450 0 -1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_607
timestamp 1300117811
transform -1 0 6450 0 -1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_608
timestamp 1300117811
transform -1 0 6450 0 -1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_609
timestamp 1300117811
transform -1 0 6450 0 -1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_610
timestamp 1300117811
transform -1 0 6450 0 -1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_611
timestamp 1300117811
transform -1 0 6450 0 -1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_612
timestamp 1300117811
transform -1 0 6450 0 -1 31906
box 0 0 6450 86
use fillpp_mt fillpp_mt_613
timestamp 1300117811
transform -1 0 6450 0 -1 31820
box 0 0 6450 86
use fillpp_mt fillpp_mt_614
timestamp 1300117811
transform -1 0 6450 0 -1 31734
box 0 0 6450 86
use fillpp_mt fillpp_mt_615
timestamp 1300117811
transform -1 0 6450 0 -1 31648
box 0 0 6450 86
use fillpp_mt fillpp_mt_616
timestamp 1300117811
transform -1 0 6450 0 -1 31562
box 0 0 6450 86
use fillpp_mt fillpp_mt_617
timestamp 1300117811
transform -1 0 6450 0 -1 31476
box 0 0 6450 86
use fillpp_mt fillpp_mt_618
timestamp 1300117811
transform -1 0 6450 0 -1 31390
box 0 0 6450 86
use fillpp_mt fillpp_mt_619
timestamp 1300117811
transform -1 0 6450 0 -1 31304
box 0 0 6450 86
use fillpp_mt fillpp_mt_620
timestamp 1300117811
transform -1 0 6450 0 -1 31218
box 0 0 6450 86
use fillpp_mt fillpp_mt_621
timestamp 1300117811
transform -1 0 6450 0 -1 31132
box 0 0 6450 86
use fillpp_mt fillpp_mt_622
timestamp 1300117811
transform -1 0 6450 0 -1 31046
box 0 0 6450 86
use fillpp_mt fillpp_mt_623
timestamp 1300117811
transform -1 0 6450 0 -1 30960
box 0 0 6450 86
use fillpp_mt fillpp_mt_624
timestamp 1300117811
transform -1 0 6450 0 -1 30874
box 0 0 6450 86
use fillpp_mt fillpp_mt_625
timestamp 1300117811
transform -1 0 6450 0 -1 30788
box 0 0 6450 86
use fillpp_mt fillpp_mt_626
timestamp 1300117811
transform -1 0 6450 0 -1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_627
timestamp 1300117811
transform -1 0 6450 0 -1 30616
box 0 0 6450 86
use obaxxcsxe04_mt SDO
timestamp 1300117393
transform -1 0 6450 0 -1 30530
box 0 0 6450 1720
use fillpp_mt fillpp_mt_628
timestamp 1300117811
transform -1 0 6450 0 -1 28810
box 0 0 6450 86
use fillpp_mt fillpp_mt_629
timestamp 1300117811
transform -1 0 6450 0 -1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_630
timestamp 1300117811
transform -1 0 6450 0 -1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_631
timestamp 1300117811
transform -1 0 6450 0 -1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_632
timestamp 1300117811
transform -1 0 6450 0 -1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_633
timestamp 1300117811
transform -1 0 6450 0 -1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_634
timestamp 1300117811
transform -1 0 6450 0 -1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_635
timestamp 1300117811
transform -1 0 6450 0 -1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_636
timestamp 1300117811
transform -1 0 6450 0 -1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_637
timestamp 1300117811
transform -1 0 6450 0 -1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_638
timestamp 1300117811
transform -1 0 6450 0 -1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_639
timestamp 1300117811
transform -1 0 6450 0 -1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_640
timestamp 1300117811
transform -1 0 6450 0 -1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_641
timestamp 1300117811
transform -1 0 6450 0 -1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_642
timestamp 1300117811
transform -1 0 6450 0 -1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_643
timestamp 1300117811
transform -1 0 6450 0 -1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_644
timestamp 1300117811
transform -1 0 6450 0 -1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_645
timestamp 1300117811
transform -1 0 6450 0 -1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_646
timestamp 1300117811
transform -1 0 6450 0 -1 27262
box 0 0 6450 86
use fillpp_mt fillpp_mt_647
timestamp 1300117811
transform -1 0 6450 0 -1 27176
box 0 0 6450 86
use fillpp_mt fillpp_mt_648
timestamp 1300117811
transform -1 0 6450 0 -1 27090
box 0 0 6450 86
use fillpp_mt fillpp_mt_649
timestamp 1300117811
transform -1 0 6450 0 -1 27004
box 0 0 6450 86
use fillpp_mt fillpp_mt_650
timestamp 1300117811
transform -1 0 6450 0 -1 26918
box 0 0 6450 86
use fillpp_mt fillpp_mt_651
timestamp 1300117811
transform -1 0 6450 0 -1 26832
box 0 0 6450 86
use fillpp_mt fillpp_mt_652
timestamp 1300117811
transform -1 0 6450 0 -1 26746
box 0 0 6450 86
use fillpp_mt fillpp_mt_653
timestamp 1300117811
transform -1 0 6450 0 -1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_654
timestamp 1300117811
transform -1 0 6450 0 -1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_655
timestamp 1300117811
transform -1 0 6450 0 -1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_656
timestamp 1300117811
transform -1 0 6450 0 -1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_657
timestamp 1300117811
transform -1 0 6450 0 -1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_658
timestamp 1300117811
transform -1 0 6450 0 -1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_659
timestamp 1300117811
transform -1 0 6450 0 -1 26144
box 0 0 6450 86
use zgppxcp_mt VDDcore
timestamp 1300120773
transform -1 0 6450 0 -1 26058
box 0 0 6450 1720
use fillpp_mt fillpp_mt_660
timestamp 1300117811
transform -1 0 6450 0 -1 24338
box 0 0 6450 86
use fillpp_mt fillpp_mt_661
timestamp 1300117811
transform -1 0 6450 0 -1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_662
timestamp 1300117811
transform -1 0 6450 0 -1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_663
timestamp 1300117811
transform -1 0 6450 0 -1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_664
timestamp 1300117811
transform -1 0 6450 0 -1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_665
timestamp 1300117811
transform -1 0 6450 0 -1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_666
timestamp 1300117811
transform -1 0 6450 0 -1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_667
timestamp 1300117811
transform -1 0 6450 0 -1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_668
timestamp 1300117811
transform -1 0 6450 0 -1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_669
timestamp 1300117811
transform -1 0 6450 0 -1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_670
timestamp 1300117811
transform -1 0 6450 0 -1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_671
timestamp 1300117811
transform -1 0 6450 0 -1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_672
timestamp 1300117811
transform -1 0 6450 0 -1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_673
timestamp 1300117811
transform -1 0 6450 0 -1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_674
timestamp 1300117811
transform -1 0 6450 0 -1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_675
timestamp 1300117811
transform -1 0 6450 0 -1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_676
timestamp 1300117811
transform -1 0 6450 0 -1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_677
timestamp 1300117811
transform -1 0 6450 0 -1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_678
timestamp 1300117811
transform -1 0 6450 0 -1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_679
timestamp 1300117811
transform -1 0 6450 0 -1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_680
timestamp 1300117811
transform -1 0 6450 0 -1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_681
timestamp 1300117811
transform -1 0 6450 0 -1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_682
timestamp 1300117811
transform -1 0 6450 0 -1 22446
box 0 0 6450 86
use fillpp_mt fillpp_mt_683
timestamp 1300117811
transform -1 0 6450 0 -1 22360
box 0 0 6450 86
use fillpp_mt fillpp_mt_684
timestamp 1300117811
transform -1 0 6450 0 -1 22274
box 0 0 6450 86
use fillpp_mt fillpp_mt_685
timestamp 1300117811
transform -1 0 6450 0 -1 22188
box 0 0 6450 86
use fillpp_mt fillpp_mt_686
timestamp 1300117811
transform -1 0 6450 0 -1 22102
box 0 0 6450 86
use fillpp_mt fillpp_mt_687
timestamp 1300117811
transform -1 0 6450 0 -1 22016
box 0 0 6450 86
use fillpp_mt fillpp_mt_688
timestamp 1300117811
transform -1 0 6450 0 -1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_689
timestamp 1300117811
transform -1 0 6450 0 -1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_690
timestamp 1300117811
transform -1 0 6450 0 -1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_691
timestamp 1300117811
transform -1 0 6450 0 -1 21672
box 0 0 6450 86
use ibacx6xx_mt SDI
timestamp 1300117536
transform -1 0 6450 0 -1 21586
box 0 0 6450 1720
use fillpp_mt fillpp_mt_692
timestamp 1300117811
transform -1 0 6450 0 -1 19866
box 0 0 6450 86
use fillpp_mt fillpp_mt_693
timestamp 1300117811
transform -1 0 6450 0 -1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_694
timestamp 1300117811
transform -1 0 6450 0 -1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_695
timestamp 1300117811
transform -1 0 6450 0 -1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_696
timestamp 1300117811
transform -1 0 6450 0 -1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_697
timestamp 1300117811
transform -1 0 6450 0 -1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_698
timestamp 1300117811
transform -1 0 6450 0 -1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_699
timestamp 1300117811
transform -1 0 6450 0 -1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_700
timestamp 1300117811
transform -1 0 6450 0 -1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_701
timestamp 1300117811
transform -1 0 6450 0 -1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_702
timestamp 1300117811
transform -1 0 6450 0 -1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_703
timestamp 1300117811
transform -1 0 6450 0 -1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_704
timestamp 1300117811
transform -1 0 6450 0 -1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_705
timestamp 1300117811
transform -1 0 6450 0 -1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_706
timestamp 1300117811
transform -1 0 6450 0 -1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_707
timestamp 1300117811
transform -1 0 6450 0 -1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_708
timestamp 1300117811
transform -1 0 6450 0 -1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_709
timestamp 1300117811
transform -1 0 6450 0 -1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_710
timestamp 1300117811
transform -1 0 6450 0 -1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_711
timestamp 1300117811
transform -1 0 6450 0 -1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_712
timestamp 1300117811
transform -1 0 6450 0 -1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_713
timestamp 1300117811
transform -1 0 6450 0 -1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_714
timestamp 1300117811
transform -1 0 6450 0 -1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_715
timestamp 1300117811
transform -1 0 6450 0 -1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_716
timestamp 1300117811
transform -1 0 6450 0 -1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_717
timestamp 1300117811
transform -1 0 6450 0 -1 17716
box 0 0 6450 86
use fillpp_mt fillpp_mt_718
timestamp 1300117811
transform -1 0 6450 0 -1 17630
box 0 0 6450 86
use fillpp_mt fillpp_mt_719
timestamp 1300117811
transform -1 0 6450 0 -1 17544
box 0 0 6450 86
use fillpp_mt fillpp_mt_720
timestamp 1300117811
transform -1 0 6450 0 -1 17458
box 0 0 6450 86
use fillpp_mt fillpp_mt_721
timestamp 1300117811
transform -1 0 6450 0 -1 17372
box 0 0 6450 86
use fillpp_mt fillpp_mt_722
timestamp 1300117811
transform -1 0 6450 0 -1 17286
box 0 0 6450 86
use fillpp_mt fillpp_mt_723
timestamp 1300117811
transform -1 0 6450 0 -1 17200
box 0 0 6450 86
use ibacx6xx_mt Test
timestamp 1300117536
transform -1 0 6450 0 -1 17114
box 0 0 6450 1720
use fillpp_mt fillpp_mt_724
timestamp 1300117811
transform -1 0 6450 0 -1 15394
box 0 0 6450 86
use fillpp_mt fillpp_mt_725
timestamp 1300117811
transform -1 0 6450 0 -1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_726
timestamp 1300117811
transform -1 0 6450 0 -1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_727
timestamp 1300117811
transform -1 0 6450 0 -1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_728
timestamp 1300117811
transform -1 0 6450 0 -1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_729
timestamp 1300117811
transform -1 0 6450 0 -1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_730
timestamp 1300117811
transform -1 0 6450 0 -1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_731
timestamp 1300117811
transform -1 0 6450 0 -1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_732
timestamp 1300117811
transform -1 0 6450 0 -1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_733
timestamp 1300117811
transform -1 0 6450 0 -1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_734
timestamp 1300117811
transform -1 0 6450 0 -1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_735
timestamp 1300117811
transform -1 0 6450 0 -1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_736
timestamp 1300117811
transform -1 0 6450 0 -1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_737
timestamp 1300117811
transform -1 0 6450 0 -1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_738
timestamp 1300117811
transform -1 0 6450 0 -1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_739
timestamp 1300117811
transform -1 0 6450 0 -1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_740
timestamp 1300117811
transform -1 0 6450 0 -1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_741
timestamp 1300117811
transform -1 0 6450 0 -1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_742
timestamp 1300117811
transform -1 0 6450 0 -1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_743
timestamp 1300117811
transform -1 0 6450 0 -1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_744
timestamp 1300117811
transform -1 0 6450 0 -1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_745
timestamp 1300117811
transform -1 0 6450 0 -1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_746
timestamp 1300117811
transform -1 0 6450 0 -1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_747
timestamp 1300117811
transform -1 0 6450 0 -1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_748
timestamp 1300117811
transform -1 0 6450 0 -1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_749
timestamp 1300117811
transform -1 0 6450 0 -1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_750
timestamp 1300117811
transform -1 0 6450 0 -1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_751
timestamp 1300117811
transform -1 0 6450 0 -1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_752
timestamp 1300117811
transform -1 0 6450 0 -1 12986
box 0 0 6450 86
use fillpp_mt fillpp_mt_753
timestamp 1300117811
transform -1 0 6450 0 -1 12900
box 0 0 6450 86
use fillpp_mt fillpp_mt_754
timestamp 1300117811
transform -1 0 6450 0 -1 12814
box 0 0 6450 86
use fillpp_mt fillpp_mt_755
timestamp 1300117811
transform -1 0 6450 0 -1 12728
box 0 0 6450 86
use ibacx6xx_mt Clock
timestamp 1300117536
transform -1 0 6450 0 -1 12642
box 0 0 6450 1720
use fillpp_mt fillpp_mt_756
timestamp 1300117811
transform -1 0 6450 0 -1 10922
box 0 0 6450 86
use fillpp_mt fillpp_mt_757
timestamp 1300117811
transform -1 0 6450 0 -1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_758
timestamp 1300117811
transform -1 0 6450 0 -1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_759
timestamp 1300117811
transform -1 0 6450 0 -1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_760
timestamp 1300117811
transform -1 0 6450 0 -1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_761
timestamp 1300117811
transform -1 0 6450 0 -1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_762
timestamp 1300117811
transform -1 0 6450 0 -1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_763
timestamp 1300117811
transform -1 0 6450 0 -1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_764
timestamp 1300117811
transform -1 0 6450 0 -1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_765
timestamp 1300117811
transform -1 0 6450 0 -1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_766
timestamp 1300117811
transform -1 0 6450 0 -1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_767
timestamp 1300117811
transform -1 0 6450 0 -1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_768
timestamp 1300117811
transform -1 0 6450 0 -1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_769
timestamp 1300117811
transform -1 0 6450 0 -1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_770
timestamp 1300117811
transform -1 0 6450 0 -1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_771
timestamp 1300117811
transform -1 0 6450 0 -1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_772
timestamp 1300117811
transform -1 0 6450 0 -1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_773
timestamp 1300117811
transform -1 0 6450 0 -1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_774
timestamp 1300117811
transform -1 0 6450 0 -1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_775
timestamp 1300117811
transform -1 0 6450 0 -1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_776
timestamp 1300117811
transform -1 0 6450 0 -1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_777
timestamp 1300117811
transform -1 0 6450 0 -1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_778
timestamp 1300117811
transform -1 0 6450 0 -1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_779
timestamp 1300117811
transform -1 0 6450 0 -1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_780
timestamp 1300117811
transform -1 0 6450 0 -1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_781
timestamp 1300117811
transform -1 0 6450 0 -1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_782
timestamp 1300117811
transform -1 0 6450 0 -1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_783
timestamp 1300117811
transform -1 0 6450 0 -1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_784
timestamp 1300117811
transform -1 0 6450 0 -1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_785
timestamp 1300117811
transform -1 0 6450 0 -1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_786
timestamp 1300117811
transform -1 0 6450 0 -1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_787
timestamp 1300117811
transform -1 0 6450 0 -1 8256
box 0 0 6450 86
use ibacx6xx_mt nReset
timestamp 1300117536
transform -1 0 6450 0 -1 8170
box 0 0 6450 1720
use ioacx6xxcsxe04_mt Data_11
timestamp 1300115302
transform 1 0 36550 0 1 37754
box 0 0 6450 1720
use fillpp_mt fillpp_mt_393
timestamp 1300117811
transform 1 0 36550 0 1 37668
box 0 0 6450 86
use fillpp_mt fillpp_mt_392
timestamp 1300117811
transform 1 0 36550 0 1 37582
box 0 0 6450 86
use fillpp_mt fillpp_mt_391
timestamp 1300117811
transform 1 0 36550 0 1 37496
box 0 0 6450 86
use fillpp_mt fillpp_mt_390
timestamp 1300117811
transform 1 0 36550 0 1 37410
box 0 0 6450 86
use fillpp_mt fillpp_mt_389
timestamp 1300117811
transform 1 0 36550 0 1 37324
box 0 0 6450 86
use fillpp_mt fillpp_mt_388
timestamp 1300117811
transform 1 0 36550 0 1 37238
box 0 0 6450 86
use fillpp_mt fillpp_mt_387
timestamp 1300117811
transform 1 0 36550 0 1 37152
box 0 0 6450 86
use fillpp_mt fillpp_mt_386
timestamp 1300117811
transform 1 0 36550 0 1 37066
box 0 0 6450 86
use fillpp_mt fillpp_mt_385
timestamp 1300117811
transform 1 0 36550 0 1 36980
box 0 0 6450 86
use fillpp_mt fillpp_mt_384
timestamp 1300117811
transform 1 0 36550 0 1 36894
box 0 0 6450 86
use fillpp_mt fillpp_mt_383
timestamp 1300117811
transform 1 0 36550 0 1 36808
box 0 0 6450 86
use fillpp_mt fillpp_mt_382
timestamp 1300117811
transform 1 0 36550 0 1 36722
box 0 0 6450 86
use fillpp_mt fillpp_mt_381
timestamp 1300117811
transform 1 0 36550 0 1 36636
box 0 0 6450 86
use fillpp_mt fillpp_mt_380
timestamp 1300117811
transform 1 0 36550 0 1 36550
box 0 0 6450 86
use fillpp_mt fillpp_mt_379
timestamp 1300117811
transform 1 0 36550 0 1 36464
box 0 0 6450 86
use fillpp_mt fillpp_mt_378
timestamp 1300117811
transform 1 0 36550 0 1 36378
box 0 0 6450 86
use fillpp_mt fillpp_mt_377
timestamp 1300117811
transform 1 0 36550 0 1 36292
box 0 0 6450 86
use fillpp_mt fillpp_mt_376
timestamp 1300117811
transform 1 0 36550 0 1 36206
box 0 0 6450 86
use fillpp_mt fillpp_mt_375
timestamp 1300117811
transform 1 0 36550 0 1 36120
box 0 0 6450 86
use fillpp_mt fillpp_mt_374
timestamp 1300117811
transform 1 0 36550 0 1 36034
box 0 0 6450 86
use fillpp_mt fillpp_mt_373
timestamp 1300117811
transform 1 0 36550 0 1 35948
box 0 0 6450 86
use fillpp_mt fillpp_mt_372
timestamp 1300117811
transform 1 0 36550 0 1 35862
box 0 0 6450 86
use fillpp_mt fillpp_mt_371
timestamp 1300117811
transform 1 0 36550 0 1 35776
box 0 0 6450 86
use fillpp_mt fillpp_mt_370
timestamp 1300117811
transform 1 0 36550 0 1 35690
box 0 0 6450 86
use fillpp_mt fillpp_mt_369
timestamp 1300117811
transform 1 0 36550 0 1 35604
box 0 0 6450 86
use fillpp_mt fillpp_mt_368
timestamp 1300117811
transform 1 0 36550 0 1 35518
box 0 0 6450 86
use fillpp_mt fillpp_mt_367
timestamp 1300117811
transform 1 0 36550 0 1 35432
box 0 0 6450 86
use fillpp_mt fillpp_mt_366
timestamp 1300117811
transform 1 0 36550 0 1 35346
box 0 0 6450 86
use fillpp_mt fillpp_mt_365
timestamp 1300117811
transform 1 0 36550 0 1 35260
box 0 0 6450 86
use fillpp_mt fillpp_mt_364
timestamp 1300117811
transform 1 0 36550 0 1 35174
box 0 0 6450 86
use fillpp_mt fillpp_mt_363
timestamp 1300117811
transform 1 0 36550 0 1 35088
box 0 0 6450 86
use fillpp_mt fillpp_mt_362
timestamp 1300117811
transform 1 0 36550 0 1 35002
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_10
timestamp 1300115302
transform 1 0 36550 0 1 33282
box 0 0 6450 1720
use fillpp_mt fillpp_mt_361
timestamp 1300117811
transform 1 0 36550 0 1 33196
box 0 0 6450 86
use fillpp_mt fillpp_mt_360
timestamp 1300117811
transform 1 0 36550 0 1 33110
box 0 0 6450 86
use fillpp_mt fillpp_mt_359
timestamp 1300117811
transform 1 0 36550 0 1 33024
box 0 0 6450 86
use fillpp_mt fillpp_mt_358
timestamp 1300117811
transform 1 0 36550 0 1 32938
box 0 0 6450 86
use fillpp_mt fillpp_mt_357
timestamp 1300117811
transform 1 0 36550 0 1 32852
box 0 0 6450 86
use fillpp_mt fillpp_mt_356
timestamp 1300117811
transform 1 0 36550 0 1 32766
box 0 0 6450 86
use fillpp_mt fillpp_mt_355
timestamp 1300117811
transform 1 0 36550 0 1 32680
box 0 0 6450 86
use fillpp_mt fillpp_mt_354
timestamp 1300117811
transform 1 0 36550 0 1 32594
box 0 0 6450 86
use fillpp_mt fillpp_mt_353
timestamp 1300117811
transform 1 0 36550 0 1 32508
box 0 0 6450 86
use fillpp_mt fillpp_mt_352
timestamp 1300117811
transform 1 0 36550 0 1 32422
box 0 0 6450 86
use fillpp_mt fillpp_mt_351
timestamp 1300117811
transform 1 0 36550 0 1 32336
box 0 0 6450 86
use fillpp_mt fillpp_mt_350
timestamp 1300117811
transform 1 0 36550 0 1 32250
box 0 0 6450 86
use fillpp_mt fillpp_mt_349
timestamp 1300117811
transform 1 0 36550 0 1 32164
box 0 0 6450 86
use fillpp_mt fillpp_mt_348
timestamp 1300117811
transform 1 0 36550 0 1 32078
box 0 0 6450 86
use fillpp_mt fillpp_mt_347
timestamp 1300117811
transform 1 0 36550 0 1 31992
box 0 0 6450 86
use fillpp_mt fillpp_mt_346
timestamp 1300117811
transform 1 0 36550 0 1 31906
box 0 0 6450 86
use fillpp_mt fillpp_mt_345
timestamp 1300117811
transform 1 0 36550 0 1 31820
box 0 0 6450 86
use fillpp_mt fillpp_mt_344
timestamp 1300117811
transform 1 0 36550 0 1 31734
box 0 0 6450 86
use fillpp_mt fillpp_mt_343
timestamp 1300117811
transform 1 0 36550 0 1 31648
box 0 0 6450 86
use fillpp_mt fillpp_mt_342
timestamp 1300117811
transform 1 0 36550 0 1 31562
box 0 0 6450 86
use fillpp_mt fillpp_mt_341
timestamp 1300117811
transform 1 0 36550 0 1 31476
box 0 0 6450 86
use fillpp_mt fillpp_mt_340
timestamp 1300117811
transform 1 0 36550 0 1 31390
box 0 0 6450 86
use fillpp_mt fillpp_mt_339
timestamp 1300117811
transform 1 0 36550 0 1 31304
box 0 0 6450 86
use fillpp_mt fillpp_mt_338
timestamp 1300117811
transform 1 0 36550 0 1 31218
box 0 0 6450 86
use fillpp_mt fillpp_mt_337
timestamp 1300117811
transform 1 0 36550 0 1 31132
box 0 0 6450 86
use fillpp_mt fillpp_mt_336
timestamp 1300117811
transform 1 0 36550 0 1 31046
box 0 0 6450 86
use fillpp_mt fillpp_mt_335
timestamp 1300117811
transform 1 0 36550 0 1 30960
box 0 0 6450 86
use fillpp_mt fillpp_mt_334
timestamp 1300117811
transform 1 0 36550 0 1 30874
box 0 0 6450 86
use fillpp_mt fillpp_mt_333
timestamp 1300117811
transform 1 0 36550 0 1 30788
box 0 0 6450 86
use fillpp_mt fillpp_mt_332
timestamp 1300117811
transform 1 0 36550 0 1 30702
box 0 0 6450 86
use fillpp_mt fillpp_mt_331
timestamp 1300117811
transform 1 0 36550 0 1 30616
box 0 0 6450 86
use fillpp_mt fillpp_mt_330
timestamp 1300117811
transform 1 0 36550 0 1 30530
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_9
timestamp 1300115302
transform 1 0 36550 0 1 28810
box 0 0 6450 1720
use fillpp_mt fillpp_mt_329
timestamp 1300117811
transform 1 0 36550 0 1 28724
box 0 0 6450 86
use fillpp_mt fillpp_mt_328
timestamp 1300117811
transform 1 0 36550 0 1 28638
box 0 0 6450 86
use fillpp_mt fillpp_mt_327
timestamp 1300117811
transform 1 0 36550 0 1 28552
box 0 0 6450 86
use fillpp_mt fillpp_mt_326
timestamp 1300117811
transform 1 0 36550 0 1 28466
box 0 0 6450 86
use fillpp_mt fillpp_mt_325
timestamp 1300117811
transform 1 0 36550 0 1 28380
box 0 0 6450 86
use fillpp_mt fillpp_mt_324
timestamp 1300117811
transform 1 0 36550 0 1 28294
box 0 0 6450 86
use fillpp_mt fillpp_mt_323
timestamp 1300117811
transform 1 0 36550 0 1 28208
box 0 0 6450 86
use fillpp_mt fillpp_mt_322
timestamp 1300117811
transform 1 0 36550 0 1 28122
box 0 0 6450 86
use fillpp_mt fillpp_mt_321
timestamp 1300117811
transform 1 0 36550 0 1 28036
box 0 0 6450 86
use fillpp_mt fillpp_mt_320
timestamp 1300117811
transform 1 0 36550 0 1 27950
box 0 0 6450 86
use fillpp_mt fillpp_mt_319
timestamp 1300117811
transform 1 0 36550 0 1 27864
box 0 0 6450 86
use fillpp_mt fillpp_mt_318
timestamp 1300117811
transform 1 0 36550 0 1 27778
box 0 0 6450 86
use fillpp_mt fillpp_mt_317
timestamp 1300117811
transform 1 0 36550 0 1 27692
box 0 0 6450 86
use fillpp_mt fillpp_mt_316
timestamp 1300117811
transform 1 0 36550 0 1 27606
box 0 0 6450 86
use fillpp_mt fillpp_mt_315
timestamp 1300117811
transform 1 0 36550 0 1 27520
box 0 0 6450 86
use fillpp_mt fillpp_mt_314
timestamp 1300117811
transform 1 0 36550 0 1 27434
box 0 0 6450 86
use fillpp_mt fillpp_mt_313
timestamp 1300117811
transform 1 0 36550 0 1 27348
box 0 0 6450 86
use fillpp_mt fillpp_mt_312
timestamp 1300117811
transform 1 0 36550 0 1 27262
box 0 0 6450 86
use fillpp_mt fillpp_mt_311
timestamp 1300117811
transform 1 0 36550 0 1 27176
box 0 0 6450 86
use fillpp_mt fillpp_mt_310
timestamp 1300117811
transform 1 0 36550 0 1 27090
box 0 0 6450 86
use fillpp_mt fillpp_mt_309
timestamp 1300117811
transform 1 0 36550 0 1 27004
box 0 0 6450 86
use fillpp_mt fillpp_mt_308
timestamp 1300117811
transform 1 0 36550 0 1 26918
box 0 0 6450 86
use fillpp_mt fillpp_mt_307
timestamp 1300117811
transform 1 0 36550 0 1 26832
box 0 0 6450 86
use fillpp_mt fillpp_mt_306
timestamp 1300117811
transform 1 0 36550 0 1 26746
box 0 0 6450 86
use fillpp_mt fillpp_mt_305
timestamp 1300117811
transform 1 0 36550 0 1 26660
box 0 0 6450 86
use fillpp_mt fillpp_mt_304
timestamp 1300117811
transform 1 0 36550 0 1 26574
box 0 0 6450 86
use fillpp_mt fillpp_mt_303
timestamp 1300117811
transform 1 0 36550 0 1 26488
box 0 0 6450 86
use fillpp_mt fillpp_mt_302
timestamp 1300117811
transform 1 0 36550 0 1 26402
box 0 0 6450 86
use fillpp_mt fillpp_mt_301
timestamp 1300117811
transform 1 0 36550 0 1 26316
box 0 0 6450 86
use fillpp_mt fillpp_mt_300
timestamp 1300117811
transform 1 0 36550 0 1 26230
box 0 0 6450 86
use fillpp_mt fillpp_mt_299
timestamp 1300117811
transform 1 0 36550 0 1 26144
box 0 0 6450 86
use fillpp_mt fillpp_mt_298
timestamp 1300117811
transform 1 0 36550 0 1 26058
box 0 0 6450 86
use zgppxcg_mt VSScore
timestamp 1300119877
transform 1 0 36550 0 1 24338
box 0 0 6450 1720
use fillpp_mt fillpp_mt_297
timestamp 1300117811
transform 1 0 36550 0 1 24252
box 0 0 6450 86
use fillpp_mt fillpp_mt_296
timestamp 1300117811
transform 1 0 36550 0 1 24166
box 0 0 6450 86
use fillpp_mt fillpp_mt_295
timestamp 1300117811
transform 1 0 36550 0 1 24080
box 0 0 6450 86
use fillpp_mt fillpp_mt_294
timestamp 1300117811
transform 1 0 36550 0 1 23994
box 0 0 6450 86
use fillpp_mt fillpp_mt_293
timestamp 1300117811
transform 1 0 36550 0 1 23908
box 0 0 6450 86
use fillpp_mt fillpp_mt_292
timestamp 1300117811
transform 1 0 36550 0 1 23822
box 0 0 6450 86
use fillpp_mt fillpp_mt_291
timestamp 1300117811
transform 1 0 36550 0 1 23736
box 0 0 6450 86
use fillpp_mt fillpp_mt_290
timestamp 1300117811
transform 1 0 36550 0 1 23650
box 0 0 6450 86
use fillpp_mt fillpp_mt_289
timestamp 1300117811
transform 1 0 36550 0 1 23564
box 0 0 6450 86
use fillpp_mt fillpp_mt_288
timestamp 1300117811
transform 1 0 36550 0 1 23478
box 0 0 6450 86
use fillpp_mt fillpp_mt_287
timestamp 1300117811
transform 1 0 36550 0 1 23392
box 0 0 6450 86
use fillpp_mt fillpp_mt_286
timestamp 1300117811
transform 1 0 36550 0 1 23306
box 0 0 6450 86
use fillpp_mt fillpp_mt_285
timestamp 1300117811
transform 1 0 36550 0 1 23220
box 0 0 6450 86
use fillpp_mt fillpp_mt_284
timestamp 1300117811
transform 1 0 36550 0 1 23134
box 0 0 6450 86
use fillpp_mt fillpp_mt_283
timestamp 1300117811
transform 1 0 36550 0 1 23048
box 0 0 6450 86
use fillpp_mt fillpp_mt_282
timestamp 1300117811
transform 1 0 36550 0 1 22962
box 0 0 6450 86
use fillpp_mt fillpp_mt_281
timestamp 1300117811
transform 1 0 36550 0 1 22876
box 0 0 6450 86
use fillpp_mt fillpp_mt_280
timestamp 1300117811
transform 1 0 36550 0 1 22790
box 0 0 6450 86
use fillpp_mt fillpp_mt_279
timestamp 1300117811
transform 1 0 36550 0 1 22704
box 0 0 6450 86
use fillpp_mt fillpp_mt_278
timestamp 1300117811
transform 1 0 36550 0 1 22618
box 0 0 6450 86
use fillpp_mt fillpp_mt_277
timestamp 1300117811
transform 1 0 36550 0 1 22532
box 0 0 6450 86
use fillpp_mt fillpp_mt_276
timestamp 1300117811
transform 1 0 36550 0 1 22446
box 0 0 6450 86
use fillpp_mt fillpp_mt_275
timestamp 1300117811
transform 1 0 36550 0 1 22360
box 0 0 6450 86
use fillpp_mt fillpp_mt_274
timestamp 1300117811
transform 1 0 36550 0 1 22274
box 0 0 6450 86
use fillpp_mt fillpp_mt_273
timestamp 1300117811
transform 1 0 36550 0 1 22188
box 0 0 6450 86
use fillpp_mt fillpp_mt_272
timestamp 1300117811
transform 1 0 36550 0 1 22102
box 0 0 6450 86
use fillpp_mt fillpp_mt_271
timestamp 1300117811
transform 1 0 36550 0 1 22016
box 0 0 6450 86
use fillpp_mt fillpp_mt_270
timestamp 1300117811
transform 1 0 36550 0 1 21930
box 0 0 6450 86
use fillpp_mt fillpp_mt_269
timestamp 1300117811
transform 1 0 36550 0 1 21844
box 0 0 6450 86
use fillpp_mt fillpp_mt_268
timestamp 1300117811
transform 1 0 36550 0 1 21758
box 0 0 6450 86
use fillpp_mt fillpp_mt_267
timestamp 1300117811
transform 1 0 36550 0 1 21672
box 0 0 6450 86
use fillpp_mt fillpp_mt_266
timestamp 1300117811
transform 1 0 36550 0 1 21586
box 0 0 6450 86
use zgppxpg_mt VSSEextra_0
timestamp 1300122446
transform 1 0 36550 0 1 19866
box 0 0 6450 1720
use fillpp_mt fillpp_mt_265
timestamp 1300117811
transform 1 0 36550 0 1 19780
box 0 0 6450 86
use fillpp_mt fillpp_mt_264
timestamp 1300117811
transform 1 0 36550 0 1 19694
box 0 0 6450 86
use fillpp_mt fillpp_mt_263
timestamp 1300117811
transform 1 0 36550 0 1 19608
box 0 0 6450 86
use fillpp_mt fillpp_mt_262
timestamp 1300117811
transform 1 0 36550 0 1 19522
box 0 0 6450 86
use fillpp_mt fillpp_mt_261
timestamp 1300117811
transform 1 0 36550 0 1 19436
box 0 0 6450 86
use fillpp_mt fillpp_mt_260
timestamp 1300117811
transform 1 0 36550 0 1 19350
box 0 0 6450 86
use fillpp_mt fillpp_mt_259
timestamp 1300117811
transform 1 0 36550 0 1 19264
box 0 0 6450 86
use fillpp_mt fillpp_mt_258
timestamp 1300117811
transform 1 0 36550 0 1 19178
box 0 0 6450 86
use fillpp_mt fillpp_mt_257
timestamp 1300117811
transform 1 0 36550 0 1 19092
box 0 0 6450 86
use fillpp_mt fillpp_mt_256
timestamp 1300117811
transform 1 0 36550 0 1 19006
box 0 0 6450 86
use fillpp_mt fillpp_mt_255
timestamp 1300117811
transform 1 0 36550 0 1 18920
box 0 0 6450 86
use fillpp_mt fillpp_mt_254
timestamp 1300117811
transform 1 0 36550 0 1 18834
box 0 0 6450 86
use fillpp_mt fillpp_mt_253
timestamp 1300117811
transform 1 0 36550 0 1 18748
box 0 0 6450 86
use fillpp_mt fillpp_mt_252
timestamp 1300117811
transform 1 0 36550 0 1 18662
box 0 0 6450 86
use fillpp_mt fillpp_mt_251
timestamp 1300117811
transform 1 0 36550 0 1 18576
box 0 0 6450 86
use fillpp_mt fillpp_mt_250
timestamp 1300117811
transform 1 0 36550 0 1 18490
box 0 0 6450 86
use fillpp_mt fillpp_mt_249
timestamp 1300117811
transform 1 0 36550 0 1 18404
box 0 0 6450 86
use fillpp_mt fillpp_mt_248
timestamp 1300117811
transform 1 0 36550 0 1 18318
box 0 0 6450 86
use fillpp_mt fillpp_mt_247
timestamp 1300117811
transform 1 0 36550 0 1 18232
box 0 0 6450 86
use fillpp_mt fillpp_mt_246
timestamp 1300117811
transform 1 0 36550 0 1 18146
box 0 0 6450 86
use fillpp_mt fillpp_mt_245
timestamp 1300117811
transform 1 0 36550 0 1 18060
box 0 0 6450 86
use fillpp_mt fillpp_mt_244
timestamp 1300117811
transform 1 0 36550 0 1 17974
box 0 0 6450 86
use fillpp_mt fillpp_mt_243
timestamp 1300117811
transform 1 0 36550 0 1 17888
box 0 0 6450 86
use fillpp_mt fillpp_mt_242
timestamp 1300117811
transform 1 0 36550 0 1 17802
box 0 0 6450 86
use fillpp_mt fillpp_mt_241
timestamp 1300117811
transform 1 0 36550 0 1 17716
box 0 0 6450 86
use fillpp_mt fillpp_mt_240
timestamp 1300117811
transform 1 0 36550 0 1 17630
box 0 0 6450 86
use fillpp_mt fillpp_mt_239
timestamp 1300117811
transform 1 0 36550 0 1 17544
box 0 0 6450 86
use fillpp_mt fillpp_mt_238
timestamp 1300117811
transform 1 0 36550 0 1 17458
box 0 0 6450 86
use fillpp_mt fillpp_mt_237
timestamp 1300117811
transform 1 0 36550 0 1 17372
box 0 0 6450 86
use fillpp_mt fillpp_mt_236
timestamp 1300117811
transform 1 0 36550 0 1 17286
box 0 0 6450 86
use fillpp_mt fillpp_mt_235
timestamp 1300117811
transform 1 0 36550 0 1 17200
box 0 0 6450 86
use fillpp_mt fillpp_mt_234
timestamp 1300117811
transform 1 0 36550 0 1 17114
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_8
timestamp 1300115302
transform 1 0 36550 0 1 15394
box 0 0 6450 1720
use fillpp_mt fillpp_mt_233
timestamp 1300117811
transform 1 0 36550 0 1 15308
box 0 0 6450 86
use fillpp_mt fillpp_mt_232
timestamp 1300117811
transform 1 0 36550 0 1 15222
box 0 0 6450 86
use fillpp_mt fillpp_mt_231
timestamp 1300117811
transform 1 0 36550 0 1 15136
box 0 0 6450 86
use fillpp_mt fillpp_mt_230
timestamp 1300117811
transform 1 0 36550 0 1 15050
box 0 0 6450 86
use fillpp_mt fillpp_mt_229
timestamp 1300117811
transform 1 0 36550 0 1 14964
box 0 0 6450 86
use fillpp_mt fillpp_mt_228
timestamp 1300117811
transform 1 0 36550 0 1 14878
box 0 0 6450 86
use fillpp_mt fillpp_mt_227
timestamp 1300117811
transform 1 0 36550 0 1 14792
box 0 0 6450 86
use fillpp_mt fillpp_mt_226
timestamp 1300117811
transform 1 0 36550 0 1 14706
box 0 0 6450 86
use fillpp_mt fillpp_mt_225
timestamp 1300117811
transform 1 0 36550 0 1 14620
box 0 0 6450 86
use fillpp_mt fillpp_mt_224
timestamp 1300117811
transform 1 0 36550 0 1 14534
box 0 0 6450 86
use fillpp_mt fillpp_mt_223
timestamp 1300117811
transform 1 0 36550 0 1 14448
box 0 0 6450 86
use fillpp_mt fillpp_mt_222
timestamp 1300117811
transform 1 0 36550 0 1 14362
box 0 0 6450 86
use fillpp_mt fillpp_mt_221
timestamp 1300117811
transform 1 0 36550 0 1 14276
box 0 0 6450 86
use fillpp_mt fillpp_mt_220
timestamp 1300117811
transform 1 0 36550 0 1 14190
box 0 0 6450 86
use fillpp_mt fillpp_mt_219
timestamp 1300117811
transform 1 0 36550 0 1 14104
box 0 0 6450 86
use fillpp_mt fillpp_mt_218
timestamp 1300117811
transform 1 0 36550 0 1 14018
box 0 0 6450 86
use fillpp_mt fillpp_mt_217
timestamp 1300117811
transform 1 0 36550 0 1 13932
box 0 0 6450 86
use fillpp_mt fillpp_mt_216
timestamp 1300117811
transform 1 0 36550 0 1 13846
box 0 0 6450 86
use fillpp_mt fillpp_mt_215
timestamp 1300117811
transform 1 0 36550 0 1 13760
box 0 0 6450 86
use fillpp_mt fillpp_mt_214
timestamp 1300117811
transform 1 0 36550 0 1 13674
box 0 0 6450 86
use fillpp_mt fillpp_mt_213
timestamp 1300117811
transform 1 0 36550 0 1 13588
box 0 0 6450 86
use fillpp_mt fillpp_mt_212
timestamp 1300117811
transform 1 0 36550 0 1 13502
box 0 0 6450 86
use fillpp_mt fillpp_mt_211
timestamp 1300117811
transform 1 0 36550 0 1 13416
box 0 0 6450 86
use fillpp_mt fillpp_mt_210
timestamp 1300117811
transform 1 0 36550 0 1 13330
box 0 0 6450 86
use fillpp_mt fillpp_mt_209
timestamp 1300117811
transform 1 0 36550 0 1 13244
box 0 0 6450 86
use fillpp_mt fillpp_mt_208
timestamp 1300117811
transform 1 0 36550 0 1 13158
box 0 0 6450 86
use fillpp_mt fillpp_mt_207
timestamp 1300117811
transform 1 0 36550 0 1 13072
box 0 0 6450 86
use fillpp_mt fillpp_mt_206
timestamp 1300117811
transform 1 0 36550 0 1 12986
box 0 0 6450 86
use fillpp_mt fillpp_mt_205
timestamp 1300117811
transform 1 0 36550 0 1 12900
box 0 0 6450 86
use fillpp_mt fillpp_mt_204
timestamp 1300117811
transform 1 0 36550 0 1 12814
box 0 0 6450 86
use fillpp_mt fillpp_mt_203
timestamp 1300117811
transform 1 0 36550 0 1 12728
box 0 0 6450 86
use fillpp_mt fillpp_mt_202
timestamp 1300117811
transform 1 0 36550 0 1 12642
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_7
timestamp 1300115302
transform 1 0 36550 0 1 10922
box 0 0 6450 1720
use fillpp_mt fillpp_mt_201
timestamp 1300117811
transform 1 0 36550 0 1 10836
box 0 0 6450 86
use fillpp_mt fillpp_mt_200
timestamp 1300117811
transform 1 0 36550 0 1 10750
box 0 0 6450 86
use fillpp_mt fillpp_mt_199
timestamp 1300117811
transform 1 0 36550 0 1 10664
box 0 0 6450 86
use fillpp_mt fillpp_mt_198
timestamp 1300117811
transform 1 0 36550 0 1 10578
box 0 0 6450 86
use fillpp_mt fillpp_mt_197
timestamp 1300117811
transform 1 0 36550 0 1 10492
box 0 0 6450 86
use fillpp_mt fillpp_mt_196
timestamp 1300117811
transform 1 0 36550 0 1 10406
box 0 0 6450 86
use fillpp_mt fillpp_mt_195
timestamp 1300117811
transform 1 0 36550 0 1 10320
box 0 0 6450 86
use fillpp_mt fillpp_mt_194
timestamp 1300117811
transform 1 0 36550 0 1 10234
box 0 0 6450 86
use fillpp_mt fillpp_mt_193
timestamp 1300117811
transform 1 0 36550 0 1 10148
box 0 0 6450 86
use fillpp_mt fillpp_mt_192
timestamp 1300117811
transform 1 0 36550 0 1 10062
box 0 0 6450 86
use fillpp_mt fillpp_mt_191
timestamp 1300117811
transform 1 0 36550 0 1 9976
box 0 0 6450 86
use fillpp_mt fillpp_mt_190
timestamp 1300117811
transform 1 0 36550 0 1 9890
box 0 0 6450 86
use fillpp_mt fillpp_mt_189
timestamp 1300117811
transform 1 0 36550 0 1 9804
box 0 0 6450 86
use fillpp_mt fillpp_mt_188
timestamp 1300117811
transform 1 0 36550 0 1 9718
box 0 0 6450 86
use fillpp_mt fillpp_mt_187
timestamp 1300117811
transform 1 0 36550 0 1 9632
box 0 0 6450 86
use fillpp_mt fillpp_mt_186
timestamp 1300117811
transform 1 0 36550 0 1 9546
box 0 0 6450 86
use fillpp_mt fillpp_mt_185
timestamp 1300117811
transform 1 0 36550 0 1 9460
box 0 0 6450 86
use fillpp_mt fillpp_mt_184
timestamp 1300117811
transform 1 0 36550 0 1 9374
box 0 0 6450 86
use fillpp_mt fillpp_mt_183
timestamp 1300117811
transform 1 0 36550 0 1 9288
box 0 0 6450 86
use fillpp_mt fillpp_mt_182
timestamp 1300117811
transform 1 0 36550 0 1 9202
box 0 0 6450 86
use fillpp_mt fillpp_mt_181
timestamp 1300117811
transform 1 0 36550 0 1 9116
box 0 0 6450 86
use fillpp_mt fillpp_mt_180
timestamp 1300117811
transform 1 0 36550 0 1 9030
box 0 0 6450 86
use fillpp_mt fillpp_mt_179
timestamp 1300117811
transform 1 0 36550 0 1 8944
box 0 0 6450 86
use fillpp_mt fillpp_mt_178
timestamp 1300117811
transform 1 0 36550 0 1 8858
box 0 0 6450 86
use fillpp_mt fillpp_mt_177
timestamp 1300117811
transform 1 0 36550 0 1 8772
box 0 0 6450 86
use fillpp_mt fillpp_mt_176
timestamp 1300117811
transform 1 0 36550 0 1 8686
box 0 0 6450 86
use fillpp_mt fillpp_mt_175
timestamp 1300117811
transform 1 0 36550 0 1 8600
box 0 0 6450 86
use fillpp_mt fillpp_mt_174
timestamp 1300117811
transform 1 0 36550 0 1 8514
box 0 0 6450 86
use fillpp_mt fillpp_mt_173
timestamp 1300117811
transform 1 0 36550 0 1 8428
box 0 0 6450 86
use fillpp_mt fillpp_mt_172
timestamp 1300117811
transform 1 0 36550 0 1 8342
box 0 0 6450 86
use fillpp_mt fillpp_mt_171
timestamp 1300117811
transform 1 0 36550 0 1 8256
box 0 0 6450 86
use fillpp_mt fillpp_mt_170
timestamp 1300117811
transform 1 0 36550 0 1 8170
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_6
timestamp 1300115302
transform 1 0 36550 0 1 6450
box 0 0 6450 1720
use corns_clamp_mt CORNER_0
timestamp 1300118495
transform 1 0 0 0 1 0
box 0 0 6450 6450
use fillpp_mt fillpp_mt_0
timestamp 1300117811
transform 0 1 6450 -1 0 6450
box 0 0 6450 86
use ibacx6c3_mt nIRQ
timestamp 1300117536
transform 0 1 6536 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_1
timestamp 1300117811
transform 0 1 8256 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_2
timestamp 1300117811
transform 0 1 8342 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_3
timestamp 1300117811
transform 0 1 8428 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_4
timestamp 1300117811
transform 0 1 8514 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_5
timestamp 1300117811
transform 0 1 8600 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_6
timestamp 1300117811
transform 0 1 8686 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_7
timestamp 1300117811
transform 0 1 8772 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_8
timestamp 1300117811
transform 0 1 8858 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_9
timestamp 1300117811
transform 0 1 8944 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_10
timestamp 1300117811
transform 0 1 9030 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_11
timestamp 1300117811
transform 0 1 9116 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_12
timestamp 1300117811
transform 0 1 9202 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_13
timestamp 1300117811
transform 0 1 9288 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_14
timestamp 1300117811
transform 0 1 9374 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_15
timestamp 1300117811
transform 0 1 9460 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_16
timestamp 1300117811
transform 0 1 9546 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_17
timestamp 1300117811
transform 0 1 9632 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_18
timestamp 1300117811
transform 0 1 9718 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_19
timestamp 1300117811
transform 0 1 9804 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_20
timestamp 1300117811
transform 0 1 9890 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_21
timestamp 1300117811
transform 0 1 9976 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_0
timestamp 1300115302
transform 0 1 10062 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_22
timestamp 1300117811
transform 0 1 11782 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_23
timestamp 1300117811
transform 0 1 11868 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_24
timestamp 1300117811
transform 0 1 11954 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_25
timestamp 1300117811
transform 0 1 12040 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_26
timestamp 1300117811
transform 0 1 12126 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_27
timestamp 1300117811
transform 0 1 12212 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_28
timestamp 1300117811
transform 0 1 12298 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_29
timestamp 1300117811
transform 0 1 12384 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_30
timestamp 1300117811
transform 0 1 12470 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_31
timestamp 1300117811
transform 0 1 12556 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_32
timestamp 1300117811
transform 0 1 12642 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_33
timestamp 1300117811
transform 0 1 12728 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_34
timestamp 1300117811
transform 0 1 12814 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_35
timestamp 1300117811
transform 0 1 12900 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_36
timestamp 1300117811
transform 0 1 12986 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_37
timestamp 1300117811
transform 0 1 13072 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_38
timestamp 1300117811
transform 0 1 13158 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_39
timestamp 1300117811
transform 0 1 13244 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_40
timestamp 1300117811
transform 0 1 13330 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_41
timestamp 1300117811
transform 0 1 13416 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_42
timestamp 1300117811
transform 0 1 13502 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_1
timestamp 1300115302
transform 0 1 13588 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_43
timestamp 1300117811
transform 0 1 15308 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_44
timestamp 1300117811
transform 0 1 15394 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_45
timestamp 1300117811
transform 0 1 15480 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_46
timestamp 1300117811
transform 0 1 15566 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_47
timestamp 1300117811
transform 0 1 15652 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_48
timestamp 1300117811
transform 0 1 15738 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_49
timestamp 1300117811
transform 0 1 15824 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_50
timestamp 1300117811
transform 0 1 15910 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_51
timestamp 1300117811
transform 0 1 15996 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_52
timestamp 1300117811
transform 0 1 16082 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_53
timestamp 1300117811
transform 0 1 16168 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_54
timestamp 1300117811
transform 0 1 16254 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_55
timestamp 1300117811
transform 0 1 16340 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_56
timestamp 1300117811
transform 0 1 16426 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_57
timestamp 1300117811
transform 0 1 16512 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_58
timestamp 1300117811
transform 0 1 16598 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_59
timestamp 1300117811
transform 0 1 16684 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_60
timestamp 1300117811
transform 0 1 16770 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_61
timestamp 1300117811
transform 0 1 16856 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_62
timestamp 1300117811
transform 0 1 16942 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_63
timestamp 1300117811
transform 0 1 17028 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_2
timestamp 1300115302
transform 0 1 17114 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_64
timestamp 1300117811
transform 0 1 18834 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_65
timestamp 1300117811
transform 0 1 18920 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_66
timestamp 1300117811
transform 0 1 19006 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_67
timestamp 1300117811
transform 0 1 19092 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_68
timestamp 1300117811
transform 0 1 19178 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_69
timestamp 1300117811
transform 0 1 19264 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_70
timestamp 1300117811
transform 0 1 19350 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_71
timestamp 1300117811
transform 0 1 19436 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_72
timestamp 1300117811
transform 0 1 19522 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_73
timestamp 1300117811
transform 0 1 19608 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_74
timestamp 1300117811
transform 0 1 19694 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_75
timestamp 1300117811
transform 0 1 19780 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_76
timestamp 1300117811
transform 0 1 19866 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_77
timestamp 1300117811
transform 0 1 19952 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_78
timestamp 1300117811
transform 0 1 20038 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_79
timestamp 1300117811
transform 0 1 20124 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_80
timestamp 1300117811
transform 0 1 20210 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_81
timestamp 1300117811
transform 0 1 20296 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_82
timestamp 1300117811
transform 0 1 20382 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_83
timestamp 1300117811
transform 0 1 20468 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_84
timestamp 1300117811
transform 0 1 20554 -1 0 6450
box 0 0 6450 86
use zgppxpp_mt VDDpads_0
timestamp 1300121810
transform 0 1 20640 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_85
timestamp 1300117811
transform 0 1 22360 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_86
timestamp 1300117811
transform 0 1 22446 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_87
timestamp 1300117811
transform 0 1 22532 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_88
timestamp 1300117811
transform 0 1 22618 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_89
timestamp 1300117811
transform 0 1 22704 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_90
timestamp 1300117811
transform 0 1 22790 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_91
timestamp 1300117811
transform 0 1 22876 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_92
timestamp 1300117811
transform 0 1 22962 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_93
timestamp 1300117811
transform 0 1 23048 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_94
timestamp 1300117811
transform 0 1 23134 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_95
timestamp 1300117811
transform 0 1 23220 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_96
timestamp 1300117811
transform 0 1 23306 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_97
timestamp 1300117811
transform 0 1 23392 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_98
timestamp 1300117811
transform 0 1 23478 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_99
timestamp 1300117811
transform 0 1 23564 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_100
timestamp 1300117811
transform 0 1 23650 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_101
timestamp 1300117811
transform 0 1 23736 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_102
timestamp 1300117811
transform 0 1 23822 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_103
timestamp 1300117811
transform 0 1 23908 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_104
timestamp 1300117811
transform 0 1 23994 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_105
timestamp 1300117811
transform 0 1 24080 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_3
timestamp 1300115302
transform 0 1 24166 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_106
timestamp 1300117811
transform 0 1 25886 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_107
timestamp 1300117811
transform 0 1 25972 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_108
timestamp 1300117811
transform 0 1 26058 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_109
timestamp 1300117811
transform 0 1 26144 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_110
timestamp 1300117811
transform 0 1 26230 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_111
timestamp 1300117811
transform 0 1 26316 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_112
timestamp 1300117811
transform 0 1 26402 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_113
timestamp 1300117811
transform 0 1 26488 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_114
timestamp 1300117811
transform 0 1 26574 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_115
timestamp 1300117811
transform 0 1 26660 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_116
timestamp 1300117811
transform 0 1 26746 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_117
timestamp 1300117811
transform 0 1 26832 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_118
timestamp 1300117811
transform 0 1 26918 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_119
timestamp 1300117811
transform 0 1 27004 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_120
timestamp 1300117811
transform 0 1 27090 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_121
timestamp 1300117811
transform 0 1 27176 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_122
timestamp 1300117811
transform 0 1 27262 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_123
timestamp 1300117811
transform 0 1 27348 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_124
timestamp 1300117811
transform 0 1 27434 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_125
timestamp 1300117811
transform 0 1 27520 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_126
timestamp 1300117811
transform 0 1 27606 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_4
timestamp 1300115302
transform 0 1 27692 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_127
timestamp 1300117811
transform 0 1 29412 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_128
timestamp 1300117811
transform 0 1 29498 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_129
timestamp 1300117811
transform 0 1 29584 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_130
timestamp 1300117811
transform 0 1 29670 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_131
timestamp 1300117811
transform 0 1 29756 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_132
timestamp 1300117811
transform 0 1 29842 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_133
timestamp 1300117811
transform 0 1 29928 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_134
timestamp 1300117811
transform 0 1 30014 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_135
timestamp 1300117811
transform 0 1 30100 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_136
timestamp 1300117811
transform 0 1 30186 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_137
timestamp 1300117811
transform 0 1 30272 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_138
timestamp 1300117811
transform 0 1 30358 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_139
timestamp 1300117811
transform 0 1 30444 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_140
timestamp 1300117811
transform 0 1 30530 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_141
timestamp 1300117811
transform 0 1 30616 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_142
timestamp 1300117811
transform 0 1 30702 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_143
timestamp 1300117811
transform 0 1 30788 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_144
timestamp 1300117811
transform 0 1 30874 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_145
timestamp 1300117811
transform 0 1 30960 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_146
timestamp 1300117811
transform 0 1 31046 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_147
timestamp 1300117811
transform 0 1 31132 -1 0 6450
box 0 0 6450 86
use ioacx6xxcsxe04_mt Data_5
timestamp 1300115302
transform 0 1 31218 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_148
timestamp 1300117811
transform 0 1 32938 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_149
timestamp 1300117811
transform 0 1 33024 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_150
timestamp 1300117811
transform 0 1 33110 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_151
timestamp 1300117811
transform 0 1 33196 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_152
timestamp 1300117811
transform 0 1 33282 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_153
timestamp 1300117811
transform 0 1 33368 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_154
timestamp 1300117811
transform 0 1 33454 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_155
timestamp 1300117811
transform 0 1 33540 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_156
timestamp 1300117811
transform 0 1 33626 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_157
timestamp 1300117811
transform 0 1 33712 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_158
timestamp 1300117811
transform 0 1 33798 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_159
timestamp 1300117811
transform 0 1 33884 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_160
timestamp 1300117811
transform 0 1 33970 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_161
timestamp 1300117811
transform 0 1 34056 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_162
timestamp 1300117811
transform 0 1 34142 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_163
timestamp 1300117811
transform 0 1 34228 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_164
timestamp 1300117811
transform 0 1 34314 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_165
timestamp 1300117811
transform 0 1 34400 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_166
timestamp 1300117811
transform 0 1 34486 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_167
timestamp 1300117811
transform 0 1 34572 -1 0 6450
box 0 0 6450 86
use fillpp_mt fillpp_mt_168
timestamp 1300117811
transform 0 1 34658 -1 0 6450
box 0 0 6450 86
use zgppxpg_mt VSSPads_1
timestamp 1300122446
transform 0 1 34744 -1 0 6450
box 0 0 6450 1720
use fillpp_mt fillpp_mt_169
timestamp 1300117811
transform 0 1 36464 -1 0 6450
box 0 0 6450 86
use corns_clamp_mt CORNER_1
timestamp 1300118495
transform 0 -1 43000 1 0 0
box 0 0 6450 6450
<< labels >>
rlabel metal4 6616 78 8176 1638 0 nIRQ
rlabel metal4 10142 78 11702 1638 0 Data[0]
rlabel metal4 13668 78 15228 1638 0 Data[1]
rlabel metal4 17194 78 18754 1638 0 Data[2]
rlabel metal4 20720 78 22280 1638 0 vdde!
rlabel metal4 24246 78 25806 1638 0 Data[3]
rlabel metal4 27772 78 29332 1638 0 Data[4]
rlabel metal4 31298 78 32858 1638 0 Data[5]
rlabel metal4 34824 78 36384 1638 0 gnde!
rlabel metal4 41362 6530 42922 8090 0 Data[6]
rlabel metal4 41362 11002 42922 12562 0 Data[7]
rlabel metal4 41362 15474 42922 17034 0 Data[8]
rlabel metal4 41362 19946 42922 21506 0 gnde!
rlabel metal4 41362 24418 42922 25978 0 GND!
rlabel metal4 41362 28890 42922 30450 0 Data[9]
rlabel metal4 41362 33362 42922 34922 0 Data[10]
rlabel metal4 41362 37834 42922 39394 0 Data[11]
rlabel metal4 34824 44286 36384 45846 0 vdde!
rlabel metal4 31298 44286 32858 45846 0 Data[12]
rlabel metal4 27772 44286 29332 45846 0 Data[13]
rlabel metal4 24246 44286 25806 45846 0 Data[14]
rlabel metal4 20720 44286 22280 45846 0 gnde!
rlabel metal4 17194 44286 18754 45846 0 Data[15]
rlabel metal4 13668 44286 15228 45846 0 ALE
rlabel metal4 10142 44286 11702 45846 0 nME
rlabel metal4 6616 44286 8176 45846 0 nWait
rlabel metal4 78 37834 1638 39394 0 nOE
rlabel metal4 78 33362 1638 34922 0 RnW
rlabel metal4 78 28890 1638 30450 0 SDO
rlabel metal4 78 24418 1638 25978 0 Vdd!
rlabel metal4 78 19946 1638 21506 0 SDI
rlabel metal4 78 15474 1638 17034 0 Test
rlabel metal4 78 11002 1638 12562 0 Clock
rlabel metal4 78 6530 1638 8090 0 nReset
<< end >>
