magic
tech c035u
timestamp 1394198348
<< metal1 >>
rect 1293 3900 1807 3910
rect 1821 3900 2647 3910
rect 2661 3900 3583 3910
rect 3597 3900 4375 3910
rect 4389 3900 5095 3910
rect 5109 3900 5863 3910
rect 5877 3900 6751 3910
rect 1269 3878 1783 3888
rect 1797 3878 2767 3888
rect 2781 3878 3487 3888
rect 3501 3878 4255 3888
rect 4269 3878 5191 3888
rect 5205 3878 5839 3888
rect 5853 3878 6631 3888
rect 1245 3855 1927 3865
rect 1941 3855 2623 3865
rect 2637 3855 3463 3865
rect 3477 3855 4231 3865
rect 4245 3855 5071 3865
rect 5085 3855 5959 3865
rect 5973 3855 6607 3865
rect 1701 3832 2407 3842
rect 2421 3832 3247 3842
rect 3261 3832 4135 3842
rect 4149 3832 4975 3842
rect 4989 3832 5647 3842
rect 5661 3832 6415 3842
rect 6429 3832 7351 3842
rect 1677 3810 2383 3820
rect 2397 3810 3367 3820
rect 3381 3810 4039 3820
rect 4053 3810 4855 3820
rect 4869 3810 5743 3820
rect 5757 3810 6391 3820
rect 6405 3810 7231 3820
rect 1653 3787 2527 3797
rect 2541 3787 3223 3797
rect 3237 3787 4015 3797
rect 4029 3787 4831 3797
rect 4845 3787 5623 3797
rect 5637 3787 6511 3797
rect 6525 3787 7207 3797
rect 1557 3764 2167 3774
rect 2181 3764 3007 3774
rect 3021 3764 3919 3774
rect 3933 3764 4735 3774
rect 4749 3764 5431 3774
rect 5445 3764 6199 3774
rect 6213 3764 7111 3774
rect 1533 3742 2143 3752
rect 2157 3742 3127 3752
rect 3141 3742 3823 3752
rect 3837 3742 4615 3752
rect 4629 3742 5527 3752
rect 5541 3742 6175 3752
rect 6189 3742 6991 3752
rect 1509 3719 2287 3729
rect 2301 3719 2983 3729
rect 2997 3719 3799 3729
rect 3813 3719 4591 3729
rect 4605 3719 5407 3729
rect 5421 3719 6295 3729
rect 6309 3719 6967 3729
rect 0 1021 73 1031
rect 88 1021 1225 1031
rect 1239 1021 2377 1031
rect 2392 1021 3529 1031
rect 3543 1021 4681 1031
rect 4695 1021 5833 1031
rect 5847 1021 6984 1031
rect 6999 1021 8137 1031
rect 664 984 793 994
rect 807 984 1009 994
rect 1814 971 1945 981
rect 1959 971 2161 981
rect 2966 971 3097 981
rect 3111 971 3313 981
rect 4118 971 4249 981
rect 4263 971 4465 981
rect 5270 971 5401 981
rect 5415 971 5617 981
rect 6422 971 6553 981
rect 6567 971 6769 981
rect 7574 971 7705 981
rect 7719 971 7921 981
rect 8726 971 8857 981
rect 8871 971 9073 981
rect 0 928 50 938
rect 9266 928 9385 938
rect 0 905 50 915
rect 9266 905 9385 915
rect 0 867 50 892
rect 9266 867 9385 892
rect 0 222 50 247
rect 9266 222 9385 247
rect 0 199 50 209
rect 9266 199 9385 209
rect 0 176 50 186
rect 9266 176 9385 186
rect 0 153 50 163
rect 9266 153 9385 163
rect 0 60 936 70
rect 951 60 2088 70
rect 2103 60 3240 70
rect 3255 60 4393 70
rect 4408 60 5543 70
rect 5561 60 6695 70
rect 6713 60 7847 70
rect 7865 60 9001 70
rect 9015 60 9385 70
rect 0 25 1153 35
rect 1167 25 2305 35
rect 2319 25 3457 35
rect 3471 25 4609 35
rect 4624 25 5760 35
rect 5778 25 6912 35
rect 6930 25 8064 35
rect 8082 25 9217 35
rect 9231 25 9385 35
<< m2contact >>
rect 1279 3898 1293 3912
rect 1807 3898 1821 3912
rect 2647 3898 2661 3912
rect 3583 3898 3597 3912
rect 4375 3898 4389 3912
rect 5095 3898 5109 3912
rect 5863 3898 5877 3912
rect 6751 3898 6765 3912
rect 1255 3876 1269 3890
rect 1783 3876 1797 3890
rect 2767 3876 2781 3890
rect 3487 3876 3501 3890
rect 4255 3876 4269 3890
rect 5191 3876 5205 3890
rect 5839 3876 5853 3890
rect 6631 3876 6645 3890
rect 1231 3853 1245 3867
rect 1927 3853 1941 3867
rect 2623 3853 2637 3867
rect 3463 3853 3477 3867
rect 4231 3853 4245 3867
rect 5071 3853 5085 3867
rect 5959 3853 5973 3867
rect 6607 3853 6621 3867
rect 1687 3830 1701 3844
rect 2407 3830 2421 3844
rect 3247 3830 3261 3844
rect 4135 3830 4149 3844
rect 4975 3830 4989 3844
rect 5647 3830 5661 3844
rect 6415 3830 6429 3844
rect 7351 3830 7365 3844
rect 1663 3808 1677 3822
rect 2383 3808 2397 3822
rect 3367 3808 3381 3822
rect 4039 3808 4053 3822
rect 4855 3808 4869 3822
rect 5743 3808 5757 3822
rect 6391 3808 6405 3822
rect 7231 3808 7245 3822
rect 1639 3785 1653 3799
rect 2527 3785 2541 3799
rect 3223 3785 3237 3799
rect 4015 3785 4029 3799
rect 4831 3785 4845 3799
rect 5623 3785 5637 3799
rect 6511 3785 6525 3799
rect 7207 3785 7221 3799
rect 1543 3762 1557 3776
rect 2167 3762 2181 3776
rect 3007 3762 3021 3776
rect 3919 3762 3933 3776
rect 4735 3762 4749 3776
rect 5431 3762 5445 3776
rect 6199 3762 6213 3776
rect 7111 3762 7125 3776
rect 1519 3740 1533 3754
rect 2143 3740 2157 3754
rect 3127 3740 3141 3754
rect 3823 3740 3837 3754
rect 4615 3740 4629 3754
rect 5527 3740 5541 3754
rect 6175 3740 6189 3754
rect 6991 3740 7005 3754
rect 1495 3717 1509 3731
rect 2287 3717 2301 3731
rect 2983 3717 2997 3731
rect 3799 3717 3813 3731
rect 4591 3717 4605 3731
rect 5407 3717 5421 3731
rect 6295 3717 6309 3731
rect 6967 3717 6981 3731
rect 73 1018 88 1034
rect 1225 1020 1239 1034
rect 2377 1020 2392 1034
rect 3529 1020 3543 1034
rect 4681 1020 4695 1034
rect 5833 1020 5847 1034
rect 6984 1019 6999 1033
rect 8137 1020 8152 1035
rect 649 983 664 997
rect 793 982 807 996
rect 1009 981 1023 995
rect 1800 969 1814 983
rect 1945 968 1959 982
rect 2161 969 2175 983
rect 2952 969 2966 983
rect 3097 968 3111 982
rect 3313 969 3327 983
rect 4104 969 4118 983
rect 4249 968 4263 982
rect 4465 969 4479 983
rect 5256 969 5270 983
rect 5401 968 5415 982
rect 5617 969 5631 983
rect 6408 969 6422 983
rect 6553 968 6567 982
rect 6769 969 6783 983
rect 7560 969 7574 983
rect 7705 968 7719 982
rect 7921 969 7935 983
rect 8712 969 8726 983
rect 8857 968 8871 982
rect 9073 969 9087 983
rect 936 58 951 72
rect 2088 58 2103 72
rect 3240 58 3255 72
rect 4393 58 4408 73
rect 5543 58 5561 73
rect 6695 58 6713 73
rect 7847 58 7865 73
rect 9001 57 9015 72
rect 1153 24 1167 38
rect 2305 24 2319 38
rect 3457 24 3471 38
rect 4609 23 4624 38
rect 5760 20 5778 35
rect 6912 20 6930 35
rect 8064 20 8082 35
rect 9217 23 9231 38
<< metal2 >>
rect 1232 3867 1244 3969
rect 1256 3890 1268 3969
rect 1280 3912 1292 3969
rect 1330 3934 1342 3969
rect 1330 3922 1489 3934
rect 1777 3922 2126 3934
rect 2606 3922 2975 3934
rect 3455 3922 3794 3934
rect 4226 3922 4582 3934
rect 5062 3922 5398 3934
rect 5830 3922 6163 3934
rect 6595 3922 6884 3934
rect 1232 3688 1244 3853
rect 1256 3688 1268 3876
rect 1280 3688 1292 3898
rect 1400 3688 1412 3922
rect 1640 3799 1652 3866
rect 1664 3822 1676 3866
rect 1688 3844 1700 3866
rect 1496 3731 1508 3798
rect 1520 3754 1532 3798
rect 1544 3776 1556 3798
rect 1496 3688 1508 3717
rect 1520 3688 1532 3740
rect 1544 3688 1556 3762
rect 1640 3688 1652 3785
rect 1664 3688 1676 3808
rect 1688 3688 1700 3830
rect 1784 3688 1796 3876
rect 1808 3688 1820 3898
rect 1928 3688 1940 3853
rect 2048 3688 2060 3922
rect 2144 3688 2156 3740
rect 2168 3688 2180 3762
rect 2288 3688 2300 3717
rect 2384 3688 2396 3808
rect 2408 3688 2420 3830
rect 2528 3688 2540 3785
rect 2624 3688 2636 3853
rect 2648 3688 2660 3898
rect 2768 3688 2780 3876
rect 2888 3688 2900 3922
rect 2984 3688 2996 3717
rect 3008 3688 3020 3762
rect 3128 3688 3140 3740
rect 3224 3688 3236 3785
rect 3248 3688 3260 3830
rect 3368 3688 3380 3808
rect 3464 3688 3476 3853
rect 3488 3688 3500 3876
rect 3584 3688 3596 3898
rect 3704 3688 3716 3922
rect 3800 3688 3812 3717
rect 3824 3688 3836 3740
rect 3920 3688 3932 3762
rect 4016 3688 4028 3785
rect 4040 3688 4052 3808
rect 4136 3688 4148 3830
rect 4232 3688 4244 3853
rect 4256 3688 4268 3876
rect 4376 3688 4388 3898
rect 4496 3688 4508 3922
rect 4592 3688 4604 3717
rect 4616 3688 4628 3740
rect 4736 3688 4748 3762
rect 4832 3688 4844 3785
rect 4856 3688 4868 3808
rect 4976 3688 4988 3830
rect 5072 3688 5084 3853
rect 5096 3688 5108 3898
rect 5192 3688 5204 3876
rect 5312 3688 5324 3922
rect 5408 3688 5420 3717
rect 5432 3688 5444 3762
rect 5528 3688 5540 3740
rect 5624 3688 5636 3785
rect 5648 3688 5660 3830
rect 5744 3688 5756 3808
rect 5840 3688 5852 3876
rect 5864 3688 5876 3898
rect 5960 3688 5972 3853
rect 6080 3688 6092 3922
rect 6176 3688 6188 3740
rect 6200 3688 6212 3762
rect 6296 3688 6308 3717
rect 6392 3688 6404 3808
rect 6416 3688 6428 3830
rect 6512 3688 6524 3785
rect 6608 3688 6620 3853
rect 6632 3688 6644 3876
rect 6752 3688 6764 3898
rect 6872 3688 6884 3922
rect 6968 3688 6980 3717
rect 6992 3688 7004 3740
rect 7112 3688 7124 3762
rect 7208 3688 7220 3785
rect 7232 3688 7244 3808
rect 7352 3688 7364 3830
rect 1328 2877 1388 2889
rect 1448 2852 1460 2889
rect 1592 2844 1604 2889
rect 1736 2844 1748 2889
rect 1856 2877 1916 2889
rect 1976 2877 2036 2889
rect 2096 2852 2108 2889
rect 2216 2877 2276 2889
rect 2336 2844 2348 2889
rect 2456 2877 2516 2889
rect 2576 2844 2588 2889
rect 2696 2877 2756 2889
rect 2816 2877 2876 2889
rect 2936 2852 2948 2890
rect 5288 2889 5300 2891
rect 6056 2889 6068 2891
rect 3056 2877 3116 2889
rect 3176 2844 3188 2889
rect 3296 2877 3356 2889
rect 3416 2844 3428 2889
rect 3512 2877 3572 2889
rect 3632 2877 3692 2889
rect 3752 2852 3764 2889
rect 3848 2877 3908 2889
rect 3968 2844 3980 2889
rect 4064 2877 4124 2889
rect 4184 2844 4196 2889
rect 4304 2877 4364 2889
rect 4424 2877 4484 2889
rect 4544 2852 4556 2889
rect 4664 2877 4724 2889
rect 4784 2844 4796 2889
rect 4904 2877 4964 2889
rect 5024 2844 5036 2889
rect 5120 2877 5180 2889
rect 5240 2877 5300 2889
rect 5360 2852 5372 2889
rect 5456 2877 5516 2889
rect 5576 2844 5588 2889
rect 5672 2877 5732 2889
rect 5792 2844 5804 2889
rect 5888 2877 5948 2889
rect 6008 2877 6068 2889
rect 6128 2852 6140 2889
rect 6224 2877 6284 2889
rect 6344 2880 6356 2889
rect 6344 2863 6359 2880
rect 6440 2877 6500 2889
rect 6347 2861 6359 2863
rect 6560 2844 6572 2889
rect 6680 2877 6740 2889
rect 6800 2877 6860 2889
rect 6920 2852 6932 2889
rect 7040 2877 7100 2889
rect 7160 2844 7172 2889
rect 7280 2877 7340 2889
rect 7400 2844 7412 2889
rect 74 945 86 1018
rect 122 945 134 1075
rect 650 945 662 983
rect 794 945 806 982
rect 866 945 878 1075
rect 1010 945 1022 981
rect 1082 945 1094 1075
rect 1226 945 1238 1020
rect 1274 945 1286 1075
rect 1802 945 1814 969
rect 1946 945 1958 968
rect 2018 945 2030 1075
rect 2162 945 2174 969
rect 2234 945 2246 1075
rect 2378 945 2390 1020
rect 2426 945 2438 1075
rect 2954 945 2966 969
rect 3098 945 3110 968
rect 3170 945 3182 1075
rect 3314 945 3326 969
rect 3386 945 3398 1075
rect 3530 945 3542 1020
rect 3578 945 3590 1075
rect 4106 945 4118 969
rect 4250 945 4262 968
rect 4322 945 4334 1075
rect 4466 945 4478 969
rect 4538 945 4550 1075
rect 4682 945 4694 1020
rect 4730 945 4742 1075
rect 5258 945 5270 969
rect 5402 945 5414 968
rect 5474 945 5486 1075
rect 5618 945 5630 969
rect 5690 945 5702 1075
rect 5834 945 5846 1020
rect 5882 945 5894 1075
rect 6410 945 6422 969
rect 6554 945 6566 968
rect 6626 945 6638 1075
rect 6770 945 6782 969
rect 6842 945 6854 1075
rect 6986 945 6998 1019
rect 7034 945 7046 1075
rect 7562 945 7574 969
rect 7706 945 7718 968
rect 7778 945 7790 1075
rect 7922 945 7934 969
rect 7994 945 8006 1075
rect 8138 945 8150 1020
rect 8186 945 8198 1075
rect 8714 945 8726 969
rect 8858 945 8870 968
rect 8930 945 8942 1075
rect 9074 945 9086 969
rect 9146 945 9158 1075
rect 122 0 134 146
rect 866 0 878 146
rect 938 72 950 146
rect 1082 0 1094 146
rect 1154 38 1166 146
rect 1274 0 1286 146
rect 2018 0 2030 146
rect 2090 72 2102 146
rect 2234 0 2246 146
rect 2306 38 2318 146
rect 2426 0 2438 146
rect 3170 0 3182 146
rect 3242 72 3254 146
rect 3386 0 3398 146
rect 3458 38 3470 146
rect 3578 0 3590 146
rect 4322 0 4334 146
rect 4394 73 4406 146
rect 4538 0 4550 146
rect 4610 38 4622 146
rect 4730 0 4742 146
rect 5474 0 5486 146
rect 5546 73 5558 146
rect 5690 0 5702 146
rect 5762 35 5774 146
rect 5882 0 5894 146
rect 6626 0 6638 146
rect 6698 73 6710 146
rect 6842 0 6854 146
rect 6914 35 6926 146
rect 7034 0 7046 146
rect 7778 0 7790 146
rect 7850 73 7862 146
rect 7994 0 8006 146
rect 8066 35 8078 146
rect 8186 0 8198 146
rect 8930 0 8942 146
rect 9002 72 9014 146
rect 9146 0 9158 146
rect 9218 38 9230 146
use nor3  nor3_2
timestamp 1386235396
transform 1 0 1208 0 1 2889
box 0 0 144 799
use and2  and2_10
timestamp 1386234845
transform 1 0 1352 0 1 2889
box 0 0 120 799
use nor3  nor3_0
timestamp 1386235396
transform 1 0 1472 0 1 2889
box 0 0 144 799
use nor3  nor3_1
timestamp 1386235396
transform 1 0 1616 0 1 2889
box 0 0 144 799
use nor2  nor2_12
timestamp 1386235306
transform 1 0 1760 0 1 2889
box 0 0 120 799
use and2  and2_11
timestamp 1386234845
transform 1 0 1880 0 1 2889
box 0 0 120 799
use and2  and2_12
timestamp 1386234845
transform 1 0 2000 0 1 2889
box 0 0 120 799
use nor2  nor2_0
timestamp 1386235306
transform 1 0 2120 0 1 2889
box 0 0 120 799
use and2  and2_0
timestamp 1386234845
transform 1 0 2240 0 1 2889
box 0 0 120 799
use nor2  nor2_6
timestamp 1386235306
transform 1 0 2360 0 1 2889
box 0 0 120 799
use and2  and2_5
timestamp 1386234845
transform 1 0 2480 0 1 2889
box 0 0 120 799
use nor2  nor2_13
timestamp 1386235306
transform 1 0 2600 0 1 2889
box 0 0 120 799
use and2  and2_13
timestamp 1386234845
transform 1 0 2720 0 1 2889
box 0 0 120 799
use and2  and2_14
timestamp 1386234845
transform 1 0 2840 0 1 2889
box 0 0 120 799
use nor2  nor2_1
timestamp 1386235306
transform 1 0 2960 0 1 2889
box 0 0 120 799
use and2  and2_1
timestamp 1386234845
transform 1 0 3080 0 1 2889
box 0 0 120 799
use nor2  nor2_7
timestamp 1386235306
transform 1 0 3200 0 1 2889
box 0 0 120 799
use and2  and2_6
timestamp 1386234845
transform 1 0 3320 0 1 2889
box 0 0 120 799
use nand2  nand2_6
timestamp 1386234792
transform 1 0 3440 0 1 2889
box 0 0 96 799
use nor2  nor2_14
timestamp 1386235306
transform 1 0 3536 0 1 2889
box 0 0 120 799
use and2  and2_15
timestamp 1386234845
transform 1 0 3656 0 1 2889
box 0 0 120 799
use nand2  nand2_0
timestamp 1386234792
transform 1 0 3776 0 1 2889
box 0 0 96 799
use nor2  nor2_2
timestamp 1386235306
transform 1 0 3872 0 1 2889
box 0 0 120 799
use nand2  nand2_3
timestamp 1386234792
transform 1 0 3992 0 1 2889
box 0 0 96 799
use nor2  nor2_8
timestamp 1386235306
transform 1 0 4088 0 1 2889
box 0 0 120 799
use nor2  nor2_15
timestamp 1386235306
transform 1 0 4208 0 1 2889
box 0 0 120 799
use and2  and2_16
timestamp 1386234845
transform 1 0 4328 0 1 2889
box 0 0 120 799
use and2  and2_17
timestamp 1386234845
transform 1 0 4448 0 1 2889
box 0 0 120 799
use nor2  nor2_3
timestamp 1386235306
transform 1 0 4568 0 1 2889
box 0 0 120 799
use and2  and2_2
timestamp 1386234845
transform 1 0 4688 0 1 2889
box 0 0 120 799
use nor2  nor2_9
timestamp 1386235306
transform 1 0 4808 0 1 2889
box 0 0 120 799
use and2  and2_7
timestamp 1386234845
transform 1 0 4928 0 1 2889
box 0 0 120 799
use nand2  nand2_7
timestamp 1386234792
transform 1 0 5048 0 1 2889
box 0 0 96 799
use nor2  nor2_16
timestamp 1386235306
transform 1 0 5144 0 1 2889
box 0 0 120 799
use and2  and2_18
timestamp 1386234845
transform 1 0 5264 0 1 2889
box 0 0 120 799
use nand2  nand2_1
timestamp 1386234792
transform 1 0 5384 0 1 2889
box 0 0 96 799
use nor2  nor2_4
timestamp 1386235306
transform 1 0 5480 0 1 2889
box 0 0 120 799
use nand2  nand2_4
timestamp 1386234792
transform 1 0 5600 0 1 2889
box 0 0 96 799
use nor2  nor2_10
timestamp 1386235306
transform 1 0 5696 0 1 2889
box 0 0 120 799
use nand2  nand2_8
timestamp 1386234792
transform 1 0 5816 0 1 2889
box 0 0 96 799
use nor2  nor2_17
timestamp 1386235306
transform 1 0 5912 0 1 2889
box 0 0 120 799
use and2  and2_19
timestamp 1386234845
transform 1 0 6032 0 1 2889
box 0 0 120 799
use nand2  nand2_2
timestamp 1386234792
transform 1 0 6152 0 1 2889
box 0 0 96 799
use nor2  nor2_5
timestamp 1386235306
transform 1 0 6248 0 1 2889
box 0 0 120 799
use nand2  nand2_5
timestamp 1386234792
transform 1 0 6368 0 1 2889
box 0 0 96 799
use nor2  nor2_11
timestamp 1386235306
transform 1 0 6464 0 1 2889
box 0 0 120 799
use and2  and2_20
timestamp 1386234845
transform 1 0 6584 0 1 2889
box 0 0 120 799
use and2  and2_21
timestamp 1386234845
transform 1 0 6704 0 1 2889
box 0 0 120 799
use and2  and2_22
timestamp 1386234845
transform 1 0 6824 0 1 2889
box 0 0 120 799
use and2  and2_3
timestamp 1386234845
transform 1 0 6944 0 1 2889
box 0 0 120 799
use and2  and2_4
timestamp 1386234845
transform 1 0 7064 0 1 2889
box 0 0 120 799
use and2  and2_8
timestamp 1386234845
transform 1 0 7184 0 1 2889
box 0 0 120 799
use and2  and2_9
timestamp 1386234845
transform 1 0 7304 0 1 2889
box 0 0 120 799
use scanreg  scanreg_1
timestamp 1386241447
transform 1 0 50 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_0
timestamp 1386237216
transform 1 0 770 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_1
timestamp 1386237216
transform 1 0 986 0 1 146
box 0 0 216 799
use scanreg  scanreg_2
timestamp 1386241447
transform 1 0 1202 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_2
timestamp 1386237216
transform 1 0 1922 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_3
timestamp 1386237216
transform 1 0 2138 0 1 146
box 0 0 216 799
use scanreg  scanreg_3
timestamp 1386241447
transform 1 0 2354 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_4
timestamp 1386237216
transform 1 0 3074 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_5
timestamp 1386237216
transform 1 0 3290 0 1 146
box 0 0 216 799
use scanreg  scanreg_4
timestamp 1386241447
transform 1 0 3506 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_6
timestamp 1386237216
transform 1 0 4226 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_7
timestamp 1386237216
transform 1 0 4442 0 1 146
box 0 0 216 799
use scanreg  scanreg_5
timestamp 1386241447
transform 1 0 4658 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_8
timestamp 1386237216
transform 1 0 5378 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_9
timestamp 1386237216
transform 1 0 5594 0 1 146
box 0 0 216 799
use scanreg  scanreg_6
timestamp 1386241447
transform 1 0 5810 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_10
timestamp 1386237216
transform 1 0 6530 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_11
timestamp 1386237216
transform 1 0 6746 0 1 146
box 0 0 216 799
use scanreg  scanreg_7
timestamp 1386241447
transform 1 0 6962 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_12
timestamp 1386237216
transform 1 0 7682 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_13
timestamp 1386237216
transform 1 0 7898 0 1 146
box 0 0 216 799
use scanreg  scanreg_8
timestamp 1386241447
transform 1 0 8114 0 1 146
box 0 0 720 799
use trisbuf  trisbuf_14
timestamp 1386237216
transform 1 0 8834 0 1 146
box 0 0 216 799
use trisbuf  trisbuf_15
timestamp 1386237216
transform 1 0 9050 0 1 146
box 0 0 216 799
<< labels >>
rlabel metal1 0 1021 0 1031 1 WData
rlabel metal1 0 60 0 70 3 Rd1
rlabel metal1 0 25 0 35 3 Rd2
rlabel metal1 0 928 0 938 3 ScanReturn
rlabel metal1 0 905 0 915 3 SDI
rlabel metal1 0 153 0 163 3 nReset
rlabel metal1 0 176 0 186 3 Test
rlabel metal1 0 199 0 209 3 Clock
rlabel metal1 0 222 0 247 3 GND!
rlabel metal1 0 867 0 892 3 Vdd!
rlabel metal2 5474 1075 5486 1075 5 Rs1[4]
rlabel metal2 4730 1075 4742 1075 5 Rw[4]
rlabel metal2 4538 1075 4550 1075 5 Rs2[3]
rlabel metal2 4322 1075 4334 1075 5 Rs1[3]
rlabel metal2 3578 1075 3590 1075 5 Rw[3]
rlabel metal2 3386 1075 3398 1075 5 Rs2[2]
rlabel metal2 3170 1075 3182 1075 5 Rs1[2]
rlabel metal2 2426 1075 2438 1075 5 Rw[2]
rlabel metal2 2234 1075 2246 1075 5 Rs2[1]
rlabel metal2 2018 1075 2030 1075 5 Rs1[1]
rlabel metal2 1274 1075 1286 1075 5 Rw[1]
rlabel metal2 1082 1075 1094 1075 5 Rs2[0]
rlabel metal2 866 1075 878 1075 5 Rs1[0]
rlabel metal2 122 0 134 0 1 Rw[0]
rlabel metal2 1082 0 1094 0 5 Rs2[0]
rlabel metal2 1274 0 1286 0 5 Rw[1]
rlabel metal2 2018 0 2030 0 5 Rs1[1]
rlabel metal2 3170 0 3182 0 5 Rs1[2]
rlabel metal2 3578 0 3590 0 5 Rw[3]
rlabel metal2 3386 0 3398 0 5 Rs2[2]
rlabel metal2 4322 0 4334 0 5 Rs1[3]
rlabel metal2 4730 0 4742 0 5 Rw[4]
rlabel metal2 4538 0 4550 0 5 Rs2[3]
rlabel metal2 5474 0 5486 0 5 Rs1[4]
rlabel metal2 2426 0 2438 0 1 Rw[2]
rlabel metal2 5690 0 5702 0 1 Rs2[4]
rlabel metal2 7778 0 7790 0 5 Rs1[6]
rlabel metal2 9146 0 9158 0 5 Rs2[7]
rlabel metal2 8930 0 8942 0 5 Rs1[7]
rlabel metal2 8186 0 8198 0 5 Rw[7]
rlabel metal2 7994 0 8006 0 5 Rs2[6]
rlabel metal2 7034 0 7046 0 5 Rw[6]
rlabel metal2 6842 0 6854 0 5 Rs2[5]
rlabel metal2 6626 0 6638 0 5 Rs1[5]
rlabel metal2 5882 0 5894 0 5 Rw[5]
rlabel metal2 5690 1075 5702 1075 5 Rs2[4]
rlabel metal2 5882 1075 5894 1075 5 Rw[5]
rlabel metal2 6626 1075 6638 1075 5 Rs1[5]
rlabel metal2 6842 1075 6854 1075 5 Rs2[5]
rlabel metal2 7034 1075 7046 1075 5 Rw[6]
rlabel metal2 7778 1075 7790 1075 5 Rs1[6]
rlabel metal2 7994 1075 8006 1075 5 Rs2[6]
rlabel metal2 8930 1075 8942 1075 5 Rs1[7]
rlabel metal2 9146 1075 9158 1075 5 Rs2[7]
rlabel metal2 8186 1075 8198 1075 5 Rw[7]
rlabel metal1 9385 25 9385 35 7 Rd2
rlabel metal1 9385 60 9385 70 7 Rd1
rlabel metal1 9385 905 9385 915 7 Scan
rlabel metal1 9385 928 9385 938 7 ScanReturn
rlabel metal1 9385 867 9385 892 7 Vdd!
rlabel metal1 9385 153 9385 163 7 nReset
rlabel metal1 9385 176 9385 186 7 Test
rlabel metal1 9385 199 9385 209 7 Clock
rlabel metal1 9385 223 9385 247 7 GND!
rlabel metal2 2234 0 2246 0 1 Rs2[1]
rlabel metal2 122 1075 134 1075 5 Rw[0]
rlabel metal2 866 0 878 0 1 Rs1[0]
rlabel metal2 1330 3969 1342 3969 5 We
rlabel metal2 1280 3969 1292 3969 5 In[2]
rlabel metal2 1256 3969 1268 3969 5 In[1]
rlabel metal2 1232 3969 1244 3969 5 In[0]
rlabel metal2 1736 2844 1748 2844 1 Out[0]
rlabel metal2 1640 3866 1652 3866 5 In[0]
rlabel metal2 1664 3866 1676 3866 5 In[1]
rlabel metal2 1688 3866 1700 3866 5 In[2]
rlabel metal2 1544 3798 1556 3798 5 In[2]
rlabel metal2 1520 3798 1532 3798 5 In[1]
rlabel metal2 1496 3798 1508 3798 5 In[0]
rlabel metal2 1592 2844 1604 2844 1 Out[0]
rlabel metal2 2336 2844 2348 2844 1 Out[1]
rlabel metal2 2576 2844 2588 2844 1 Out[1]
rlabel metal2 3176 2844 3188 2844 1 Out[2]
rlabel metal2 3416 2844 3428 2844 1 Out[2]
rlabel metal2 3968 2844 3980 2844 1 Out[3]
rlabel metal2 4184 2844 4196 2844 1 Out[3]
rlabel metal2 4784 2844 4796 2844 1 Out[4]
rlabel metal2 5024 2844 5036 2844 1 Out[4]
rlabel metal2 5576 2844 5588 2844 1 Out[5]
rlabel metal2 5792 2844 5804 2844 1 Out[5]
rlabel metal2 6347 2861 6359 2861 1 Out[6]
rlabel metal2 6560 2844 6572 2844 1 Out[6]
rlabel metal2 7160 2844 7172 2844 1 Out[7]
rlabel metal2 7400 2844 7412 2844 1 Out[7]
<< end >>
