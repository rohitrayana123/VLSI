magic
tech c035u
timestamp 1394121372
<< metal1 >>
rect 0 1021 73 1031
rect 88 1021 1225 1031
rect 1239 1021 2377 1031
rect 2392 1021 3529 1031
rect 3543 1021 4681 1031
rect 4695 1021 5833 1031
rect 5847 1021 6984 1031
rect 6999 1021 8137 1031
rect 664 984 793 994
rect 807 984 1009 994
rect 1814 971 1945 981
rect 1959 971 2161 981
rect 2966 971 3097 981
rect 3111 971 3313 981
rect 4118 971 4249 981
rect 4263 971 4465 981
rect 5270 971 5401 981
rect 5415 971 5617 981
rect 6422 971 6553 981
rect 6567 971 6769 981
rect 7574 971 7705 981
rect 7719 971 7921 981
rect 8726 971 8857 981
rect 8871 971 9073 981
rect 0 928 50 938
rect 9266 928 9385 938
rect 0 905 50 915
rect 9266 905 9385 915
rect 0 867 50 892
rect 9266 867 9385 892
rect 0 222 50 247
rect 9266 222 9385 247
rect 0 199 50 209
rect 9266 199 9385 209
rect 0 176 50 186
rect 9266 176 9385 186
rect 0 153 50 163
rect 9266 153 9385 163
rect 0 60 936 70
rect 951 60 2088 70
rect 2103 60 3240 70
rect 3255 60 4393 70
rect 4408 60 5543 70
rect 5561 60 6695 70
rect 6713 60 7847 70
rect 7865 60 9001 70
rect 9015 60 9385 70
rect 0 25 1153 35
rect 1167 25 2305 35
rect 2319 25 3457 35
rect 3471 25 4609 35
rect 4624 25 5760 35
rect 5778 25 6912 35
rect 6930 25 8064 35
rect 8082 25 9217 35
rect 9231 25 9385 35
<< m2contact >>
rect 73 1018 88 1034
rect 1225 1020 1239 1034
rect 2377 1020 2392 1034
rect 3529 1020 3543 1034
rect 4681 1020 4695 1034
rect 5833 1020 5847 1034
rect 6984 1019 6999 1033
rect 8137 1020 8152 1035
rect 649 983 664 997
rect 793 982 807 996
rect 1009 981 1023 995
rect 1800 969 1814 983
rect 1945 968 1959 982
rect 2161 969 2175 983
rect 2952 969 2966 983
rect 3097 968 3111 982
rect 3313 969 3327 983
rect 4104 969 4118 983
rect 4249 968 4263 982
rect 4465 969 4479 983
rect 5256 969 5270 983
rect 5401 968 5415 982
rect 5617 969 5631 983
rect 6408 969 6422 983
rect 6553 968 6567 982
rect 6769 969 6783 983
rect 7560 969 7574 983
rect 7705 968 7719 982
rect 7921 969 7935 983
rect 8712 969 8726 983
rect 8857 968 8871 982
rect 9073 969 9087 983
rect 936 58 951 72
rect 2088 58 2103 72
rect 3240 58 3255 72
rect 4393 58 4408 73
rect 5543 58 5561 73
rect 6695 58 6713 73
rect 7847 58 7865 73
rect 9001 57 9015 72
rect 1153 24 1167 38
rect 2305 24 2319 38
rect 3457 24 3471 38
rect 4609 23 4624 38
rect 5760 20 5778 35
rect 6912 20 6930 35
rect 8064 20 8082 35
rect 9217 23 9231 38
<< metal2 >>
rect 74 945 86 1018
rect 122 945 134 1075
rect 650 945 662 983
rect 794 945 806 982
rect 866 945 878 1075
rect 1010 945 1022 981
rect 1082 945 1094 1075
rect 1226 945 1238 1020
rect 1274 945 1286 1075
rect 1802 945 1814 969
rect 1946 945 1958 968
rect 2018 945 2030 1075
rect 2162 945 2174 969
rect 2234 945 2246 1075
rect 2378 945 2390 1020
rect 2426 945 2438 1075
rect 2954 945 2966 969
rect 3098 945 3110 968
rect 3170 945 3182 1075
rect 3314 945 3326 969
rect 3386 945 3398 1075
rect 3530 945 3542 1020
rect 3578 945 3590 1075
rect 4106 945 4118 969
rect 4250 945 4262 968
rect 4322 945 4334 1075
rect 4466 945 4478 969
rect 4538 945 4550 1075
rect 4682 945 4694 1020
rect 4730 945 4742 1075
rect 5258 945 5270 969
rect 5402 945 5414 968
rect 5474 945 5486 1075
rect 5618 945 5630 969
rect 5690 945 5702 1075
rect 5834 945 5846 1020
rect 5882 945 5894 1075
rect 6410 945 6422 969
rect 6554 945 6566 968
rect 6626 945 6638 1075
rect 6770 945 6782 969
rect 6842 945 6854 1075
rect 6986 945 6998 1019
rect 7034 945 7046 1075
rect 7562 945 7574 969
rect 7706 945 7718 968
rect 7778 945 7790 1075
rect 7922 945 7934 969
rect 7994 945 8006 1075
rect 8138 945 8150 1020
rect 8186 945 8198 1075
rect 8714 945 8726 969
rect 8858 945 8870 968
rect 8930 945 8942 1075
rect 9074 945 9086 969
rect 9146 945 9158 1075
rect 122 0 134 146
rect 866 0 878 146
rect 938 72 950 146
rect 1082 0 1094 146
rect 1154 38 1166 146
rect 1274 0 1286 146
rect 2018 0 2030 146
rect 2090 72 2102 146
rect 2234 0 2246 146
rect 2306 38 2318 146
rect 2426 0 2438 146
rect 3170 0 3182 146
rect 3242 72 3254 146
rect 3386 0 3398 146
rect 3458 38 3470 146
rect 3578 0 3590 146
rect 4322 0 4334 146
rect 4394 73 4406 146
rect 4538 0 4550 146
rect 4610 38 4622 146
rect 4730 0 4742 146
rect 5474 0 5486 146
rect 5546 73 5558 146
rect 5690 0 5702 146
rect 5762 35 5774 146
rect 5882 0 5894 146
rect 6626 0 6638 146
rect 6698 73 6710 146
rect 6842 0 6854 146
rect 6914 35 6926 146
rect 7034 0 7046 146
rect 7778 0 7790 146
rect 7850 73 7862 146
rect 7994 0 8006 146
rect 8066 35 8078 146
rect 8186 0 8198 146
rect 8930 0 8942 146
rect 9002 72 9014 146
rect 9146 0 9158 146
rect 9218 38 9230 146
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 50 0 1 146
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 770 0 1 146
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 986 0 1 146
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 1202 0 1 146
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 1922 0 1 146
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 2138 0 1 146
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 2354 0 1 146
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 3074 0 1 146
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 3290 0 1 146
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 3506 0 1 146
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 4226 0 1 146
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 4442 0 1 146
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 4658 0 1 146
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 5378 0 1 146
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 5594 0 1 146
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 5810 0 1 146
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 6530 0 1 146
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 6746 0 1 146
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 6962 0 1 146
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 7682 0 1 146
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 7898 0 1 146
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 8114 0 1 146
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 8834 0 1 146
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 9050 0 1 146
box 0 0 216 799
<< labels >>
rlabel metal1 0 1021 0 1031 1 WData
rlabel metal1 0 60 0 70 3 Rd1
rlabel metal1 0 25 0 35 3 Rd2
rlabel metal1 0 928 0 938 3 ScanReturn
rlabel metal1 0 905 0 915 3 SDI
rlabel metal1 0 153 0 163 3 nReset
rlabel metal1 0 176 0 186 3 Test
rlabel metal1 0 199 0 209 3 Clock
rlabel metal1 0 222 0 247 3 GND!
rlabel metal1 0 867 0 892 3 Vdd!
rlabel metal2 5474 1075 5486 1075 5 Rs1[4]
rlabel metal2 4730 1075 4742 1075 5 Rw[4]
rlabel metal2 4538 1075 4550 1075 5 Rs2[3]
rlabel metal2 4322 1075 4334 1075 5 Rs1[3]
rlabel metal2 3578 1075 3590 1075 5 Rw[3]
rlabel metal2 3386 1075 3398 1075 5 Rs2[2]
rlabel metal2 3170 1075 3182 1075 5 Rs1[2]
rlabel metal2 2426 1075 2438 1075 5 Rw[2]
rlabel metal2 2234 1075 2246 1075 5 Rs2[1]
rlabel metal2 2018 1075 2030 1075 5 Rs1[1]
rlabel metal2 1274 1075 1286 1075 5 Rw[1]
rlabel metal2 1082 1075 1094 1075 5 Rs2[0]
rlabel metal2 866 1075 878 1075 5 Rs1[0]
rlabel metal2 122 0 134 0 1 Rw[0]
rlabel metal2 1082 0 1094 0 5 Rs2[0]
rlabel metal2 1274 0 1286 0 5 Rw[1]
rlabel metal2 2018 0 2030 0 5 Rs1[1]
rlabel metal2 3170 0 3182 0 5 Rs1[2]
rlabel metal2 3578 0 3590 0 5 Rw[3]
rlabel metal2 3386 0 3398 0 5 Rs2[2]
rlabel metal2 4322 0 4334 0 5 Rs1[3]
rlabel metal2 4730 0 4742 0 5 Rw[4]
rlabel metal2 4538 0 4550 0 5 Rs2[3]
rlabel metal2 5474 0 5486 0 5 Rs1[4]
rlabel metal2 2426 0 2438 0 1 Rw[2]
rlabel metal2 5690 0 5702 0 1 Rs2[4]
rlabel metal2 7778 0 7790 0 5 Rs1[6]
rlabel metal2 9146 0 9158 0 5 Rs2[7]
rlabel metal2 8930 0 8942 0 5 Rs1[7]
rlabel metal2 8186 0 8198 0 5 Rw[7]
rlabel metal2 7994 0 8006 0 5 Rs2[6]
rlabel metal2 7034 0 7046 0 5 Rw[6]
rlabel metal2 6842 0 6854 0 5 Rs2[5]
rlabel metal2 6626 0 6638 0 5 Rs1[5]
rlabel metal2 5882 0 5894 0 5 Rw[5]
rlabel metal2 5690 1075 5702 1075 5 Rs2[4]
rlabel metal2 5882 1075 5894 1075 5 Rw[5]
rlabel metal2 6626 1075 6638 1075 5 Rs1[5]
rlabel metal2 6842 1075 6854 1075 5 Rs2[5]
rlabel metal2 7034 1075 7046 1075 5 Rw[6]
rlabel metal2 7778 1075 7790 1075 5 Rs1[6]
rlabel metal2 7994 1075 8006 1075 5 Rs2[6]
rlabel metal2 8930 1075 8942 1075 5 Rs1[7]
rlabel metal2 9146 1075 9158 1075 5 Rs2[7]
rlabel metal2 8186 1075 8198 1075 5 Rw[7]
rlabel metal1 9385 25 9385 35 7 Rd2
rlabel metal1 9385 60 9385 70 7 Rd1
rlabel metal1 9385 905 9385 915 7 Scan
rlabel metal1 9385 928 9385 938 7 ScanReturn
rlabel metal1 9385 867 9385 892 7 Vdd!
rlabel metal1 9385 153 9385 163 7 nReset
rlabel metal1 9385 176 9385 186 7 Test
rlabel metal1 9385 199 9385 209 7 Clock
rlabel metal1 9385 223 9385 247 7 GND!
rlabel metal2 2234 0 2246 0 1 Rs2[1]
rlabel metal2 122 1075 134 1075 5 Rw[0]
rlabel metal2 866 0 878 0 1 Rs1[0]
<< end >>
