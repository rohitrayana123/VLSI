magic
tech c035u
timestamp 1394133196
<< metal1 >>
rect 5161 16721 5195 16731
rect 5209 16721 5243 16731
rect 5257 16721 5291 16731
rect 5305 16721 5603 16731
rect 5617 16721 5651 16731
rect 5665 16721 5699 16731
rect 5713 16721 6011 16731
rect 6025 16721 6059 16731
rect 6073 16721 6371 16731
rect 2 16563 12 16573
rect 2 16541 12 16551
rect 6972 15722 6982 15732
rect 2 15521 12 15531
rect 2 15499 12 15509
rect 6972 14680 6982 14690
rect 2 14479 12 14489
rect 2 14457 12 14467
rect 6972 13638 6982 13648
rect 2 13437 12 13447
rect 2 13415 12 13425
rect 6972 12596 6982 12606
rect 2 12395 12 12405
rect 2 12373 12 12383
rect 6972 11554 6982 11564
rect 2 11353 12 11363
rect 2 11331 12 11341
rect 6972 10512 6982 10522
rect 2 10311 12 10321
rect 2 10289 12 10299
rect 6972 9470 6982 9480
rect 2 9269 12 9279
rect 2 9247 12 9257
rect 6972 8428 6982 8438
rect 2 8227 12 8237
rect 2 8205 12 8215
rect 6972 7386 6982 7396
rect 2 7185 12 7195
rect 2 7163 12 7173
rect 6972 6344 6982 6354
rect 2 6143 12 6153
rect 2 6121 12 6131
rect 6972 5302 6982 5312
rect 2 5101 12 5111
rect 2 5079 12 5089
rect 6972 4260 6982 4270
rect 2 4059 12 4069
rect 2 4037 12 4047
rect 6972 3218 6982 3228
rect 2 3017 12 3027
rect 2 2995 12 3005
rect 6972 2176 6982 2186
rect 2 1975 12 1985
rect 2 1953 12 1963
rect 6972 1134 6982 1144
rect 2 933 12 943
rect 2 911 12 921
rect 6972 92 6982 102
rect 14 24 947 34
rect 961 24 3611 34
rect 3625 24 3659 34
rect 3673 24 3707 34
rect 3721 24 3755 34
rect 3769 24 4067 34
rect 4081 24 4115 34
rect 4129 24 4163 34
rect 4177 24 4475 34
rect 4489 24 4523 34
rect 4537 24 4907 34
rect 481 2 659 12
<< m2contact >>
rect 5147 16719 5161 16733
rect 5195 16719 5209 16733
rect 5243 16719 5257 16733
rect 5291 16719 5305 16733
rect 5603 16719 5617 16733
rect 5651 16719 5665 16733
rect 5699 16719 5713 16733
rect 6011 16719 6025 16733
rect 6059 16719 6073 16733
rect 6371 16719 6385 16733
rect 0 24 14 38
rect 947 22 961 36
rect 3611 22 3625 36
rect 3659 22 3673 36
rect 3707 22 3721 36
rect 3755 22 3769 36
rect 4067 22 4081 36
rect 4115 22 4129 36
rect 4163 22 4177 36
rect 4475 22 4489 36
rect 4523 22 4537 36
rect 4907 22 4921 36
rect 467 0 481 14
rect 659 0 673 14
<< metal2 >>
rect 36 16713 48 16785
rect 300 16713 312 16785
rect 468 16713 480 16785
rect 636 16713 648 16785
rect 660 16713 672 16785
rect 732 16713 744 16785
rect 948 16713 960 16785
rect 1092 16713 1104 16785
rect 1428 16713 1440 16785
rect 1788 16713 1800 16785
rect 2196 16713 2208 16785
rect 2532 16713 2544 16785
rect 2844 16713 2856 16785
rect 3180 16713 3192 16785
rect 3300 16713 3312 16785
rect 3348 16713 3360 16785
rect 3516 16713 3528 16785
rect 5076 16713 5088 16785
rect 5101 16713 5113 16785
rect 5148 16713 5160 16719
rect 5196 16713 5208 16719
rect 5244 16713 5256 16719
rect 5292 16713 5304 16719
rect 5532 16713 5544 16785
rect 5700 16733 5712 16785
rect 5604 16713 5616 16719
rect 5652 16713 5664 16719
rect 5700 16713 5712 16719
rect 5940 16713 5952 16785
rect 6012 16713 6024 16719
rect 6060 16713 6072 16719
rect 6300 16713 6312 16785
rect 6372 16713 6384 16719
rect 6660 16713 6672 16785
rect 6828 16713 6840 16785
rect 468 14 480 41
rect 660 14 672 41
rect 948 36 960 41
rect 3612 36 3624 41
rect 3660 36 3672 41
rect 3708 36 3720 41
rect 3756 36 3768 41
rect 4068 36 4080 41
rect 4116 36 4128 41
rect 4164 36 4176 41
rect 4476 36 4488 41
rect 4524 36 4536 41
rect 4908 36 4920 41
use ALUSlice ALUSlice_15
timestamp 1394128665
transform 1 0 12 0 1 15671
box 0 0 6768 1042
use LLIcell_U LLIcell_U_7
timestamp 1393855556
transform 1 0 6780 0 1 15671
box 0 0 192 1042
use ALUSlice ALUSlice_14
timestamp 1394128665
transform 1 0 12 0 1 14629
box 0 0 6768 1042
use LLIcell_U LLIcell_U_6
timestamp 1393855556
transform 1 0 6780 0 1 14629
box 0 0 192 1042
use ALUSlice ALUSlice_13
timestamp 1394128665
transform 1 0 12 0 1 13587
box 0 0 6768 1042
use LLIcell_U LLIcell_U_5
timestamp 1393855556
transform 1 0 6780 0 1 13587
box 0 0 192 1042
use ALUSlice ALUSlice_12
timestamp 1394128665
transform 1 0 12 0 1 12545
box 0 0 6768 1042
use LLIcell_U LLIcell_U_4
timestamp 1393855556
transform 1 0 6780 0 1 12545
box 0 0 192 1042
use ALUSlice ALUSlice_11
timestamp 1394128665
transform 1 0 12 0 1 11503
box 0 0 6768 1042
use LLIcell_U LLIcell_U_3
timestamp 1393855556
transform 1 0 6780 0 1 11503
box 0 0 192 1042
use ALUSlice ALUSlice_10
timestamp 1394128665
transform 1 0 12 0 1 10461
box 0 0 6768 1042
use LLIcell_U LLIcell_U_2
timestamp 1393855556
transform 1 0 6780 0 1 10461
box 0 0 192 1042
use ALUSlice ALUSlice_9
timestamp 1394128665
transform 1 0 12 0 1 9419
box 0 0 6768 1042
use LLIcell_U LLIcell_U_1
timestamp 1393855556
transform 1 0 6780 0 1 9419
box 0 0 192 1042
use ALUSlice ALUSlice_8
timestamp 1394128665
transform 1 0 12 0 1 8377
box 0 0 6768 1042
use LLIcell_U LLIcell_U_0
timestamp 1393855556
transform 1 0 6780 0 1 8377
box 0 0 192 1042
use ALUSlice ALUSlice_7
timestamp 1394128665
transform 1 0 12 0 1 7335
box 0 0 6768 1042
use LLIcell_L LLIcell_L_3
timestamp 1393855517
transform 1 0 6780 0 1 7335
box 0 0 192 1042
use ALUSlice ALUSlice_6
timestamp 1394128665
transform 1 0 12 0 1 6293
box 0 0 6768 1042
use LLIcell_L LLIcell_L_7
timestamp 1393855517
transform 1 0 6780 0 1 6293
box 0 0 192 1042
use ALUSlice ALUSlice_5
timestamp 1394128665
transform 1 0 12 0 1 5251
box 0 0 6768 1042
use LLIcell_L LLIcell_L_6
timestamp 1393855517
transform 1 0 6780 0 1 5251
box 0 0 192 1042
use ALUSlice ALUSlice_4
timestamp 1394128665
transform 1 0 12 0 1 4209
box 0 0 6768 1042
use LLIcell_L LLIcell_L_5
timestamp 1393855517
transform 1 0 6780 0 1 4209
box 0 0 192 1042
use ALUSlice ALUSlice_3
timestamp 1394128665
transform 1 0 12 0 1 3167
box 0 0 6768 1042
use LLIcell_L LLIcell_L_4
timestamp 1393855517
transform 1 0 6780 0 1 3167
box 0 0 192 1042
use ALUSlice ALUSlice_2
timestamp 1394128665
transform 1 0 12 0 1 2125
box 0 0 6768 1042
use LLIcell_L LLIcell_L_2
timestamp 1393855517
transform 1 0 6780 0 1 2125
box 0 0 192 1042
use ALUSlice ALUSlice_1
timestamp 1394128665
transform 1 0 12 0 1 1083
box 0 0 6768 1042
use LLIcell_L LLIcell_L_1
timestamp 1393855517
transform 1 0 6780 0 1 1083
box 0 0 192 1042
use ALUSlice ALUSlice_0
timestamp 1394128665
transform 1 0 12 0 1 41
box 0 0 6768 1042
use LLIcell_L LLIcell_L_0
timestamp 1393855517
transform 1 0 6780 0 1 41
box 0 0 192 1042
<< labels >>
rlabel metal1 2 16563 2 16573 3 B[15]
rlabel metal1 2 16541 2 16551 3 A[15]
rlabel metal1 2 15521 2 15531 3 B[14]
rlabel metal1 2 15499 2 15509 3 A[14]
rlabel metal1 2 14457 2 14467 3 A[13]
rlabel metal1 2 14479 2 14489 3 B[13]
rlabel metal1 2 13415 2 13425 3 A[12]
rlabel metal1 2 13437 2 13447 3 B[12]
rlabel metal1 2 12373 2 12383 3 A[11]
rlabel metal1 2 12395 2 12405 3 B[11]
rlabel metal1 2 11331 2 11341 3 A[10]
rlabel metal1 2 11353 2 11363 3 B[10]
rlabel metal1 2 10289 2 10299 3 A[9]
rlabel metal1 2 10311 2 10321 3 B[9]
rlabel metal1 2 9247 2 9257 3 A[8]
rlabel metal1 2 9269 2 9279 3 B[8]
rlabel metal1 2 8205 2 8215 3 A[7]
rlabel metal1 2 8227 2 8237 3 B[7]
rlabel metal1 2 7163 2 7173 3 A[6]
rlabel metal1 2 7185 2 7195 3 B[6]
rlabel metal1 2 6143 2 6153 3 B[5]
rlabel metal1 2 6121 2 6131 3 A[5]
rlabel metal1 2 5079 2 5089 3 A[4]
rlabel metal1 2 5101 2 5111 3 B[4]
rlabel metal1 2 4037 2 4047 3 A[3]
rlabel metal1 2 4059 2 4069 3 B[3]
rlabel metal1 2 3017 2 3027 3 B[2]
rlabel metal1 2 2995 2 3005 3 A[2]
rlabel metal1 2 1975 2 1984 3 B[1]
rlabel metal1 2 1953 2 1963 3 A[1]
rlabel metal1 2 933 2 943 3 B[0]
rlabel metal1 2 911 2 921 3 A[0]
rlabel metal1 6982 92 6982 102 7 ALUOut[0]
rlabel metal1 6982 1134 6982 1144 7 ALUOut[1]
rlabel metal1 6982 2176 6982 2186 7 ALUOut[2]
rlabel metal1 6982 3218 6982 3228 7 ALUOut[3]
rlabel metal1 6982 4260 6982 4270 7 ALUOut[4]
rlabel metal1 6982 5302 6982 5312 7 ALUOut[5]
rlabel metal1 6982 6344 6982 6354 7 ALUOut[6]
rlabel metal1 6982 7386 6982 7396 7 ALUOut[7]
rlabel metal1 6982 8428 6982 8438 7 ALUOut[8]
rlabel metal1 6982 9470 6982 9480 7 ALUOut[9]
rlabel metal1 6982 10512 6982 10522 7 ALUOut[10]
rlabel metal1 6982 11554 6982 11564 7 ALUOut[11]
rlabel metal1 6982 12596 6982 12606 7 ALUOut[12]
rlabel metal1 6982 13638 6982 13648 7 ALUOut[13]
rlabel metal1 6982 14680 6982 14690 7 ALUOut[14]
rlabel metal1 6982 15722 6982 15732 7 ALUOut[15]
rlabel metal2 636 16785 648 16785 5 CIn_Slice
rlabel metal2 3516 16785 3528 16785 5 ShL
rlabel metal2 5101 16785 5113 16785 5 ShR
rlabel metal2 6660 16785 6672 16785 5 ShOut
rlabel metal2 5076 16785 5088 16785 5 Sh8
rlabel metal2 5532 16785 5544 16785 5 Sh4
rlabel metal2 5940 16785 5952 16785 5 Sh2
rlabel metal2 6300 16785 6312 16785 5 Sh1
rlabel metal2 1092 16785 1104 16785 5 FAOut
rlabel metal2 948 16785 960 16785 5 nZ
rlabel metal2 300 16785 312 16785 5 SUB
rlabel metal2 1428 16785 1440 16785 5 AND
rlabel metal2 1788 16785 1800 16785 5 OR
rlabel metal2 2196 16785 2208 16785 5 XOR
rlabel metal2 2532 16785 2544 16785 5 NOT
rlabel metal2 2844 16785 2856 16785 5 NAND
rlabel metal2 3180 16785 3192 16785 5 NOR
rlabel metal2 3348 16785 3360 16785 5 ShB
rlabel metal2 660 16785 672 16785 5 COut
rlabel metal2 732 16785 744 16785 5 Sum
rlabel metal2 468 16785 480 16785 5 CIn
rlabel metal2 3300 16785 3312 16785 5 A
rlabel metal2 36 16785 48 16785 5 ZeroA
rlabel metal2 6828 16785 6840 16785 5 LLI
rlabel metal2 5700 16785 5712 16785 5 ShSignIn
<< end >>
