magic
tech c035u
timestamp 1396390011
<< nwell >>
rect 0 513 192 911
<< pwell >>
rect 0 112 192 513
<< pohmic >>
rect 0 188 6 198
rect 186 188 192 198
<< nohmic >>
rect 0 848 6 858
rect 186 848 192 858
<< psubstratetap >>
rect 6 188 186 204
<< nsubstratetap >>
rect 6 842 186 858
<< metal1 >>
rect 0 1094 192 1104
rect 0 894 192 904
rect 0 871 192 881
rect 0 842 6 858
rect 186 842 192 858
rect 0 833 192 842
rect 0 204 192 213
rect 0 188 6 204
rect 186 188 192 204
rect 0 165 192 175
rect 0 142 192 152
rect 0 119 192 129
rect 0 97 192 107
rect 0 29 192 39
<< metal2 >>
rect 48 0 60 1111
<< labels >>
rlabel metal1 0 833 0 858 1 Vdd!
rlabel metal1 0 871 0 881 1 Scan
rlabel metal1 0 894 0 904 1 ScanReturn
rlabel metal1 192 894 192 904 7 ScanReturn
rlabel metal1 0 97 0 107 3 ALUOut
rlabel metal1 192 97 192 107 7 ALUOut
rlabel metal1 192 188 192 213 7 GND!
rlabel metal1 192 165 192 175 7 Clock
rlabel metal1 192 142 192 152 7 Test
rlabel metal1 192 119 192 129 7 nReset
rlabel metal1 0 188 0 213 1 GND!
rlabel metal1 0 165 0 175 1 Clock
rlabel metal1 0 142 0 152 1 Test
rlabel metal1 0 119 0 129 1 nReset
rlabel metal1 192 833 192 858 7 Vdd!
rlabel metal1 192 871 192 881 7 Scan
rlabel metal1 0 29 0 39 3 SysBus
rlabel metal1 192 29 192 39 7 SysBus
rlabel metal2 48 1111 60 1111 5 LLI
rlabel metal1 0 1094 0 1104 3 ALUOut
rlabel metal1 192 1094 192 1104 7 ALUOut
rlabel metal2 48 0 60 0 1 LLI
<< end >>
