magic
tech c035u
timestamp 1394615469
<< metal1 >>
rect 0 1234 10 1919
rect 120 1258 130 1919
rect 240 1282 250 1919
rect 360 1306 370 1919
rect 480 1330 490 1919
rect 6120 1906 6130 1919
rect 1248 1896 6130 1906
rect 1248 1573 1258 1896
rect 6456 1906 6466 1919
rect 6576 1906 6586 1919
rect 6157 1896 6466 1906
rect 6480 1896 6586 1906
rect 1560 1872 6335 1882
rect 1560 1621 1570 1872
rect 6480 1882 6490 1896
rect 6360 1872 6490 1882
rect 6360 1858 6370 1872
rect 1800 1848 6370 1858
rect 1800 1621 1810 1848
rect 1920 1824 6143 1834
rect 1920 1621 1930 1824
rect 4261 1752 4295 1762
rect 4333 1752 4391 1762
rect 3565 1728 3623 1738
rect 3805 1728 3863 1738
rect 4237 1728 4511 1738
rect 3421 1704 3922 1714
rect 2845 1680 2903 1690
rect 3301 1680 3887 1690
rect 3912 1690 3922 1704
rect 4045 1704 4079 1714
rect 4117 1704 4607 1714
rect 3912 1680 4487 1690
rect 4549 1680 4703 1690
rect 2701 1656 2999 1666
rect 3061 1656 3143 1666
rect 3181 1656 4775 1666
rect 2389 1632 2447 1642
rect 2485 1632 2519 1642
rect 2581 1632 4679 1642
rect 4717 1632 4799 1642
rect 4909 1632 4943 1642
rect 5005 1632 5039 1642
rect 1669 1608 1703 1618
rect 2029 1608 2183 1618
rect 2245 1608 3119 1618
rect 3157 1608 4415 1618
rect 4429 1608 4847 1618
rect 4885 1608 5146 1618
rect 1477 1584 4583 1594
rect 4621 1584 5111 1594
rect 5136 1594 5146 1608
rect 5136 1584 5231 1594
rect 1453 1560 4055 1570
rect 4093 1560 4463 1570
rect 4525 1560 4655 1570
rect 4669 1560 4727 1570
rect 4741 1560 5375 1570
rect 1165 1536 1199 1546
rect 1237 1536 1295 1546
rect 1357 1536 4439 1546
rect 4453 1536 4631 1546
rect 4645 1536 5063 1546
rect 5077 1536 5447 1546
rect 1141 1512 1319 1522
rect 1333 1512 2975 1522
rect 3013 1512 4271 1522
rect 4309 1512 5183 1522
rect 5197 1512 5255 1522
rect 5269 1512 5351 1522
rect 5389 1512 5567 1522
rect 1069 1488 2879 1498
rect 2917 1488 3071 1498
rect 3085 1488 5639 1498
rect 901 1464 935 1474
rect 1021 1464 5015 1474
rect 5053 1464 5591 1474
rect 5605 1464 5783 1474
rect 829 1440 2159 1450
rect 2197 1440 4367 1450
rect 4405 1440 5927 1450
rect 805 1416 1271 1426
rect 1309 1416 1535 1426
rect 1549 1416 1775 1426
rect 1789 1416 1895 1426
rect 1909 1416 3839 1426
rect 3877 1416 5711 1426
rect 5725 1416 6023 1426
rect 733 1392 1031 1402
rect 1045 1392 5543 1402
rect 5581 1392 5759 1402
rect 5797 1392 6095 1402
rect 685 1368 1175 1378
rect 1213 1368 6178 1378
rect 661 1344 4919 1354
rect 4957 1344 6143 1354
rect 6168 1354 6178 1368
rect 6168 1344 6191 1354
rect 480 1320 911 1330
rect 949 1320 2423 1330
rect 2461 1320 3527 1330
rect 3541 1320 3647 1330
rect 3661 1320 3767 1330
rect 3781 1320 4007 1330
rect 4021 1320 5423 1330
rect 5461 1320 6311 1330
rect 360 1296 1679 1306
rect 1717 1296 3599 1306
rect 3637 1296 5903 1306
rect 5941 1296 6167 1306
rect 6205 1296 6263 1306
rect 6277 1296 6335 1306
rect 240 1272 4823 1282
rect 4837 1272 5519 1282
rect 5533 1272 6071 1282
rect 6109 1272 6287 1282
rect 6325 1272 6407 1282
rect 120 1248 2591 1258
rect 2605 1248 2711 1258
rect 2725 1248 4127 1258
rect 4141 1248 4751 1258
rect 4789 1248 5207 1258
rect 5245 1248 5495 1258
rect 5509 1248 6538 1258
rect 0 1224 2506 1234
rect 2496 1213 2506 1224
rect 2533 1224 4786 1234
rect 2928 1213 2938 1224
rect 4776 1213 4786 1224
rect 4813 1224 6010 1234
rect 6000 1213 6010 1224
rect 6528 1234 6538 1248
rect 6037 1224 6514 1234
rect 6528 1224 6562 1234
rect 6504 1213 6514 1224
rect 6552 1213 6562 1224
rect 1392 322 1402 335
rect 0 312 1402 322
rect 0 -443 10 312
rect 2280 322 2290 335
rect 1429 312 2290 322
rect 4176 322 4186 335
rect 2317 312 4186 322
rect 5376 322 5386 335
rect 6576 322 6586 335
rect 6816 322 6826 335
rect 6936 322 6946 335
rect 4213 312 6946 322
rect 7032 322 7042 335
rect 7344 322 7354 335
rect 6997 312 7354 322
rect 7632 322 7642 335
rect 7381 312 7642 322
rect 7704 322 7714 335
rect 7752 322 7762 335
rect 7669 312 7714 322
rect 7728 312 7762 322
rect 277 288 575 298
rect 613 288 743 298
rect 781 288 2063 298
rect 2101 288 4967 298
rect 4981 288 6623 298
rect 6661 288 7391 298
rect 7429 288 7463 298
rect 7501 288 7583 298
rect 7728 298 7738 312
rect 7621 288 7738 298
rect 24 -422 34 287
rect 192 -398 202 287
rect 264 264 455 274
rect 264 -371 274 264
rect 469 264 1079 274
rect 1117 264 2519 274
rect 2557 264 2639 274
rect 2677 264 3095 274
rect 3109 264 6359 274
rect 6373 264 6911 274
rect 6925 264 7007 274
rect 7021 264 7655 274
rect 432 240 599 250
rect 288 -374 298 239
rect 432 -347 442 240
rect 709 240 767 250
rect 925 240 3311 250
rect 3325 240 4031 250
rect 4069 240 6095 250
rect 6109 240 6239 250
rect 6253 240 6455 250
rect 6469 240 7511 250
rect 7536 240 7607 250
rect 480 -350 490 215
rect 480 -360 634 -350
rect 624 -371 634 -360
rect 288 -384 599 -374
rect 840 -398 850 239
rect 912 216 7223 226
rect 912 -371 922 216
rect 7536 226 7546 240
rect 7261 216 7546 226
rect 1056 192 1103 202
rect 960 -374 970 191
rect 1056 -347 1066 192
rect 1392 192 1415 202
rect 1392 -347 1402 192
rect 1693 192 2855 202
rect 2869 192 6479 202
rect 6493 192 6791 202
rect 6805 192 7127 202
rect 7141 192 7487 202
rect 1488 -350 1498 191
rect 1608 -326 1618 191
rect 1752 168 3455 178
rect 1728 -302 1738 167
rect 1752 -275 1762 168
rect 3493 168 3719 178
rect 3757 168 5087 178
rect 5101 168 5159 178
rect 5173 168 5471 178
rect 5485 168 7175 178
rect 7213 168 7415 178
rect 2053 144 2087 154
rect 2160 144 2303 154
rect 1848 -278 1858 143
rect 1968 -254 1978 143
rect 2112 -230 2122 143
rect 2160 -203 2170 144
rect 2365 144 4343 154
rect 4357 144 4559 154
rect 4573 144 7367 154
rect 2509 120 2663 130
rect 2725 120 2807 130
rect 2821 120 3191 130
rect 3216 120 3239 130
rect 2400 -206 2410 119
rect 2496 96 2543 106
rect 2496 -179 2506 96
rect 3216 106 3226 120
rect 3312 120 3359 130
rect 3144 96 3226 106
rect 2760 -182 2770 95
rect 3144 -179 3154 96
rect 2760 -192 2807 -182
rect 2400 -216 3263 -206
rect 3312 -227 3322 120
rect 3685 120 3743 130
rect 3901 120 5303 130
rect 5341 120 6719 130
rect 6757 120 6959 130
rect 7021 120 7247 130
rect 3480 -227 3490 119
rect 3925 96 4055 106
rect 4141 96 4199 106
rect 4477 96 5855 106
rect 5869 96 7103 106
rect 7117 96 7199 106
rect 4861 72 5279 82
rect 5293 72 6863 82
rect 6901 72 7055 82
rect 2112 -240 3311 -230
rect 3960 -230 3970 71
rect 5269 48 5327 58
rect 5509 48 7007 58
rect 5533 24 6983 34
rect 5845 0 5951 10
rect 5965 0 6671 10
rect 6685 0 6887 10
rect 5989 -24 6743 -14
rect 6349 -48 6647 -38
rect 3960 -240 5327 -230
rect 1968 -264 5351 -254
rect 1848 -288 5687 -278
rect 1728 -312 5303 -302
rect 5365 -312 5962 -302
rect 1608 -336 5927 -326
rect 5952 -326 5962 -312
rect 5952 -336 6383 -326
rect 1488 -360 6778 -350
rect 960 -384 5663 -374
rect 5701 -384 6743 -374
rect 6768 -374 6778 -360
rect 6768 -384 7103 -374
rect 192 -408 730 -398
rect 840 -408 5279 -398
rect 720 -422 730 -408
rect 5341 -408 7271 -398
rect 24 -432 706 -422
rect 720 -432 7522 -422
rect 696 -443 706 -432
rect 7512 -443 7522 -432
<< m2contact >>
rect -1 1919 13 1933
rect 119 1919 133 1933
rect 239 1919 253 1933
rect 359 1919 373 1933
rect 479 1919 493 1933
rect 6119 1919 6133 1933
rect 6455 1919 6469 1933
rect 6575 1919 6589 1933
rect 6143 1895 6157 1909
rect 6335 1871 6349 1885
rect 6143 1823 6157 1837
rect 4247 1751 4261 1765
rect 4295 1751 4309 1765
rect 4319 1751 4333 1765
rect 4391 1751 4405 1765
rect 3551 1727 3565 1741
rect 3623 1727 3637 1741
rect 3791 1727 3805 1741
rect 3863 1727 3877 1741
rect 4223 1727 4237 1741
rect 4511 1727 4525 1741
rect 3407 1703 3421 1717
rect 2831 1679 2845 1693
rect 2903 1679 2917 1693
rect 3287 1679 3301 1693
rect 3887 1679 3901 1693
rect 4031 1703 4045 1717
rect 4079 1703 4093 1717
rect 4103 1703 4117 1717
rect 4607 1703 4621 1717
rect 4487 1679 4501 1693
rect 4535 1679 4549 1693
rect 4703 1679 4717 1693
rect 2687 1655 2701 1669
rect 2999 1655 3013 1669
rect 3047 1655 3061 1669
rect 3143 1655 3157 1669
rect 3167 1655 3181 1669
rect 4775 1655 4789 1669
rect 2375 1631 2389 1645
rect 2447 1631 2461 1645
rect 2471 1631 2485 1645
rect 2519 1631 2533 1645
rect 2567 1631 2581 1645
rect 4679 1631 4693 1645
rect 4703 1631 4717 1645
rect 4799 1631 4813 1645
rect 4895 1631 4909 1645
rect 4943 1631 4957 1645
rect 4991 1631 5005 1645
rect 5039 1631 5053 1645
rect 1559 1607 1573 1621
rect 1655 1607 1669 1621
rect 1703 1607 1717 1621
rect 1799 1607 1813 1621
rect 1919 1607 1933 1621
rect 2015 1607 2029 1621
rect 2183 1607 2197 1621
rect 2231 1607 2245 1621
rect 3119 1607 3133 1621
rect 3143 1607 3157 1621
rect 4415 1607 4429 1621
rect 4847 1607 4861 1621
rect 4871 1607 4885 1621
rect 1463 1583 1477 1597
rect 4583 1583 4597 1597
rect 4607 1583 4621 1597
rect 5111 1583 5125 1597
rect 5231 1583 5245 1597
rect 1247 1559 1261 1573
rect 1439 1559 1453 1573
rect 4055 1559 4069 1573
rect 4079 1559 4093 1573
rect 4463 1559 4477 1573
rect 4511 1559 4525 1573
rect 4655 1559 4669 1573
rect 4727 1559 4741 1573
rect 5375 1559 5389 1573
rect 1151 1535 1165 1549
rect 1199 1535 1213 1549
rect 1223 1535 1237 1549
rect 1295 1535 1309 1549
rect 1343 1535 1357 1549
rect 4439 1535 4453 1549
rect 4631 1535 4645 1549
rect 5063 1535 5077 1549
rect 5447 1535 5461 1549
rect 1127 1511 1141 1525
rect 1319 1511 1333 1525
rect 2975 1511 2989 1525
rect 2999 1511 3013 1525
rect 4271 1511 4285 1525
rect 4295 1511 4309 1525
rect 5183 1511 5197 1525
rect 5255 1511 5269 1525
rect 5351 1511 5365 1525
rect 5375 1511 5389 1525
rect 5567 1511 5581 1525
rect 1055 1487 1069 1501
rect 2879 1487 2893 1501
rect 2903 1487 2917 1501
rect 3071 1487 3085 1501
rect 5639 1487 5653 1501
rect 887 1463 901 1477
rect 935 1463 949 1477
rect 1007 1463 1021 1477
rect 5015 1463 5029 1477
rect 5039 1463 5053 1477
rect 5591 1463 5605 1477
rect 5783 1463 5797 1477
rect 815 1439 829 1453
rect 2159 1439 2173 1453
rect 2183 1439 2197 1453
rect 4367 1439 4381 1453
rect 4391 1439 4405 1453
rect 5927 1439 5941 1453
rect 791 1415 805 1429
rect 1271 1415 1285 1429
rect 1295 1415 1309 1429
rect 1535 1415 1549 1429
rect 1775 1415 1789 1429
rect 1895 1415 1909 1429
rect 3839 1415 3853 1429
rect 3863 1415 3877 1429
rect 5711 1415 5725 1429
rect 6023 1415 6037 1429
rect 719 1391 733 1405
rect 1031 1391 1045 1405
rect 5543 1391 5557 1405
rect 5567 1391 5581 1405
rect 5759 1391 5773 1405
rect 5783 1391 5797 1405
rect 6095 1391 6109 1405
rect 671 1367 685 1381
rect 1175 1367 1189 1381
rect 1199 1367 1213 1381
rect 647 1343 661 1357
rect 4919 1343 4933 1357
rect 4943 1343 4957 1357
rect 6143 1343 6157 1357
rect 6191 1343 6205 1357
rect 911 1319 925 1333
rect 935 1319 949 1333
rect 2423 1319 2437 1333
rect 2447 1319 2461 1333
rect 3527 1319 3541 1333
rect 3647 1319 3661 1333
rect 3767 1319 3781 1333
rect 4007 1319 4021 1333
rect 5423 1319 5437 1333
rect 5447 1319 5461 1333
rect 6311 1319 6325 1333
rect 1679 1295 1693 1309
rect 1703 1295 1717 1309
rect 3599 1295 3613 1309
rect 3623 1295 3637 1309
rect 5903 1295 5917 1309
rect 5927 1295 5941 1309
rect 6167 1295 6181 1309
rect 6191 1295 6205 1309
rect 6263 1295 6277 1309
rect 6335 1295 6349 1309
rect 4823 1271 4837 1285
rect 5519 1271 5533 1285
rect 6071 1271 6085 1285
rect 6095 1271 6109 1285
rect 6287 1271 6301 1285
rect 6311 1271 6325 1285
rect 6407 1271 6421 1285
rect 2591 1247 2605 1261
rect 2711 1247 2725 1261
rect 4127 1247 4141 1261
rect 4751 1247 4765 1261
rect 4775 1247 4789 1261
rect 5207 1247 5221 1261
rect 5231 1247 5245 1261
rect 5495 1247 5509 1261
rect 2519 1223 2533 1237
rect 4799 1223 4813 1237
rect 6023 1223 6037 1237
rect 2495 1199 2509 1213
rect 2927 1199 2941 1213
rect 4775 1199 4789 1213
rect 5999 1199 6013 1213
rect 6503 1199 6517 1213
rect 6551 1199 6565 1213
rect 1391 335 1405 349
rect 2279 335 2293 349
rect 4175 335 4189 349
rect 5375 335 5389 349
rect 6575 335 6589 349
rect 6815 335 6829 349
rect 6935 335 6949 349
rect 7031 335 7045 349
rect 7343 335 7357 349
rect 7631 335 7645 349
rect 7703 335 7717 349
rect 7751 335 7765 349
rect 1415 311 1429 325
rect 2303 311 2317 325
rect 4199 311 4213 325
rect 6959 311 6973 325
rect 6983 311 6997 325
rect 7367 311 7381 325
rect 7655 311 7669 325
rect 23 287 37 301
rect 191 287 205 301
rect 263 287 277 301
rect 575 287 589 301
rect 599 287 613 301
rect 743 287 757 301
rect 767 287 781 301
rect 2063 287 2077 301
rect 2087 287 2101 301
rect 4967 287 4981 301
rect 6623 287 6637 301
rect 6647 287 6661 301
rect 7391 287 7405 301
rect 7415 287 7429 301
rect 7463 287 7477 301
rect 7487 287 7501 301
rect 7583 287 7597 301
rect 7607 287 7621 301
rect 455 263 469 277
rect 1079 263 1093 277
rect 1103 263 1117 277
rect 2519 263 2533 277
rect 2543 263 2557 277
rect 2639 263 2653 277
rect 2663 263 2677 277
rect 3095 263 3109 277
rect 6359 263 6373 277
rect 6911 263 6925 277
rect 7007 263 7021 277
rect 7655 263 7669 277
rect 287 239 301 253
rect 263 -385 277 -371
rect 599 239 613 253
rect 695 239 709 253
rect 767 239 781 253
rect 839 239 853 253
rect 911 239 925 253
rect 3311 239 3325 253
rect 4031 239 4045 253
rect 4055 239 4069 253
rect 6095 239 6109 253
rect 6239 239 6253 253
rect 6455 239 6469 253
rect 7511 239 7525 253
rect 479 215 493 229
rect 431 -361 445 -347
rect 599 -385 613 -371
rect 623 -385 637 -371
rect 7223 215 7237 229
rect 7247 215 7261 229
rect 7607 239 7621 253
rect 959 191 973 205
rect 911 -385 925 -371
rect 1103 191 1117 205
rect 1415 191 1429 205
rect 1487 191 1501 205
rect 1607 191 1621 205
rect 1679 191 1693 205
rect 2855 191 2869 205
rect 6479 191 6493 205
rect 6791 191 6805 205
rect 7127 191 7141 205
rect 7487 191 7501 205
rect 1055 -361 1069 -347
rect 1391 -361 1405 -347
rect 1727 167 1741 181
rect 3455 167 3469 181
rect 3479 167 3493 181
rect 3719 167 3733 181
rect 3743 167 3757 181
rect 5087 167 5101 181
rect 5159 167 5173 181
rect 5471 167 5485 181
rect 7175 167 7189 181
rect 7199 167 7213 181
rect 7415 167 7429 181
rect 1847 143 1861 157
rect 1967 143 1981 157
rect 2039 143 2053 157
rect 2087 143 2101 157
rect 2111 143 2125 157
rect 1751 -289 1765 -275
rect 2303 143 2317 157
rect 2351 143 2365 157
rect 4343 143 4357 157
rect 4559 143 4573 157
rect 7367 143 7381 157
rect 2399 119 2413 133
rect 2495 119 2509 133
rect 2663 119 2677 133
rect 2711 119 2725 133
rect 2807 119 2821 133
rect 3191 119 3205 133
rect 2159 -217 2173 -203
rect 2543 95 2557 109
rect 2759 95 2773 109
rect 3239 119 3253 133
rect 2495 -193 2509 -179
rect 2807 -193 2821 -179
rect 3143 -193 3157 -179
rect 3263 -217 3277 -203
rect 3359 119 3373 133
rect 3479 119 3493 133
rect 3671 119 3685 133
rect 3743 119 3757 133
rect 3887 119 3901 133
rect 5303 119 5317 133
rect 5327 119 5341 133
rect 6719 119 6733 133
rect 6743 119 6757 133
rect 6959 119 6973 133
rect 7007 119 7021 133
rect 7247 119 7261 133
rect 3911 95 3925 109
rect 4055 95 4069 109
rect 4127 95 4141 109
rect 4199 95 4213 109
rect 4463 95 4477 109
rect 5855 95 5869 109
rect 7103 95 7117 109
rect 7199 95 7213 109
rect 3959 71 3973 85
rect 4847 71 4861 85
rect 5279 71 5293 85
rect 6863 71 6877 85
rect 6887 71 6901 85
rect 7055 71 7069 85
rect 3311 -241 3325 -227
rect 3479 -241 3493 -227
rect 5255 47 5269 61
rect 5327 47 5341 61
rect 5495 47 5509 61
rect 7007 47 7021 61
rect 5519 23 5533 37
rect 6983 23 6997 37
rect 5831 -1 5845 13
rect 5951 -1 5965 13
rect 6671 -1 6685 13
rect 6887 -1 6901 13
rect 5975 -25 5989 -11
rect 6743 -25 6757 -11
rect 6335 -49 6349 -35
rect 6647 -49 6661 -35
rect 5327 -241 5341 -227
rect 5351 -265 5365 -251
rect 5687 -289 5701 -275
rect 5303 -313 5317 -299
rect 5351 -313 5365 -299
rect 5927 -337 5941 -323
rect 6383 -337 6397 -323
rect 5663 -385 5677 -371
rect 5687 -385 5701 -371
rect 6743 -385 6757 -371
rect 7103 -385 7117 -371
rect 5279 -409 5293 -395
rect 5327 -409 5341 -395
rect 7271 -409 7285 -395
rect -1 -457 13 -443
rect 695 -457 709 -443
rect 7511 -457 7525 -443
<< metal2 >>
rect 0 1933 12 1959
rect 120 1933 132 1959
rect 240 1933 252 1959
rect 360 1933 372 1959
rect 480 1933 492 1959
rect 6120 1933 6132 1959
rect 6144 1837 6156 1895
rect 6336 1885 6348 1959
rect 6456 1933 6468 1959
rect 6576 1933 6588 1959
rect 6960 1800 6972 1963
rect 144 1788 6972 1800
rect 144 1173 156 1788
rect 648 1173 660 1343
rect 672 1173 684 1367
rect 720 1173 732 1391
rect 792 1173 804 1415
rect 816 1173 828 1439
rect 888 1173 900 1463
rect 936 1333 948 1463
rect 912 1173 924 1319
rect 1008 1173 1020 1463
rect 1032 1173 1044 1391
rect 1056 1173 1068 1487
rect 1128 1173 1140 1511
rect 1152 1173 1164 1535
rect 1200 1381 1212 1535
rect 1176 1173 1188 1367
rect 1224 1173 1236 1535
rect 1248 1173 1260 1559
rect 1296 1429 1308 1535
rect 1272 1173 1284 1415
rect 1320 1173 1332 1511
rect 1344 1173 1356 1535
rect 1440 1173 1452 1559
rect 1464 1173 1476 1583
rect 1536 1173 1548 1415
rect 1560 1173 1572 1607
rect 1656 1173 1668 1607
rect 1704 1309 1716 1607
rect 1680 1173 1692 1295
rect 1776 1173 1788 1415
rect 1800 1173 1812 1607
rect 1896 1173 1908 1415
rect 1920 1173 1932 1607
rect 2016 1173 2028 1607
rect 2184 1453 2196 1607
rect 2160 1173 2172 1439
rect 2232 1173 2244 1607
rect 2376 1173 2388 1631
rect 2448 1333 2460 1631
rect 2424 1173 2436 1319
rect 2472 1173 2484 1631
rect 2520 1237 2532 1631
rect 2496 1173 2508 1199
rect 2568 1173 2580 1631
rect 2592 1173 2604 1247
rect 2688 1173 2700 1655
rect 2712 1173 2724 1247
rect 2832 1173 2844 1679
rect 2904 1501 2916 1679
rect 3000 1525 3012 1655
rect 2880 1173 2892 1487
rect 2928 1173 2940 1199
rect 2976 1173 2988 1511
rect 3048 1173 3060 1655
rect 3144 1621 3156 1655
rect 3072 1173 3084 1487
rect 3120 1173 3132 1607
rect 3168 1173 3180 1655
rect 3288 1173 3300 1679
rect 3408 1173 3420 1703
rect 3528 1173 3540 1319
rect 3552 1173 3564 1727
rect 3624 1309 3636 1727
rect 3600 1173 3612 1295
rect 3648 1173 3660 1319
rect 3768 1173 3780 1319
rect 3792 1173 3804 1727
rect 3864 1429 3876 1727
rect 3840 1173 3852 1415
rect 3888 1173 3900 1679
rect 4008 1173 4020 1319
rect 4032 1173 4044 1703
rect 4080 1573 4092 1703
rect 4056 1173 4068 1559
rect 4104 1173 4116 1703
rect 4128 1173 4140 1247
rect 4224 1173 4236 1727
rect 4248 1173 4260 1751
rect 4296 1525 4308 1751
rect 4272 1173 4284 1511
rect 4320 1173 4332 1751
rect 4392 1453 4404 1751
rect 4368 1173 4380 1439
rect 4416 1173 4428 1607
rect 4440 1173 4452 1535
rect 4464 1173 4476 1559
rect 4488 1173 4500 1679
rect 4512 1573 4524 1727
rect 4536 1173 4548 1679
rect 4608 1597 4620 1703
rect 4704 1645 4716 1679
rect 4584 1173 4596 1583
rect 4632 1173 4644 1535
rect 4656 1173 4668 1559
rect 4680 1173 4692 1631
rect 4728 1173 4740 1559
rect 4776 1261 4788 1655
rect 4752 1173 4764 1247
rect 4800 1237 4812 1631
rect 4776 1173 4788 1199
rect 4824 1173 4836 1271
rect 4848 1173 4860 1607
rect 4872 1173 4884 1607
rect 4896 1173 4908 1631
rect 4944 1357 4956 1631
rect 4920 1173 4932 1343
rect 4992 1173 5004 1631
rect 5040 1477 5052 1631
rect 5016 1173 5028 1463
rect 5064 1173 5076 1535
rect 5112 1173 5124 1583
rect 5184 1173 5196 1511
rect 5232 1261 5244 1583
rect 5376 1525 5388 1559
rect 5208 1173 5220 1247
rect 5256 1173 5268 1511
rect 5352 1173 5364 1511
rect 5448 1333 5460 1535
rect 5568 1405 5580 1511
rect 5424 1173 5436 1319
rect 5496 1173 5508 1247
rect 5520 1173 5532 1271
rect 5544 1173 5556 1391
rect 5592 1173 5604 1463
rect 5640 1173 5652 1487
rect 5712 1173 5724 1415
rect 5784 1405 5796 1463
rect 5760 1173 5772 1391
rect 5928 1309 5940 1439
rect 5904 1173 5916 1295
rect 6024 1237 6036 1415
rect 6096 1285 6108 1391
rect 6000 1173 6012 1199
rect 6072 1173 6084 1271
rect 6144 1173 6156 1343
rect 6192 1309 6204 1343
rect 6168 1173 6180 1295
rect 6264 1173 6276 1295
rect 6312 1285 6324 1319
rect 6288 1173 6300 1271
rect 6336 1173 6348 1295
rect 6408 1173 6420 1271
rect 6504 1173 6516 1199
rect 6552 1173 6564 1199
rect 24 301 36 374
rect 192 301 204 374
rect 264 301 276 374
rect 288 253 300 374
rect 456 277 468 374
rect 480 229 492 374
rect 576 301 588 374
rect 600 253 612 287
rect 696 253 708 374
rect 744 301 756 374
rect 768 253 780 287
rect 840 253 852 374
rect 912 253 924 374
rect 960 205 972 374
rect 1080 277 1092 374
rect 1392 349 1404 374
rect 1104 205 1116 263
rect 1416 205 1428 311
rect 1488 205 1500 374
rect 1608 205 1620 374
rect 1680 205 1692 374
rect 1728 181 1740 374
rect 1848 157 1860 374
rect 1968 157 1980 374
rect 2040 157 2052 374
rect 2064 301 2076 374
rect 2088 157 2100 287
rect 2112 157 2124 374
rect 2280 349 2292 374
rect 2304 157 2316 311
rect 2352 157 2364 374
rect 2400 133 2412 374
rect 2496 133 2508 374
rect 2520 277 2532 374
rect 2640 277 2652 374
rect 2544 109 2556 263
rect 2664 133 2676 263
rect 2712 133 2724 374
rect 2760 109 2772 374
rect 2808 133 2820 374
rect 2856 205 2868 374
rect 3096 277 3108 374
rect 3192 133 3204 374
rect 3240 133 3252 374
rect 3312 253 3324 374
rect 3360 133 3372 374
rect 3456 181 3468 374
rect 3480 133 3492 167
rect 3672 133 3684 374
rect 3720 181 3732 374
rect 3744 133 3756 167
rect 3888 133 3900 374
rect 3912 109 3924 374
rect 3960 85 3972 374
rect 4032 253 4044 374
rect 4056 109 4068 239
rect 4128 109 4140 374
rect 4176 349 4188 374
rect 4200 109 4212 311
rect 4344 157 4356 374
rect 4464 109 4476 374
rect 4560 157 4572 374
rect 4848 85 4860 374
rect 4968 301 4980 374
rect 5088 181 5100 374
rect 5160 181 5172 374
rect 5256 61 5268 374
rect 5280 85 5292 374
rect 5304 133 5316 374
rect 5376 349 5388 374
rect 5472 181 5484 374
rect 5328 61 5340 119
rect 5496 61 5508 374
rect 5520 37 5532 374
rect 5832 13 5844 374
rect 5856 109 5868 374
rect 5952 13 5964 374
rect 5976 -11 5988 374
rect 6096 253 6108 374
rect 6240 253 6252 374
rect 6336 -35 6348 374
rect 6360 277 6372 374
rect 6456 253 6468 374
rect 6480 205 6492 374
rect 6576 349 6588 374
rect 6624 301 6636 374
rect 6648 -35 6660 287
rect 6672 13 6684 374
rect 6720 133 6732 374
rect 6792 205 6804 374
rect 6816 349 6828 374
rect 6744 -11 6756 119
rect 6864 85 6876 374
rect 6912 277 6924 374
rect 6936 349 6948 374
rect 6960 325 6972 374
rect 6960 133 6972 311
rect 6888 13 6900 71
rect 6984 37 6996 311
rect 7008 277 7020 374
rect 7032 349 7044 374
rect 7008 61 7020 119
rect 7056 85 7068 374
rect 7104 109 7116 374
rect 7128 205 7140 374
rect 7176 181 7188 374
rect 7224 229 7236 374
rect 7344 349 7356 374
rect 7200 109 7212 167
rect 7248 133 7260 215
rect 7368 157 7380 311
rect 7392 301 7404 374
rect 7464 301 7476 374
rect 7416 181 7428 287
rect 7488 205 7500 287
rect 7512 253 7524 374
rect 7584 301 7596 374
rect 7632 349 7644 374
rect 7704 349 7716 374
rect 7752 349 7764 374
rect 7608 253 7620 287
rect 7656 277 7668 311
rect 0 -488 12 -457
rect 264 -488 276 -385
rect 432 -488 444 -361
rect 600 -488 612 -385
rect 624 -488 636 -385
rect 696 -488 708 -457
rect 912 -488 924 -385
rect 1056 -488 1068 -361
rect 1392 -488 1404 -361
rect 1752 -488 1764 -289
rect 2160 -488 2172 -217
rect 2496 -488 2508 -193
rect 2808 -488 2820 -193
rect 3144 -488 3156 -193
rect 3264 -488 3276 -217
rect 3312 -488 3324 -241
rect 3480 -488 3492 -241
rect 5280 -488 5292 -409
rect 5304 -444 5316 -313
rect 5328 -395 5340 -241
rect 5352 -299 5364 -265
rect 5688 -371 5700 -289
rect 5304 -456 5317 -444
rect 5305 -488 5317 -456
rect 5664 -488 5676 -385
rect 5928 -488 5940 -337
rect 6384 -488 6396 -337
rect 6744 -488 6756 -385
rect 7104 -488 7116 -385
rect 7272 -488 7284 -409
rect 7512 -488 7524 -457
use buffer rm_assigns_buf_N
timestamp 1386236986
transform 1 0 0 0 1 374
box 0 0 120 799
use buffer rm_assigns_buf_OutEn_slice
timestamp 1386236986
transform 1 0 120 0 1 374
box 0 0 120 799
use xor2 g2055
timestamp 1386237344
transform 1 0 240 0 1 374
box 0 0 192 799
use xor2 g2057
timestamp 1386237344
transform 1 0 432 0 1 374
box 0 0 192 799
use nand4 g2056
timestamp 1386234936
transform 1 0 624 0 1 374
box 0 0 144 799
use nand2 g2058
timestamp 1386234792
transform 1 0 768 0 1 374
box 0 0 96 799
use nor2 g2059
timestamp 1386235306
transform 1 0 864 0 1 374
box 0 0 120 799
use nand3 g2060
timestamp 1386234893
transform 1 0 984 0 1 374
box 0 0 120 799
use nand2 g2070
timestamp 1386234792
transform 1 0 1104 0 1 374
box 0 0 96 799
use nand2 g2063
timestamp 1386234792
transform 1 0 1200 0 1 374
box 0 0 96 799
use and2 g2077
timestamp 1386234845
transform 1 0 1296 0 1 374
box 0 0 120 799
use nand2 g2062
timestamp 1386234792
transform 1 0 1416 0 1 374
box 0 0 96 799
use and2 g2064
timestamp 1386234845
transform 1 0 1512 0 1 374
box 0 0 120 799
use nor2 g2061
timestamp 1386235306
transform 1 0 1632 0 1 374
box 0 0 120 799
use and2 g2066
timestamp 1386234845
transform 1 0 1752 0 1 374
box 0 0 120 799
use and2 g2065
timestamp 1386234845
transform 1 0 1872 0 1 374
box 0 0 120 799
use nand2 g2067
timestamp 1386234792
transform 1 0 1992 0 1 374
box 0 0 96 799
use inv g2072
timestamp 1386238110
transform 1 0 2088 0 1 374
box 0 0 120 799
use inv g2088
timestamp 1386238110
transform 1 0 2208 0 1 374
box 0 0 120 799
use nand3 g2068
timestamp 1386234893
transform 1 0 2328 0 1 374
box 0 0 120 799
use nand2 g2086
timestamp 1386234792
transform 1 0 2448 0 1 374
box 0 0 96 799
use nor2 g2079
timestamp 1386235306
transform 1 0 2544 0 1 374
box 0 0 120 799
use nor2 g2083
timestamp 1386235306
transform 1 0 2664 0 1 374
box 0 0 120 799
use nand3 g2087
timestamp 1386234893
transform 1 0 2784 0 1 374
box 0 0 120 799
use inv g2096
timestamp 1386238110
transform 1 0 2904 0 1 374
box 0 0 120 799
use nand3 g2089
timestamp 1386234893
transform 1 0 3024 0 1 374
box 0 0 120 799
use nor2 g2084
timestamp 1386235306
transform 1 0 3144 0 1 374
box 0 0 120 799
use nor2 g2073
timestamp 1386235306
transform 1 0 3264 0 1 374
box 0 0 120 799
use inv g2090
timestamp 1386238110
transform 1 0 3384 0 1 374
box 0 0 120 799
use nor2 g2075
timestamp 1386235306
transform 1 0 3504 0 1 374
box 0 0 120 799
use and2 g2082
timestamp 1386234845
transform 1 0 3624 0 1 374
box 0 0 120 799
use and2 g2080
timestamp 1386234845
transform 1 0 3744 0 1 374
box 0 0 120 799
use nor2 g2076
timestamp 1386235306
transform 1 0 3864 0 1 374
box 0 0 120 799
use nand2 g2081
timestamp 1386234792
transform 1 0 3984 0 1 374
box 0 0 96 799
use nor2 g2078
timestamp 1386235306
transform 1 0 4080 0 1 374
box 0 0 120 799
use nand2 g2098
timestamp 1386234792
transform 1 0 4200 0 1 374
box 0 0 96 799
use nand2 g2071
timestamp 1386234792
transform 1 0 4296 0 1 374
box 0 0 96 799
use nand3 g2091
timestamp 1386234893
transform 1 0 4392 0 1 374
box 0 0 120 799
use nand2 g2074
timestamp 1386234792
transform 1 0 4512 0 1 374
box 0 0 96 799
use nand2 g2095
timestamp 1386234792
transform 1 0 4608 0 1 374
box 0 0 96 799
use nand2 g2097
timestamp 1386234792
transform 1 0 4704 0 1 374
box 0 0 96 799
use nand4 g2069
timestamp 1386234936
transform 1 0 4800 0 1 374
box 0 0 144 799
use nand2 g2092
timestamp 1386234792
transform 1 0 4944 0 1 374
box 0 0 96 799
use nand2 g2094
timestamp 1386234792
transform 1 0 5040 0 1 374
box 0 0 96 799
use nand2 g2099
timestamp 1386234792
transform 1 0 5136 0 1 374
box 0 0 96 799
use nand2 g2100
timestamp 1386234792
transform 1 0 5232 0 1 374
box 0 0 96 799
use and2 g2101
timestamp 1386234845
transform 1 0 5328 0 1 374
box 0 0 120 799
use nand3 g2085
timestamp 1386234893
transform 1 0 5448 0 1 374
box 0 0 120 799
use inv g2104
timestamp 1386238110
transform 1 0 5568 0 1 374
box 0 0 120 799
use inv g2108
timestamp 1386238110
transform 1 0 5688 0 1 374
box 0 0 120 799
use nor2 g2093
timestamp 1386235306
transform 1 0 5808 0 1 374
box 0 0 120 799
use nand2 g2102
timestamp 1386234792
transform 1 0 5928 0 1 374
box 0 0 96 799
use mux2 g2103
timestamp 1386235218
transform 1 0 6024 0 1 374
box 0 0 192 799
use nand2 g2105
timestamp 1386234792
transform 1 0 6216 0 1 374
box 0 0 96 799
use and2 g2107
timestamp 1386234845
transform 1 0 6312 0 1 374
box 0 0 120 799
use nand2 g2109
timestamp 1386234792
transform 1 0 6432 0 1 374
box 0 0 96 799
use and2 g2110
timestamp 1386234845
transform 1 0 6528 0 1 374
box 0 0 120 799
use inv g2112
timestamp 1386238110
transform 1 0 6648 0 1 374
box 0 0 120 799
use nor2 g2106
timestamp 1386235306
transform 1 0 6768 0 1 374
box 0 0 120 799
use nand2 g2111
timestamp 1386234792
transform 1 0 6888 0 1 374
box 0 0 96 799
use nand2 g2113
timestamp 1386234792
transform 1 0 6984 0 1 374
box 0 0 96 799
use and2 g2114
timestamp 1386234845
transform 1 0 7080 0 1 374
box 0 0 120 799
use inv g2116
timestamp 1386238110
transform 1 0 7200 0 1 374
box 0 0 120 799
use inv g2117
timestamp 1386238110
transform 1 0 7320 0 1 374
box 0 0 120 799
use inv g2118
timestamp 1386238110
transform 1 0 7440 0 1 374
box 0 0 120 799
use inv g2115
timestamp 1386238110
transform 1 0 7560 0 1 374
box 0 0 120 799
use inv g2119
timestamp 1386238110
transform 1 0 7680 0 1 374
box 0 0 120 799
<< labels >>
rlabel metal2 0 1959 12 1959 5 OpCode[4]
rlabel metal2 120 1959 132 1959 5 OpCode[3]
rlabel metal2 240 1959 252 1959 5 OpCode[2]
rlabel metal2 360 1959 372 1959 5 OpCode[1]
rlabel metal2 480 1959 492 1959 5 OpCode[0]
rlabel metal2 6120 1959 6132 1959 5 imm4[3]
rlabel metal2 6336 1959 6348 1959 5 imm4[2]
rlabel metal2 6456 1959 6468 1959 5 imm4[1]
rlabel metal2 6576 1959 6588 1959 5 imm4[0]
rlabel metal2 600 -488 612 -488 1 LastCIn
rlabel metal2 624 -488 636 -488 1 COut
rlabel metal2 696 -488 708 -488 1 N_slice
rlabel metal2 912 -488 924 -488 1 nZ
rlabel metal2 3264 -488 3276 -488 1 ASign
rlabel metal2 0 -488 12 -488 1 ZeroA
rlabel metal2 264 -488 276 -488 1 SUB
rlabel metal2 1056 -488 1068 -488 1 FAOut
rlabel metal2 1392 -488 1404 -488 1 AND
rlabel metal2 1752 -488 1764 -488 1 OR
rlabel metal2 2496 -488 2508 -488 1 NOT
rlabel metal2 2808 -488 2820 -488 1 NAND
rlabel metal2 5280 -488 5292 -488 1 Sh8
rlabel metal2 5664 -488 5676 -488 1 ShInBit
rlabel metal2 432 -488 444 -488 1 CIn_slice
rlabel metal2 2160 -488 2172 -488 1 XOR
rlabel metal2 3144 -488 3156 -488 1 NOR
rlabel metal2 3312 -488 3324 -488 1 ShB
rlabel metal2 3480 -488 3492 -488 1 ShL
rlabel metal2 5305 -488 5317 -488 1 ShR
rlabel metal2 5928 -488 5940 -488 1 Sh4
rlabel metal2 6384 -488 6396 -488 1 Sh2
rlabel metal2 6744 -488 6756 -488 1 Sh1
rlabel metal2 7104 -488 7116 -488 1 ShOut
rlabel metal2 7272 -488 7284 -488 1 LLI
rlabel metal2 7512 -488 7524 -488 1 OutEn_slice
<< end >>
