magic
tech c035u
timestamp 1393710283
<< metal1 >>
rect 2677 1309 3719 1319
rect 2557 1287 3623 1297
rect 2317 1265 3431 1275
rect 2077 1244 3239 1254
rect 1957 1222 3143 1232
rect 709 1200 1103 1210
rect 2797 1200 3047 1210
rect 3061 1200 3815 1210
rect 829 1178 1079 1188
rect 1165 1178 1320 1188
rect 1381 1178 1439 1188
rect 2437 1178 2951 1188
rect 2965 1178 3527 1188
rect 925 1156 960 1166
rect 1045 1156 1199 1166
rect 1285 1156 1415 1166
rect 2197 1156 2855 1166
rect 2869 1156 3335 1166
rect 3565 1156 5255 1166
rect 517 1134 671 1144
rect 685 1134 863 1144
rect 877 1134 2039 1144
rect 2053 1134 2279 1144
rect 2293 1134 2519 1144
rect 2533 1134 2759 1144
rect 2773 1134 3935 1144
rect 3949 1134 4271 1144
rect 397 1112 1343 1122
rect 1357 1112 2135 1122
rect 2149 1112 2255 1122
rect 2269 1112 2615 1122
rect 2629 1112 2735 1122
rect 2749 1112 3911 1122
rect 3925 1112 4151 1122
rect 4165 1112 4247 1122
rect 4261 1112 4775 1122
rect 4789 1112 5759 1122
rect 277 1090 647 1100
rect 661 1090 983 1100
rect 997 1090 1559 1100
rect 1573 1090 2351 1100
rect 2365 1090 2471 1100
rect 2485 1090 2591 1100
rect 2605 1090 2711 1100
rect 2725 1090 5735 1100
rect 5965 1090 6023 1100
rect 157 1068 791 1078
rect 805 1068 1223 1078
rect 1237 1068 1799 1078
rect 1813 1068 3887 1078
rect 3973 1068 4006 1078
rect 4333 1068 4391 1078
rect 4717 1068 4895 1078
rect 4957 1068 4991 1078
rect 5101 1068 5135 1078
rect 5149 1068 5351 1078
rect 5365 1068 5471 1078
rect 5485 1068 5591 1078
rect 5821 1068 5999 1078
rect 6277 1068 6575 1078
rect 37 1046 1535 1056
rect 1549 1046 1679 1056
rect 1693 1046 1775 1056
rect 1789 1046 4031 1056
rect 4213 1046 4367 1056
rect 4453 1046 4487 1056
rect 4837 1046 4871 1056
rect 4885 1046 6047 1056
rect 6109 1046 6143 1056
rect 6349 1046 6383 1056
rect 6613 1046 6887 1056
rect 7032 963 7042 988
rect 7032 318 7042 343
rect 85 227 623 237
rect 637 227 1247 237
rect 1261 227 4511 237
rect 4525 227 5015 237
rect 5029 227 6167 237
rect 6421 229 6767 239
rect 205 205 1703 215
rect 1717 205 4127 215
rect 4141 205 5039 215
rect 5053 205 5711 215
rect 5725 205 5855 215
rect 325 183 767 193
rect 781 183 887 193
rect 901 183 1583 193
rect 1597 183 1871 193
rect 1885 183 1991 193
rect 2005 183 2111 193
rect 2125 183 2231 193
rect 2245 183 4535 193
rect 4549 183 4631 193
rect 4645 183 4751 193
rect 4765 183 5879 193
rect 445 161 1895 171
rect 1909 161 2015 171
rect 2029 161 2375 171
rect 2389 161 2495 171
rect 3133 161 3215 171
rect 3229 161 3311 171
rect 3325 161 3407 171
rect 3421 161 3503 171
rect 3517 161 3599 171
rect 3613 161 3695 171
rect 3709 161 3791 171
rect 5189 161 5223 171
rect 565 139 743 149
rect 757 139 1919 149
rect 1933 139 2159 149
rect 2173 139 2399 149
rect 2413 139 2639 149
rect 2653 139 4655 149
rect 4669 139 5903 149
rect 1837 116 2831 126
rect 2845 116 2927 126
rect 2941 116 3023 126
rect 3085 117 4202 127
rect 1741 94 3119 104
rect 3321 95 3455 105
rect 3565 95 4146 105
rect 1576 72 2879 82
rect 3661 73 6349 83
rect 2989 51 4656 61
rect 1501 29 6407 39
rect 1645 7 6287 17
<< m2contact >>
rect 2663 1307 2677 1321
rect 3719 1307 3733 1321
rect 2543 1285 2557 1299
rect 3623 1285 3637 1299
rect 2303 1264 2317 1278
rect 3431 1263 3445 1277
rect 2063 1242 2077 1256
rect 3239 1241 3253 1255
rect 1943 1220 1957 1234
rect 3143 1220 3157 1234
rect 695 1198 709 1212
rect 1103 1198 1117 1212
rect 2783 1198 2797 1212
rect 3047 1198 3061 1212
rect 3815 1198 3829 1212
rect 815 1176 829 1190
rect 1079 1176 1093 1190
rect 1151 1176 1165 1190
rect 1320 1176 1334 1190
rect 1367 1176 1381 1190
rect 1439 1176 1453 1190
rect 2423 1176 2437 1190
rect 2951 1176 2965 1190
rect 3527 1176 3541 1190
rect 911 1154 925 1168
rect 960 1154 974 1168
rect 1031 1154 1045 1168
rect 1199 1154 1213 1168
rect 1271 1154 1285 1168
rect 1415 1154 1429 1168
rect 2183 1154 2197 1168
rect 2855 1154 2869 1168
rect 3335 1154 3349 1168
rect 3551 1154 3565 1168
rect 5255 1154 5269 1168
rect 503 1132 517 1146
rect 671 1132 685 1146
rect 863 1132 877 1146
rect 2039 1132 2053 1146
rect 2279 1132 2293 1146
rect 2519 1132 2533 1146
rect 2759 1132 2773 1146
rect 3935 1132 3949 1146
rect 4271 1132 4285 1146
rect 383 1110 397 1124
rect 1343 1110 1357 1124
rect 2135 1110 2149 1124
rect 2255 1110 2269 1124
rect 2615 1110 2629 1124
rect 2735 1110 2749 1124
rect 3911 1110 3925 1124
rect 4151 1110 4165 1124
rect 4247 1110 4261 1124
rect 4775 1110 4789 1124
rect 5759 1110 5773 1124
rect 263 1088 277 1102
rect 647 1088 661 1102
rect 983 1088 997 1102
rect 1559 1088 1573 1102
rect 2351 1088 2365 1102
rect 2471 1088 2485 1102
rect 2591 1088 2605 1102
rect 2711 1088 2725 1102
rect 5735 1088 5749 1102
rect 5951 1088 5965 1102
rect 6023 1088 6037 1102
rect 143 1066 157 1080
rect 791 1066 805 1080
rect 1223 1066 1237 1080
rect 1799 1066 1813 1080
rect 3887 1066 3901 1080
rect 3959 1066 3973 1080
rect 4006 1066 4020 1080
rect 4319 1066 4333 1080
rect 4391 1066 4405 1080
rect 4703 1066 4717 1080
rect 4895 1066 4909 1080
rect 4943 1066 4957 1080
rect 4991 1066 5005 1080
rect 5087 1066 5101 1080
rect 5135 1066 5149 1080
rect 5351 1066 5365 1080
rect 5471 1066 5485 1080
rect 5591 1066 5605 1080
rect 5807 1066 5821 1080
rect 5999 1066 6013 1080
rect 6263 1066 6277 1080
rect 6575 1066 6589 1080
rect 23 1044 37 1058
rect 1535 1044 1549 1058
rect 1679 1044 1693 1058
rect 1775 1044 1789 1058
rect 4031 1044 4045 1058
rect 4199 1044 4213 1058
rect 4367 1044 4381 1058
rect 4439 1044 4453 1058
rect 4487 1044 4501 1058
rect 4823 1044 4837 1058
rect 4871 1044 4885 1058
rect 6047 1044 6061 1058
rect 6095 1044 6109 1058
rect 6143 1044 6157 1058
rect 6335 1044 6349 1058
rect 6383 1044 6397 1058
rect 6599 1044 6613 1058
rect 6887 1044 6901 1058
rect 71 225 85 239
rect 623 225 637 239
rect 1247 225 1261 239
rect 4511 225 4525 239
rect 5015 225 5029 239
rect 6167 225 6181 239
rect 6407 227 6421 241
rect 6767 227 6781 241
rect 191 203 205 217
rect 1703 203 1717 217
rect 4127 203 4141 217
rect 5039 203 5053 217
rect 5711 203 5725 217
rect 5855 203 5869 217
rect 311 181 325 195
rect 767 181 781 195
rect 887 181 901 195
rect 1583 181 1597 195
rect 1871 181 1885 195
rect 1991 181 2005 195
rect 2111 181 2125 195
rect 2231 181 2245 195
rect 4535 181 4549 195
rect 4631 181 4645 195
rect 4751 181 4765 195
rect 5879 181 5893 195
rect 431 159 445 173
rect 1895 159 1909 173
rect 2015 159 2029 173
rect 2375 159 2389 173
rect 2495 159 2509 173
rect 3119 159 3133 173
rect 3215 159 3229 173
rect 3311 159 3325 173
rect 3407 159 3421 173
rect 3503 159 3517 173
rect 3599 159 3613 173
rect 3695 159 3709 173
rect 3791 159 3805 173
rect 5175 159 5189 173
rect 5223 159 5237 173
rect 551 137 565 151
rect 743 137 757 151
rect 1919 137 1933 151
rect 2159 137 2173 151
rect 2399 137 2413 151
rect 2639 137 2653 151
rect 4655 137 4669 151
rect 5903 136 5917 150
rect 1823 114 1837 128
rect 2831 114 2845 128
rect 2927 114 2941 128
rect 3023 114 3037 128
rect 3071 115 3085 129
rect 4202 115 4216 129
rect 1727 92 1741 106
rect 3119 92 3133 106
rect 3307 93 3321 107
rect 3455 93 3469 107
rect 3551 93 3565 107
rect 4146 93 4160 107
rect 1562 70 1576 84
rect 2879 70 2893 84
rect 3647 71 3661 85
rect 6349 71 6363 85
rect 2975 49 2989 63
rect 4656 49 4670 63
rect 1487 27 1501 41
rect 6407 27 6421 41
rect 1631 5 1645 19
rect 6287 5 6301 19
<< metal2 >>
rect 24 1058 36 1326
rect 144 1080 156 1326
rect 264 1102 276 1326
rect 384 1124 396 1326
rect 504 1146 516 1326
rect 24 1041 36 1044
rect 144 1041 156 1066
rect 264 1041 276 1088
rect 384 1041 396 1110
rect 504 1041 516 1132
rect 648 1041 660 1088
rect 672 1041 684 1132
rect 696 1041 708 1198
rect 792 1041 804 1066
rect 816 1041 828 1176
rect 864 1041 876 1132
rect 912 1041 924 1154
rect 960 1041 972 1154
rect 984 1041 996 1088
rect 1032 1041 1044 1154
rect 1080 1041 1092 1176
rect 1104 1041 1116 1198
rect 1152 1041 1164 1176
rect 1200 1041 1212 1154
rect 1224 1041 1236 1066
rect 1272 1041 1284 1154
rect 1320 1041 1332 1176
rect 1344 1041 1356 1110
rect 1368 1041 1380 1176
rect 1416 1041 1428 1154
rect 1440 1041 1452 1176
rect 1536 1041 1548 1044
rect 1560 1041 1572 1088
rect 1680 1041 1692 1044
rect 1776 1041 1788 1044
rect 1800 1041 1812 1066
rect 1944 1041 1956 1220
rect 2040 1041 2052 1132
rect 2064 1041 2076 1242
rect 2136 1041 2148 1110
rect 2184 1041 2196 1154
rect 2256 1041 2268 1110
rect 2280 1041 2292 1132
rect 2304 1041 2316 1264
rect 2352 1041 2364 1088
rect 2424 1041 2436 1176
rect 2472 1041 2484 1088
rect 2520 1041 2532 1132
rect 2544 1041 2556 1285
rect 2592 1041 2604 1088
rect 2616 1041 2628 1110
rect 2664 1041 2676 1307
rect 2712 1041 2724 1088
rect 2736 1041 2748 1110
rect 2760 1041 2772 1132
rect 2784 1041 2796 1198
rect 2856 1041 2868 1154
rect 2952 1041 2964 1176
rect 3048 1041 3060 1198
rect 3144 1041 3156 1220
rect 3240 1041 3252 1241
rect 3336 1041 3348 1154
rect 3432 1041 3444 1263
rect 3528 1041 3540 1176
rect 3552 1041 3564 1154
rect 3624 1041 3636 1285
rect 3720 1041 3732 1307
rect 3816 1041 3828 1198
rect 3888 1041 3900 1066
rect 3912 1041 3924 1110
rect 3936 1041 3948 1132
rect 3960 1041 3972 1066
rect 4008 1041 4020 1066
rect 4032 1041 4044 1044
rect 4152 1041 4164 1110
rect 4200 1041 4212 1044
rect 4248 1041 4260 1110
rect 4272 1041 4284 1132
rect 4320 1041 4332 1066
rect 4368 1041 4380 1044
rect 4392 1041 4404 1066
rect 4440 1041 4452 1044
rect 4488 1041 4500 1044
rect 4704 1041 4716 1066
rect 4776 1041 4788 1110
rect 4824 1041 4836 1044
rect 4872 1041 4884 1044
rect 4896 1041 4908 1066
rect 4944 1041 4956 1066
rect 4992 1041 5004 1066
rect 5088 1041 5100 1066
rect 5136 1041 5148 1066
rect 5160 1041 5172 1326
rect 5256 1041 5268 1154
rect 5352 1041 5364 1066
rect 5376 1041 5388 1326
rect 5472 1041 5484 1066
rect 5496 1041 5508 1326
rect 5592 1041 5604 1066
rect 5616 1041 5628 1326
rect 5736 1041 5748 1088
rect 5760 1041 5772 1110
rect 5808 1041 5820 1066
rect 5952 1041 5964 1088
rect 6000 1041 6012 1066
rect 6024 1041 6036 1088
rect 6264 1080 6276 1326
rect 6048 1041 6060 1044
rect 6096 1041 6108 1044
rect 6144 1041 6156 1044
rect 6264 1041 6276 1066
rect 6336 1041 6348 1044
rect 6384 1041 6396 1044
rect 6576 1041 6588 1066
rect 6600 1041 6612 1044
rect 6696 1041 6708 1326
rect 6792 1041 6804 1326
rect 6888 1041 6900 1044
rect 6960 1041 6972 1326
rect 7008 1041 7020 1326
rect 72 239 84 242
rect 192 217 204 242
rect 312 195 324 242
rect 432 173 444 242
rect 552 151 564 242
rect 624 239 636 242
rect 744 151 756 242
rect 768 195 780 242
rect 888 195 900 242
rect 1248 239 1260 242
rect 1488 41 1500 242
rect 1584 195 1596 242
rect 1488 0 1500 27
rect 1563 0 1575 70
rect 1632 19 1644 242
rect 1704 217 1716 242
rect 1728 106 1740 242
rect 1824 128 1836 242
rect 1872 195 1884 242
rect 1896 173 1908 242
rect 1920 151 1932 242
rect 1992 195 2004 242
rect 2016 173 2028 242
rect 2112 195 2124 242
rect 2160 151 2172 242
rect 2232 195 2244 242
rect 2376 173 2388 242
rect 2400 151 2412 242
rect 2496 173 2508 242
rect 2640 151 2652 242
rect 2832 128 2844 242
rect 2880 84 2892 242
rect 2928 128 2940 242
rect 2976 63 2988 242
rect 3024 128 3036 242
rect 3072 129 3084 242
rect 3120 173 3132 242
rect 3120 106 3132 159
rect 1632 0 1644 5
rect 3168 0 3180 242
rect 3216 173 3228 242
rect 3264 0 3276 242
rect 3312 173 3324 242
rect 3308 0 3320 93
rect 3360 0 3372 242
rect 3408 173 3420 242
rect 3456 107 3468 242
rect 3504 173 3516 242
rect 3552 107 3564 242
rect 3600 173 3612 242
rect 3648 85 3660 242
rect 3696 173 3708 242
rect 3744 0 3756 242
rect 3792 173 3804 242
rect 3840 0 3852 242
rect 4080 0 4092 242
rect 4128 217 4140 242
rect 4512 239 4524 242
rect 4536 195 4548 242
rect 4147 0 4159 93
rect 4203 0 4215 115
rect 4584 0 4596 242
rect 4632 195 4644 242
rect 4656 151 4668 242
rect 4752 195 4764 242
rect 5016 239 5028 242
rect 5040 217 5052 242
rect 5176 173 5188 242
rect 5224 173 5236 242
rect 4657 0 4669 49
rect 5304 0 5316 242
rect 5424 0 5436 242
rect 5544 0 5556 242
rect 5664 0 5676 242
rect 5712 217 5724 242
rect 5856 217 5868 242
rect 5880 195 5892 242
rect 5904 150 5916 242
rect 6168 239 6180 242
rect 6216 0 6228 242
rect 6288 19 6300 242
rect 6408 241 6420 242
rect 6350 0 6362 71
rect 6408 41 6420 227
rect 6504 0 6516 242
rect 6768 241 6780 242
rect 6768 225 6780 227
rect 6792 0 6804 242
rect 6960 0 6972 242
rect 7008 0 7020 242
use inv inv_0
timestamp 1386238110
transform 1 0 0 0 1 242
box 0 0 120 799
use inv inv_1
timestamp 1386238110
transform 1 0 120 0 1 242
box 0 0 120 799
use inv inv_2
timestamp 1386238110
transform 1 0 240 0 1 242
box 0 0 120 799
use inv inv_3
timestamp 1386238110
transform 1 0 360 0 1 242
box 0 0 120 799
use inv inv_4
timestamp 1386238110
transform 1 0 480 0 1 242
box 0 0 120 799
use nand3 nand3_0
timestamp 1386234893
transform 1 0 600 0 1 242
box 0 0 120 799
use nand3 nand3_1
timestamp 1386234893
transform 1 0 720 0 1 242
box 0 0 120 799
use nand2 nand2_0
timestamp 1386234792
transform 1 0 840 0 1 242
box 0 0 96 799
use nor2 nor2_0
timestamp 1386235306
transform 1 0 936 0 1 242
box 0 0 120 799
use nor2 nor2_1
timestamp 1386235306
transform 1 0 1056 0 1 242
box 0 0 120 799
use nand3 nand3_2
timestamp 1386234893
transform 1 0 1176 0 1 242
box 0 0 120 799
use nand2 nand2_1
timestamp 1386234792
transform 1 0 1296 0 1 242
box 0 0 96 799
use nor2 nor2_2
timestamp 1386235306
transform 1 0 1392 0 1 242
box 0 0 120 799
use nor3 nor3_0
timestamp 1386235396
transform 1 0 1512 0 1 242
box 0 0 144 799
use nand2 nand2_2
timestamp 1386234792
transform 1 0 1656 0 1 242
box 0 0 96 799
use nand2 nand2_3
timestamp 1386234792
transform 1 0 1752 0 1 242
box 0 0 96 799
use nand3 nand3_4
timestamp 1386234893
transform 1 0 1848 0 1 242
box 0 0 120 799
use nand3 nand3_5
timestamp 1386234893
transform 1 0 1968 0 1 242
box 0 0 120 799
use nand3 nand3_6
timestamp 1386234893
transform 1 0 2088 0 1 242
box 0 0 120 799
use nand3 nand3_7
timestamp 1386234893
transform 1 0 2208 0 1 242
box 0 0 120 799
use nand3 nand3_8
timestamp 1386234893
transform 1 0 2328 0 1 242
box 0 0 120 799
use nand3 nand3_9
timestamp 1386234893
transform 1 0 2448 0 1 242
box 0 0 120 799
use nand3 nand3_10
timestamp 1386234893
transform 1 0 2568 0 1 242
box 0 0 120 799
use nand3 nand3_11
timestamp 1386234893
transform 1 0 2688 0 1 242
box 0 0 120 799
use nand2 nand2_4
timestamp 1386234792
transform 1 0 2808 0 1 242
box 0 0 96 799
use nand2 nand2_5
timestamp 1386234792
transform 1 0 2904 0 1 242
box 0 0 96 799
use nand2 nand2_6
timestamp 1386234792
transform 1 0 3000 0 1 242
box 0 0 96 799
use nand2 nand2_7
timestamp 1386234792
transform 1 0 3096 0 1 242
box 0 0 96 799
use nand2 nand2_8
timestamp 1386234792
transform 1 0 3192 0 1 242
box 0 0 96 799
use nand2 nand2_9
timestamp 1386234792
transform 1 0 3288 0 1 242
box 0 0 96 799
use nand2 nand2_10
timestamp 1386234792
transform 1 0 3384 0 1 242
box 0 0 96 799
use nand2 nand2_11
timestamp 1386234792
transform 1 0 3480 0 1 242
box 0 0 96 799
use nand2 nand2_12
timestamp 1386234792
transform 1 0 3576 0 1 242
box 0 0 96 799
use nand2 nand2_13
timestamp 1386234792
transform 1 0 3672 0 1 242
box 0 0 96 799
use nand2 nand2_14
timestamp 1386234792
transform 1 0 3768 0 1 242
box 0 0 96 799
use nand3 nand3_3
timestamp 1386234893
transform 1 0 3864 0 1 242
box 0 0 120 799
use nor2 nor2_3
timestamp 1386235306
transform 1 0 3984 0 1 242
box 0 0 120 799
use nor2 nor2_4
timestamp 1386235306
transform 1 0 4104 0 1 242
box 0 0 120 799
use nor2 nor2_5
timestamp 1386235306
transform 1 0 4224 0 1 242
box 0 0 120 799
use nor2 nor2_6
timestamp 1386235306
transform 1 0 4344 0 1 242
box 0 0 120 799
use nor3 nor3_1
timestamp 1386235396
transform 1 0 4464 0 1 242
box 0 0 144 799
use nor2 nor2_7
timestamp 1386235306
transform 1 0 4608 0 1 242
box 0 0 120 799
use nor2 nor2_8
timestamp 1386235306
transform 1 0 4728 0 1 242
box 0 0 120 799
use nor2 nor2_9
timestamp 1386235306
transform 1 0 4848 0 1 242
box 0 0 120 799
use nor3 nor3_2
timestamp 1386235396
transform 1 0 4968 0 1 242
box 0 0 144 799
use nand2 nand2_15
timestamp 1386234792
transform 1 0 5112 0 1 242
box 0 0 96 799
use nor2 nor2_10
timestamp 1386235306
transform 1 0 5208 0 1 242
box 0 0 120 799
use and2 and2_0
timestamp 1386234845
transform 1 0 5328 0 1 242
box 0 0 120 799
use and2 and2_1
timestamp 1386234845
transform 1 0 5448 0 1 242
box 0 0 120 799
use and2 and2_2
timestamp 1386234845
transform 1 0 5568 0 1 242
box 0 0 120 799
use nor3 nor3_3
timestamp 1386235396
transform 1 0 5688 0 1 242
box 0 0 144 799
use nor3 nor3_4
timestamp 1386235396
transform 1 0 5832 0 1 242
box 0 0 144 799
use nor3 nor3_5
timestamp 1386235396
transform 1 0 5976 0 1 242
box 0 0 144 799
use nor2 nor2_11
timestamp 1386235306
transform 1 0 6120 0 1 242
box 0 0 120 799
use and2 and2_3
timestamp 1386234845
transform 1 0 6240 0 1 242
box 0 0 120 799
use xor2 xor2_0
timestamp 1386237344
transform 1 0 6360 0 1 242
box 0 0 192 799
use xor2 xor2_1
timestamp 1386237344
transform 1 0 6552 0 1 242
box 0 0 192 799
use xor2 xor2_2
timestamp 1386237344
transform 1 0 6744 0 1 242
box 0 0 192 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 6936 0 1 242
box 0 0 48 799
use rowcrosser rowcrosser_1
timestamp 1386086759
transform 1 0 6984 0 1 242
box 0 0 48 799
<< labels >>
rlabel metal1 336 189 336 189 1 nC
rlabel metal1 579 142 579 142 1 nE
rlabel metal2 5093 1043 5093 1043 1 N
rlabel metal1 104 231 104 231 1 nA
rlabel metal1 210 209 210 209 1 nB
rlabel metal1 459 164 459 164 1 nD
rlabel metal2 24 1326 36 1326 5 OpCode[4]
rlabel metal2 144 1326 156 1326 5 OpCode[3]
rlabel metal2 264 1326 276 1326 5 OpCode[2]
rlabel metal2 384 1326 396 1326 5 OpCode[1]
rlabel metal2 504 1326 516 1326 5 OpCode[0]
rlabel metal2 5160 1326 5172 1326 5 imm4[3]
rlabel metal2 5376 1326 5388 1326 5 imm4[2]
rlabel metal2 5496 1326 5508 1326 5 imm4[1]
rlabel metal2 5616 1326 5628 1326 5 imm4[0]
rlabel metal2 6264 1326 6276 1326 5 Cin
rlabel metal2 6696 1326 6708 1326 5 V
rlabel metal2 6792 1326 6804 1326 5 C
rlabel metal2 6960 1326 6972 1326 5 N
rlabel metal2 7008 1326 7020 1326 5 Z
rlabel metal2 7008 0 7020 0 1 Z
rlabel metal2 6960 0 6972 0 1 N
rlabel metal2 6792 0 6804 0 1 C
rlabel metal2 6504 0 6516 0 1 Cin_slice
rlabel metal2 1488 0 1500 0 1 SUB
rlabel metal2 1563 0 1575 0 1 ZeroA
rlabel metal2 1632 0 1644 0 1 UseC
rlabel metal2 3168 0 3180 0 1 AND
rlabel metal2 3264 0 3276 0 1 OR
rlabel metal2 3308 0 3320 0 1 XOR
rlabel metal2 3360 0 3372 0 1 NOT
rlabel metal2 3744 0 3756 0 1 NAND
rlabel metal2 3840 0 3852 0 1 NOR
rlabel metal2 4080 0 4092 0 1 FAOut
rlabel metal2 4147 0 4159 0 1 ShB
rlabel metal2 4203 0 4215 0 1 ShL
rlabel metal2 4584 0 4596 0 1 ShR
rlabel metal2 4657 0 4669 0 1 ShSign
rlabel metal2 5304 0 5316 0 1 Sh8
rlabel metal2 5424 0 5436 0 1 Sh4
rlabel metal2 5544 0 5556 0 1 Sh2
rlabel metal2 5664 0 5676 0 1 Sh1
rlabel metal2 6216 0 6228 0 1 ShOut
rlabel metal2 6350 0 6362 0 1 LLI
rlabel metal1 7042 318 7042 343 7 GND!
rlabel metal1 7042 963 7042 988 7 Vdd!
<< end >>
